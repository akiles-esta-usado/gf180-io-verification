* NGSPICE file created from gf180mcu_fd_io__asig_5p0_pex.ext - technology: gf180mcuD

.subckt gf180mcu_fd_io__asig_5p0_pex VSS VDD DVSS DVDD ASIG5V
X0 DVDD.t1 DVSS.t36 cap_nmos_06v0 c_width=15u c_length=15u
X1 DVDD.t2 DVSS.t35 cap_nmos_06v0 c_width=15u c_length=15u
X2 DVDD.t3 DVSS.t34 cap_nmos_06v0 c_width=15u c_length=15u
X3 DVDD.t4 DVSS.t33 cap_nmos_06v0 c_width=15u c_length=15u
X4 DVDD.t5 DVSS.t32 cap_nmos_06v0 c_width=15u c_length=15u
D0 DVSS.t3 DVDD.t6 diode_nd2ps_06v0 pj=82u area=40p
X5 DVDD.t7 DVSS.t31 cap_nmos_06v0 c_width=15u c_length=15u
X6 DVDD.t8 DVSS.t30 cap_nmos_06v0 c_width=15u c_length=15u
X7 DVDD.t9 DVSS.t29 cap_nmos_06v0 c_width=15u c_length=15u
X8 DVDD.t10 DVSS.t28 cap_nmos_06v0 c_width=15u c_length=15u
X9 DVDD.t11 DVSS.t27 cap_nmos_06v0 c_width=15u c_length=15u
X10 DVDD.t12 DVSS.t26 cap_nmos_06v0 c_width=15u c_length=15u
X11 DVDD.t13 DVSS.t25 cap_nmos_06v0 c_width=15u c_length=15u
X12 DVDD.t14 DVSS.t24 cap_nmos_06v0 c_width=15u c_length=15u
X13 DVDD.t15 DVSS.t23 cap_nmos_06v0 c_width=15u c_length=15u
X14 DVDD.t16 DVSS.t22 cap_nmos_06v0 c_width=15u c_length=15u
D1 DVSS.t37 ASIG5V.t0 diode_nd2ps_06v0 pj=0.106m area=0.15n
X15 DVDD.t17 DVSS.t21 cap_nmos_06v0 c_width=15u c_length=15u
X16 DVDD.t18 DVSS.t20 cap_nmos_06v0 c_width=15u c_length=15u
X17 DVDD.t19 DVSS.t19 cap_nmos_06v0 c_width=15u c_length=15u
D2 DVSS.t37 ASIG5V.t1 diode_nd2ps_06v0 pj=0.106m area=0.15n
D3 ASIG5V.t2 DVDD.t0 diode_pd2nw_06v0 pj=0.106m area=0.15n
X18 DVDD.t20 DVSS.t18 cap_nmos_06v0 c_width=15u c_length=15u
X19 DVDD.t21 DVSS.t17 cap_nmos_06v0 c_width=15u c_length=15u
D4 ASIG5V.t3 DVDD.t0 diode_pd2nw_06v0 pj=0.106m area=0.15n
D5 DVSS.t37 ASIG5V.t4 diode_nd2ps_06v0 pj=0.106m area=0.15n
X20 DVDD.t22 DVSS.t16 cap_nmos_06v0 c_width=15u c_length=15u
D6 ASIG5V.t5 DVDD.t0 diode_pd2nw_06v0 pj=0.106m area=0.15n
X21 DVDD.t23 DVSS.t15 cap_nmos_06v0 c_width=15u c_length=15u
X22 DVDD.t24 DVSS.t14 cap_nmos_06v0 c_width=15u c_length=15u
D7 DVSS.t3 DVDD.t25 diode_nd2ps_06v0 pj=82u area=40p
X23 DVDD.t26 DVSS.t13 cap_nmos_06v0 c_width=15u c_length=15u
X24 DVDD.t27 DVSS.t12 cap_nmos_06v0 c_width=15u c_length=15u
X25 DVDD.t28 DVSS.t11 cap_nmos_06v0 c_width=15u c_length=15u
X26 DVDD.t29 DVSS.t10 cap_nmos_06v0 c_width=15u c_length=15u
X27 DVDD.t30 DVSS.t9 cap_nmos_06v0 c_width=15u c_length=15u
D8 DVSS.t3 DVDD.t31 diode_nd2ps_06v0 pj=82u area=40p
X28 DVDD.t32 DVSS.t8 cap_nmos_06v0 c_width=15u c_length=15u
D9 DVSS.t37 ASIG5V.t6 diode_nd2ps_06v0 pj=0.106m area=0.15n
X29 DVDD.t33 DVSS.t7 cap_nmos_06v0 c_width=15u c_length=15u
X30 DVDD.t34 DVSS.t6 cap_nmos_06v0 c_width=15u c_length=15u
X31 DVDD.t35 DVSS.t5 cap_nmos_06v0 c_width=15u c_length=15u
X32 DVDD.t36 DVSS.t4 cap_nmos_06v0 c_width=15u c_length=15u
D10 DVSS.t3 DVDD.t37 diode_nd2ps_06v0 pj=82u area=40p
D11 ASIG5V.t7 DVDD.t0 diode_pd2nw_06v0 pj=0.106m area=0.15n
X33 DVDD.t38 DVSS.t2 cap_nmos_06v0 c_width=15u c_length=15u
X34 DVDD.t39 DVSS.t1 cap_nmos_06v0 c_width=15u c_length=15u
X35 DVDD.t40 DVSS.t0 cap_nmos_06v0 c_width=15u c_length=15u
R0 DVDD.n1305 DVDD.n1304 13378
R1 DVDD.n8641 DVDD.n1304 13378
R2 DVDD.n8641 DVDD.n8640 13378
R3 DVDD.n8640 DVDD.n1305 13378
R4 DVDD.n2343 DVDD.n2342 12277
R5 DVDD.n7728 DVDD.n2342 12277
R6 DVDD.n7728 DVDD.n7727 12277
R7 DVDD.n7727 DVDD.n2343 12277
R8 DVDD.n8587 DVDD.t0 893.734
R9 DVDD.n8616 DVDD.t0 893.734
R10 DVDD.n1372 DVDD.n1340 150.477
R11 DVDD.n8588 DVDD.n1372 150.477
R12 DVDD.n8618 DVDD.n1336 150.477
R13 DVDD.n8618 DVDD.n8617 150.477
R14 DVDD.n8590 DVDD.n8589 84.2907
R15 DVDD.n8590 DVDD.n1343 84.2907
R16 DVDD.n8502 DVDD.n1376 84.2907
R17 DVDD.n8502 DVDD.n1342 84.2907
R18 DVDD.n8429 DVDD.n1375 84.2907
R19 DVDD.n8429 DVDD.n1337 84.2907
R20 DVDD.n8587 DVDD.n1374 26.3372
R21 DVDD.n8616 DVDD.n1341 26.3372
R22 DVDD.n1343 DVDD.n1340 12.9878
R23 DVDD.n1376 DVDD.n1371 12.9878
R24 DVDD.n8589 DVDD.n1371 12.9878
R25 DVDD.n8589 DVDD.n8588 12.9878
R26 DVDD.n1339 DVDD.n1337 12.9878
R27 DVDD.n1342 DVDD.n1339 12.9878
R28 DVDD.n8615 DVDD.n1342 12.9878
R29 DVDD.n8615 DVDD.n1343 12.9878
R30 DVDD.n1375 DVDD.n1336 12.9878
R31 DVDD.n8586 DVDD.n1375 12.9878
R32 DVDD.n8586 DVDD.n1376 12.9878
R33 DVDD.n8617 DVDD.n1337 12.9878
R34 DVDD.n5377 DVDD.n4472 4.5005
R35 DVDD.n5377 DVDD.n4470 4.5005
R36 DVDD.n5466 DVDD.n5377 4.5005
R37 DVDD.n5419 DVDD.n4472 4.5005
R38 DVDD.n5466 DVDD.n5419 4.5005
R39 DVDD.n4483 DVDD.n4472 4.5005
R40 DVDD.n5466 DVDD.n4483 4.5005
R41 DVDD.n5422 DVDD.n4472 4.5005
R42 DVDD.n5422 DVDD.n4470 4.5005
R43 DVDD.n5466 DVDD.n5422 4.5005
R44 DVDD.n4482 DVDD.n4471 4.5005
R45 DVDD.n4482 DVDD.n4472 4.5005
R46 DVDD.n4482 DVDD.n4470 4.5005
R47 DVDD.n5466 DVDD.n4482 4.5005
R48 DVDD.n5423 DVDD.n4471 4.5005
R49 DVDD.n5423 DVDD.n4472 4.5005
R50 DVDD.n5423 DVDD.n4470 4.5005
R51 DVDD.n5466 DVDD.n5423 4.5005
R52 DVDD.n4481 DVDD.n4471 4.5005
R53 DVDD.n4481 DVDD.n4472 4.5005
R54 DVDD.n4481 DVDD.n4470 4.5005
R55 DVDD.n5466 DVDD.n4481 4.5005
R56 DVDD.n5424 DVDD.n4471 4.5005
R57 DVDD.n5424 DVDD.n4472 4.5005
R58 DVDD.n5424 DVDD.n4470 4.5005
R59 DVDD.n5466 DVDD.n5424 4.5005
R60 DVDD.n4480 DVDD.n4471 4.5005
R61 DVDD.n4480 DVDD.n4472 4.5005
R62 DVDD.n4480 DVDD.n4470 4.5005
R63 DVDD.n5466 DVDD.n4480 4.5005
R64 DVDD.n5425 DVDD.n4471 4.5005
R65 DVDD.n5425 DVDD.n4472 4.5005
R66 DVDD.n5425 DVDD.n4470 4.5005
R67 DVDD.n5466 DVDD.n5425 4.5005
R68 DVDD.n4479 DVDD.n4471 4.5005
R69 DVDD.n4479 DVDD.n4472 4.5005
R70 DVDD.n4479 DVDD.n4470 4.5005
R71 DVDD.n5466 DVDD.n4479 4.5005
R72 DVDD.n5426 DVDD.n4471 4.5005
R73 DVDD.n5426 DVDD.n4472 4.5005
R74 DVDD.n5426 DVDD.n4470 4.5005
R75 DVDD.n5466 DVDD.n5426 4.5005
R76 DVDD.n4478 DVDD.n4471 4.5005
R77 DVDD.n4478 DVDD.n4472 4.5005
R78 DVDD.n4478 DVDD.n4470 4.5005
R79 DVDD.n5466 DVDD.n4478 4.5005
R80 DVDD.n5427 DVDD.n4471 4.5005
R81 DVDD.n5427 DVDD.n4472 4.5005
R82 DVDD.n5427 DVDD.n4470 4.5005
R83 DVDD.n5466 DVDD.n5427 4.5005
R84 DVDD.n4477 DVDD.n4471 4.5005
R85 DVDD.n4477 DVDD.n4472 4.5005
R86 DVDD.n4477 DVDD.n4470 4.5005
R87 DVDD.n5466 DVDD.n4477 4.5005
R88 DVDD.n5428 DVDD.n4471 4.5005
R89 DVDD.n5428 DVDD.n4472 4.5005
R90 DVDD.n5428 DVDD.n4470 4.5005
R91 DVDD.n5466 DVDD.n5428 4.5005
R92 DVDD.n4476 DVDD.n4471 4.5005
R93 DVDD.n4476 DVDD.n4472 4.5005
R94 DVDD.n4476 DVDD.n4470 4.5005
R95 DVDD.n5466 DVDD.n4476 4.5005
R96 DVDD.n5429 DVDD.n4471 4.5005
R97 DVDD.n5429 DVDD.n4472 4.5005
R98 DVDD.n5429 DVDD.n4470 4.5005
R99 DVDD.n5466 DVDD.n5429 4.5005
R100 DVDD.n4475 DVDD.n4471 4.5005
R101 DVDD.n4475 DVDD.n4472 4.5005
R102 DVDD.n4475 DVDD.n4470 4.5005
R103 DVDD.n5466 DVDD.n4475 4.5005
R104 DVDD.n5430 DVDD.n4471 4.5005
R105 DVDD.n5430 DVDD.n4472 4.5005
R106 DVDD.n5430 DVDD.n4470 4.5005
R107 DVDD.n5466 DVDD.n5430 4.5005
R108 DVDD.n4474 DVDD.n4471 4.5005
R109 DVDD.n4474 DVDD.n4472 4.5005
R110 DVDD.n4474 DVDD.n4470 4.5005
R111 DVDD.n5466 DVDD.n4474 4.5005
R112 DVDD.n5465 DVDD.n4471 4.5005
R113 DVDD.n5465 DVDD.n4472 4.5005
R114 DVDD.n5465 DVDD.n4470 4.5005
R115 DVDD.n5466 DVDD.n5465 4.5005
R116 DVDD.n5467 DVDD.n4471 4.5005
R117 DVDD.n5467 DVDD.n4472 4.5005
R118 DVDD.n5467 DVDD.n4470 4.5005
R119 DVDD.n5467 DVDD.n5466 4.5005
R120 DVDD.n4471 DVDD.n4467 4.5005
R121 DVDD.n4472 DVDD.n4467 4.5005
R122 DVDD.n4470 DVDD.n4467 4.5005
R123 DVDD.n5466 DVDD.n4467 4.5005
R124 DVDD.n5659 DVDD.n4465 4.5005
R125 DVDD.n4465 DVDD.n4459 4.5005
R126 DVDD.n5483 DVDD.n4465 4.5005
R127 DVDD.n5657 DVDD.n4465 4.5005
R128 DVDD.n5659 DVDD.n4464 4.5005
R129 DVDD.n4464 DVDD.n4459 4.5005
R130 DVDD.n5483 DVDD.n4464 4.5005
R131 DVDD.n5657 DVDD.n4464 4.5005
R132 DVDD.n5659 DVDD.n5480 4.5005
R133 DVDD.n5480 DVDD.n4459 4.5005
R134 DVDD.n5483 DVDD.n5480 4.5005
R135 DVDD.n5657 DVDD.n5480 4.5005
R136 DVDD.n5659 DVDD.n4463 4.5005
R137 DVDD.n4463 DVDD.n4459 4.5005
R138 DVDD.n5657 DVDD.n4463 4.5005
R139 DVDD.n5652 DVDD.n4459 4.5005
R140 DVDD.n5657 DVDD.n5652 4.5005
R141 DVDD.n5643 DVDD.n4459 4.5005
R142 DVDD.n5657 DVDD.n5643 4.5005
R143 DVDD.n5654 DVDD.n4459 4.5005
R144 DVDD.n5657 DVDD.n5654 4.5005
R145 DVDD.n5642 DVDD.n4459 4.5005
R146 DVDD.n5657 DVDD.n5642 4.5005
R147 DVDD.n5656 DVDD.n4459 4.5005
R148 DVDD.n5657 DVDD.n5656 4.5005
R149 DVDD.n5641 DVDD.n4459 4.5005
R150 DVDD.n5641 DVDD.n5483 4.5005
R151 DVDD.n5657 DVDD.n5641 4.5005
R152 DVDD.n5659 DVDD.n5658 4.5005
R153 DVDD.n5658 DVDD.n4459 4.5005
R154 DVDD.n5658 DVDD.n5483 4.5005
R155 DVDD.n5658 DVDD.n5657 4.5005
R156 DVDD.n5615 DVDD.n5493 4.5005
R157 DVDD.n5615 DVDD.n5495 4.5005
R158 DVDD.n5615 DVDD.n5492 4.5005
R159 DVDD.n5615 DVDD.n5614 4.5005
R160 DVDD.n5531 DVDD.n5493 4.5005
R161 DVDD.n5531 DVDD.n5495 4.5005
R162 DVDD.n5531 DVDD.n5492 4.5005
R163 DVDD.n5614 DVDD.n5531 4.5005
R164 DVDD.n5507 DVDD.n5493 4.5005
R165 DVDD.n5507 DVDD.n5495 4.5005
R166 DVDD.n5507 DVDD.n5492 4.5005
R167 DVDD.n5614 DVDD.n5507 4.5005
R168 DVDD.n5532 DVDD.n5493 4.5005
R169 DVDD.n5532 DVDD.n5495 4.5005
R170 DVDD.n5532 DVDD.n5492 4.5005
R171 DVDD.n5614 DVDD.n5532 4.5005
R172 DVDD.n5506 DVDD.n5493 4.5005
R173 DVDD.n5506 DVDD.n5495 4.5005
R174 DVDD.n5506 DVDD.n5492 4.5005
R175 DVDD.n5614 DVDD.n5506 4.5005
R176 DVDD.n5533 DVDD.n5493 4.5005
R177 DVDD.n5533 DVDD.n5495 4.5005
R178 DVDD.n5533 DVDD.n5492 4.5005
R179 DVDD.n5614 DVDD.n5533 4.5005
R180 DVDD.n5505 DVDD.n5493 4.5005
R181 DVDD.n5505 DVDD.n5495 4.5005
R182 DVDD.n5505 DVDD.n5492 4.5005
R183 DVDD.n5614 DVDD.n5505 4.5005
R184 DVDD.n5549 DVDD.n5493 4.5005
R185 DVDD.n5549 DVDD.n5495 4.5005
R186 DVDD.n5549 DVDD.n5492 4.5005
R187 DVDD.n5614 DVDD.n5549 4.5005
R188 DVDD.n5504 DVDD.n5493 4.5005
R189 DVDD.n5504 DVDD.n5495 4.5005
R190 DVDD.n5504 DVDD.n5492 4.5005
R191 DVDD.n5614 DVDD.n5504 4.5005
R192 DVDD.n5552 DVDD.n5493 4.5005
R193 DVDD.n5552 DVDD.n5495 4.5005
R194 DVDD.n5614 DVDD.n5552 4.5005
R195 DVDD.n5503 DVDD.n5495 4.5005
R196 DVDD.n5614 DVDD.n5503 4.5005
R197 DVDD.n5555 DVDD.n5495 4.5005
R198 DVDD.n5614 DVDD.n5555 4.5005
R199 DVDD.n5502 DVDD.n5495 4.5005
R200 DVDD.n5614 DVDD.n5502 4.5005
R201 DVDD.n5558 DVDD.n5495 4.5005
R202 DVDD.n5614 DVDD.n5558 4.5005
R203 DVDD.n5501 DVDD.n5495 4.5005
R204 DVDD.n5614 DVDD.n5501 4.5005
R205 DVDD.n5561 DVDD.n5495 4.5005
R206 DVDD.n5561 DVDD.n5492 4.5005
R207 DVDD.n5614 DVDD.n5561 4.5005
R208 DVDD.n5500 DVDD.n5493 4.5005
R209 DVDD.n5500 DVDD.n5495 4.5005
R210 DVDD.n5500 DVDD.n5492 4.5005
R211 DVDD.n5614 DVDD.n5500 4.5005
R212 DVDD.n5562 DVDD.n5493 4.5005
R213 DVDD.n5562 DVDD.n5495 4.5005
R214 DVDD.n5562 DVDD.n5492 4.5005
R215 DVDD.n5614 DVDD.n5562 4.5005
R216 DVDD.n5499 DVDD.n5493 4.5005
R217 DVDD.n5499 DVDD.n5495 4.5005
R218 DVDD.n5499 DVDD.n5492 4.5005
R219 DVDD.n5614 DVDD.n5499 4.5005
R220 DVDD.n5563 DVDD.n5493 4.5005
R221 DVDD.n5563 DVDD.n5495 4.5005
R222 DVDD.n5563 DVDD.n5492 4.5005
R223 DVDD.n5614 DVDD.n5563 4.5005
R224 DVDD.n5498 DVDD.n5493 4.5005
R225 DVDD.n5498 DVDD.n5495 4.5005
R226 DVDD.n5498 DVDD.n5492 4.5005
R227 DVDD.n5614 DVDD.n5498 4.5005
R228 DVDD.n5564 DVDD.n5493 4.5005
R229 DVDD.n5564 DVDD.n5495 4.5005
R230 DVDD.n5564 DVDD.n5492 4.5005
R231 DVDD.n5614 DVDD.n5564 4.5005
R232 DVDD.n5497 DVDD.n5493 4.5005
R233 DVDD.n5497 DVDD.n5495 4.5005
R234 DVDD.n5497 DVDD.n5492 4.5005
R235 DVDD.n5614 DVDD.n5497 4.5005
R236 DVDD.n5613 DVDD.n5493 4.5005
R237 DVDD.n5613 DVDD.n5495 4.5005
R238 DVDD.n5613 DVDD.n5492 4.5005
R239 DVDD.n5614 DVDD.n5613 4.5005
R240 DVDD.n7024 DVDD.n2535 4.5005
R241 DVDD.n7020 DVDD.n2535 4.5005
R242 DVDD.n2535 DVDD.n2522 4.5005
R243 DVDD.n2535 DVDD.n2521 4.5005
R244 DVDD.n7024 DVDD.n2537 4.5005
R245 DVDD.n7020 DVDD.n2537 4.5005
R246 DVDD.n2537 DVDD.n2522 4.5005
R247 DVDD.n2537 DVDD.n2521 4.5005
R248 DVDD.n7024 DVDD.n2534 4.5005
R249 DVDD.n7020 DVDD.n2534 4.5005
R250 DVDD.n2534 DVDD.n2522 4.5005
R251 DVDD.n2534 DVDD.n2521 4.5005
R252 DVDD.n7024 DVDD.n2538 4.5005
R253 DVDD.n7020 DVDD.n2538 4.5005
R254 DVDD.n2538 DVDD.n2522 4.5005
R255 DVDD.n2538 DVDD.n2521 4.5005
R256 DVDD.n7024 DVDD.n2533 4.5005
R257 DVDD.n7020 DVDD.n2533 4.5005
R258 DVDD.n2533 DVDD.n2522 4.5005
R259 DVDD.n2533 DVDD.n2521 4.5005
R260 DVDD.n7024 DVDD.n2539 4.5005
R261 DVDD.n7020 DVDD.n2539 4.5005
R262 DVDD.n2539 DVDD.n2522 4.5005
R263 DVDD.n2539 DVDD.n2521 4.5005
R264 DVDD.n7024 DVDD.n2532 4.5005
R265 DVDD.n7020 DVDD.n2532 4.5005
R266 DVDD.n2532 DVDD.n2522 4.5005
R267 DVDD.n2532 DVDD.n2521 4.5005
R268 DVDD.n7024 DVDD.n2540 4.5005
R269 DVDD.n7020 DVDD.n2540 4.5005
R270 DVDD.n2540 DVDD.n2522 4.5005
R271 DVDD.n2540 DVDD.n2521 4.5005
R272 DVDD.n7024 DVDD.n2531 4.5005
R273 DVDD.n7020 DVDD.n2531 4.5005
R274 DVDD.n2531 DVDD.n2522 4.5005
R275 DVDD.n2531 DVDD.n2521 4.5005
R276 DVDD.n7024 DVDD.n2541 4.5005
R277 DVDD.n7020 DVDD.n2541 4.5005
R278 DVDD.n2541 DVDD.n2522 4.5005
R279 DVDD.n2541 DVDD.n2521 4.5005
R280 DVDD.n7024 DVDD.n2530 4.5005
R281 DVDD.n7020 DVDD.n2530 4.5005
R282 DVDD.n2530 DVDD.n2522 4.5005
R283 DVDD.n2530 DVDD.n2521 4.5005
R284 DVDD.n7024 DVDD.n2542 4.5005
R285 DVDD.n7020 DVDD.n2542 4.5005
R286 DVDD.n2542 DVDD.n2522 4.5005
R287 DVDD.n2542 DVDD.n2521 4.5005
R288 DVDD.n7024 DVDD.n2529 4.5005
R289 DVDD.n7020 DVDD.n2529 4.5005
R290 DVDD.n2529 DVDD.n2522 4.5005
R291 DVDD.n2529 DVDD.n2521 4.5005
R292 DVDD.n7024 DVDD.n2543 4.5005
R293 DVDD.n7020 DVDD.n2543 4.5005
R294 DVDD.n2543 DVDD.n2522 4.5005
R295 DVDD.n2543 DVDD.n2521 4.5005
R296 DVDD.n7024 DVDD.n2528 4.5005
R297 DVDD.n7020 DVDD.n2528 4.5005
R298 DVDD.n2528 DVDD.n2522 4.5005
R299 DVDD.n2528 DVDD.n2521 4.5005
R300 DVDD.n7024 DVDD.n2545 4.5005
R301 DVDD.n7020 DVDD.n2545 4.5005
R302 DVDD.n2545 DVDD.n2521 4.5005
R303 DVDD.n2527 DVDD.n2521 4.5005
R304 DVDD.n7024 DVDD.n2527 4.5005
R305 DVDD.n2547 DVDD.n2522 4.5005
R306 DVDD.n7024 DVDD.n2547 4.5005
R307 DVDD.n2526 DVDD.n2522 4.5005
R308 DVDD.n7024 DVDD.n2526 4.5005
R309 DVDD.n2549 DVDD.n2522 4.5005
R310 DVDD.n7024 DVDD.n2549 4.5005
R311 DVDD.n2525 DVDD.n2522 4.5005
R312 DVDD.n7024 DVDD.n2525 4.5005
R313 DVDD.n7023 DVDD.n2522 4.5005
R314 DVDD.n7024 DVDD.n7023 4.5005
R315 DVDD.n2524 DVDD.n2522 4.5005
R316 DVDD.n7024 DVDD.n2524 4.5005
R317 DVDD.n7025 DVDD.n2521 4.5005
R318 DVDD.n7025 DVDD.n2522 4.5005
R319 DVDD.n7025 DVDD.n7024 4.5005
R320 DVDD.n7550 DVDD.n7026 4.5005
R321 DVDD.n7026 DVDD.n2508 4.5005
R322 DVDD.n7548 DVDD.n7026 4.5005
R323 DVDD.n7524 DVDD.n2508 4.5005
R324 DVDD.n7548 DVDD.n7524 4.5005
R325 DVDD.n7521 DVDD.n2508 4.5005
R326 DVDD.n7548 DVDD.n7521 4.5005
R327 DVDD.n7525 DVDD.n2508 4.5005
R328 DVDD.n7548 DVDD.n7525 4.5005
R329 DVDD.n7520 DVDD.n2508 4.5005
R330 DVDD.n7548 DVDD.n7520 4.5005
R331 DVDD.n7526 DVDD.n2508 4.5005
R332 DVDD.n7548 DVDD.n7526 4.5005
R333 DVDD.n7519 DVDD.n2508 4.5005
R334 DVDD.n7548 DVDD.n7519 4.5005
R335 DVDD.n7527 DVDD.n2508 4.5005
R336 DVDD.n7548 DVDD.n7527 4.5005
R337 DVDD.n7518 DVDD.n2508 4.5005
R338 DVDD.n7548 DVDD.n7518 4.5005
R339 DVDD.n7528 DVDD.n2508 4.5005
R340 DVDD.n7548 DVDD.n7528 4.5005
R341 DVDD.n7517 DVDD.n2508 4.5005
R342 DVDD.n7548 DVDD.n7517 4.5005
R343 DVDD.n7529 DVDD.n2508 4.5005
R344 DVDD.n7548 DVDD.n7529 4.5005
R345 DVDD.n7516 DVDD.n2508 4.5005
R346 DVDD.n7548 DVDD.n7516 4.5005
R347 DVDD.n7530 DVDD.n2508 4.5005
R348 DVDD.n7548 DVDD.n7530 4.5005
R349 DVDD.n7515 DVDD.n2508 4.5005
R350 DVDD.n7548 DVDD.n7515 4.5005
R351 DVDD.n7531 DVDD.n2508 4.5005
R352 DVDD.n7548 DVDD.n7531 4.5005
R353 DVDD.n7514 DVDD.n2508 4.5005
R354 DVDD.n7548 DVDD.n7514 4.5005
R355 DVDD.n7532 DVDD.n2508 4.5005
R356 DVDD.n7548 DVDD.n7532 4.5005
R357 DVDD.n7513 DVDD.n2508 4.5005
R358 DVDD.n7548 DVDD.n7513 4.5005
R359 DVDD.n7533 DVDD.n2508 4.5005
R360 DVDD.n7548 DVDD.n7533 4.5005
R361 DVDD.n7512 DVDD.n2508 4.5005
R362 DVDD.n7548 DVDD.n7512 4.5005
R363 DVDD.n7547 DVDD.n2508 4.5005
R364 DVDD.n7548 DVDD.n7547 4.5005
R365 DVDD.n7511 DVDD.n2508 4.5005
R366 DVDD.n7548 DVDD.n7511 4.5005
R367 DVDD.n7550 DVDD.n7549 4.5005
R368 DVDD.n7549 DVDD.n2508 4.5005
R369 DVDD.n7549 DVDD.n7548 4.5005
R370 DVDD.n7509 DVDD.n7029 4.5005
R371 DVDD.n7509 DVDD.n7030 4.5005
R372 DVDD.n7509 DVDD.n7508 4.5005
R373 DVDD.n7045 DVDD.n7030 4.5005
R374 DVDD.n7508 DVDD.n7045 4.5005
R375 DVDD.n7042 DVDD.n7030 4.5005
R376 DVDD.n7508 DVDD.n7042 4.5005
R377 DVDD.n7047 DVDD.n7030 4.5005
R378 DVDD.n7508 DVDD.n7047 4.5005
R379 DVDD.n7041 DVDD.n7030 4.5005
R380 DVDD.n7508 DVDD.n7041 4.5005
R381 DVDD.n7049 DVDD.n7030 4.5005
R382 DVDD.n7508 DVDD.n7049 4.5005
R383 DVDD.n7040 DVDD.n7030 4.5005
R384 DVDD.n7508 DVDD.n7040 4.5005
R385 DVDD.n7051 DVDD.n7030 4.5005
R386 DVDD.n7508 DVDD.n7051 4.5005
R387 DVDD.n7039 DVDD.n7030 4.5005
R388 DVDD.n7508 DVDD.n7039 4.5005
R389 DVDD.n7053 DVDD.n7030 4.5005
R390 DVDD.n7508 DVDD.n7053 4.5005
R391 DVDD.n7038 DVDD.n7030 4.5005
R392 DVDD.n7508 DVDD.n7038 4.5005
R393 DVDD.n7055 DVDD.n7030 4.5005
R394 DVDD.n7508 DVDD.n7055 4.5005
R395 DVDD.n7037 DVDD.n7030 4.5005
R396 DVDD.n7508 DVDD.n7037 4.5005
R397 DVDD.n7057 DVDD.n7030 4.5005
R398 DVDD.n7508 DVDD.n7057 4.5005
R399 DVDD.n7036 DVDD.n7030 4.5005
R400 DVDD.n7508 DVDD.n7036 4.5005
R401 DVDD.n7059 DVDD.n7030 4.5005
R402 DVDD.n7508 DVDD.n7059 4.5005
R403 DVDD.n7035 DVDD.n7030 4.5005
R404 DVDD.n7508 DVDD.n7035 4.5005
R405 DVDD.n7061 DVDD.n7030 4.5005
R406 DVDD.n7508 DVDD.n7061 4.5005
R407 DVDD.n7034 DVDD.n7030 4.5005
R408 DVDD.n7508 DVDD.n7034 4.5005
R409 DVDD.n7063 DVDD.n7030 4.5005
R410 DVDD.n7508 DVDD.n7063 4.5005
R411 DVDD.n7033 DVDD.n7030 4.5005
R412 DVDD.n7508 DVDD.n7033 4.5005
R413 DVDD.n7065 DVDD.n7030 4.5005
R414 DVDD.n7508 DVDD.n7065 4.5005
R415 DVDD.n7032 DVDD.n7030 4.5005
R416 DVDD.n7508 DVDD.n7032 4.5005
R417 DVDD.n7507 DVDD.n7029 4.5005
R418 DVDD.n7507 DVDD.n7030 4.5005
R419 DVDD.n7508 DVDD.n7507 4.5005
R420 DVDD.n6543 DVDD.n6542 4.5005
R421 DVDD.n6541 DVDD.n6540 4.5005
R422 DVDD.n6539 DVDD.n6538 4.5005
R423 DVDD.n6537 DVDD.n6536 4.5005
R424 DVDD.n6535 DVDD.n6534 4.5005
R425 DVDD.n6533 DVDD.n6532 4.5005
R426 DVDD.n6531 DVDD.n6530 4.5005
R427 DVDD.n6529 DVDD.n6528 4.5005
R428 DVDD.n6527 DVDD.n3356 4.5005
R429 DVDD.n6526 DVDD.n3358 4.5005
R430 DVDD.n6525 DVDD.n6524 4.5005
R431 DVDD.n6523 DVDD.n6522 4.5005
R432 DVDD.n6521 DVDD.n6520 4.5005
R433 DVDD.n6519 DVDD.n6518 4.5005
R434 DVDD.n6517 DVDD.n6516 4.5005
R435 DVDD.n6515 DVDD.n6514 4.5005
R436 DVDD.n6513 DVDD.n6512 4.5005
R437 DVDD.n6511 DVDD.n6510 4.5005
R438 DVDD.n6509 DVDD.n6508 4.5005
R439 DVDD.n6507 DVDD.n6506 4.5005
R440 DVDD.n6505 DVDD.n6504 4.5005
R441 DVDD.n6503 DVDD.n6502 4.5005
R442 DVDD.n6501 DVDD.n6500 4.5005
R443 DVDD.n6499 DVDD.n6498 4.5005
R444 DVDD.n6497 DVDD.n6496 4.5005
R445 DVDD.n6495 DVDD.n6494 4.5005
R446 DVDD.n6493 DVDD.n6492 4.5005
R447 DVDD.n6491 DVDD.n6490 4.5005
R448 DVDD.n6489 DVDD.n6488 4.5005
R449 DVDD.n6300 DVDD.n3417 4.5005
R450 DVDD.n6298 DVDD.n6297 4.5005
R451 DVDD.n6296 DVDD.n6245 4.5005
R452 DVDD.n6295 DVDD.n6294 4.5005
R453 DVDD.n6293 DVDD.n6246 4.5005
R454 DVDD.n6292 DVDD.n6291 4.5005
R455 DVDD.n6290 DVDD.n6247 4.5005
R456 DVDD.n6289 DVDD.n6288 4.5005
R457 DVDD.n6287 DVDD.n6248 4.5005
R458 DVDD.n6286 DVDD.n6285 4.5005
R459 DVDD.n6284 DVDD.n6249 4.5005
R460 DVDD.n6283 DVDD.n6282 4.5005
R461 DVDD.n6281 DVDD.n6250 4.5005
R462 DVDD.n6280 DVDD.n6279 4.5005
R463 DVDD.n6278 DVDD.n6251 4.5005
R464 DVDD.n6277 DVDD.n6276 4.5005
R465 DVDD.n6275 DVDD.n6252 4.5005
R466 DVDD.n6274 DVDD.n6273 4.5005
R467 DVDD.n6272 DVDD.n6253 4.5005
R468 DVDD.n6271 DVDD.n6270 4.5005
R469 DVDD.n6269 DVDD.n6268 4.5005
R470 DVDD.n6267 DVDD.n6266 4.5005
R471 DVDD.n6265 DVDD.n6264 4.5005
R472 DVDD.n6263 DVDD.n6262 4.5005
R473 DVDD.n6261 DVDD.n6260 4.5005
R474 DVDD.n6259 DVDD.n6258 4.5005
R475 DVDD.n6257 DVDD.n6256 4.5005
R476 DVDD.n6255 DVDD.n6254 4.5005
R477 DVDD.n3416 DVDD.n3415 4.5005
R478 DVDD.n6337 DVDD.n6336 4.5005
R479 DVDD.n3559 DVDD.n3555 4.5005
R480 DVDD.n3821 DVDD.n3820 4.5005
R481 DVDD.n3823 DVDD.n3822 4.5005
R482 DVDD.n3825 DVDD.n3824 4.5005
R483 DVDD.n3827 DVDD.n3826 4.5005
R484 DVDD.n3829 DVDD.n3828 4.5005
R485 DVDD.n3831 DVDD.n3830 4.5005
R486 DVDD.n3833 DVDD.n3832 4.5005
R487 DVDD.n3835 DVDD.n3834 4.5005
R488 DVDD.n3837 DVDD.n3836 4.5005
R489 DVDD.n3839 DVDD.n3838 4.5005
R490 DVDD.n3841 DVDD.n3840 4.5005
R491 DVDD.n3843 DVDD.n3842 4.5005
R492 DVDD.n3845 DVDD.n3844 4.5005
R493 DVDD.n3847 DVDD.n3846 4.5005
R494 DVDD.n3849 DVDD.n3848 4.5005
R495 DVDD.n3851 DVDD.n3850 4.5005
R496 DVDD.n3853 DVDD.n3852 4.5005
R497 DVDD.n3855 DVDD.n3854 4.5005
R498 DVDD.n3857 DVDD.n3856 4.5005
R499 DVDD.n3859 DVDD.n3858 4.5005
R500 DVDD.n3860 DVDD.n3818 4.5005
R501 DVDD.n6332 DVDD.n6331 4.5005
R502 DVDD.n6330 DVDD.n3819 4.5005
R503 DVDD.n6329 DVDD.n6328 4.5005
R504 DVDD.n3863 DVDD.n3861 4.5005
R505 DVDD.n6323 DVDD.n6322 4.5005
R506 DVDD.n3867 DVDD.n3554 4.5005
R507 DVDD.n3702 DVDD.n3577 4.5005
R508 DVDD.n3701 DVDD.n3700 4.5005
R509 DVDD.n3699 DVDD.n3650 4.5005
R510 DVDD.n3698 DVDD.n3697 4.5005
R511 DVDD.n3696 DVDD.n3651 4.5005
R512 DVDD.n3695 DVDD.n3694 4.5005
R513 DVDD.n3693 DVDD.n3652 4.5005
R514 DVDD.n3692 DVDD.n3691 4.5005
R515 DVDD.n3690 DVDD.n3653 4.5005
R516 DVDD.n3689 DVDD.n3688 4.5005
R517 DVDD.n3687 DVDD.n3654 4.5005
R518 DVDD.n3686 DVDD.n3685 4.5005
R519 DVDD.n3684 DVDD.n3655 4.5005
R520 DVDD.n3683 DVDD.n3682 4.5005
R521 DVDD.n3681 DVDD.n3656 4.5005
R522 DVDD.n3680 DVDD.n3679 4.5005
R523 DVDD.n3678 DVDD.n3657 4.5005
R524 DVDD.n3677 DVDD.n3676 4.5005
R525 DVDD.n3675 DVDD.n3658 4.5005
R526 DVDD.n3674 DVDD.n3673 4.5005
R527 DVDD.n3672 DVDD.n3659 4.5005
R528 DVDD.n3671 DVDD.n3670 4.5005
R529 DVDD.n3669 DVDD.n3660 4.5005
R530 DVDD.n3668 DVDD.n3667 4.5005
R531 DVDD.n3666 DVDD.n3661 4.5005
R532 DVDD.n3665 DVDD.n3664 4.5005
R533 DVDD.n3663 DVDD.n3662 4.5005
R534 DVDD.n3575 DVDD.n3574 4.5005
R535 DVDD.n3804 DVDD.n3803 4.5005
R536 DVDD.n3582 DVDD.n1010 4.5005
R537 DVDD.n3637 DVDD.n1041 4.5005
R538 DVDD.n3638 DVDD.n1042 4.5005
R539 DVDD.n3740 DVDD.n3739 4.5005
R540 DVDD.n3738 DVDD.n3636 4.5005
R541 DVDD.n3737 DVDD.n1049 4.5005
R542 DVDD.n3736 DVDD.n1050 4.5005
R543 DVDD.n3735 DVDD.n3734 4.5005
R544 DVDD.n3733 DVDD.n3639 4.5005
R545 DVDD.n3732 DVDD.n3731 4.5005
R546 DVDD.n3730 DVDD.n3641 4.5005
R547 DVDD.n3729 DVDD.n3728 4.5005
R548 DVDD.n3727 DVDD.n3642 4.5005
R549 DVDD.n3726 DVDD.n3725 4.5005
R550 DVDD.n3724 DVDD.n3643 4.5005
R551 DVDD.n3723 DVDD.n3722 4.5005
R552 DVDD.n3721 DVDD.n3644 4.5005
R553 DVDD.n3720 DVDD.n3719 4.5005
R554 DVDD.n3718 DVDD.n3645 4.5005
R555 DVDD.n3717 DVDD.n3716 4.5005
R556 DVDD.n3715 DVDD.n3646 4.5005
R557 DVDD.n3714 DVDD.n3713 4.5005
R558 DVDD.n3712 DVDD.n3647 4.5005
R559 DVDD.n3711 DVDD.n3710 4.5005
R560 DVDD.n3709 DVDD.n3648 4.5005
R561 DVDD.n3708 DVDD.n3707 4.5005
R562 DVDD.n3706 DVDD.n3649 4.5005
R563 DVDD.n3705 DVDD.n3704 4.5005
R564 DVDD.n3703 DVDD.n3581 4.5005
R565 DVDD.n9633 DVDD.n9632 4.5005
R566 DVDD.n9631 DVDD.n79 4.5005
R567 DVDD.n9630 DVDD.n9629 4.5005
R568 DVDD.n82 DVDD.n80 4.5005
R569 DVDD.n844 DVDD.n843 4.5005
R570 DVDD.n845 DVDD.n91 4.5005
R571 DVDD.n846 DVDD.n92 4.5005
R572 DVDD.n8770 DVDD.n8769 4.5005
R573 DVDD.n8768 DVDD.n8767 4.5005
R574 DVDD.n848 DVDD.n847 4.5005
R575 DVDD.n930 DVDD.n855 4.5005
R576 DVDD.n940 DVDD.n939 4.5005
R577 DVDD.n938 DVDD.n864 4.5005
R578 DVDD.n937 DVDD.n865 4.5005
R579 DVDD.n936 DVDD.n935 4.5005
R580 DVDD.n934 DVDD.n932 4.5005
R581 DVDD.n931 DVDD.n873 4.5005
R582 DVDD.n878 DVDD.n874 4.5005
R583 DVDD.n8744 DVDD.n8743 4.5005
R584 DVDD.n8742 DVDD.n8741 4.5005
R585 DVDD.n8740 DVDD.n879 4.5005
R586 DVDD.n887 DVDD.n880 4.5005
R587 DVDD.n8723 DVDD.n8722 4.5005
R588 DVDD.n8721 DVDD.n8720 4.5005
R589 DVDD.n889 DVDD.n888 4.5005
R590 DVDD.n914 DVDD.n896 4.5005
R591 DVDD.n916 DVDD.n915 4.5005
R592 DVDD.n998 DVDD.n997 4.5005
R593 DVDD.n999 DVDD.n904 4.5005
R594 DVDD.n8835 DVDD.n8834 4.5005
R595 DVDD.n8833 DVDD.n789 4.5005
R596 DVDD.n8832 DVDD.n8831 4.5005
R597 DVDD.n8830 DVDD.n8797 4.5005
R598 DVDD.n8829 DVDD.n8828 4.5005
R599 DVDD.n8827 DVDD.n8798 4.5005
R600 DVDD.n8826 DVDD.n8825 4.5005
R601 DVDD.n8824 DVDD.n8799 4.5005
R602 DVDD.n8823 DVDD.n8822 4.5005
R603 DVDD.n8821 DVDD.n8820 4.5005
R604 DVDD.n8819 DVDD.n8818 4.5005
R605 DVDD.n8817 DVDD.n8816 4.5005
R606 DVDD.n8815 DVDD.n8814 4.5005
R607 DVDD.n8813 DVDD.n8812 4.5005
R608 DVDD.n8811 DVDD.n8810 4.5005
R609 DVDD.n8809 DVDD.n8808 4.5005
R610 DVDD.n8807 DVDD.n8806 4.5005
R611 DVDD.n8805 DVDD.n8804 4.5005
R612 DVDD.n8803 DVDD.n8802 4.5005
R613 DVDD.n8801 DVDD.n8800 4.5005
R614 DVDD.n75 DVDD.n71 4.5005
R615 DVDD.n9645 DVDD.n9644 4.5005
R616 DVDD.n9643 DVDD.n74 4.5005
R617 DVDD.n9642 DVDD.n9641 4.5005
R618 DVDD.n9640 DVDD.n76 4.5005
R619 DVDD.n9639 DVDD.n9638 4.5005
R620 DVDD.n9637 DVDD.n77 4.5005
R621 DVDD.n9636 DVDD.n9635 4.5005
R622 DVDD.n9634 DVDD.n78 4.5005
R623 DVDD.n748 DVDD.n747 4.5005
R624 DVDD.n749 DVDD.n686 4.5005
R625 DVDD.n751 DVDD.n750 4.5005
R626 DVDD.n752 DVDD.n685 4.5005
R627 DVDD.n754 DVDD.n753 4.5005
R628 DVDD.n755 DVDD.n684 4.5005
R629 DVDD.n757 DVDD.n756 4.5005
R630 DVDD.n758 DVDD.n683 4.5005
R631 DVDD.n760 DVDD.n759 4.5005
R632 DVDD.n761 DVDD.n682 4.5005
R633 DVDD.n763 DVDD.n762 4.5005
R634 DVDD.n764 DVDD.n681 4.5005
R635 DVDD.n766 DVDD.n765 4.5005
R636 DVDD.n767 DVDD.n680 4.5005
R637 DVDD.n769 DVDD.n768 4.5005
R638 DVDD.n770 DVDD.n679 4.5005
R639 DVDD.n772 DVDD.n771 4.5005
R640 DVDD.n773 DVDD.n678 4.5005
R641 DVDD.n775 DVDD.n774 4.5005
R642 DVDD.n776 DVDD.n677 4.5005
R643 DVDD.n778 DVDD.n777 4.5005
R644 DVDD.n779 DVDD.n676 4.5005
R645 DVDD.n781 DVDD.n780 4.5005
R646 DVDD.n782 DVDD.n675 4.5005
R647 DVDD.n784 DVDD.n783 4.5005
R648 DVDD.n785 DVDD.n674 4.5005
R649 DVDD.n787 DVDD.n786 4.5005
R650 DVDD.n788 DVDD.n673 4.5005
R651 DVDD.n8837 DVDD.n8836 4.5005
R652 DVDD.n724 DVDD.n723 4.5005
R653 DVDD.n722 DVDD.n721 4.5005
R654 DVDD.n720 DVDD.n719 4.5005
R655 DVDD.n718 DVDD.n717 4.5005
R656 DVDD.n716 DVDD.n715 4.5005
R657 DVDD.n714 DVDD.n713 4.5005
R658 DVDD.n712 DVDD.n711 4.5005
R659 DVDD.n710 DVDD.n709 4.5005
R660 DVDD.n708 DVDD.n707 4.5005
R661 DVDD.n706 DVDD.n705 4.5005
R662 DVDD.n704 DVDD.n703 4.5005
R663 DVDD.n6334 DVDD.n3807 4.5005
R664 DVDD.n3807 DVDD.n3558 4.5005
R665 DVDD.n3807 DVDD.n3557 4.5005
R666 DVDD.n3805 DVDD.n3558 4.5005
R667 DVDD.n3805 DVDD.n3557 4.5005
R668 DVDD.n3572 DVDD.n3558 4.5005
R669 DVDD.n3572 DVDD.n3557 4.5005
R670 DVDD.n6334 DVDD.n3556 4.5005
R671 DVDD.n3558 DVDD.n3556 4.5005
R672 DVDD.n3557 DVDD.n3556 4.5005
R673 DVDD.n6335 DVDD.n3558 4.5005
R674 DVDD.n6335 DVDD.n3560 4.5005
R675 DVDD.n6335 DVDD.n3557 4.5005
R676 DVDD.n6335 DVDD.n6334 4.5005
R677 DVDD.n6334 DVDD.n3809 4.5005
R678 DVDD.n3809 DVDD.n3558 4.5005
R679 DVDD.n3809 DVDD.n3560 4.5005
R680 DVDD.n3809 DVDD.n3557 4.5005
R681 DVDD.n6334 DVDD.n3570 4.5005
R682 DVDD.n3570 DVDD.n3558 4.5005
R683 DVDD.n3570 DVDD.n3560 4.5005
R684 DVDD.n3570 DVDD.n3557 4.5005
R685 DVDD.n6334 DVDD.n3810 4.5005
R686 DVDD.n3810 DVDD.n3558 4.5005
R687 DVDD.n3810 DVDD.n3560 4.5005
R688 DVDD.n3810 DVDD.n3557 4.5005
R689 DVDD.n6334 DVDD.n3569 4.5005
R690 DVDD.n3569 DVDD.n3558 4.5005
R691 DVDD.n3569 DVDD.n3560 4.5005
R692 DVDD.n3569 DVDD.n3557 4.5005
R693 DVDD.n3811 DVDD.n3558 4.5005
R694 DVDD.n3811 DVDD.n3560 4.5005
R695 DVDD.n3811 DVDD.n3557 4.5005
R696 DVDD.n6334 DVDD.n3811 4.5005
R697 DVDD.n3568 DVDD.n3558 4.5005
R698 DVDD.n3568 DVDD.n3560 4.5005
R699 DVDD.n3568 DVDD.n3557 4.5005
R700 DVDD.n6334 DVDD.n3568 4.5005
R701 DVDD.n3812 DVDD.n3558 4.5005
R702 DVDD.n3812 DVDD.n3560 4.5005
R703 DVDD.n3812 DVDD.n3557 4.5005
R704 DVDD.n6334 DVDD.n3812 4.5005
R705 DVDD.n6334 DVDD.n3567 4.5005
R706 DVDD.n3567 DVDD.n3558 4.5005
R707 DVDD.n3567 DVDD.n3560 4.5005
R708 DVDD.n3567 DVDD.n3557 4.5005
R709 DVDD.n6334 DVDD.n3813 4.5005
R710 DVDD.n3813 DVDD.n3558 4.5005
R711 DVDD.n3813 DVDD.n3560 4.5005
R712 DVDD.n3813 DVDD.n3557 4.5005
R713 DVDD.n6334 DVDD.n3566 4.5005
R714 DVDD.n3566 DVDD.n3558 4.5005
R715 DVDD.n3566 DVDD.n3560 4.5005
R716 DVDD.n3566 DVDD.n3557 4.5005
R717 DVDD.n3814 DVDD.n3558 4.5005
R718 DVDD.n3814 DVDD.n3560 4.5005
R719 DVDD.n3814 DVDD.n3557 4.5005
R720 DVDD.n6334 DVDD.n3814 4.5005
R721 DVDD.n3565 DVDD.n3558 4.5005
R722 DVDD.n3565 DVDD.n3560 4.5005
R723 DVDD.n3565 DVDD.n3557 4.5005
R724 DVDD.n6334 DVDD.n3565 4.5005
R725 DVDD.n3815 DVDD.n3558 4.5005
R726 DVDD.n3815 DVDD.n3560 4.5005
R727 DVDD.n3815 DVDD.n3557 4.5005
R728 DVDD.n6334 DVDD.n3815 4.5005
R729 DVDD.n3564 DVDD.n3558 4.5005
R730 DVDD.n3564 DVDD.n3560 4.5005
R731 DVDD.n3564 DVDD.n3557 4.5005
R732 DVDD.n6334 DVDD.n3564 4.5005
R733 DVDD.n6334 DVDD.n3816 4.5005
R734 DVDD.n3816 DVDD.n3558 4.5005
R735 DVDD.n3816 DVDD.n3560 4.5005
R736 DVDD.n3816 DVDD.n3557 4.5005
R737 DVDD.n6334 DVDD.n3563 4.5005
R738 DVDD.n3563 DVDD.n3558 4.5005
R739 DVDD.n3563 DVDD.n3560 4.5005
R740 DVDD.n3563 DVDD.n3557 4.5005
R741 DVDD.n6334 DVDD.n3817 4.5005
R742 DVDD.n3817 DVDD.n3558 4.5005
R743 DVDD.n3817 DVDD.n3560 4.5005
R744 DVDD.n3817 DVDD.n3557 4.5005
R745 DVDD.n3562 DVDD.n3558 4.5005
R746 DVDD.n3562 DVDD.n3560 4.5005
R747 DVDD.n3562 DVDD.n3557 4.5005
R748 DVDD.n6334 DVDD.n3562 4.5005
R749 DVDD.n6333 DVDD.n3558 4.5005
R750 DVDD.n6333 DVDD.n3560 4.5005
R751 DVDD.n6333 DVDD.n3557 4.5005
R752 DVDD.n6334 DVDD.n6333 4.5005
R753 DVDD.n6327 DVDD.n3862 4.5005
R754 DVDD.n6327 DVDD.n3864 4.5005
R755 DVDD.n6324 DVDD.n3862 4.5005
R756 DVDD.n6324 DVDD.n3864 4.5005
R757 DVDD.n6321 DVDD.n3862 4.5005
R758 DVDD.n6321 DVDD.n3864 4.5005
R759 DVDD.n3874 DVDD.n3864 4.5005
R760 DVDD.n6301 DVDD.n3862 4.5005
R761 DVDD.n6299 DVDD.n3864 4.5005
R762 DVDD.n6299 DVDD.n3862 4.5005
R763 DVDD.n6648 DVDD.n3343 4.5005
R764 DVDD.n3357 DVDD.n3343 4.5005
R765 DVDD.n3362 DVDD.n3343 4.5005
R766 DVDD.n6650 DVDD.n3343 4.5005
R767 DVDD.n6648 DVDD.n3345 4.5005
R768 DVDD.n3357 DVDD.n3345 4.5005
R769 DVDD.n3362 DVDD.n3345 4.5005
R770 DVDD.n6650 DVDD.n3345 4.5005
R771 DVDD.n6648 DVDD.n3342 4.5005
R772 DVDD.n3357 DVDD.n3342 4.5005
R773 DVDD.n3362 DVDD.n3342 4.5005
R774 DVDD.n6650 DVDD.n3342 4.5005
R775 DVDD.n6648 DVDD.n3346 4.5005
R776 DVDD.n3357 DVDD.n3346 4.5005
R777 DVDD.n3362 DVDD.n3346 4.5005
R778 DVDD.n6650 DVDD.n3346 4.5005
R779 DVDD.n3357 DVDD.n3341 4.5005
R780 DVDD.n3362 DVDD.n3341 4.5005
R781 DVDD.n6650 DVDD.n3341 4.5005
R782 DVDD.n6648 DVDD.n3341 4.5005
R783 DVDD.n3357 DVDD.n3347 4.5005
R784 DVDD.n3362 DVDD.n3347 4.5005
R785 DVDD.n6650 DVDD.n3347 4.5005
R786 DVDD.n6648 DVDD.n3347 4.5005
R787 DVDD.n3357 DVDD.n3340 4.5005
R788 DVDD.n3362 DVDD.n3340 4.5005
R789 DVDD.n6650 DVDD.n3340 4.5005
R790 DVDD.n6648 DVDD.n3340 4.5005
R791 DVDD.n6648 DVDD.n3348 4.5005
R792 DVDD.n3357 DVDD.n3348 4.5005
R793 DVDD.n3362 DVDD.n3348 4.5005
R794 DVDD.n6650 DVDD.n3348 4.5005
R795 DVDD.n6648 DVDD.n3339 4.5005
R796 DVDD.n3357 DVDD.n3339 4.5005
R797 DVDD.n3362 DVDD.n3339 4.5005
R798 DVDD.n6650 DVDD.n3339 4.5005
R799 DVDD.n6648 DVDD.n3349 4.5005
R800 DVDD.n3357 DVDD.n3349 4.5005
R801 DVDD.n6650 DVDD.n3349 4.5005
R802 DVDD.n3357 DVDD.n3338 4.5005
R803 DVDD.n6650 DVDD.n3338 4.5005
R804 DVDD.n3357 DVDD.n3350 4.5005
R805 DVDD.n6650 DVDD.n3350 4.5005
R806 DVDD.n3357 DVDD.n3337 4.5005
R807 DVDD.n6650 DVDD.n3337 4.5005
R808 DVDD.n3357 DVDD.n3351 4.5005
R809 DVDD.n6650 DVDD.n3351 4.5005
R810 DVDD.n3357 DVDD.n3336 4.5005
R811 DVDD.n6650 DVDD.n3336 4.5005
R812 DVDD.n3357 DVDD.n3352 4.5005
R813 DVDD.n3362 DVDD.n3352 4.5005
R814 DVDD.n6650 DVDD.n3352 4.5005
R815 DVDD.n3357 DVDD.n3335 4.5005
R816 DVDD.n3362 DVDD.n3335 4.5005
R817 DVDD.n6650 DVDD.n3335 4.5005
R818 DVDD.n6648 DVDD.n3335 4.5005
R819 DVDD.n3357 DVDD.n3353 4.5005
R820 DVDD.n3362 DVDD.n3353 4.5005
R821 DVDD.n6650 DVDD.n3353 4.5005
R822 DVDD.n6648 DVDD.n3353 4.5005
R823 DVDD.n6648 DVDD.n3334 4.5005
R824 DVDD.n3357 DVDD.n3334 4.5005
R825 DVDD.n3362 DVDD.n3334 4.5005
R826 DVDD.n6650 DVDD.n3334 4.5005
R827 DVDD.n6648 DVDD.n3354 4.5005
R828 DVDD.n3357 DVDD.n3354 4.5005
R829 DVDD.n3362 DVDD.n3354 4.5005
R830 DVDD.n6650 DVDD.n3354 4.5005
R831 DVDD.n6648 DVDD.n3333 4.5005
R832 DVDD.n3357 DVDD.n3333 4.5005
R833 DVDD.n3362 DVDD.n3333 4.5005
R834 DVDD.n6650 DVDD.n3333 4.5005
R835 DVDD.n3357 DVDD.n3355 4.5005
R836 DVDD.n3362 DVDD.n3355 4.5005
R837 DVDD.n6650 DVDD.n3355 4.5005
R838 DVDD.n6648 DVDD.n3355 4.5005
R839 DVDD.n3357 DVDD.n3332 4.5005
R840 DVDD.n3362 DVDD.n3332 4.5005
R841 DVDD.n6650 DVDD.n3332 4.5005
R842 DVDD.n6648 DVDD.n3332 4.5005
R843 DVDD.n6649 DVDD.n3357 4.5005
R844 DVDD.n6649 DVDD.n3362 4.5005
R845 DVDD.n6650 DVDD.n6649 4.5005
R846 DVDD.n6649 DVDD.n6648 4.5005
R847 DVDD.n7893 DVDD.n2082 4.5005
R848 DVDD.n2096 DVDD.n2082 4.5005
R849 DVDD.n7886 DVDD.n2082 4.5005
R850 DVDD.n7890 DVDD.n2082 4.5005
R851 DVDD.n7893 DVDD.n2083 4.5005
R852 DVDD.n2096 DVDD.n2083 4.5005
R853 DVDD.n7886 DVDD.n2083 4.5005
R854 DVDD.n7890 DVDD.n2083 4.5005
R855 DVDD.n7893 DVDD.n2081 4.5005
R856 DVDD.n2096 DVDD.n2081 4.5005
R857 DVDD.n7886 DVDD.n2081 4.5005
R858 DVDD.n7890 DVDD.n2081 4.5005
R859 DVDD.n2096 DVDD.n2084 4.5005
R860 DVDD.n7886 DVDD.n2084 4.5005
R861 DVDD.n7890 DVDD.n2084 4.5005
R862 DVDD.n7893 DVDD.n2084 4.5005
R863 DVDD.n2096 DVDD.n2080 4.5005
R864 DVDD.n7886 DVDD.n2080 4.5005
R865 DVDD.n7890 DVDD.n2080 4.5005
R866 DVDD.n7893 DVDD.n2080 4.5005
R867 DVDD.n2096 DVDD.n2085 4.5005
R868 DVDD.n7886 DVDD.n2085 4.5005
R869 DVDD.n7890 DVDD.n2085 4.5005
R870 DVDD.n7893 DVDD.n2085 4.5005
R871 DVDD.n2096 DVDD.n2079 4.5005
R872 DVDD.n7886 DVDD.n2079 4.5005
R873 DVDD.n7890 DVDD.n2079 4.5005
R874 DVDD.n7893 DVDD.n2079 4.5005
R875 DVDD.n7893 DVDD.n2086 4.5005
R876 DVDD.n2096 DVDD.n2086 4.5005
R877 DVDD.n7886 DVDD.n2086 4.5005
R878 DVDD.n7890 DVDD.n2086 4.5005
R879 DVDD.n7893 DVDD.n2078 4.5005
R880 DVDD.n2096 DVDD.n2078 4.5005
R881 DVDD.n7886 DVDD.n2078 4.5005
R882 DVDD.n7890 DVDD.n2078 4.5005
R883 DVDD.n7893 DVDD.n2087 4.5005
R884 DVDD.n2096 DVDD.n2087 4.5005
R885 DVDD.n7886 DVDD.n2087 4.5005
R886 DVDD.n7890 DVDD.n2087 4.5005
R887 DVDD.n2096 DVDD.n2077 4.5005
R888 DVDD.n7886 DVDD.n2077 4.5005
R889 DVDD.n7890 DVDD.n2077 4.5005
R890 DVDD.n7893 DVDD.n2077 4.5005
R891 DVDD.n2096 DVDD.n2088 4.5005
R892 DVDD.n7886 DVDD.n2088 4.5005
R893 DVDD.n7890 DVDD.n2088 4.5005
R894 DVDD.n7893 DVDD.n2088 4.5005
R895 DVDD.n2096 DVDD.n2076 4.5005
R896 DVDD.n7886 DVDD.n2076 4.5005
R897 DVDD.n7890 DVDD.n2076 4.5005
R898 DVDD.n7893 DVDD.n2076 4.5005
R899 DVDD.n7893 DVDD.n2089 4.5005
R900 DVDD.n2096 DVDD.n2089 4.5005
R901 DVDD.n7886 DVDD.n2089 4.5005
R902 DVDD.n7890 DVDD.n2089 4.5005
R903 DVDD.n7893 DVDD.n2075 4.5005
R904 DVDD.n2096 DVDD.n2075 4.5005
R905 DVDD.n7886 DVDD.n2075 4.5005
R906 DVDD.n7890 DVDD.n2075 4.5005
R907 DVDD.n7893 DVDD.n2090 4.5005
R908 DVDD.n2096 DVDD.n2090 4.5005
R909 DVDD.n7890 DVDD.n2090 4.5005
R910 DVDD.n2100 DVDD.n2096 4.5005
R911 DVDD.n7890 DVDD.n2100 4.5005
R912 DVDD.n2102 DVDD.n2096 4.5005
R913 DVDD.n7890 DVDD.n2102 4.5005
R914 DVDD.n2099 DVDD.n2096 4.5005
R915 DVDD.n7890 DVDD.n2099 4.5005
R916 DVDD.n7888 DVDD.n2096 4.5005
R917 DVDD.n7890 DVDD.n7888 4.5005
R918 DVDD.n2098 DVDD.n2096 4.5005
R919 DVDD.n7890 DVDD.n2098 4.5005
R920 DVDD.n7889 DVDD.n2096 4.5005
R921 DVDD.n7890 DVDD.n7889 4.5005
R922 DVDD.n7891 DVDD.n2096 4.5005
R923 DVDD.n7891 DVDD.n7890 4.5005
R924 DVDD.n2096 DVDD.n2094 4.5005
R925 DVDD.n7886 DVDD.n2094 4.5005
R926 DVDD.n7890 DVDD.n2094 4.5005
R927 DVDD.n8052 DVDD.n1972 4.5005
R928 DVDD.n8054 DVDD.n1972 4.5005
R929 DVDD.n1972 DVDD.n1947 4.5005
R930 DVDD.n8054 DVDD.n1974 4.5005
R931 DVDD.n1974 DVDD.n1947 4.5005
R932 DVDD.n8054 DVDD.n1971 4.5005
R933 DVDD.n1971 DVDD.n1947 4.5005
R934 DVDD.n8054 DVDD.n1975 4.5005
R935 DVDD.n1975 DVDD.n1947 4.5005
R936 DVDD.n8054 DVDD.n1970 4.5005
R937 DVDD.n1970 DVDD.n1947 4.5005
R938 DVDD.n8052 DVDD.n1976 4.5005
R939 DVDD.n8054 DVDD.n1976 4.5005
R940 DVDD.n1976 DVDD.n1947 4.5005
R941 DVDD.n8052 DVDD.n1953 4.5005
R942 DVDD.n8054 DVDD.n1953 4.5005
R943 DVDD.n8056 DVDD.n1953 4.5005
R944 DVDD.n1953 DVDD.n1947 4.5005
R945 DVDD.n8052 DVDD.n1977 4.5005
R946 DVDD.n8054 DVDD.n1977 4.5005
R947 DVDD.n1977 DVDD.n1947 4.5005
R948 DVDD.n8054 DVDD.n1969 4.5005
R949 DVDD.n1969 DVDD.n1947 4.5005
R950 DVDD.n8054 DVDD.n1978 4.5005
R951 DVDD.n1978 DVDD.n1947 4.5005
R952 DVDD.n8054 DVDD.n1968 4.5005
R953 DVDD.n1968 DVDD.n1947 4.5005
R954 DVDD.n8054 DVDD.n1979 4.5005
R955 DVDD.n1979 DVDD.n1947 4.5005
R956 DVDD.n8052 DVDD.n1967 4.5005
R957 DVDD.n8054 DVDD.n1967 4.5005
R958 DVDD.n1967 DVDD.n1947 4.5005
R959 DVDD.n8052 DVDD.n1958 4.5005
R960 DVDD.n8054 DVDD.n1958 4.5005
R961 DVDD.n8056 DVDD.n1958 4.5005
R962 DVDD.n1958 DVDD.n1947 4.5005
R963 DVDD.n8052 DVDD.n1966 4.5005
R964 DVDD.n8054 DVDD.n1966 4.5005
R965 DVDD.n1966 DVDD.n1947 4.5005
R966 DVDD.n8054 DVDD.n1980 4.5005
R967 DVDD.n1980 DVDD.n1947 4.5005
R968 DVDD.n8054 DVDD.n1965 4.5005
R969 DVDD.n1965 DVDD.n1947 4.5005
R970 DVDD.n8054 DVDD.n1981 4.5005
R971 DVDD.n1981 DVDD.n1947 4.5005
R972 DVDD.n8054 DVDD.n1964 4.5005
R973 DVDD.n1964 DVDD.n1947 4.5005
R974 DVDD.n8052 DVDD.n1982 4.5005
R975 DVDD.n8054 DVDD.n1982 4.5005
R976 DVDD.n1982 DVDD.n1947 4.5005
R977 DVDD.n8052 DVDD.n1949 4.5005
R978 DVDD.n8054 DVDD.n1949 4.5005
R979 DVDD.n8056 DVDD.n1949 4.5005
R980 DVDD.n1949 DVDD.n1947 4.5005
R981 DVDD.n8053 DVDD.n8052 4.5005
R982 DVDD.n8054 DVDD.n8053 4.5005
R983 DVDD.n8053 DVDD.n1947 4.5005
R984 DVDD.n8054 DVDD.n1963 4.5005
R985 DVDD.n1963 DVDD.n1947 4.5005
R986 DVDD.n8055 DVDD.n8054 4.5005
R987 DVDD.n8056 DVDD.n8055 4.5005
R988 DVDD.n8055 DVDD.n1947 4.5005
R989 DVDD.n8120 DVDD.n1865 4.5005
R990 DVDD.n1891 DVDD.n1865 4.5005
R991 DVDD.n8115 DVDD.n1865 4.5005
R992 DVDD.n8118 DVDD.n1865 4.5005
R993 DVDD.n8118 DVDD.n1885 4.5005
R994 DVDD.n8115 DVDD.n1885 4.5005
R995 DVDD.n1891 DVDD.n1885 4.5005
R996 DVDD.n8120 DVDD.n1885 4.5005
R997 DVDD.n8120 DVDD.n1864 4.5005
R998 DVDD.n1891 DVDD.n1864 4.5005
R999 DVDD.n8118 DVDD.n1864 4.5005
R1000 DVDD.n1900 DVDD.n1891 4.5005
R1001 DVDD.n8118 DVDD.n1900 4.5005
R1002 DVDD.n1898 DVDD.n1891 4.5005
R1003 DVDD.n8118 DVDD.n1898 4.5005
R1004 DVDD.n1901 DVDD.n1891 4.5005
R1005 DVDD.n8118 DVDD.n1901 4.5005
R1006 DVDD.n1897 DVDD.n1891 4.5005
R1007 DVDD.n8118 DVDD.n1897 4.5005
R1008 DVDD.n8120 DVDD.n1886 4.5005
R1009 DVDD.n1891 DVDD.n1886 4.5005
R1010 DVDD.n8118 DVDD.n1886 4.5005
R1011 DVDD.n8118 DVDD.n1861 4.5005
R1012 DVDD.n8115 DVDD.n1861 4.5005
R1013 DVDD.n1891 DVDD.n1861 4.5005
R1014 DVDD.n8120 DVDD.n1861 4.5005
R1015 DVDD.n8118 DVDD.n1887 4.5005
R1016 DVDD.n8115 DVDD.n1887 4.5005
R1017 DVDD.n1891 DVDD.n1887 4.5005
R1018 DVDD.n8120 DVDD.n1887 4.5005
R1019 DVDD.n8120 DVDD.n1860 4.5005
R1020 DVDD.n1891 DVDD.n1860 4.5005
R1021 DVDD.n8118 DVDD.n1860 4.5005
R1022 DVDD.n1902 DVDD.n1891 4.5005
R1023 DVDD.n8118 DVDD.n1902 4.5005
R1024 DVDD.n1896 DVDD.n1891 4.5005
R1025 DVDD.n8118 DVDD.n1896 4.5005
R1026 DVDD.n1903 DVDD.n1891 4.5005
R1027 DVDD.n8118 DVDD.n1903 4.5005
R1028 DVDD.n1895 DVDD.n1891 4.5005
R1029 DVDD.n8115 DVDD.n1895 4.5005
R1030 DVDD.n8118 DVDD.n1895 4.5005
R1031 DVDD.n8120 DVDD.n1888 4.5005
R1032 DVDD.n1891 DVDD.n1888 4.5005
R1033 DVDD.n8115 DVDD.n1888 4.5005
R1034 DVDD.n8118 DVDD.n1888 4.5005
R1035 DVDD.n8120 DVDD.n1857 4.5005
R1036 DVDD.n1891 DVDD.n1857 4.5005
R1037 DVDD.n8115 DVDD.n1857 4.5005
R1038 DVDD.n8118 DVDD.n1857 4.5005
R1039 DVDD.n8120 DVDD.n1889 4.5005
R1040 DVDD.n1891 DVDD.n1889 4.5005
R1041 DVDD.n8115 DVDD.n1889 4.5005
R1042 DVDD.n8118 DVDD.n1889 4.5005
R1043 DVDD.n8120 DVDD.n1856 4.5005
R1044 DVDD.n1891 DVDD.n1856 4.5005
R1045 DVDD.n8118 DVDD.n1856 4.5005
R1046 DVDD.n1904 DVDD.n1891 4.5005
R1047 DVDD.n8118 DVDD.n1904 4.5005
R1048 DVDD.n1894 DVDD.n1891 4.5005
R1049 DVDD.n8118 DVDD.n1894 4.5005
R1050 DVDD.n8117 DVDD.n1891 4.5005
R1051 DVDD.n8118 DVDD.n8117 4.5005
R1052 DVDD.n1893 DVDD.n1891 4.5005
R1053 DVDD.n8118 DVDD.n1893 4.5005
R1054 DVDD.n8120 DVDD.n8119 4.5005
R1055 DVDD.n8119 DVDD.n1891 4.5005
R1056 DVDD.n8119 DVDD.n8118 4.5005
R1057 DVDD.n702 DVDD.n588 4.5005
R1058 DVDD.n701 DVDD.n590 4.5005
R1059 DVDD.n700 DVDD.n699 4.5005
R1060 DVDD.n698 DVDD.n689 4.5005
R1061 DVDD.n697 DVDD.n696 4.5005
R1062 DVDD.n695 DVDD.n690 4.5005
R1063 DVDD.n694 DVDD.n693 4.5005
R1064 DVDD.n692 DVDD.n691 4.5005
R1065 DVDD.n688 DVDD.n687 4.5005
R1066 DVDD.n746 DVDD.n745 4.5005
R1067 DVDD.n8538 DVDD.n1360 4.5005
R1068 DVDD.n8532 DVDD.n1360 4.5005
R1069 DVDD.n8535 DVDD.n8522 4.5005
R1070 DVDD.n8532 DVDD.n8522 4.5005
R1071 DVDD.n1450 DVDD.n1328 4.5005
R1072 DVDD.n8440 DVDD.n1328 4.5005
R1073 DVDD.n8627 DVDD.n1324 4.5005
R1074 DVDD.n8627 DVDD.n8626 4.5005
R1075 DVDD.n8625 DVDD.n8624 4.5005
R1076 DVDD.n8626 DVDD.n8625 4.5005
R1077 DVDD.n8440 DVDD.n8439 4.5005
R1078 DVDD.n8439 DVDD.n1450 4.5005
R1079 DVDD.n8439 DVDD.n8438 4.5005
R1080 DVDD.n1450 DVDD.n1432 4.5005
R1081 DVDD.n8438 DVDD.n1432 4.5005
R1082 DVDD.n8495 DVDD.n1434 4.5005
R1083 DVDD.n8495 DVDD.n8494 4.5005
R1084 DVDD.n8494 DVDD.n1429 4.5005
R1085 DVDD.n1434 DVDD.n1429 4.5005
R1086 DVDD.n8497 DVDD.n1429 4.5005
R1087 DVDD.n1434 DVDD.n1354 4.5005
R1088 DVDD.n8497 DVDD.n1354 4.5005
R1089 DVDD.n8600 DVDD.n8599 4.5005
R1090 DVDD.n8601 DVDD.n8600 4.5005
R1091 DVDD.n8601 DVDD.n1353 4.5005
R1092 DVDD.n8599 DVDD.n1353 4.5005
R1093 DVDD.n8597 DVDD.n1353 4.5005
R1094 DVDD.n8599 DVDD.n8598 4.5005
R1095 DVDD.n8598 DVDD.n8597 4.5005
R1096 DVDD.n1876 DVDD.n1677 4.5005
R1097 DVDD.n1687 DVDD.n1678 4.5005
R1098 DVDD.n8290 DVDD.n1687 4.5005
R1099 DVDD.n1687 DVDD.n1660 4.5005
R1100 DVDD.n8290 DVDD.n1690 4.5005
R1101 DVDD.n1690 DVDD.n1660 4.5005
R1102 DVDD.n8290 DVDD.n1686 4.5005
R1103 DVDD.n1686 DVDD.n1660 4.5005
R1104 DVDD.n8290 DVDD.n1692 4.5005
R1105 DVDD.n1692 DVDD.n1660 4.5005
R1106 DVDD.n8290 DVDD.n1685 4.5005
R1107 DVDD.n1685 DVDD.n1660 4.5005
R1108 DVDD.n1693 DVDD.n1678 4.5005
R1109 DVDD.n8290 DVDD.n1693 4.5005
R1110 DVDD.n1693 DVDD.n1660 4.5005
R1111 DVDD.n1664 DVDD.n1660 4.5005
R1112 DVDD.n8292 DVDD.n1664 4.5005
R1113 DVDD.n8290 DVDD.n1664 4.5005
R1114 DVDD.n1678 DVDD.n1664 4.5005
R1115 DVDD.n1669 DVDD.n1660 4.5005
R1116 DVDD.n8292 DVDD.n1669 4.5005
R1117 DVDD.n8290 DVDD.n1669 4.5005
R1118 DVDD.n1678 DVDD.n1669 4.5005
R1119 DVDD.n1684 DVDD.n1678 4.5005
R1120 DVDD.n8290 DVDD.n1684 4.5005
R1121 DVDD.n1684 DVDD.n1660 4.5005
R1122 DVDD.n8290 DVDD.n1695 4.5005
R1123 DVDD.n1695 DVDD.n1660 4.5005
R1124 DVDD.n8290 DVDD.n1683 4.5005
R1125 DVDD.n1683 DVDD.n1660 4.5005
R1126 DVDD.n8290 DVDD.n1697 4.5005
R1127 DVDD.n1697 DVDD.n1660 4.5005
R1128 DVDD.n8290 DVDD.n1663 4.5005
R1129 DVDD.n8292 DVDD.n1663 4.5005
R1130 DVDD.n1663 DVDD.n1660 4.5005
R1131 DVDD.n1678 DVDD.n1672 4.5005
R1132 DVDD.n8290 DVDD.n1672 4.5005
R1133 DVDD.n8292 DVDD.n1672 4.5005
R1134 DVDD.n1672 DVDD.n1660 4.5005
R1135 DVDD.n1678 DVDD.n1662 4.5005
R1136 DVDD.n8290 DVDD.n1662 4.5005
R1137 DVDD.n8292 DVDD.n1662 4.5005
R1138 DVDD.n1662 DVDD.n1660 4.5005
R1139 DVDD.n1678 DVDD.n1673 4.5005
R1140 DVDD.n8290 DVDD.n1673 4.5005
R1141 DVDD.n8292 DVDD.n1673 4.5005
R1142 DVDD.n1673 DVDD.n1660 4.5005
R1143 DVDD.n1682 DVDD.n1678 4.5005
R1144 DVDD.n8290 DVDD.n1682 4.5005
R1145 DVDD.n1682 DVDD.n1660 4.5005
R1146 DVDD.n8290 DVDD.n1699 4.5005
R1147 DVDD.n1699 DVDD.n1660 4.5005
R1148 DVDD.n8290 DVDD.n1681 4.5005
R1149 DVDD.n1681 DVDD.n1660 4.5005
R1150 DVDD.n8290 DVDD.n1701 4.5005
R1151 DVDD.n1701 DVDD.n1660 4.5005
R1152 DVDD.n8290 DVDD.n1680 4.5005
R1153 DVDD.n1680 DVDD.n1660 4.5005
R1154 DVDD.n8289 DVDD.n1678 4.5005
R1155 DVDD.n8290 DVDD.n8289 4.5005
R1156 DVDD.n8289 DVDD.n1660 4.5005
R1157 DVDD.n1661 DVDD.n1660 4.5005
R1158 DVDD.n8292 DVDD.n1661 4.5005
R1159 DVDD.n8290 DVDD.n1661 4.5005
R1160 DVDD.n1678 DVDD.n1661 4.5005
R1161 DVDD.n7749 DVDD.n2284 4.5005
R1162 DVDD.n2294 DVDD.n2284 4.5005
R1163 DVDD.n7747 DVDD.n2284 4.5005
R1164 DVDD.n2318 DVDD.n2294 4.5005
R1165 DVDD.n7747 DVDD.n2318 4.5005
R1166 DVDD.n2306 DVDD.n2294 4.5005
R1167 DVDD.n2306 DVDD.n2292 4.5005
R1168 DVDD.n7747 DVDD.n2306 4.5005
R1169 DVDD.n2320 DVDD.n2294 4.5005
R1170 DVDD.n7747 DVDD.n2320 4.5005
R1171 DVDD.n2305 DVDD.n2294 4.5005
R1172 DVDD.n7747 DVDD.n2305 4.5005
R1173 DVDD.n2322 DVDD.n2294 4.5005
R1174 DVDD.n7747 DVDD.n2322 4.5005
R1175 DVDD.n2304 DVDD.n2294 4.5005
R1176 DVDD.n7747 DVDD.n2304 4.5005
R1177 DVDD.n2323 DVDD.n2294 4.5005
R1178 DVDD.n2323 DVDD.n2292 4.5005
R1179 DVDD.n7747 DVDD.n2323 4.5005
R1180 DVDD.n2303 DVDD.n2294 4.5005
R1181 DVDD.n7747 DVDD.n2303 4.5005
R1182 DVDD.n2325 DVDD.n2294 4.5005
R1183 DVDD.n7747 DVDD.n2325 4.5005
R1184 DVDD.n2302 DVDD.n2294 4.5005
R1185 DVDD.n7747 DVDD.n2302 4.5005
R1186 DVDD.n2327 DVDD.n2294 4.5005
R1187 DVDD.n7747 DVDD.n2327 4.5005
R1188 DVDD.n2301 DVDD.n2294 4.5005
R1189 DVDD.n2301 DVDD.n2292 4.5005
R1190 DVDD.n7747 DVDD.n2301 4.5005
R1191 DVDD.n2329 DVDD.n2294 4.5005
R1192 DVDD.n7747 DVDD.n2329 4.5005
R1193 DVDD.n2300 DVDD.n2294 4.5005
R1194 DVDD.n7747 DVDD.n2300 4.5005
R1195 DVDD.n2331 DVDD.n2294 4.5005
R1196 DVDD.n7747 DVDD.n2331 4.5005
R1197 DVDD.n2299 DVDD.n2294 4.5005
R1198 DVDD.n7747 DVDD.n2299 4.5005
R1199 DVDD.n7746 DVDD.n2294 4.5005
R1200 DVDD.n7746 DVDD.n2292 4.5005
R1201 DVDD.n7747 DVDD.n7746 4.5005
R1202 DVDD.n7851 DVDD.n2132 4.5005
R1203 DVDD.n7853 DVDD.n2132 4.5005
R1204 DVDD.n7851 DVDD.n2133 4.5005
R1205 DVDD.n7853 DVDD.n2133 4.5005
R1206 DVDD.n7851 DVDD.n2131 4.5005
R1207 DVDD.n7853 DVDD.n2131 4.5005
R1208 DVDD.n7851 DVDD.n2134 4.5005
R1209 DVDD.n7853 DVDD.n2134 4.5005
R1210 DVDD.n7851 DVDD.n2130 4.5005
R1211 DVDD.n7853 DVDD.n2130 4.5005
R1212 DVDD.n7851 DVDD.n2135 4.5005
R1213 DVDD.n7853 DVDD.n2135 4.5005
R1214 DVDD.n7851 DVDD.n2129 4.5005
R1215 DVDD.n7853 DVDD.n2129 4.5005
R1216 DVDD.n7842 DVDD.n2136 4.5005
R1217 DVDD.n7851 DVDD.n2136 4.5005
R1218 DVDD.n7853 DVDD.n2136 4.5005
R1219 DVDD.n7851 DVDD.n2128 4.5005
R1220 DVDD.n2149 DVDD.n2128 4.5005
R1221 DVDD.n7853 DVDD.n2128 4.5005
R1222 DVDD.n7851 DVDD.n2137 4.5005
R1223 DVDD.n2149 DVDD.n2137 4.5005
R1224 DVDD.n7853 DVDD.n2137 4.5005
R1225 DVDD.n7842 DVDD.n2127 4.5005
R1226 DVDD.n7851 DVDD.n2127 4.5005
R1227 DVDD.n2149 DVDD.n2127 4.5005
R1228 DVDD.n7853 DVDD.n2127 4.5005
R1229 DVDD.n7842 DVDD.n2138 4.5005
R1230 DVDD.n7851 DVDD.n2138 4.5005
R1231 DVDD.n2149 DVDD.n2138 4.5005
R1232 DVDD.n7853 DVDD.n2138 4.5005
R1233 DVDD.n7842 DVDD.n2126 4.5005
R1234 DVDD.n7851 DVDD.n2126 4.5005
R1235 DVDD.n2149 DVDD.n2126 4.5005
R1236 DVDD.n7853 DVDD.n2126 4.5005
R1237 DVDD.n7851 DVDD.n2139 4.5005
R1238 DVDD.n2149 DVDD.n2139 4.5005
R1239 DVDD.n7853 DVDD.n2139 4.5005
R1240 DVDD.n7851 DVDD.n2125 4.5005
R1241 DVDD.n2149 DVDD.n2125 4.5005
R1242 DVDD.n7853 DVDD.n2125 4.5005
R1243 DVDD.n7851 DVDD.n2140 4.5005
R1244 DVDD.n2149 DVDD.n2140 4.5005
R1245 DVDD.n7853 DVDD.n2140 4.5005
R1246 DVDD.n7842 DVDD.n2124 4.5005
R1247 DVDD.n7851 DVDD.n2124 4.5005
R1248 DVDD.n2149 DVDD.n2124 4.5005
R1249 DVDD.n7853 DVDD.n2124 4.5005
R1250 DVDD.n7842 DVDD.n2141 4.5005
R1251 DVDD.n7851 DVDD.n2141 4.5005
R1252 DVDD.n2149 DVDD.n2141 4.5005
R1253 DVDD.n7853 DVDD.n2141 4.5005
R1254 DVDD.n7842 DVDD.n2123 4.5005
R1255 DVDD.n7851 DVDD.n2123 4.5005
R1256 DVDD.n2149 DVDD.n2123 4.5005
R1257 DVDD.n7853 DVDD.n2123 4.5005
R1258 DVDD.n7842 DVDD.n2142 4.5005
R1259 DVDD.n7851 DVDD.n2142 4.5005
R1260 DVDD.n2149 DVDD.n2142 4.5005
R1261 DVDD.n7853 DVDD.n2142 4.5005
R1262 DVDD.n7851 DVDD.n2122 4.5005
R1263 DVDD.n2149 DVDD.n2122 4.5005
R1264 DVDD.n7853 DVDD.n2122 4.5005
R1265 DVDD.n7851 DVDD.n2143 4.5005
R1266 DVDD.n2149 DVDD.n2143 4.5005
R1267 DVDD.n7853 DVDD.n2143 4.5005
R1268 DVDD.n7851 DVDD.n2121 4.5005
R1269 DVDD.n2149 DVDD.n2121 4.5005
R1270 DVDD.n7853 DVDD.n2121 4.5005
R1271 DVDD.n6676 DVDD.n3226 4.5005
R1272 DVDD.n3238 DVDD.n3226 4.5005
R1273 DVDD.n6674 DVDD.n3226 4.5005
R1274 DVDD.n3237 DVDD.n3226 4.5005
R1275 DVDD.n6676 DVDD.n3228 4.5005
R1276 DVDD.n3238 DVDD.n3228 4.5005
R1277 DVDD.n6674 DVDD.n3228 4.5005
R1278 DVDD.n3237 DVDD.n3228 4.5005
R1279 DVDD.n6676 DVDD.n3225 4.5005
R1280 DVDD.n3238 DVDD.n3225 4.5005
R1281 DVDD.n6674 DVDD.n3225 4.5005
R1282 DVDD.n3237 DVDD.n3225 4.5005
R1283 DVDD.n6675 DVDD.n3238 4.5005
R1284 DVDD.n6675 DVDD.n6674 4.5005
R1285 DVDD.n6675 DVDD.n3237 4.5005
R1286 DVDD.n3238 DVDD.n3215 4.5005
R1287 DVDD.n6674 DVDD.n3215 4.5005
R1288 DVDD.n3237 DVDD.n3215 4.5005
R1289 DVDD.n3238 DVDD.n3235 4.5005
R1290 DVDD.n6674 DVDD.n3235 4.5005
R1291 DVDD.n3237 DVDD.n3235 4.5005
R1292 DVDD.n6676 DVDD.n3229 4.5005
R1293 DVDD.n3238 DVDD.n3229 4.5005
R1294 DVDD.n6674 DVDD.n3229 4.5005
R1295 DVDD.n3237 DVDD.n3229 4.5005
R1296 DVDD.n6676 DVDD.n3224 4.5005
R1297 DVDD.n3238 DVDD.n3224 4.5005
R1298 DVDD.n6674 DVDD.n3224 4.5005
R1299 DVDD.n3237 DVDD.n3224 4.5005
R1300 DVDD.n6676 DVDD.n3230 4.5005
R1301 DVDD.n3238 DVDD.n3230 4.5005
R1302 DVDD.n3237 DVDD.n3230 4.5005
R1303 DVDD.n3305 DVDD.n3238 4.5005
R1304 DVDD.n3305 DVDD.n3237 4.5005
R1305 DVDD.n3303 DVDD.n3238 4.5005
R1306 DVDD.n3303 DVDD.n3237 4.5005
R1307 DVDD.n3302 DVDD.n3238 4.5005
R1308 DVDD.n3302 DVDD.n3237 4.5005
R1309 DVDD.n3300 DVDD.n3238 4.5005
R1310 DVDD.n3300 DVDD.n3237 4.5005
R1311 DVDD.n3299 DVDD.n3238 4.5005
R1312 DVDD.n3299 DVDD.n3237 4.5005
R1313 DVDD.n3298 DVDD.n3238 4.5005
R1314 DVDD.n6674 DVDD.n3298 4.5005
R1315 DVDD.n3298 DVDD.n3237 4.5005
R1316 DVDD.n3238 DVDD.n3216 4.5005
R1317 DVDD.n6674 DVDD.n3216 4.5005
R1318 DVDD.n3237 DVDD.n3216 4.5005
R1319 DVDD.n3238 DVDD.n3234 4.5005
R1320 DVDD.n6674 DVDD.n3234 4.5005
R1321 DVDD.n3237 DVDD.n3234 4.5005
R1322 DVDD.n6676 DVDD.n3220 4.5005
R1323 DVDD.n3238 DVDD.n3220 4.5005
R1324 DVDD.n6674 DVDD.n3220 4.5005
R1325 DVDD.n3237 DVDD.n3220 4.5005
R1326 DVDD.n6676 DVDD.n3231 4.5005
R1327 DVDD.n3238 DVDD.n3231 4.5005
R1328 DVDD.n6674 DVDD.n3231 4.5005
R1329 DVDD.n3237 DVDD.n3231 4.5005
R1330 DVDD.n6676 DVDD.n3219 4.5005
R1331 DVDD.n3238 DVDD.n3219 4.5005
R1332 DVDD.n6674 DVDD.n3219 4.5005
R1333 DVDD.n3237 DVDD.n3219 4.5005
R1334 DVDD.n3238 DVDD.n3217 4.5005
R1335 DVDD.n6674 DVDD.n3217 4.5005
R1336 DVDD.n3237 DVDD.n3217 4.5005
R1337 DVDD.n3238 DVDD.n3233 4.5005
R1338 DVDD.n6674 DVDD.n3233 4.5005
R1339 DVDD.n3237 DVDD.n3233 4.5005
R1340 DVDD.n3238 DVDD.n3218 4.5005
R1341 DVDD.n6674 DVDD.n3218 4.5005
R1342 DVDD.n3237 DVDD.n3218 4.5005
R1343 DVDD.n3238 DVDD.n3232 4.5005
R1344 DVDD.n6674 DVDD.n3232 4.5005
R1345 DVDD.n3237 DVDD.n3232 4.5005
R1346 DVDD.n5929 DVDD.n5917 4.5005
R1347 DVDD.n5929 DVDD.n5922 4.5005
R1348 DVDD.n6062 DVDD.n5929 4.5005
R1349 DVDD.n6002 DVDD.n5929 4.5005
R1350 DVDD.n5993 DVDD.n5917 4.5005
R1351 DVDD.n5993 DVDD.n5922 4.5005
R1352 DVDD.n6002 DVDD.n5993 4.5005
R1353 DVDD.n5997 DVDD.n5922 4.5005
R1354 DVDD.n6002 DVDD.n5997 4.5005
R1355 DVDD.n5933 DVDD.n5922 4.5005
R1356 DVDD.n6002 DVDD.n5933 4.5005
R1357 DVDD.n5999 DVDD.n5922 4.5005
R1358 DVDD.n6002 DVDD.n5999 4.5005
R1359 DVDD.n5932 DVDD.n5922 4.5005
R1360 DVDD.n6002 DVDD.n5932 4.5005
R1361 DVDD.n6001 DVDD.n5922 4.5005
R1362 DVDD.n6002 DVDD.n6001 4.5005
R1363 DVDD.n5924 DVDD.n5922 4.5005
R1364 DVDD.n6062 DVDD.n5924 4.5005
R1365 DVDD.n6002 DVDD.n5924 4.5005
R1366 DVDD.n5930 DVDD.n5922 4.5005
R1367 DVDD.n6062 DVDD.n5930 4.5005
R1368 DVDD.n6002 DVDD.n5930 4.5005
R1369 DVDD.n5923 DVDD.n5922 4.5005
R1370 DVDD.n6062 DVDD.n5923 4.5005
R1371 DVDD.n6002 DVDD.n5923 4.5005
R1372 DVDD.n6061 DVDD.n5922 4.5005
R1373 DVDD.n6062 DVDD.n6061 4.5005
R1374 DVDD.n6061 DVDD.n6002 4.5005
R1375 DVDD.n4282 DVDD.n3958 4.5005
R1376 DVDD.n6153 DVDD.n3958 4.5005
R1377 DVDD.n4285 DVDD.n3958 4.5005
R1378 DVDD.n6155 DVDD.n3958 4.5005
R1379 DVDD.n4282 DVDD.n3959 4.5005
R1380 DVDD.n6153 DVDD.n3959 4.5005
R1381 DVDD.n4285 DVDD.n3959 4.5005
R1382 DVDD.n6155 DVDD.n3959 4.5005
R1383 DVDD.n6153 DVDD.n3957 4.5005
R1384 DVDD.n4285 DVDD.n3957 4.5005
R1385 DVDD.n6155 DVDD.n3957 4.5005
R1386 DVDD.n6153 DVDD.n3960 4.5005
R1387 DVDD.n4285 DVDD.n3960 4.5005
R1388 DVDD.n6155 DVDD.n3960 4.5005
R1389 DVDD.n6153 DVDD.n3956 4.5005
R1390 DVDD.n4285 DVDD.n3956 4.5005
R1391 DVDD.n6155 DVDD.n3956 4.5005
R1392 DVDD.n4282 DVDD.n3961 4.5005
R1393 DVDD.n6153 DVDD.n3961 4.5005
R1394 DVDD.n4285 DVDD.n3961 4.5005
R1395 DVDD.n6155 DVDD.n3961 4.5005
R1396 DVDD.n4282 DVDD.n3955 4.5005
R1397 DVDD.n6153 DVDD.n3955 4.5005
R1398 DVDD.n4285 DVDD.n3955 4.5005
R1399 DVDD.n6155 DVDD.n3955 4.5005
R1400 DVDD.n4282 DVDD.n3962 4.5005
R1401 DVDD.n6153 DVDD.n3962 4.5005
R1402 DVDD.n4285 DVDD.n3962 4.5005
R1403 DVDD.n6155 DVDD.n3962 4.5005
R1404 DVDD.n4282 DVDD.n3954 4.5005
R1405 DVDD.n6153 DVDD.n3954 4.5005
R1406 DVDD.n4285 DVDD.n3954 4.5005
R1407 DVDD.n6155 DVDD.n3954 4.5005
R1408 DVDD.n6153 DVDD.n3963 4.5005
R1409 DVDD.n4285 DVDD.n3963 4.5005
R1410 DVDD.n6155 DVDD.n3963 4.5005
R1411 DVDD.n6153 DVDD.n3953 4.5005
R1412 DVDD.n4285 DVDD.n3953 4.5005
R1413 DVDD.n6155 DVDD.n3953 4.5005
R1414 DVDD.n6153 DVDD.n3964 4.5005
R1415 DVDD.n4285 DVDD.n3964 4.5005
R1416 DVDD.n6155 DVDD.n3964 4.5005
R1417 DVDD.n4282 DVDD.n3952 4.5005
R1418 DVDD.n6153 DVDD.n3952 4.5005
R1419 DVDD.n4285 DVDD.n3952 4.5005
R1420 DVDD.n6155 DVDD.n3952 4.5005
R1421 DVDD.n4282 DVDD.n3965 4.5005
R1422 DVDD.n6153 DVDD.n3965 4.5005
R1423 DVDD.n4285 DVDD.n3965 4.5005
R1424 DVDD.n6155 DVDD.n3965 4.5005
R1425 DVDD.n4282 DVDD.n3951 4.5005
R1426 DVDD.n6153 DVDD.n3951 4.5005
R1427 DVDD.n4285 DVDD.n3951 4.5005
R1428 DVDD.n6155 DVDD.n3951 4.5005
R1429 DVDD.n4282 DVDD.n3966 4.5005
R1430 DVDD.n6153 DVDD.n3966 4.5005
R1431 DVDD.n4285 DVDD.n3966 4.5005
R1432 DVDD.n6155 DVDD.n3966 4.5005
R1433 DVDD.n6153 DVDD.n3950 4.5005
R1434 DVDD.n4285 DVDD.n3950 4.5005
R1435 DVDD.n6155 DVDD.n3950 4.5005
R1436 DVDD.n6153 DVDD.n3967 4.5005
R1437 DVDD.n4285 DVDD.n3967 4.5005
R1438 DVDD.n6155 DVDD.n3967 4.5005
R1439 DVDD.n6153 DVDD.n3949 4.5005
R1440 DVDD.n4285 DVDD.n3949 4.5005
R1441 DVDD.n6155 DVDD.n3949 4.5005
R1442 DVDD.n4282 DVDD.n3968 4.5005
R1443 DVDD.n6153 DVDD.n3968 4.5005
R1444 DVDD.n4285 DVDD.n3968 4.5005
R1445 DVDD.n6155 DVDD.n3968 4.5005
R1446 DVDD.n4282 DVDD.n3948 4.5005
R1447 DVDD.n6153 DVDD.n3948 4.5005
R1448 DVDD.n6155 DVDD.n3948 4.5005
R1449 DVDD.n6153 DVDD.n3969 4.5005
R1450 DVDD.n6155 DVDD.n3969 4.5005
R1451 DVDD.n6153 DVDD.n3947 4.5005
R1452 DVDD.n6155 DVDD.n3947 4.5005
R1453 DVDD.n6154 DVDD.n4282 4.5005
R1454 DVDD.n6154 DVDD.n6153 4.5005
R1455 DVDD.n6155 DVDD.n6154 4.5005
R1456 DVDD.n4282 DVDD.n3949 4.5005
R1457 DVDD.n4282 DVDD.n3967 4.5005
R1458 DVDD.n4282 DVDD.n3950 4.5005
R1459 DVDD.n4282 DVDD.n3964 4.5005
R1460 DVDD.n4282 DVDD.n3953 4.5005
R1461 DVDD.n4282 DVDD.n3963 4.5005
R1462 DVDD.n4282 DVDD.n3956 4.5005
R1463 DVDD.n4282 DVDD.n3960 4.5005
R1464 DVDD.n4282 DVDD.n3957 4.5005
R1465 DVDD.n6061 DVDD.n5917 4.5005
R1466 DVDD.n5923 DVDD.n5917 4.5005
R1467 DVDD.n5930 DVDD.n5917 4.5005
R1468 DVDD.n6676 DVDD.n3232 4.5005
R1469 DVDD.n6676 DVDD.n3218 4.5005
R1470 DVDD.n6676 DVDD.n3233 4.5005
R1471 DVDD.n6676 DVDD.n3217 4.5005
R1472 DVDD.n6676 DVDD.n3234 4.5005
R1473 DVDD.n6676 DVDD.n3216 4.5005
R1474 DVDD.n6676 DVDD.n3235 4.5005
R1475 DVDD.n6676 DVDD.n3215 4.5005
R1476 DVDD.n6676 DVDD.n6675 4.5005
R1477 DVDD.n7842 DVDD.n2121 4.5005
R1478 DVDD.n7842 DVDD.n2143 4.5005
R1479 DVDD.n7842 DVDD.n2122 4.5005
R1480 DVDD.n7842 DVDD.n2140 4.5005
R1481 DVDD.n7842 DVDD.n2125 4.5005
R1482 DVDD.n7842 DVDD.n2139 4.5005
R1483 DVDD.n7842 DVDD.n2137 4.5005
R1484 DVDD.n7842 DVDD.n2128 4.5005
R1485 DVDD.n7852 DVDD.n7851 4.5005
R1486 DVDD.n7852 DVDD.n2149 4.5005
R1487 DVDD.n7853 DVDD.n7852 4.5005
R1488 DVDD.n2298 DVDD.n2294 4.5005
R1489 DVDD.n2298 DVDD.n2292 4.5005
R1490 DVDD.n7747 DVDD.n2298 4.5005
R1491 DVDD.n7749 DVDD.n2289 4.5005
R1492 DVDD.n2294 DVDD.n2289 4.5005
R1493 DVDD.n2292 DVDD.n2289 4.5005
R1494 DVDD.n7747 DVDD.n2289 4.5005
R1495 DVDD.n2297 DVDD.n2294 4.5005
R1496 DVDD.n2297 DVDD.n2292 4.5005
R1497 DVDD.n7747 DVDD.n2297 4.5005
R1498 DVDD.n7749 DVDD.n2290 4.5005
R1499 DVDD.n2294 DVDD.n2290 4.5005
R1500 DVDD.n2292 DVDD.n2290 4.5005
R1501 DVDD.n7747 DVDD.n2290 4.5005
R1502 DVDD.n2296 DVDD.n2294 4.5005
R1503 DVDD.n2296 DVDD.n2292 4.5005
R1504 DVDD.n7747 DVDD.n2296 4.5005
R1505 DVDD.n7749 DVDD.n7748 4.5005
R1506 DVDD.n7748 DVDD.n2294 4.5005
R1507 DVDD.n7748 DVDD.n2292 4.5005
R1508 DVDD.n7748 DVDD.n7747 4.5005
R1509 DVDD.n8291 DVDD.n1678 4.5005
R1510 DVDD.n8291 DVDD.n8290 4.5005
R1511 DVDD.n8291 DVDD.n1660 4.5005
R1512 DVDD.n8292 DVDD.n8291 4.5005
R1513 DVDD.n1878 DVDD.n1677 4.5005
R1514 DVDD.n1882 DVDD.n1677 4.5005
R1515 DVDD.n1879 DVDD.n1679 4.5005
R1516 DVDD.n7666 DVDD.n2291 4.5005
R1517 DVDD.n7671 DVDD.n2293 4.5005
R1518 DVDD.n2436 DVDD.n2435 4.5005
R1519 DVDD.n2440 DVDD.n2439 4.5005
R1520 DVDD.n2413 DVDD.n2412 4.5005
R1521 DVDD.n2417 DVDD.n2416 4.5005
R1522 DVDD.n3249 DVDD.n3248 4.5005
R1523 DVDD.n3247 DVDD.n3246 4.5005
R1524 DVDD.n3245 DVDD.n3244 4.5005
R1525 DVDD.n3243 DVDD.n3242 4.5005
R1526 DVDD.n3240 DVDD.n3236 4.5005
R1527 DVDD.n3296 DVDD.n3295 4.5005
R1528 DVDD.n3294 DVDD.n3239 4.5005
R1529 DVDD.n3293 DVDD.n3292 4.5005
R1530 DVDD.n3291 DVDD.n3290 4.5005
R1531 DVDD.n3289 DVDD.n3288 4.5005
R1532 DVDD.n3287 DVDD.n3241 4.5005
R1533 DVDD.n3286 DVDD.n3285 4.5005
R1534 DVDD.n3284 DVDD.n3283 4.5005
R1535 DVDD.n3282 DVDD.n3281 4.5005
R1536 DVDD.n3280 DVDD.n3279 4.5005
R1537 DVDD.n3278 DVDD.n3277 4.5005
R1538 DVDD.n3276 DVDD.n3275 4.5005
R1539 DVDD.n3274 DVDD.n3273 4.5005
R1540 DVDD.n3272 DVDD.n3271 4.5005
R1541 DVDD.n3270 DVDD.n3269 4.5005
R1542 DVDD.n3268 DVDD.n3267 4.5005
R1543 DVDD.n3266 DVDD.n3265 4.5005
R1544 DVDD.n3264 DVDD.n3263 4.5005
R1545 DVDD.n3262 DVDD.n3261 4.5005
R1546 DVDD.n3260 DVDD.n3259 4.5005
R1547 DVDD.n3258 DVDD.n3257 4.5005
R1548 DVDD.n3256 DVDD.n3255 4.5005
R1549 DVDD.n3254 DVDD.n3253 4.5005
R1550 DVDD.n3252 DVDD.n3251 4.5005
R1551 DVDD.n5992 DVDD.n5991 4.5005
R1552 DVDD.n5990 DVDD.n5989 4.5005
R1553 DVDD.n5988 DVDD.n5934 4.5005
R1554 DVDD.n5987 DVDD.n5986 4.5005
R1555 DVDD.n5985 DVDD.n5935 4.5005
R1556 DVDD.n5984 DVDD.n5983 4.5005
R1557 DVDD.n5982 DVDD.n5936 4.5005
R1558 DVDD.n5981 DVDD.n5980 4.5005
R1559 DVDD.n5979 DVDD.n5937 4.5005
R1560 DVDD.n5978 DVDD.n5977 4.5005
R1561 DVDD.n5976 DVDD.n5938 4.5005
R1562 DVDD.n5975 DVDD.n5974 4.5005
R1563 DVDD.n5973 DVDD.n5939 4.5005
R1564 DVDD.n5972 DVDD.n5971 4.5005
R1565 DVDD.n5970 DVDD.n5940 4.5005
R1566 DVDD.n5969 DVDD.n5968 4.5005
R1567 DVDD.n5967 DVDD.n5941 4.5005
R1568 DVDD.n5966 DVDD.n5965 4.5005
R1569 DVDD.n5964 DVDD.n5963 4.5005
R1570 DVDD.n5962 DVDD.n5961 4.5005
R1571 DVDD.n5960 DVDD.n5959 4.5005
R1572 DVDD.n5958 DVDD.n5957 4.5005
R1573 DVDD.n5956 DVDD.n5955 4.5005
R1574 DVDD.n5954 DVDD.n5953 4.5005
R1575 DVDD.n5952 DVDD.n5951 4.5005
R1576 DVDD.n5950 DVDD.n5949 4.5005
R1577 DVDD.n5948 DVDD.n5947 4.5005
R1578 DVDD.n5946 DVDD.n5945 4.5005
R1579 DVDD.n5944 DVDD.n5943 4.5005
R1580 DVDD.n6053 DVDD.n6052 4.5005
R1581 DVDD.n6051 DVDD.n6050 4.5005
R1582 DVDD.n6049 DVDD.n6048 4.5005
R1583 DVDD.n6047 DVDD.n6046 4.5005
R1584 DVDD.n6045 DVDD.n6044 4.5005
R1585 DVDD.n6043 DVDD.n6042 4.5005
R1586 DVDD.n6041 DVDD.n6040 4.5005
R1587 DVDD.n6039 DVDD.n6038 4.5005
R1588 DVDD.n6037 DVDD.n6036 4.5005
R1589 DVDD.n6035 DVDD.n6034 4.5005
R1590 DVDD.n6033 DVDD.n6032 4.5005
R1591 DVDD.n6031 DVDD.n6030 4.5005
R1592 DVDD.n6029 DVDD.n6028 4.5005
R1593 DVDD.n6027 DVDD.n6026 4.5005
R1594 DVDD.n6025 DVDD.n6024 4.5005
R1595 DVDD.n6023 DVDD.n6022 4.5005
R1596 DVDD.n6021 DVDD.n6020 4.5005
R1597 DVDD.n6019 DVDD.n6018 4.5005
R1598 DVDD.n6017 DVDD.n6016 4.5005
R1599 DVDD.n6015 DVDD.n6014 4.5005
R1600 DVDD.n6013 DVDD.n6012 4.5005
R1601 DVDD.n6011 DVDD.n6010 4.5005
R1602 DVDD.n6009 DVDD.n6008 4.5005
R1603 DVDD.n6007 DVDD.n6006 4.5005
R1604 DVDD.n6005 DVDD.n6004 4.5005
R1605 DVDD.n6003 DVDD.n5931 4.5005
R1606 DVDD.n6060 DVDD.n6059 4.5005
R1607 DVDD.n6058 DVDD.n6057 4.5005
R1608 DVDD.n6056 DVDD.n6055 4.5005
R1609 DVDD.n4276 DVDD.n4275 4.5005
R1610 DVDD.n4274 DVDD.n3972 4.5005
R1611 DVDD.n4273 DVDD.n4272 4.5005
R1612 DVDD.n4271 DVDD.n4224 4.5005
R1613 DVDD.n4270 DVDD.n4269 4.5005
R1614 DVDD.n4268 DVDD.n4225 4.5005
R1615 DVDD.n4267 DVDD.n4266 4.5005
R1616 DVDD.n4265 DVDD.n4226 4.5005
R1617 DVDD.n4264 DVDD.n4263 4.5005
R1618 DVDD.n4262 DVDD.n4227 4.5005
R1619 DVDD.n4261 DVDD.n4260 4.5005
R1620 DVDD.n4259 DVDD.n4228 4.5005
R1621 DVDD.n4258 DVDD.n4257 4.5005
R1622 DVDD.n4256 DVDD.n4229 4.5005
R1623 DVDD.n4255 DVDD.n4254 4.5005
R1624 DVDD.n4253 DVDD.n4230 4.5005
R1625 DVDD.n4252 DVDD.n4251 4.5005
R1626 DVDD.n4250 DVDD.n4231 4.5005
R1627 DVDD.n4249 DVDD.n4248 4.5005
R1628 DVDD.n4247 DVDD.n4232 4.5005
R1629 DVDD.n4246 DVDD.n4245 4.5005
R1630 DVDD.n4244 DVDD.n4233 4.5005
R1631 DVDD.n4243 DVDD.n4242 4.5005
R1632 DVDD.n4241 DVDD.n4234 4.5005
R1633 DVDD.n4240 DVDD.n4239 4.5005
R1634 DVDD.n4238 DVDD.n4235 4.5005
R1635 DVDD.n4237 DVDD.n4236 4.5005
R1636 DVDD.n3971 DVDD.n3970 4.5005
R1637 DVDD.n4279 DVDD.n4278 4.5005
R1638 DVDD.n4220 DVDD.n4219 4.5005
R1639 DVDD.n4217 DVDD.n3975 4.5005
R1640 DVDD.n4156 DVDD.n4147 4.5005
R1641 DVDD.n4159 DVDD.n4157 4.5005
R1642 DVDD.n4162 DVDD.n4161 4.5005
R1643 DVDD.n4163 DVDD.n4154 4.5005
R1644 DVDD.n4205 DVDD.n4204 4.5005
R1645 DVDD.n4203 DVDD.n4202 4.5005
R1646 DVDD.n4201 DVDD.n4164 4.5005
R1647 DVDD.n4200 DVDD.n4199 4.5005
R1648 DVDD.n4198 DVDD.n4165 4.5005
R1649 DVDD.n4197 DVDD.n4196 4.5005
R1650 DVDD.n4195 DVDD.n4166 4.5005
R1651 DVDD.n4194 DVDD.n4193 4.5005
R1652 DVDD.n4192 DVDD.n4167 4.5005
R1653 DVDD.n4191 DVDD.n4190 4.5005
R1654 DVDD.n4189 DVDD.n4168 4.5005
R1655 DVDD.n4188 DVDD.n4187 4.5005
R1656 DVDD.n4186 DVDD.n4169 4.5005
R1657 DVDD.n4185 DVDD.n4184 4.5005
R1658 DVDD.n4183 DVDD.n4170 4.5005
R1659 DVDD.n4182 DVDD.n4181 4.5005
R1660 DVDD.n4180 DVDD.n4171 4.5005
R1661 DVDD.n4179 DVDD.n4178 4.5005
R1662 DVDD.n4177 DVDD.n4172 4.5005
R1663 DVDD.n4176 DVDD.n4175 4.5005
R1664 DVDD.n4174 DVDD.n4173 4.5005
R1665 DVDD.n3974 DVDD.n3973 4.5005
R1666 DVDD.n4223 DVDD.n4222 4.5005
R1667 DVDD.n4115 DVDD.n4114 4.5005
R1668 DVDD.n4113 DVDD.n3996 4.5005
R1669 DVDD.n4005 DVDD.n3997 4.5005
R1670 DVDD.n4007 DVDD.n4006 4.5005
R1671 DVDD.n4008 DVDD.n4003 4.5005
R1672 DVDD.n4013 DVDD.n4012 4.5005
R1673 DVDD.n4014 DVDD.n4002 4.5005
R1674 DVDD.n4100 DVDD.n4099 4.5005
R1675 DVDD.n4098 DVDD.n4097 4.5005
R1676 DVDD.n4016 DVDD.n4015 4.5005
R1677 DVDD.n4038 DVDD.n4037 4.5005
R1678 DVDD.n4040 DVDD.n4039 4.5005
R1679 DVDD.n4044 DVDD.n4035 4.5005
R1680 DVDD.n4049 DVDD.n4048 4.5005
R1681 DVDD.n4051 DVDD.n4050 4.5005
R1682 DVDD.n4052 DVDD.n4033 4.5005
R1683 DVDD.n4054 DVDD.n4053 4.5005
R1684 DVDD.n4057 DVDD.n4056 4.5005
R1685 DVDD.n4055 DVDD.n4030 4.5005
R1686 DVDD.n4063 DVDD.n4029 4.5005
R1687 DVDD.n4066 DVDD.n4065 4.5005
R1688 DVDD.n4067 DVDD.n4028 4.5005
R1689 DVDD.n4077 DVDD.n4076 4.5005
R1690 DVDD.n4075 DVDD.n4074 4.5005
R1691 DVDD.n4070 DVDD.n4068 4.5005
R1692 DVDD.n3995 DVDD.n3993 4.5005
R1693 DVDD.n4121 DVDD.n4120 4.5005
R1694 DVDD.n4119 DVDD.n4118 4.5005
R1695 DVDD.n4117 DVDD.n3984 4.5005
R1696 DVDD.n9107 DVDD.n9106 4.5005
R1697 DVDD.n9105 DVDD.n541 4.5005
R1698 DVDD.n9104 DVDD.n9103 4.5005
R1699 DVDD.n9102 DVDD.n9075 4.5005
R1700 DVDD.n9101 DVDD.n9100 4.5005
R1701 DVDD.n9099 DVDD.n9076 4.5005
R1702 DVDD.n9098 DVDD.n9097 4.5005
R1703 DVDD.n9096 DVDD.n9077 4.5005
R1704 DVDD.n9095 DVDD.n9094 4.5005
R1705 DVDD.n9093 DVDD.n9092 4.5005
R1706 DVDD.n9091 DVDD.n9090 4.5005
R1707 DVDD.n9089 DVDD.n9088 4.5005
R1708 DVDD.n9087 DVDD.n9086 4.5005
R1709 DVDD.n9085 DVDD.n9084 4.5005
R1710 DVDD.n9083 DVDD.n9082 4.5005
R1711 DVDD.n9081 DVDD.n9080 4.5005
R1712 DVDD.n9079 DVDD.n9078 4.5005
R1713 DVDD.n536 DVDD.n532 4.5005
R1714 DVDD.n9125 DVDD.n9124 4.5005
R1715 DVDD.n9123 DVDD.n535 4.5005
R1716 DVDD.n9122 DVDD.n9121 4.5005
R1717 DVDD.n9120 DVDD.n9119 4.5005
R1718 DVDD.n9118 DVDD.n537 4.5005
R1719 DVDD.n9117 DVDD.n9116 4.5005
R1720 DVDD.n9115 DVDD.n538 4.5005
R1721 DVDD.n9114 DVDD.n9113 4.5005
R1722 DVDD.n9112 DVDD.n539 4.5005
R1723 DVDD.n9111 DVDD.n9110 4.5005
R1724 DVDD.n9109 DVDD.n540 4.5005
R1725 DVDD.n9071 DVDD.n9070 4.5005
R1726 DVDD.n9069 DVDD.n544 4.5005
R1727 DVDD.n9068 DVDD.n9067 4.5005
R1728 DVDD.n9066 DVDD.n9019 4.5005
R1729 DVDD.n9065 DVDD.n9064 4.5005
R1730 DVDD.n9063 DVDD.n9020 4.5005
R1731 DVDD.n9062 DVDD.n9061 4.5005
R1732 DVDD.n9060 DVDD.n9021 4.5005
R1733 DVDD.n9059 DVDD.n9058 4.5005
R1734 DVDD.n9057 DVDD.n9022 4.5005
R1735 DVDD.n9056 DVDD.n9055 4.5005
R1736 DVDD.n9054 DVDD.n9023 4.5005
R1737 DVDD.n9053 DVDD.n9052 4.5005
R1738 DVDD.n9051 DVDD.n9024 4.5005
R1739 DVDD.n9050 DVDD.n9049 4.5005
R1740 DVDD.n9048 DVDD.n9025 4.5005
R1741 DVDD.n9047 DVDD.n9046 4.5005
R1742 DVDD.n9045 DVDD.n9026 4.5005
R1743 DVDD.n9044 DVDD.n9043 4.5005
R1744 DVDD.n9042 DVDD.n9027 4.5005
R1745 DVDD.n9041 DVDD.n9040 4.5005
R1746 DVDD.n9039 DVDD.n9028 4.5005
R1747 DVDD.n9038 DVDD.n9037 4.5005
R1748 DVDD.n9036 DVDD.n9029 4.5005
R1749 DVDD.n9035 DVDD.n9034 4.5005
R1750 DVDD.n9033 DVDD.n9030 4.5005
R1751 DVDD.n9032 DVDD.n9031 4.5005
R1752 DVDD.n543 DVDD.n542 4.5005
R1753 DVDD.n9074 DVDD.n9073 4.5005
R1754 DVDD.n550 DVDD.n547 4.5005
R1755 DVDD.n8978 DVDD.n8977 4.5005
R1756 DVDD.n8980 DVDD.n8979 4.5005
R1757 DVDD.n8982 DVDD.n8981 4.5005
R1758 DVDD.n8984 DVDD.n8983 4.5005
R1759 DVDD.n8986 DVDD.n8985 4.5005
R1760 DVDD.n8988 DVDD.n8987 4.5005
R1761 DVDD.n8989 DVDD.n8976 4.5005
R1762 DVDD.n9011 DVDD.n9010 4.5005
R1763 DVDD.n9009 DVDD.n9008 4.5005
R1764 DVDD.n9007 DVDD.n9006 4.5005
R1765 DVDD.n9005 DVDD.n9004 4.5005
R1766 DVDD.n9003 DVDD.n9002 4.5005
R1767 DVDD.n9001 DVDD.n8990 4.5005
R1768 DVDD.n9000 DVDD.n8999 4.5005
R1769 DVDD.n8998 DVDD.n8991 4.5005
R1770 DVDD.n8997 DVDD.n8996 4.5005
R1771 DVDD.n8995 DVDD.n8992 4.5005
R1772 DVDD.n8994 DVDD.n8993 4.5005
R1773 DVDD.n546 DVDD.n545 4.5005
R1774 DVDD.n9018 DVDD.n9017 4.5005
R1775 DVDD.n8520 DVDD.n1369 4.5005
R1776 DVDD.n8539 DVDD.n1369 4.5005
R1777 DVDD.n8541 DVDD.n8540 4.5005
R1778 DVDD.n8540 DVDD.n8539 4.5005
R1779 DVDD.n1455 DVDD.n1334 4.5005
R1780 DVDD.n8435 DVDD.n1334 4.5005
R1781 DVDD.n1332 DVDD.n1330 4.5005
R1782 DVDD.n8623 DVDD.n1330 4.5005
R1783 DVDD.n8622 DVDD.n8621 4.5005
R1784 DVDD.n8623 DVDD.n8622 4.5005
R1785 DVDD.n8435 DVDD.n8434 4.5005
R1786 DVDD.n8434 DVDD.n1455 4.5005
R1787 DVDD.n8434 DVDD.n8433 4.5005
R1788 DVDD.n1455 DVDD.n1424 4.5005
R1789 DVDD.n8433 DVDD.n1424 4.5005
R1790 DVDD.n8499 DVDD.n1426 4.5005
R1791 DVDD.n8499 DVDD.n8498 4.5005
R1792 DVDD.n8498 DVDD.n1421 4.5005
R1793 DVDD.n1426 DVDD.n1421 4.5005
R1794 DVDD.n8501 DVDD.n1421 4.5005
R1795 DVDD.n1426 DVDD.n1363 4.5005
R1796 DVDD.n8501 DVDD.n1363 4.5005
R1797 DVDD.n8595 DVDD.n8594 4.5005
R1798 DVDD.n8596 DVDD.n8595 4.5005
R1799 DVDD.n8596 DVDD.n1362 4.5005
R1800 DVDD.n8594 DVDD.n1362 4.5005
R1801 DVDD.n8592 DVDD.n1362 4.5005
R1802 DVDD.n8594 DVDD.n8593 4.5005
R1803 DVDD.n8593 DVDD.n8592 4.5005
R1804 DVDD.n7733 DVDD.n7732 4.5005
R1805 DVDD.n7734 DVDD.n7733 4.5005
R1806 DVDD.n7743 DVDD.n7742 4.5005
R1807 DVDD.n7736 DVDD.n2336 4.5005
R1808 DVDD.n7732 DVDD.n2336 4.5005
R1809 DVDD.n7734 DVDD.n2336 4.5005
R1810 DVDD.n7743 DVDD.n2150 4.5005
R1811 DVDD.n2334 DVDD.n2150 4.5005
R1812 DVDD.n7740 DVDD.n2150 4.5005
R1813 DVDD.n7737 DVDD.n2150 4.5005
R1814 DVDD.n7736 DVDD.n7735 4.5005
R1815 DVDD.n7735 DVDD.n7734 4.5005
R1816 DVDD.n7723 DVDD.n7722 4.5005
R1817 DVDD.n7716 DVDD.n2341 4.5005
R1818 DVDD.n7725 DVDD.n7703 4.5005
R1819 DVDD.n7720 DVDD.n7710 4.5005
R1820 DVDD.n7725 DVDD.n7724 4.5005
R1821 DVDD.n7724 DVDD.n7706 4.5005
R1822 DVDD.n7724 DVDD.n7708 4.5005
R1823 DVDD.n7724 DVDD.n7705 4.5005
R1824 DVDD.n7724 DVDD.n7723 4.5005
R1825 DVDD.n7720 DVDD.n7719 4.5005
R1826 DVDD.n7719 DVDD.n7714 4.5005
R1827 DVDD.n7719 DVDD.n7718 4.5005
R1828 DVDD.n7719 DVDD.n7713 4.5005
R1829 DVDD.n7719 DVDD.n2341 4.5005
R1830 DVDD.n7696 DVDD.n2345 4.5005
R1831 DVDD.n2348 DVDD.n2345 4.5005
R1832 DVDD.n7702 DVDD.n2345 4.5005
R1833 DVDD.n7697 DVDD.n7696 4.5005
R1834 DVDD.n7701 DVDD.n7700 4.5005
R1835 DVDD.n7701 DVDD.n2346 4.5005
R1836 DVDD.n7702 DVDD.n7701 4.5005
R1837 DVDD.n1875 DVDD.n1874 4.5005
R1838 DVDD.n1872 DVDD.n1871 4.5005
R1839 DVDD.n7673 DVDD.n7672 4.5005
R1840 DVDD.n7675 DVDD.n2246 4.5005
R1841 DVDD.n2442 DVDD.n2441 4.5005
R1842 DVDD.n2446 DVDD.n2445 4.5005
R1843 DVDD.n2419 DVDD.n2418 4.5005
R1844 DVDD.n2423 DVDD.n2422 4.5005
R1845 DVDD.n2367 DVDD.n2366 4.5005
R1846 DVDD.n2368 DVDD.n2367 4.5005
R1847 DVDD.n2370 DVDD.n2359 4.5005
R1848 DVDD.n2366 DVDD.n2359 4.5005
R1849 DVDD.n2368 DVDD.n2359 4.5005
R1850 DVDD.n2370 DVDD.n2369 4.5005
R1851 DVDD.n2369 DVDD.n2368 4.5005
R1852 DVDD.n3140 DVDD.n3139 4.5005
R1853 DVDD.n3143 DVDD.n3142 4.5005
R1854 DVDD.n3145 DVDD.n3144 4.5005
R1855 DVDD.n3147 DVDD.n3146 4.5005
R1856 DVDD.n3149 DVDD.n3148 4.5005
R1857 DVDD.n3151 DVDD.n3150 4.5005
R1858 DVDD.n3153 DVDD.n3152 4.5005
R1859 DVDD.n3155 DVDD.n3154 4.5005
R1860 DVDD.n3157 DVDD.n3156 4.5005
R1861 DVDD.n3159 DVDD.n3158 4.5005
R1862 DVDD.n3161 DVDD.n3160 4.5005
R1863 DVDD.n3163 DVDD.n3162 4.5005
R1864 DVDD.n3165 DVDD.n3164 4.5005
R1865 DVDD.n3167 DVDD.n3166 4.5005
R1866 DVDD.n3169 DVDD.n3168 4.5005
R1867 DVDD.n3171 DVDD.n3170 4.5005
R1868 DVDD.n3173 DVDD.n3172 4.5005
R1869 DVDD.n3175 DVDD.n3174 4.5005
R1870 DVDD.n3177 DVDD.n3176 4.5005
R1871 DVDD.n3178 DVDD.n3123 4.5005
R1872 DVDD.n3180 DVDD.n3179 4.5005
R1873 DVDD.n3124 DVDD.n3121 4.5005
R1874 DVDD.n3126 DVDD.n3125 4.5005
R1875 DVDD.n3128 DVDD.n3127 4.5005
R1876 DVDD.n3130 DVDD.n3129 4.5005
R1877 DVDD.n3132 DVDD.n3131 4.5005
R1878 DVDD.n3134 DVDD.n3133 4.5005
R1879 DVDD.n3136 DVDD.n3135 4.5005
R1880 DVDD.n3138 DVDD.n3137 4.5005
R1881 DVDD.n5831 DVDD.n5828 4.5005
R1882 DVDD.n5842 DVDD.n5841 4.5005
R1883 DVDD.n5844 DVDD.n5843 4.5005
R1884 DVDD.n5846 DVDD.n5845 4.5005
R1885 DVDD.n5848 DVDD.n5847 4.5005
R1886 DVDD.n5850 DVDD.n5849 4.5005
R1887 DVDD.n5852 DVDD.n5851 4.5005
R1888 DVDD.n5854 DVDD.n5853 4.5005
R1889 DVDD.n5856 DVDD.n5855 4.5005
R1890 DVDD.n5858 DVDD.n5857 4.5005
R1891 DVDD.n5860 DVDD.n5859 4.5005
R1892 DVDD.n5861 DVDD.n5839 4.5005
R1893 DVDD.n5863 DVDD.n5862 4.5005
R1894 DVDD.n5864 DVDD.n5838 4.5005
R1895 DVDD.n5866 DVDD.n5865 4.5005
R1896 DVDD.n5867 DVDD.n5837 4.5005
R1897 DVDD.n5869 DVDD.n5868 4.5005
R1898 DVDD.n5870 DVDD.n5836 4.5005
R1899 DVDD.n5872 DVDD.n5871 4.5005
R1900 DVDD.n5873 DVDD.n5835 4.5005
R1901 DVDD.n5875 DVDD.n5874 4.5005
R1902 DVDD.n5876 DVDD.n5834 4.5005
R1903 DVDD.n5878 DVDD.n5877 4.5005
R1904 DVDD.n5879 DVDD.n5833 4.5005
R1905 DVDD.n5881 DVDD.n5880 4.5005
R1906 DVDD.n5882 DVDD.n5832 4.5005
R1907 DVDD.n5884 DVDD.n5883 4.5005
R1908 DVDD.n5885 DVDD.n5830 4.5005
R1909 DVDD.n5887 DVDD.n5886 4.5005
R1910 DVDD.n5820 DVDD.n5819 4.5005
R1911 DVDD.n5823 DVDD.n5822 4.5005
R1912 DVDD.n5768 DVDD.n5767 4.5005
R1913 DVDD.n5770 DVDD.n5769 4.5005
R1914 DVDD.n5772 DVDD.n5771 4.5005
R1915 DVDD.n5774 DVDD.n5773 4.5005
R1916 DVDD.n5775 DVDD.n4389 4.5005
R1917 DVDD.n5776 DVDD.n4387 4.5005
R1918 DVDD.n5778 DVDD.n5777 4.5005
R1919 DVDD.n5780 DVDD.n5779 4.5005
R1920 DVDD.n5782 DVDD.n5781 4.5005
R1921 DVDD.n5784 DVDD.n5783 4.5005
R1922 DVDD.n5786 DVDD.n5785 4.5005
R1923 DVDD.n5788 DVDD.n5787 4.5005
R1924 DVDD.n5790 DVDD.n5789 4.5005
R1925 DVDD.n5792 DVDD.n5791 4.5005
R1926 DVDD.n5794 DVDD.n5793 4.5005
R1927 DVDD.n5796 DVDD.n5795 4.5005
R1928 DVDD.n5798 DVDD.n5797 4.5005
R1929 DVDD.n5800 DVDD.n5799 4.5005
R1930 DVDD.n5802 DVDD.n5801 4.5005
R1931 DVDD.n5804 DVDD.n5803 4.5005
R1932 DVDD.n5806 DVDD.n5805 4.5005
R1933 DVDD.n5808 DVDD.n5807 4.5005
R1934 DVDD.n5810 DVDD.n5809 4.5005
R1935 DVDD.n5812 DVDD.n5811 4.5005
R1936 DVDD.n5814 DVDD.n5813 4.5005
R1937 DVDD.n5816 DVDD.n5815 4.5005
R1938 DVDD.n5818 DVDD.n5817 4.5005
R1939 DVDD.n4372 DVDD.n4371 4.5005
R1940 DVDD.n4375 DVDD.n4374 4.5005
R1941 DVDD.n4318 DVDD.n4317 4.5005
R1942 DVDD.n4333 DVDD.n4332 4.5005
R1943 DVDD.n4334 DVDD.n4331 4.5005
R1944 DVDD.n4336 DVDD.n4335 4.5005
R1945 DVDD.n4337 DVDD.n4330 4.5005
R1946 DVDD.n4339 DVDD.n4338 4.5005
R1947 DVDD.n4340 DVDD.n4329 4.5005
R1948 DVDD.n4342 DVDD.n4341 4.5005
R1949 DVDD.n4343 DVDD.n4328 4.5005
R1950 DVDD.n4345 DVDD.n4344 4.5005
R1951 DVDD.n4346 DVDD.n4327 4.5005
R1952 DVDD.n4348 DVDD.n4347 4.5005
R1953 DVDD.n4349 DVDD.n4326 4.5005
R1954 DVDD.n4351 DVDD.n4350 4.5005
R1955 DVDD.n4352 DVDD.n4325 4.5005
R1956 DVDD.n4354 DVDD.n4353 4.5005
R1957 DVDD.n4355 DVDD.n4324 4.5005
R1958 DVDD.n4357 DVDD.n4356 4.5005
R1959 DVDD.n4358 DVDD.n4323 4.5005
R1960 DVDD.n4360 DVDD.n4359 4.5005
R1961 DVDD.n4361 DVDD.n4322 4.5005
R1962 DVDD.n4363 DVDD.n4362 4.5005
R1963 DVDD.n4364 DVDD.n4321 4.5005
R1964 DVDD.n4366 DVDD.n4365 4.5005
R1965 DVDD.n4367 DVDD.n4320 4.5005
R1966 DVDD.n4369 DVDD.n4368 4.5005
R1967 DVDD.n4370 DVDD.n4319 4.5005
R1968 DVDD.n9511 DVDD.n9510 4.5005
R1969 DVDD.n9513 DVDD.n265 4.5005
R1970 DVDD.n9515 DVDD.n9514 4.5005
R1971 DVDD.n9516 DVDD.n264 4.5005
R1972 DVDD.n9518 DVDD.n9517 4.5005
R1973 DVDD.n9519 DVDD.n263 4.5005
R1974 DVDD.n9521 DVDD.n9520 4.5005
R1975 DVDD.n9522 DVDD.n262 4.5005
R1976 DVDD.n9524 DVDD.n9523 4.5005
R1977 DVDD.n9525 DVDD.n261 4.5005
R1978 DVDD.n9527 DVDD.n9526 4.5005
R1979 DVDD.n9528 DVDD.n260 4.5005
R1980 DVDD.n9530 DVDD.n9529 4.5005
R1981 DVDD.n9531 DVDD.n259 4.5005
R1982 DVDD.n9533 DVDD.n9532 4.5005
R1983 DVDD.n9534 DVDD.n258 4.5005
R1984 DVDD.n9536 DVDD.n9535 4.5005
R1985 DVDD.n9537 DVDD.n257 4.5005
R1986 DVDD.n9539 DVDD.n9538 4.5005
R1987 DVDD.n9540 DVDD.n256 4.5005
R1988 DVDD.n9542 DVDD.n9541 4.5005
R1989 DVDD.n9543 DVDD.n255 4.5005
R1990 DVDD.n9545 DVDD.n9544 4.5005
R1991 DVDD.n250 DVDD.n248 4.5005
R1992 DVDD.n9551 DVDD.n9550 4.5005
R1993 DVDD.n9552 DVDD.n246 4.5005
R1994 DVDD.n9554 DVDD.n9553 4.5005
R1995 DVDD.n247 DVDD.n245 4.5005
R1996 DVDD.n9508 DVDD.n266 4.5005
R1997 DVDD.n9475 DVDD.n9474 4.5005
R1998 DVDD.n9477 DVDD.n275 4.5005
R1999 DVDD.n9479 DVDD.n9478 4.5005
R2000 DVDD.n9481 DVDD.n9480 4.5005
R2001 DVDD.n285 DVDD.n283 4.5005
R2002 DVDD.n367 DVDD.n366 4.5005
R2003 DVDD.n369 DVDD.n368 4.5005
R2004 DVDD.n345 DVDD.n343 4.5005
R2005 DVDD.n9434 DVDD.n9433 4.5005
R2006 DVDD.n9435 DVDD.n332 4.5005
R2007 DVDD.n9437 DVDD.n9436 4.5005
R2008 DVDD.n342 DVDD.n331 4.5005
R2009 DVDD.n341 DVDD.n340 4.5005
R2010 DVDD.n336 DVDD.n333 4.5005
R2011 DVDD.n335 DVDD.n334 4.5005
R2012 DVDD.n321 DVDD.n320 4.5005
R2013 DVDD.n9448 DVDD.n9447 4.5005
R2014 DVDD.n9450 DVDD.n9449 4.5005
R2015 DVDD.n319 DVDD.n314 4.5005
R2016 DVDD.n318 DVDD.n317 4.5005
R2017 DVDD.n307 DVDD.n306 4.5005
R2018 DVDD.n9460 DVDD.n9459 4.5005
R2019 DVDD.n9462 DVDD.n9461 4.5005
R2020 DVDD.n9464 DVDD.n9463 4.5005
R2021 DVDD.n305 DVDD.n295 4.5005
R2022 DVDD.n304 DVDD.n303 4.5005
R2023 DVDD.n301 DVDD.n299 4.5005
R2024 DVDD.n298 DVDD.n288 4.5005
R2025 DVDD.n9473 DVDD.n286 4.5005
R2026 DVDD.n4950 DVDD.n4949 4.5005
R2027 DVDD.n4902 DVDD.n287 4.5005
R2028 DVDD.n4904 DVDD.n4903 4.5005
R2029 DVDD.n4906 DVDD.n4905 4.5005
R2030 DVDD.n4907 DVDD.n4900 4.5005
R2031 DVDD.n4909 DVDD.n4908 4.5005
R2032 DVDD.n4910 DVDD.n4899 4.5005
R2033 DVDD.n4912 DVDD.n4911 4.5005
R2034 DVDD.n4913 DVDD.n497 4.5005
R2035 DVDD.n4914 DVDD.n495 4.5005
R2036 DVDD.n4916 DVDD.n4915 4.5005
R2037 DVDD.n4918 DVDD.n4917 4.5005
R2038 DVDD.n4920 DVDD.n4919 4.5005
R2039 DVDD.n4922 DVDD.n4921 4.5005
R2040 DVDD.n4924 DVDD.n4923 4.5005
R2041 DVDD.n4926 DVDD.n4925 4.5005
R2042 DVDD.n4928 DVDD.n4927 4.5005
R2043 DVDD.n4930 DVDD.n4929 4.5005
R2044 DVDD.n4932 DVDD.n4931 4.5005
R2045 DVDD.n4934 DVDD.n4933 4.5005
R2046 DVDD.n4936 DVDD.n4935 4.5005
R2047 DVDD.n4938 DVDD.n4937 4.5005
R2048 DVDD.n4939 DVDD.n4898 4.5005
R2049 DVDD.n4941 DVDD.n4940 4.5005
R2050 DVDD.n4942 DVDD.n4897 4.5005
R2051 DVDD.n4944 DVDD.n4943 4.5005
R2052 DVDD.n4945 DVDD.n4896 4.5005
R2053 DVDD.n4947 DVDD.n4946 4.5005
R2054 DVDD.n4948 DVDD.n4895 4.5005
R2055 DVDD.n4995 DVDD.n4994 4.5005
R2056 DVDD.n4953 DVDD.n4952 4.5005
R2057 DVDD.n4954 DVDD.n4894 4.5005
R2058 DVDD.n4956 DVDD.n4955 4.5005
R2059 DVDD.n4957 DVDD.n4893 4.5005
R2060 DVDD.n4959 DVDD.n4958 4.5005
R2061 DVDD.n4960 DVDD.n4892 4.5005
R2062 DVDD.n4962 DVDD.n4961 4.5005
R2063 DVDD.n4963 DVDD.n4891 4.5005
R2064 DVDD.n4965 DVDD.n4964 4.5005
R2065 DVDD.n4966 DVDD.n4890 4.5005
R2066 DVDD.n4968 DVDD.n4967 4.5005
R2067 DVDD.n4969 DVDD.n4889 4.5005
R2068 DVDD.n4971 DVDD.n4970 4.5005
R2069 DVDD.n4972 DVDD.n4888 4.5005
R2070 DVDD.n4974 DVDD.n4973 4.5005
R2071 DVDD.n4975 DVDD.n4887 4.5005
R2072 DVDD.n4977 DVDD.n4976 4.5005
R2073 DVDD.n4978 DVDD.n4886 4.5005
R2074 DVDD.n4980 DVDD.n4979 4.5005
R2075 DVDD.n4981 DVDD.n4885 4.5005
R2076 DVDD.n4983 DVDD.n4982 4.5005
R2077 DVDD.n4984 DVDD.n4884 4.5005
R2078 DVDD.n4986 DVDD.n4985 4.5005
R2079 DVDD.n4987 DVDD.n4883 4.5005
R2080 DVDD.n4989 DVDD.n4988 4.5005
R2081 DVDD.n4990 DVDD.n4882 4.5005
R2082 DVDD.n4992 DVDD.n4991 4.5005
R2083 DVDD.n4993 DVDD.n4881 4.5005
R2084 DVDD.n4997 DVDD.n4996 4.5005
R2085 DVDD.n4998 DVDD.n4874 4.5005
R2086 DVDD.n5000 DVDD.n4999 4.5005
R2087 DVDD.n5001 DVDD.n4873 4.5005
R2088 DVDD.n5003 DVDD.n5002 4.5005
R2089 DVDD.n5004 DVDD.n4872 4.5005
R2090 DVDD.n5006 DVDD.n5005 4.5005
R2091 DVDD.n5007 DVDD.n4871 4.5005
R2092 DVDD.n5009 DVDD.n5008 4.5005
R2093 DVDD.n5011 DVDD.n5010 4.5005
R2094 DVDD.n5013 DVDD.n5012 4.5005
R2095 DVDD.n5015 DVDD.n5014 4.5005
R2096 DVDD.n5017 DVDD.n5016 4.5005
R2097 DVDD.n5019 DVDD.n5018 4.5005
R2098 DVDD.n5021 DVDD.n5020 4.5005
R2099 DVDD.n5023 DVDD.n5022 4.5005
R2100 DVDD.n5025 DVDD.n5024 4.5005
R2101 DVDD.n5027 DVDD.n5026 4.5005
R2102 DVDD.n6113 DVDD.n4376 4.5005
R2103 DVDD.n4376 DVDD.n4305 4.5005
R2104 DVDD.n4388 DVDD.n4376 4.5005
R2105 DVDD.n6107 DVDD.n4305 4.5005
R2106 DVDD.n6107 DVDD.n4388 4.5005
R2107 DVDD.n6109 DVDD.n4305 4.5005
R2108 DVDD.n6109 DVDD.n4388 4.5005
R2109 DVDD.n6113 DVDD.n4377 4.5005
R2110 DVDD.n4377 DVDD.n4305 4.5005
R2111 DVDD.n4388 DVDD.n4377 4.5005
R2112 DVDD.n4315 DVDD.n4305 4.5005
R2113 DVDD.n6111 DVDD.n4315 4.5005
R2114 DVDD.n4388 DVDD.n4315 4.5005
R2115 DVDD.n6113 DVDD.n4315 4.5005
R2116 DVDD.n6113 DVDD.n4378 4.5005
R2117 DVDD.n4378 DVDD.n4305 4.5005
R2118 DVDD.n6111 DVDD.n4378 4.5005
R2119 DVDD.n4388 DVDD.n4378 4.5005
R2120 DVDD.n6113 DVDD.n4314 4.5005
R2121 DVDD.n4314 DVDD.n4305 4.5005
R2122 DVDD.n6111 DVDD.n4314 4.5005
R2123 DVDD.n4388 DVDD.n4314 4.5005
R2124 DVDD.n6113 DVDD.n4379 4.5005
R2125 DVDD.n4379 DVDD.n4305 4.5005
R2126 DVDD.n6111 DVDD.n4379 4.5005
R2127 DVDD.n4388 DVDD.n4379 4.5005
R2128 DVDD.n6113 DVDD.n4313 4.5005
R2129 DVDD.n4313 DVDD.n4305 4.5005
R2130 DVDD.n6111 DVDD.n4313 4.5005
R2131 DVDD.n4388 DVDD.n4313 4.5005
R2132 DVDD.n4380 DVDD.n4305 4.5005
R2133 DVDD.n6111 DVDD.n4380 4.5005
R2134 DVDD.n4388 DVDD.n4380 4.5005
R2135 DVDD.n6113 DVDD.n4380 4.5005
R2136 DVDD.n4312 DVDD.n4305 4.5005
R2137 DVDD.n6111 DVDD.n4312 4.5005
R2138 DVDD.n4388 DVDD.n4312 4.5005
R2139 DVDD.n6113 DVDD.n4312 4.5005
R2140 DVDD.n4381 DVDD.n4305 4.5005
R2141 DVDD.n6111 DVDD.n4381 4.5005
R2142 DVDD.n4388 DVDD.n4381 4.5005
R2143 DVDD.n6113 DVDD.n4381 4.5005
R2144 DVDD.n6113 DVDD.n4311 4.5005
R2145 DVDD.n4311 DVDD.n4305 4.5005
R2146 DVDD.n6111 DVDD.n4311 4.5005
R2147 DVDD.n4388 DVDD.n4311 4.5005
R2148 DVDD.n6113 DVDD.n4382 4.5005
R2149 DVDD.n4382 DVDD.n4305 4.5005
R2150 DVDD.n6111 DVDD.n4382 4.5005
R2151 DVDD.n4388 DVDD.n4382 4.5005
R2152 DVDD.n6113 DVDD.n4310 4.5005
R2153 DVDD.n4310 DVDD.n4305 4.5005
R2154 DVDD.n6111 DVDD.n4310 4.5005
R2155 DVDD.n4388 DVDD.n4310 4.5005
R2156 DVDD.n4383 DVDD.n4305 4.5005
R2157 DVDD.n6111 DVDD.n4383 4.5005
R2158 DVDD.n4388 DVDD.n4383 4.5005
R2159 DVDD.n6113 DVDD.n4383 4.5005
R2160 DVDD.n4309 DVDD.n4305 4.5005
R2161 DVDD.n6111 DVDD.n4309 4.5005
R2162 DVDD.n4388 DVDD.n4309 4.5005
R2163 DVDD.n6113 DVDD.n4309 4.5005
R2164 DVDD.n4384 DVDD.n4305 4.5005
R2165 DVDD.n6111 DVDD.n4384 4.5005
R2166 DVDD.n4388 DVDD.n4384 4.5005
R2167 DVDD.n6113 DVDD.n4384 4.5005
R2168 DVDD.n4308 DVDD.n4305 4.5005
R2169 DVDD.n6111 DVDD.n4308 4.5005
R2170 DVDD.n4388 DVDD.n4308 4.5005
R2171 DVDD.n6113 DVDD.n4308 4.5005
R2172 DVDD.n6113 DVDD.n4385 4.5005
R2173 DVDD.n4385 DVDD.n4305 4.5005
R2174 DVDD.n6111 DVDD.n4385 4.5005
R2175 DVDD.n4388 DVDD.n4385 4.5005
R2176 DVDD.n6113 DVDD.n4307 4.5005
R2177 DVDD.n4307 DVDD.n4305 4.5005
R2178 DVDD.n6111 DVDD.n4307 4.5005
R2179 DVDD.n4388 DVDD.n4307 4.5005
R2180 DVDD.n6113 DVDD.n4386 4.5005
R2181 DVDD.n4386 DVDD.n4305 4.5005
R2182 DVDD.n6111 DVDD.n4386 4.5005
R2183 DVDD.n4388 DVDD.n4386 4.5005
R2184 DVDD.n4306 DVDD.n4305 4.5005
R2185 DVDD.n6111 DVDD.n4306 4.5005
R2186 DVDD.n4388 DVDD.n4306 4.5005
R2187 DVDD.n6113 DVDD.n4306 4.5005
R2188 DVDD.n6112 DVDD.n4305 4.5005
R2189 DVDD.n6112 DVDD.n6111 4.5005
R2190 DVDD.n6112 DVDD.n4388 4.5005
R2191 DVDD.n6113 DVDD.n6112 4.5005
R2192 DVDD.n6095 DVDD.n5766 4.5005
R2193 DVDD.n5829 DVDD.n5766 4.5005
R2194 DVDD.n5891 DVDD.n5766 4.5005
R2195 DVDD.n6097 DVDD.n5766 4.5005
R2196 DVDD.n6095 DVDD.n5764 4.5005
R2197 DVDD.n5829 DVDD.n5764 4.5005
R2198 DVDD.n5891 DVDD.n5764 4.5005
R2199 DVDD.n6097 DVDD.n5764 4.5005
R2200 DVDD.n6095 DVDD.n5824 4.5005
R2201 DVDD.n5829 DVDD.n5824 4.5005
R2202 DVDD.n5891 DVDD.n5824 4.5005
R2203 DVDD.n6097 DVDD.n5824 4.5005
R2204 DVDD.n6095 DVDD.n5763 4.5005
R2205 DVDD.n5829 DVDD.n5763 4.5005
R2206 DVDD.n6097 DVDD.n5763 4.5005
R2207 DVDD.n5829 DVDD.n5825 4.5005
R2208 DVDD.n6097 DVDD.n5825 4.5005
R2209 DVDD.n5829 DVDD.n5762 4.5005
R2210 DVDD.n6097 DVDD.n5762 4.5005
R2211 DVDD.n5829 DVDD.n5826 4.5005
R2212 DVDD.n6097 DVDD.n5826 4.5005
R2213 DVDD.n5829 DVDD.n5761 4.5005
R2214 DVDD.n6097 DVDD.n5761 4.5005
R2215 DVDD.n5829 DVDD.n5827 4.5005
R2216 DVDD.n6097 DVDD.n5827 4.5005
R2217 DVDD.n5829 DVDD.n5760 4.5005
R2218 DVDD.n5891 DVDD.n5760 4.5005
R2219 DVDD.n6097 DVDD.n5760 4.5005
R2220 DVDD.n6096 DVDD.n5829 4.5005
R2221 DVDD.n6096 DVDD.n5891 4.5005
R2222 DVDD.n6097 DVDD.n6096 4.5005
R2223 DVDD.n6096 DVDD.n6095 4.5005
R2224 DVDD.n6704 DVDD.n3108 4.5005
R2225 DVDD.n3122 DVDD.n3108 4.5005
R2226 DVDD.n3184 DVDD.n3108 4.5005
R2227 DVDD.n6706 DVDD.n3108 4.5005
R2228 DVDD.n6704 DVDD.n3110 4.5005
R2229 DVDD.n3122 DVDD.n3110 4.5005
R2230 DVDD.n3184 DVDD.n3110 4.5005
R2231 DVDD.n6706 DVDD.n3110 4.5005
R2232 DVDD.n6704 DVDD.n3107 4.5005
R2233 DVDD.n3122 DVDD.n3107 4.5005
R2234 DVDD.n3184 DVDD.n3107 4.5005
R2235 DVDD.n6706 DVDD.n3107 4.5005
R2236 DVDD.n6704 DVDD.n3111 4.5005
R2237 DVDD.n3122 DVDD.n3111 4.5005
R2238 DVDD.n3184 DVDD.n3111 4.5005
R2239 DVDD.n6706 DVDD.n3111 4.5005
R2240 DVDD.n3122 DVDD.n3106 4.5005
R2241 DVDD.n3184 DVDD.n3106 4.5005
R2242 DVDD.n6706 DVDD.n3106 4.5005
R2243 DVDD.n6704 DVDD.n3106 4.5005
R2244 DVDD.n3122 DVDD.n3112 4.5005
R2245 DVDD.n3184 DVDD.n3112 4.5005
R2246 DVDD.n6706 DVDD.n3112 4.5005
R2247 DVDD.n6704 DVDD.n3112 4.5005
R2248 DVDD.n3122 DVDD.n3105 4.5005
R2249 DVDD.n3184 DVDD.n3105 4.5005
R2250 DVDD.n6706 DVDD.n3105 4.5005
R2251 DVDD.n6704 DVDD.n3105 4.5005
R2252 DVDD.n6704 DVDD.n3113 4.5005
R2253 DVDD.n3122 DVDD.n3113 4.5005
R2254 DVDD.n3184 DVDD.n3113 4.5005
R2255 DVDD.n6706 DVDD.n3113 4.5005
R2256 DVDD.n6704 DVDD.n3104 4.5005
R2257 DVDD.n3122 DVDD.n3104 4.5005
R2258 DVDD.n3184 DVDD.n3104 4.5005
R2259 DVDD.n6706 DVDD.n3104 4.5005
R2260 DVDD.n6704 DVDD.n3114 4.5005
R2261 DVDD.n3122 DVDD.n3114 4.5005
R2262 DVDD.n6706 DVDD.n3114 4.5005
R2263 DVDD.n3122 DVDD.n3103 4.5005
R2264 DVDD.n6706 DVDD.n3103 4.5005
R2265 DVDD.n3122 DVDD.n3115 4.5005
R2266 DVDD.n6706 DVDD.n3115 4.5005
R2267 DVDD.n3122 DVDD.n3102 4.5005
R2268 DVDD.n6706 DVDD.n3102 4.5005
R2269 DVDD.n3122 DVDD.n3116 4.5005
R2270 DVDD.n6706 DVDD.n3116 4.5005
R2271 DVDD.n3122 DVDD.n3101 4.5005
R2272 DVDD.n6706 DVDD.n3101 4.5005
R2273 DVDD.n3122 DVDD.n3117 4.5005
R2274 DVDD.n3184 DVDD.n3117 4.5005
R2275 DVDD.n6706 DVDD.n3117 4.5005
R2276 DVDD.n3122 DVDD.n3100 4.5005
R2277 DVDD.n3184 DVDD.n3100 4.5005
R2278 DVDD.n6706 DVDD.n3100 4.5005
R2279 DVDD.n6704 DVDD.n3100 4.5005
R2280 DVDD.n3122 DVDD.n3118 4.5005
R2281 DVDD.n3184 DVDD.n3118 4.5005
R2282 DVDD.n6706 DVDD.n3118 4.5005
R2283 DVDD.n6704 DVDD.n3118 4.5005
R2284 DVDD.n6704 DVDD.n3099 4.5005
R2285 DVDD.n3122 DVDD.n3099 4.5005
R2286 DVDD.n3184 DVDD.n3099 4.5005
R2287 DVDD.n6706 DVDD.n3099 4.5005
R2288 DVDD.n6704 DVDD.n3119 4.5005
R2289 DVDD.n3122 DVDD.n3119 4.5005
R2290 DVDD.n3184 DVDD.n3119 4.5005
R2291 DVDD.n6706 DVDD.n3119 4.5005
R2292 DVDD.n6704 DVDD.n3098 4.5005
R2293 DVDD.n3122 DVDD.n3098 4.5005
R2294 DVDD.n3184 DVDD.n3098 4.5005
R2295 DVDD.n6706 DVDD.n3098 4.5005
R2296 DVDD.n3122 DVDD.n3120 4.5005
R2297 DVDD.n3184 DVDD.n3120 4.5005
R2298 DVDD.n6706 DVDD.n3120 4.5005
R2299 DVDD.n6704 DVDD.n3120 4.5005
R2300 DVDD.n3122 DVDD.n3097 4.5005
R2301 DVDD.n3184 DVDD.n3097 4.5005
R2302 DVDD.n6706 DVDD.n3097 4.5005
R2303 DVDD.n6704 DVDD.n3097 4.5005
R2304 DVDD.n6705 DVDD.n3122 4.5005
R2305 DVDD.n6705 DVDD.n3184 4.5005
R2306 DVDD.n6706 DVDD.n6705 4.5005
R2307 DVDD.n6705 DVDD.n6704 4.5005
R2308 DVDD.n7806 DVDD.n2179 4.5005
R2309 DVDD.n2179 DVDD.n2171 4.5005
R2310 DVDD.n7799 DVDD.n2179 4.5005
R2311 DVDD.n7803 DVDD.n2179 4.5005
R2312 DVDD.n7806 DVDD.n2180 4.5005
R2313 DVDD.n2180 DVDD.n2171 4.5005
R2314 DVDD.n7799 DVDD.n2180 4.5005
R2315 DVDD.n7803 DVDD.n2180 4.5005
R2316 DVDD.n7806 DVDD.n2178 4.5005
R2317 DVDD.n2178 DVDD.n2171 4.5005
R2318 DVDD.n7799 DVDD.n2178 4.5005
R2319 DVDD.n7803 DVDD.n2178 4.5005
R2320 DVDD.n2181 DVDD.n2171 4.5005
R2321 DVDD.n7799 DVDD.n2181 4.5005
R2322 DVDD.n7803 DVDD.n2181 4.5005
R2323 DVDD.n7806 DVDD.n2181 4.5005
R2324 DVDD.n2177 DVDD.n2171 4.5005
R2325 DVDD.n7799 DVDD.n2177 4.5005
R2326 DVDD.n7803 DVDD.n2177 4.5005
R2327 DVDD.n7806 DVDD.n2177 4.5005
R2328 DVDD.n2182 DVDD.n2171 4.5005
R2329 DVDD.n7799 DVDD.n2182 4.5005
R2330 DVDD.n7803 DVDD.n2182 4.5005
R2331 DVDD.n7806 DVDD.n2182 4.5005
R2332 DVDD.n2176 DVDD.n2171 4.5005
R2333 DVDD.n7799 DVDD.n2176 4.5005
R2334 DVDD.n7803 DVDD.n2176 4.5005
R2335 DVDD.n7806 DVDD.n2176 4.5005
R2336 DVDD.n7806 DVDD.n2183 4.5005
R2337 DVDD.n2183 DVDD.n2171 4.5005
R2338 DVDD.n7799 DVDD.n2183 4.5005
R2339 DVDD.n7803 DVDD.n2183 4.5005
R2340 DVDD.n7806 DVDD.n2175 4.5005
R2341 DVDD.n2175 DVDD.n2171 4.5005
R2342 DVDD.n7799 DVDD.n2175 4.5005
R2343 DVDD.n7803 DVDD.n2175 4.5005
R2344 DVDD.n7806 DVDD.n2184 4.5005
R2345 DVDD.n2184 DVDD.n2171 4.5005
R2346 DVDD.n7799 DVDD.n2184 4.5005
R2347 DVDD.n7803 DVDD.n2184 4.5005
R2348 DVDD.n2174 DVDD.n2171 4.5005
R2349 DVDD.n7799 DVDD.n2174 4.5005
R2350 DVDD.n7803 DVDD.n2174 4.5005
R2351 DVDD.n7806 DVDD.n2174 4.5005
R2352 DVDD.n2185 DVDD.n2171 4.5005
R2353 DVDD.n7799 DVDD.n2185 4.5005
R2354 DVDD.n7803 DVDD.n2185 4.5005
R2355 DVDD.n7806 DVDD.n2185 4.5005
R2356 DVDD.n2173 DVDD.n2171 4.5005
R2357 DVDD.n7799 DVDD.n2173 4.5005
R2358 DVDD.n7803 DVDD.n2173 4.5005
R2359 DVDD.n7806 DVDD.n2173 4.5005
R2360 DVDD.n7806 DVDD.n2186 4.5005
R2361 DVDD.n2186 DVDD.n2171 4.5005
R2362 DVDD.n7799 DVDD.n2186 4.5005
R2363 DVDD.n7803 DVDD.n2186 4.5005
R2364 DVDD.n7806 DVDD.n2172 4.5005
R2365 DVDD.n2172 DVDD.n2171 4.5005
R2366 DVDD.n7799 DVDD.n2172 4.5005
R2367 DVDD.n7803 DVDD.n2172 4.5005
R2368 DVDD.n7806 DVDD.n2187 4.5005
R2369 DVDD.n2187 DVDD.n2171 4.5005
R2370 DVDD.n7803 DVDD.n2187 4.5005
R2371 DVDD.n2196 DVDD.n2171 4.5005
R2372 DVDD.n7803 DVDD.n2196 4.5005
R2373 DVDD.n7795 DVDD.n2171 4.5005
R2374 DVDD.n7803 DVDD.n7795 4.5005
R2375 DVDD.n2195 DVDD.n2171 4.5005
R2376 DVDD.n7803 DVDD.n2195 4.5005
R2377 DVDD.n7801 DVDD.n2171 4.5005
R2378 DVDD.n7803 DVDD.n7801 4.5005
R2379 DVDD.n2194 DVDD.n2171 4.5005
R2380 DVDD.n7803 DVDD.n2194 4.5005
R2381 DVDD.n7802 DVDD.n2171 4.5005
R2382 DVDD.n7803 DVDD.n7802 4.5005
R2383 DVDD.n7804 DVDD.n2171 4.5005
R2384 DVDD.n7804 DVDD.n7803 4.5005
R2385 DVDD.n2191 DVDD.n2171 4.5005
R2386 DVDD.n7799 DVDD.n2191 4.5005
R2387 DVDD.n7803 DVDD.n2191 4.5005
R2388 DVDD.n7776 DVDD.n2235 4.5005
R2389 DVDD.n7778 DVDD.n2235 4.5005
R2390 DVDD.n2235 DVDD.n2207 4.5005
R2391 DVDD.n7778 DVDD.n2237 4.5005
R2392 DVDD.n2237 DVDD.n2207 4.5005
R2393 DVDD.n7778 DVDD.n2234 4.5005
R2394 DVDD.n2234 DVDD.n2207 4.5005
R2395 DVDD.n7778 DVDD.n2238 4.5005
R2396 DVDD.n2238 DVDD.n2207 4.5005
R2397 DVDD.n7778 DVDD.n2233 4.5005
R2398 DVDD.n2233 DVDD.n2207 4.5005
R2399 DVDD.n7776 DVDD.n2239 4.5005
R2400 DVDD.n7778 DVDD.n2239 4.5005
R2401 DVDD.n2239 DVDD.n2207 4.5005
R2402 DVDD.n7776 DVDD.n2216 4.5005
R2403 DVDD.n7778 DVDD.n2216 4.5005
R2404 DVDD.n7780 DVDD.n2216 4.5005
R2405 DVDD.n2216 DVDD.n2207 4.5005
R2406 DVDD.n7776 DVDD.n2240 4.5005
R2407 DVDD.n7778 DVDD.n2240 4.5005
R2408 DVDD.n2240 DVDD.n2207 4.5005
R2409 DVDD.n7778 DVDD.n2232 4.5005
R2410 DVDD.n2232 DVDD.n2207 4.5005
R2411 DVDD.n7778 DVDD.n2241 4.5005
R2412 DVDD.n2241 DVDD.n2207 4.5005
R2413 DVDD.n7778 DVDD.n2231 4.5005
R2414 DVDD.n2231 DVDD.n2207 4.5005
R2415 DVDD.n7778 DVDD.n2242 4.5005
R2416 DVDD.n2242 DVDD.n2207 4.5005
R2417 DVDD.n7776 DVDD.n2230 4.5005
R2418 DVDD.n7778 DVDD.n2230 4.5005
R2419 DVDD.n2230 DVDD.n2207 4.5005
R2420 DVDD.n7776 DVDD.n2221 4.5005
R2421 DVDD.n7778 DVDD.n2221 4.5005
R2422 DVDD.n7780 DVDD.n2221 4.5005
R2423 DVDD.n2221 DVDD.n2207 4.5005
R2424 DVDD.n7776 DVDD.n2229 4.5005
R2425 DVDD.n7778 DVDD.n2229 4.5005
R2426 DVDD.n2229 DVDD.n2207 4.5005
R2427 DVDD.n7778 DVDD.n2243 4.5005
R2428 DVDD.n2243 DVDD.n2207 4.5005
R2429 DVDD.n7778 DVDD.n2228 4.5005
R2430 DVDD.n2228 DVDD.n2207 4.5005
R2431 DVDD.n7778 DVDD.n2244 4.5005
R2432 DVDD.n2244 DVDD.n2207 4.5005
R2433 DVDD.n7778 DVDD.n2227 4.5005
R2434 DVDD.n2227 DVDD.n2207 4.5005
R2435 DVDD.n7776 DVDD.n2245 4.5005
R2436 DVDD.n7778 DVDD.n2245 4.5005
R2437 DVDD.n2245 DVDD.n2207 4.5005
R2438 DVDD.n7776 DVDD.n2212 4.5005
R2439 DVDD.n7778 DVDD.n2212 4.5005
R2440 DVDD.n7780 DVDD.n2212 4.5005
R2441 DVDD.n2212 DVDD.n2207 4.5005
R2442 DVDD.n7777 DVDD.n7776 4.5005
R2443 DVDD.n7778 DVDD.n7777 4.5005
R2444 DVDD.n7777 DVDD.n2207 4.5005
R2445 DVDD.n7778 DVDD.n2226 4.5005
R2446 DVDD.n2226 DVDD.n2207 4.5005
R2447 DVDD.n7779 DVDD.n7778 4.5005
R2448 DVDD.n7780 DVDD.n7779 4.5005
R2449 DVDD.n7779 DVDD.n2207 4.5005
R2450 DVDD.n1619 DVDD.n1599 4.5005
R2451 DVDD.n8321 DVDD.n1599 4.5005
R2452 DVDD.n1628 DVDD.n1599 4.5005
R2453 DVDD.n8323 DVDD.n1599 4.5005
R2454 DVDD.n8323 DVDD.n1601 4.5005
R2455 DVDD.n1628 DVDD.n1601 4.5005
R2456 DVDD.n8321 DVDD.n1601 4.5005
R2457 DVDD.n1619 DVDD.n1601 4.5005
R2458 DVDD.n1619 DVDD.n1598 4.5005
R2459 DVDD.n8321 DVDD.n1598 4.5005
R2460 DVDD.n8323 DVDD.n1598 4.5005
R2461 DVDD.n8321 DVDD.n1602 4.5005
R2462 DVDD.n8323 DVDD.n1602 4.5005
R2463 DVDD.n8321 DVDD.n1597 4.5005
R2464 DVDD.n8323 DVDD.n1597 4.5005
R2465 DVDD.n8321 DVDD.n1603 4.5005
R2466 DVDD.n8323 DVDD.n1603 4.5005
R2467 DVDD.n8321 DVDD.n1596 4.5005
R2468 DVDD.n8323 DVDD.n1596 4.5005
R2469 DVDD.n1619 DVDD.n1604 4.5005
R2470 DVDD.n8321 DVDD.n1604 4.5005
R2471 DVDD.n8323 DVDD.n1604 4.5005
R2472 DVDD.n8323 DVDD.n1595 4.5005
R2473 DVDD.n1628 DVDD.n1595 4.5005
R2474 DVDD.n8321 DVDD.n1595 4.5005
R2475 DVDD.n1619 DVDD.n1595 4.5005
R2476 DVDD.n8323 DVDD.n1605 4.5005
R2477 DVDD.n1628 DVDD.n1605 4.5005
R2478 DVDD.n8321 DVDD.n1605 4.5005
R2479 DVDD.n1619 DVDD.n1605 4.5005
R2480 DVDD.n1619 DVDD.n1594 4.5005
R2481 DVDD.n8321 DVDD.n1594 4.5005
R2482 DVDD.n8323 DVDD.n1594 4.5005
R2483 DVDD.n8321 DVDD.n1606 4.5005
R2484 DVDD.n8323 DVDD.n1606 4.5005
R2485 DVDD.n8321 DVDD.n1593 4.5005
R2486 DVDD.n8323 DVDD.n1593 4.5005
R2487 DVDD.n8321 DVDD.n1607 4.5005
R2488 DVDD.n8323 DVDD.n1607 4.5005
R2489 DVDD.n8321 DVDD.n1592 4.5005
R2490 DVDD.n1628 DVDD.n1592 4.5005
R2491 DVDD.n8323 DVDD.n1592 4.5005
R2492 DVDD.n1619 DVDD.n1608 4.5005
R2493 DVDD.n8321 DVDD.n1608 4.5005
R2494 DVDD.n1628 DVDD.n1608 4.5005
R2495 DVDD.n8323 DVDD.n1608 4.5005
R2496 DVDD.n1619 DVDD.n1591 4.5005
R2497 DVDD.n8321 DVDD.n1591 4.5005
R2498 DVDD.n1628 DVDD.n1591 4.5005
R2499 DVDD.n8323 DVDD.n1591 4.5005
R2500 DVDD.n1619 DVDD.n1609 4.5005
R2501 DVDD.n8321 DVDD.n1609 4.5005
R2502 DVDD.n1628 DVDD.n1609 4.5005
R2503 DVDD.n8323 DVDD.n1609 4.5005
R2504 DVDD.n1619 DVDD.n1590 4.5005
R2505 DVDD.n8321 DVDD.n1590 4.5005
R2506 DVDD.n8323 DVDD.n1590 4.5005
R2507 DVDD.n8321 DVDD.n1610 4.5005
R2508 DVDD.n8323 DVDD.n1610 4.5005
R2509 DVDD.n8321 DVDD.n1589 4.5005
R2510 DVDD.n8323 DVDD.n1589 4.5005
R2511 DVDD.n8321 DVDD.n1611 4.5005
R2512 DVDD.n8323 DVDD.n1611 4.5005
R2513 DVDD.n8321 DVDD.n1588 4.5005
R2514 DVDD.n8323 DVDD.n1588 4.5005
R2515 DVDD.n8322 DVDD.n1619 4.5005
R2516 DVDD.n8322 DVDD.n8321 4.5005
R2517 DVDD.n8323 DVDD.n8322 4.5005
R2518 DVDD.n4870 DVDD.n4868 4.5005
R2519 DVDD.n4876 DVDD.n4875 4.5005
R2520 DVDD.n4878 DVDD.n4877 4.5005
R2521 DVDD.n8516 DVDD.n8515 4.5005
R2522 DVDD.n8543 DVDD.n8516 4.5005
R2523 DVDD.n8545 DVDD.n8544 4.5005
R2524 DVDD.n8544 DVDD.n8543 4.5005
R2525 DVDD.n8427 DVDD.n8426 4.5005
R2526 DVDD.n8428 DVDD.n8427 4.5005
R2527 DVDD.n7358 DVDD.n7357 4.5005
R2528 DVDD.n7358 DVDD.n1335 4.5005
R2529 DVDD.n7353 DVDD.n1458 4.5005
R2530 DVDD.n1458 DVDD.n1335 4.5005
R2531 DVDD.n8428 DVDD.n1457 4.5005
R2532 DVDD.n8426 DVDD.n1457 4.5005
R2533 DVDD.n8421 DVDD.n1457 4.5005
R2534 DVDD.n8426 DVDD.n1418 4.5005
R2535 DVDD.n8421 DVDD.n1418 4.5005
R2536 DVDD.n8505 DVDD.n1414 4.5005
R2537 DVDD.n8505 DVDD.n8504 4.5005
R2538 DVDD.n8504 DVDD.n1416 4.5005
R2539 DVDD.n1416 DVDD.n1414 4.5005
R2540 DVDD.n8507 DVDD.n1416 4.5005
R2541 DVDD.n8508 DVDD.n1414 4.5005
R2542 DVDD.n8508 DVDD.n8507 4.5005
R2543 DVDD.n8511 DVDD.n1408 4.5005
R2544 DVDD.n8511 DVDD.n1370 4.5005
R2545 DVDD.n1410 DVDD.n1370 4.5005
R2546 DVDD.n1410 DVDD.n1408 4.5005
R2547 DVDD.n8513 DVDD.n1410 4.5005
R2548 DVDD.n8514 DVDD.n1408 4.5005
R2549 DVDD.n8514 DVDD.n8513 4.5005
R2550 DVDD.n7182 DVDD.n7152 4.5005
R2551 DVDD.n7180 DVDD.n7152 4.5005
R2552 DVDD.n7177 DVDD.n7158 4.5005
R2553 DVDD.n7175 DVDD.n7158 4.5005
R2554 DVDD.n7186 DVDD.n7145 4.5005
R2555 DVDD.n7184 DVDD.n7145 4.5005
R2556 DVDD.n7186 DVDD.n7143 4.5005
R2557 DVDD.n7148 DVDD.n7143 4.5005
R2558 DVDD.n7146 DVDD.n7143 4.5005
R2559 DVDD.n7184 DVDD.n7143 4.5005
R2560 DVDD.n7182 DVDD.n7151 4.5005
R2561 DVDD.n7156 DVDD.n7151 4.5005
R2562 DVDD.n7154 DVDD.n7151 4.5005
R2563 DVDD.n7180 DVDD.n7151 4.5005
R2564 DVDD.n7177 DVDD.n7157 4.5005
R2565 DVDD.n7162 DVDD.n7157 4.5005
R2566 DVDD.n7160 DVDD.n7157 4.5005
R2567 DVDD.n7175 DVDD.n7157 4.5005
R2568 DVDD.n7186 DVDD.n7185 4.5005
R2569 DVDD.n7185 DVDD.n7148 4.5005
R2570 DVDD.n7185 DVDD.n7146 4.5005
R2571 DVDD.n7185 DVDD.n7184 4.5005
R2572 DVDD.n7182 DVDD.n7181 4.5005
R2573 DVDD.n7181 DVDD.n7156 4.5005
R2574 DVDD.n7181 DVDD.n7154 4.5005
R2575 DVDD.n7181 DVDD.n7180 4.5005
R2576 DVDD.n7177 DVDD.n7176 4.5005
R2577 DVDD.n7176 DVDD.n7162 4.5005
R2578 DVDD.n7176 DVDD.n7160 4.5005
R2579 DVDD.n7176 DVDD.n7175 4.5005
R2580 DVDD.n7359 DVDD.n1306 4.5005
R2581 DVDD.n8636 DVDD.n1314 4.5005
R2582 DVDD.n8631 DVDD.n8628 4.5005
R2583 DVDD.n7362 DVDD.n7361 4.5005
R2584 DVDD.n7361 DVDD.n1306 4.5005
R2585 DVDD.n8635 DVDD.n1311 4.5005
R2586 DVDD.n8636 DVDD.n8635 4.5005
R2587 DVDD.n8630 DVDD.n1319 4.5005
R2588 DVDD.n8631 DVDD.n8630 4.5005
R2589 DVDD.n7362 DVDD.n7342 4.5005
R2590 DVDD.n7342 DVDD.n1306 4.5005
R2591 DVDD.n1313 DVDD.n1311 4.5005
R2592 DVDD.n8636 DVDD.n1313 4.5005
R2593 DVDD.n1321 DVDD.n1319 4.5005
R2594 DVDD.n8631 DVDD.n1321 4.5005
R2595 DVDD.n7363 DVDD.n1508 4.5005
R2596 DVDD.n7363 DVDD.n7362 4.5005
R2597 DVDD.n7363 DVDD.n1306 4.5005
R2598 DVDD.n8638 DVDD.n8637 4.5005
R2599 DVDD.n8637 DVDD.n1311 4.5005
R2600 DVDD.n8637 DVDD.n8636 4.5005
R2601 DVDD.n8633 DVDD.n8632 4.5005
R2602 DVDD.n8632 DVDD.n1319 4.5005
R2603 DVDD.n8632 DVDD.n8631 4.5005
R2604 DVDD.n8378 DVDD.n8377 4.5005
R2605 DVDD.n8377 DVDD.n1507 4.5005
R2606 DVDD.n8377 DVDD.n8376 4.5005
R2607 DVDD.n8371 DVDD.n1507 4.5005
R2608 DVDD.n7191 DVDD.n7138 4.5005
R2609 DVDD.n7189 DVDD.n7138 4.5005
R2610 DVDD.n7191 DVDD.n7137 4.5005
R2611 DVDD.n7142 DVDD.n7137 4.5005
R2612 DVDD.n7140 DVDD.n7137 4.5005
R2613 DVDD.n7189 DVDD.n7137 4.5005
R2614 DVDD.n7191 DVDD.n7190 4.5005
R2615 DVDD.n7190 DVDD.n7142 4.5005
R2616 DVDD.n7190 DVDD.n7140 4.5005
R2617 DVDD.n7190 DVDD.n7189 4.5005
R2618 DVDD.n7695 DVDD.n2350 4.5005
R2619 DVDD.n7690 DVDD.n7689 4.5005
R2620 DVDD.n7694 DVDD.n7689 4.5005
R2621 DVDD.n7694 DVDD.n2352 4.5005
R2622 DVDD.n7694 DVDD.n7693 4.5005
R2623 DVDD.n7694 DVDD.n2351 4.5005
R2624 DVDD.n7695 DVDD.n7694 4.5005
R2625 DVDD.n1543 DVDD.n1529 4.5005
R2626 DVDD.n1543 DVDD.n1530 4.5005
R2627 DVDD.n8358 DVDD.n1543 4.5005
R2628 DVDD.n1546 DVDD.n1530 4.5005
R2629 DVDD.n8358 DVDD.n1546 4.5005
R2630 DVDD.n1542 DVDD.n1530 4.5005
R2631 DVDD.n8358 DVDD.n1542 4.5005
R2632 DVDD.n1548 DVDD.n1530 4.5005
R2633 DVDD.n8358 DVDD.n1548 4.5005
R2634 DVDD.n1541 DVDD.n1530 4.5005
R2635 DVDD.n8358 DVDD.n1541 4.5005
R2636 DVDD.n1549 DVDD.n1529 4.5005
R2637 DVDD.n1549 DVDD.n1530 4.5005
R2638 DVDD.n8358 DVDD.n1549 4.5005
R2639 DVDD.n8358 DVDD.n1540 4.5005
R2640 DVDD.n8356 DVDD.n1540 4.5005
R2641 DVDD.n1540 DVDD.n1530 4.5005
R2642 DVDD.n1540 DVDD.n1529 4.5005
R2643 DVDD.n8358 DVDD.n1550 4.5005
R2644 DVDD.n8356 DVDD.n1550 4.5005
R2645 DVDD.n1550 DVDD.n1530 4.5005
R2646 DVDD.n1550 DVDD.n1529 4.5005
R2647 DVDD.n1539 DVDD.n1529 4.5005
R2648 DVDD.n1539 DVDD.n1530 4.5005
R2649 DVDD.n8358 DVDD.n1539 4.5005
R2650 DVDD.n1552 DVDD.n1530 4.5005
R2651 DVDD.n8358 DVDD.n1552 4.5005
R2652 DVDD.n1538 DVDD.n1530 4.5005
R2653 DVDD.n8358 DVDD.n1538 4.5005
R2654 DVDD.n1554 DVDD.n1530 4.5005
R2655 DVDD.n8358 DVDD.n1554 4.5005
R2656 DVDD.n1537 DVDD.n1530 4.5005
R2657 DVDD.n8356 DVDD.n1537 4.5005
R2658 DVDD.n8358 DVDD.n1537 4.5005
R2659 DVDD.n1555 DVDD.n1529 4.5005
R2660 DVDD.n1555 DVDD.n1530 4.5005
R2661 DVDD.n8356 DVDD.n1555 4.5005
R2662 DVDD.n8358 DVDD.n1555 4.5005
R2663 DVDD.n1536 DVDD.n1529 4.5005
R2664 DVDD.n1536 DVDD.n1530 4.5005
R2665 DVDD.n8356 DVDD.n1536 4.5005
R2666 DVDD.n8358 DVDD.n1536 4.5005
R2667 DVDD.n1556 DVDD.n1529 4.5005
R2668 DVDD.n1556 DVDD.n1530 4.5005
R2669 DVDD.n8356 DVDD.n1556 4.5005
R2670 DVDD.n8358 DVDD.n1556 4.5005
R2671 DVDD.n1535 DVDD.n1529 4.5005
R2672 DVDD.n1535 DVDD.n1530 4.5005
R2673 DVDD.n8358 DVDD.n1535 4.5005
R2674 DVDD.n1558 DVDD.n1530 4.5005
R2675 DVDD.n8358 DVDD.n1558 4.5005
R2676 DVDD.n1534 DVDD.n1530 4.5005
R2677 DVDD.n8358 DVDD.n1534 4.5005
R2678 DVDD.n1560 DVDD.n1530 4.5005
R2679 DVDD.n8358 DVDD.n1560 4.5005
R2680 DVDD.n1533 DVDD.n1530 4.5005
R2681 DVDD.n8358 DVDD.n1533 4.5005
R2682 DVDD.n8359 DVDD.n1529 4.5005
R2683 DVDD.n8359 DVDD.n1530 4.5005
R2684 DVDD.n8359 DVDD.n8358 4.5005
R2685 DVDD.n8358 DVDD.n1532 4.5005
R2686 DVDD.n8356 DVDD.n1532 4.5005
R2687 DVDD.n1532 DVDD.n1530 4.5005
R2688 DVDD.n1532 DVDD.n1529 4.5005
R2689 DVDD.n7660 DVDD.n2387 4.5005
R2690 DVDD.n2387 DVDD.n2374 4.5005
R2691 DVDD.n7679 DVDD.n2387 4.5005
R2692 DVDD.n2390 DVDD.n2374 4.5005
R2693 DVDD.n7679 DVDD.n2390 4.5005
R2694 DVDD.n2386 DVDD.n2374 4.5005
R2695 DVDD.n2386 DVDD.n2372 4.5005
R2696 DVDD.n7679 DVDD.n2386 4.5005
R2697 DVDD.n2392 DVDD.n2374 4.5005
R2698 DVDD.n7679 DVDD.n2392 4.5005
R2699 DVDD.n2385 DVDD.n2374 4.5005
R2700 DVDD.n7679 DVDD.n2385 4.5005
R2701 DVDD.n2394 DVDD.n2374 4.5005
R2702 DVDD.n7679 DVDD.n2394 4.5005
R2703 DVDD.n2384 DVDD.n2374 4.5005
R2704 DVDD.n7679 DVDD.n2384 4.5005
R2705 DVDD.n2395 DVDD.n2374 4.5005
R2706 DVDD.n2395 DVDD.n2372 4.5005
R2707 DVDD.n7679 DVDD.n2395 4.5005
R2708 DVDD.n2383 DVDD.n2374 4.5005
R2709 DVDD.n7679 DVDD.n2383 4.5005
R2710 DVDD.n2397 DVDD.n2374 4.5005
R2711 DVDD.n7679 DVDD.n2397 4.5005
R2712 DVDD.n2382 DVDD.n2374 4.5005
R2713 DVDD.n7679 DVDD.n2382 4.5005
R2714 DVDD.n2399 DVDD.n2374 4.5005
R2715 DVDD.n7679 DVDD.n2399 4.5005
R2716 DVDD.n2381 DVDD.n2374 4.5005
R2717 DVDD.n2381 DVDD.n2372 4.5005
R2718 DVDD.n7679 DVDD.n2381 4.5005
R2719 DVDD.n2401 DVDD.n2374 4.5005
R2720 DVDD.n7679 DVDD.n2401 4.5005
R2721 DVDD.n2380 DVDD.n2374 4.5005
R2722 DVDD.n7679 DVDD.n2380 4.5005
R2723 DVDD.n2403 DVDD.n2374 4.5005
R2724 DVDD.n7679 DVDD.n2403 4.5005
R2725 DVDD.n2379 DVDD.n2374 4.5005
R2726 DVDD.n7679 DVDD.n2379 4.5005
R2727 DVDD.n7680 DVDD.n2374 4.5005
R2728 DVDD.n7680 DVDD.n2372 4.5005
R2729 DVDD.n7680 DVDD.n7679 4.5005
R2730 DVDD.n6983 DVDD.n6934 4.5005
R2731 DVDD.n6983 DVDD.n6982 4.5005
R2732 DVDD.n6940 DVDD.n6934 4.5005
R2733 DVDD.n6982 DVDD.n6940 4.5005
R2734 DVDD.n6938 DVDD.n6934 4.5005
R2735 DVDD.n6982 DVDD.n6938 4.5005
R2736 DVDD.n6941 DVDD.n6934 4.5005
R2737 DVDD.n6982 DVDD.n6941 4.5005
R2738 DVDD.n6937 DVDD.n6934 4.5005
R2739 DVDD.n6982 DVDD.n6937 4.5005
R2740 DVDD.n6981 DVDD.n6934 4.5005
R2741 DVDD.n6982 DVDD.n6981 4.5005
R2742 DVDD.n6936 DVDD.n6934 4.5005
R2743 DVDD.n6982 DVDD.n6936 4.5005
R2744 DVDD.n6985 DVDD.n2642 4.5005
R2745 DVDD.n6934 DVDD.n2642 4.5005
R2746 DVDD.n6982 DVDD.n2642 4.5005
R2747 DVDD.n6934 DVDD.n2630 4.5005
R2748 DVDD.n6979 DVDD.n2630 4.5005
R2749 DVDD.n6982 DVDD.n2630 4.5005
R2750 DVDD.n6934 DVDD.n6932 4.5005
R2751 DVDD.n6979 DVDD.n6932 4.5005
R2752 DVDD.n6982 DVDD.n6932 4.5005
R2753 DVDD.n6985 DVDD.n2637 4.5005
R2754 DVDD.n6934 DVDD.n2637 4.5005
R2755 DVDD.n6979 DVDD.n2637 4.5005
R2756 DVDD.n6982 DVDD.n2637 4.5005
R2757 DVDD.n6985 DVDD.n2643 4.5005
R2758 DVDD.n6934 DVDD.n2643 4.5005
R2759 DVDD.n6979 DVDD.n2643 4.5005
R2760 DVDD.n6982 DVDD.n2643 4.5005
R2761 DVDD.n6985 DVDD.n2636 4.5005
R2762 DVDD.n6934 DVDD.n2636 4.5005
R2763 DVDD.n6979 DVDD.n2636 4.5005
R2764 DVDD.n6982 DVDD.n2636 4.5005
R2765 DVDD.n6934 DVDD.n2631 4.5005
R2766 DVDD.n6979 DVDD.n2631 4.5005
R2767 DVDD.n6982 DVDD.n2631 4.5005
R2768 DVDD.n6934 DVDD.n2648 4.5005
R2769 DVDD.n6979 DVDD.n2648 4.5005
R2770 DVDD.n6982 DVDD.n2648 4.5005
R2771 DVDD.n6934 DVDD.n2632 4.5005
R2772 DVDD.n6979 DVDD.n2632 4.5005
R2773 DVDD.n6982 DVDD.n2632 4.5005
R2774 DVDD.n6985 DVDD.n2644 4.5005
R2775 DVDD.n6934 DVDD.n2644 4.5005
R2776 DVDD.n6979 DVDD.n2644 4.5005
R2777 DVDD.n6982 DVDD.n2644 4.5005
R2778 DVDD.n6985 DVDD.n2635 4.5005
R2779 DVDD.n6934 DVDD.n2635 4.5005
R2780 DVDD.n6979 DVDD.n2635 4.5005
R2781 DVDD.n6982 DVDD.n2635 4.5005
R2782 DVDD.n6985 DVDD.n2645 4.5005
R2783 DVDD.n6934 DVDD.n2645 4.5005
R2784 DVDD.n6979 DVDD.n2645 4.5005
R2785 DVDD.n6982 DVDD.n2645 4.5005
R2786 DVDD.n6985 DVDD.n2634 4.5005
R2787 DVDD.n6934 DVDD.n2634 4.5005
R2788 DVDD.n6979 DVDD.n2634 4.5005
R2789 DVDD.n6982 DVDD.n2634 4.5005
R2790 DVDD.n6934 DVDD.n2647 4.5005
R2791 DVDD.n6979 DVDD.n2647 4.5005
R2792 DVDD.n6982 DVDD.n2647 4.5005
R2793 DVDD.n6934 DVDD.n2633 4.5005
R2794 DVDD.n6979 DVDD.n2633 4.5005
R2795 DVDD.n6982 DVDD.n2633 4.5005
R2796 DVDD.n6934 DVDD.n2646 4.5005
R2797 DVDD.n6979 DVDD.n2646 4.5005
R2798 DVDD.n6982 DVDD.n2646 4.5005
R2799 DVDD.n2671 DVDD.n2657 4.5005
R2800 DVDD.n2671 DVDD.n2659 4.5005
R2801 DVDD.n2671 DVDD.n2656 4.5005
R2802 DVDD.n6924 DVDD.n2671 4.5005
R2803 DVDD.n2673 DVDD.n2657 4.5005
R2804 DVDD.n2673 DVDD.n2659 4.5005
R2805 DVDD.n2673 DVDD.n2656 4.5005
R2806 DVDD.n6924 DVDD.n2673 4.5005
R2807 DVDD.n2670 DVDD.n2657 4.5005
R2808 DVDD.n2670 DVDD.n2659 4.5005
R2809 DVDD.n2670 DVDD.n2656 4.5005
R2810 DVDD.n6924 DVDD.n2670 4.5005
R2811 DVDD.n2674 DVDD.n2659 4.5005
R2812 DVDD.n2674 DVDD.n2656 4.5005
R2813 DVDD.n6924 DVDD.n2674 4.5005
R2814 DVDD.n2669 DVDD.n2659 4.5005
R2815 DVDD.n2669 DVDD.n2656 4.5005
R2816 DVDD.n6924 DVDD.n2669 4.5005
R2817 DVDD.n2723 DVDD.n2659 4.5005
R2818 DVDD.n2723 DVDD.n2656 4.5005
R2819 DVDD.n6924 DVDD.n2723 4.5005
R2820 DVDD.n2668 DVDD.n2657 4.5005
R2821 DVDD.n2668 DVDD.n2659 4.5005
R2822 DVDD.n2668 DVDD.n2656 4.5005
R2823 DVDD.n6924 DVDD.n2668 4.5005
R2824 DVDD.n6925 DVDD.n2657 4.5005
R2825 DVDD.n6925 DVDD.n2659 4.5005
R2826 DVDD.n6925 DVDD.n2656 4.5005
R2827 DVDD.n6925 DVDD.n6924 4.5005
R2828 DVDD.n2657 DVDD.n2655 4.5005
R2829 DVDD.n2659 DVDD.n2655 4.5005
R2830 DVDD.n6924 DVDD.n2655 4.5005
R2831 DVDD.n2726 DVDD.n2659 4.5005
R2832 DVDD.n6924 DVDD.n2726 4.5005
R2833 DVDD.n2667 DVDD.n2659 4.5005
R2834 DVDD.n6924 DVDD.n2667 4.5005
R2835 DVDD.n2729 DVDD.n2659 4.5005
R2836 DVDD.n6924 DVDD.n2729 4.5005
R2837 DVDD.n2666 DVDD.n2659 4.5005
R2838 DVDD.n6924 DVDD.n2666 4.5005
R2839 DVDD.n2732 DVDD.n2659 4.5005
R2840 DVDD.n6924 DVDD.n2732 4.5005
R2841 DVDD.n2665 DVDD.n2659 4.5005
R2842 DVDD.n2665 DVDD.n2656 4.5005
R2843 DVDD.n6924 DVDD.n2665 4.5005
R2844 DVDD.n2733 DVDD.n2659 4.5005
R2845 DVDD.n2733 DVDD.n2656 4.5005
R2846 DVDD.n6924 DVDD.n2733 4.5005
R2847 DVDD.n2664 DVDD.n2659 4.5005
R2848 DVDD.n2664 DVDD.n2656 4.5005
R2849 DVDD.n6924 DVDD.n2664 4.5005
R2850 DVDD.n2734 DVDD.n2657 4.5005
R2851 DVDD.n2734 DVDD.n2659 4.5005
R2852 DVDD.n2734 DVDD.n2656 4.5005
R2853 DVDD.n6924 DVDD.n2734 4.5005
R2854 DVDD.n2663 DVDD.n2657 4.5005
R2855 DVDD.n2663 DVDD.n2659 4.5005
R2856 DVDD.n2663 DVDD.n2656 4.5005
R2857 DVDD.n6924 DVDD.n2663 4.5005
R2858 DVDD.n2735 DVDD.n2657 4.5005
R2859 DVDD.n2735 DVDD.n2659 4.5005
R2860 DVDD.n2735 DVDD.n2656 4.5005
R2861 DVDD.n6924 DVDD.n2735 4.5005
R2862 DVDD.n2662 DVDD.n2659 4.5005
R2863 DVDD.n2662 DVDD.n2656 4.5005
R2864 DVDD.n6924 DVDD.n2662 4.5005
R2865 DVDD.n2736 DVDD.n2659 4.5005
R2866 DVDD.n2736 DVDD.n2656 4.5005
R2867 DVDD.n6924 DVDD.n2736 4.5005
R2868 DVDD.n2661 DVDD.n2659 4.5005
R2869 DVDD.n2661 DVDD.n2656 4.5005
R2870 DVDD.n6924 DVDD.n2661 4.5005
R2871 DVDD.n6923 DVDD.n2659 4.5005
R2872 DVDD.n6923 DVDD.n2656 4.5005
R2873 DVDD.n6924 DVDD.n6923 4.5005
R2874 DVDD.n6900 DVDD.n2743 4.5005
R2875 DVDD.n6900 DVDD.n2777 4.5005
R2876 DVDD.n2777 DVDD.n2742 4.5005
R2877 DVDD.n6873 DVDD.n2743 4.5005
R2878 DVDD.n6861 DVDD.n2777 4.5005
R2879 DVDD.n2798 DVDD.n2777 4.5005
R2880 DVDD.n6866 DVDD.n2777 4.5005
R2881 DVDD.n2819 DVDD.n2805 4.5005
R2882 DVDD.n2819 DVDD.n2807 4.5005
R2883 DVDD.n2819 DVDD.n2804 4.5005
R2884 DVDD.n6856 DVDD.n2819 4.5005
R2885 DVDD.n2821 DVDD.n2805 4.5005
R2886 DVDD.n2821 DVDD.n2807 4.5005
R2887 DVDD.n2821 DVDD.n2804 4.5005
R2888 DVDD.n6856 DVDD.n2821 4.5005
R2889 DVDD.n2818 DVDD.n2807 4.5005
R2890 DVDD.n2818 DVDD.n2804 4.5005
R2891 DVDD.n6856 DVDD.n2818 4.5005
R2892 DVDD.n2822 DVDD.n2807 4.5005
R2893 DVDD.n2822 DVDD.n2804 4.5005
R2894 DVDD.n6856 DVDD.n2822 4.5005
R2895 DVDD.n2817 DVDD.n2807 4.5005
R2896 DVDD.n2817 DVDD.n2804 4.5005
R2897 DVDD.n6856 DVDD.n2817 4.5005
R2898 DVDD.n2823 DVDD.n2805 4.5005
R2899 DVDD.n2823 DVDD.n2807 4.5005
R2900 DVDD.n2823 DVDD.n2804 4.5005
R2901 DVDD.n6856 DVDD.n2823 4.5005
R2902 DVDD.n2816 DVDD.n2805 4.5005
R2903 DVDD.n2816 DVDD.n2807 4.5005
R2904 DVDD.n2816 DVDD.n2804 4.5005
R2905 DVDD.n6856 DVDD.n2816 4.5005
R2906 DVDD.n2824 DVDD.n2805 4.5005
R2907 DVDD.n2824 DVDD.n2807 4.5005
R2908 DVDD.n2824 DVDD.n2804 4.5005
R2909 DVDD.n6856 DVDD.n2824 4.5005
R2910 DVDD.n2815 DVDD.n2805 4.5005
R2911 DVDD.n2815 DVDD.n2807 4.5005
R2912 DVDD.n2815 DVDD.n2804 4.5005
R2913 DVDD.n6856 DVDD.n2815 4.5005
R2914 DVDD.n2825 DVDD.n2807 4.5005
R2915 DVDD.n2825 DVDD.n2804 4.5005
R2916 DVDD.n6856 DVDD.n2825 4.5005
R2917 DVDD.n2814 DVDD.n2807 4.5005
R2918 DVDD.n2814 DVDD.n2804 4.5005
R2919 DVDD.n6856 DVDD.n2814 4.5005
R2920 DVDD.n2826 DVDD.n2807 4.5005
R2921 DVDD.n2826 DVDD.n2804 4.5005
R2922 DVDD.n6856 DVDD.n2826 4.5005
R2923 DVDD.n2813 DVDD.n2805 4.5005
R2924 DVDD.n2813 DVDD.n2807 4.5005
R2925 DVDD.n2813 DVDD.n2804 4.5005
R2926 DVDD.n6856 DVDD.n2813 4.5005
R2927 DVDD.n2827 DVDD.n2805 4.5005
R2928 DVDD.n2827 DVDD.n2807 4.5005
R2929 DVDD.n2827 DVDD.n2804 4.5005
R2930 DVDD.n6856 DVDD.n2827 4.5005
R2931 DVDD.n2812 DVDD.n2805 4.5005
R2932 DVDD.n2812 DVDD.n2807 4.5005
R2933 DVDD.n2812 DVDD.n2804 4.5005
R2934 DVDD.n6856 DVDD.n2812 4.5005
R2935 DVDD.n2828 DVDD.n2805 4.5005
R2936 DVDD.n2828 DVDD.n2807 4.5005
R2937 DVDD.n2828 DVDD.n2804 4.5005
R2938 DVDD.n6856 DVDD.n2828 4.5005
R2939 DVDD.n2811 DVDD.n2807 4.5005
R2940 DVDD.n2811 DVDD.n2804 4.5005
R2941 DVDD.n6856 DVDD.n2811 4.5005
R2942 DVDD.n2875 DVDD.n2807 4.5005
R2943 DVDD.n2875 DVDD.n2804 4.5005
R2944 DVDD.n6856 DVDD.n2875 4.5005
R2945 DVDD.n2810 DVDD.n2807 4.5005
R2946 DVDD.n2810 DVDD.n2804 4.5005
R2947 DVDD.n6856 DVDD.n2810 4.5005
R2948 DVDD.n6857 DVDD.n2805 4.5005
R2949 DVDD.n6857 DVDD.n2807 4.5005
R2950 DVDD.n6857 DVDD.n2804 4.5005
R2951 DVDD.n6857 DVDD.n6856 4.5005
R2952 DVDD.n2805 DVDD.n2803 4.5005
R2953 DVDD.n2807 DVDD.n2803 4.5005
R2954 DVDD.n6856 DVDD.n2803 4.5005
R2955 DVDD.n2878 DVDD.n2807 4.5005
R2956 DVDD.n6856 DVDD.n2878 4.5005
R2957 DVDD.n2809 DVDD.n2807 4.5005
R2958 DVDD.n6856 DVDD.n2809 4.5005
R2959 DVDD.n6855 DVDD.n2805 4.5005
R2960 DVDD.n6855 DVDD.n2807 4.5005
R2961 DVDD.n6856 DVDD.n6855 4.5005
R2962 DVDD.n2810 DVDD.n2805 4.5005
R2963 DVDD.n2875 DVDD.n2805 4.5005
R2964 DVDD.n2811 DVDD.n2805 4.5005
R2965 DVDD.n2826 DVDD.n2805 4.5005
R2966 DVDD.n2814 DVDD.n2805 4.5005
R2967 DVDD.n2825 DVDD.n2805 4.5005
R2968 DVDD.n2817 DVDD.n2805 4.5005
R2969 DVDD.n2822 DVDD.n2805 4.5005
R2970 DVDD.n2818 DVDD.n2805 4.5005
R2971 DVDD.n6866 DVDD.n2743 4.5005
R2972 DVDD.n2798 DVDD.n2743 4.5005
R2973 DVDD.n6861 DVDD.n2743 4.5005
R2974 DVDD.n6923 DVDD.n2657 4.5005
R2975 DVDD.n2661 DVDD.n2657 4.5005
R2976 DVDD.n2736 DVDD.n2657 4.5005
R2977 DVDD.n2662 DVDD.n2657 4.5005
R2978 DVDD.n2664 DVDD.n2657 4.5005
R2979 DVDD.n2733 DVDD.n2657 4.5005
R2980 DVDD.n2723 DVDD.n2657 4.5005
R2981 DVDD.n2669 DVDD.n2657 4.5005
R2982 DVDD.n2674 DVDD.n2657 4.5005
R2983 DVDD.n6985 DVDD.n2646 4.5005
R2984 DVDD.n6985 DVDD.n2633 4.5005
R2985 DVDD.n6985 DVDD.n2647 4.5005
R2986 DVDD.n6985 DVDD.n2632 4.5005
R2987 DVDD.n6985 DVDD.n2648 4.5005
R2988 DVDD.n6985 DVDD.n2631 4.5005
R2989 DVDD.n6985 DVDD.n6932 4.5005
R2990 DVDD.n6985 DVDD.n2630 4.5005
R2991 DVDD.n6934 DVDD.n2355 4.5005
R2992 DVDD.n6979 DVDD.n2355 4.5005
R2993 DVDD.n6982 DVDD.n2355 4.5005
R2994 DVDD.n2378 DVDD.n2374 4.5005
R2995 DVDD.n2378 DVDD.n2372 4.5005
R2996 DVDD.n7679 DVDD.n2378 4.5005
R2997 DVDD.n7660 DVDD.n2426 4.5005
R2998 DVDD.n2426 DVDD.n2374 4.5005
R2999 DVDD.n2426 DVDD.n2372 4.5005
R3000 DVDD.n7679 DVDD.n2426 4.5005
R3001 DVDD.n2377 DVDD.n2374 4.5005
R3002 DVDD.n2377 DVDD.n2372 4.5005
R3003 DVDD.n7679 DVDD.n2377 4.5005
R3004 DVDD.n7660 DVDD.n2449 4.5005
R3005 DVDD.n2449 DVDD.n2374 4.5005
R3006 DVDD.n2449 DVDD.n2372 4.5005
R3007 DVDD.n7679 DVDD.n2449 4.5005
R3008 DVDD.n2376 DVDD.n2374 4.5005
R3009 DVDD.n2376 DVDD.n2372 4.5005
R3010 DVDD.n7679 DVDD.n2376 4.5005
R3011 DVDD.n7678 DVDD.n7660 4.5005
R3012 DVDD.n7678 DVDD.n2374 4.5005
R3013 DVDD.n7678 DVDD.n2372 4.5005
R3014 DVDD.n7679 DVDD.n7678 4.5005
R3015 DVDD.n8357 DVDD.n1529 4.5005
R3016 DVDD.n8357 DVDD.n1530 4.5005
R3017 DVDD.n8358 DVDD.n8357 4.5005
R3018 DVDD.n8357 DVDD.n8356 4.5005
R3019 DVDD.n7683 DVDD.n7682 4.5005
R3020 DVDD.n7684 DVDD.n7683 4.5005
R3021 DVDD.n7686 DVDD.n2353 4.5005
R3022 DVDD.n7682 DVDD.n2353 4.5005
R3023 DVDD.n7684 DVDD.n2353 4.5005
R3024 DVDD.n7686 DVDD.n7685 4.5005
R3025 DVDD.n7685 DVDD.n7684 4.5005
R3026 DVDD.n6927 DVDD.n6926 4.5005
R3027 DVDD.n6929 DVDD.n6928 4.5005
R3028 DVDD.n6931 DVDD.n6930 4.5005
R3029 DVDD.n2650 DVDD.n2649 4.5005
R3030 DVDD.n2679 DVDD.n2678 4.5005
R3031 DVDD.n2681 DVDD.n2680 4.5005
R3032 DVDD.n2683 DVDD.n2682 4.5005
R3033 DVDD.n2685 DVDD.n2684 4.5005
R3034 DVDD.n2687 DVDD.n2686 4.5005
R3035 DVDD.n2689 DVDD.n2688 4.5005
R3036 DVDD.n2691 DVDD.n2690 4.5005
R3037 DVDD.n2693 DVDD.n2692 4.5005
R3038 DVDD.n2695 DVDD.n2694 4.5005
R3039 DVDD.n2697 DVDD.n2696 4.5005
R3040 DVDD.n2699 DVDD.n2698 4.5005
R3041 DVDD.n2701 DVDD.n2700 4.5005
R3042 DVDD.n2703 DVDD.n2702 4.5005
R3043 DVDD.n2705 DVDD.n2704 4.5005
R3044 DVDD.n2707 DVDD.n2706 4.5005
R3045 DVDD.n2708 DVDD.n2677 4.5005
R3046 DVDD.n2710 DVDD.n2709 4.5005
R3047 DVDD.n2712 DVDD.n2711 4.5005
R3048 DVDD.n2714 DVDD.n2713 4.5005
R3049 DVDD.n2716 DVDD.n2715 4.5005
R3050 DVDD.n2718 DVDD.n2717 4.5005
R3051 DVDD.n2720 DVDD.n2719 4.5005
R3052 DVDD.n2722 DVDD.n2721 4.5005
R3053 DVDD.n2676 DVDD.n2675 4.5005
R3054 DVDD.n2658 DVDD.n2654 4.5005
R3055 DVDD.n6902 DVDD.n6901 4.5005
R3056 DVDD.n6904 DVDD.n6903 4.5005
R3057 DVDD.n6906 DVDD.n6905 4.5005
R3058 DVDD.n6908 DVDD.n6907 4.5005
R3059 DVDD.n6910 DVDD.n6909 4.5005
R3060 DVDD.n6912 DVDD.n6911 4.5005
R3061 DVDD.n6914 DVDD.n6913 4.5005
R3062 DVDD.n6916 DVDD.n6915 4.5005
R3063 DVDD.n6918 DVDD.n6917 4.5005
R3064 DVDD.n6920 DVDD.n6919 4.5005
R3065 DVDD.n6922 DVDD.n6921 4.5005
R3066 DVDD.n2738 DVDD.n2737 4.5005
R3067 DVDD.n2752 DVDD.n2751 4.5005
R3068 DVDD.n2754 DVDD.n2753 4.5005
R3069 DVDD.n2755 DVDD.n2750 4.5005
R3070 DVDD.n2757 DVDD.n2756 4.5005
R3071 DVDD.n2758 DVDD.n2749 4.5005
R3072 DVDD.n2760 DVDD.n2759 4.5005
R3073 DVDD.n2761 DVDD.n2748 4.5005
R3074 DVDD.n2763 DVDD.n2762 4.5005
R3075 DVDD.n2764 DVDD.n2747 4.5005
R3076 DVDD.n2766 DVDD.n2765 4.5005
R3077 DVDD.n2767 DVDD.n2746 4.5005
R3078 DVDD.n2769 DVDD.n2768 4.5005
R3079 DVDD.n2770 DVDD.n2745 4.5005
R3080 DVDD.n2772 DVDD.n2771 4.5005
R3081 DVDD.n2773 DVDD.n2744 4.5005
R3082 DVDD.n2775 DVDD.n2774 4.5005
R3083 DVDD.n2776 DVDD.n2741 4.5005
R3084 DVDD.n6859 DVDD.n6858 4.5005
R3085 DVDD.n6860 DVDD.n2792 4.5005
R3086 DVDD.n6863 DVDD.n6862 4.5005
R3087 DVDD.n6865 DVDD.n6864 4.5005
R3088 DVDD.n2799 DVDD.n2797 4.5005
R3089 DVDD.n2832 DVDD.n2831 4.5005
R3090 DVDD.n2834 DVDD.n2833 4.5005
R3091 DVDD.n2836 DVDD.n2835 4.5005
R3092 DVDD.n2838 DVDD.n2837 4.5005
R3093 DVDD.n2840 DVDD.n2839 4.5005
R3094 DVDD.n2842 DVDD.n2841 4.5005
R3095 DVDD.n2844 DVDD.n2843 4.5005
R3096 DVDD.n2846 DVDD.n2845 4.5005
R3097 DVDD.n2848 DVDD.n2847 4.5005
R3098 DVDD.n2850 DVDD.n2849 4.5005
R3099 DVDD.n2852 DVDD.n2851 4.5005
R3100 DVDD.n2854 DVDD.n2853 4.5005
R3101 DVDD.n2856 DVDD.n2855 4.5005
R3102 DVDD.n2858 DVDD.n2857 4.5005
R3103 DVDD.n2860 DVDD.n2859 4.5005
R3104 DVDD.n2862 DVDD.n2861 4.5005
R3105 DVDD.n2864 DVDD.n2863 4.5005
R3106 DVDD.n2866 DVDD.n2865 4.5005
R3107 DVDD.n2868 DVDD.n2867 4.5005
R3108 DVDD.n2870 DVDD.n2869 4.5005
R3109 DVDD.n2872 DVDD.n2871 4.5005
R3110 DVDD.n2874 DVDD.n2873 4.5005
R3111 DVDD.n2830 DVDD.n2829 4.5005
R3112 DVDD.n2806 DVDD.n2802 4.5005
R3113 DVDD.n6851 DVDD.n6850 4.5005
R3114 DVDD.n6853 DVDD.n6852 4.5005
R3115 DVDD.n2880 DVDD.n2879 4.5005
R3116 DVDD.n6812 DVDD.n6811 4.5005
R3117 DVDD.n6813 DVDD.n6810 4.5005
R3118 DVDD.n6815 DVDD.n6814 4.5005
R3119 DVDD.n6816 DVDD.n6809 4.5005
R3120 DVDD.n6818 DVDD.n6817 4.5005
R3121 DVDD.n6819 DVDD.n6808 4.5005
R3122 DVDD.n6821 DVDD.n6820 4.5005
R3123 DVDD.n6822 DVDD.n6807 4.5005
R3124 DVDD.n6824 DVDD.n6823 4.5005
R3125 DVDD.n6825 DVDD.n6806 4.5005
R3126 DVDD.n6827 DVDD.n6826 4.5005
R3127 DVDD.n6828 DVDD.n6805 4.5005
R3128 DVDD.n6830 DVDD.n6829 4.5005
R3129 DVDD.n6831 DVDD.n6804 4.5005
R3130 DVDD.n6833 DVDD.n6832 4.5005
R3131 DVDD.n6834 DVDD.n6803 4.5005
R3132 DVDD.n6836 DVDD.n6835 4.5005
R3133 DVDD.n6837 DVDD.n6802 4.5005
R3134 DVDD.n6839 DVDD.n6838 4.5005
R3135 DVDD.n6840 DVDD.n6801 4.5005
R3136 DVDD.n6842 DVDD.n6841 4.5005
R3137 DVDD.n6843 DVDD.n6800 4.5005
R3138 DVDD.n6845 DVDD.n6844 4.5005
R3139 DVDD.n6846 DVDD.n6799 4.5005
R3140 DVDD.n6848 DVDD.n6847 4.5005
R3141 DVDD.n6849 DVDD.n2883 4.5005
R3142 DVDD.n6796 DVDD.n6795 4.5005
R3143 DVDD.n6798 DVDD.n6797 4.5005
R3144 DVDD.n2885 DVDD.n2884 4.5005
R3145 DVDD.n2927 DVDD.n2926 4.5005
R3146 DVDD.n2929 DVDD.n2928 4.5005
R3147 DVDD.n2930 DVDD.n2925 4.5005
R3148 DVDD.n2932 DVDD.n2931 4.5005
R3149 DVDD.n2933 DVDD.n2924 4.5005
R3150 DVDD.n2935 DVDD.n2934 4.5005
R3151 DVDD.n2936 DVDD.n2923 4.5005
R3152 DVDD.n2938 DVDD.n2937 4.5005
R3153 DVDD.n2939 DVDD.n2922 4.5005
R3154 DVDD.n2941 DVDD.n2940 4.5005
R3155 DVDD.n2942 DVDD.n2921 4.5005
R3156 DVDD.n2944 DVDD.n2943 4.5005
R3157 DVDD.n2945 DVDD.n2920 4.5005
R3158 DVDD.n2947 DVDD.n2946 4.5005
R3159 DVDD.n2948 DVDD.n2919 4.5005
R3160 DVDD.n2950 DVDD.n2949 4.5005
R3161 DVDD.n2951 DVDD.n2918 4.5005
R3162 DVDD.n2953 DVDD.n2952 4.5005
R3163 DVDD.n2954 DVDD.n2917 4.5005
R3164 DVDD.n2956 DVDD.n2955 4.5005
R3165 DVDD.n2905 DVDD.n2903 4.5005
R3166 DVDD.n6783 DVDD.n6782 4.5005
R3167 DVDD.n6784 DVDD.n2901 4.5005
R3168 DVDD.n6786 DVDD.n6785 4.5005
R3169 DVDD.n2902 DVDD.n2892 4.5005
R3170 DVDD.n6793 DVDD.n2888 4.5005
R3171 DVDD.n9302 DVDD.n445 4.5005
R3172 DVDD.n9409 DVDD.n391 4.5005
R3173 DVDD.n9411 DVDD.n9410 4.5005
R3174 DVDD.n9413 DVDD.n9412 4.5005
R3175 DVDD.n390 DVDD.n387 4.5005
R3176 DVDD.n9397 DVDD.n9396 4.5005
R3177 DVDD.n9395 DVDD.n401 4.5005
R3178 DVDD.n9394 DVDD.n9393 4.5005
R3179 DVDD.n403 DVDD.n173 4.5005
R3180 DVDD.n402 DVDD.n172 4.5005
R3181 DVDD.n165 DVDD.n163 4.5005
R3182 DVDD.n9592 DVDD.n9591 4.5005
R3183 DVDD.n9594 DVDD.n9593 4.5005
R3184 DVDD.n162 DVDD.n154 4.5005
R3185 DVDD.n161 DVDD.n160 4.5005
R3186 DVDD.n159 DVDD.n143 4.5005
R3187 DVDD.n158 DVDD.n142 4.5005
R3188 DVDD.n157 DVDD.n136 4.5005
R3189 DVDD.n9607 DVDD.n135 4.5005
R3190 DVDD.n9609 DVDD.n9608 4.5005
R3191 DVDD.n9611 DVDD.n9610 4.5005
R3192 DVDD.n134 DVDD.n131 4.5005
R3193 DVDD.n9308 DVDD.n411 4.5005
R3194 DVDD.n9309 DVDD.n410 4.5005
R3195 DVDD.n9311 DVDD.n9310 4.5005
R3196 DVDD.n9307 DVDD.n443 4.5005
R3197 DVDD.n9306 DVDD.n437 4.5005
R3198 DVDD.n9305 DVDD.n436 4.5005
R3199 DVDD.n9304 DVDD.n9303 4.5005
R3200 DVDD.n9299 DVDD.n9298 4.5005
R3201 DVDD.n9301 DVDD.n9300 4.5005
R3202 DVDD.n447 DVDD.n446 4.5005
R3203 DVDD.n9269 DVDD.n9268 4.5005
R3204 DVDD.n9271 DVDD.n9270 4.5005
R3205 DVDD.n9272 DVDD.n9267 4.5005
R3206 DVDD.n9274 DVDD.n9273 4.5005
R3207 DVDD.n9275 DVDD.n9266 4.5005
R3208 DVDD.n9277 DVDD.n9276 4.5005
R3209 DVDD.n9279 DVDD.n9278 4.5005
R3210 DVDD.n9280 DVDD.n9250 4.5005
R3211 DVDD.n9282 DVDD.n9281 4.5005
R3212 DVDD.n9265 DVDD.n9249 4.5005
R3213 DVDD.n9264 DVDD.n9263 4.5005
R3214 DVDD.n9262 DVDD.n9261 4.5005
R3215 DVDD.n9260 DVDD.n9259 4.5005
R3216 DVDD.n9258 DVDD.n9257 4.5005
R3217 DVDD.n9256 DVDD.n9255 4.5005
R3218 DVDD.n9254 DVDD.n9253 4.5005
R3219 DVDD.n9252 DVDD.n9251 4.5005
R3220 DVDD.n458 DVDD.n455 4.5005
R3221 DVDD.n9287 DVDD.n9286 4.5005
R3222 DVDD.n9288 DVDD.n454 4.5005
R3223 DVDD.n9290 DVDD.n9289 4.5005
R3224 DVDD.n9291 DVDD.n453 4.5005
R3225 DVDD.n9293 DVDD.n9292 4.5005
R3226 DVDD.n9294 DVDD.n452 4.5005
R3227 DVDD.n9296 DVDD.n9295 4.5005
R3228 DVDD.n9297 DVDD.n450 4.5005
R3229 DVDD.n5216 DVDD.n5215 4.5005
R3230 DVDD.n4562 DVDD.n451 4.5005
R3231 DVDD.n5175 DVDD.n5174 4.5005
R3232 DVDD.n5177 DVDD.n5176 4.5005
R3233 DVDD.n5178 DVDD.n5173 4.5005
R3234 DVDD.n5180 DVDD.n5179 4.5005
R3235 DVDD.n5181 DVDD.n5172 4.5005
R3236 DVDD.n5183 DVDD.n5182 4.5005
R3237 DVDD.n5184 DVDD.n5171 4.5005
R3238 DVDD.n5186 DVDD.n5185 4.5005
R3239 DVDD.n5187 DVDD.n5170 4.5005
R3240 DVDD.n5189 DVDD.n5188 4.5005
R3241 DVDD.n5190 DVDD.n5169 4.5005
R3242 DVDD.n5192 DVDD.n5191 4.5005
R3243 DVDD.n5193 DVDD.n5168 4.5005
R3244 DVDD.n5195 DVDD.n5194 4.5005
R3245 DVDD.n5196 DVDD.n5167 4.5005
R3246 DVDD.n5198 DVDD.n5197 4.5005
R3247 DVDD.n5199 DVDD.n5166 4.5005
R3248 DVDD.n5201 DVDD.n5200 4.5005
R3249 DVDD.n5202 DVDD.n5165 4.5005
R3250 DVDD.n5204 DVDD.n5203 4.5005
R3251 DVDD.n5205 DVDD.n5164 4.5005
R3252 DVDD.n5207 DVDD.n5206 4.5005
R3253 DVDD.n5208 DVDD.n5163 4.5005
R3254 DVDD.n5210 DVDD.n5209 4.5005
R3255 DVDD.n5211 DVDD.n5162 4.5005
R3256 DVDD.n5213 DVDD.n5212 4.5005
R3257 DVDD.n5214 DVDD.n4564 4.5005
R3258 DVDD.n5161 DVDD.n5160 4.5005
R3259 DVDD.n4566 DVDD.n4565 4.5005
R3260 DVDD.n5138 DVDD.n5137 4.5005
R3261 DVDD.n5139 DVDD.n5136 4.5005
R3262 DVDD.n5141 DVDD.n5140 4.5005
R3263 DVDD.n5142 DVDD.n5135 4.5005
R3264 DVDD.n5144 DVDD.n5143 4.5005
R3265 DVDD.n5145 DVDD.n5134 4.5005
R3266 DVDD.n5147 DVDD.n5146 4.5005
R3267 DVDD.n5149 DVDD.n5148 4.5005
R3268 DVDD.n5151 DVDD.n5150 4.5005
R3269 DVDD.n5153 DVDD.n5152 4.5005
R3270 DVDD.n5155 DVDD.n5154 4.5005
R3271 DVDD.n5133 DVDD.n5120 4.5005
R3272 DVDD.n5132 DVDD.n5131 4.5005
R3273 DVDD.n5130 DVDD.n5129 4.5005
R3274 DVDD.n5128 DVDD.n5127 4.5005
R3275 DVDD.n5126 DVDD.n5125 4.5005
R3276 DVDD.n5124 DVDD.n5123 4.5005
R3277 DVDD.n5122 DVDD.n5121 4.5005
R3278 DVDD.n4572 DVDD.n4569 4.5005
R3279 DVDD.n1401 DVDD.n1400 4.5005
R3280 DVDD.n8546 DVDD.n1401 4.5005
R3281 DVDD.n8548 DVDD.n8547 4.5005
R3282 DVDD.n8547 DVDD.n8546 4.5005
R3283 DVDD.n8419 DVDD.n8418 4.5005
R3284 DVDD.n8420 DVDD.n8419 4.5005
R3285 DVDD.n7349 DVDD.n1506 4.5005
R3286 DVDD.n7352 DVDD.n1506 4.5005
R3287 DVDD.n1497 DVDD.n1462 4.5005
R3288 DVDD.n7352 DVDD.n1462 4.5005
R3289 DVDD.n8420 DVDD.n1461 4.5005
R3290 DVDD.n8418 DVDD.n1461 4.5005
R3291 DVDD.n8416 DVDD.n1461 4.5005
R3292 DVDD.n8418 DVDD.n8417 4.5005
R3293 DVDD.n8417 DVDD.n8416 4.5005
R3294 DVDD.n1488 DVDD.n1487 4.5005
R3295 DVDD.n1488 DVDD.n1415 4.5005
R3296 DVDD.n1471 DVDD.n1415 4.5005
R3297 DVDD.n1487 DVDD.n1471 4.5005
R3298 DVDD.n1485 DVDD.n1471 4.5005
R3299 DVDD.n1487 DVDD.n1486 4.5005
R3300 DVDD.n1486 DVDD.n1485 4.5005
R3301 DVDD.n1483 DVDD.n1482 4.5005
R3302 DVDD.n1483 DVDD.n1409 4.5005
R3303 DVDD.n1477 DVDD.n1409 4.5005
R3304 DVDD.n1482 DVDD.n1477 4.5005
R3305 DVDD.n1477 DVDD.n1393 4.5005
R3306 DVDD.n1482 DVDD.n1481 4.5005
R3307 DVDD.n1481 DVDD.n1393 4.5005
R3308 DVDD.n8360 DVDD.n1512 4.5005
R3309 DVDD.n8360 DVDD.n1513 4.5005
R3310 DVDD.n8365 DVDD.n8360 4.5005
R3311 DVDD.n8361 DVDD.n1512 4.5005
R3312 DVDD.n8361 DVDD.n1513 4.5005
R3313 DVDD.n1522 DVDD.n1513 4.5005
R3314 DVDD.n8369 DVDD.n1522 4.5005
R3315 DVDD.n1518 DVDD.n1513 4.5005
R3316 DVDD.n8369 DVDD.n1518 4.5005
R3317 DVDD.n1524 DVDD.n1513 4.5005
R3318 DVDD.n8369 DVDD.n1524 4.5005
R3319 DVDD.n1517 DVDD.n1513 4.5005
R3320 DVDD.n8369 DVDD.n1517 4.5005
R3321 DVDD.n1526 DVDD.n1513 4.5005
R3322 DVDD.n8369 DVDD.n1526 4.5005
R3323 DVDD.n1516 DVDD.n1513 4.5005
R3324 DVDD.n8369 DVDD.n1516 4.5005
R3325 DVDD.n8368 DVDD.n1513 4.5005
R3326 DVDD.n8369 DVDD.n8368 4.5005
R3327 DVDD.n1515 DVDD.n1513 4.5005
R3328 DVDD.n8369 DVDD.n1515 4.5005
R3329 DVDD.n8370 DVDD.n1512 4.5005
R3330 DVDD.n8370 DVDD.n1513 4.5005
R3331 DVDD.n8370 DVDD.n8369 4.5005
R3332 DVDD.n8288 DVDD.n1703 4.5005
R3333 DVDD.n8288 DVDD.n1704 4.5005
R3334 DVDD.n8288 DVDD.n8287 4.5005
R3335 DVDD.n1711 DVDD.n1704 4.5005
R3336 DVDD.n8287 DVDD.n1711 4.5005
R3337 DVDD.n1714 DVDD.n1704 4.5005
R3338 DVDD.n8287 DVDD.n1714 4.5005
R3339 DVDD.n1710 DVDD.n1704 4.5005
R3340 DVDD.n8287 DVDD.n1710 4.5005
R3341 DVDD.n1716 DVDD.n1704 4.5005
R3342 DVDD.n8287 DVDD.n1716 4.5005
R3343 DVDD.n1709 DVDD.n1704 4.5005
R3344 DVDD.n8287 DVDD.n1709 4.5005
R3345 DVDD.n1718 DVDD.n1704 4.5005
R3346 DVDD.n8287 DVDD.n1718 4.5005
R3347 DVDD.n1708 DVDD.n1704 4.5005
R3348 DVDD.n8287 DVDD.n1708 4.5005
R3349 DVDD.n8286 DVDD.n1704 4.5005
R3350 DVDD.n8287 DVDD.n8286 4.5005
R3351 DVDD.n1707 DVDD.n1704 4.5005
R3352 DVDD.n8287 DVDD.n1707 4.5005
R3353 DVDD.n1704 DVDD.n1309 4.5005
R3354 DVDD.n8284 DVDD.n1309 4.5005
R3355 DVDD.n8287 DVDD.n1309 4.5005
R3356 DVDD.n7506 DVDD.n7068 4.5005
R3357 DVDD.n7506 DVDD.n7069 4.5005
R3358 DVDD.n7506 DVDD.n7505 4.5005
R3359 DVDD.n7075 DVDD.n7069 4.5005
R3360 DVDD.n7505 DVDD.n7075 4.5005
R3361 DVDD.n7078 DVDD.n7069 4.5005
R3362 DVDD.n7505 DVDD.n7078 4.5005
R3363 DVDD.n7074 DVDD.n7069 4.5005
R3364 DVDD.n7505 DVDD.n7074 4.5005
R3365 DVDD.n7080 DVDD.n7069 4.5005
R3366 DVDD.n7505 DVDD.n7080 4.5005
R3367 DVDD.n7073 DVDD.n7069 4.5005
R3368 DVDD.n7505 DVDD.n7073 4.5005
R3369 DVDD.n7082 DVDD.n7069 4.5005
R3370 DVDD.n7505 DVDD.n7082 4.5005
R3371 DVDD.n7072 DVDD.n7069 4.5005
R3372 DVDD.n7505 DVDD.n7072 4.5005
R3373 DVDD.n7084 DVDD.n7069 4.5005
R3374 DVDD.n7505 DVDD.n7084 4.5005
R3375 DVDD.n7071 DVDD.n7069 4.5005
R3376 DVDD.n7505 DVDD.n7071 4.5005
R3377 DVDD.n7504 DVDD.n7069 4.5005
R3378 DVDD.n7504 DVDD.n7503 4.5005
R3379 DVDD.n7505 DVDD.n7504 4.5005
R3380 DVDD.n7425 DVDD.n1620 4.5005
R3381 DVDD.n7428 DVDD.n1620 4.5005
R3382 DVDD.n7333 DVDD.n1620 4.5005
R3383 DVDD.n7428 DVDD.n7368 4.5005
R3384 DVDD.n7368 DVDD.n7333 4.5005
R3385 DVDD.n7428 DVDD.n7370 4.5005
R3386 DVDD.n7370 DVDD.n7333 4.5005
R3387 DVDD.n7428 DVDD.n7367 4.5005
R3388 DVDD.n7367 DVDD.n7333 4.5005
R3389 DVDD.n7428 DVDD.n7371 4.5005
R3390 DVDD.n7371 DVDD.n7333 4.5005
R3391 DVDD.n7428 DVDD.n7366 4.5005
R3392 DVDD.n7366 DVDD.n7333 4.5005
R3393 DVDD.n7428 DVDD.n7372 4.5005
R3394 DVDD.n7372 DVDD.n7333 4.5005
R3395 DVDD.n7428 DVDD.n7365 4.5005
R3396 DVDD.n7365 DVDD.n7333 4.5005
R3397 DVDD.n7428 DVDD.n7427 4.5005
R3398 DVDD.n7427 DVDD.n7333 4.5005
R3399 DVDD.n7428 DVDD.n7364 4.5005
R3400 DVDD.n7364 DVDD.n7333 4.5005
R3401 DVDD.n7429 DVDD.n7428 4.5005
R3402 DVDD.n7430 DVDD.n7429 4.5005
R3403 DVDD.n7429 DVDD.n7333 4.5005
R3404 DVDD.n1763 DVDD.n1747 4.5005
R3405 DVDD.n8250 DVDD.n1747 4.5005
R3406 DVDD.n8252 DVDD.n1747 4.5005
R3407 DVDD.n8250 DVDD.n1745 4.5005
R3408 DVDD.n8252 DVDD.n1745 4.5005
R3409 DVDD.n8250 DVDD.n1748 4.5005
R3410 DVDD.n8252 DVDD.n1748 4.5005
R3411 DVDD.n8250 DVDD.n1744 4.5005
R3412 DVDD.n8252 DVDD.n1744 4.5005
R3413 DVDD.n8250 DVDD.n1749 4.5005
R3414 DVDD.n8252 DVDD.n1749 4.5005
R3415 DVDD.n8250 DVDD.n1743 4.5005
R3416 DVDD.n8252 DVDD.n1743 4.5005
R3417 DVDD.n8250 DVDD.n1750 4.5005
R3418 DVDD.n8252 DVDD.n1750 4.5005
R3419 DVDD.n8250 DVDD.n1742 4.5005
R3420 DVDD.n8252 DVDD.n1742 4.5005
R3421 DVDD.n8251 DVDD.n8250 4.5005
R3422 DVDD.n8252 DVDD.n8251 4.5005
R3423 DVDD.n8250 DVDD.n1741 4.5005
R3424 DVDD.n8252 DVDD.n1741 4.5005
R3425 DVDD.n8250 DVDD.n1317 4.5005
R3426 DVDD.n1757 DVDD.n1317 4.5005
R3427 DVDD.n8252 DVDD.n1317 4.5005
R3428 DVDD.n8205 DVDD.n8193 4.5005
R3429 DVDD.n8208 DVDD.n8193 4.5005
R3430 DVDD.n8193 DVDD.n1784 4.5005
R3431 DVDD.n8208 DVDD.n1796 4.5005
R3432 DVDD.n1796 DVDD.n1784 4.5005
R3433 DVDD.n8208 DVDD.n8194 4.5005
R3434 DVDD.n8194 DVDD.n1784 4.5005
R3435 DVDD.n8208 DVDD.n1795 4.5005
R3436 DVDD.n1795 DVDD.n1784 4.5005
R3437 DVDD.n8208 DVDD.n8195 4.5005
R3438 DVDD.n8195 DVDD.n1784 4.5005
R3439 DVDD.n8208 DVDD.n1794 4.5005
R3440 DVDD.n1794 DVDD.n1784 4.5005
R3441 DVDD.n8208 DVDD.n8196 4.5005
R3442 DVDD.n8196 DVDD.n1784 4.5005
R3443 DVDD.n8208 DVDD.n1793 4.5005
R3444 DVDD.n1793 DVDD.n1784 4.5005
R3445 DVDD.n8208 DVDD.n8207 4.5005
R3446 DVDD.n8207 DVDD.n1784 4.5005
R3447 DVDD.n8208 DVDD.n1792 4.5005
R3448 DVDD.n1792 DVDD.n1784 4.5005
R3449 DVDD.n8209 DVDD.n8208 4.5005
R3450 DVDD.n8210 DVDD.n8209 4.5005
R3451 DVDD.n8209 DVDD.n1784 4.5005
R3452 DVDD.n1813 DVDD.n1799 4.5005
R3453 DVDD.n1813 DVDD.n1800 4.5005
R3454 DVDD.n8191 DVDD.n1813 4.5005
R3455 DVDD.n1816 DVDD.n1800 4.5005
R3456 DVDD.n8191 DVDD.n1816 4.5005
R3457 DVDD.n1812 DVDD.n1800 4.5005
R3458 DVDD.n8191 DVDD.n1812 4.5005
R3459 DVDD.n1818 DVDD.n1800 4.5005
R3460 DVDD.n8191 DVDD.n1818 4.5005
R3461 DVDD.n1811 DVDD.n1800 4.5005
R3462 DVDD.n8191 DVDD.n1811 4.5005
R3463 DVDD.n1820 DVDD.n1800 4.5005
R3464 DVDD.n8191 DVDD.n1820 4.5005
R3465 DVDD.n1810 DVDD.n1800 4.5005
R3466 DVDD.n8191 DVDD.n1810 4.5005
R3467 DVDD.n1822 DVDD.n1800 4.5005
R3468 DVDD.n8191 DVDD.n1822 4.5005
R3469 DVDD.n1809 DVDD.n1800 4.5005
R3470 DVDD.n8191 DVDD.n1809 4.5005
R3471 DVDD.n1824 DVDD.n1800 4.5005
R3472 DVDD.n8191 DVDD.n1824 4.5005
R3473 DVDD.n1808 DVDD.n1800 4.5005
R3474 DVDD.n8191 DVDD.n1808 4.5005
R3475 DVDD.n1826 DVDD.n1800 4.5005
R3476 DVDD.n8191 DVDD.n1826 4.5005
R3477 DVDD.n1807 DVDD.n1800 4.5005
R3478 DVDD.n8191 DVDD.n1807 4.5005
R3479 DVDD.n1828 DVDD.n1800 4.5005
R3480 DVDD.n8191 DVDD.n1828 4.5005
R3481 DVDD.n1806 DVDD.n1800 4.5005
R3482 DVDD.n8191 DVDD.n1806 4.5005
R3483 DVDD.n1830 DVDD.n1800 4.5005
R3484 DVDD.n8191 DVDD.n1830 4.5005
R3485 DVDD.n1805 DVDD.n1800 4.5005
R3486 DVDD.n8191 DVDD.n1805 4.5005
R3487 DVDD.n1832 DVDD.n1800 4.5005
R3488 DVDD.n8191 DVDD.n1832 4.5005
R3489 DVDD.n1804 DVDD.n1800 4.5005
R3490 DVDD.n8191 DVDD.n1804 4.5005
R3491 DVDD.n1834 DVDD.n1800 4.5005
R3492 DVDD.n8191 DVDD.n1834 4.5005
R3493 DVDD.n1803 DVDD.n1800 4.5005
R3494 DVDD.n8191 DVDD.n1803 4.5005
R3495 DVDD.n8190 DVDD.n1800 4.5005
R3496 DVDD.n8191 DVDD.n8190 4.5005
R3497 DVDD.n1802 DVDD.n1800 4.5005
R3498 DVDD.n8191 DVDD.n1802 4.5005
R3499 DVDD.n8192 DVDD.n1799 4.5005
R3500 DVDD.n8192 DVDD.n1800 4.5005
R3501 DVDD.n8192 DVDD.n8191 4.5005
R3502 DVDD.n7985 DVDD.n7960 4.5005
R3503 DVDD.n8008 DVDD.n7960 4.5005
R3504 DVDD.n8010 DVDD.n7960 4.5005
R3505 DVDD.n8008 DVDD.n7962 4.5005
R3506 DVDD.n8010 DVDD.n7962 4.5005
R3507 DVDD.n8008 DVDD.n2026 4.5005
R3508 DVDD.n8010 DVDD.n2026 4.5005
R3509 DVDD.n8008 DVDD.n7963 4.5005
R3510 DVDD.n8010 DVDD.n7963 4.5005
R3511 DVDD.n8008 DVDD.n2025 4.5005
R3512 DVDD.n8010 DVDD.n2025 4.5005
R3513 DVDD.n8008 DVDD.n7964 4.5005
R3514 DVDD.n8010 DVDD.n7964 4.5005
R3515 DVDD.n8008 DVDD.n2024 4.5005
R3516 DVDD.n8010 DVDD.n2024 4.5005
R3517 DVDD.n8008 DVDD.n7965 4.5005
R3518 DVDD.n8010 DVDD.n7965 4.5005
R3519 DVDD.n8008 DVDD.n2023 4.5005
R3520 DVDD.n8010 DVDD.n2023 4.5005
R3521 DVDD.n8008 DVDD.n7966 4.5005
R3522 DVDD.n8010 DVDD.n7966 4.5005
R3523 DVDD.n8008 DVDD.n2022 4.5005
R3524 DVDD.n8010 DVDD.n2022 4.5005
R3525 DVDD.n8008 DVDD.n7967 4.5005
R3526 DVDD.n8010 DVDD.n7967 4.5005
R3527 DVDD.n8008 DVDD.n2021 4.5005
R3528 DVDD.n8010 DVDD.n2021 4.5005
R3529 DVDD.n8008 DVDD.n7968 4.5005
R3530 DVDD.n8010 DVDD.n7968 4.5005
R3531 DVDD.n8008 DVDD.n2020 4.5005
R3532 DVDD.n8010 DVDD.n2020 4.5005
R3533 DVDD.n8008 DVDD.n7969 4.5005
R3534 DVDD.n8010 DVDD.n7969 4.5005
R3535 DVDD.n8008 DVDD.n2019 4.5005
R3536 DVDD.n8010 DVDD.n2019 4.5005
R3537 DVDD.n8008 DVDD.n7970 4.5005
R3538 DVDD.n8010 DVDD.n7970 4.5005
R3539 DVDD.n8008 DVDD.n2018 4.5005
R3540 DVDD.n8010 DVDD.n2018 4.5005
R3541 DVDD.n8008 DVDD.n7971 4.5005
R3542 DVDD.n8010 DVDD.n7971 4.5005
R3543 DVDD.n8008 DVDD.n2017 4.5005
R3544 DVDD.n8010 DVDD.n2017 4.5005
R3545 DVDD.n8008 DVDD.n7972 4.5005
R3546 DVDD.n8010 DVDD.n7972 4.5005
R3547 DVDD.n8008 DVDD.n2016 4.5005
R3548 DVDD.n8010 DVDD.n2016 4.5005
R3549 DVDD.n8009 DVDD.n7985 4.5005
R3550 DVDD.n8009 DVDD.n8008 4.5005
R3551 DVDD.n8010 DVDD.n8009 4.5005
R3552 DVDD.n7958 DVDD.n2042 4.5005
R3553 DVDD.n7954 DVDD.n2042 4.5005
R3554 DVDD.n2042 DVDD.n2029 4.5005
R3555 DVDD.n2042 DVDD.n2028 4.5005
R3556 DVDD.n7958 DVDD.n2044 4.5005
R3557 DVDD.n7954 DVDD.n2044 4.5005
R3558 DVDD.n2044 DVDD.n2029 4.5005
R3559 DVDD.n2044 DVDD.n2028 4.5005
R3560 DVDD.n7958 DVDD.n2041 4.5005
R3561 DVDD.n7954 DVDD.n2041 4.5005
R3562 DVDD.n2041 DVDD.n2029 4.5005
R3563 DVDD.n2041 DVDD.n2028 4.5005
R3564 DVDD.n7958 DVDD.n2045 4.5005
R3565 DVDD.n7954 DVDD.n2045 4.5005
R3566 DVDD.n2045 DVDD.n2029 4.5005
R3567 DVDD.n2045 DVDD.n2028 4.5005
R3568 DVDD.n7958 DVDD.n2040 4.5005
R3569 DVDD.n7954 DVDD.n2040 4.5005
R3570 DVDD.n2040 DVDD.n2029 4.5005
R3571 DVDD.n2040 DVDD.n2028 4.5005
R3572 DVDD.n7958 DVDD.n2046 4.5005
R3573 DVDD.n7954 DVDD.n2046 4.5005
R3574 DVDD.n2046 DVDD.n2029 4.5005
R3575 DVDD.n2046 DVDD.n2028 4.5005
R3576 DVDD.n7958 DVDD.n2039 4.5005
R3577 DVDD.n7954 DVDD.n2039 4.5005
R3578 DVDD.n2039 DVDD.n2029 4.5005
R3579 DVDD.n2039 DVDD.n2028 4.5005
R3580 DVDD.n7958 DVDD.n2047 4.5005
R3581 DVDD.n7954 DVDD.n2047 4.5005
R3582 DVDD.n2047 DVDD.n2029 4.5005
R3583 DVDD.n2047 DVDD.n2028 4.5005
R3584 DVDD.n7958 DVDD.n2038 4.5005
R3585 DVDD.n7954 DVDD.n2038 4.5005
R3586 DVDD.n2038 DVDD.n2029 4.5005
R3587 DVDD.n2038 DVDD.n2028 4.5005
R3588 DVDD.n7958 DVDD.n2048 4.5005
R3589 DVDD.n7954 DVDD.n2048 4.5005
R3590 DVDD.n2048 DVDD.n2029 4.5005
R3591 DVDD.n2048 DVDD.n2028 4.5005
R3592 DVDD.n7958 DVDD.n2037 4.5005
R3593 DVDD.n7954 DVDD.n2037 4.5005
R3594 DVDD.n2037 DVDD.n2029 4.5005
R3595 DVDD.n2037 DVDD.n2028 4.5005
R3596 DVDD.n7958 DVDD.n2049 4.5005
R3597 DVDD.n7954 DVDD.n2049 4.5005
R3598 DVDD.n2049 DVDD.n2029 4.5005
R3599 DVDD.n2049 DVDD.n2028 4.5005
R3600 DVDD.n7958 DVDD.n2036 4.5005
R3601 DVDD.n7954 DVDD.n2036 4.5005
R3602 DVDD.n2036 DVDD.n2029 4.5005
R3603 DVDD.n2036 DVDD.n2028 4.5005
R3604 DVDD.n7958 DVDD.n2050 4.5005
R3605 DVDD.n7954 DVDD.n2050 4.5005
R3606 DVDD.n2050 DVDD.n2029 4.5005
R3607 DVDD.n2050 DVDD.n2028 4.5005
R3608 DVDD.n7958 DVDD.n2035 4.5005
R3609 DVDD.n7954 DVDD.n2035 4.5005
R3610 DVDD.n2035 DVDD.n2029 4.5005
R3611 DVDD.n2035 DVDD.n2028 4.5005
R3612 DVDD.n7958 DVDD.n2052 4.5005
R3613 DVDD.n7954 DVDD.n2052 4.5005
R3614 DVDD.n2052 DVDD.n2028 4.5005
R3615 DVDD.n2034 DVDD.n2028 4.5005
R3616 DVDD.n7958 DVDD.n2034 4.5005
R3617 DVDD.n2054 DVDD.n2029 4.5005
R3618 DVDD.n7958 DVDD.n2054 4.5005
R3619 DVDD.n2033 DVDD.n2029 4.5005
R3620 DVDD.n7958 DVDD.n2033 4.5005
R3621 DVDD.n2056 DVDD.n2029 4.5005
R3622 DVDD.n7958 DVDD.n2056 4.5005
R3623 DVDD.n2032 DVDD.n2029 4.5005
R3624 DVDD.n7958 DVDD.n2032 4.5005
R3625 DVDD.n7957 DVDD.n2029 4.5005
R3626 DVDD.n7958 DVDD.n7957 4.5005
R3627 DVDD.n2031 DVDD.n2029 4.5005
R3628 DVDD.n7958 DVDD.n2031 4.5005
R3629 DVDD.n7959 DVDD.n2028 4.5005
R3630 DVDD.n7959 DVDD.n2029 4.5005
R3631 DVDD.n7959 DVDD.n7958 4.5005
R3632 DVDD.n6485 DVDD.n3407 4.5005
R3633 DVDD.n6603 DVDD.n3407 4.5005
R3634 DVDD.n6481 DVDD.n3407 4.5005
R3635 DVDD.n6605 DVDD.n3407 4.5005
R3636 DVDD.n6485 DVDD.n3409 4.5005
R3637 DVDD.n6603 DVDD.n3409 4.5005
R3638 DVDD.n6481 DVDD.n3409 4.5005
R3639 DVDD.n6605 DVDD.n3409 4.5005
R3640 DVDD.n6485 DVDD.n3406 4.5005
R3641 DVDD.n6603 DVDD.n3406 4.5005
R3642 DVDD.n6481 DVDD.n3406 4.5005
R3643 DVDD.n6605 DVDD.n3406 4.5005
R3644 DVDD.n6485 DVDD.n3410 4.5005
R3645 DVDD.n6603 DVDD.n3410 4.5005
R3646 DVDD.n6481 DVDD.n3410 4.5005
R3647 DVDD.n6605 DVDD.n3410 4.5005
R3648 DVDD.n6485 DVDD.n3405 4.5005
R3649 DVDD.n6603 DVDD.n3405 4.5005
R3650 DVDD.n6481 DVDD.n3405 4.5005
R3651 DVDD.n6605 DVDD.n3405 4.5005
R3652 DVDD.n6485 DVDD.n3411 4.5005
R3653 DVDD.n6603 DVDD.n3411 4.5005
R3654 DVDD.n6481 DVDD.n3411 4.5005
R3655 DVDD.n6605 DVDD.n3411 4.5005
R3656 DVDD.n6485 DVDD.n3404 4.5005
R3657 DVDD.n6603 DVDD.n3404 4.5005
R3658 DVDD.n6481 DVDD.n3404 4.5005
R3659 DVDD.n6605 DVDD.n3404 4.5005
R3660 DVDD.n6485 DVDD.n3412 4.5005
R3661 DVDD.n6603 DVDD.n3412 4.5005
R3662 DVDD.n6481 DVDD.n3412 4.5005
R3663 DVDD.n6605 DVDD.n3412 4.5005
R3664 DVDD.n6485 DVDD.n3403 4.5005
R3665 DVDD.n6603 DVDD.n3403 4.5005
R3666 DVDD.n6481 DVDD.n3403 4.5005
R3667 DVDD.n6605 DVDD.n3403 4.5005
R3668 DVDD.n6485 DVDD.n6470 4.5005
R3669 DVDD.n6603 DVDD.n6470 4.5005
R3670 DVDD.n6605 DVDD.n6470 4.5005
R3671 DVDD.n6603 DVDD.n3402 4.5005
R3672 DVDD.n6605 DVDD.n3402 4.5005
R3673 DVDD.n6603 DVDD.n6471 4.5005
R3674 DVDD.n6605 DVDD.n6471 4.5005
R3675 DVDD.n6603 DVDD.n3401 4.5005
R3676 DVDD.n6605 DVDD.n3401 4.5005
R3677 DVDD.n6603 DVDD.n6472 4.5005
R3678 DVDD.n6605 DVDD.n6472 4.5005
R3679 DVDD.n6603 DVDD.n3400 4.5005
R3680 DVDD.n6605 DVDD.n3400 4.5005
R3681 DVDD.n6603 DVDD.n6473 4.5005
R3682 DVDD.n6481 DVDD.n6473 4.5005
R3683 DVDD.n6605 DVDD.n6473 4.5005
R3684 DVDD.n6485 DVDD.n3399 4.5005
R3685 DVDD.n6603 DVDD.n3399 4.5005
R3686 DVDD.n6481 DVDD.n3399 4.5005
R3687 DVDD.n6605 DVDD.n3399 4.5005
R3688 DVDD.n6485 DVDD.n6474 4.5005
R3689 DVDD.n6603 DVDD.n6474 4.5005
R3690 DVDD.n6481 DVDD.n6474 4.5005
R3691 DVDD.n6605 DVDD.n6474 4.5005
R3692 DVDD.n6485 DVDD.n3398 4.5005
R3693 DVDD.n6603 DVDD.n3398 4.5005
R3694 DVDD.n6481 DVDD.n3398 4.5005
R3695 DVDD.n6605 DVDD.n3398 4.5005
R3696 DVDD.n6485 DVDD.n6475 4.5005
R3697 DVDD.n6603 DVDD.n6475 4.5005
R3698 DVDD.n6481 DVDD.n6475 4.5005
R3699 DVDD.n6605 DVDD.n6475 4.5005
R3700 DVDD.n6485 DVDD.n3397 4.5005
R3701 DVDD.n6603 DVDD.n3397 4.5005
R3702 DVDD.n6481 DVDD.n3397 4.5005
R3703 DVDD.n6605 DVDD.n3397 4.5005
R3704 DVDD.n6485 DVDD.n6476 4.5005
R3705 DVDD.n6603 DVDD.n6476 4.5005
R3706 DVDD.n6481 DVDD.n6476 4.5005
R3707 DVDD.n6605 DVDD.n6476 4.5005
R3708 DVDD.n6485 DVDD.n3396 4.5005
R3709 DVDD.n6603 DVDD.n3396 4.5005
R3710 DVDD.n6481 DVDD.n3396 4.5005
R3711 DVDD.n6605 DVDD.n3396 4.5005
R3712 DVDD.n6604 DVDD.n6485 4.5005
R3713 DVDD.n6604 DVDD.n6603 4.5005
R3714 DVDD.n6604 DVDD.n6481 4.5005
R3715 DVDD.n6605 DVDD.n6604 4.5005
R3716 DVDD.n3492 DVDD.n3474 4.5005
R3717 DVDD.n3474 DVDD.n3467 4.5005
R3718 DVDD.n3474 DVDD.n3420 4.5005
R3719 DVDD.n6464 DVDD.n3474 4.5005
R3720 DVDD.n3493 DVDD.n3472 4.5005
R3721 DVDD.n3472 DVDD.n3467 4.5005
R3722 DVDD.n3472 DVDD.n3420 4.5005
R3723 DVDD.n6464 DVDD.n3472 4.5005
R3724 DVDD.n3495 DVDD.n3475 4.5005
R3725 DVDD.n3475 DVDD.n3467 4.5005
R3726 DVDD.n3475 DVDD.n3420 4.5005
R3727 DVDD.n6464 DVDD.n3475 4.5005
R3728 DVDD.n3497 DVDD.n3471 4.5005
R3729 DVDD.n3471 DVDD.n3467 4.5005
R3730 DVDD.n6464 DVDD.n3471 4.5005
R3731 DVDD.n3487 DVDD.n3478 4.5005
R3732 DVDD.n6464 DVDD.n3478 4.5005
R3733 DVDD.n6449 DVDD.n3470 4.5005
R3734 DVDD.n6464 DVDD.n3470 4.5005
R3735 DVDD.n6451 DVDD.n3481 4.5005
R3736 DVDD.n6464 DVDD.n3481 4.5005
R3737 DVDD.n6452 DVDD.n3469 4.5005
R3738 DVDD.n6464 DVDD.n3469 4.5005
R3739 DVDD.n6463 DVDD.n6461 4.5005
R3740 DVDD.n6464 DVDD.n6463 4.5005
R3741 DVDD.n6460 DVDD.n3419 4.5005
R3742 DVDD.n3420 DVDD.n3419 4.5005
R3743 DVDD.n6464 DVDD.n3419 4.5005
R3744 DVDD.n6465 DVDD.n3421 4.5005
R3745 DVDD.n6465 DVDD.n3467 4.5005
R3746 DVDD.n6465 DVDD.n3420 4.5005
R3747 DVDD.n6465 DVDD.n6464 4.5005
R3748 DVDD.n3551 DVDD.n3533 4.5005
R3749 DVDD.n6397 DVDD.n3533 4.5005
R3750 DVDD.n6399 DVDD.n3533 4.5005
R3751 DVDD.n6397 DVDD.n3535 4.5005
R3752 DVDD.n6399 DVDD.n3535 4.5005
R3753 DVDD.n6397 DVDD.n3532 4.5005
R3754 DVDD.n6399 DVDD.n3532 4.5005
R3755 DVDD.n3551 DVDD.n3536 4.5005
R3756 DVDD.n6397 DVDD.n3536 4.5005
R3757 DVDD.n6399 DVDD.n3536 4.5005
R3758 DVDD.n3551 DVDD.n3531 4.5005
R3759 DVDD.n6397 DVDD.n3531 4.5005
R3760 DVDD.n3549 DVDD.n3531 4.5005
R3761 DVDD.n6399 DVDD.n3531 4.5005
R3762 DVDD.n3551 DVDD.n3537 4.5005
R3763 DVDD.n6397 DVDD.n3537 4.5005
R3764 DVDD.n3549 DVDD.n3537 4.5005
R3765 DVDD.n6399 DVDD.n3537 4.5005
R3766 DVDD.n3551 DVDD.n3530 4.5005
R3767 DVDD.n6397 DVDD.n3530 4.5005
R3768 DVDD.n3549 DVDD.n3530 4.5005
R3769 DVDD.n6399 DVDD.n3530 4.5005
R3770 DVDD.n3551 DVDD.n3538 4.5005
R3771 DVDD.n6397 DVDD.n3538 4.5005
R3772 DVDD.n3549 DVDD.n3538 4.5005
R3773 DVDD.n6399 DVDD.n3538 4.5005
R3774 DVDD.n3551 DVDD.n3529 4.5005
R3775 DVDD.n6397 DVDD.n3529 4.5005
R3776 DVDD.n3549 DVDD.n3529 4.5005
R3777 DVDD.n6399 DVDD.n3529 4.5005
R3778 DVDD.n3551 DVDD.n3539 4.5005
R3779 DVDD.n6397 DVDD.n3539 4.5005
R3780 DVDD.n3549 DVDD.n3539 4.5005
R3781 DVDD.n6399 DVDD.n3539 4.5005
R3782 DVDD.n3551 DVDD.n3528 4.5005
R3783 DVDD.n6397 DVDD.n3528 4.5005
R3784 DVDD.n3549 DVDD.n3528 4.5005
R3785 DVDD.n6399 DVDD.n3528 4.5005
R3786 DVDD.n3551 DVDD.n3540 4.5005
R3787 DVDD.n6397 DVDD.n3540 4.5005
R3788 DVDD.n3549 DVDD.n3540 4.5005
R3789 DVDD.n6399 DVDD.n3540 4.5005
R3790 DVDD.n3551 DVDD.n3527 4.5005
R3791 DVDD.n6397 DVDD.n3527 4.5005
R3792 DVDD.n3549 DVDD.n3527 4.5005
R3793 DVDD.n6399 DVDD.n3527 4.5005
R3794 DVDD.n3551 DVDD.n3541 4.5005
R3795 DVDD.n6397 DVDD.n3541 4.5005
R3796 DVDD.n3549 DVDD.n3541 4.5005
R3797 DVDD.n6399 DVDD.n3541 4.5005
R3798 DVDD.n3551 DVDD.n3526 4.5005
R3799 DVDD.n6397 DVDD.n3526 4.5005
R3800 DVDD.n3549 DVDD.n3526 4.5005
R3801 DVDD.n6399 DVDD.n3526 4.5005
R3802 DVDD.n3551 DVDD.n3542 4.5005
R3803 DVDD.n6397 DVDD.n3542 4.5005
R3804 DVDD.n3549 DVDD.n3542 4.5005
R3805 DVDD.n6399 DVDD.n3542 4.5005
R3806 DVDD.n3551 DVDD.n3525 4.5005
R3807 DVDD.n6397 DVDD.n3525 4.5005
R3808 DVDD.n3549 DVDD.n3525 4.5005
R3809 DVDD.n6399 DVDD.n3525 4.5005
R3810 DVDD.n3551 DVDD.n3543 4.5005
R3811 DVDD.n6397 DVDD.n3543 4.5005
R3812 DVDD.n3549 DVDD.n3543 4.5005
R3813 DVDD.n6399 DVDD.n3543 4.5005
R3814 DVDD.n3551 DVDD.n3524 4.5005
R3815 DVDD.n6397 DVDD.n3524 4.5005
R3816 DVDD.n3549 DVDD.n3524 4.5005
R3817 DVDD.n6399 DVDD.n3524 4.5005
R3818 DVDD.n3551 DVDD.n3544 4.5005
R3819 DVDD.n6397 DVDD.n3544 4.5005
R3820 DVDD.n3549 DVDD.n3544 4.5005
R3821 DVDD.n6399 DVDD.n3544 4.5005
R3822 DVDD.n3551 DVDD.n3523 4.5005
R3823 DVDD.n6397 DVDD.n3523 4.5005
R3824 DVDD.n3549 DVDD.n3523 4.5005
R3825 DVDD.n6399 DVDD.n3523 4.5005
R3826 DVDD.n3551 DVDD.n3545 4.5005
R3827 DVDD.n6397 DVDD.n3545 4.5005
R3828 DVDD.n3549 DVDD.n3545 4.5005
R3829 DVDD.n6399 DVDD.n3545 4.5005
R3830 DVDD.n3551 DVDD.n3522 4.5005
R3831 DVDD.n6397 DVDD.n3522 4.5005
R3832 DVDD.n3549 DVDD.n3522 4.5005
R3833 DVDD.n6399 DVDD.n3522 4.5005
R3834 DVDD.n6398 DVDD.n3551 4.5005
R3835 DVDD.n6398 DVDD.n6397 4.5005
R3836 DVDD.n6398 DVDD.n3549 4.5005
R3837 DVDD.n6399 DVDD.n6398 4.5005
R3838 DVDD.n8667 DVDD.n1056 4.5005
R3839 DVDD.n8667 DVDD.n1057 4.5005
R3840 DVDD.n8667 DVDD.n8666 4.5005
R3841 DVDD.n1072 DVDD.n1057 4.5005
R3842 DVDD.n8666 DVDD.n1072 4.5005
R3843 DVDD.n1069 DVDD.n1057 4.5005
R3844 DVDD.n8666 DVDD.n1069 4.5005
R3845 DVDD.n1074 DVDD.n1057 4.5005
R3846 DVDD.n8666 DVDD.n1074 4.5005
R3847 DVDD.n1068 DVDD.n1057 4.5005
R3848 DVDD.n8666 DVDD.n1068 4.5005
R3849 DVDD.n1076 DVDD.n1057 4.5005
R3850 DVDD.n8666 DVDD.n1076 4.5005
R3851 DVDD.n1067 DVDD.n1057 4.5005
R3852 DVDD.n8666 DVDD.n1067 4.5005
R3853 DVDD.n1078 DVDD.n1057 4.5005
R3854 DVDD.n8666 DVDD.n1078 4.5005
R3855 DVDD.n1066 DVDD.n1057 4.5005
R3856 DVDD.n8666 DVDD.n1066 4.5005
R3857 DVDD.n1080 DVDD.n1057 4.5005
R3858 DVDD.n8666 DVDD.n1080 4.5005
R3859 DVDD.n1065 DVDD.n1057 4.5005
R3860 DVDD.n8666 DVDD.n1065 4.5005
R3861 DVDD.n1082 DVDD.n1057 4.5005
R3862 DVDD.n8666 DVDD.n1082 4.5005
R3863 DVDD.n1064 DVDD.n1057 4.5005
R3864 DVDD.n8666 DVDD.n1064 4.5005
R3865 DVDD.n1084 DVDD.n1057 4.5005
R3866 DVDD.n8666 DVDD.n1084 4.5005
R3867 DVDD.n1063 DVDD.n1057 4.5005
R3868 DVDD.n8666 DVDD.n1063 4.5005
R3869 DVDD.n1086 DVDD.n1057 4.5005
R3870 DVDD.n8666 DVDD.n1086 4.5005
R3871 DVDD.n1062 DVDD.n1057 4.5005
R3872 DVDD.n8666 DVDD.n1062 4.5005
R3873 DVDD.n1088 DVDD.n1057 4.5005
R3874 DVDD.n8666 DVDD.n1088 4.5005
R3875 DVDD.n1061 DVDD.n1057 4.5005
R3876 DVDD.n8666 DVDD.n1061 4.5005
R3877 DVDD.n1090 DVDD.n1057 4.5005
R3878 DVDD.n8666 DVDD.n1090 4.5005
R3879 DVDD.n1060 DVDD.n1057 4.5005
R3880 DVDD.n8666 DVDD.n1060 4.5005
R3881 DVDD.n1092 DVDD.n1057 4.5005
R3882 DVDD.n8666 DVDD.n1092 4.5005
R3883 DVDD.n1059 DVDD.n1057 4.5005
R3884 DVDD.n8666 DVDD.n1059 4.5005
R3885 DVDD.n8665 DVDD.n1056 4.5005
R3886 DVDD.n8665 DVDD.n1057 4.5005
R3887 DVDD.n8666 DVDD.n8665 4.5005
R3888 DVDD.n8664 DVDD.n1095 4.5005
R3889 DVDD.n8664 DVDD.n1096 4.5005
R3890 DVDD.n8664 DVDD.n8663 4.5005
R3891 DVDD.n1101 DVDD.n1096 4.5005
R3892 DVDD.n8663 DVDD.n1101 4.5005
R3893 DVDD.n1104 DVDD.n1096 4.5005
R3894 DVDD.n8663 DVDD.n1104 4.5005
R3895 DVDD.n1100 DVDD.n1096 4.5005
R3896 DVDD.n8663 DVDD.n1100 4.5005
R3897 DVDD.n1106 DVDD.n1096 4.5005
R3898 DVDD.n8663 DVDD.n1106 4.5005
R3899 DVDD.n1099 DVDD.n1096 4.5005
R3900 DVDD.n8663 DVDD.n1099 4.5005
R3901 DVDD.n1108 DVDD.n1096 4.5005
R3902 DVDD.n8663 DVDD.n1108 4.5005
R3903 DVDD.n1098 DVDD.n1096 4.5005
R3904 DVDD.n8663 DVDD.n1098 4.5005
R3905 DVDD.n1110 DVDD.n1096 4.5005
R3906 DVDD.n8663 DVDD.n1110 4.5005
R3907 DVDD.n1097 DVDD.n1096 4.5005
R3908 DVDD.n8663 DVDD.n1097 4.5005
R3909 DVDD.n8662 DVDD.n1096 4.5005
R3910 DVDD.n8662 DVDD.n1116 4.5005
R3911 DVDD.n8663 DVDD.n8662 4.5005
R3912 DVDD.n8661 DVDD.n1118 4.5005
R3913 DVDD.n8661 DVDD.n1119 4.5005
R3914 DVDD.n8661 DVDD.n8660 4.5005
R3915 DVDD.n1134 DVDD.n1119 4.5005
R3916 DVDD.n8660 DVDD.n1134 4.5005
R3917 DVDD.n1131 DVDD.n1119 4.5005
R3918 DVDD.n8660 DVDD.n1131 4.5005
R3919 DVDD.n1136 DVDD.n1119 4.5005
R3920 DVDD.n8660 DVDD.n1136 4.5005
R3921 DVDD.n1130 DVDD.n1119 4.5005
R3922 DVDD.n8660 DVDD.n1130 4.5005
R3923 DVDD.n1138 DVDD.n1119 4.5005
R3924 DVDD.n8660 DVDD.n1138 4.5005
R3925 DVDD.n1129 DVDD.n1119 4.5005
R3926 DVDD.n8660 DVDD.n1129 4.5005
R3927 DVDD.n1140 DVDD.n1119 4.5005
R3928 DVDD.n8660 DVDD.n1140 4.5005
R3929 DVDD.n1128 DVDD.n1119 4.5005
R3930 DVDD.n8660 DVDD.n1128 4.5005
R3931 DVDD.n1142 DVDD.n1119 4.5005
R3932 DVDD.n8660 DVDD.n1142 4.5005
R3933 DVDD.n1127 DVDD.n1119 4.5005
R3934 DVDD.n8660 DVDD.n1127 4.5005
R3935 DVDD.n1144 DVDD.n1119 4.5005
R3936 DVDD.n8660 DVDD.n1144 4.5005
R3937 DVDD.n1126 DVDD.n1119 4.5005
R3938 DVDD.n8660 DVDD.n1126 4.5005
R3939 DVDD.n1146 DVDD.n1119 4.5005
R3940 DVDD.n8660 DVDD.n1146 4.5005
R3941 DVDD.n1125 DVDD.n1119 4.5005
R3942 DVDD.n8660 DVDD.n1125 4.5005
R3943 DVDD.n1148 DVDD.n1119 4.5005
R3944 DVDD.n8660 DVDD.n1148 4.5005
R3945 DVDD.n1124 DVDD.n1119 4.5005
R3946 DVDD.n8660 DVDD.n1124 4.5005
R3947 DVDD.n1150 DVDD.n1119 4.5005
R3948 DVDD.n8660 DVDD.n1150 4.5005
R3949 DVDD.n1123 DVDD.n1119 4.5005
R3950 DVDD.n8660 DVDD.n1123 4.5005
R3951 DVDD.n1152 DVDD.n1119 4.5005
R3952 DVDD.n8660 DVDD.n1152 4.5005
R3953 DVDD.n1122 DVDD.n1119 4.5005
R3954 DVDD.n8660 DVDD.n1122 4.5005
R3955 DVDD.n1154 DVDD.n1119 4.5005
R3956 DVDD.n8660 DVDD.n1154 4.5005
R3957 DVDD.n1121 DVDD.n1119 4.5005
R3958 DVDD.n8660 DVDD.n1121 4.5005
R3959 DVDD.n8659 DVDD.n1118 4.5005
R3960 DVDD.n8659 DVDD.n1119 4.5005
R3961 DVDD.n8660 DVDD.n8659 4.5005
R3962 DVDD.n8658 DVDD.n1157 4.5005
R3963 DVDD.n8658 DVDD.n1158 4.5005
R3964 DVDD.n8658 DVDD.n8657 4.5005
R3965 DVDD.n1173 DVDD.n1158 4.5005
R3966 DVDD.n8657 DVDD.n1173 4.5005
R3967 DVDD.n1170 DVDD.n1158 4.5005
R3968 DVDD.n8657 DVDD.n1170 4.5005
R3969 DVDD.n1175 DVDD.n1158 4.5005
R3970 DVDD.n8657 DVDD.n1175 4.5005
R3971 DVDD.n1169 DVDD.n1158 4.5005
R3972 DVDD.n8657 DVDD.n1169 4.5005
R3973 DVDD.n1177 DVDD.n1158 4.5005
R3974 DVDD.n8657 DVDD.n1177 4.5005
R3975 DVDD.n1168 DVDD.n1158 4.5005
R3976 DVDD.n8657 DVDD.n1168 4.5005
R3977 DVDD.n1179 DVDD.n1158 4.5005
R3978 DVDD.n8657 DVDD.n1179 4.5005
R3979 DVDD.n1167 DVDD.n1158 4.5005
R3980 DVDD.n8657 DVDD.n1167 4.5005
R3981 DVDD.n1181 DVDD.n1158 4.5005
R3982 DVDD.n8657 DVDD.n1181 4.5005
R3983 DVDD.n1166 DVDD.n1158 4.5005
R3984 DVDD.n8657 DVDD.n1166 4.5005
R3985 DVDD.n1183 DVDD.n1158 4.5005
R3986 DVDD.n8657 DVDD.n1183 4.5005
R3987 DVDD.n1165 DVDD.n1158 4.5005
R3988 DVDD.n8657 DVDD.n1165 4.5005
R3989 DVDD.n1185 DVDD.n1158 4.5005
R3990 DVDD.n8657 DVDD.n1185 4.5005
R3991 DVDD.n1164 DVDD.n1158 4.5005
R3992 DVDD.n8657 DVDD.n1164 4.5005
R3993 DVDD.n1187 DVDD.n1158 4.5005
R3994 DVDD.n8657 DVDD.n1187 4.5005
R3995 DVDD.n1163 DVDD.n1158 4.5005
R3996 DVDD.n8657 DVDD.n1163 4.5005
R3997 DVDD.n1189 DVDD.n1158 4.5005
R3998 DVDD.n8657 DVDD.n1189 4.5005
R3999 DVDD.n1162 DVDD.n1158 4.5005
R4000 DVDD.n8657 DVDD.n1162 4.5005
R4001 DVDD.n1191 DVDD.n1158 4.5005
R4002 DVDD.n8657 DVDD.n1191 4.5005
R4003 DVDD.n1161 DVDD.n1158 4.5005
R4004 DVDD.n8657 DVDD.n1161 4.5005
R4005 DVDD.n1193 DVDD.n1158 4.5005
R4006 DVDD.n8657 DVDD.n1193 4.5005
R4007 DVDD.n1160 DVDD.n1158 4.5005
R4008 DVDD.n8657 DVDD.n1160 4.5005
R4009 DVDD.n8656 DVDD.n1157 4.5005
R4010 DVDD.n8656 DVDD.n1158 4.5005
R4011 DVDD.n8657 DVDD.n8656 4.5005
R4012 DVDD.n8655 DVDD.n1196 4.5005
R4013 DVDD.n8655 DVDD.n1197 4.5005
R4014 DVDD.n8655 DVDD.n8654 4.5005
R4015 DVDD.n1212 DVDD.n1197 4.5005
R4016 DVDD.n8654 DVDD.n1212 4.5005
R4017 DVDD.n1209 DVDD.n1197 4.5005
R4018 DVDD.n8654 DVDD.n1209 4.5005
R4019 DVDD.n1214 DVDD.n1197 4.5005
R4020 DVDD.n8654 DVDD.n1214 4.5005
R4021 DVDD.n1208 DVDD.n1197 4.5005
R4022 DVDD.n8654 DVDD.n1208 4.5005
R4023 DVDD.n1216 DVDD.n1197 4.5005
R4024 DVDD.n8654 DVDD.n1216 4.5005
R4025 DVDD.n1207 DVDD.n1197 4.5005
R4026 DVDD.n8654 DVDD.n1207 4.5005
R4027 DVDD.n1218 DVDD.n1197 4.5005
R4028 DVDD.n8654 DVDD.n1218 4.5005
R4029 DVDD.n1206 DVDD.n1197 4.5005
R4030 DVDD.n8654 DVDD.n1206 4.5005
R4031 DVDD.n1220 DVDD.n1197 4.5005
R4032 DVDD.n8654 DVDD.n1220 4.5005
R4033 DVDD.n1205 DVDD.n1197 4.5005
R4034 DVDD.n8654 DVDD.n1205 4.5005
R4035 DVDD.n1222 DVDD.n1197 4.5005
R4036 DVDD.n8654 DVDD.n1222 4.5005
R4037 DVDD.n1204 DVDD.n1197 4.5005
R4038 DVDD.n8654 DVDD.n1204 4.5005
R4039 DVDD.n1224 DVDD.n1197 4.5005
R4040 DVDD.n8654 DVDD.n1224 4.5005
R4041 DVDD.n1203 DVDD.n1197 4.5005
R4042 DVDD.n8654 DVDD.n1203 4.5005
R4043 DVDD.n1226 DVDD.n1197 4.5005
R4044 DVDD.n8654 DVDD.n1226 4.5005
R4045 DVDD.n1202 DVDD.n1197 4.5005
R4046 DVDD.n8654 DVDD.n1202 4.5005
R4047 DVDD.n1228 DVDD.n1197 4.5005
R4048 DVDD.n8654 DVDD.n1228 4.5005
R4049 DVDD.n1201 DVDD.n1197 4.5005
R4050 DVDD.n8654 DVDD.n1201 4.5005
R4051 DVDD.n1230 DVDD.n1197 4.5005
R4052 DVDD.n8654 DVDD.n1230 4.5005
R4053 DVDD.n1200 DVDD.n1197 4.5005
R4054 DVDD.n8654 DVDD.n1200 4.5005
R4055 DVDD.n1232 DVDD.n1197 4.5005
R4056 DVDD.n8654 DVDD.n1232 4.5005
R4057 DVDD.n1199 DVDD.n1197 4.5005
R4058 DVDD.n8654 DVDD.n1199 4.5005
R4059 DVDD.n8653 DVDD.n1196 4.5005
R4060 DVDD.n8653 DVDD.n1197 4.5005
R4061 DVDD.n8654 DVDD.n8653 4.5005
R4062 DVDD.n8652 DVDD.n1235 4.5005
R4063 DVDD.n8652 DVDD.n1236 4.5005
R4064 DVDD.n8652 DVDD.n8651 4.5005
R4065 DVDD.n1251 DVDD.n1236 4.5005
R4066 DVDD.n8651 DVDD.n1251 4.5005
R4067 DVDD.n1248 DVDD.n1236 4.5005
R4068 DVDD.n8651 DVDD.n1248 4.5005
R4069 DVDD.n1253 DVDD.n1236 4.5005
R4070 DVDD.n8651 DVDD.n1253 4.5005
R4071 DVDD.n1247 DVDD.n1236 4.5005
R4072 DVDD.n8651 DVDD.n1247 4.5005
R4073 DVDD.n1255 DVDD.n1236 4.5005
R4074 DVDD.n8651 DVDD.n1255 4.5005
R4075 DVDD.n1246 DVDD.n1236 4.5005
R4076 DVDD.n8651 DVDD.n1246 4.5005
R4077 DVDD.n1257 DVDD.n1236 4.5005
R4078 DVDD.n8651 DVDD.n1257 4.5005
R4079 DVDD.n1245 DVDD.n1236 4.5005
R4080 DVDD.n8651 DVDD.n1245 4.5005
R4081 DVDD.n1259 DVDD.n1236 4.5005
R4082 DVDD.n8651 DVDD.n1259 4.5005
R4083 DVDD.n1244 DVDD.n1236 4.5005
R4084 DVDD.n8651 DVDD.n1244 4.5005
R4085 DVDD.n1261 DVDD.n1236 4.5005
R4086 DVDD.n8651 DVDD.n1261 4.5005
R4087 DVDD.n1243 DVDD.n1236 4.5005
R4088 DVDD.n8651 DVDD.n1243 4.5005
R4089 DVDD.n1263 DVDD.n1236 4.5005
R4090 DVDD.n8651 DVDD.n1263 4.5005
R4091 DVDD.n1242 DVDD.n1236 4.5005
R4092 DVDD.n8151 DVDD.n1242 4.5005
R4093 DVDD.n8651 DVDD.n1242 4.5005
R4094 DVDD.n1264 DVDD.n1235 4.5005
R4095 DVDD.n1264 DVDD.n1236 4.5005
R4096 DVDD.n8151 DVDD.n1264 4.5005
R4097 DVDD.n8651 DVDD.n1264 4.5005
R4098 DVDD.n1241 DVDD.n1235 4.5005
R4099 DVDD.n1241 DVDD.n1236 4.5005
R4100 DVDD.n8151 DVDD.n1241 4.5005
R4101 DVDD.n8651 DVDD.n1241 4.5005
R4102 DVDD.n1265 DVDD.n1235 4.5005
R4103 DVDD.n1265 DVDD.n1236 4.5005
R4104 DVDD.n8151 DVDD.n1265 4.5005
R4105 DVDD.n8651 DVDD.n1265 4.5005
R4106 DVDD.n1240 DVDD.n1235 4.5005
R4107 DVDD.n1240 DVDD.n1236 4.5005
R4108 DVDD.n8651 DVDD.n1240 4.5005
R4109 DVDD.n1267 DVDD.n1236 4.5005
R4110 DVDD.n8651 DVDD.n1267 4.5005
R4111 DVDD.n1239 DVDD.n1236 4.5005
R4112 DVDD.n8651 DVDD.n1239 4.5005
R4113 DVDD.n1269 DVDD.n1236 4.5005
R4114 DVDD.n8651 DVDD.n1269 4.5005
R4115 DVDD.n1238 DVDD.n1236 4.5005
R4116 DVDD.n8651 DVDD.n1238 4.5005
R4117 DVDD.n8650 DVDD.n1235 4.5005
R4118 DVDD.n8650 DVDD.n1236 4.5005
R4119 DVDD.n8651 DVDD.n8650 4.5005
R4120 DVDD.n8649 DVDD.n1272 4.5005
R4121 DVDD.n8649 DVDD.n1273 4.5005
R4122 DVDD.n8649 DVDD.n8648 4.5005
R4123 DVDD.n1279 DVDD.n1273 4.5005
R4124 DVDD.n8648 DVDD.n1279 4.5005
R4125 DVDD.n1282 DVDD.n1273 4.5005
R4126 DVDD.n8648 DVDD.n1282 4.5005
R4127 DVDD.n1278 DVDD.n1273 4.5005
R4128 DVDD.n8648 DVDD.n1278 4.5005
R4129 DVDD.n1284 DVDD.n1273 4.5005
R4130 DVDD.n8648 DVDD.n1284 4.5005
R4131 DVDD.n1277 DVDD.n1273 4.5005
R4132 DVDD.n8648 DVDD.n1277 4.5005
R4133 DVDD.n1286 DVDD.n1273 4.5005
R4134 DVDD.n8648 DVDD.n1286 4.5005
R4135 DVDD.n1276 DVDD.n1273 4.5005
R4136 DVDD.n8648 DVDD.n1276 4.5005
R4137 DVDD.n1288 DVDD.n1273 4.5005
R4138 DVDD.n8648 DVDD.n1288 4.5005
R4139 DVDD.n1275 DVDD.n1273 4.5005
R4140 DVDD.n8648 DVDD.n1275 4.5005
R4141 DVDD.n8647 DVDD.n1273 4.5005
R4142 DVDD.n8647 DVDD.n1294 4.5005
R4143 DVDD.n8648 DVDD.n8647 4.5005
R4144 DVDD.n8644 DVDD.n1299 4.5005
R4145 DVDD.n8644 DVDD.n1295 4.5005
R4146 DVDD.n8646 DVDD.n1296 4.5005
R4147 DVDD.n8646 DVDD.n1299 4.5005
R4148 DVDD.n8646 DVDD.n1295 4.5005
R4149 DVDD.n7172 DVDD.n7164 4.5005
R4150 DVDD.n7172 DVDD.n7165 4.5005
R4151 DVDD.n7170 DVDD.n7165 4.5005
R4152 DVDD.n7168 DVDD.n7165 4.5005
R4153 DVDD.n7172 DVDD.n7171 4.5005
R4154 DVDD.n7171 DVDD.n7170 4.5005
R4155 DVDD.n7171 DVDD.n7168 4.5005
R4156 DVDD.n8645 DVDD.n1302 4.5005
R4157 DVDD.n8645 DVDD.n8644 4.5005
R4158 DVDD.n8646 DVDD.n8645 4.5005
R4159 DVDD.n7164 DVDD.n1303 4.5005
R4160 DVDD.n7165 DVDD.n1303 4.5005
R4161 DVDD.n7171 DVDD.n1303 4.5005
R4162 DVDD.n8450 DVDD.n8449 4.5005
R4163 DVDD.n8451 DVDD.n8450 4.5005
R4164 DVDD.n8467 DVDD.n8466 4.5005
R4165 DVDD.n8467 DVDD.n1444 4.5005
R4166 DVDD.n8491 DVDD.n8490 4.5005
R4167 DVDD.n8490 DVDD.n8489 4.5005
R4168 DVDD.n8606 DVDD.n8605 4.5005
R4169 DVDD.n8605 DVDD.n8604 4.5005
R4170 DVDD.n8910 DVDD.n619 4.5005
R4171 DVDD.n8912 DVDD.n619 4.5005
R4172 DVDD.n619 DVDD.n611 4.5005
R4173 DVDD.n8910 DVDD.n616 4.5005
R4174 DVDD.n8912 DVDD.n616 4.5005
R4175 DVDD.n8912 DVDD.n621 4.5005
R4176 DVDD.n621 DVDD.n606 4.5005
R4177 DVDD.n8912 DVDD.n615 4.5005
R4178 DVDD.n615 DVDD.n606 4.5005
R4179 DVDD.n8912 DVDD.n623 4.5005
R4180 DVDD.n623 DVDD.n606 4.5005
R4181 DVDD.n8912 DVDD.n614 4.5005
R4182 DVDD.n614 DVDD.n606 4.5005
R4183 DVDD.n8912 DVDD.n625 4.5005
R4184 DVDD.n625 DVDD.n606 4.5005
R4185 DVDD.n8912 DVDD.n613 4.5005
R4186 DVDD.n613 DVDD.n606 4.5005
R4187 DVDD.n8912 DVDD.n627 4.5005
R4188 DVDD.n627 DVDD.n606 4.5005
R4189 DVDD.n8912 DVDD.n612 4.5005
R4190 DVDD.n612 DVDD.n606 4.5005
R4191 DVDD.n8911 DVDD.n8910 4.5005
R4192 DVDD.n8912 DVDD.n8911 4.5005
R4193 DVDD.n8911 DVDD.n606 4.5005
R4194 DVDD.n649 DVDD.n637 4.5005
R4195 DVDD.n649 DVDD.n642 4.5005
R4196 DVDD.n8894 DVDD.n649 4.5005
R4197 DVDD.n8892 DVDD.n649 4.5005
R4198 DVDD.n647 DVDD.n637 4.5005
R4199 DVDD.n647 DVDD.n642 4.5005
R4200 DVDD.n8894 DVDD.n647 4.5005
R4201 DVDD.n8892 DVDD.n647 4.5005
R4202 DVDD.n650 DVDD.n637 4.5005
R4203 DVDD.n650 DVDD.n642 4.5005
R4204 DVDD.n8894 DVDD.n650 4.5005
R4205 DVDD.n8892 DVDD.n650 4.5005
R4206 DVDD.n646 DVDD.n637 4.5005
R4207 DVDD.n646 DVDD.n642 4.5005
R4208 DVDD.n8894 DVDD.n646 4.5005
R4209 DVDD.n8892 DVDD.n646 4.5005
R4210 DVDD.n651 DVDD.n637 4.5005
R4211 DVDD.n651 DVDD.n642 4.5005
R4212 DVDD.n8894 DVDD.n651 4.5005
R4213 DVDD.n8892 DVDD.n651 4.5005
R4214 DVDD.n645 DVDD.n637 4.5005
R4215 DVDD.n645 DVDD.n642 4.5005
R4216 DVDD.n8894 DVDD.n645 4.5005
R4217 DVDD.n8892 DVDD.n645 4.5005
R4218 DVDD.n652 DVDD.n637 4.5005
R4219 DVDD.n652 DVDD.n642 4.5005
R4220 DVDD.n8894 DVDD.n652 4.5005
R4221 DVDD.n8892 DVDD.n652 4.5005
R4222 DVDD.n644 DVDD.n637 4.5005
R4223 DVDD.n644 DVDD.n642 4.5005
R4224 DVDD.n8894 DVDD.n644 4.5005
R4225 DVDD.n8892 DVDD.n644 4.5005
R4226 DVDD.n653 DVDD.n637 4.5005
R4227 DVDD.n653 DVDD.n642 4.5005
R4228 DVDD.n8894 DVDD.n653 4.5005
R4229 DVDD.n8892 DVDD.n653 4.5005
R4230 DVDD.n643 DVDD.n637 4.5005
R4231 DVDD.n643 DVDD.n642 4.5005
R4232 DVDD.n8894 DVDD.n643 4.5005
R4233 DVDD.n8892 DVDD.n643 4.5005
R4234 DVDD.n8893 DVDD.n637 4.5005
R4235 DVDD.n8893 DVDD.n642 4.5005
R4236 DVDD.n8894 DVDD.n8893 4.5005
R4237 DVDD.n8893 DVDD.n8892 4.5005
R4238 DVDD.n5157 DVDD.n5116 4.5005
R4239 DVDD.n5116 DVDD.n4571 4.5005
R4240 DVDD.n5116 DVDD.n4573 4.5005
R4241 DVDD.n5116 DVDD.n4570 4.5005
R4242 DVDD.n5157 DVDD.n4579 4.5005
R4243 DVDD.n4579 DVDD.n4571 4.5005
R4244 DVDD.n4579 DVDD.n4573 4.5005
R4245 DVDD.n4579 DVDD.n4570 4.5005
R4246 DVDD.n5157 DVDD.n5117 4.5005
R4247 DVDD.n5117 DVDD.n4571 4.5005
R4248 DVDD.n5117 DVDD.n4573 4.5005
R4249 DVDD.n5117 DVDD.n4570 4.5005
R4250 DVDD.n5156 DVDD.n4571 4.5005
R4251 DVDD.n5156 DVDD.n4573 4.5005
R4252 DVDD.n5156 DVDD.n4570 4.5005
R4253 DVDD.n4575 DVDD.n4571 4.5005
R4254 DVDD.n4575 DVDD.n4573 4.5005
R4255 DVDD.n4575 DVDD.n4570 4.5005
R4256 DVDD.n5119 DVDD.n4571 4.5005
R4257 DVDD.n5119 DVDD.n4573 4.5005
R4258 DVDD.n5119 DVDD.n4570 4.5005
R4259 DVDD.n5157 DVDD.n4578 4.5005
R4260 DVDD.n4578 DVDD.n4571 4.5005
R4261 DVDD.n4578 DVDD.n4573 4.5005
R4262 DVDD.n4578 DVDD.n4570 4.5005
R4263 DVDD.n5157 DVDD.n5118 4.5005
R4264 DVDD.n5118 DVDD.n4571 4.5005
R4265 DVDD.n5118 DVDD.n4573 4.5005
R4266 DVDD.n5118 DVDD.n4570 4.5005
R4267 DVDD.n5157 DVDD.n4577 4.5005
R4268 DVDD.n4577 DVDD.n4571 4.5005
R4269 DVDD.n4577 DVDD.n4573 4.5005
R4270 DVDD.n4577 DVDD.n4570 4.5005
R4271 DVDD.n4576 DVDD.n4571 4.5005
R4272 DVDD.n4576 DVDD.n4573 4.5005
R4273 DVDD.n4576 DVDD.n4570 4.5005
R4274 DVDD.n5158 DVDD.n4571 4.5005
R4275 DVDD.n5158 DVDD.n4573 4.5005
R4276 DVDD.n5158 DVDD.n4570 4.5005
R4277 DVDD.n5158 DVDD.n5157 4.5005
R4278 DVDD.n5157 DVDD.n4576 4.5005
R4279 DVDD.n5157 DVDD.n5119 4.5005
R4280 DVDD.n5157 DVDD.n4575 4.5005
R4281 DVDD.n5157 DVDD.n5156 4.5005
R4282 DVDD.n9013 DVDD.n8972 4.5005
R4283 DVDD.n8972 DVDD.n549 4.5005
R4284 DVDD.n8972 DVDD.n551 4.5005
R4285 DVDD.n8972 DVDD.n548 4.5005
R4286 DVDD.n9013 DVDD.n557 4.5005
R4287 DVDD.n557 DVDD.n549 4.5005
R4288 DVDD.n557 DVDD.n551 4.5005
R4289 DVDD.n557 DVDD.n548 4.5005
R4290 DVDD.n9013 DVDD.n8973 4.5005
R4291 DVDD.n8973 DVDD.n549 4.5005
R4292 DVDD.n8973 DVDD.n551 4.5005
R4293 DVDD.n8973 DVDD.n548 4.5005
R4294 DVDD.n9012 DVDD.n549 4.5005
R4295 DVDD.n9012 DVDD.n551 4.5005
R4296 DVDD.n9012 DVDD.n548 4.5005
R4297 DVDD.n553 DVDD.n549 4.5005
R4298 DVDD.n553 DVDD.n551 4.5005
R4299 DVDD.n553 DVDD.n548 4.5005
R4300 DVDD.n8975 DVDD.n549 4.5005
R4301 DVDD.n8975 DVDD.n551 4.5005
R4302 DVDD.n8975 DVDD.n548 4.5005
R4303 DVDD.n9013 DVDD.n556 4.5005
R4304 DVDD.n556 DVDD.n549 4.5005
R4305 DVDD.n556 DVDD.n551 4.5005
R4306 DVDD.n556 DVDD.n548 4.5005
R4307 DVDD.n9013 DVDD.n8974 4.5005
R4308 DVDD.n8974 DVDD.n549 4.5005
R4309 DVDD.n8974 DVDD.n551 4.5005
R4310 DVDD.n8974 DVDD.n548 4.5005
R4311 DVDD.n9013 DVDD.n555 4.5005
R4312 DVDD.n555 DVDD.n549 4.5005
R4313 DVDD.n555 DVDD.n551 4.5005
R4314 DVDD.n555 DVDD.n548 4.5005
R4315 DVDD.n554 DVDD.n549 4.5005
R4316 DVDD.n554 DVDD.n551 4.5005
R4317 DVDD.n554 DVDD.n548 4.5005
R4318 DVDD.n9014 DVDD.n549 4.5005
R4319 DVDD.n9014 DVDD.n551 4.5005
R4320 DVDD.n9014 DVDD.n548 4.5005
R4321 DVDD.n9014 DVDD.n9013 4.5005
R4322 DVDD.n9013 DVDD.n554 4.5005
R4323 DVDD.n9013 DVDD.n8975 4.5005
R4324 DVDD.n9013 DVDD.n553 4.5005
R4325 DVDD.n9013 DVDD.n9012 4.5005
R4326 DVDD.n4625 DVDD.n4619 4.5005
R4327 DVDD.n4711 DVDD.n4619 4.5005
R4328 DVDD.n4619 DVDD.n4613 4.5005
R4329 DVDD.n4713 DVDD.n4619 4.5005
R4330 DVDD.n4625 DVDD.n4618 4.5005
R4331 DVDD.n4711 DVDD.n4618 4.5005
R4332 DVDD.n4618 DVDD.n4613 4.5005
R4333 DVDD.n4713 DVDD.n4618 4.5005
R4334 DVDD.n4625 DVDD.n4620 4.5005
R4335 DVDD.n4711 DVDD.n4620 4.5005
R4336 DVDD.n4620 DVDD.n4613 4.5005
R4337 DVDD.n4713 DVDD.n4620 4.5005
R4338 DVDD.n4625 DVDD.n4617 4.5005
R4339 DVDD.n4711 DVDD.n4617 4.5005
R4340 DVDD.n4617 DVDD.n4613 4.5005
R4341 DVDD.n4713 DVDD.n4617 4.5005
R4342 DVDD.n4625 DVDD.n4621 4.5005
R4343 DVDD.n4711 DVDD.n4621 4.5005
R4344 DVDD.n4621 DVDD.n4613 4.5005
R4345 DVDD.n4713 DVDD.n4621 4.5005
R4346 DVDD.n4625 DVDD.n4616 4.5005
R4347 DVDD.n4711 DVDD.n4616 4.5005
R4348 DVDD.n4616 DVDD.n4613 4.5005
R4349 DVDD.n4713 DVDD.n4616 4.5005
R4350 DVDD.n4625 DVDD.n4622 4.5005
R4351 DVDD.n4711 DVDD.n4622 4.5005
R4352 DVDD.n4622 DVDD.n4613 4.5005
R4353 DVDD.n4713 DVDD.n4622 4.5005
R4354 DVDD.n4625 DVDD.n4615 4.5005
R4355 DVDD.n4711 DVDD.n4615 4.5005
R4356 DVDD.n4615 DVDD.n4613 4.5005
R4357 DVDD.n4713 DVDD.n4615 4.5005
R4358 DVDD.n4625 DVDD.n4623 4.5005
R4359 DVDD.n4711 DVDD.n4623 4.5005
R4360 DVDD.n4623 DVDD.n4613 4.5005
R4361 DVDD.n4713 DVDD.n4623 4.5005
R4362 DVDD.n4625 DVDD.n4614 4.5005
R4363 DVDD.n4711 DVDD.n4614 4.5005
R4364 DVDD.n4614 DVDD.n4613 4.5005
R4365 DVDD.n4713 DVDD.n4614 4.5005
R4366 DVDD.n4713 DVDD.n4712 4.5005
R4367 DVDD.n4712 DVDD.n4613 4.5005
R4368 DVDD.n4712 DVDD.n4625 4.5005
R4369 DVDD.n4712 DVDD.n4711 4.5005
R4370 DVDD.n4869 DVDD.n4863 4.5005
R4371 DVDD.n5028 DVDD.n4863 4.5005
R4372 DVDD.n5082 DVDD.n4863 4.5005
R4373 DVDD.n5080 DVDD.n4863 4.5005
R4374 DVDD.n4869 DVDD.n4861 4.5005
R4375 DVDD.n5028 DVDD.n4861 4.5005
R4376 DVDD.n5082 DVDD.n4861 4.5005
R4377 DVDD.n5080 DVDD.n4861 4.5005
R4378 DVDD.n5080 DVDD.n4864 4.5005
R4379 DVDD.n4869 DVDD.n4864 4.5005
R4380 DVDD.n5028 DVDD.n4864 4.5005
R4381 DVDD.n5082 DVDD.n4864 4.5005
R4382 DVDD.n5080 DVDD.n4860 4.5005
R4383 DVDD.n4869 DVDD.n4860 4.5005
R4384 DVDD.n5028 DVDD.n4860 4.5005
R4385 DVDD.n5082 DVDD.n4860 4.5005
R4386 DVDD.n5080 DVDD.n4865 4.5005
R4387 DVDD.n4869 DVDD.n4865 4.5005
R4388 DVDD.n5028 DVDD.n4865 4.5005
R4389 DVDD.n5082 DVDD.n4865 4.5005
R4390 DVDD.n5080 DVDD.n4859 4.5005
R4391 DVDD.n4869 DVDD.n4859 4.5005
R4392 DVDD.n5028 DVDD.n4859 4.5005
R4393 DVDD.n5082 DVDD.n4859 4.5005
R4394 DVDD.n4869 DVDD.n4866 4.5005
R4395 DVDD.n5028 DVDD.n4866 4.5005
R4396 DVDD.n5082 DVDD.n4866 4.5005
R4397 DVDD.n5080 DVDD.n4866 4.5005
R4398 DVDD.n4869 DVDD.n4858 4.5005
R4399 DVDD.n5028 DVDD.n4858 4.5005
R4400 DVDD.n5082 DVDD.n4858 4.5005
R4401 DVDD.n5080 DVDD.n4858 4.5005
R4402 DVDD.n5080 DVDD.n4857 4.5005
R4403 DVDD.n5080 DVDD.n4867 4.5005
R4404 DVDD.n4869 DVDD.n4867 4.5005
R4405 DVDD.n5028 DVDD.n4867 4.5005
R4406 DVDD.n5082 DVDD.n4867 4.5005
R4407 DVDD.n4869 DVDD.n4857 4.5005
R4408 DVDD.n5028 DVDD.n4857 4.5005
R4409 DVDD.n5082 DVDD.n4857 4.5005
R4410 DVDD.n5082 DVDD.n5081 4.5005
R4411 DVDD.n5081 DVDD.n5028 4.5005
R4412 DVDD.n5081 DVDD.n4869 4.5005
R4413 DVDD.n5081 DVDD.n5080 4.5005
R4414 DVDD.n8938 DVDD.n583 4.5005
R4415 DVDD.n591 DVDD.n583 4.5005
R4416 DVDD.n589 DVDD.n583 4.5005
R4417 DVDD.n8936 DVDD.n583 4.5005
R4418 DVDD.n8938 DVDD.n581 4.5005
R4419 DVDD.n591 DVDD.n581 4.5005
R4420 DVDD.n589 DVDD.n581 4.5005
R4421 DVDD.n8936 DVDD.n581 4.5005
R4422 DVDD.n8936 DVDD.n577 4.5005
R4423 DVDD.n8936 DVDD.n587 4.5005
R4424 DVDD.n8936 DVDD.n578 4.5005
R4425 DVDD.n8938 DVDD.n584 4.5005
R4426 DVDD.n591 DVDD.n584 4.5005
R4427 DVDD.n589 DVDD.n584 4.5005
R4428 DVDD.n8936 DVDD.n584 4.5005
R4429 DVDD.n8938 DVDD.n580 4.5005
R4430 DVDD.n591 DVDD.n580 4.5005
R4431 DVDD.n589 DVDD.n580 4.5005
R4432 DVDD.n8936 DVDD.n580 4.5005
R4433 DVDD.n8938 DVDD.n585 4.5005
R4434 DVDD.n591 DVDD.n585 4.5005
R4435 DVDD.n589 DVDD.n585 4.5005
R4436 DVDD.n8936 DVDD.n585 4.5005
R4437 DVDD.n8936 DVDD.n586 4.5005
R4438 DVDD.n8936 DVDD.n579 4.5005
R4439 DVDD.n589 DVDD.n579 4.5005
R4440 DVDD.n591 DVDD.n579 4.5005
R4441 DVDD.n8938 DVDD.n579 4.5005
R4442 DVDD.n589 DVDD.n586 4.5005
R4443 DVDD.n591 DVDD.n586 4.5005
R4444 DVDD.n8938 DVDD.n586 4.5005
R4445 DVDD.n589 DVDD.n578 4.5005
R4446 DVDD.n591 DVDD.n578 4.5005
R4447 DVDD.n8938 DVDD.n578 4.5005
R4448 DVDD.n589 DVDD.n587 4.5005
R4449 DVDD.n591 DVDD.n587 4.5005
R4450 DVDD.n8938 DVDD.n587 4.5005
R4451 DVDD.n589 DVDD.n577 4.5005
R4452 DVDD.n591 DVDD.n577 4.5005
R4453 DVDD.n8938 DVDD.n577 4.5005
R4454 DVDD.n8938 DVDD.n8937 4.5005
R4455 DVDD.n8937 DVDD.n591 4.5005
R4456 DVDD.n8937 DVDD.n589 4.5005
R4457 DVDD.n8937 DVDD.n8936 4.5005
R4458 DVDD.n4821 DVDD.n4820 4.5005
R4459 DVDD.n4820 DVDD.n4593 4.5005
R4460 DVDD.n4820 DVDD.n4819 4.5005
R4461 DVDD.n4605 DVDD.n4593 4.5005
R4462 DVDD.n4819 DVDD.n4605 4.5005
R4463 DVDD.n4729 DVDD.n4593 4.5005
R4464 DVDD.n4819 DVDD.n4729 4.5005
R4465 DVDD.n4604 DVDD.n4593 4.5005
R4466 DVDD.n4819 DVDD.n4604 4.5005
R4467 DVDD.n4730 DVDD.n4593 4.5005
R4468 DVDD.n4819 DVDD.n4730 4.5005
R4469 DVDD.n4603 DVDD.n4593 4.5005
R4470 DVDD.n4819 DVDD.n4603 4.5005
R4471 DVDD.n4731 DVDD.n4593 4.5005
R4472 DVDD.n4819 DVDD.n4731 4.5005
R4473 DVDD.n4602 DVDD.n4593 4.5005
R4474 DVDD.n4819 DVDD.n4602 4.5005
R4475 DVDD.n4732 DVDD.n4593 4.5005
R4476 DVDD.n4819 DVDD.n4732 4.5005
R4477 DVDD.n4601 DVDD.n4593 4.5005
R4478 DVDD.n4819 DVDD.n4601 4.5005
R4479 DVDD.n4818 DVDD.n4593 4.5005
R4480 DVDD.n4818 DVDD.n4738 4.5005
R4481 DVDD.n4819 DVDD.n4818 4.5005
R4482 DVDD.n6775 DVDD.n2961 4.5005
R4483 DVDD.n6775 DVDD.n2962 4.5005
R4484 DVDD.n6775 DVDD.n6774 4.5005
R4485 DVDD.n2977 DVDD.n2962 4.5005
R4486 DVDD.n6774 DVDD.n2977 4.5005
R4487 DVDD.n2974 DVDD.n2962 4.5005
R4488 DVDD.n6774 DVDD.n2974 4.5005
R4489 DVDD.n2979 DVDD.n2962 4.5005
R4490 DVDD.n6774 DVDD.n2979 4.5005
R4491 DVDD.n2973 DVDD.n2962 4.5005
R4492 DVDD.n6774 DVDD.n2973 4.5005
R4493 DVDD.n2981 DVDD.n2962 4.5005
R4494 DVDD.n6774 DVDD.n2981 4.5005
R4495 DVDD.n2972 DVDD.n2962 4.5005
R4496 DVDD.n6774 DVDD.n2972 4.5005
R4497 DVDD.n2983 DVDD.n2962 4.5005
R4498 DVDD.n6774 DVDD.n2983 4.5005
R4499 DVDD.n2971 DVDD.n2962 4.5005
R4500 DVDD.n6774 DVDD.n2971 4.5005
R4501 DVDD.n2985 DVDD.n2962 4.5005
R4502 DVDD.n6774 DVDD.n2985 4.5005
R4503 DVDD.n2970 DVDD.n2962 4.5005
R4504 DVDD.n6774 DVDD.n2970 4.5005
R4505 DVDD.n2987 DVDD.n2962 4.5005
R4506 DVDD.n6774 DVDD.n2987 4.5005
R4507 DVDD.n2969 DVDD.n2962 4.5005
R4508 DVDD.n6774 DVDD.n2969 4.5005
R4509 DVDD.n2989 DVDD.n2962 4.5005
R4510 DVDD.n6774 DVDD.n2989 4.5005
R4511 DVDD.n2968 DVDD.n2962 4.5005
R4512 DVDD.n6774 DVDD.n2968 4.5005
R4513 DVDD.n2991 DVDD.n2962 4.5005
R4514 DVDD.n6774 DVDD.n2991 4.5005
R4515 DVDD.n2967 DVDD.n2962 4.5005
R4516 DVDD.n6774 DVDD.n2967 4.5005
R4517 DVDD.n2993 DVDD.n2962 4.5005
R4518 DVDD.n6774 DVDD.n2993 4.5005
R4519 DVDD.n2966 DVDD.n2962 4.5005
R4520 DVDD.n6774 DVDD.n2966 4.5005
R4521 DVDD.n2995 DVDD.n2962 4.5005
R4522 DVDD.n6774 DVDD.n2995 4.5005
R4523 DVDD.n2965 DVDD.n2962 4.5005
R4524 DVDD.n6774 DVDD.n2965 4.5005
R4525 DVDD.n2997 DVDD.n2962 4.5005
R4526 DVDD.n6774 DVDD.n2997 4.5005
R4527 DVDD.n2964 DVDD.n2962 4.5005
R4528 DVDD.n6774 DVDD.n2964 4.5005
R4529 DVDD.n6773 DVDD.n2961 4.5005
R4530 DVDD.n6773 DVDD.n2962 4.5005
R4531 DVDD.n6774 DVDD.n6773 4.5005
R4532 DVDD.n6772 DVDD.n3000 4.5005
R4533 DVDD.n6772 DVDD.n3001 4.5005
R4534 DVDD.n6772 DVDD.n6771 4.5005
R4535 DVDD.n3007 DVDD.n3001 4.5005
R4536 DVDD.n6771 DVDD.n3007 4.5005
R4537 DVDD.n3010 DVDD.n3001 4.5005
R4538 DVDD.n6771 DVDD.n3010 4.5005
R4539 DVDD.n3006 DVDD.n3001 4.5005
R4540 DVDD.n6771 DVDD.n3006 4.5005
R4541 DVDD.n3012 DVDD.n3001 4.5005
R4542 DVDD.n6771 DVDD.n3012 4.5005
R4543 DVDD.n3005 DVDD.n3001 4.5005
R4544 DVDD.n6771 DVDD.n3005 4.5005
R4545 DVDD.n3014 DVDD.n3001 4.5005
R4546 DVDD.n6771 DVDD.n3014 4.5005
R4547 DVDD.n3004 DVDD.n3001 4.5005
R4548 DVDD.n6771 DVDD.n3004 4.5005
R4549 DVDD.n3016 DVDD.n3001 4.5005
R4550 DVDD.n6771 DVDD.n3016 4.5005
R4551 DVDD.n3003 DVDD.n3001 4.5005
R4552 DVDD.n6771 DVDD.n3003 4.5005
R4553 DVDD.n6770 DVDD.n3001 4.5005
R4554 DVDD.n6770 DVDD.n3022 4.5005
R4555 DVDD.n6771 DVDD.n6770 4.5005
R4556 DVDD.n6769 DVDD.n3024 4.5005
R4557 DVDD.n6769 DVDD.n3025 4.5005
R4558 DVDD.n6769 DVDD.n6768 4.5005
R4559 DVDD.n3040 DVDD.n3025 4.5005
R4560 DVDD.n6768 DVDD.n3040 4.5005
R4561 DVDD.n3037 DVDD.n3025 4.5005
R4562 DVDD.n6768 DVDD.n3037 4.5005
R4563 DVDD.n3042 DVDD.n3025 4.5005
R4564 DVDD.n6768 DVDD.n3042 4.5005
R4565 DVDD.n3036 DVDD.n3025 4.5005
R4566 DVDD.n6768 DVDD.n3036 4.5005
R4567 DVDD.n3044 DVDD.n3025 4.5005
R4568 DVDD.n6768 DVDD.n3044 4.5005
R4569 DVDD.n3035 DVDD.n3025 4.5005
R4570 DVDD.n6768 DVDD.n3035 4.5005
R4571 DVDD.n3046 DVDD.n3025 4.5005
R4572 DVDD.n6768 DVDD.n3046 4.5005
R4573 DVDD.n3034 DVDD.n3025 4.5005
R4574 DVDD.n6768 DVDD.n3034 4.5005
R4575 DVDD.n3048 DVDD.n3025 4.5005
R4576 DVDD.n6768 DVDD.n3048 4.5005
R4577 DVDD.n3033 DVDD.n3025 4.5005
R4578 DVDD.n6768 DVDD.n3033 4.5005
R4579 DVDD.n3050 DVDD.n3025 4.5005
R4580 DVDD.n6768 DVDD.n3050 4.5005
R4581 DVDD.n3032 DVDD.n3025 4.5005
R4582 DVDD.n6768 DVDD.n3032 4.5005
R4583 DVDD.n3052 DVDD.n3025 4.5005
R4584 DVDD.n6768 DVDD.n3052 4.5005
R4585 DVDD.n3031 DVDD.n3025 4.5005
R4586 DVDD.n6768 DVDD.n3031 4.5005
R4587 DVDD.n3054 DVDD.n3025 4.5005
R4588 DVDD.n6768 DVDD.n3054 4.5005
R4589 DVDD.n3030 DVDD.n3025 4.5005
R4590 DVDD.n6768 DVDD.n3030 4.5005
R4591 DVDD.n3056 DVDD.n3025 4.5005
R4592 DVDD.n6768 DVDD.n3056 4.5005
R4593 DVDD.n3029 DVDD.n3025 4.5005
R4594 DVDD.n6768 DVDD.n3029 4.5005
R4595 DVDD.n3058 DVDD.n3025 4.5005
R4596 DVDD.n6768 DVDD.n3058 4.5005
R4597 DVDD.n3028 DVDD.n3025 4.5005
R4598 DVDD.n6768 DVDD.n3028 4.5005
R4599 DVDD.n3060 DVDD.n3025 4.5005
R4600 DVDD.n6768 DVDD.n3060 4.5005
R4601 DVDD.n3027 DVDD.n3025 4.5005
R4602 DVDD.n6768 DVDD.n3027 4.5005
R4603 DVDD.n6767 DVDD.n3024 4.5005
R4604 DVDD.n6767 DVDD.n3025 4.5005
R4605 DVDD.n6768 DVDD.n6767 4.5005
R4606 DVDD.n2597 DVDD.n2572 4.5005
R4607 DVDD.n7003 DVDD.n2572 4.5005
R4608 DVDD.n7005 DVDD.n2572 4.5005
R4609 DVDD.n7003 DVDD.n2574 4.5005
R4610 DVDD.n7005 DVDD.n2574 4.5005
R4611 DVDD.n7003 DVDD.n2571 4.5005
R4612 DVDD.n7005 DVDD.n2571 4.5005
R4613 DVDD.n7003 DVDD.n2575 4.5005
R4614 DVDD.n7005 DVDD.n2575 4.5005
R4615 DVDD.n7003 DVDD.n2570 4.5005
R4616 DVDD.n7005 DVDD.n2570 4.5005
R4617 DVDD.n7003 DVDD.n2576 4.5005
R4618 DVDD.n7005 DVDD.n2576 4.5005
R4619 DVDD.n7003 DVDD.n2569 4.5005
R4620 DVDD.n7005 DVDD.n2569 4.5005
R4621 DVDD.n7003 DVDD.n2577 4.5005
R4622 DVDD.n7005 DVDD.n2577 4.5005
R4623 DVDD.n7003 DVDD.n2568 4.5005
R4624 DVDD.n7005 DVDD.n2568 4.5005
R4625 DVDD.n7003 DVDD.n2578 4.5005
R4626 DVDD.n7005 DVDD.n2578 4.5005
R4627 DVDD.n7003 DVDD.n2567 4.5005
R4628 DVDD.n7005 DVDD.n2567 4.5005
R4629 DVDD.n7003 DVDD.n2579 4.5005
R4630 DVDD.n7005 DVDD.n2579 4.5005
R4631 DVDD.n7003 DVDD.n2566 4.5005
R4632 DVDD.n7005 DVDD.n2566 4.5005
R4633 DVDD.n7003 DVDD.n2580 4.5005
R4634 DVDD.n7005 DVDD.n2580 4.5005
R4635 DVDD.n7003 DVDD.n2565 4.5005
R4636 DVDD.n7005 DVDD.n2565 4.5005
R4637 DVDD.n7003 DVDD.n2581 4.5005
R4638 DVDD.n7005 DVDD.n2581 4.5005
R4639 DVDD.n7003 DVDD.n2564 4.5005
R4640 DVDD.n7005 DVDD.n2564 4.5005
R4641 DVDD.n7003 DVDD.n2582 4.5005
R4642 DVDD.n7005 DVDD.n2582 4.5005
R4643 DVDD.n7003 DVDD.n2563 4.5005
R4644 DVDD.n7005 DVDD.n2563 4.5005
R4645 DVDD.n7003 DVDD.n2583 4.5005
R4646 DVDD.n7005 DVDD.n2583 4.5005
R4647 DVDD.n7003 DVDD.n2562 4.5005
R4648 DVDD.n7005 DVDD.n2562 4.5005
R4649 DVDD.n7003 DVDD.n2584 4.5005
R4650 DVDD.n7005 DVDD.n2584 4.5005
R4651 DVDD.n7003 DVDD.n2561 4.5005
R4652 DVDD.n7005 DVDD.n2561 4.5005
R4653 DVDD.n7004 DVDD.n2597 4.5005
R4654 DVDD.n7004 DVDD.n7003 4.5005
R4655 DVDD.n7005 DVDD.n7004 4.5005
R4656 DVDD.n7592 DVDD.n2486 4.5005
R4657 DVDD.n2486 DVDD.n2472 4.5005
R4658 DVDD.n7590 DVDD.n2486 4.5005
R4659 DVDD.n7566 DVDD.n2472 4.5005
R4660 DVDD.n7590 DVDD.n7566 4.5005
R4661 DVDD.n2500 DVDD.n2472 4.5005
R4662 DVDD.n7590 DVDD.n2500 4.5005
R4663 DVDD.n7567 DVDD.n2472 4.5005
R4664 DVDD.n7590 DVDD.n7567 4.5005
R4665 DVDD.n2499 DVDD.n2472 4.5005
R4666 DVDD.n7590 DVDD.n2499 4.5005
R4667 DVDD.n7568 DVDD.n2472 4.5005
R4668 DVDD.n7590 DVDD.n7568 4.5005
R4669 DVDD.n2498 DVDD.n2472 4.5005
R4670 DVDD.n7590 DVDD.n2498 4.5005
R4671 DVDD.n7569 DVDD.n2472 4.5005
R4672 DVDD.n7590 DVDD.n7569 4.5005
R4673 DVDD.n2497 DVDD.n2472 4.5005
R4674 DVDD.n7590 DVDD.n2497 4.5005
R4675 DVDD.n7570 DVDD.n2472 4.5005
R4676 DVDD.n7590 DVDD.n7570 4.5005
R4677 DVDD.n2496 DVDD.n2472 4.5005
R4678 DVDD.n7590 DVDD.n2496 4.5005
R4679 DVDD.n7571 DVDD.n2472 4.5005
R4680 DVDD.n7590 DVDD.n7571 4.5005
R4681 DVDD.n2495 DVDD.n2472 4.5005
R4682 DVDD.n7590 DVDD.n2495 4.5005
R4683 DVDD.n7572 DVDD.n2472 4.5005
R4684 DVDD.n7590 DVDD.n7572 4.5005
R4685 DVDD.n2494 DVDD.n2472 4.5005
R4686 DVDD.n7590 DVDD.n2494 4.5005
R4687 DVDD.n7573 DVDD.n2472 4.5005
R4688 DVDD.n7590 DVDD.n7573 4.5005
R4689 DVDD.n2493 DVDD.n2472 4.5005
R4690 DVDD.n7590 DVDD.n2493 4.5005
R4691 DVDD.n7574 DVDD.n2472 4.5005
R4692 DVDD.n7590 DVDD.n7574 4.5005
R4693 DVDD.n2492 DVDD.n2472 4.5005
R4694 DVDD.n7590 DVDD.n2492 4.5005
R4695 DVDD.n7575 DVDD.n2472 4.5005
R4696 DVDD.n7590 DVDD.n7575 4.5005
R4697 DVDD.n2491 DVDD.n2472 4.5005
R4698 DVDD.n7590 DVDD.n2491 4.5005
R4699 DVDD.n7589 DVDD.n2472 4.5005
R4700 DVDD.n7590 DVDD.n7589 4.5005
R4701 DVDD.n2490 DVDD.n2472 4.5005
R4702 DVDD.n7590 DVDD.n2490 4.5005
R4703 DVDD.n7592 DVDD.n7591 4.5005
R4704 DVDD.n7591 DVDD.n2472 4.5005
R4705 DVDD.n7591 DVDD.n7590 4.5005
R4706 DVDD.n7106 DVDD.n2488 4.5005
R4707 DVDD.n7107 DVDD.n2488 4.5005
R4708 DVDD.n7285 DVDD.n2488 4.5005
R4709 DVDD.n7122 DVDD.n7107 4.5005
R4710 DVDD.n7285 DVDD.n7122 4.5005
R4711 DVDD.n7119 DVDD.n7107 4.5005
R4712 DVDD.n7285 DVDD.n7119 4.5005
R4713 DVDD.n7124 DVDD.n7107 4.5005
R4714 DVDD.n7285 DVDD.n7124 4.5005
R4715 DVDD.n7118 DVDD.n7107 4.5005
R4716 DVDD.n7285 DVDD.n7118 4.5005
R4717 DVDD.n7126 DVDD.n7107 4.5005
R4718 DVDD.n7285 DVDD.n7126 4.5005
R4719 DVDD.n7117 DVDD.n7107 4.5005
R4720 DVDD.n7285 DVDD.n7117 4.5005
R4721 DVDD.n7128 DVDD.n7107 4.5005
R4722 DVDD.n7285 DVDD.n7128 4.5005
R4723 DVDD.n7116 DVDD.n7107 4.5005
R4724 DVDD.n7285 DVDD.n7116 4.5005
R4725 DVDD.n7130 DVDD.n7107 4.5005
R4726 DVDD.n7285 DVDD.n7130 4.5005
R4727 DVDD.n7115 DVDD.n7107 4.5005
R4728 DVDD.n7285 DVDD.n7115 4.5005
R4729 DVDD.n7132 DVDD.n7107 4.5005
R4730 DVDD.n7285 DVDD.n7132 4.5005
R4731 DVDD.n7114 DVDD.n7107 4.5005
R4732 DVDD.n7285 DVDD.n7114 4.5005
R4733 DVDD.n7134 DVDD.n7107 4.5005
R4734 DVDD.n7285 DVDD.n7134 4.5005
R4735 DVDD.n7113 DVDD.n7107 4.5005
R4736 DVDD.n7281 DVDD.n7113 4.5005
R4737 DVDD.n7285 DVDD.n7113 4.5005
R4738 DVDD.n7135 DVDD.n7106 4.5005
R4739 DVDD.n7135 DVDD.n7107 4.5005
R4740 DVDD.n7281 DVDD.n7135 4.5005
R4741 DVDD.n7285 DVDD.n7135 4.5005
R4742 DVDD.n7112 DVDD.n7106 4.5005
R4743 DVDD.n7112 DVDD.n7107 4.5005
R4744 DVDD.n7281 DVDD.n7112 4.5005
R4745 DVDD.n7285 DVDD.n7112 4.5005
R4746 DVDD.n7202 DVDD.n7106 4.5005
R4747 DVDD.n7202 DVDD.n7107 4.5005
R4748 DVDD.n7281 DVDD.n7202 4.5005
R4749 DVDD.n7285 DVDD.n7202 4.5005
R4750 DVDD.n7111 DVDD.n7106 4.5005
R4751 DVDD.n7111 DVDD.n7107 4.5005
R4752 DVDD.n7285 DVDD.n7111 4.5005
R4753 DVDD.n7204 DVDD.n7107 4.5005
R4754 DVDD.n7285 DVDD.n7204 4.5005
R4755 DVDD.n7110 DVDD.n7107 4.5005
R4756 DVDD.n7285 DVDD.n7110 4.5005
R4757 DVDD.n7284 DVDD.n7107 4.5005
R4758 DVDD.n7285 DVDD.n7284 4.5005
R4759 DVDD.n7109 DVDD.n7107 4.5005
R4760 DVDD.n7285 DVDD.n7109 4.5005
R4761 DVDD.n7286 DVDD.n7106 4.5005
R4762 DVDD.n7286 DVDD.n7107 4.5005
R4763 DVDD.n7286 DVDD.n7285 4.5005
R4764 DVDD.n7304 DVDD.n7287 4.5005
R4765 DVDD.n7485 DVDD.n7287 4.5005
R4766 DVDD.n7487 DVDD.n7287 4.5005
R4767 DVDD.n7485 DVDD.n7103 4.5005
R4768 DVDD.n7487 DVDD.n7103 4.5005
R4769 DVDD.n7485 DVDD.n7288 4.5005
R4770 DVDD.n7487 DVDD.n7288 4.5005
R4771 DVDD.n7485 DVDD.n7102 4.5005
R4772 DVDD.n7487 DVDD.n7102 4.5005
R4773 DVDD.n7485 DVDD.n7289 4.5005
R4774 DVDD.n7487 DVDD.n7289 4.5005
R4775 DVDD.n7485 DVDD.n7101 4.5005
R4776 DVDD.n7487 DVDD.n7101 4.5005
R4777 DVDD.n7485 DVDD.n7290 4.5005
R4778 DVDD.n7487 DVDD.n7290 4.5005
R4779 DVDD.n7485 DVDD.n7100 4.5005
R4780 DVDD.n7487 DVDD.n7100 4.5005
R4781 DVDD.n7485 DVDD.n7291 4.5005
R4782 DVDD.n7487 DVDD.n7291 4.5005
R4783 DVDD.n7485 DVDD.n7099 4.5005
R4784 DVDD.n7487 DVDD.n7099 4.5005
R4785 DVDD.n7486 DVDD.n7485 4.5005
R4786 DVDD.n7486 DVDD.n7298 4.5005
R4787 DVDD.n7487 DVDD.n7486 4.5005
R4788 DVDD.n8383 DVDD.n1501 4.5005
R4789 DVDD.n8380 DVDD.n1501 4.5005
R4790 DVDD.n8383 DVDD.n1502 4.5005
R4791 DVDD.n8380 DVDD.n1502 4.5005
R4792 DVDD.n8379 DVDD.n1502 4.5005
R4793 DVDD.n7201 DVDD.n7192 4.5005
R4794 DVDD.n7198 DVDD.n7136 4.5005
R4795 DVDD.n7195 DVDD.n7136 4.5005
R4796 DVDD.n7192 DVDD.n7136 4.5005
R4797 DVDD.n7198 DVDD.n7194 4.5005
R4798 DVDD.n7195 DVDD.n7194 4.5005
R4799 DVDD.n7194 DVDD.n7192 4.5005
R4800 DVDD.n7200 DVDD.n7194 4.5005
R4801 DVDD.n7200 DVDD.n7136 4.5005
R4802 DVDD.n7201 DVDD.n7200 4.5005
R4803 DVDD.n8385 DVDD.n1502 4.5005
R4804 DVDD.n8385 DVDD.n1501 4.5005
R4805 DVDD.n8386 DVDD.n8385 4.5005
R4806 DVDD.n8388 DVDD.n1495 4.5005
R4807 DVDD.n8415 DVDD.n8404 4.5005
R4808 DVDD.n8388 DVDD.n8387 4.5005
R4809 DVDD.n8415 DVDD.n8414 4.5005
R4810 DVDD.n8577 DVDD.n1382 4.5005
R4811 DVDD.n8573 DVDD.n1382 4.5005
R4812 DVDD.n8557 DVDD.n1388 4.5005
R4813 DVDD.n8557 DVDD.n8556 4.5005
R4814 DVDD.n4817 DVDD.n4816 4.5005
R4815 DVDD.n4817 DVDD.n4741 4.5005
R4816 DVDD.n4817 DVDD.n4740 4.5005
R4817 DVDD.n4816 DVDD.n4747 4.5005
R4818 DVDD.n4747 DVDD.n4741 4.5005
R4819 DVDD.n4780 DVDD.n4741 4.5005
R4820 DVDD.n4787 DVDD.n4780 4.5005
R4821 DVDD.n4778 DVDD.n4741 4.5005
R4822 DVDD.n4787 DVDD.n4778 4.5005
R4823 DVDD.n4782 DVDD.n4741 4.5005
R4824 DVDD.n4787 DVDD.n4782 4.5005
R4825 DVDD.n4777 DVDD.n4741 4.5005
R4826 DVDD.n4787 DVDD.n4777 4.5005
R4827 DVDD.n4784 DVDD.n4741 4.5005
R4828 DVDD.n4787 DVDD.n4784 4.5005
R4829 DVDD.n4776 DVDD.n4741 4.5005
R4830 DVDD.n4787 DVDD.n4776 4.5005
R4831 DVDD.n4786 DVDD.n4741 4.5005
R4832 DVDD.n4787 DVDD.n4786 4.5005
R4833 DVDD.n4775 DVDD.n4741 4.5005
R4834 DVDD.n4787 DVDD.n4775 4.5005
R4835 DVDD.n4816 DVDD.n432 4.5005
R4836 DVDD.n4741 DVDD.n432 4.5005
R4837 DVDD.n4787 DVDD.n432 4.5005
R4838 DVDD.n32 DVDD.n20 4.5005
R4839 DVDD.n9674 DVDD.n32 4.5005
R4840 DVDD.n9672 DVDD.n32 4.5005
R4841 DVDD.n9674 DVDD.n29 4.5005
R4842 DVDD.n9672 DVDD.n29 4.5005
R4843 DVDD.n9674 DVDD.n35 4.5005
R4844 DVDD.n9672 DVDD.n35 4.5005
R4845 DVDD.n9674 DVDD.n28 4.5005
R4846 DVDD.n9672 DVDD.n28 4.5005
R4847 DVDD.n9674 DVDD.n38 4.5005
R4848 DVDD.n9672 DVDD.n38 4.5005
R4849 DVDD.n9674 DVDD.n27 4.5005
R4850 DVDD.n9672 DVDD.n27 4.5005
R4851 DVDD.n9674 DVDD.n41 4.5005
R4852 DVDD.n9672 DVDD.n41 4.5005
R4853 DVDD.n9674 DVDD.n26 4.5005
R4854 DVDD.n9672 DVDD.n26 4.5005
R4855 DVDD.n9674 DVDD.n44 4.5005
R4856 DVDD.n9672 DVDD.n44 4.5005
R4857 DVDD.n9674 DVDD.n25 4.5005
R4858 DVDD.n9672 DVDD.n25 4.5005
R4859 DVDD.n9674 DVDD.n9673 4.5005
R4860 DVDD.n9673 DVDD.n24 4.5005
R4861 DVDD.n9673 DVDD.n9672 4.5005
R4862 DVDD.n9693 DVDD.n9 4.5005
R4863 DVDD.n9691 DVDD.n9 4.5005
R4864 DVDD.n9693 DVDD.n8 4.5005
R4865 DVDD.n9691 DVDD.n8 4.5005
R4866 DVDD.n9693 DVDD.n10 4.5005
R4867 DVDD.n9691 DVDD.n10 4.5005
R4868 DVDD.n9693 DVDD.n7 4.5005
R4869 DVDD.n9691 DVDD.n7 4.5005
R4870 DVDD.n9693 DVDD.n11 4.5005
R4871 DVDD.n9691 DVDD.n11 4.5005
R4872 DVDD.n9693 DVDD.n6 4.5005
R4873 DVDD.n9691 DVDD.n6 4.5005
R4874 DVDD.n9693 DVDD.n12 4.5005
R4875 DVDD.n9691 DVDD.n12 4.5005
R4876 DVDD.n9693 DVDD.n5 4.5005
R4877 DVDD.n9691 DVDD.n5 4.5005
R4878 DVDD.n9693 DVDD.n13 4.5005
R4879 DVDD.n9691 DVDD.n13 4.5005
R4880 DVDD.n9693 DVDD.n4 4.5005
R4881 DVDD.n9691 DVDD.n4 4.5005
R4882 DVDD.n9693 DVDD.n9692 4.5005
R4883 DVDD.n9692 DVDD.n9691 4.5005
R4884 DVDD.n9284 DVDD.n9244 4.5005
R4885 DVDD.n9244 DVDD.n457 4.5005
R4886 DVDD.n9244 DVDD.n459 4.5005
R4887 DVDD.n9244 DVDD.n456 4.5005
R4888 DVDD.n9284 DVDD.n464 4.5005
R4889 DVDD.n464 DVDD.n457 4.5005
R4890 DVDD.n464 DVDD.n459 4.5005
R4891 DVDD.n464 DVDD.n456 4.5005
R4892 DVDD.n9283 DVDD.n457 4.5005
R4893 DVDD.n9283 DVDD.n459 4.5005
R4894 DVDD.n9283 DVDD.n456 4.5005
R4895 DVDD.n461 DVDD.n457 4.5005
R4896 DVDD.n461 DVDD.n459 4.5005
R4897 DVDD.n461 DVDD.n456 4.5005
R4898 DVDD.n9248 DVDD.n457 4.5005
R4899 DVDD.n9248 DVDD.n459 4.5005
R4900 DVDD.n9248 DVDD.n456 4.5005
R4901 DVDD.n462 DVDD.n457 4.5005
R4902 DVDD.n462 DVDD.n459 4.5005
R4903 DVDD.n462 DVDD.n456 4.5005
R4904 DVDD.n9284 DVDD.n9245 4.5005
R4905 DVDD.n9245 DVDD.n457 4.5005
R4906 DVDD.n9245 DVDD.n459 4.5005
R4907 DVDD.n9245 DVDD.n456 4.5005
R4908 DVDD.n9284 DVDD.n463 4.5005
R4909 DVDD.n463 DVDD.n457 4.5005
R4910 DVDD.n463 DVDD.n459 4.5005
R4911 DVDD.n463 DVDD.n456 4.5005
R4912 DVDD.n9284 DVDD.n9246 4.5005
R4913 DVDD.n9246 DVDD.n457 4.5005
R4914 DVDD.n9246 DVDD.n459 4.5005
R4915 DVDD.n9246 DVDD.n456 4.5005
R4916 DVDD.n9247 DVDD.n457 4.5005
R4917 DVDD.n9247 DVDD.n459 4.5005
R4918 DVDD.n9247 DVDD.n456 4.5005
R4919 DVDD.n9285 DVDD.n457 4.5005
R4920 DVDD.n9285 DVDD.n459 4.5005
R4921 DVDD.n9285 DVDD.n456 4.5005
R4922 DVDD.n9285 DVDD.n9284 4.5005
R4923 DVDD.n9284 DVDD.n9247 4.5005
R4924 DVDD.n9284 DVDD.n462 4.5005
R4925 DVDD.n9284 DVDD.n9248 4.5005
R4926 DVDD.n9284 DVDD.n461 4.5005
R4927 DVDD.n9284 DVDD.n9283 4.5005
R4928 DVDD.n9175 DVDD.n527 4.5005
R4929 DVDD.n534 DVDD.n527 4.5005
R4930 DVDD.n9173 DVDD.n527 4.5005
R4931 DVDD.n533 DVDD.n527 4.5005
R4932 DVDD.n9175 DVDD.n525 4.5005
R4933 DVDD.n534 DVDD.n525 4.5005
R4934 DVDD.n9173 DVDD.n525 4.5005
R4935 DVDD.n533 DVDD.n525 4.5005
R4936 DVDD.n9174 DVDD.n534 4.5005
R4937 DVDD.n9174 DVDD.n9173 4.5005
R4938 DVDD.n9174 DVDD.n533 4.5005
R4939 DVDD.n534 DVDD.n521 4.5005
R4940 DVDD.n9173 DVDD.n521 4.5005
R4941 DVDD.n533 DVDD.n521 4.5005
R4942 DVDD.n534 DVDD.n531 4.5005
R4943 DVDD.n9173 DVDD.n531 4.5005
R4944 DVDD.n533 DVDD.n531 4.5005
R4945 DVDD.n534 DVDD.n522 4.5005
R4946 DVDD.n9173 DVDD.n522 4.5005
R4947 DVDD.n533 DVDD.n522 4.5005
R4948 DVDD.n9175 DVDD.n528 4.5005
R4949 DVDD.n534 DVDD.n528 4.5005
R4950 DVDD.n9173 DVDD.n528 4.5005
R4951 DVDD.n533 DVDD.n528 4.5005
R4952 DVDD.n9175 DVDD.n524 4.5005
R4953 DVDD.n534 DVDD.n524 4.5005
R4954 DVDD.n9173 DVDD.n524 4.5005
R4955 DVDD.n533 DVDD.n524 4.5005
R4956 DVDD.n9175 DVDD.n529 4.5005
R4957 DVDD.n534 DVDD.n529 4.5005
R4958 DVDD.n9173 DVDD.n529 4.5005
R4959 DVDD.n533 DVDD.n529 4.5005
R4960 DVDD.n534 DVDD.n530 4.5005
R4961 DVDD.n9173 DVDD.n530 4.5005
R4962 DVDD.n533 DVDD.n530 4.5005
R4963 DVDD.n534 DVDD.n523 4.5005
R4964 DVDD.n9173 DVDD.n523 4.5005
R4965 DVDD.n533 DVDD.n523 4.5005
R4966 DVDD.n9175 DVDD.n523 4.5005
R4967 DVDD.n9175 DVDD.n530 4.5005
R4968 DVDD.n9175 DVDD.n522 4.5005
R4969 DVDD.n9175 DVDD.n531 4.5005
R4970 DVDD.n9175 DVDD.n521 4.5005
R4971 DVDD.n9175 DVDD.n9174 4.5005
R4972 DVDD.n4552 DVDD.n4543 4.5005
R4973 DVDD.n4552 DVDD.n4544 4.5005
R4974 DVDD.n4552 DVDD.n4542 4.5005
R4975 DVDD.n5249 DVDD.n4552 4.5005
R4976 DVDD.n4550 DVDD.n4543 4.5005
R4977 DVDD.n4550 DVDD.n4544 4.5005
R4978 DVDD.n4550 DVDD.n4542 4.5005
R4979 DVDD.n5249 DVDD.n4550 4.5005
R4980 DVDD.n4553 DVDD.n4543 4.5005
R4981 DVDD.n4553 DVDD.n4544 4.5005
R4982 DVDD.n4553 DVDD.n4542 4.5005
R4983 DVDD.n5249 DVDD.n4553 4.5005
R4984 DVDD.n4549 DVDD.n4543 4.5005
R4985 DVDD.n4549 DVDD.n4544 4.5005
R4986 DVDD.n4549 DVDD.n4542 4.5005
R4987 DVDD.n5249 DVDD.n4549 4.5005
R4988 DVDD.n4554 DVDD.n4543 4.5005
R4989 DVDD.n4554 DVDD.n4544 4.5005
R4990 DVDD.n4554 DVDD.n4542 4.5005
R4991 DVDD.n5249 DVDD.n4554 4.5005
R4992 DVDD.n4548 DVDD.n4543 4.5005
R4993 DVDD.n4548 DVDD.n4544 4.5005
R4994 DVDD.n4548 DVDD.n4542 4.5005
R4995 DVDD.n5249 DVDD.n4548 4.5005
R4996 DVDD.n4555 DVDD.n4543 4.5005
R4997 DVDD.n4555 DVDD.n4544 4.5005
R4998 DVDD.n4555 DVDD.n4542 4.5005
R4999 DVDD.n5249 DVDD.n4555 4.5005
R5000 DVDD.n4547 DVDD.n4543 4.5005
R5001 DVDD.n4547 DVDD.n4544 4.5005
R5002 DVDD.n4547 DVDD.n4542 4.5005
R5003 DVDD.n5249 DVDD.n4547 4.5005
R5004 DVDD.n5248 DVDD.n4543 4.5005
R5005 DVDD.n5248 DVDD.n4544 4.5005
R5006 DVDD.n5248 DVDD.n4542 4.5005
R5007 DVDD.n5249 DVDD.n5248 4.5005
R5008 DVDD.n4546 DVDD.n4543 4.5005
R5009 DVDD.n4546 DVDD.n4544 4.5005
R5010 DVDD.n4546 DVDD.n4542 4.5005
R5011 DVDD.n5249 DVDD.n4546 4.5005
R5012 DVDD.n5250 DVDD.n4543 4.5005
R5013 DVDD.n5250 DVDD.n4544 4.5005
R5014 DVDD.n5250 DVDD.n4542 4.5005
R5015 DVDD.n5250 DVDD.n5249 4.5005
R5016 DVDD.n9208 DVDD.n490 4.5005
R5017 DVDD.n496 DVDD.n490 4.5005
R5018 DVDD.n498 DVDD.n490 4.5005
R5019 DVDD.n9210 DVDD.n490 4.5005
R5020 DVDD.n9208 DVDD.n488 4.5005
R5021 DVDD.n496 DVDD.n488 4.5005
R5022 DVDD.n498 DVDD.n488 4.5005
R5023 DVDD.n9210 DVDD.n488 4.5005
R5024 DVDD.n496 DVDD.n491 4.5005
R5025 DVDD.n498 DVDD.n491 4.5005
R5026 DVDD.n9210 DVDD.n491 4.5005
R5027 DVDD.n9208 DVDD.n491 4.5005
R5028 DVDD.n496 DVDD.n487 4.5005
R5029 DVDD.n498 DVDD.n487 4.5005
R5030 DVDD.n9210 DVDD.n487 4.5005
R5031 DVDD.n9208 DVDD.n487 4.5005
R5032 DVDD.n496 DVDD.n492 4.5005
R5033 DVDD.n498 DVDD.n492 4.5005
R5034 DVDD.n9210 DVDD.n492 4.5005
R5035 DVDD.n9208 DVDD.n492 4.5005
R5036 DVDD.n9208 DVDD.n486 4.5005
R5037 DVDD.n496 DVDD.n486 4.5005
R5038 DVDD.n498 DVDD.n486 4.5005
R5039 DVDD.n9210 DVDD.n486 4.5005
R5040 DVDD.n9208 DVDD.n493 4.5005
R5041 DVDD.n496 DVDD.n493 4.5005
R5042 DVDD.n498 DVDD.n493 4.5005
R5043 DVDD.n9210 DVDD.n493 4.5005
R5044 DVDD.n9208 DVDD.n485 4.5005
R5045 DVDD.n496 DVDD.n485 4.5005
R5046 DVDD.n498 DVDD.n485 4.5005
R5047 DVDD.n9210 DVDD.n485 4.5005
R5048 DVDD.n9208 DVDD.n494 4.5005
R5049 DVDD.n496 DVDD.n494 4.5005
R5050 DVDD.n498 DVDD.n494 4.5005
R5051 DVDD.n9210 DVDD.n494 4.5005
R5052 DVDD.n496 DVDD.n484 4.5005
R5053 DVDD.n498 DVDD.n484 4.5005
R5054 DVDD.n9210 DVDD.n484 4.5005
R5055 DVDD.n9208 DVDD.n484 4.5005
R5056 DVDD.n9209 DVDD.n496 4.5005
R5057 DVDD.n9209 DVDD.n498 4.5005
R5058 DVDD.n9210 DVDD.n9209 4.5005
R5059 DVDD.n9209 DVDD.n9208 4.5005
R5060 DVDD.n66 DVDD.n55 4.5005
R5061 DVDD.n9647 DVDD.n66 4.5005
R5062 DVDD.n66 DVDD.n59 4.5005
R5063 DVDD.n73 DVDD.n66 4.5005
R5064 DVDD.n64 DVDD.n55 4.5005
R5065 DVDD.n9647 DVDD.n64 4.5005
R5066 DVDD.n64 DVDD.n59 4.5005
R5067 DVDD.n73 DVDD.n64 4.5005
R5068 DVDD.n9647 DVDD.n67 4.5005
R5069 DVDD.n67 DVDD.n59 4.5005
R5070 DVDD.n73 DVDD.n67 4.5005
R5071 DVDD.n67 DVDD.n55 4.5005
R5072 DVDD.n9647 DVDD.n63 4.5005
R5073 DVDD.n63 DVDD.n59 4.5005
R5074 DVDD.n73 DVDD.n63 4.5005
R5075 DVDD.n63 DVDD.n55 4.5005
R5076 DVDD.n9647 DVDD.n68 4.5005
R5077 DVDD.n68 DVDD.n59 4.5005
R5078 DVDD.n73 DVDD.n68 4.5005
R5079 DVDD.n68 DVDD.n55 4.5005
R5080 DVDD.n62 DVDD.n55 4.5005
R5081 DVDD.n9647 DVDD.n62 4.5005
R5082 DVDD.n62 DVDD.n59 4.5005
R5083 DVDD.n73 DVDD.n62 4.5005
R5084 DVDD.n69 DVDD.n55 4.5005
R5085 DVDD.n9647 DVDD.n69 4.5005
R5086 DVDD.n69 DVDD.n59 4.5005
R5087 DVDD.n73 DVDD.n69 4.5005
R5088 DVDD.n61 DVDD.n55 4.5005
R5089 DVDD.n9647 DVDD.n61 4.5005
R5090 DVDD.n61 DVDD.n59 4.5005
R5091 DVDD.n73 DVDD.n61 4.5005
R5092 DVDD.n70 DVDD.n55 4.5005
R5093 DVDD.n9647 DVDD.n70 4.5005
R5094 DVDD.n70 DVDD.n59 4.5005
R5095 DVDD.n73 DVDD.n70 4.5005
R5096 DVDD.n9647 DVDD.n60 4.5005
R5097 DVDD.n60 DVDD.n59 4.5005
R5098 DVDD.n73 DVDD.n60 4.5005
R5099 DVDD.n60 DVDD.n55 4.5005
R5100 DVDD.n9647 DVDD.n9646 4.5005
R5101 DVDD.n9646 DVDD.n59 4.5005
R5102 DVDD.n9646 DVDD.n73 4.5005
R5103 DVDD.n9646 DVDD.n55 4.5005
R5104 DVDD.t1 DVDD 4.04483
R5105 DVDD DVDD.t1 4.04483
R5106 DVDD.t7 DVDD 4.04483
R5107 DVDD DVDD.t7 4.04483
R5108 DVDD.t32 DVDD 4.04483
R5109 DVDD DVDD.t32 4.04483
R5110 DVDD.t33 DVDD 4.04483
R5111 DVDD DVDD.t33 4.04483
R5112 DVDD.t12 DVDD 4.04483
R5113 DVDD DVDD.t12 4.04483
R5114 DVDD.t40 DVDD 4.04483
R5115 DVDD DVDD.t40 4.04483
R5116 DVDD.t18 DVDD 4.04483
R5117 DVDD DVDD.t18 4.04483
R5118 DVDD.t28 DVDD 4.04483
R5119 DVDD DVDD.t28 4.04483
R5120 DVDD.t5 DVDD 4.04483
R5121 DVDD DVDD.t5 4.04483
R5122 DVDD.t9 DVDD 4.04483
R5123 DVDD DVDD.t9 4.04483
R5124 DVDD.t14 DVDD 4.04483
R5125 DVDD DVDD.t14 4.04483
R5126 DVDD DVDD.t38 4.04483
R5127 DVDD.t38 DVDD 4.04483
R5128 DVDD.t4 DVDD 4.04483
R5129 DVDD DVDD.t4 4.04483
R5130 DVDD.t19 DVDD 4.04483
R5131 DVDD DVDD.t19 4.04483
R5132 DVDD.t11 DVDD 4.04483
R5133 DVDD DVDD.t11 4.04483
R5134 DVDD.t20 DVDD 4.04483
R5135 DVDD DVDD.t20 4.04483
R5136 DVDD.t35 DVDD 4.04483
R5137 DVDD DVDD.t35 4.04483
R5138 DVDD.t16 DVDD 4.04483
R5139 DVDD DVDD.t16 4.04483
R5140 DVDD.n8389 DVDD.n1496 2.26366
R5141 DVDD.n96 DVDD.n81 2.2505
R5142 DVDD.n9628 DVDD.n83 2.2505
R5143 DVDD.n842 DVDD.n841 2.2505
R5144 DVDD.n9622 DVDD.n9621 2.2505
R5145 DVDD.n8771 DVDD.n94 2.2505
R5146 DVDD.n8766 DVDD.n849 2.2505
R5147 DVDD.n8761 DVDD.n8760 2.2505
R5148 DVDD.n941 DVDD.n857 2.2505
R5149 DVDD.n8755 DVDD.n8754 2.2505
R5150 DVDD.n933 DVDD.n863 2.2505
R5151 DVDD.n8748 DVDD.n8747 2.2505
R5152 DVDD.n8746 DVDD.n8745 2.2505
R5153 DVDD.n8725 DVDD.n877 2.2505
R5154 DVDD.n8739 DVDD.n881 2.2505
R5155 DVDD.n8734 DVDD.n8733 2.2505
R5156 DVDD.n8719 DVDD.n890 2.2505
R5157 DVDD.n8714 DVDD.n8713 2.2505
R5158 DVDD.n918 DVDD.n898 2.2505
R5159 DVDD.n996 DVDD.n917 2.2505
R5160 DVDD.n8708 DVDD.n8707 2.2505
R5161 DVDD.n8691 DVDD.n905 2.2505
R5162 DVDD.n8699 DVDD.n8698 2.2505
R5163 DVDD.n8697 DVDD.n1004 2.2505
R5164 DVDD.n1009 DVDD.n1006 2.2505
R5165 DVDD.n8688 DVDD.n8687 2.2505
R5166 DVDD.n8681 DVDD.n8680 2.2505
R5167 DVDD.n3741 DVDD.n1044 2.2505
R5168 DVDD.n3635 DVDD.n1048 2.2505
R5169 DVDD.n8672 DVDD.n8671 2.2505
R5170 DVDD.n3640 DVDD.n1046 2.2505
R5171 DVDD.n6327 DVDD.n6326 2.2505
R5172 DVDD.n6325 DVDD.n6324 2.2505
R5173 DVDD.n6321 DVDD.n6320 2.2505
R5174 DVDD.n3874 DVDD.n3868 2.2505
R5175 DVDD.n6315 DVDD.n6314 2.2505
R5176 DVDD.n6312 DVDD.n3876 2.2505
R5177 DVDD.n6310 DVDD.n6309 2.2505
R5178 DVDD.n6240 DVDD.n3879 2.2505
R5179 DVDD.n6304 DVDD.n6303 2.2505
R5180 DVDD.n6301 DVDD.n6239 2.2505
R5181 DVDD.n6299 DVDD.n6244 2.2505
R5182 DVDD.n6900 DVDD.n6899 2.2505
R5183 DVDD.n2783 DVDD.n2742 2.2505
R5184 DVDD.n6894 DVDD.n6893 2.2505
R5185 DVDD.n6890 DVDD.n2782 2.2505
R5186 DVDD.n6888 DVDD.n6887 2.2505
R5187 DVDD.n6875 DVDD.n2785 2.2505
R5188 DVDD.n6878 DVDD.n6877 2.2505
R5189 DVDD.n6873 DVDD.n6872 2.2505
R5190 DVDD.n6861 DVDD.n2793 2.2505
R5191 DVDD.n2798 DVDD.n2796 2.2505
R5192 DVDD.n6867 DVDD.n6866 2.2505
R5193 DVDD.n6778 DVDD.n6777 2.2505
R5194 DVDD.n6779 DVDD.n6778 2.2505
R5195 DVDD.n6781 DVDD.n2906 2.2505
R5196 DVDD.n6781 DVDD.n6780 2.2505
R5197 DVDD.n5303 DVDD.n2904 2.2505
R5198 DVDD.n2912 DVDD.n2904 2.2505
R5199 DVDD.n6787 DVDD.n2900 2.2505
R5200 DVDD.n6792 DVDD.n2891 2.2505
R5201 DVDD.n4512 DVDD.n2889 2.2505
R5202 DVDD.n5284 DVDD.n5283 2.2505
R5203 DVDD.n5283 DVDD.n5282 2.2505
R5204 DVDD.n4516 DVDD.n4509 2.2505
R5205 DVDD.n4515 DVDD.n4509 2.2505
R5206 DVDD.n5273 DVDD.n5272 2.2505
R5207 DVDD.n5274 DVDD.n5273 2.2505
R5208 DVDD.n5269 DVDD.n392 2.2505
R5209 DVDD.n4514 DVDD.n392 2.2505
R5210 DVDD.n9408 DVDD.n394 2.2505
R5211 DVDD.n9408 DVDD.n9407 2.2505
R5212 DVDD.n389 DVDD.n385 2.2505
R5213 DVDD.n395 DVDD.n389 2.2505
R5214 DVDD.n9414 DVDD.n388 2.2505
R5215 DVDD.n9402 DVDD.n382 2.2505
R5216 DVDD.n9400 DVDD.n9399 2.2505
R5217 DVDD.n9392 DVDD.n9391 2.2505
R5218 DVDD.n9392 DVDD.n175 2.2505
R5219 DVDD.n9586 DVDD.n9585 2.2505
R5220 DVDD.n9585 DVDD.n9584 2.2505
R5221 DVDD.n9590 DVDD.n164 2.2505
R5222 DVDD.n178 DVDD.n156 2.2505
R5223 DVDD.n9595 DVDD.n155 2.2505
R5224 DVDD.n9600 DVDD.n9599 2.2505
R5225 DVDD.n9601 DVDD.n9600 2.2505
R5226 DVDD.n145 DVDD.n144 2.2505
R5227 DVDD.n144 DVDD.n139 2.2505
R5228 DVDD.n9606 DVDD.n137 2.2505
R5229 DVDD.n9606 DVDD.n9605 2.2505
R5230 DVDD.n9349 DVDD.n133 2.2505
R5231 DVDD.n9612 DVDD.n132 2.2505
R5232 DVDD.n9361 DVDD.n9360 2.2505
R5233 DVDD.n9360 DVDD.n9359 2.2505
R5234 DVDD.n4528 DVDD.n444 2.2505
R5235 DVDD.n444 DVDD.n412 2.2505
R5236 DVDD.n9312 DVDD.n434 2.2505
R5237 DVDD.n9313 DVDD.n9312 2.2505
R5238 DVDD.n9316 DVDD.n9315 2.2505
R5239 DVDD.n9315 DVDD.n9314 2.2505
R5240 DVDD.n438 DVDD.n431 2.2505
R5241 DVDD.n9319 DVDD.n431 2.2505
R5242 DVDD.n9613 DVDD.n9612 2.2505
R5243 DVDD.n9327 DVDD.n133 2.2505
R5244 DVDD.n9596 DVDD.n9595 2.2505
R5245 DVDD.n156 DVDD.n152 2.2505
R5246 DVDD.n9590 DVDD.n9589 2.2505
R5247 DVDD.n9399 DVDD.n9398 2.2505
R5248 DVDD.n9418 DVDD.n382 2.2505
R5249 DVDD.n9415 DVDD.n9414 2.2505
R5250 DVDD.n5287 DVDD.n2889 2.2505
R5251 DVDD.n6792 DVDD.n6791 2.2505
R5252 DVDD.n6788 DVDD.n6787 2.2505
R5253 DVDD.n3580 DVDD.n3579 2.2505
R5254 DVDD.n3602 DVDD.n3601 2.2505
R5255 DVDD.n3603 DVDD.n3600 2.2505
R5256 DVDD.n3605 DVDD.n3604 2.2505
R5257 DVDD.n3606 DVDD.n3599 2.2505
R5258 DVDD.n3608 DVDD.n3607 2.2505
R5259 DVDD.n3609 DVDD.n3598 2.2505
R5260 DVDD.n3611 DVDD.n3610 2.2505
R5261 DVDD.n3612 DVDD.n3597 2.2505
R5262 DVDD.n3614 DVDD.n3613 2.2505
R5263 DVDD.n3615 DVDD.n3596 2.2505
R5264 DVDD.n3617 DVDD.n3616 2.2505
R5265 DVDD.n3618 DVDD.n3595 2.2505
R5266 DVDD.n3620 DVDD.n3619 2.2505
R5267 DVDD.n3621 DVDD.n3594 2.2505
R5268 DVDD.n3623 DVDD.n3622 2.2505
R5269 DVDD.n3624 DVDD.n3593 2.2505
R5270 DVDD.n3626 DVDD.n3625 2.2505
R5271 DVDD.n3627 DVDD.n3592 2.2505
R5272 DVDD.n3630 DVDD.n3629 2.2505
R5273 DVDD.n3632 DVDD.n3631 2.2505
R5274 DVDD.n3584 DVDD.n3583 2.2505
R5275 DVDD.n3745 DVDD.n3744 2.2505
R5276 DVDD.n3747 DVDD.n3746 2.2505
R5277 DVDD.n3750 DVDD.n3749 2.2505
R5278 DVDD.n3752 DVDD.n3751 2.2505
R5279 DVDD.n993 DVDD.n913 2.2505
R5280 DVDD.n992 DVDD.n991 2.2505
R5281 DVDD.n990 DVDD.n989 2.2505
R5282 DVDD.n988 DVDD.n987 2.2505
R5283 DVDD.n986 DVDD.n985 2.2505
R5284 DVDD.n984 DVDD.n983 2.2505
R5285 DVDD.n982 DVDD.n981 2.2505
R5286 DVDD.n980 DVDD.n979 2.2505
R5287 DVDD.n956 DVDD.n921 2.2505
R5288 DVDD.n954 DVDD.n953 2.2505
R5289 DVDD.n952 DVDD.n951 2.2505
R5290 DVDD.n950 DVDD.n922 2.2505
R5291 DVDD.n949 DVDD.n948 2.2505
R5292 DVDD.n947 DVDD.n946 2.2505
R5293 DVDD.n945 DVDD.n944 2.2505
R5294 DVDD.n929 DVDD.n928 2.2505
R5295 DVDD.n927 DVDD.n926 2.2505
R5296 DVDD.n925 DVDD.n924 2.2505
R5297 DVDD.n840 DVDD.n839 2.2505
R5298 DVDD.n8775 DVDD.n8774 2.2505
R5299 DVDD.n8777 DVDD.n8776 2.2505
R5300 DVDD.n8780 DVDD.n8779 2.2505
R5301 DVDD.n8791 DVDD.n8790 2.2505
R5302 DVDD.n8792 DVDD.n838 2.2505
R5303 DVDD.n8794 DVDD.n8793 2.2505
R5304 DVDD.n1001 DVDD.n1000 2.2505
R5305 DVDD.n837 DVDD.n791 2.2505
R5306 DVDD.n836 DVDD.n835 2.2505
R5307 DVDD.n834 DVDD.n792 2.2505
R5308 DVDD.n833 DVDD.n832 2.2505
R5309 DVDD.n831 DVDD.n793 2.2505
R5310 DVDD.n830 DVDD.n829 2.2505
R5311 DVDD.n828 DVDD.n15 2.2505
R5312 DVDD.n827 DVDD.n14 2.2505
R5313 DVDD.n826 DVDD.n825 2.2505
R5314 DVDD.n824 DVDD.n823 2.2505
R5315 DVDD.n822 DVDD.n821 2.2505
R5316 DVDD.n820 DVDD.n819 2.2505
R5317 DVDD.n818 DVDD.n817 2.2505
R5318 DVDD.n816 DVDD.n815 2.2505
R5319 DVDD.n814 DVDD.n813 2.2505
R5320 DVDD.n812 DVDD.n811 2.2505
R5321 DVDD.n810 DVDD.n809 2.2505
R5322 DVDD.n808 DVDD.n807 2.2505
R5323 DVDD.n806 DVDD.n794 2.2505
R5324 DVDD.n805 DVDD.n804 2.2505
R5325 DVDD.n803 DVDD.n795 2.2505
R5326 DVDD.n802 DVDD.n801 2.2505
R5327 DVDD.n800 DVDD.n796 2.2505
R5328 DVDD.n799 DVDD.n798 2.2505
R5329 DVDD.n797 DVDD.n790 2.2505
R5330 DVDD.n8796 DVDD.n8795 2.2505
R5331 DVDD.n8840 DVDD.n8839 2.2505
R5332 DVDD.n8841 DVDD.n671 2.2505
R5333 DVDD.n8843 DVDD.n8842 2.2505
R5334 DVDD.n8844 DVDD.n670 2.2505
R5335 DVDD.n8846 DVDD.n8845 2.2505
R5336 DVDD.n8847 DVDD.n669 2.2505
R5337 DVDD.n8849 DVDD.n8848 2.2505
R5338 DVDD.n8850 DVDD.n668 2.2505
R5339 DVDD.n8852 DVDD.n8851 2.2505
R5340 DVDD.n8853 DVDD.n667 2.2505
R5341 DVDD.n8855 DVDD.n8854 2.2505
R5342 DVDD.n8856 DVDD.n666 2.2505
R5343 DVDD.n8858 DVDD.n8857 2.2505
R5344 DVDD.n8859 DVDD.n665 2.2505
R5345 DVDD.n8861 DVDD.n8860 2.2505
R5346 DVDD.n8862 DVDD.n664 2.2505
R5347 DVDD.n8864 DVDD.n8863 2.2505
R5348 DVDD.n8865 DVDD.n663 2.2505
R5349 DVDD.n8867 DVDD.n8866 2.2505
R5350 DVDD.n8868 DVDD.n662 2.2505
R5351 DVDD.n8870 DVDD.n8869 2.2505
R5352 DVDD.n8871 DVDD.n661 2.2505
R5353 DVDD.n8873 DVDD.n8872 2.2505
R5354 DVDD.n8874 DVDD.n660 2.2505
R5355 DVDD.n8876 DVDD.n8875 2.2505
R5356 DVDD.n8838 DVDD.n672 2.2505
R5357 DVDD.n8789 DVDD.n8788 2.2505
R5358 DVDD.n9627 DVDD.n86 2.2505
R5359 DVDD.n8778 DVDD.n85 2.2505
R5360 DVDD.n9623 DVDD.n90 2.2505
R5361 DVDD.n8773 DVDD.n8772 2.2505
R5362 DVDD.n9616 DVDD.n115 2.2505
R5363 DVDD.n8765 DVDD.n851 2.2505
R5364 DVDD.n8762 DVDD.n854 2.2505
R5365 DVDD.n943 DVDD.n942 2.2505
R5366 DVDD.n8753 DVDD.n868 2.2505
R5367 DVDD.n923 DVDD.n867 2.2505
R5368 DVDD.n8749 DVDD.n872 2.2505
R5369 DVDD.n955 DVDD.n871 2.2505
R5370 DVDD.n978 DVDD.n977 2.2505
R5371 DVDD.n8738 DVDD.n884 2.2505
R5372 DVDD.n8735 DVDD.n886 2.2505
R5373 DVDD.n9425 DVDD.n350 2.2505
R5374 DVDD.n8718 DVDD.n892 2.2505
R5375 DVDD.n8715 DVDD.n895 2.2505
R5376 DVDD.n920 DVDD.n919 2.2505
R5377 DVDD.n995 DVDD.n994 2.2505
R5378 DVDD.n8706 DVDD.n908 2.2505
R5379 DVDD.n8703 DVDD.n8702 2.2505
R5380 DVDD.n8701 DVDD.n8700 2.2505
R5381 DVDD.n1003 DVDD.n1002 2.2505
R5382 DVDD.n1034 DVDD.n1033 2.2505
R5383 DVDD.n8686 DVDD.n1013 2.2505
R5384 DVDD.n3748 DVDD.n228 2.2505
R5385 DVDD.n8682 DVDD.n1039 2.2505
R5386 DVDD.n3743 DVDD.n3742 2.2505
R5387 DVDD.n3634 DVDD.n3633 2.2505
R5388 DVDD.n8670 DVDD.n1053 2.2505
R5389 DVDD.n3628 DVDD.n1052 2.2505
R5390 DVDD.n8788 DVDD.n81 2.2505
R5391 DVDD.n9628 DVDD.n9627 2.2505
R5392 DVDD.n842 DVDD.n85 2.2505
R5393 DVDD.n9623 DVDD.n9622 2.2505
R5394 DVDD.n8772 DVDD.n8771 2.2505
R5395 DVDD.n8766 DVDD.n8765 2.2505
R5396 DVDD.n8762 DVDD.n8761 2.2505
R5397 DVDD.n942 DVDD.n941 2.2505
R5398 DVDD.n8754 DVDD.n8753 2.2505
R5399 DVDD.n933 DVDD.n867 2.2505
R5400 DVDD.n8749 DVDD.n8748 2.2505
R5401 DVDD.n8745 DVDD.n871 2.2505
R5402 DVDD.n977 DVDD.n877 2.2505
R5403 DVDD.n8739 DVDD.n8738 2.2505
R5404 DVDD.n8735 DVDD.n8734 2.2505
R5405 DVDD.n8719 DVDD.n8718 2.2505
R5406 DVDD.n8715 DVDD.n8714 2.2505
R5407 DVDD.n919 DVDD.n918 2.2505
R5408 DVDD.n996 DVDD.n995 2.2505
R5409 DVDD.n8707 DVDD.n8706 2.2505
R5410 DVDD.n8703 DVDD.n905 2.2505
R5411 DVDD.n8700 DVDD.n8699 2.2505
R5412 DVDD.n1004 DVDD.n1003 2.2505
R5413 DVDD.n1034 DVDD.n1009 2.2505
R5414 DVDD.n8687 DVDD.n8686 2.2505
R5415 DVDD.n8682 DVDD.n8681 2.2505
R5416 DVDD.n3742 DVDD.n3741 2.2505
R5417 DVDD.n3635 DVDD.n3634 2.2505
R5418 DVDD.n8671 DVDD.n8670 2.2505
R5419 DVDD.n3640 DVDD.n1052 2.2505
R5420 DVDD.n8452 DVDD.n8446 2.2505
R5421 DVDD.n8454 DVDD.n8453 2.2505
R5422 DVDD.n8455 DVDD.n8445 2.2505
R5423 DVDD.n8457 DVDD.n8456 2.2505
R5424 DVDD.n8458 DVDD.n1338 2.2505
R5425 DVDD.n8460 DVDD.n8459 2.2505
R5426 DVDD.n8461 DVDD.n8444 2.2505
R5427 DVDD.n8463 DVDD.n8462 2.2505
R5428 DVDD.n8464 DVDD.n1445 2.2505
R5429 DVDD.n8470 DVDD.n8469 2.2505
R5430 DVDD.n8471 DVDD.n1443 2.2505
R5431 DVDD.n8473 DVDD.n8472 2.2505
R5432 DVDD.n8474 DVDD.n1442 2.2505
R5433 DVDD.n8476 DVDD.n8475 2.2505
R5434 DVDD.n8477 DVDD.n1441 2.2505
R5435 DVDD.n8479 DVDD.n8478 2.2505
R5436 DVDD.n8480 DVDD.n1440 2.2505
R5437 DVDD.n8482 DVDD.n8481 2.2505
R5438 DVDD.n8488 DVDD.n8487 2.2505
R5439 DVDD.n8486 DVDD.n8483 2.2505
R5440 DVDD.n8485 DVDD.n8484 2.2505
R5441 DVDD.n1346 DVDD.n1344 2.2505
R5442 DVDD.n8614 DVDD.n8613 2.2505
R5443 DVDD.n8612 DVDD.n1345 2.2505
R5444 DVDD.n8611 DVDD.n8610 2.2505
R5445 DVDD.n8609 DVDD.n1347 2.2505
R5446 DVDD.n8608 DVDD.n8607 2.2505
R5447 DVDD.n8530 DVDD.n8529 2.2505
R5448 DVDD.n8528 DVDD.n8524 2.2505
R5449 DVDD.n8527 DVDD.n8526 2.2505
R5450 DVDD.n8525 DVDD.n1351 2.2505
R5451 DVDD.n8551 DVDD.n8550 2.2505
R5452 DVDD.n8552 DVDD.n1395 2.2505
R5453 DVDD.n8554 DVDD.n8553 2.2505
R5454 DVDD.n8555 DVDD.n1389 2.2505
R5455 DVDD.n8560 DVDD.n8559 2.2505
R5456 DVDD.n8561 DVDD.n1387 2.2505
R5457 DVDD.n8563 DVDD.n8562 2.2505
R5458 DVDD.n8564 DVDD.n1386 2.2505
R5459 DVDD.n8566 DVDD.n8565 2.2505
R5460 DVDD.n8567 DVDD.n1385 2.2505
R5461 DVDD.n8569 DVDD.n8568 2.2505
R5462 DVDD.n8570 DVDD.n1384 2.2505
R5463 DVDD.n8572 DVDD.n8571 2.2505
R5464 DVDD.n8579 DVDD.n8578 2.2505
R5465 DVDD.n8580 DVDD.n1380 2.2505
R5466 DVDD.n8582 DVDD.n8581 2.2505
R5467 DVDD.n8583 DVDD.n1378 2.2505
R5468 DVDD.n8585 DVDD.n8584 2.2505
R5469 DVDD.n1379 DVDD.n1377 2.2505
R5470 DVDD.n8410 DVDD.n8409 2.2505
R5471 DVDD.n8411 DVDD.n8408 2.2505
R5472 DVDD.n8413 DVDD.n8412 2.2505
R5473 DVDD.n8403 DVDD.n8402 2.2505
R5474 DVDD.n8401 DVDD.n1491 2.2505
R5475 DVDD.n8400 DVDD.n8399 2.2505
R5476 DVDD.n8398 DVDD.n1492 2.2505
R5477 DVDD.n8397 DVDD.n8396 2.2505
R5478 DVDD.n8395 DVDD.n1493 2.2505
R5479 DVDD.n8394 DVDD.n8393 2.2505
R5480 DVDD.n8392 DVDD.n1494 2.2505
R5481 DVDD.n8391 DVDD.n8390 2.2505
R5482 DVDD.n8534 DVDD.n8533 2.24623
R5483 DVDD.n1325 DVDD.n1322 2.24623
R5484 DVDD.n1449 DVDD.n1447 2.24623
R5485 DVDD.n8436 DVDD.n1448 2.24623
R5486 DVDD.n1435 DVDD.n1433 2.24623
R5487 DVDD.n1431 DVDD.n1430 2.24623
R5488 DVDD.n1358 DVDD.n1355 2.24623
R5489 DVDD.n1359 DVDD.n1357 2.24623
R5490 DVDD.n8521 DVDD.n8518 2.24623
R5491 DVDD.n1331 DVDD.n1329 2.24623
R5492 DVDD.n1454 DVDD.n1452 2.24623
R5493 DVDD.n8431 DVDD.n1453 2.24623
R5494 DVDD.n1427 DVDD.n1425 2.24623
R5495 DVDD.n1423 DVDD.n1422 2.24623
R5496 DVDD.n1367 DVDD.n1364 2.24623
R5497 DVDD.n1368 DVDD.n1366 2.24623
R5498 DVDD.n7737 DVDD.n2332 2.24623
R5499 DVDD.n7730 DVDD.n2340 2.24623
R5500 DVDD.n7739 DVDD.n7738 2.24623
R5501 DVDD.n7731 DVDD.n2338 2.24623
R5502 DVDD.n2364 DVDD.n2363 2.24623
R5503 DVDD.n2365 DVDD.n2361 2.24623
R5504 DVDD.n1405 DVDD.n1403 2.24623
R5505 DVDD.n7355 DVDD.n7346 2.24623
R5506 DVDD.n8425 DVDD.n1459 2.24623
R5507 DVDD.n8424 DVDD.n8423 2.24623
R5508 DVDD.n1420 DVDD.n1419 2.24623
R5509 DVDD.n1417 DVDD.n1412 2.24623
R5510 DVDD.n8510 DVDD.n8509 2.24623
R5511 DVDD.n1411 DVDD.n1406 2.24623
R5512 DVDD.n2371 DVDD.n2358 2.24623
R5513 DVDD.n7681 DVDD.n2356 2.24623
R5514 DVDD.n1399 DVDD.n1397 2.24623
R5515 DVDD.n7351 DVDD.n7350 2.24623
R5516 DVDD.n1466 DVDD.n1463 2.24623
R5517 DVDD.n1467 DVDD.n1465 2.24623
R5518 DVDD.n1472 DVDD.n1468 2.24623
R5519 DVDD.n1473 DVDD.n1470 2.24623
R5520 DVDD.n1478 DVDD.n1474 2.24623
R5521 DVDD.n1479 DVDD.n1476 2.24623
R5522 DVDD.n8447 DVDD.n1326 2.24623
R5523 DVDD.n8465 DVDD.n8441 2.24623
R5524 DVDD.n8467 DVDD.n8443 2.24623
R5525 DVDD.n8442 DVDD.n8441 2.24623
R5526 DVDD.n8493 DVDD.n8492 2.24623
R5527 DVDD.n8490 DVDD.n1439 2.24623
R5528 DVDD.n8493 DVDD.n1437 2.24623
R5529 DVDD.n8602 DVDD.n1349 2.24623
R5530 DVDD.n8605 DVDD.n1350 2.24623
R5531 DVDD.n8603 DVDD.n8602 2.24623
R5532 DVDD.n8415 DVDD.n1490 2.24623
R5533 DVDD.n8575 DVDD.n1382 2.24623
R5534 DVDD.n8557 DVDD.n1392 2.24623
R5535 DVDD.n1394 DVDD.n1390 2.24623
R5536 DVDD.n1391 DVDD.n1390 2.24623
R5537 DVDD.n8574 DVDD.n1383 2.24623
R5538 DVDD.n8576 DVDD.n1383 2.24623
R5539 DVDD.n8407 DVDD.n8406 2.24623
R5540 DVDD.n8406 DVDD.n8405 2.24623
R5541 DVDD.n5417 DVDD.n4471 2.24552
R5542 DVDD.n5418 DVDD.n4470 2.24552
R5543 DVDD.n5420 DVDD.n4471 2.24552
R5544 DVDD.n5651 DVDD.n5483 2.24552
R5545 DVDD.n5659 DVDD.n4462 2.24552
R5546 DVDD.n5653 DVDD.n5483 2.24552
R5547 DVDD.n5659 DVDD.n4461 2.24552
R5548 DVDD.n5655 DVDD.n5483 2.24552
R5549 DVDD.n5659 DVDD.n4460 2.24552
R5550 DVDD.n5551 DVDD.n5492 2.24552
R5551 DVDD.n5553 DVDD.n5493 2.24552
R5552 DVDD.n5554 DVDD.n5492 2.24552
R5553 DVDD.n5556 DVDD.n5493 2.24552
R5554 DVDD.n5557 DVDD.n5492 2.24552
R5555 DVDD.n5559 DVDD.n5493 2.24552
R5556 DVDD.n2544 DVDD.n2522 2.24552
R5557 DVDD.n7020 DVDD.n7018 2.24552
R5558 DVDD.n2546 DVDD.n2521 2.24552
R5559 DVDD.n7020 DVDD.n7019 2.24552
R5560 DVDD.n2548 DVDD.n2521 2.24552
R5561 DVDD.n7021 DVDD.n7020 2.24552
R5562 DVDD.n7022 DVDD.n2521 2.24552
R5563 DVDD.n7020 DVDD.n2520 2.24552
R5564 DVDD.n7545 DVDD.n7535 2.24552
R5565 DVDD.n7550 DVDD.n2519 2.24552
R5566 DVDD.n7545 DVDD.n7536 2.24552
R5567 DVDD.n7550 DVDD.n2518 2.24552
R5568 DVDD.n7545 DVDD.n7537 2.24552
R5569 DVDD.n7550 DVDD.n2517 2.24552
R5570 DVDD.n7545 DVDD.n7538 2.24552
R5571 DVDD.n7550 DVDD.n2516 2.24552
R5572 DVDD.n7545 DVDD.n7539 2.24552
R5573 DVDD.n7550 DVDD.n2515 2.24552
R5574 DVDD.n7545 DVDD.n7540 2.24552
R5575 DVDD.n7550 DVDD.n2514 2.24552
R5576 DVDD.n7545 DVDD.n7541 2.24552
R5577 DVDD.n7550 DVDD.n2513 2.24552
R5578 DVDD.n7545 DVDD.n7542 2.24552
R5579 DVDD.n7550 DVDD.n2512 2.24552
R5580 DVDD.n7545 DVDD.n7543 2.24552
R5581 DVDD.n7550 DVDD.n2511 2.24552
R5582 DVDD.n7545 DVDD.n7544 2.24552
R5583 DVDD.n7550 DVDD.n2510 2.24552
R5584 DVDD.n7546 DVDD.n7545 2.24552
R5585 DVDD.n7550 DVDD.n2509 2.24552
R5586 DVDD.n7545 DVDD.n7027 2.24552
R5587 DVDD.n7222 DVDD.n7028 2.24552
R5588 DVDD.n7044 DVDD.n7029 2.24552
R5589 DVDD.n7222 DVDD.n7212 2.24552
R5590 DVDD.n7046 DVDD.n7029 2.24552
R5591 DVDD.n7222 DVDD.n7213 2.24552
R5592 DVDD.n7048 DVDD.n7029 2.24552
R5593 DVDD.n7222 DVDD.n7214 2.24552
R5594 DVDD.n7050 DVDD.n7029 2.24552
R5595 DVDD.n7222 DVDD.n7215 2.24552
R5596 DVDD.n7052 DVDD.n7029 2.24552
R5597 DVDD.n7222 DVDD.n7216 2.24552
R5598 DVDD.n7054 DVDD.n7029 2.24552
R5599 DVDD.n7222 DVDD.n7217 2.24552
R5600 DVDD.n7056 DVDD.n7029 2.24552
R5601 DVDD.n7222 DVDD.n7218 2.24552
R5602 DVDD.n7058 DVDD.n7029 2.24552
R5603 DVDD.n7222 DVDD.n7219 2.24552
R5604 DVDD.n7060 DVDD.n7029 2.24552
R5605 DVDD.n7222 DVDD.n7220 2.24552
R5606 DVDD.n7062 DVDD.n7029 2.24552
R5607 DVDD.n7222 DVDD.n7221 2.24552
R5608 DVDD.n7064 DVDD.n7029 2.24552
R5609 DVDD.n7222 DVDD.n7066 2.24552
R5610 DVDD.n3806 DVDD.n3560 2.24552
R5611 DVDD.n6334 DVDD.n3573 2.24552
R5612 DVDD.n3571 DVDD.n3560 2.24552
R5613 DVDD.n3875 DVDD.n3862 2.24552
R5614 DVDD.n6313 DVDD.n3864 2.24552
R5615 DVDD.n6311 DVDD.n3862 2.24552
R5616 DVDD.n3877 DVDD.n3864 2.24552
R5617 DVDD.n6241 DVDD.n3862 2.24552
R5618 DVDD.n6302 DVDD.n3864 2.24552
R5619 DVDD.n3362 DVDD.n3361 2.24552
R5620 DVDD.n6648 DVDD.n6645 2.24552
R5621 DVDD.n3362 DVDD.n3360 2.24552
R5622 DVDD.n6648 DVDD.n6646 2.24552
R5623 DVDD.n3362 DVDD.n3359 2.24552
R5624 DVDD.n6648 DVDD.n6647 2.24552
R5625 DVDD.n7886 DVDD.n2104 2.24552
R5626 DVDD.n7893 DVDD.n2091 2.24552
R5627 DVDD.n7886 DVDD.n2103 2.24552
R5628 DVDD.n7893 DVDD.n2092 2.24552
R5629 DVDD.n7887 DVDD.n7886 2.24552
R5630 DVDD.n7893 DVDD.n2093 2.24552
R5631 DVDD.n7886 DVDD.n2095 2.24552
R5632 DVDD.n7893 DVDD.n7892 2.24552
R5633 DVDD.n8056 DVDD.n1955 2.24552
R5634 DVDD.n8052 DVDD.n1987 2.24552
R5635 DVDD.n8056 DVDD.n1956 2.24552
R5636 DVDD.n8052 DVDD.n1986 2.24552
R5637 DVDD.n8056 DVDD.n1957 2.24552
R5638 DVDD.n8056 DVDD.n1952 2.24552
R5639 DVDD.n8052 DVDD.n8050 2.24552
R5640 DVDD.n8056 DVDD.n1951 2.24552
R5641 DVDD.n8052 DVDD.n8051 2.24552
R5642 DVDD.n8056 DVDD.n1950 2.24552
R5643 DVDD.n8056 DVDD.n1959 2.24552
R5644 DVDD.n8052 DVDD.n1985 2.24552
R5645 DVDD.n8056 DVDD.n1960 2.24552
R5646 DVDD.n8052 DVDD.n1984 2.24552
R5647 DVDD.n8056 DVDD.n1961 2.24552
R5648 DVDD.n8056 DVDD.n1948 2.24552
R5649 DVDD.n8052 DVDD.n1962 2.24552
R5650 DVDD.n8115 DVDD.n8109 2.24552
R5651 DVDD.n8120 DVDD.n1863 2.24552
R5652 DVDD.n8115 DVDD.n8110 2.24552
R5653 DVDD.n8120 DVDD.n1862 2.24552
R5654 DVDD.n8115 DVDD.n8111 2.24552
R5655 DVDD.n8115 DVDD.n8112 2.24552
R5656 DVDD.n8120 DVDD.n1859 2.24552
R5657 DVDD.n8115 DVDD.n8113 2.24552
R5658 DVDD.n8120 DVDD.n1858 2.24552
R5659 DVDD.n8115 DVDD.n8114 2.24552
R5660 DVDD.n8120 DVDD.n1855 2.24552
R5661 DVDD.n8116 DVDD.n8115 2.24552
R5662 DVDD.n8120 DVDD.n1854 2.24552
R5663 DVDD.n8115 DVDD.n1890 2.24552
R5664 DVDD.n8292 DVDD.n1666 2.24552
R5665 DVDD.n1689 DVDD.n1678 2.24552
R5666 DVDD.n8292 DVDD.n1667 2.24552
R5667 DVDD.n1691 DVDD.n1678 2.24552
R5668 DVDD.n8292 DVDD.n1668 2.24552
R5669 DVDD.n8292 DVDD.n1670 2.24552
R5670 DVDD.n1694 DVDD.n1678 2.24552
R5671 DVDD.n8292 DVDD.n1671 2.24552
R5672 DVDD.n1696 DVDD.n1678 2.24552
R5673 DVDD.n8292 DVDD.n1674 2.24552
R5674 DVDD.n1698 DVDD.n1678 2.24552
R5675 DVDD.n8292 DVDD.n1675 2.24552
R5676 DVDD.n1700 DVDD.n1678 2.24552
R5677 DVDD.n8292 DVDD.n1676 2.24552
R5678 DVDD.n2317 DVDD.n2292 2.24552
R5679 DVDD.n7749 DVDD.n2286 2.24552
R5680 DVDD.n2319 DVDD.n2292 2.24552
R5681 DVDD.n7749 DVDD.n2283 2.24552
R5682 DVDD.n2321 DVDD.n2292 2.24552
R5683 DVDD.n7749 DVDD.n2282 2.24552
R5684 DVDD.n2324 DVDD.n2292 2.24552
R5685 DVDD.n7749 DVDD.n2287 2.24552
R5686 DVDD.n2326 DVDD.n2292 2.24552
R5687 DVDD.n7749 DVDD.n2288 2.24552
R5688 DVDD.n2328 DVDD.n2292 2.24552
R5689 DVDD.n7749 DVDD.n2281 2.24552
R5690 DVDD.n2330 DVDD.n2292 2.24552
R5691 DVDD.n7749 DVDD.n2280 2.24552
R5692 DVDD.n2149 DVDD.n2148 2.24552
R5693 DVDD.n7842 DVDD.n7839 2.24552
R5694 DVDD.n2149 DVDD.n2147 2.24552
R5695 DVDD.n7842 DVDD.n7840 2.24552
R5696 DVDD.n2149 DVDD.n2146 2.24552
R5697 DVDD.n7842 DVDD.n7841 2.24552
R5698 DVDD.n2149 DVDD.n2145 2.24552
R5699 DVDD.n6674 DVDD.n3306 2.24552
R5700 DVDD.n6676 DVDD.n3223 2.24552
R5701 DVDD.n6674 DVDD.n3304 2.24552
R5702 DVDD.n6676 DVDD.n3222 2.24552
R5703 DVDD.n6674 DVDD.n3301 2.24552
R5704 DVDD.n6676 DVDD.n3221 2.24552
R5705 DVDD.n6062 DVDD.n5927 2.24552
R5706 DVDD.n5996 DVDD.n5917 2.24552
R5707 DVDD.n6062 DVDD.n5926 2.24552
R5708 DVDD.n5998 DVDD.n5917 2.24552
R5709 DVDD.n6062 DVDD.n5925 2.24552
R5710 DVDD.n6000 DVDD.n5917 2.24552
R5711 DVDD.n4285 DVDD.n4284 2.24552
R5712 DVDD.n4282 DVDD.n4281 2.24552
R5713 DVDD.n4285 DVDD.n4280 2.24552
R5714 DVDD.n7842 DVDD.n2144 2.24552
R5715 DVDD.n7749 DVDD.n2279 2.24552
R5716 DVDD.n7749 DVDD.n2278 2.24552
R5717 DVDD.n7749 DVDD.n2277 2.24552
R5718 DVDD.n6111 DVDD.n6108 2.24552
R5719 DVDD.n6113 DVDD.n4316 2.24552
R5720 DVDD.n6111 DVDD.n6110 2.24552
R5721 DVDD.n5891 DVDD.n5888 2.24552
R5722 DVDD.n6095 DVDD.n5895 2.24552
R5723 DVDD.n5891 DVDD.n5889 2.24552
R5724 DVDD.n6095 DVDD.n5894 2.24552
R5725 DVDD.n5891 DVDD.n5890 2.24552
R5726 DVDD.n6095 DVDD.n5893 2.24552
R5727 DVDD.n3184 DVDD.n3183 2.24552
R5728 DVDD.n6704 DVDD.n6701 2.24552
R5729 DVDD.n3184 DVDD.n3182 2.24552
R5730 DVDD.n6704 DVDD.n6702 2.24552
R5731 DVDD.n3184 DVDD.n3181 2.24552
R5732 DVDD.n6704 DVDD.n6703 2.24552
R5733 DVDD.n7799 DVDD.n7797 2.24552
R5734 DVDD.n7806 DVDD.n2188 2.24552
R5735 DVDD.n7799 DVDD.n7796 2.24552
R5736 DVDD.n7806 DVDD.n2189 2.24552
R5737 DVDD.n7800 DVDD.n7799 2.24552
R5738 DVDD.n7806 DVDD.n2190 2.24552
R5739 DVDD.n7799 DVDD.n2192 2.24552
R5740 DVDD.n7806 DVDD.n7805 2.24552
R5741 DVDD.n7780 DVDD.n2218 2.24552
R5742 DVDD.n7776 DVDD.n2250 2.24552
R5743 DVDD.n7780 DVDD.n2219 2.24552
R5744 DVDD.n7776 DVDD.n2249 2.24552
R5745 DVDD.n7780 DVDD.n2220 2.24552
R5746 DVDD.n7780 DVDD.n2215 2.24552
R5747 DVDD.n7776 DVDD.n7774 2.24552
R5748 DVDD.n7780 DVDD.n2214 2.24552
R5749 DVDD.n7776 DVDD.n7775 2.24552
R5750 DVDD.n7780 DVDD.n2213 2.24552
R5751 DVDD.n7780 DVDD.n2222 2.24552
R5752 DVDD.n7776 DVDD.n2248 2.24552
R5753 DVDD.n7780 DVDD.n2223 2.24552
R5754 DVDD.n7776 DVDD.n2247 2.24552
R5755 DVDD.n7780 DVDD.n2224 2.24552
R5756 DVDD.n7780 DVDD.n2211 2.24552
R5757 DVDD.n7776 DVDD.n2225 2.24552
R5758 DVDD.n1628 DVDD.n1621 2.24552
R5759 DVDD.n1619 DVDD.n1618 2.24552
R5760 DVDD.n1628 DVDD.n1622 2.24552
R5761 DVDD.n1619 DVDD.n1617 2.24552
R5762 DVDD.n1628 DVDD.n1623 2.24552
R5763 DVDD.n1628 DVDD.n1624 2.24552
R5764 DVDD.n1619 DVDD.n1616 2.24552
R5765 DVDD.n1628 DVDD.n1625 2.24552
R5766 DVDD.n1619 DVDD.n1615 2.24552
R5767 DVDD.n1628 DVDD.n1626 2.24552
R5768 DVDD.n1619 DVDD.n1614 2.24552
R5769 DVDD.n1628 DVDD.n1627 2.24552
R5770 DVDD.n1619 DVDD.n1613 2.24552
R5771 DVDD.n1628 DVDD.n1612 2.24552
R5772 DVDD.n7360 DVDD.n7344 2.24552
R5773 DVDD.n8634 DVDD.n1312 2.24552
R5774 DVDD.n8629 DVDD.n1320 2.24552
R5775 DVDD.n7345 DVDD.n1508 2.24552
R5776 DVDD.n8638 DVDD.n1308 2.24552
R5777 DVDD.n8633 DVDD.n1316 2.24552
R5778 DVDD.n7344 DVDD.n7341 2.24552
R5779 DVDD.n1312 DVDD.n1310 2.24552
R5780 DVDD.n1320 DVDD.n1318 2.24552
R5781 DVDD.n8374 DVDD.n1505 2.24552
R5782 DVDD.n8376 DVDD.n1510 2.24552
R5783 DVDD.n8378 DVDD.n1503 2.24552
R5784 DVDD.n8356 DVDD.n8349 2.24552
R5785 DVDD.n1545 DVDD.n1529 2.24552
R5786 DVDD.n8356 DVDD.n8350 2.24552
R5787 DVDD.n1547 DVDD.n1529 2.24552
R5788 DVDD.n8356 DVDD.n8351 2.24552
R5789 DVDD.n8356 DVDD.n8352 2.24552
R5790 DVDD.n1551 DVDD.n1529 2.24552
R5791 DVDD.n8356 DVDD.n8353 2.24552
R5792 DVDD.n1553 DVDD.n1529 2.24552
R5793 DVDD.n8356 DVDD.n8354 2.24552
R5794 DVDD.n1557 DVDD.n1529 2.24552
R5795 DVDD.n8356 DVDD.n8355 2.24552
R5796 DVDD.n1559 DVDD.n1529 2.24552
R5797 DVDD.n8356 DVDD.n1528 2.24552
R5798 DVDD.n2389 DVDD.n2372 2.24552
R5799 DVDD.n7660 DVDD.n7657 2.24552
R5800 DVDD.n2391 DVDD.n2372 2.24552
R5801 DVDD.n7660 DVDD.n2457 2.24552
R5802 DVDD.n2393 DVDD.n2372 2.24552
R5803 DVDD.n7660 DVDD.n2456 2.24552
R5804 DVDD.n2396 DVDD.n2372 2.24552
R5805 DVDD.n7660 DVDD.n7658 2.24552
R5806 DVDD.n2398 DVDD.n2372 2.24552
R5807 DVDD.n7660 DVDD.n7659 2.24552
R5808 DVDD.n2400 DVDD.n2372 2.24552
R5809 DVDD.n7660 DVDD.n2455 2.24552
R5810 DVDD.n2402 DVDD.n2372 2.24552
R5811 DVDD.n7660 DVDD.n2373 2.24552
R5812 DVDD.n6979 DVDD.n6933 2.24552
R5813 DVDD.n6985 DVDD.n2639 2.24552
R5814 DVDD.n6979 DVDD.n6978 2.24552
R5815 DVDD.n6985 DVDD.n2640 2.24552
R5816 DVDD.n6980 DVDD.n6979 2.24552
R5817 DVDD.n6985 DVDD.n2641 2.24552
R5818 DVDD.n6979 DVDD.n6977 2.24552
R5819 DVDD.n2725 DVDD.n2656 2.24552
R5820 DVDD.n2724 DVDD.n2657 2.24552
R5821 DVDD.n2728 DVDD.n2656 2.24552
R5822 DVDD.n2727 DVDD.n2657 2.24552
R5823 DVDD.n2731 DVDD.n2656 2.24552
R5824 DVDD.n2730 DVDD.n2657 2.24552
R5825 DVDD.n6892 DVDD.n2743 2.24552
R5826 DVDD.n6891 DVDD.n2777 2.24552
R5827 DVDD.n6889 DVDD.n2743 2.24552
R5828 DVDD.n2784 DVDD.n2777 2.24552
R5829 DVDD.n6876 DVDD.n2743 2.24552
R5830 DVDD.n6874 DVDD.n2777 2.24552
R5831 DVDD.n2877 DVDD.n2804 2.24552
R5832 DVDD.n2876 DVDD.n2805 2.24552
R5833 DVDD.n6854 DVDD.n2804 2.24552
R5834 DVDD.n6985 DVDD.n6984 2.24552
R5835 DVDD.n7660 DVDD.n2454 2.24552
R5836 DVDD.n7660 DVDD.n2453 2.24552
R5837 DVDD.n7660 DVDD.n2452 2.24552
R5838 DVDD.n8369 DVDD.n1519 2.24552
R5839 DVDD.n8365 DVDD.n8362 2.24552
R5840 DVDD.n1521 DVDD.n1512 2.24552
R5841 DVDD.n8365 DVDD.n8363 2.24552
R5842 DVDD.n1523 DVDD.n1512 2.24552
R5843 DVDD.n8365 DVDD.n8364 2.24552
R5844 DVDD.n1525 DVDD.n1512 2.24552
R5845 DVDD.n8366 DVDD.n8365 2.24552
R5846 DVDD.n8367 DVDD.n1512 2.24552
R5847 DVDD.n8365 DVDD.n1511 2.24552
R5848 DVDD.n8284 DVDD.n1702 2.24552
R5849 DVDD.n1713 DVDD.n1703 2.24552
R5850 DVDD.n8284 DVDD.n1722 2.24552
R5851 DVDD.n1715 DVDD.n1703 2.24552
R5852 DVDD.n8284 DVDD.n1721 2.24552
R5853 DVDD.n1717 DVDD.n1703 2.24552
R5854 DVDD.n8284 DVDD.n1720 2.24552
R5855 DVDD.n1719 DVDD.n1703 2.24552
R5856 DVDD.n8285 DVDD.n8284 2.24552
R5857 DVDD.n1706 DVDD.n1703 2.24552
R5858 DVDD.n7503 DVDD.n7067 2.24552
R5859 DVDD.n7077 DVDD.n7068 2.24552
R5860 DVDD.n7503 DVDD.n7089 2.24552
R5861 DVDD.n7079 DVDD.n7068 2.24552
R5862 DVDD.n7503 DVDD.n7088 2.24552
R5863 DVDD.n7081 DVDD.n7068 2.24552
R5864 DVDD.n7503 DVDD.n7087 2.24552
R5865 DVDD.n7083 DVDD.n7068 2.24552
R5866 DVDD.n7503 DVDD.n7086 2.24552
R5867 DVDD.n7085 DVDD.n7068 2.24552
R5868 DVDD.n7430 DVDD.n7338 2.24552
R5869 DVDD.n7425 DVDD.n7422 2.24552
R5870 DVDD.n7430 DVDD.n7337 2.24552
R5871 DVDD.n7425 DVDD.n7423 2.24552
R5872 DVDD.n7430 DVDD.n7336 2.24552
R5873 DVDD.n7425 DVDD.n7424 2.24552
R5874 DVDD.n7430 DVDD.n7335 2.24552
R5875 DVDD.n7426 DVDD.n7425 2.24552
R5876 DVDD.n7430 DVDD.n7334 2.24552
R5877 DVDD.n7425 DVDD.n7340 2.24552
R5878 DVDD.n1757 DVDD.n1756 2.24552
R5879 DVDD.n1763 DVDD.n1759 2.24552
R5880 DVDD.n1757 DVDD.n1755 2.24552
R5881 DVDD.n1763 DVDD.n1760 2.24552
R5882 DVDD.n1757 DVDD.n1754 2.24552
R5883 DVDD.n1763 DVDD.n1761 2.24552
R5884 DVDD.n1757 DVDD.n1753 2.24552
R5885 DVDD.n1763 DVDD.n1751 2.24552
R5886 DVDD.n1757 DVDD.n1752 2.24552
R5887 DVDD.n1763 DVDD.n1762 2.24552
R5888 DVDD.n6420 DVDD.n1055 2.24552
R5889 DVDD.n1071 DVDD.n1056 2.24552
R5890 DVDD.n6420 DVDD.n6410 2.24552
R5891 DVDD.n1073 DVDD.n1056 2.24552
R5892 DVDD.n6420 DVDD.n6411 2.24552
R5893 DVDD.n1075 DVDD.n1056 2.24552
R5894 DVDD.n6420 DVDD.n6412 2.24552
R5895 DVDD.n1077 DVDD.n1056 2.24552
R5896 DVDD.n6420 DVDD.n6413 2.24552
R5897 DVDD.n1079 DVDD.n1056 2.24552
R5898 DVDD.n6420 DVDD.n6414 2.24552
R5899 DVDD.n1081 DVDD.n1056 2.24552
R5900 DVDD.n6420 DVDD.n6415 2.24552
R5901 DVDD.n1083 DVDD.n1056 2.24552
R5902 DVDD.n6420 DVDD.n6416 2.24552
R5903 DVDD.n1085 DVDD.n1056 2.24552
R5904 DVDD.n6420 DVDD.n6417 2.24552
R5905 DVDD.n1087 DVDD.n1056 2.24552
R5906 DVDD.n6420 DVDD.n6418 2.24552
R5907 DVDD.n1089 DVDD.n1056 2.24552
R5908 DVDD.n6420 DVDD.n6419 2.24552
R5909 DVDD.n1091 DVDD.n1056 2.24552
R5910 DVDD.n6420 DVDD.n1093 2.24552
R5911 DVDD.n1116 DVDD.n1094 2.24552
R5912 DVDD.n1103 DVDD.n1095 2.24552
R5913 DVDD.n1116 DVDD.n1115 2.24552
R5914 DVDD.n1105 DVDD.n1095 2.24552
R5915 DVDD.n1116 DVDD.n1114 2.24552
R5916 DVDD.n1107 DVDD.n1095 2.24552
R5917 DVDD.n1116 DVDD.n1113 2.24552
R5918 DVDD.n1109 DVDD.n1095 2.24552
R5919 DVDD.n1116 DVDD.n1112 2.24552
R5920 DVDD.n1111 DVDD.n1095 2.24552
R5921 DVDD.n6626 DVDD.n1117 2.24552
R5922 DVDD.n1133 DVDD.n1118 2.24552
R5923 DVDD.n6626 DVDD.n6616 2.24552
R5924 DVDD.n1135 DVDD.n1118 2.24552
R5925 DVDD.n6626 DVDD.n6617 2.24552
R5926 DVDD.n1137 DVDD.n1118 2.24552
R5927 DVDD.n6626 DVDD.n6618 2.24552
R5928 DVDD.n1139 DVDD.n1118 2.24552
R5929 DVDD.n6626 DVDD.n6619 2.24552
R5930 DVDD.n1141 DVDD.n1118 2.24552
R5931 DVDD.n6626 DVDD.n6620 2.24552
R5932 DVDD.n1143 DVDD.n1118 2.24552
R5933 DVDD.n6626 DVDD.n6621 2.24552
R5934 DVDD.n1145 DVDD.n1118 2.24552
R5935 DVDD.n6626 DVDD.n6622 2.24552
R5936 DVDD.n1147 DVDD.n1118 2.24552
R5937 DVDD.n6626 DVDD.n6623 2.24552
R5938 DVDD.n1149 DVDD.n1118 2.24552
R5939 DVDD.n6626 DVDD.n6624 2.24552
R5940 DVDD.n1151 DVDD.n1118 2.24552
R5941 DVDD.n6626 DVDD.n6625 2.24552
R5942 DVDD.n1153 DVDD.n1118 2.24552
R5943 DVDD.n6626 DVDD.n1155 2.24552
R5944 DVDD.n7926 DVDD.n1156 2.24552
R5945 DVDD.n1172 DVDD.n1157 2.24552
R5946 DVDD.n7926 DVDD.n7916 2.24552
R5947 DVDD.n1174 DVDD.n1157 2.24552
R5948 DVDD.n7926 DVDD.n7917 2.24552
R5949 DVDD.n1176 DVDD.n1157 2.24552
R5950 DVDD.n7926 DVDD.n7918 2.24552
R5951 DVDD.n1178 DVDD.n1157 2.24552
R5952 DVDD.n7926 DVDD.n7919 2.24552
R5953 DVDD.n1180 DVDD.n1157 2.24552
R5954 DVDD.n7926 DVDD.n7920 2.24552
R5955 DVDD.n1182 DVDD.n1157 2.24552
R5956 DVDD.n7926 DVDD.n7921 2.24552
R5957 DVDD.n1184 DVDD.n1157 2.24552
R5958 DVDD.n7926 DVDD.n7922 2.24552
R5959 DVDD.n1186 DVDD.n1157 2.24552
R5960 DVDD.n7926 DVDD.n7923 2.24552
R5961 DVDD.n1188 DVDD.n1157 2.24552
R5962 DVDD.n7926 DVDD.n7924 2.24552
R5963 DVDD.n1190 DVDD.n1157 2.24552
R5964 DVDD.n7926 DVDD.n7925 2.24552
R5965 DVDD.n1192 DVDD.n1157 2.24552
R5966 DVDD.n7926 DVDD.n1194 2.24552
R5967 DVDD.n8031 DVDD.n1195 2.24552
R5968 DVDD.n1211 DVDD.n1196 2.24552
R5969 DVDD.n8031 DVDD.n8021 2.24552
R5970 DVDD.n1213 DVDD.n1196 2.24552
R5971 DVDD.n8031 DVDD.n8022 2.24552
R5972 DVDD.n1215 DVDD.n1196 2.24552
R5973 DVDD.n8031 DVDD.n8023 2.24552
R5974 DVDD.n1217 DVDD.n1196 2.24552
R5975 DVDD.n8031 DVDD.n8024 2.24552
R5976 DVDD.n1219 DVDD.n1196 2.24552
R5977 DVDD.n8031 DVDD.n8025 2.24552
R5978 DVDD.n1221 DVDD.n1196 2.24552
R5979 DVDD.n8031 DVDD.n8026 2.24552
R5980 DVDD.n1223 DVDD.n1196 2.24552
R5981 DVDD.n8031 DVDD.n8027 2.24552
R5982 DVDD.n1225 DVDD.n1196 2.24552
R5983 DVDD.n8031 DVDD.n8028 2.24552
R5984 DVDD.n1227 DVDD.n1196 2.24552
R5985 DVDD.n8031 DVDD.n8029 2.24552
R5986 DVDD.n1229 DVDD.n1196 2.24552
R5987 DVDD.n8031 DVDD.n8030 2.24552
R5988 DVDD.n1231 DVDD.n1196 2.24552
R5989 DVDD.n8031 DVDD.n1233 2.24552
R5990 DVDD.n8151 DVDD.n1234 2.24552
R5991 DVDD.n1250 DVDD.n1235 2.24552
R5992 DVDD.n8151 DVDD.n8143 2.24552
R5993 DVDD.n1252 DVDD.n1235 2.24552
R5994 DVDD.n8151 DVDD.n8144 2.24552
R5995 DVDD.n1254 DVDD.n1235 2.24552
R5996 DVDD.n8151 DVDD.n8145 2.24552
R5997 DVDD.n1256 DVDD.n1235 2.24552
R5998 DVDD.n8151 DVDD.n8146 2.24552
R5999 DVDD.n1258 DVDD.n1235 2.24552
R6000 DVDD.n8151 DVDD.n8147 2.24552
R6001 DVDD.n1260 DVDD.n1235 2.24552
R6002 DVDD.n8151 DVDD.n8148 2.24552
R6003 DVDD.n1262 DVDD.n1235 2.24552
R6004 DVDD.n8151 DVDD.n8149 2.24552
R6005 DVDD.n1266 DVDD.n1235 2.24552
R6006 DVDD.n8151 DVDD.n8150 2.24552
R6007 DVDD.n1268 DVDD.n1235 2.24552
R6008 DVDD.n8151 DVDD.n1270 2.24552
R6009 DVDD.n1294 DVDD.n1271 2.24552
R6010 DVDD.n1281 DVDD.n1272 2.24552
R6011 DVDD.n1294 DVDD.n1293 2.24552
R6012 DVDD.n1283 DVDD.n1272 2.24552
R6013 DVDD.n1294 DVDD.n1292 2.24552
R6014 DVDD.n1285 DVDD.n1272 2.24552
R6015 DVDD.n1294 DVDD.n1291 2.24552
R6016 DVDD.n1287 DVDD.n1272 2.24552
R6017 DVDD.n1294 DVDD.n1290 2.24552
R6018 DVDD.n1289 DVDD.n1272 2.24552
R6019 DVDD.n8643 DVDD.n1296 2.24552
R6020 DVDD.n618 DVDD.n606 2.24552
R6021 DVDD.n620 DVDD.n611 2.24552
R6022 DVDD.n8910 DVDD.n632 2.24552
R6023 DVDD.n622 DVDD.n611 2.24552
R6024 DVDD.n8910 DVDD.n631 2.24552
R6025 DVDD.n624 DVDD.n611 2.24552
R6026 DVDD.n8910 DVDD.n630 2.24552
R6027 DVDD.n626 DVDD.n611 2.24552
R6028 DVDD.n8910 DVDD.n629 2.24552
R6029 DVDD.n628 DVDD.n611 2.24552
R6030 DVDD.n4738 DVDD.n4599 2.24552
R6031 DVDD.n4821 DVDD.n4598 2.24552
R6032 DVDD.n4738 DVDD.n4736 2.24552
R6033 DVDD.n4821 DVDD.n4597 2.24552
R6034 DVDD.n4738 DVDD.n4735 2.24552
R6035 DVDD.n4821 DVDD.n4596 2.24552
R6036 DVDD.n4738 DVDD.n4734 2.24552
R6037 DVDD.n4821 DVDD.n4595 2.24552
R6038 DVDD.n4738 DVDD.n4733 2.24552
R6039 DVDD.n4821 DVDD.n4594 2.24552
R6040 DVDD.n5400 DVDD.n2960 2.24552
R6041 DVDD.n2976 DVDD.n2961 2.24552
R6042 DVDD.n5400 DVDD.n5390 2.24552
R6043 DVDD.n2978 DVDD.n2961 2.24552
R6044 DVDD.n5400 DVDD.n5391 2.24552
R6045 DVDD.n2980 DVDD.n2961 2.24552
R6046 DVDD.n5400 DVDD.n5392 2.24552
R6047 DVDD.n2982 DVDD.n2961 2.24552
R6048 DVDD.n5400 DVDD.n5393 2.24552
R6049 DVDD.n2984 DVDD.n2961 2.24552
R6050 DVDD.n5400 DVDD.n5394 2.24552
R6051 DVDD.n2986 DVDD.n2961 2.24552
R6052 DVDD.n5400 DVDD.n5395 2.24552
R6053 DVDD.n2988 DVDD.n2961 2.24552
R6054 DVDD.n5400 DVDD.n5396 2.24552
R6055 DVDD.n2990 DVDD.n2961 2.24552
R6056 DVDD.n5400 DVDD.n5397 2.24552
R6057 DVDD.n2992 DVDD.n2961 2.24552
R6058 DVDD.n5400 DVDD.n5398 2.24552
R6059 DVDD.n2994 DVDD.n2961 2.24552
R6060 DVDD.n5400 DVDD.n5399 2.24552
R6061 DVDD.n2996 DVDD.n2961 2.24552
R6062 DVDD.n5400 DVDD.n2998 2.24552
R6063 DVDD.n3022 DVDD.n2999 2.24552
R6064 DVDD.n3009 DVDD.n3000 2.24552
R6065 DVDD.n3022 DVDD.n3021 2.24552
R6066 DVDD.n3011 DVDD.n3000 2.24552
R6067 DVDD.n3022 DVDD.n3020 2.24552
R6068 DVDD.n3013 DVDD.n3000 2.24552
R6069 DVDD.n3022 DVDD.n3019 2.24552
R6070 DVDD.n3015 DVDD.n3000 2.24552
R6071 DVDD.n3022 DVDD.n3018 2.24552
R6072 DVDD.n3017 DVDD.n3000 2.24552
R6073 DVDD.n6765 DVDD.n3023 2.24552
R6074 DVDD.n3039 DVDD.n3024 2.24552
R6075 DVDD.n6765 DVDD.n6755 2.24552
R6076 DVDD.n3041 DVDD.n3024 2.24552
R6077 DVDD.n6765 DVDD.n6756 2.24552
R6078 DVDD.n3043 DVDD.n3024 2.24552
R6079 DVDD.n6765 DVDD.n6757 2.24552
R6080 DVDD.n3045 DVDD.n3024 2.24552
R6081 DVDD.n6765 DVDD.n6758 2.24552
R6082 DVDD.n3047 DVDD.n3024 2.24552
R6083 DVDD.n6765 DVDD.n6759 2.24552
R6084 DVDD.n3049 DVDD.n3024 2.24552
R6085 DVDD.n6765 DVDD.n6760 2.24552
R6086 DVDD.n3051 DVDD.n3024 2.24552
R6087 DVDD.n6765 DVDD.n6761 2.24552
R6088 DVDD.n3053 DVDD.n3024 2.24552
R6089 DVDD.n6765 DVDD.n6762 2.24552
R6090 DVDD.n3055 DVDD.n3024 2.24552
R6091 DVDD.n6765 DVDD.n6763 2.24552
R6092 DVDD.n3057 DVDD.n3024 2.24552
R6093 DVDD.n6765 DVDD.n6764 2.24552
R6094 DVDD.n3059 DVDD.n3024 2.24552
R6095 DVDD.n6766 DVDD.n6765 2.24552
R6096 DVDD.n2609 DVDD.n2598 2.24552
R6097 DVDD.n2597 DVDD.n2596 2.24552
R6098 DVDD.n2609 DVDD.n2599 2.24552
R6099 DVDD.n2597 DVDD.n2595 2.24552
R6100 DVDD.n2609 DVDD.n2600 2.24552
R6101 DVDD.n2597 DVDD.n2594 2.24552
R6102 DVDD.n2609 DVDD.n2601 2.24552
R6103 DVDD.n2597 DVDD.n2593 2.24552
R6104 DVDD.n2609 DVDD.n2602 2.24552
R6105 DVDD.n2597 DVDD.n2592 2.24552
R6106 DVDD.n2609 DVDD.n2603 2.24552
R6107 DVDD.n2597 DVDD.n2591 2.24552
R6108 DVDD.n2609 DVDD.n2604 2.24552
R6109 DVDD.n2597 DVDD.n2590 2.24552
R6110 DVDD.n2609 DVDD.n2605 2.24552
R6111 DVDD.n2597 DVDD.n2589 2.24552
R6112 DVDD.n2609 DVDD.n2606 2.24552
R6113 DVDD.n2597 DVDD.n2588 2.24552
R6114 DVDD.n2609 DVDD.n2607 2.24552
R6115 DVDD.n2597 DVDD.n2587 2.24552
R6116 DVDD.n2609 DVDD.n2608 2.24552
R6117 DVDD.n2597 DVDD.n2586 2.24552
R6118 DVDD.n2609 DVDD.n2585 2.24552
R6119 DVDD.n7587 DVDD.n7577 2.24552
R6120 DVDD.n7592 DVDD.n2485 2.24552
R6121 DVDD.n7587 DVDD.n7578 2.24552
R6122 DVDD.n7592 DVDD.n2484 2.24552
R6123 DVDD.n7587 DVDD.n7579 2.24552
R6124 DVDD.n7592 DVDD.n2483 2.24552
R6125 DVDD.n7587 DVDD.n7580 2.24552
R6126 DVDD.n7592 DVDD.n2482 2.24552
R6127 DVDD.n7587 DVDD.n7581 2.24552
R6128 DVDD.n7592 DVDD.n2481 2.24552
R6129 DVDD.n7587 DVDD.n7582 2.24552
R6130 DVDD.n7592 DVDD.n2480 2.24552
R6131 DVDD.n7587 DVDD.n7583 2.24552
R6132 DVDD.n7592 DVDD.n2479 2.24552
R6133 DVDD.n7587 DVDD.n7584 2.24552
R6134 DVDD.n7592 DVDD.n2478 2.24552
R6135 DVDD.n7587 DVDD.n7585 2.24552
R6136 DVDD.n7592 DVDD.n2477 2.24552
R6137 DVDD.n7587 DVDD.n7586 2.24552
R6138 DVDD.n7592 DVDD.n2476 2.24552
R6139 DVDD.n7588 DVDD.n7587 2.24552
R6140 DVDD.n7592 DVDD.n2475 2.24552
R6141 DVDD.n7587 DVDD.n2487 2.24552
R6142 DVDD.n7281 DVDD.n7273 2.24552
R6143 DVDD.n7121 DVDD.n7106 2.24552
R6144 DVDD.n7281 DVDD.n7274 2.24552
R6145 DVDD.n7123 DVDD.n7106 2.24552
R6146 DVDD.n7281 DVDD.n7275 2.24552
R6147 DVDD.n7125 DVDD.n7106 2.24552
R6148 DVDD.n7281 DVDD.n7276 2.24552
R6149 DVDD.n7127 DVDD.n7106 2.24552
R6150 DVDD.n7281 DVDD.n7277 2.24552
R6151 DVDD.n7129 DVDD.n7106 2.24552
R6152 DVDD.n7281 DVDD.n7278 2.24552
R6153 DVDD.n7131 DVDD.n7106 2.24552
R6154 DVDD.n7281 DVDD.n7279 2.24552
R6155 DVDD.n7133 DVDD.n7106 2.24552
R6156 DVDD.n7281 DVDD.n7280 2.24552
R6157 DVDD.n7203 DVDD.n7106 2.24552
R6158 DVDD.n7282 DVDD.n7281 2.24552
R6159 DVDD.n7283 DVDD.n7106 2.24552
R6160 DVDD.n7281 DVDD.n7105 2.24552
R6161 DVDD.n7298 DVDD.n7297 2.24552
R6162 DVDD.n7304 DVDD.n7300 2.24552
R6163 DVDD.n7298 DVDD.n7296 2.24552
R6164 DVDD.n7304 DVDD.n7301 2.24552
R6165 DVDD.n7298 DVDD.n7295 2.24552
R6166 DVDD.n7304 DVDD.n7302 2.24552
R6167 DVDD.n7298 DVDD.n7294 2.24552
R6168 DVDD.n7304 DVDD.n7303 2.24552
R6169 DVDD.n7298 DVDD.n7293 2.24552
R6170 DVDD.n7304 DVDD.n7292 2.24552
R6171 DVDD.n8379 DVDD.n1498 2.24552
R6172 DVDD.n4787 DVDD.n4739 2.24552
R6173 DVDD.n4779 DVDD.n4740 2.24552
R6174 DVDD.n4816 DVDD.n4746 2.24552
R6175 DVDD.n4781 DVDD.n4740 2.24552
R6176 DVDD.n4816 DVDD.n4745 2.24552
R6177 DVDD.n4783 DVDD.n4740 2.24552
R6178 DVDD.n4816 DVDD.n4744 2.24552
R6179 DVDD.n4785 DVDD.n4740 2.24552
R6180 DVDD.n4816 DVDD.n4743 2.24552
R6181 DVDD.n4774 DVDD.n4740 2.24552
R6182 DVDD.n31 DVDD.n24 2.24552
R6183 DVDD.n33 DVDD.n20 2.24552
R6184 DVDD.n34 DVDD.n24 2.24552
R6185 DVDD.n36 DVDD.n20 2.24552
R6186 DVDD.n37 DVDD.n24 2.24552
R6187 DVDD.n39 DVDD.n20 2.24552
R6188 DVDD.n40 DVDD.n24 2.24552
R6189 DVDD.n42 DVDD.n20 2.24552
R6190 DVDD.n43 DVDD.n24 2.24552
R6191 DVDD.n45 DVDD.n20 2.24552
R6192 DVDD.n8210 DVDD.n1789 2.24518
R6193 DVDD.n8205 DVDD.n8199 2.24518
R6194 DVDD.n8210 DVDD.n1788 2.24518
R6195 DVDD.n8205 DVDD.n8198 2.24518
R6196 DVDD.n8210 DVDD.n1787 2.24518
R6197 DVDD.n8205 DVDD.n8197 2.24518
R6198 DVDD.n8210 DVDD.n1786 2.24518
R6199 DVDD.n8206 DVDD.n8205 2.24518
R6200 DVDD.n8210 DVDD.n1785 2.24518
R6201 DVDD.n8205 DVDD.n1791 2.24518
R6202 DVDD.n8187 DVDD.n8177 2.24518
R6203 DVDD.n1815 DVDD.n1799 2.24518
R6204 DVDD.n8187 DVDD.n8178 2.24518
R6205 DVDD.n1817 DVDD.n1799 2.24518
R6206 DVDD.n8187 DVDD.n8179 2.24518
R6207 DVDD.n1819 DVDD.n1799 2.24518
R6208 DVDD.n8187 DVDD.n8180 2.24518
R6209 DVDD.n1821 DVDD.n1799 2.24518
R6210 DVDD.n8187 DVDD.n8181 2.24518
R6211 DVDD.n1823 DVDD.n1799 2.24518
R6212 DVDD.n8187 DVDD.n8182 2.24518
R6213 DVDD.n1825 DVDD.n1799 2.24518
R6214 DVDD.n8187 DVDD.n8183 2.24518
R6215 DVDD.n1827 DVDD.n1799 2.24518
R6216 DVDD.n8187 DVDD.n8184 2.24518
R6217 DVDD.n1829 DVDD.n1799 2.24518
R6218 DVDD.n8187 DVDD.n8185 2.24518
R6219 DVDD.n1831 DVDD.n1799 2.24518
R6220 DVDD.n8187 DVDD.n8186 2.24518
R6221 DVDD.n1833 DVDD.n1799 2.24518
R6222 DVDD.n8188 DVDD.n8187 2.24518
R6223 DVDD.n8189 DVDD.n1799 2.24518
R6224 DVDD.n8187 DVDD.n1798 2.24518
R6225 DVDD.n7997 DVDD.n7986 2.24518
R6226 DVDD.n7985 DVDD.n7984 2.24518
R6227 DVDD.n7997 DVDD.n7987 2.24518
R6228 DVDD.n7985 DVDD.n7983 2.24518
R6229 DVDD.n7997 DVDD.n7988 2.24518
R6230 DVDD.n7985 DVDD.n7982 2.24518
R6231 DVDD.n7997 DVDD.n7989 2.24518
R6232 DVDD.n7985 DVDD.n7981 2.24518
R6233 DVDD.n7997 DVDD.n7990 2.24518
R6234 DVDD.n7985 DVDD.n7980 2.24518
R6235 DVDD.n7997 DVDD.n7991 2.24518
R6236 DVDD.n7985 DVDD.n7979 2.24518
R6237 DVDD.n7997 DVDD.n7992 2.24518
R6238 DVDD.n7985 DVDD.n7978 2.24518
R6239 DVDD.n7997 DVDD.n7993 2.24518
R6240 DVDD.n7985 DVDD.n7977 2.24518
R6241 DVDD.n7997 DVDD.n7994 2.24518
R6242 DVDD.n7985 DVDD.n7976 2.24518
R6243 DVDD.n7997 DVDD.n7995 2.24518
R6244 DVDD.n7985 DVDD.n7975 2.24518
R6245 DVDD.n7997 DVDD.n7996 2.24518
R6246 DVDD.n7985 DVDD.n7974 2.24518
R6247 DVDD.n7997 DVDD.n7973 2.24518
R6248 DVDD.n2051 DVDD.n2029 2.24518
R6249 DVDD.n7954 DVDD.n7952 2.24518
R6250 DVDD.n2053 DVDD.n2028 2.24518
R6251 DVDD.n7954 DVDD.n7953 2.24518
R6252 DVDD.n2055 DVDD.n2028 2.24518
R6253 DVDD.n7955 DVDD.n7954 2.24518
R6254 DVDD.n7956 DVDD.n2028 2.24518
R6255 DVDD.n7954 DVDD.n2027 2.24518
R6256 DVDD.n6481 DVDD.n6480 2.24518
R6257 DVDD.n6485 DVDD.n6482 2.24518
R6258 DVDD.n6481 DVDD.n6479 2.24518
R6259 DVDD.n6485 DVDD.n6483 2.24518
R6260 DVDD.n6481 DVDD.n6478 2.24518
R6261 DVDD.n6485 DVDD.n6484 2.24518
R6262 DVDD.n3477 DVDD.n3467 2.24518
R6263 DVDD.n3476 DVDD.n3420 2.24518
R6264 DVDD.n3480 DVDD.n3467 2.24518
R6265 DVDD.n3479 DVDD.n3420 2.24518
R6266 DVDD.n6462 DVDD.n3467 2.24518
R6267 DVDD.n3482 DVDD.n3420 2.24518
R6268 DVDD.n3549 DVDD.n3547 2.24518
R6269 DVDD.n3551 DVDD.n3550 2.24518
R6270 DVDD.n3549 DVDD.n3548 2.24518
R6271 DVDD.n7149 DVDD.n7144 2.24505
R6272 DVDD.n7150 DVDD.n7149 2.24505
R6273 DVDD.n7155 DVDD.n7152 2.24505
R6274 DVDD.n7161 DVDD.n7158 2.24505
R6275 DVDD.n7147 DVDD.n7145 2.24505
R6276 DVDD.n7178 DVDD.n7153 2.24505
R6277 DVDD.n7179 DVDD.n7178 2.24505
R6278 DVDD.n7173 DVDD.n7159 2.24505
R6279 DVDD.n7174 DVDD.n7173 2.24505
R6280 DVDD.n7359 DVDD.n7343 2.24505
R6281 DVDD.n1314 DVDD.n1307 2.24505
R6282 DVDD.n8628 DVDD.n1315 2.24505
R6283 DVDD.n1509 DVDD.n1504 2.24505
R6284 DVDD.n8373 DVDD.n8372 2.24505
R6285 DVDD.n8375 DVDD.n8371 2.24505
R6286 DVDD.n7141 DVDD.n7138 2.24505
R6287 DVDD.n7187 DVDD.n7139 2.24505
R6288 DVDD.n7188 DVDD.n7187 2.24505
R6289 DVDD.n1302 DVDD.n1301 2.24505
R6290 DVDD.n1298 DVDD.n1297 2.24505
R6291 DVDD.n7169 DVDD.n7164 2.24505
R6292 DVDD.n7166 DVDD.n7163 2.24505
R6293 DVDD.n1300 DVDD.n1297 2.24505
R6294 DVDD.n7167 DVDD.n7166 2.24505
R6295 DVDD.n8386 DVDD.n1499 2.24505
R6296 DVDD.n8384 DVDD.n8382 2.24505
R6297 DVDD.n8382 DVDD.n8381 2.24505
R6298 DVDD.n7201 DVDD.n7193 2.24505
R6299 DVDD.n7199 DVDD.n7197 2.24505
R6300 DVDD.n7197 DVDD.n7196 2.24505
R6301 DVDD.n8437 DVDD.n1328 2.24456
R6302 DVDD.n8496 DVDD.n8495 2.24456
R6303 DVDD.n8600 DVDD.n1356 2.24456
R6304 DVDD.n8432 DVDD.n1334 2.24456
R6305 DVDD.n8500 DVDD.n8499 2.24456
R6306 DVDD.n8595 DVDD.n1365 2.24456
R6307 DVDD.n8427 DVDD.n8422 2.24456
R6308 DVDD.n8506 DVDD.n8505 2.24456
R6309 DVDD.n8512 DVDD.n8511 2.24456
R6310 DVDD.n8419 DVDD.n1464 2.24456
R6311 DVDD.n1488 DVDD.n1469 2.24456
R6312 DVDD.n1483 DVDD.n1475 2.24456
R6313 DVDD.n1446 DVDD.n1432 2.24456
R6314 DVDD.n1436 DVDD.n1354 2.24456
R6315 DVDD.n8598 DVDD.n1352 2.24456
R6316 DVDD.n1451 DVDD.n1424 2.24456
R6317 DVDD.n1428 DVDD.n1363 2.24456
R6318 DVDD.n8593 DVDD.n1361 2.24456
R6319 DVDD.n1456 DVDD.n1418 2.24456
R6320 DVDD.n8508 DVDD.n1413 2.24456
R6321 DVDD.n8514 DVDD.n1407 2.24456
R6322 DVDD.n8417 DVDD.n1460 2.24456
R6323 DVDD.n1486 DVDD.n1484 2.24456
R6324 DVDD.n1481 DVDD.n1480 2.24456
R6325 DVDD.n7745 DVDD.n7744 2.24442
R6326 DVDD.n7745 DVDD.n2333 2.24442
R6327 DVDD.n7733 DVDD.n2337 2.24442
R6328 DVDD.n7742 DVDD.n7741 2.24442
R6329 DVDD.n7735 DVDD.n2339 2.24442
R6330 DVDD.n7722 DVDD.n7704 2.24442
R6331 DVDD.n7722 DVDD.n7721 2.24442
R6332 DVDD.n7716 DVDD.n7711 2.24442
R6333 DVDD.n7717 DVDD.n7716 2.24442
R6334 DVDD.n7707 DVDD.n7703 2.24442
R6335 DVDD.n7709 DVDD.n7703 2.24442
R6336 DVDD.n7715 DVDD.n7710 2.24442
R6337 DVDD.n7712 DVDD.n7710 2.24442
R6338 DVDD.n7699 DVDD.n2345 2.24442
R6339 DVDD.n7698 DVDD.n7697 2.24442
R6340 DVDD.n7697 DVDD.n2344 2.24442
R6341 DVDD.n7701 DVDD.n2347 2.24442
R6342 DVDD.n2367 DVDD.n2360 2.24442
R6343 DVDD.n2369 DVDD.n2362 2.24442
R6344 DVDD.n7688 DVDD.n2350 2.24442
R6345 DVDD.n7692 DVDD.n2350 2.24442
R6346 DVDD.n7691 DVDD.n7690 2.24442
R6347 DVDD.n7690 DVDD.n2349 2.24442
R6348 DVDD.n7683 DVDD.n2354 2.24442
R6349 DVDD.n7685 DVDD.n2357 2.24442
R6350 DVDD.n8537 DVDD.n8522 2.24011
R6351 DVDD.n8625 DVDD.n1327 2.24011
R6352 DVDD.n8540 DVDD.n8519 2.24011
R6353 DVDD.n8622 DVDD.n1333 2.24011
R6354 DVDD.n8544 DVDD.n1404 2.24011
R6355 DVDD.n7356 DVDD.n1458 2.24011
R6356 DVDD.n8547 DVDD.n1398 2.24011
R6357 DVDD.n7348 DVDD.n1462 2.24011
R6358 DVDD.n8536 DVDD.n1360 2.24011
R6359 DVDD.n8627 DVDD.n1323 2.24011
R6360 DVDD.n8517 DVDD.n1369 2.24011
R6361 DVDD.n8620 DVDD.n1330 2.24011
R6362 DVDD.n8516 DVDD.n1402 2.24011
R6363 DVDD.n7358 DVDD.n7354 2.24011
R6364 DVDD.n1401 DVDD.n1396 2.24011
R6365 DVDD.n7347 DVDD.n1506 2.24011
R6366 DVDD.n1880 DVDD.n1677 2.23892
R6367 DVDD.n1881 DVDD.n1679 2.23892
R6368 DVDD.n1877 DVDD.n1679 2.23892
R6369 DVDD.n7670 DVDD.n2291 2.23892
R6370 DVDD.n7668 DVDD.n2291 2.23892
R6371 DVDD.n7667 DVDD.n2293 2.23892
R6372 DVDD.n7669 DVDD.n2293 2.23892
R6373 DVDD.n2436 DVDD.n2430 2.23892
R6374 DVDD.n2437 DVDD.n2436 2.23892
R6375 DVDD.n2439 DVDD.n2431 2.23892
R6376 DVDD.n2439 DVDD.n2438 2.23892
R6377 DVDD.n2413 DVDD.n2407 2.23892
R6378 DVDD.n2414 DVDD.n2413 2.23892
R6379 DVDD.n2416 DVDD.n2408 2.23892
R6380 DVDD.n2416 DVDD.n2415 2.23892
R6381 DVDD.n1874 DVDD.n1873 2.23892
R6382 DVDD.n1874 DVDD.n1868 2.23892
R6383 DVDD.n1871 DVDD.n1867 2.23892
R6384 DVDD.n1871 DVDD.n1869 2.23892
R6385 DVDD.n7674 DVDD.n7673 2.23892
R6386 DVDD.n7673 DVDD.n7662 2.23892
R6387 DVDD.n7663 DVDD.n2246 2.23892
R6388 DVDD.n7661 DVDD.n2246 2.23892
R6389 DVDD.n2442 DVDD.n2428 2.23892
R6390 DVDD.n2443 DVDD.n2442 2.23892
R6391 DVDD.n2445 DVDD.n2429 2.23892
R6392 DVDD.n2445 DVDD.n2444 2.23892
R6393 DVDD.n2419 DVDD.n2405 2.23892
R6394 DVDD.n2420 DVDD.n2419 2.23892
R6395 DVDD.n2422 DVDD.n2406 2.23892
R6396 DVDD.n2422 DVDD.n2421 2.23892
R6397 DVDD.n4880 DVDD.t10 1.70818
R6398 DVDD.n4951 DVDD.t15 1.70818
R6399 DVDD.n4901 DVDD.t39 1.70818
R6400 DVDD.n9476 DVDD.t2 1.70818
R6401 DVDD.n9512 DVDD.t17 1.70818
R6402 DVDD.n4373 DVDD.t8 1.70818
R6403 DVDD.n5821 DVDD.t21 1.70818
R6404 DVDD.n5840 DVDD.t36 1.70818
R6405 DVDD.n3141 DVDD.t13 1.70818
R6406 DVDD.n9016 DVDD.t26 1.70818
R6407 DVDD.n9072 DVDD.t29 1.70818
R6408 DVDD.n9108 DVDD.t23 1.70818
R6409 DVDD.n4116 DVDD.t24 1.70818
R6410 DVDD.n4221 DVDD.t34 1.70818
R6411 DVDD.n4277 DVDD.t27 1.70818
R6412 DVDD.n6054 DVDD.t3 1.70818
R6413 DVDD.n5942 DVDD.t22 1.70818
R6414 DVDD.n3250 DVDD.t30 1.70818
R6415 DVDD.n9407 DVDD.n9406 1.52335
R6416 DVDD.n8709 DVDD.n8708 1.52335
R6417 DVDD.n8692 DVDD.n8691 1.52209
R6418 DVDD.n6244 DVDD.n6243 1.52209
R6419 DVDD.n6899 DVDD.n6898 1.52209
R6420 DVDD.n5277 DVDD.n4514 1.52209
R6421 DVDD.n439 DVDD.n438 1.52209
R6422 DVDD.n99 DVDD.n96 1.52209
R6423 DVDD.n9602 DVDD.n9601 1.52155
R6424 DVDD.n8675 DVDD.n1046 1.52029
R6425 DVDD.n8747 DVDD.n875 1.52029
R6426 DVDD.n6326 DVDD.n3865 1.52029
R6427 DVDD.n6868 DVDD.n6867 1.52029
R6428 DVDD.n181 DVDD.n155 1.52029
R6429 DVDD.n6779 DVDD.n2916 1.52029
R6430 DVDD.n863 DVDD.n862 1.52029
R6431 DVDD.n1043 DVDD.n217 1.5005
R6432 DVDD.n1008 DVDD.n214 1.5005
R6433 DVDD.n8690 DVDD.n8689 1.5005
R6434 DVDD.n8696 DVDD.n8695 1.5005
R6435 DVDD.n1007 DVDD.n1005 1.5005
R6436 DVDD.n8679 DVDD.n8678 1.5005
R6437 DVDD.n1047 DVDD.n1045 1.5005
R6438 DVDD.n8674 DVDD.n8673 1.5005
R6439 DVDD.n6306 DVDD.n6237 1.5005
R6440 DVDD.n6307 DVDD.n6236 1.5005
R6441 DVDD.n6235 DVDD.n3880 1.5005
R6442 DVDD.n3881 DVDD.n3872 1.5005
R6443 DVDD.n6317 DVDD.n3871 1.5005
R6444 DVDD.n6318 DVDD.n3870 1.5005
R6445 DVDD.n6242 DVDD.n6238 1.5005
R6446 DVDD.n3873 DVDD.n3872 1.5005
R6447 DVDD.n6317 DVDD.n6316 1.5005
R6448 DVDD.n6319 DVDD.n6318 1.5005
R6449 DVDD.n3869 DVDD.n3866 1.5005
R6450 DVDD.n3880 DVDD.n3878 1.5005
R6451 DVDD.n6308 DVDD.n6307 1.5005
R6452 DVDD.n6306 DVDD.n6305 1.5005
R6453 DVDD.n2779 DVDD.n2778 1.5005
R6454 DVDD.n6880 DVDD.n6879 1.5005
R6455 DVDD.n2791 DVDD.n2790 1.5005
R6456 DVDD.n6871 DVDD.n6870 1.5005
R6457 DVDD.n2795 DVDD.n2794 1.5005
R6458 DVDD.n6885 DVDD.n6884 1.5005
R6459 DVDD.n6886 DVDD.n2781 1.5005
R6460 DVDD.n6896 DVDD.n6895 1.5005
R6461 DVDD.n6897 DVDD.n6896 1.5005
R6462 DVDD.n2781 DVDD.n2780 1.5005
R6463 DVDD.n6884 DVDD.n6883 1.5005
R6464 DVDD.n6881 DVDD.n6880 1.5005
R6465 DVDD.n2790 DVDD.n2789 1.5005
R6466 DVDD.n6870 DVDD.n6869 1.5005
R6467 DVDD.n5560 DVDD.n2653 1.5005
R6468 DVDD.n5568 DVDD.n5567 1.5005
R6469 DVDD.n5570 DVDD.n5569 1.5005
R6470 DVDD.n5572 DVDD.n5571 1.5005
R6471 DVDD.n5574 DVDD.n5573 1.5005
R6472 DVDD.n5576 DVDD.n5575 1.5005
R6473 DVDD.n5578 DVDD.n5577 1.5005
R6474 DVDD.n5579 DVDD.n5565 1.5005
R6475 DVDD.n5612 DVDD.n5611 1.5005
R6476 DVDD.n5610 DVDD.n5566 1.5005
R6477 DVDD.n5609 DVDD.n5608 1.5005
R6478 DVDD.n5607 DVDD.n5606 1.5005
R6479 DVDD.n5605 DVDD.n5604 1.5005
R6480 DVDD.n5603 DVDD.n5602 1.5005
R6481 DVDD.n5601 DVDD.n5600 1.5005
R6482 DVDD.n5599 DVDD.n5598 1.5005
R6483 DVDD.n5597 DVDD.n5596 1.5005
R6484 DVDD.n5595 DVDD.n5594 1.5005
R6485 DVDD.n5593 DVDD.n5592 1.5005
R6486 DVDD.n5591 DVDD.n5590 1.5005
R6487 DVDD.n5589 DVDD.n5588 1.5005
R6488 DVDD.n5587 DVDD.n5586 1.5005
R6489 DVDD.n5585 DVDD.n5584 1.5005
R6490 DVDD.n5583 DVDD.n5582 1.5005
R6491 DVDD.n5581 DVDD.n5580 1.5005
R6492 DVDD.n2652 DVDD.n2651 1.5005
R6493 DVDD.n5481 DVDD.n2740 1.5005
R6494 DVDD.n5639 DVDD.n5638 1.5005
R6495 DVDD.n5637 DVDD.n5484 1.5005
R6496 DVDD.n5636 DVDD.n5635 1.5005
R6497 DVDD.n5634 DVDD.n5485 1.5005
R6498 DVDD.n5633 DVDD.n5632 1.5005
R6499 DVDD.n5631 DVDD.n5486 1.5005
R6500 DVDD.n5630 DVDD.n5629 1.5005
R6501 DVDD.n5628 DVDD.n5487 1.5005
R6502 DVDD.n5627 DVDD.n5626 1.5005
R6503 DVDD.n5625 DVDD.n5488 1.5005
R6504 DVDD.n5624 DVDD.n5623 1.5005
R6505 DVDD.n5622 DVDD.n5489 1.5005
R6506 DVDD.n5621 DVDD.n5620 1.5005
R6507 DVDD.n5619 DVDD.n5490 1.5005
R6508 DVDD.n5618 DVDD.n5617 1.5005
R6509 DVDD.n5616 DVDD.n5491 1.5005
R6510 DVDD.n5535 DVDD.n5494 1.5005
R6511 DVDD.n5537 DVDD.n5536 1.5005
R6512 DVDD.n5539 DVDD.n5538 1.5005
R6513 DVDD.n5541 DVDD.n5540 1.5005
R6514 DVDD.n5543 DVDD.n5542 1.5005
R6515 DVDD.n5545 DVDD.n5544 1.5005
R6516 DVDD.n5546 DVDD.n5534 1.5005
R6517 DVDD.n5548 DVDD.n5547 1.5005
R6518 DVDD.n5550 DVDD.n2739 1.5005
R6519 DVDD.n5421 DVDD.n2801 1.5005
R6520 DVDD.n5432 DVDD.n5431 1.5005
R6521 DVDD.n5434 DVDD.n5433 1.5005
R6522 DVDD.n5436 DVDD.n5435 1.5005
R6523 DVDD.n5438 DVDD.n5437 1.5005
R6524 DVDD.n5440 DVDD.n5439 1.5005
R6525 DVDD.n5442 DVDD.n5441 1.5005
R6526 DVDD.n5444 DVDD.n5443 1.5005
R6527 DVDD.n5446 DVDD.n5445 1.5005
R6528 DVDD.n5448 DVDD.n5447 1.5005
R6529 DVDD.n5450 DVDD.n5449 1.5005
R6530 DVDD.n5452 DVDD.n5451 1.5005
R6531 DVDD.n5454 DVDD.n5453 1.5005
R6532 DVDD.n5456 DVDD.n5455 1.5005
R6533 DVDD.n5458 DVDD.n5457 1.5005
R6534 DVDD.n5460 DVDD.n5459 1.5005
R6535 DVDD.n5462 DVDD.n5461 1.5005
R6536 DVDD.n5464 DVDD.n5463 1.5005
R6537 DVDD.n4469 DVDD.n4468 1.5005
R6538 DVDD.n5469 DVDD.n5468 1.5005
R6539 DVDD.n5471 DVDD.n5470 1.5005
R6540 DVDD.n5472 DVDD.n4466 1.5005
R6541 DVDD.n5474 DVDD.n5473 1.5005
R6542 DVDD.n5476 DVDD.n5475 1.5005
R6543 DVDD.n5478 DVDD.n5477 1.5005
R6544 DVDD.n5479 DVDD.n2800 1.5005
R6545 DVDD.n5339 DVDD.n2882 1.5005
R6546 DVDD.n5340 DVDD.n4495 1.5005
R6547 DVDD.n5342 DVDD.n5341 1.5005
R6548 DVDD.n5343 DVDD.n4494 1.5005
R6549 DVDD.n5345 DVDD.n5344 1.5005
R6550 DVDD.n5346 DVDD.n4493 1.5005
R6551 DVDD.n5348 DVDD.n5347 1.5005
R6552 DVDD.n5349 DVDD.n4492 1.5005
R6553 DVDD.n5351 DVDD.n5350 1.5005
R6554 DVDD.n5352 DVDD.n4491 1.5005
R6555 DVDD.n5354 DVDD.n5353 1.5005
R6556 DVDD.n5355 DVDD.n4490 1.5005
R6557 DVDD.n5357 DVDD.n5356 1.5005
R6558 DVDD.n5358 DVDD.n4489 1.5005
R6559 DVDD.n5360 DVDD.n5359 1.5005
R6560 DVDD.n5361 DVDD.n4488 1.5005
R6561 DVDD.n5363 DVDD.n5362 1.5005
R6562 DVDD.n5364 DVDD.n4487 1.5005
R6563 DVDD.n5366 DVDD.n5365 1.5005
R6564 DVDD.n5367 DVDD.n4486 1.5005
R6565 DVDD.n5369 DVDD.n5368 1.5005
R6566 DVDD.n5370 DVDD.n4485 1.5005
R6567 DVDD.n5372 DVDD.n5371 1.5005
R6568 DVDD.n5373 DVDD.n4484 1.5005
R6569 DVDD.n5375 DVDD.n5374 1.5005
R6570 DVDD.n5376 DVDD.n2881 1.5005
R6571 DVDD.n5289 DVDD.n2887 1.5005
R6572 DVDD.n5292 DVDD.n5291 1.5005
R6573 DVDD.n5294 DVDD.n5293 1.5005
R6574 DVDD.n5296 DVDD.n5295 1.5005
R6575 DVDD.n5305 DVDD.n4505 1.5005
R6576 DVDD.n5308 DVDD.n5307 1.5005
R6577 DVDD.n5310 DVDD.n5309 1.5005
R6578 DVDD.n5311 DVDD.n4504 1.5005
R6579 DVDD.n5313 DVDD.n5312 1.5005
R6580 DVDD.n5314 DVDD.n4503 1.5005
R6581 DVDD.n5316 DVDD.n5315 1.5005
R6582 DVDD.n5317 DVDD.n4502 1.5005
R6583 DVDD.n5319 DVDD.n5318 1.5005
R6584 DVDD.n5320 DVDD.n4501 1.5005
R6585 DVDD.n5322 DVDD.n5321 1.5005
R6586 DVDD.n5323 DVDD.n4500 1.5005
R6587 DVDD.n5325 DVDD.n5324 1.5005
R6588 DVDD.n5326 DVDD.n4499 1.5005
R6589 DVDD.n5328 DVDD.n5327 1.5005
R6590 DVDD.n5329 DVDD.n4498 1.5005
R6591 DVDD.n5331 DVDD.n5330 1.5005
R6592 DVDD.n5332 DVDD.n4497 1.5005
R6593 DVDD.n5334 DVDD.n5333 1.5005
R6594 DVDD.n5335 DVDD.n4496 1.5005
R6595 DVDD.n5337 DVDD.n5336 1.5005
R6596 DVDD.n5338 DVDD.n2886 1.5005
R6597 DVDD.n5265 DVDD.n5264 1.5005
R6598 DVDD.n5263 DVDD.n4536 1.5005
R6599 DVDD.n4535 DVDD.n4534 1.5005
R6600 DVDD.n4533 DVDD.n4532 1.5005
R6601 DVDD.n4530 DVDD.n4526 1.5005
R6602 DVDD.n408 DVDD.n407 1.5005
R6603 DVDD.n9364 DVDD.n9363 1.5005
R6604 DVDD.n9366 DVDD.n9365 1.5005
R6605 DVDD.n9368 DVDD.n9367 1.5005
R6606 DVDD.n9370 DVDD.n9369 1.5005
R6607 DVDD.n9372 DVDD.n405 1.5005
R6608 DVDD.n9375 DVDD.n9374 1.5005
R6609 DVDD.n9377 DVDD.n9376 1.5005
R6610 DVDD.n9378 DVDD.n404 1.5005
R6611 DVDD.n9380 DVDD.n9379 1.5005
R6612 DVDD.n9382 DVDD.n9381 1.5005
R6613 DVDD.n9385 DVDD.n9384 1.5005
R6614 DVDD.n9387 DVDD.n9386 1.5005
R6615 DVDD.n9389 DVDD.n9388 1.5005
R6616 DVDD.n379 DVDD.n377 1.5005
R6617 DVDD.n9423 DVDD.n9422 1.5005
R6618 DVDD.n9421 DVDD.n9420 1.5005
R6619 DVDD.n381 DVDD.n380 1.5005
R6620 DVDD.n4522 DVDD.n4521 1.5005
R6621 DVDD.n4525 DVDD.n4524 1.5005
R6622 DVDD.n5267 DVDD.n5266 1.5005
R6623 DVDD.n5219 DVDD.n449 1.5005
R6624 DVDD.n5221 DVDD.n5220 1.5005
R6625 DVDD.n5222 DVDD.n4559 1.5005
R6626 DVDD.n5224 DVDD.n5223 1.5005
R6627 DVDD.n5225 DVDD.n4558 1.5005
R6628 DVDD.n5227 DVDD.n5226 1.5005
R6629 DVDD.n5228 DVDD.n4557 1.5005
R6630 DVDD.n5230 DVDD.n5229 1.5005
R6631 DVDD.n5232 DVDD.n5231 1.5005
R6632 DVDD.n5234 DVDD.n5233 1.5005
R6633 DVDD.n5236 DVDD.n5235 1.5005
R6634 DVDD.n5238 DVDD.n5237 1.5005
R6635 DVDD.n5240 DVDD.n5239 1.5005
R6636 DVDD.n5242 DVDD.n5241 1.5005
R6637 DVDD.n5244 DVDD.n5243 1.5005
R6638 DVDD.n5245 DVDD.n4556 1.5005
R6639 DVDD.n5247 DVDD.n5246 1.5005
R6640 DVDD.n4541 DVDD.n4540 1.5005
R6641 DVDD.n5252 DVDD.n5251 1.5005
R6642 DVDD.n5253 DVDD.n4539 1.5005
R6643 DVDD.n5255 DVDD.n5254 1.5005
R6644 DVDD.n5256 DVDD.n4538 1.5005
R6645 DVDD.n5258 DVDD.n5257 1.5005
R6646 DVDD.n5259 DVDD.n4537 1.5005
R6647 DVDD.n5261 DVDD.n5260 1.5005
R6648 DVDD.n5262 DVDD.n448 1.5005
R6649 DVDD.n4694 DVDD.n4563 1.5005
R6650 DVDD.n4693 DVDD.n4692 1.5005
R6651 DVDD.n4691 DVDD.n4648 1.5005
R6652 DVDD.n4690 DVDD.n4689 1.5005
R6653 DVDD.n4688 DVDD.n4649 1.5005
R6654 DVDD.n4687 DVDD.n4686 1.5005
R6655 DVDD.n4685 DVDD.n4650 1.5005
R6656 DVDD.n4684 DVDD.n4683 1.5005
R6657 DVDD.n4682 DVDD.n4651 1.5005
R6658 DVDD.n4681 DVDD.n4680 1.5005
R6659 DVDD.n4679 DVDD.n4652 1.5005
R6660 DVDD.n4678 DVDD.n4677 1.5005
R6661 DVDD.n4676 DVDD.n4653 1.5005
R6662 DVDD.n4675 DVDD.n4674 1.5005
R6663 DVDD.n4673 DVDD.n4654 1.5005
R6664 DVDD.n4672 DVDD.n4671 1.5005
R6665 DVDD.n4670 DVDD.n4655 1.5005
R6666 DVDD.n4669 DVDD.n4668 1.5005
R6667 DVDD.n4667 DVDD.n4656 1.5005
R6668 DVDD.n4666 DVDD.n4665 1.5005
R6669 DVDD.n4664 DVDD.n4657 1.5005
R6670 DVDD.n4663 DVDD.n4662 1.5005
R6671 DVDD.n4661 DVDD.n4658 1.5005
R6672 DVDD.n4660 DVDD.n4659 1.5005
R6673 DVDD.n4561 DVDD.n4560 1.5005
R6674 DVDD.n5218 DVDD.n5217 1.5005
R6675 DVDD.n4628 DVDD.n4627 1.5005
R6676 DVDD.n4630 DVDD.n4629 1.5005
R6677 DVDD.n4632 DVDD.n4631 1.5005
R6678 DVDD.n4634 DVDD.n4633 1.5005
R6679 DVDD.n4636 DVDD.n4635 1.5005
R6680 DVDD.n4638 DVDD.n4637 1.5005
R6681 DVDD.n4640 DVDD.n4639 1.5005
R6682 DVDD.n4642 DVDD.n4641 1.5005
R6683 DVDD.n4644 DVDD.n4643 1.5005
R6684 DVDD.n4645 DVDD.n4624 1.5005
R6685 DVDD.n4706 DVDD.n4705 1.5005
R6686 DVDD.n4704 DVDD.n4626 1.5005
R6687 DVDD.n4703 DVDD.n4702 1.5005
R6688 DVDD.n4701 DVDD.n4646 1.5005
R6689 DVDD.n4700 DVDD.n4699 1.5005
R6690 DVDD.n4698 DVDD.n4647 1.5005
R6691 DVDD.n4697 DVDD.n4696 1.5005
R6692 DVDD.n4695 DVDD.n4567 1.5005
R6693 DVDD.n397 DVDD.n396 1.5005
R6694 DVDD.n376 DVDD.n177 1.5005
R6695 DVDD.n9583 DVDD.n9582 1.5005
R6696 DVDD.n176 DVDD.n174 1.5005
R6697 DVDD.n180 DVDD.n179 1.5005
R6698 DVDD.n399 DVDD.n374 1.5005
R6699 DVDD.n9401 DVDD.n400 1.5005
R6700 DVDD.n9404 DVDD.n9403 1.5005
R6701 DVDD.n9405 DVDD.n9404 1.5005
R6702 DVDD.n400 DVDD.n398 1.5005
R6703 DVDD.n399 DVDD.n197 1.5005
R6704 DVDD.n9580 DVDD.n177 1.5005
R6705 DVDD.n9582 DVDD.n9581 1.5005
R6706 DVDD.n182 DVDD.n176 1.5005
R6707 DVDD.n8676 DVDD.n1045 1.5005
R6708 DVDD.n8678 DVDD.n8677 1.5005
R6709 DVDD.n233 DVDD.n217 1.5005
R6710 DVDD.n230 DVDD.n214 1.5005
R6711 DVDD.n8693 DVDD.n8690 1.5005
R6712 DVDD.n8695 DVDD.n8694 1.5005
R6713 DVDD.n2890 DVDD.n224 1.5005
R6714 DVDD.n4511 DVDD.n225 1.5005
R6715 DVDD.n5281 DVDD.n5280 1.5005
R6716 DVDD.n4513 DVDD.n4510 1.5005
R6717 DVDD.n5276 DVDD.n5275 1.5005
R6718 DVDD.n2911 DVDD.n2910 1.5005
R6719 DVDD.n2914 DVDD.n2913 1.5005
R6720 DVDD.n2908 DVDD.n2907 1.5005
R6721 DVDD.n2915 DVDD.n2914 1.5005
R6722 DVDD.n2911 DVDD.n2909 1.5005
R6723 DVDD.n238 DVDD.n224 1.5005
R6724 DVDD.n236 DVDD.n225 1.5005
R6725 DVDD.n5280 DVDD.n5279 1.5005
R6726 DVDD.n5278 DVDD.n4513 1.5005
R6727 DVDD.n9352 DVDD.n110 1.5005
R6728 DVDD.n414 DVDD.n109 1.5005
R6729 DVDD.n9358 DVDD.n9357 1.5005
R6730 DVDD.n442 DVDD.n413 1.5005
R6731 DVDD.n441 DVDD.n440 1.5005
R6732 DVDD.n9351 DVDD.n9350 1.5005
R6733 DVDD.n140 DVDD.n138 1.5005
R6734 DVDD.n9604 DVDD.n9603 1.5005
R6735 DVDD.n141 DVDD.n140 1.5005
R6736 DVDD.n9351 DVDD.n9348 1.5005
R6737 DVDD.n9353 DVDD.n9352 1.5005
R6738 DVDD.n9355 DVDD.n414 1.5005
R6739 DVDD.n9357 DVDD.n9356 1.5005
R6740 DVDD.n415 DVDD.n413 1.5005
R6741 DVDD.n903 DVDD.n901 1.5005
R6742 DVDD.n8728 DVDD.n348 1.5005
R6743 DVDD.n8732 DVDD.n8731 1.5005
R6744 DVDD.n8727 DVDD.n8726 1.5005
R6745 DVDD.n8724 DVDD.n876 1.5005
R6746 DVDD.n899 DVDD.n357 1.5005
R6747 DVDD.n900 DVDD.n897 1.5005
R6748 DVDD.n8712 DVDD.n8711 1.5005
R6749 DVDD.n8711 DVDD.n8710 1.5005
R6750 DVDD.n902 DVDD.n900 1.5005
R6751 DVDD.n899 DVDD.n189 1.5005
R6752 DVDD.n8728 DVDD.n194 1.5005
R6753 DVDD.n8731 DVDD.n8730 1.5005
R6754 DVDD.n8729 DVDD.n8727 1.5005
R6755 DVDD.n8758 DVDD.n861 1.5005
R6756 DVDD.n860 DVDD.n859 1.5005
R6757 DVDD.n858 DVDD.n421 1.5005
R6758 DVDD.n9618 DVDD.n102 1.5005
R6759 DVDD.n9619 DVDD.n101 1.5005
R6760 DVDD.n100 DVDD.n95 1.5005
R6761 DVDD.n858 DVDD.n118 1.5005
R6762 DVDD.n9618 DVDD.n9617 1.5005
R6763 DVDD.n9620 DVDD.n9619 1.5005
R6764 DVDD.n95 DVDD.n93 1.5005
R6765 DVDD.n98 DVDD.n97 1.5005
R6766 DVDD.n859 DVDD.n856 1.5005
R6767 DVDD.n8759 DVDD.n8758 1.5005
R6768 DVDD.n8757 DVDD.n8756 1.5005
R6769 DVDD.n8879 DVDD.n8878 1.5005
R6770 DVDD.n8880 DVDD.n658 1.5005
R6771 DVDD.n8882 DVDD.n8881 1.5005
R6772 DVDD.n8883 DVDD.n657 1.5005
R6773 DVDD.n8885 DVDD.n8884 1.5005
R6774 DVDD.n8886 DVDD.n655 1.5005
R6775 DVDD.n8888 DVDD.n8887 1.5005
R6776 DVDD.n656 DVDD.n654 1.5005
R6777 DVDD.n727 DVDD.n726 1.5005
R6778 DVDD.n729 DVDD.n728 1.5005
R6779 DVDD.n731 DVDD.n730 1.5005
R6780 DVDD.n733 DVDD.n732 1.5005
R6781 DVDD.n735 DVDD.n734 1.5005
R6782 DVDD.n737 DVDD.n736 1.5005
R6783 DVDD.n739 DVDD.n738 1.5005
R6784 DVDD.n741 DVDD.n740 1.5005
R6785 DVDD.n743 DVDD.n742 1.5005
R6786 DVDD.n8877 DVDD.n659 1.5005
R6787 DVDD.n6561 DVDD.n6560 1.5005
R6788 DVDD.n6563 DVDD.n6562 1.5005
R6789 DVDD.n6565 DVDD.n6564 1.5005
R6790 DVDD.n6567 DVDD.n6566 1.5005
R6791 DVDD.n6569 DVDD.n6568 1.5005
R6792 DVDD.n6571 DVDD.n6570 1.5005
R6793 DVDD.n6573 DVDD.n6572 1.5005
R6794 DVDD.n6575 DVDD.n6574 1.5005
R6795 DVDD.n6577 DVDD.n6576 1.5005
R6796 DVDD.n6579 DVDD.n6578 1.5005
R6797 DVDD.n6581 DVDD.n6580 1.5005
R6798 DVDD.n6583 DVDD.n6582 1.5005
R6799 DVDD.n6585 DVDD.n6584 1.5005
R6800 DVDD.n6587 DVDD.n6586 1.5005
R6801 DVDD.n6559 DVDD.n6558 1.5005
R6802 DVDD.n6589 DVDD.n6588 1.5005
R6803 DVDD.n6590 DVDD.n6486 1.5005
R6804 DVDD.n6592 DVDD.n6591 1.5005
R6805 DVDD.n6487 DVDD.n6477 1.5005
R6806 DVDD.n6545 DVDD.n6544 1.5005
R6807 DVDD.n6547 DVDD.n6546 1.5005
R6808 DVDD.n6549 DVDD.n6548 1.5005
R6809 DVDD.n6551 DVDD.n6550 1.5005
R6810 DVDD.n6553 DVDD.n6552 1.5005
R6811 DVDD.n6555 DVDD.n6554 1.5005
R6812 DVDD.n6557 DVDD.n6556 1.5005
R6813 DVDD.n3414 DVDD.n3413 1.5005
R6814 DVDD.n3430 DVDD.n3429 1.5005
R6815 DVDD.n3432 DVDD.n3431 1.5005
R6816 DVDD.n3434 DVDD.n3433 1.5005
R6817 DVDD.n3436 DVDD.n3435 1.5005
R6818 DVDD.n3438 DVDD.n3437 1.5005
R6819 DVDD.n3440 DVDD.n3439 1.5005
R6820 DVDD.n3442 DVDD.n3441 1.5005
R6821 DVDD.n6469 DVDD.n6468 1.5005
R6822 DVDD.n3444 DVDD.n3443 1.5005
R6823 DVDD.n3445 DVDD.n3428 1.5005
R6824 DVDD.n3447 DVDD.n3446 1.5005
R6825 DVDD.n3448 DVDD.n3427 1.5005
R6826 DVDD.n3450 DVDD.n3449 1.5005
R6827 DVDD.n3451 DVDD.n3426 1.5005
R6828 DVDD.n3453 DVDD.n3452 1.5005
R6829 DVDD.n3454 DVDD.n3425 1.5005
R6830 DVDD.n3456 DVDD.n3455 1.5005
R6831 DVDD.n3457 DVDD.n3424 1.5005
R6832 DVDD.n3459 DVDD.n3458 1.5005
R6833 DVDD.n3460 DVDD.n3423 1.5005
R6834 DVDD.n3462 DVDD.n3461 1.5005
R6835 DVDD.n3463 DVDD.n3422 1.5005
R6836 DVDD.n3465 DVDD.n3464 1.5005
R6837 DVDD.n3466 DVDD.n3418 1.5005
R6838 DVDD.n6467 DVDD.n6466 1.5005
R6839 DVDD.n6379 DVDD.n6378 1.5005
R6840 DVDD.n6381 DVDD.n6380 1.5005
R6841 DVDD.n6377 DVDD.n6376 1.5005
R6842 DVDD.n6383 DVDD.n6382 1.5005
R6843 DVDD.n6384 DVDD.n3552 1.5005
R6844 DVDD.n6386 DVDD.n6385 1.5005
R6845 DVDD.n3553 DVDD.n3546 1.5005
R6846 DVDD.n6339 DVDD.n6338 1.5005
R6847 DVDD.n6341 DVDD.n6340 1.5005
R6848 DVDD.n6343 DVDD.n6342 1.5005
R6849 DVDD.n6345 DVDD.n6344 1.5005
R6850 DVDD.n6347 DVDD.n6346 1.5005
R6851 DVDD.n6349 DVDD.n6348 1.5005
R6852 DVDD.n6351 DVDD.n6350 1.5005
R6853 DVDD.n6353 DVDD.n6352 1.5005
R6854 DVDD.n6355 DVDD.n6354 1.5005
R6855 DVDD.n6357 DVDD.n6356 1.5005
R6856 DVDD.n6359 DVDD.n6358 1.5005
R6857 DVDD.n6361 DVDD.n6360 1.5005
R6858 DVDD.n6363 DVDD.n6362 1.5005
R6859 DVDD.n6365 DVDD.n6364 1.5005
R6860 DVDD.n6367 DVDD.n6366 1.5005
R6861 DVDD.n6369 DVDD.n6368 1.5005
R6862 DVDD.n6371 DVDD.n6370 1.5005
R6863 DVDD.n6373 DVDD.n6372 1.5005
R6864 DVDD.n6375 DVDD.n6374 1.5005
R6865 DVDD.n3766 DVDD.n3765 1.5005
R6866 DVDD.n3767 DVDD.n3763 1.5005
R6867 DVDD.n3769 DVDD.n3768 1.5005
R6868 DVDD.n3770 DVDD.n3762 1.5005
R6869 DVDD.n3772 DVDD.n3771 1.5005
R6870 DVDD.n3773 DVDD.n3761 1.5005
R6871 DVDD.n3775 DVDD.n3774 1.5005
R6872 DVDD.n3776 DVDD.n3760 1.5005
R6873 DVDD.n3778 DVDD.n3777 1.5005
R6874 DVDD.n3779 DVDD.n3759 1.5005
R6875 DVDD.n3781 DVDD.n3780 1.5005
R6876 DVDD.n3782 DVDD.n3758 1.5005
R6877 DVDD.n3784 DVDD.n3783 1.5005
R6878 DVDD.n3785 DVDD.n3757 1.5005
R6879 DVDD.n3787 DVDD.n3786 1.5005
R6880 DVDD.n3788 DVDD.n3756 1.5005
R6881 DVDD.n3790 DVDD.n3789 1.5005
R6882 DVDD.n3791 DVDD.n3755 1.5005
R6883 DVDD.n3793 DVDD.n3792 1.5005
R6884 DVDD.n3794 DVDD.n3754 1.5005
R6885 DVDD.n3796 DVDD.n3795 1.5005
R6886 DVDD.n3797 DVDD.n3753 1.5005
R6887 DVDD.n3799 DVDD.n3798 1.5005
R6888 DVDD.n3800 DVDD.n3578 1.5005
R6889 DVDD.n3802 DVDD.n3801 1.5005
R6890 DVDD.n3764 DVDD.n3576 1.5005
R6891 DVDD.n1376 DVDD.n1374 1.21934
R6892 DVDD.n1342 DVDD.n1341 1.21934
R6893 DVDD.n8911 DVDD.n32 1.19814
R6894 DVDD.n4818 DVDD.n4817 1.19814
R6895 DVDD.n8668 DVDD.n8667 1.19707
R6896 DVDD.n6776 DVDD.n6775 1.19707
R6897 DVDD.n9319 DVDD.n429 1.1255
R6898 DVDD.n9316 DVDD.n435 1.1255
R6899 DVDD.n4531 DVDD.n434 1.1255
R6900 DVDD.n4529 DVDD.n4528 1.1255
R6901 DVDD.n9362 DVDD.n9361 1.1255
R6902 DVDD.n9616 DVDD.n107 1.1255
R6903 DVDD.n9613 DVDD.n130 1.1255
R6904 DVDD.n9327 DVDD.n406 1.1255
R6905 DVDD.n9371 DVDD.n137 1.1255
R6906 DVDD.n9373 DVDD.n145 1.1255
R6907 DVDD.n9599 DVDD.n147 1.1255
R6908 DVDD.n9596 DVDD.n153 1.1255
R6909 DVDD.n9383 DVDD.n152 1.1255
R6910 DVDD.n9589 DVDD.n168 1.1255
R6911 DVDD.n9586 DVDD.n171 1.1255
R6912 DVDD.n9391 DVDD.n9390 1.1255
R6913 DVDD.n9425 DVDD.n9424 1.1255
R6914 DVDD.n9398 DVDD.n378 1.1255
R6915 DVDD.n9419 DVDD.n9418 1.1255
R6916 DVDD.n9415 DVDD.n386 1.1255
R6917 DVDD.n4523 DVDD.n385 1.1255
R6918 DVDD.n4520 DVDD.n394 1.1255
R6919 DVDD.n5269 DVDD.n5268 1.1255
R6920 DVDD.n5272 DVDD.n4518 1.1255
R6921 DVDD.n4517 DVDD.n4516 1.1255
R6922 DVDD.n5284 DVDD.n4506 1.1255
R6923 DVDD.n5288 DVDD.n5287 1.1255
R6924 DVDD.n5290 DVDD.n228 1.1255
R6925 DVDD.n6791 DVDD.n2895 1.1255
R6926 DVDD.n6788 DVDD.n2899 1.1255
R6927 DVDD.n5304 DVDD.n5303 1.1255
R6928 DVDD.n5306 DVDD.n2906 1.1255
R6929 DVDD.n6777 DVDD.n2958 1.1255
R6930 DVDD.n9425 DVDD.n356 1.1255
R6931 DVDD.n4155 DVDD.n4151 1.1255
R6932 DVDD.n4207 DVDD.n4206 1.1255
R6933 DVDD.n4160 DVDD.n4153 1.1255
R6934 DVDD.n3977 DVDD.n3976 1.1255
R6935 DVDD.n4134 DVDD.n3983 1.1255
R6936 DVDD.n4136 DVDD.n4135 1.1255
R6937 DVDD.n4133 DVDD.n3981 1.1255
R6938 DVDD.n4132 DVDD.n4131 1.1255
R6939 DVDD.n3994 DVDD.n3992 1.1255
R6940 DVDD.n9425 DVDD.n372 1.1255
R6941 DVDD.n4079 DVDD.n4078 1.1255
R6942 DVDD.n4064 DVDD.n4027 1.1255
R6943 DVDD.n4045 DVDD.n4034 1.1255
R6944 DVDD.n4047 DVDD.n4046 1.1255
R6945 DVDD.n4043 DVDD.n4042 1.1255
R6946 DVDD.n4102 DVDD.n4101 1.1255
R6947 DVDD.n4011 DVDD.n4001 1.1255
R6948 DVDD.n4010 DVDD.n4009 1.1255
R6949 DVDD.n4004 DVDD.n3999 1.1255
R6950 DVDD.n4112 DVDD.n4111 1.1255
R6951 DVDD.n9616 DVDD.n112 1.1255
R6952 DVDD.n4096 DVDD.n4095 1.1255
R6953 DVDD.n4036 DVDD.n4017 1.1255
R6954 DVDD.n4032 DVDD.n4031 1.1255
R6955 DVDD.n4059 DVDD.n4058 1.1255
R6956 DVDD.n4062 DVDD.n4061 1.1255
R6957 DVDD.n4073 DVDD.n4072 1.1255
R6958 DVDD.n4069 DVDD.n3991 1.1255
R6959 DVDD.n4123 DVDD.n4122 1.1255
R6960 DVDD.n4146 DVDD.n4145 1.1255
R6961 DVDD.n4218 DVDD.n228 1.1255
R6962 DVDD.n4216 DVDD.n4215 1.1255
R6963 DVDD.n4158 DVDD.n4149 1.1255
R6964 DVDD.n9472 DVDD.n9471 1.1255
R6965 DVDD.n300 DVDD.n290 1.1255
R6966 DVDD.n302 DVDD.n293 1.1255
R6967 DVDD.n9466 DVDD.n9465 1.1255
R6968 DVDD.n297 DVDD.n296 1.1255
R6969 DVDD.n9616 DVDD.n125 1.1255
R6970 DVDD.n9458 DVDD.n9457 1.1255
R6971 DVDD.n316 DVDD.n308 1.1255
R6972 DVDD.n9452 DVDD.n9451 1.1255
R6973 DVDD.n322 DVDD.n315 1.1255
R6974 DVDD.n9446 DVDD.n9445 1.1255
R6975 DVDD.n338 DVDD.n337 1.1255
R6976 DVDD.n339 DVDD.n329 1.1255
R6977 DVDD.n9439 DVDD.n9438 1.1255
R6978 DVDD.n346 DVDD.n344 1.1255
R6979 DVDD.n9432 DVDD.n9431 1.1255
R6980 DVDD.n9425 DVDD.n370 1.1255
R6981 DVDD.n364 DVDD.n363 1.1255
R6982 DVDD.n365 DVDD.n281 1.1255
R6983 DVDD.n9483 DVDD.n9482 1.1255
R6984 DVDD.n284 DVDD.n282 1.1255
R6985 DVDD.n9492 DVDD.n9491 1.1255
R6986 DVDD.n9493 DVDD.n272 1.1255
R6987 DVDD.n9496 DVDD.n9495 1.1255
R6988 DVDD.n9494 DVDD.n274 1.1255
R6989 DVDD.n268 DVDD.n267 1.1255
R6990 DVDD.n9506 DVDD.n9505 1.1255
R6991 DVDD.n9509 DVDD.n228 1.1255
R6992 DVDD.n9507 DVDD.n243 1.1255
R6993 DVDD.n9556 DVDD.n9555 1.1255
R6994 DVDD.n251 DVDD.n249 1.1255
R6995 DVDD.n9549 DVDD.n9548 1.1255
R6996 DVDD.n9547 DVDD.n9546 1.1255
R6997 DVDD.n9425 DVDD.n375 1.1255
R6998 DVDD.n9616 DVDD.n126 1.1255
R6999 DVDD.n6794 DVDD.n228 1.1255
R7000 DVDD.n9616 DVDD.n114 1.1255
R7001 DVDD.n1040 DVDD.n228 1.1255
R7002 DVDD.n8788 DVDD.n46 1.1255
R7003 DVDD.n9627 DVDD.n9626 1.1255
R7004 DVDD.n9625 DVDD.n85 1.1255
R7005 DVDD.n9624 DVDD.n9623 1.1255
R7006 DVDD.n8772 DVDD.n87 1.1255
R7007 DVDD.n9616 DVDD.n113 1.1255
R7008 DVDD.n8765 DVDD.n8764 1.1255
R7009 DVDD.n8763 DVDD.n8762 1.1255
R7010 DVDD.n942 DVDD.n852 1.1255
R7011 DVDD.n8753 DVDD.n8752 1.1255
R7012 DVDD.n8751 DVDD.n867 1.1255
R7013 DVDD.n8750 DVDD.n8749 1.1255
R7014 DVDD.n871 DVDD.n869 1.1255
R7015 DVDD.n977 DVDD.n885 1.1255
R7016 DVDD.n8738 DVDD.n8737 1.1255
R7017 DVDD.n8736 DVDD.n8735 1.1255
R7018 DVDD.n9425 DVDD.n351 1.1255
R7019 DVDD.n8718 DVDD.n8717 1.1255
R7020 DVDD.n8716 DVDD.n8715 1.1255
R7021 DVDD.n919 DVDD.n893 1.1255
R7022 DVDD.n995 DVDD.n909 1.1255
R7023 DVDD.n8706 DVDD.n8705 1.1255
R7024 DVDD.n8704 DVDD.n8703 1.1255
R7025 DVDD.n8700 DVDD.n910 1.1255
R7026 DVDD.n1014 DVDD.n1003 1.1255
R7027 DVDD.n1035 DVDD.n1034 1.1255
R7028 DVDD.n8686 DVDD.n8685 1.1255
R7029 DVDD.n8684 DVDD.n228 1.1255
R7030 DVDD.n8683 DVDD.n8682 1.1255
R7031 DVDD.n3742 DVDD.n1036 1.1255
R7032 DVDD.n3634 DVDD.n1054 1.1255
R7033 DVDD.n8670 DVDD.n8669 1.1255
R7034 DVDD.n8668 DVDD.n1052 1.1255
R7035 DVDD.n9319 DVDD.n9318 1.1255
R7036 DVDD.n9317 DVDD.n9316 1.1255
R7037 DVDD.n434 DVDD.n433 1.1255
R7038 DVDD.n4528 DVDD.n4527 1.1255
R7039 DVDD.n9361 DVDD.n127 1.1255
R7040 DVDD.n9616 DVDD.n9615 1.1255
R7041 DVDD.n9614 DVDD.n9613 1.1255
R7042 DVDD.n9327 DVDD.n128 1.1255
R7043 DVDD.n148 DVDD.n137 1.1255
R7044 DVDD.n149 DVDD.n145 1.1255
R7045 DVDD.n9599 DVDD.n9598 1.1255
R7046 DVDD.n9597 DVDD.n9596 1.1255
R7047 DVDD.n152 DVDD.n150 1.1255
R7048 DVDD.n9589 DVDD.n9588 1.1255
R7049 DVDD.n9587 DVDD.n9586 1.1255
R7050 DVDD.n9391 DVDD.n169 1.1255
R7051 DVDD.n9425 DVDD.n359 1.1255
R7052 DVDD.n9398 DVDD.n383 1.1255
R7053 DVDD.n9418 DVDD.n9417 1.1255
R7054 DVDD.n9416 DVDD.n9415 1.1255
R7055 DVDD.n385 DVDD.n384 1.1255
R7056 DVDD.n4519 DVDD.n394 1.1255
R7057 DVDD.n5270 DVDD.n5269 1.1255
R7058 DVDD.n5272 DVDD.n5271 1.1255
R7059 DVDD.n4516 DVDD.n4507 1.1255
R7060 DVDD.n5285 DVDD.n5284 1.1255
R7061 DVDD.n5287 DVDD.n5286 1.1255
R7062 DVDD.n2896 DVDD.n228 1.1255
R7063 DVDD.n6791 DVDD.n6790 1.1255
R7064 DVDD.n6789 DVDD.n6788 1.1255
R7065 DVDD.n5303 DVDD.n2897 1.1255
R7066 DVDD.n2959 DVDD.n2906 1.1255
R7067 DVDD.n6777 DVDD.n6776 1.1255
R7068 DVDD.n1884 DVDD.n1883 0.902365
R7069 DVDD.n1883 DVDD.n1866 0.902314
R7070 DVDD.n1870 DVDD.n1562 0.902208
R7071 DVDD.n7677 DVDD.n7676 0.902208
R7072 DVDD.n2448 DVDD.n2447 0.902208
R7073 DVDD.n2425 DVDD.n2424 0.902208
R7074 DVDD.n7665 DVDD.n1983 0.902195
R7075 DVDD.n2434 DVDD.n2432 0.902195
R7076 DVDD.n2411 DVDD.n2409 0.902195
R7077 DVDD.n7665 DVDD.n7664 0.902164
R7078 DVDD.n2434 DVDD.n2433 0.902164
R7079 DVDD.n2411 DVDD.n2410 0.902164
R7080 DVDD.n2424 DVDD.n2404 0.901912
R7081 DVDD.n2447 DVDD.n2427 0.901912
R7082 DVDD.n7676 DVDD.n2450 0.901912
R7083 DVDD.n1870 DVDD.n1561 0.901912
R7084 DVDD.n1872 DVDD.n1870 0.886486
R7085 DVDD.n7676 DVDD.n7675 0.886486
R7086 DVDD.n2447 DVDD.n2446 0.886486
R7087 DVDD.n2424 DVDD.n2423 0.886486
R7088 DVDD.n2412 DVDD.n2411 0.886311
R7089 DVDD.n2435 DVDD.n2434 0.886311
R7090 DVDD.n7666 DVDD.n7665 0.886311
R7091 DVDD.n1883 DVDD.n1882 0.88609
R7092 DVDD.n8193 DVDD.n8192 0.85991
R7093 DVDD.n9406 DVDD.n9405 0.770072
R7094 DVDD.n9602 DVDD.n141 0.770072
R7095 DVDD.n8710 DVDD.n8709 0.770072
R7096 DVDD.n3870 DVDD.n3865 0.769684
R7097 DVDD.n6243 DVDD.n6237 0.769684
R7098 DVDD.n6869 DVDD.n6868 0.769684
R7099 DVDD.n6898 DVDD.n6897 0.769684
R7100 DVDD.n182 DVDD.n181 0.769684
R7101 DVDD.n8694 DVDD.n8692 0.769684
R7102 DVDD.n8676 DVDD.n8675 0.769684
R7103 DVDD.n5278 DVDD.n5277 0.769684
R7104 DVDD.n2916 DVDD.n2915 0.769684
R7105 DVDD.n439 DVDD.n415 0.769684
R7106 DVDD.n8729 DVDD.n875 0.769684
R7107 DVDD.n100 DVDD.n99 0.769684
R7108 DVDD.n862 DVDD.n861 0.769684
R7109 DVDD.n6457 DVDD.n3421 0.760008
R7110 DVDD.n3492 DVDD.n3490 0.75924
R7111 DVDD.n7687 DVDD.n7686 0.757185
R7112 DVDD.n7689 DVDD.n7687 0.757185
R7113 DVDD.n7734 DVDD.n7729 0.757185
R7114 DVDD.n7729 DVDD.n2341 0.757185
R7115 DVDD.n6459 DVDD.n6458 0.7505
R7116 DVDD.n6448 DVDD.n6447 0.7505
R7117 DVDD.n3496 DVDD.n3488 0.7505
R7118 DVDD.n3499 DVDD.n3498 0.7505
R7119 DVDD.n3494 DVDD.n3491 0.7505
R7120 DVDD.n6450 DVDD.n3486 0.7505
R7121 DVDD.n6454 DVDD.n6453 0.7505
R7122 DVDD.n3484 DVDD.n3483 0.7505
R7123 DVDD.n6456 DVDD.n3484 0.7505
R7124 DVDD.n6455 DVDD.n6454 0.7505
R7125 DVDD.n3486 DVDD.n3485 0.7505
R7126 DVDD.n6447 DVDD.n6446 0.7505
R7127 DVDD.n3501 DVDD.n3488 0.7505
R7128 DVDD.n3500 DVDD.n3499 0.7505
R7129 DVDD.n355 DVDD.n354 0.7505
R7130 DVDD.n354 DVDD.n193 0.7505
R7131 DVDD.n7353 DVDD.n7352 0.746446
R7132 DVDD.n8624 DVDD.n8623 0.746446
R7133 DVDD.n8546 DVDD.n8545 0.746446
R7134 DVDD.n8539 DVDD.n8538 0.746446
R7135 DVDD.n8549 DVDD.n8548 0.690924
R7136 DVDD.n8532 DVDD.n8531 0.690922
R7137 DVDD DVDD.n744 0.654219
R7138 DVDD DVDD.n4568 0.652634
R7139 DVDD DVDD.n9015 0.649902
R7140 DVDD DVDD.n725 0.649902
R7141 DVDD DVDD.n4879 0.649902
R7142 DVDD DVDD.n5159 0.649902
R7143 DVDD.n7200 DVDD.n1500 0.648577
R7144 DVDD.n8385 DVDD.n1500 0.648577
R7145 DVDD.n8642 DVDD.n1303 0.648577
R7146 DVDD.n8645 DVDD.n8642 0.648577
R7147 DVDD DVDD.n4880 0.630979
R7148 DVDD.n4880 DVDD 0.630979
R7149 DVDD DVDD.n4951 0.630979
R7150 DVDD.n4951 DVDD 0.630979
R7151 DVDD DVDD.n4901 0.630979
R7152 DVDD.n4901 DVDD 0.630979
R7153 DVDD DVDD.n9476 0.630979
R7154 DVDD.n9476 DVDD 0.630979
R7155 DVDD DVDD.n9512 0.630979
R7156 DVDD.n9512 DVDD 0.630979
R7157 DVDD DVDD.n4373 0.630979
R7158 DVDD.n4373 DVDD 0.630979
R7159 DVDD DVDD.n5821 0.630979
R7160 DVDD.n5821 DVDD 0.630979
R7161 DVDD DVDD.n5840 0.630979
R7162 DVDD.n5840 DVDD 0.630979
R7163 DVDD DVDD.n3141 0.630979
R7164 DVDD.n3141 DVDD 0.630979
R7165 DVDD DVDD.n9016 0.630979
R7166 DVDD.n9016 DVDD 0.630979
R7167 DVDD DVDD.n9072 0.630979
R7168 DVDD.n9072 DVDD 0.630979
R7169 DVDD DVDD.n9108 0.630979
R7170 DVDD.n9108 DVDD 0.630979
R7171 DVDD DVDD.n4116 0.630979
R7172 DVDD.n4116 DVDD 0.630979
R7173 DVDD DVDD.n4221 0.630979
R7174 DVDD.n4221 DVDD 0.630979
R7175 DVDD DVDD.n4277 0.630979
R7176 DVDD.n4277 DVDD 0.630979
R7177 DVDD DVDD.n6054 0.630979
R7178 DVDD.n6054 DVDD 0.630979
R7179 DVDD DVDD.n5942 0.630979
R7180 DVDD.n5942 DVDD 0.630979
R7181 DVDD DVDD.n3250 0.630979
R7182 DVDD.n3250 DVDD 0.630979
R7183 DVDD.n4997 DVDD 0.610636
R7184 DVDD.n4994 DVDD 0.610636
R7185 DVDD.n4952 DVDD 0.610636
R7186 DVDD.n4949 DVDD 0.610636
R7187 DVDD.n4902 DVDD 0.610636
R7188 DVDD DVDD.n9475 0.610636
R7189 DVDD.n9477 DVDD 0.610636
R7190 DVDD DVDD.n9511 0.610636
R7191 DVDD.n9513 DVDD 0.610636
R7192 DVDD DVDD.n4372 0.610636
R7193 DVDD.n4374 DVDD 0.610636
R7194 DVDD DVDD.n5820 0.610636
R7195 DVDD.n5822 DVDD 0.610636
R7196 DVDD DVDD.n5831 0.610636
R7197 DVDD.n5842 DVDD 0.610636
R7198 DVDD DVDD.n3140 0.610636
R7199 DVDD.n3143 DVDD 0.610636
R7200 DVDD.n9017 DVDD 0.610636
R7201 DVDD.n9073 DVDD 0.610636
R7202 DVDD DVDD.n9071 0.610636
R7203 DVDD.n9109 DVDD 0.610636
R7204 DVDD DVDD.n9107 0.610636
R7205 DVDD.n4117 DVDD 0.610636
R7206 DVDD DVDD.n4115 0.610636
R7207 DVDD.n4222 DVDD 0.610636
R7208 DVDD DVDD.n4220 0.610636
R7209 DVDD.n4278 DVDD 0.610636
R7210 DVDD DVDD.n4276 0.610636
R7211 DVDD.n6056 DVDD 0.610636
R7212 DVDD DVDD.n6053 0.610636
R7213 DVDD.n5944 DVDD 0.610636
R7214 DVDD.n5991 DVDD 0.610636
R7215 DVDD.n3252 DVDD 0.610636
R7216 DVDD DVDD.n3249 0.610636
R7217 DVDD.n5160 DVDD 0.610636
R7218 DVDD DVDD.n4562 0.610636
R7219 DVDD DVDD.n5216 0.610636
R7220 DVDD.n9300 DVDD 0.610636
R7221 DVDD DVDD.n9299 0.610636
R7222 DVDD DVDD.n391 0.610636
R7223 DVDD DVDD.n445 0.610636
R7224 DVDD.n6797 DVDD 0.610636
R7225 DVDD DVDD.n6796 0.610636
R7226 DVDD.n6852 DVDD 0.610636
R7227 DVDD DVDD.n6851 0.610636
R7228 DVDD.n6860 DVDD 0.610636
R7229 DVDD DVDD.n6859 0.610636
R7230 DVDD.n6904 DVDD 0.610636
R7231 DVDD DVDD.n6902 0.610636
R7232 DVDD.n6929 DVDD 0.610636
R7233 DVDD DVDD.n6927 0.610636
R7234 DVDD.n745 DVDD 0.610636
R7235 DVDD DVDD.n8837 0.610636
R7236 DVDD.n748 DVDD 0.610636
R7237 DVDD DVDD.n78 0.610636
R7238 DVDD.n8834 DVDD 0.610636
R7239 DVDD DVDD.n999 0.610636
R7240 DVDD.n9632 DVDD 0.610636
R7241 DVDD DVDD.n3581 0.610636
R7242 DVDD DVDD.n3582 0.610636
R7243 DVDD.n3803 DVDD 0.610636
R7244 DVDD DVDD.n3577 0.610636
R7245 DVDD DVDD.n3554 0.610636
R7246 DVDD DVDD.n6337 0.610636
R7247 DVDD DVDD.n3416 0.610636
R7248 DVDD DVDD.n3417 0.610636
R7249 DVDD DVDD.n6489 0.610636
R7250 DVDD DVDD.n6543 0.610636
R7251 DVDD.n725 DVDD.n579 0.607735
R7252 DVDD.n9015 DVDD.n9014 0.607735
R7253 DVDD.n4879 DVDD.n4867 0.607735
R7254 DVDD.n5159 DVDD.n5158 0.607735
R7255 DVDD DVDD.n4567 0.607216
R7256 DVDD.n5217 DVDD 0.607216
R7257 DVDD DVDD.n4563 0.607216
R7258 DVDD DVDD.n448 0.607216
R7259 DVDD DVDD.n449 0.607216
R7260 DVDD.n5266 DVDD 0.607216
R7261 DVDD DVDD.n5265 0.607216
R7262 DVDD DVDD.n2886 0.607216
R7263 DVDD DVDD.n2887 0.607216
R7264 DVDD DVDD.n2881 0.607216
R7265 DVDD DVDD.n2882 0.607216
R7266 DVDD DVDD.n2800 0.607216
R7267 DVDD DVDD.n2801 0.607216
R7268 DVDD DVDD.n2739 0.607216
R7269 DVDD DVDD.n2740 0.607216
R7270 DVDD DVDD.n2652 0.607216
R7271 DVDD DVDD.n2653 0.607216
R7272 DVDD DVDD.n659 0.607216
R7273 DVDD.n8838 DVDD 0.607216
R7274 DVDD.n8875 DVDD 0.607216
R7275 DVDD DVDD.n8796 0.607216
R7276 DVDD DVDD.n790 0.607216
R7277 DVDD.n1000 DVDD 0.607216
R7278 DVDD.n8793 DVDD 0.607216
R7279 DVDD.n3751 DVDD 0.607216
R7280 DVDD DVDD.n3750 0.607216
R7281 DVDD DVDD.n3576 0.607216
R7282 DVDD DVDD.n3802 0.607216
R7283 DVDD.n6377 DVDD 0.607216
R7284 DVDD DVDD.n6375 0.607216
R7285 DVDD.n6468 DVDD 0.607216
R7286 DVDD DVDD.n6467 0.607216
R7287 DVDD.n6559 DVDD 0.607216
R7288 DVDD DVDD.n6557 0.607216
R7289 DVDD.n8388 DVDD.n1497 0.581851
R7290 DVDD.n8626 DVDD.n1326 0.581851
R7291 DVDD.n8617 DVDD.n1338 0.5255
R7292 DVDD.n8617 DVDD.n8616 0.5255
R7293 DVDD.n8396 DVDD.n1336 0.5255
R7294 DVDD.n8587 DVDD.n1336 0.5255
R7295 DVDD.n8586 DVDD.n8585 0.5255
R7296 DVDD.n8587 DVDD.n8586 0.5255
R7297 DVDD.n8475 DVDD.n1339 0.5255
R7298 DVDD.n8616 DVDD.n1339 0.5255
R7299 DVDD.n8615 DVDD.n8614 0.5255
R7300 DVDD.n8616 DVDD.n8615 0.5255
R7301 DVDD.n8565 DVDD.n1371 0.5255
R7302 DVDD.n8587 DVDD.n1371 0.5255
R7303 DVDD.n8588 DVDD.n1373 0.5255
R7304 DVDD.n8588 DVDD.n8587 0.5255
R7305 DVDD.n8523 DVDD.n1340 0.5255
R7306 DVDD.n8616 DVDD.n1340 0.5255
R7307 DVDD.n2418 DVDD 0.5054
R7308 DVDD DVDD.n2417 0.5054
R7309 DVDD.n2441 DVDD 0.5054
R7310 DVDD DVDD.n2440 0.5054
R7311 DVDD.n7672 DVDD 0.5054
R7312 DVDD DVDD.n7671 0.5054
R7313 DVDD DVDD.n1875 0.5054
R7314 DVDD.n1876 DVDD 0.5054
R7315 DVDD.n8619 DVDD.n1335 0.455365
R7316 DVDD.n8621 DVDD.n8619 0.455365
R7317 DVDD.n8543 DVDD.n8542 0.455365
R7318 DVDD.n8542 DVDD.n8541 0.455365
R7319 DVDD.n598 DVDD.n597 0.4505
R7320 DVDD.n599 DVDD.n594 0.4505
R7321 DVDD.n8934 DVDD.n8933 0.4505
R7322 DVDD.n8932 DVDD.n595 0.4505
R7323 DVDD.n8931 DVDD.n8930 0.4505
R7324 DVDD.n601 DVDD.n600 0.4505
R7325 DVDD.n8926 DVDD.n8925 0.4505
R7326 DVDD.n8924 DVDD.n603 0.4505
R7327 DVDD.n8923 DVDD.n8922 0.4505
R7328 DVDD.n605 DVDD.n604 0.4505
R7329 DVDD.n8918 DVDD.n8917 0.4505
R7330 DVDD.n8916 DVDD.n607 0.4505
R7331 DVDD.n8915 DVDD.n8914 0.4505
R7332 DVDD.n609 DVDD.n608 0.4505
R7333 DVDD.n8908 DVDD.n8907 0.4505
R7334 DVDD.n8906 DVDD.n634 0.4505
R7335 DVDD.n8905 DVDD.n8904 0.4505
R7336 DVDD.n636 DVDD.n635 0.4505
R7337 DVDD.n8900 DVDD.n8899 0.4505
R7338 DVDD.n8898 DVDD.n638 0.4505
R7339 DVDD.n8897 DVDD.n8896 0.4505
R7340 DVDD.n640 DVDD.n639 0.4505
R7341 DVDD.n8890 DVDD.n8889 0.4505
R7342 DVDD.n4612 DVDD.n4611 0.4505
R7343 DVDD.n4716 DVDD.n4715 0.4505
R7344 DVDD.n4717 DVDD.n4610 0.4505
R7345 DVDD.n4719 DVDD.n4718 0.4505
R7346 DVDD.n4608 DVDD.n4607 0.4505
R7347 DVDD.n4724 DVDD.n4723 0.4505
R7348 DVDD.n4725 DVDD.n4606 0.4505
R7349 DVDD.n4727 DVDD.n4726 0.4505
R7350 DVDD.n4592 DVDD.n4591 0.4505
R7351 DVDD.n4824 DVDD.n4823 0.4505
R7352 DVDD.n4825 DVDD.n4590 0.4505
R7353 DVDD.n4827 DVDD.n4826 0.4505
R7354 DVDD.n4588 DVDD.n4587 0.4505
R7355 DVDD.n4832 DVDD.n4831 0.4505
R7356 DVDD.n4833 DVDD.n4586 0.4505
R7357 DVDD.n4835 DVDD.n4834 0.4505
R7358 DVDD.n4584 DVDD.n4583 0.4505
R7359 DVDD.n4840 DVDD.n4839 0.4505
R7360 DVDD.n4841 DVDD.n4580 0.4505
R7361 DVDD.n5114 DVDD.n5113 0.4505
R7362 DVDD.n5112 DVDD.n4582 0.4505
R7363 DVDD.n5111 DVDD.n5110 0.4505
R7364 DVDD.n5108 DVDD.n4842 0.4505
R7365 DVDD.n4846 DVDD.n4843 0.4505
R7366 DVDD.n5104 DVDD.n5103 0.4505
R7367 DVDD.n5102 DVDD.n4845 0.4505
R7368 DVDD.n5101 DVDD.n5100 0.4505
R7369 DVDD.n4848 DVDD.n4847 0.4505
R7370 DVDD.n5096 DVDD.n5095 0.4505
R7371 DVDD.n5094 DVDD.n4850 0.4505
R7372 DVDD.n5093 DVDD.n5092 0.4505
R7373 DVDD.n4852 DVDD.n4851 0.4505
R7374 DVDD.n5088 DVDD.n5087 0.4505
R7375 DVDD.n5086 DVDD.n4854 0.4505
R7376 DVDD.n5085 DVDD.n5084 0.4505
R7377 DVDD.n4856 DVDD.n4855 0.4505
R7378 DVDD.n5035 DVDD.n5034 0.4505
R7379 DVDD.n5036 DVDD.n5031 0.4505
R7380 DVDD.n5078 DVDD.n5077 0.4505
R7381 DVDD.n5076 DVDD.n5032 0.4505
R7382 DVDD.n5075 DVDD.n5074 0.4505
R7383 DVDD.n5038 DVDD.n5037 0.4505
R7384 DVDD.n5070 DVDD.n5069 0.4505
R7385 DVDD.n5068 DVDD.n5040 0.4505
R7386 DVDD.n5067 DVDD.n5066 0.4505
R7387 DVDD.n5042 DVDD.n5041 0.4505
R7388 DVDD.n5062 DVDD.n5061 0.4505
R7389 DVDD.n5060 DVDD.n5044 0.4505
R7390 DVDD.n5059 DVDD.n5058 0.4505
R7391 DVDD.n5046 DVDD.n5045 0.4505
R7392 DVDD.n5054 DVDD.n5053 0.4505
R7393 DVDD.n5052 DVDD.n5048 0.4505
R7394 DVDD.n5051 DVDD.n5050 0.4505
R7395 DVDD.n561 DVDD.n558 0.4505
R7396 DVDD.n8970 DVDD.n8969 0.4505
R7397 DVDD.n8968 DVDD.n560 0.4505
R7398 DVDD.n8967 DVDD.n8966 0.4505
R7399 DVDD.n8964 DVDD.n562 0.4505
R7400 DVDD.n566 DVDD.n563 0.4505
R7401 DVDD.n8960 DVDD.n8959 0.4505
R7402 DVDD.n8958 DVDD.n565 0.4505
R7403 DVDD.n8957 DVDD.n8956 0.4505
R7404 DVDD.n568 DVDD.n567 0.4505
R7405 DVDD.n8952 DVDD.n8951 0.4505
R7406 DVDD.n8950 DVDD.n570 0.4505
R7407 DVDD.n8949 DVDD.n8948 0.4505
R7408 DVDD.n572 DVDD.n571 0.4505
R7409 DVDD.n8944 DVDD.n8943 0.4505
R7410 DVDD.n8942 DVDD.n574 0.4505
R7411 DVDD.n8941 DVDD.n8940 0.4505
R7412 DVDD.n576 DVDD.n575 0.4505
R7413 DVDD.n1766 DVDD.n1764 0.4505
R7414 DVDD.n8248 DVDD.n8247 0.4505
R7415 DVDD.n8246 DVDD.n1765 0.4505
R7416 DVDD.n8245 DVDD.n8244 0.4505
R7417 DVDD.n1768 DVDD.n1767 0.4505
R7418 DVDD.n8240 DVDD.n8239 0.4505
R7419 DVDD.n8238 DVDD.n1771 0.4505
R7420 DVDD.n8237 DVDD.n8236 0.4505
R7421 DVDD.n1773 DVDD.n1772 0.4505
R7422 DVDD.n8232 DVDD.n8231 0.4505
R7423 DVDD.n8230 DVDD.n1774 0.4505
R7424 DVDD.n8229 DVDD.n8228 0.4505
R7425 DVDD.n8227 DVDD.n1775 0.4505
R7426 DVDD.n8225 DVDD.n8223 0.4505
R7427 DVDD.n8222 DVDD.n1776 0.4505
R7428 DVDD.n8221 DVDD.n8220 0.4505
R7429 DVDD.n1778 DVDD.n1777 0.4505
R7430 DVDD.n8216 DVDD.n8215 0.4505
R7431 DVDD.n8214 DVDD.n1781 0.4505
R7432 DVDD.n8213 DVDD.n8212 0.4505
R7433 DVDD.n1783 DVDD.n1782 0.4505
R7434 DVDD.n8201 DVDD.n8200 0.4505
R7435 DVDD.n8203 DVDD.n8202 0.4505
R7436 DVDD.n7501 DVDD.n7500 0.4505
R7437 DVDD.n7499 DVDD.n7092 0.4505
R7438 DVDD.n7498 DVDD.n7497 0.4505
R7439 DVDD.n7094 DVDD.n7093 0.4505
R7440 DVDD.n7493 DVDD.n7492 0.4505
R7441 DVDD.n7491 DVDD.n7096 0.4505
R7442 DVDD.n7490 DVDD.n7489 0.4505
R7443 DVDD.n7098 DVDD.n7097 0.4505
R7444 DVDD.n7307 DVDD.n7305 0.4505
R7445 DVDD.n7483 DVDD.n7482 0.4505
R7446 DVDD.n7481 DVDD.n7306 0.4505
R7447 DVDD.n7480 DVDD.n7479 0.4505
R7448 DVDD.n7309 DVDD.n7308 0.4505
R7449 DVDD.n7475 DVDD.n7474 0.4505
R7450 DVDD.n7473 DVDD.n7312 0.4505
R7451 DVDD.n7472 DVDD.n7471 0.4505
R7452 DVDD.n7314 DVDD.n7313 0.4505
R7453 DVDD.n7467 DVDD.n7466 0.4505
R7454 DVDD.n7465 DVDD.n7315 0.4505
R7455 DVDD.n7464 DVDD.n7463 0.4505
R7456 DVDD.n7462 DVDD.n7316 0.4505
R7457 DVDD.n7461 DVDD.n7459 0.4505
R7458 DVDD.n7458 DVDD.n7317 0.4505
R7459 DVDD.n7457 DVDD.n7456 0.4505
R7460 DVDD.n7319 DVDD.n7318 0.4505
R7461 DVDD.n7452 DVDD.n7451 0.4505
R7462 DVDD.n7450 DVDD.n7322 0.4505
R7463 DVDD.n7449 DVDD.n7448 0.4505
R7464 DVDD.n7324 DVDD.n7323 0.4505
R7465 DVDD.n7444 DVDD.n7443 0.4505
R7466 DVDD.n7442 DVDD.n7326 0.4505
R7467 DVDD.n7441 DVDD.n7440 0.4505
R7468 DVDD.n7328 DVDD.n7327 0.4505
R7469 DVDD.n7436 DVDD.n7435 0.4505
R7470 DVDD.n7434 DVDD.n7330 0.4505
R7471 DVDD.n7433 DVDD.n7432 0.4505
R7472 DVDD.n7332 DVDD.n7331 0.4505
R7473 DVDD.n7376 DVDD.n7374 0.4505
R7474 DVDD.n7420 DVDD.n7419 0.4505
R7475 DVDD.n7418 DVDD.n7375 0.4505
R7476 DVDD.n7417 DVDD.n7416 0.4505
R7477 DVDD.n7378 DVDD.n7377 0.4505
R7478 DVDD.n7412 DVDD.n7411 0.4505
R7479 DVDD.n7410 DVDD.n7380 0.4505
R7480 DVDD.n7409 DVDD.n7408 0.4505
R7481 DVDD.n7382 DVDD.n7381 0.4505
R7482 DVDD.n7404 DVDD.n7403 0.4505
R7483 DVDD.n7402 DVDD.n7384 0.4505
R7484 DVDD.n7401 DVDD.n7400 0.4505
R7485 DVDD.n7386 DVDD.n7385 0.4505
R7486 DVDD.n7396 DVDD.n7395 0.4505
R7487 DVDD.n7394 DVDD.n7388 0.4505
R7488 DVDD.n7393 DVDD.n7392 0.4505
R7489 DVDD.n7390 DVDD.n7389 0.4505
R7490 DVDD.n1726 DVDD.n1723 0.4505
R7491 DVDD.n8282 DVDD.n8281 0.4505
R7492 DVDD.n8280 DVDD.n1725 0.4505
R7493 DVDD.n8279 DVDD.n8278 0.4505
R7494 DVDD.n1728 DVDD.n1727 0.4505
R7495 DVDD.n8274 DVDD.n8273 0.4505
R7496 DVDD.n8272 DVDD.n1730 0.4505
R7497 DVDD.n8271 DVDD.n8270 0.4505
R7498 DVDD.n1732 DVDD.n1731 0.4505
R7499 DVDD.n8266 DVDD.n8265 0.4505
R7500 DVDD.n8264 DVDD.n1734 0.4505
R7501 DVDD.n8263 DVDD.n8262 0.4505
R7502 DVDD.n1736 DVDD.n1735 0.4505
R7503 DVDD.n8258 DVDD.n8257 0.4505
R7504 DVDD.n8256 DVDD.n1738 0.4505
R7505 DVDD.n8255 DVDD.n8254 0.4505
R7506 DVDD.n1740 DVDD.n1739 0.4505
R7507 DVDD.n6232 DVDD.n3885 0.4505
R7508 DVDD.n6443 DVDD.n6442 0.4505
R7509 DVDD.n6441 DVDD.n3473 0.4505
R7510 DVDD.n6440 DVDD.n3468 0.4505
R7511 DVDD.n6434 DVDD.n3503 0.4505
R7512 DVDD.n6436 DVDD.n6435 0.4505
R7513 DVDD.n6433 DVDD.n3505 0.4505
R7514 DVDD.n6432 DVDD.n6431 0.4505
R7515 DVDD.n3507 DVDD.n3506 0.4505
R7516 DVDD.n6427 DVDD.n6426 0.4505
R7517 DVDD.n6425 DVDD.n1102 0.4505
R7518 DVDD.n6214 DVDD.n3509 0.4505
R7519 DVDD.n6215 DVDD.n6213 0.4505
R7520 DVDD.n6217 DVDD.n6216 0.4505
R7521 DVDD.n3892 DVDD.n3891 0.4505
R7522 DVDD.n6222 DVDD.n6221 0.4505
R7523 DVDD.n6223 DVDD.n3889 0.4505
R7524 DVDD.n6225 DVDD.n6224 0.4505
R7525 DVDD.n3890 DVDD.n3886 0.4505
R7526 DVDD.n6229 DVDD.n3887 0.4505
R7527 DVDD.n6231 DVDD.n6230 0.4505
R7528 DVDD.n6233 DVDD.n6232 0.4505
R7529 DVDD.n6231 DVDD.n3883 0.4505
R7530 DVDD.n6229 DVDD.n6228 0.4505
R7531 DVDD.n6227 DVDD.n3886 0.4505
R7532 DVDD.n6226 DVDD.n6225 0.4505
R7533 DVDD.n3889 DVDD.n3888 0.4505
R7534 DVDD.n6221 DVDD.n6220 0.4505
R7535 DVDD.n6219 DVDD.n3892 0.4505
R7536 DVDD.n6218 DVDD.n6217 0.4505
R7537 DVDD.n6213 DVDD.n6212 0.4505
R7538 DVDD.n6211 DVDD.n3509 0.4505
R7539 DVDD.n6425 DVDD.n3508 0.4505
R7540 DVDD.n6428 DVDD.n6427 0.4505
R7541 DVDD.n6429 DVDD.n3507 0.4505
R7542 DVDD.n6431 DVDD.n6430 0.4505
R7543 DVDD.n3505 DVDD.n3504 0.4505
R7544 DVDD.n6437 DVDD.n6436 0.4505
R7545 DVDD.n6438 DVDD.n3503 0.4505
R7546 DVDD.n6440 DVDD.n6439 0.4505
R7547 DVDD.n6441 DVDD.n3502 0.4505
R7548 DVDD.n6444 DVDD.n6443 0.4505
R7549 DVDD.n6080 DVDD.n6079 0.4505
R7550 DVDD.n6078 DVDD.n5911 0.4505
R7551 DVDD.n6077 DVDD.n6076 0.4505
R7552 DVDD.n5914 DVDD.n5913 0.4505
R7553 DVDD.n6072 DVDD.n6071 0.4505
R7554 DVDD.n6070 DVDD.n5916 0.4505
R7555 DVDD.n6069 DVDD.n6068 0.4505
R7556 DVDD.n5921 DVDD.n5918 0.4505
R7557 DVDD.n6064 DVDD.n6063 0.4505
R7558 DVDD.n5928 DVDD.n5920 0.4505
R7559 DVDD.n5995 DVDD.n5994 0.4505
R7560 DVDD.n3942 DVDD.n3941 0.4505
R7561 DVDD.n3940 DVDD.n3916 0.4505
R7562 DVDD.n3939 DVDD.n3938 0.4505
R7563 DVDD.n3918 DVDD.n3917 0.4505
R7564 DVDD.n3934 DVDD.n3933 0.4505
R7565 DVDD.n3932 DVDD.n3920 0.4505
R7566 DVDD.n3931 DVDD.n3930 0.4505
R7567 DVDD.n3922 DVDD.n3921 0.4505
R7568 DVDD.n3926 DVDD.n3925 0.4505
R7569 DVDD.n3924 DVDD.n3923 0.4505
R7570 DVDD.n6081 DVDD.n6080 0.4505
R7571 DVDD.n5911 DVDD.n5909 0.4505
R7572 DVDD.n6076 DVDD.n6075 0.4505
R7573 DVDD.n6074 DVDD.n5914 0.4505
R7574 DVDD.n6073 DVDD.n6072 0.4505
R7575 DVDD.n5916 DVDD.n5915 0.4505
R7576 DVDD.n6068 DVDD.n6067 0.4505
R7577 DVDD.n6066 DVDD.n5918 0.4505
R7578 DVDD.n6065 DVDD.n6064 0.4505
R7579 DVDD.n5920 DVDD.n5919 0.4505
R7580 DVDD.n5994 DVDD.n3914 0.4505
R7581 DVDD.n3943 DVDD.n3942 0.4505
R7582 DVDD.n3916 DVDD.n3915 0.4505
R7583 DVDD.n3938 DVDD.n3937 0.4505
R7584 DVDD.n3936 DVDD.n3918 0.4505
R7585 DVDD.n3935 DVDD.n3934 0.4505
R7586 DVDD.n3920 DVDD.n3919 0.4505
R7587 DVDD.n3930 DVDD.n3929 0.4505
R7588 DVDD.n3928 DVDD.n3922 0.4505
R7589 DVDD.n3927 DVDD.n3926 0.4505
R7590 DVDD.n3923 DVDD.n3882 0.4505
R7591 DVDD.n4405 DVDD.n4404 0.4505
R7592 DVDD.n4408 DVDD.n4407 0.4505
R7593 DVDD.n4409 DVDD.n4403 0.4505
R7594 DVDD.n4411 DVDD.n4410 0.4505
R7595 DVDD.n4401 DVDD.n4400 0.4505
R7596 DVDD.n4416 DVDD.n4415 0.4505
R7597 DVDD.n4417 DVDD.n4399 0.4505
R7598 DVDD.n4420 DVDD.n4419 0.4505
R7599 DVDD.n4418 DVDD.n4397 0.4505
R7600 DVDD.n4424 DVDD.n4396 0.4505
R7601 DVDD.n4426 DVDD.n4425 0.4505
R7602 DVDD.n6099 DVDD.n6098 0.4505
R7603 DVDD.n5765 DVDD.n4395 0.4505
R7604 DVDD.n5900 DVDD.n5899 0.4505
R7605 DVDD.n5897 DVDD.n5892 0.4505
R7606 DVDD.n6094 DVDD.n6093 0.4505
R7607 DVDD.n5898 DVDD.n5896 0.4505
R7608 DVDD.n6089 DVDD.n6088 0.4505
R7609 DVDD.n6087 DVDD.n5904 0.4505
R7610 DVDD.n6086 DVDD.n6085 0.4505
R7611 DVDD.n5906 DVDD.n5905 0.4505
R7612 DVDD.n4405 DVDD.n2787 0.4505
R7613 DVDD.n4407 DVDD.n4406 0.4505
R7614 DVDD.n4403 DVDD.n4402 0.4505
R7615 DVDD.n4412 DVDD.n4411 0.4505
R7616 DVDD.n4413 DVDD.n4401 0.4505
R7617 DVDD.n4415 DVDD.n4414 0.4505
R7618 DVDD.n4399 DVDD.n4398 0.4505
R7619 DVDD.n4421 DVDD.n4420 0.4505
R7620 DVDD.n4422 DVDD.n4397 0.4505
R7621 DVDD.n4424 DVDD.n4423 0.4505
R7622 DVDD.n4425 DVDD.n4392 0.4505
R7623 DVDD.n6100 DVDD.n6099 0.4505
R7624 DVDD.n4395 DVDD.n4393 0.4505
R7625 DVDD.n5901 DVDD.n5900 0.4505
R7626 DVDD.n5902 DVDD.n5897 0.4505
R7627 DVDD.n6093 DVDD.n6092 0.4505
R7628 DVDD.n6091 DVDD.n5898 0.4505
R7629 DVDD.n6090 DVDD.n6089 0.4505
R7630 DVDD.n5904 DVDD.n5903 0.4505
R7631 DVDD.n6085 DVDD.n6084 0.4505
R7632 DVDD.n6083 DVDD.n5906 0.4505
R7633 DVDD.n5649 DVDD.n5648 0.4505
R7634 DVDD.n4458 DVDD.n4457 0.4505
R7635 DVDD.n5662 DVDD.n5661 0.4505
R7636 DVDD.n5663 DVDD.n4456 0.4505
R7637 DVDD.n5666 DVDD.n5665 0.4505
R7638 DVDD.n5664 DVDD.n4453 0.4505
R7639 DVDD.n5670 DVDD.n4454 0.4505
R7640 DVDD.n5671 DVDD.n4452 0.4505
R7641 DVDD.n5673 DVDD.n5672 0.4505
R7642 DVDD.n5674 DVDD.n4451 0.4505
R7643 DVDD.n5679 DVDD.n5675 0.4505
R7644 DVDD.n5708 DVDD.n5681 0.4505
R7645 DVDD.n5684 DVDD.n5680 0.4505
R7646 DVDD.n5704 DVDD.n5703 0.4505
R7647 DVDD.n5702 DVDD.n5683 0.4505
R7648 DVDD.n5701 DVDD.n5700 0.4505
R7649 DVDD.n5686 DVDD.n5685 0.4505
R7650 DVDD.n5696 DVDD.n5695 0.4505
R7651 DVDD.n5694 DVDD.n5688 0.4505
R7652 DVDD.n5693 DVDD.n5692 0.4505
R7653 DVDD.n5690 DVDD.n2788 0.4505
R7654 DVDD.n5650 DVDD.n5649 0.4505
R7655 DVDD.n5482 DVDD.n4458 0.4505
R7656 DVDD.n5661 DVDD.n5660 0.4505
R7657 DVDD.n4456 DVDD.n4455 0.4505
R7658 DVDD.n5667 DVDD.n5666 0.4505
R7659 DVDD.n5668 DVDD.n4453 0.4505
R7660 DVDD.n5670 DVDD.n5669 0.4505
R7661 DVDD.n5671 DVDD.n3002 0.4505
R7662 DVDD.n5672 DVDD.n3008 0.4505
R7663 DVDD.n4451 DVDD.n4450 0.4505
R7664 DVDD.n5679 DVDD.n5678 0.4505
R7665 DVDD.n5708 DVDD.n5707 0.4505
R7666 DVDD.n5706 DVDD.n5680 0.4505
R7667 DVDD.n5705 DVDD.n5704 0.4505
R7668 DVDD.n5683 DVDD.n5682 0.4505
R7669 DVDD.n5700 DVDD.n5699 0.4505
R7670 DVDD.n5698 DVDD.n5686 0.4505
R7671 DVDD.n5697 DVDD.n5696 0.4505
R7672 DVDD.n5688 DVDD.n5687 0.4505
R7673 DVDD.n5692 DVDD.n5691 0.4505
R7674 DVDD.n5690 DVDD.n5689 0.4505
R7675 DVDD.n7684 DVDD.n2370 0.4505
R7676 DVDD.n7737 DVDD.n7736 0.4505
R7677 DVDD.n7696 DVDD.n7695 0.4505
R7678 DVDD.n7723 DVDD.n7720 0.4505
R7679 DVDD.n8200 DVDD.n1797 0.4505
R7680 DVDD.n1790 DVDD.n1783 0.4505
R7681 DVDD.n8212 DVDD.n8211 0.4505
R7682 DVDD.n1781 DVDD.n1780 0.4505
R7683 DVDD.n8217 DVDD.n8216 0.4505
R7684 DVDD.n8218 DVDD.n1778 0.4505
R7685 DVDD.n8220 DVDD.n8219 0.4505
R7686 DVDD.n1779 DVDD.n1776 0.4505
R7687 DVDD.n8225 DVDD.n8224 0.4505
R7688 DVDD.n8227 DVDD.n8226 0.4505
R7689 DVDD.n8228 DVDD.n1280 0.4505
R7690 DVDD.n1774 DVDD.n1274 0.4505
R7691 DVDD.n8233 DVDD.n8232 0.4505
R7692 DVDD.n8234 DVDD.n1773 0.4505
R7693 DVDD.n8236 DVDD.n8235 0.4505
R7694 DVDD.n1771 DVDD.n1770 0.4505
R7695 DVDD.n8241 DVDD.n8240 0.4505
R7696 DVDD.n8242 DVDD.n1768 0.4505
R7697 DVDD.n8244 DVDD.n8243 0.4505
R7698 DVDD.n1769 DVDD.n1765 0.4505
R7699 DVDD.n8249 DVDD.n8248 0.4505
R7700 DVDD.n1764 DVDD.n1758 0.4505
R7701 DVDD.n7090 DVDD.n7076 0.4505
R7702 DVDD.n7502 DVDD.n7501 0.4505
R7703 DVDD.n7092 DVDD.n7091 0.4505
R7704 DVDD.n7497 DVDD.n7496 0.4505
R7705 DVDD.n7495 DVDD.n7094 0.4505
R7706 DVDD.n7494 DVDD.n7493 0.4505
R7707 DVDD.n7096 DVDD.n7095 0.4505
R7708 DVDD.n7489 DVDD.n7488 0.4505
R7709 DVDD.n7104 DVDD.n7098 0.4505
R7710 DVDD.n7305 DVDD.n7299 0.4505
R7711 DVDD.n7484 DVDD.n7483 0.4505
R7712 DVDD.n7310 DVDD.n7306 0.4505
R7713 DVDD.n7479 DVDD.n7478 0.4505
R7714 DVDD.n7477 DVDD.n7309 0.4505
R7715 DVDD.n7476 DVDD.n7475 0.4505
R7716 DVDD.n7312 DVDD.n7311 0.4505
R7717 DVDD.n7471 DVDD.n7470 0.4505
R7718 DVDD.n7469 DVDD.n7314 0.4505
R7719 DVDD.n7468 DVDD.n7467 0.4505
R7720 DVDD.n7315 DVDD.n1514 0.4505
R7721 DVDD.n7463 DVDD.n1520 0.4505
R7722 DVDD.n7462 DVDD.n1527 0.4505
R7723 DVDD.n7461 DVDD.n7460 0.4505
R7724 DVDD.n7320 DVDD.n7317 0.4505
R7725 DVDD.n7456 DVDD.n7455 0.4505
R7726 DVDD.n7454 DVDD.n7319 0.4505
R7727 DVDD.n7453 DVDD.n7452 0.4505
R7728 DVDD.n7322 DVDD.n7321 0.4505
R7729 DVDD.n7448 DVDD.n7447 0.4505
R7730 DVDD.n7446 DVDD.n7324 0.4505
R7731 DVDD.n7445 DVDD.n7444 0.4505
R7732 DVDD.n7326 DVDD.n7325 0.4505
R7733 DVDD.n7440 DVDD.n7439 0.4505
R7734 DVDD.n7438 DVDD.n7328 0.4505
R7735 DVDD.n7437 DVDD.n7436 0.4505
R7736 DVDD.n7330 DVDD.n7329 0.4505
R7737 DVDD.n7432 DVDD.n7431 0.4505
R7738 DVDD.n7339 DVDD.n7332 0.4505
R7739 DVDD.n7374 DVDD.n7369 0.4505
R7740 DVDD.n7421 DVDD.n7420 0.4505
R7741 DVDD.n7375 DVDD.n7373 0.4505
R7742 DVDD.n7416 DVDD.n7415 0.4505
R7743 DVDD.n7414 DVDD.n7378 0.4505
R7744 DVDD.n7413 DVDD.n7412 0.4505
R7745 DVDD.n7380 DVDD.n7379 0.4505
R7746 DVDD.n7408 DVDD.n7407 0.4505
R7747 DVDD.n7406 DVDD.n7382 0.4505
R7748 DVDD.n7405 DVDD.n7404 0.4505
R7749 DVDD.n7384 DVDD.n7383 0.4505
R7750 DVDD.n7400 DVDD.n7399 0.4505
R7751 DVDD.n7398 DVDD.n7386 0.4505
R7752 DVDD.n7397 DVDD.n7396 0.4505
R7753 DVDD.n7388 DVDD.n7387 0.4505
R7754 DVDD.n7392 DVDD.n7391 0.4505
R7755 DVDD.n7390 DVDD.n1705 0.4505
R7756 DVDD.n1723 DVDD.n1712 0.4505
R7757 DVDD.n8283 DVDD.n8282 0.4505
R7758 DVDD.n1725 DVDD.n1724 0.4505
R7759 DVDD.n8278 DVDD.n8277 0.4505
R7760 DVDD.n8276 DVDD.n1728 0.4505
R7761 DVDD.n8275 DVDD.n8274 0.4505
R7762 DVDD.n1730 DVDD.n1729 0.4505
R7763 DVDD.n8270 DVDD.n8269 0.4505
R7764 DVDD.n8268 DVDD.n1732 0.4505
R7765 DVDD.n8267 DVDD.n8266 0.4505
R7766 DVDD.n1734 DVDD.n1733 0.4505
R7767 DVDD.n8262 DVDD.n8261 0.4505
R7768 DVDD.n8260 DVDD.n1736 0.4505
R7769 DVDD.n8259 DVDD.n8258 0.4505
R7770 DVDD.n1738 DVDD.n1737 0.4505
R7771 DVDD.n8254 DVDD.n8253 0.4505
R7772 DVDD.n1746 DVDD.n1740 0.4505
R7773 DVDD.n648 DVDD.n640 0.4505
R7774 DVDD.n8896 DVDD.n8895 0.4505
R7775 DVDD.n641 DVDD.n638 0.4505
R7776 DVDD.n8901 DVDD.n8900 0.4505
R7777 DVDD.n8902 DVDD.n636 0.4505
R7778 DVDD.n8904 DVDD.n8903 0.4505
R7779 DVDD.n634 DVDD.n633 0.4505
R7780 DVDD.n8909 DVDD.n8908 0.4505
R7781 DVDD.n617 DVDD.n609 0.4505
R7782 DVDD.n8914 DVDD.n8913 0.4505
R7783 DVDD.n610 DVDD.n607 0.4505
R7784 DVDD.n8919 DVDD.n8918 0.4505
R7785 DVDD.n8920 DVDD.n605 0.4505
R7786 DVDD.n8922 DVDD.n8921 0.4505
R7787 DVDD.n603 DVDD.n602 0.4505
R7788 DVDD.n8927 DVDD.n8926 0.4505
R7789 DVDD.n8928 DVDD.n601 0.4505
R7790 DVDD.n8930 DVDD.n8929 0.4505
R7791 DVDD.n595 DVDD.n593 0.4505
R7792 DVDD.n8935 DVDD.n8934 0.4505
R7793 DVDD.n594 DVDD.n592 0.4505
R7794 DVDD.n597 DVDD.n596 0.4505
R7795 DVDD.n4709 DVDD.n4708 0.4505
R7796 DVDD.n4710 DVDD.n4612 0.4505
R7797 DVDD.n4715 DVDD.n4714 0.4505
R7798 DVDD.n4610 DVDD.n4609 0.4505
R7799 DVDD.n4720 DVDD.n4719 0.4505
R7800 DVDD.n4721 DVDD.n4608 0.4505
R7801 DVDD.n4723 DVDD.n4722 0.4505
R7802 DVDD.n4606 DVDD.n4600 0.4505
R7803 DVDD.n4728 DVDD.n4727 0.4505
R7804 DVDD.n4737 DVDD.n4592 0.4505
R7805 DVDD.n4823 DVDD.n4822 0.4505
R7806 DVDD.n4590 DVDD.n4589 0.4505
R7807 DVDD.n4828 DVDD.n4827 0.4505
R7808 DVDD.n4829 DVDD.n4588 0.4505
R7809 DVDD.n4831 DVDD.n4830 0.4505
R7810 DVDD.n4586 DVDD.n4585 0.4505
R7811 DVDD.n4836 DVDD.n4835 0.4505
R7812 DVDD.n4837 DVDD.n4584 0.4505
R7813 DVDD.n4839 DVDD.n4838 0.4505
R7814 DVDD.n4580 DVDD.n4574 0.4505
R7815 DVDD.n5115 DVDD.n5114 0.4505
R7816 DVDD.n4582 DVDD.n4581 0.4505
R7817 DVDD.n5110 DVDD.n5109 0.4505
R7818 DVDD.n5108 DVDD.n5107 0.4505
R7819 DVDD.n5106 DVDD.n4843 0.4505
R7820 DVDD.n5105 DVDD.n5104 0.4505
R7821 DVDD.n4845 DVDD.n4844 0.4505
R7822 DVDD.n5100 DVDD.n5099 0.4505
R7823 DVDD.n5098 DVDD.n4848 0.4505
R7824 DVDD.n5097 DVDD.n5096 0.4505
R7825 DVDD.n4850 DVDD.n4849 0.4505
R7826 DVDD.n5092 DVDD.n5091 0.4505
R7827 DVDD.n5090 DVDD.n4852 0.4505
R7828 DVDD.n5089 DVDD.n5088 0.4505
R7829 DVDD.n4854 DVDD.n4853 0.4505
R7830 DVDD.n5084 DVDD.n5083 0.4505
R7831 DVDD.n4862 DVDD.n4856 0.4505
R7832 DVDD.n5034 DVDD.n5033 0.4505
R7833 DVDD.n5031 DVDD.n5029 0.4505
R7834 DVDD.n5079 DVDD.n5078 0.4505
R7835 DVDD.n5032 DVDD.n5030 0.4505
R7836 DVDD.n5074 DVDD.n5073 0.4505
R7837 DVDD.n5072 DVDD.n5038 0.4505
R7838 DVDD.n5071 DVDD.n5070 0.4505
R7839 DVDD.n5040 DVDD.n5039 0.4505
R7840 DVDD.n5066 DVDD.n5065 0.4505
R7841 DVDD.n5064 DVDD.n5042 0.4505
R7842 DVDD.n5063 DVDD.n5062 0.4505
R7843 DVDD.n5044 DVDD.n5043 0.4505
R7844 DVDD.n5058 DVDD.n5057 0.4505
R7845 DVDD.n5056 DVDD.n5046 0.4505
R7846 DVDD.n5055 DVDD.n5054 0.4505
R7847 DVDD.n5048 DVDD.n5047 0.4505
R7848 DVDD.n5050 DVDD.n5049 0.4505
R7849 DVDD.n558 DVDD.n552 0.4505
R7850 DVDD.n8971 DVDD.n8970 0.4505
R7851 DVDD.n560 DVDD.n559 0.4505
R7852 DVDD.n8966 DVDD.n8965 0.4505
R7853 DVDD.n8964 DVDD.n8963 0.4505
R7854 DVDD.n8962 DVDD.n563 0.4505
R7855 DVDD.n8961 DVDD.n8960 0.4505
R7856 DVDD.n565 DVDD.n564 0.4505
R7857 DVDD.n8956 DVDD.n8955 0.4505
R7858 DVDD.n8954 DVDD.n568 0.4505
R7859 DVDD.n8953 DVDD.n8952 0.4505
R7860 DVDD.n570 DVDD.n569 0.4505
R7861 DVDD.n8948 DVDD.n8947 0.4505
R7862 DVDD.n8946 DVDD.n572 0.4505
R7863 DVDD.n8945 DVDD.n8944 0.4505
R7864 DVDD.n574 DVDD.n573 0.4505
R7865 DVDD.n8940 DVDD.n8939 0.4505
R7866 DVDD.n582 DVDD.n576 0.4505
R7867 DVDD.n9695 DVDD.n9694 0.4505
R7868 DVDD.n9696 DVDD.n0 0.4505
R7869 DVDD.n3 DVDD.n2 0.4505
R7870 DVDD.n9690 DVDD.n9689 0.4505
R7871 DVDD.n17 DVDD.n16 0.4505
R7872 DVDD.n9684 DVDD.n9683 0.4505
R7873 DVDD.n9682 DVDD.n19 0.4505
R7874 DVDD.n9681 DVDD.n9680 0.4505
R7875 DVDD.n30 DVDD.n21 0.4505
R7876 DVDD.n9676 DVDD.n9675 0.4505
R7877 DVDD.n9671 DVDD.n23 0.4505
R7878 DVDD.n9670 DVDD.n9669 0.4505
R7879 DVDD.n48 DVDD.n47 0.4505
R7880 DVDD.n9665 DVDD.n9664 0.4505
R7881 DVDD.n9663 DVDD.n50 0.4505
R7882 DVDD.n9662 DVDD.n9661 0.4505
R7883 DVDD.n52 DVDD.n51 0.4505
R7884 DVDD.n9657 DVDD.n9656 0.4505
R7885 DVDD.n9655 DVDD.n54 0.4505
R7886 DVDD.n9654 DVDD.n9653 0.4505
R7887 DVDD.n65 DVDD.n56 0.4505
R7888 DVDD.n9649 DVDD.n9648 0.4505
R7889 DVDD.n4756 DVDD.n4551 0.4505
R7890 DVDD.n4758 DVDD.n4757 0.4505
R7891 DVDD.n4762 DVDD.n4759 0.4505
R7892 DVDD.n4764 DVDD.n4763 0.4505
R7893 DVDD.n4766 DVDD.n4765 0.4505
R7894 DVDD.n4754 DVDD.n4753 0.4505
R7895 DVDD.n4772 DVDD.n4771 0.4505
R7896 DVDD.n4773 DVDD.n4752 0.4505
R7897 DVDD.n4789 DVDD.n4788 0.4505
R7898 DVDD.n4791 DVDD.n4790 0.4505
R7899 DVDD.n4749 DVDD.n4742 0.4505
R7900 DVDD.n4815 DVDD.n4814 0.4505
R7901 DVDD.n4750 DVDD.n4748 0.4505
R7902 DVDD.n4810 DVDD.n4809 0.4505
R7903 DVDD.n4808 DVDD.n4795 0.4505
R7904 DVDD.n4807 DVDD.n4806 0.4505
R7905 DVDD.n4797 DVDD.n4796 0.4505
R7906 DVDD.n4802 DVDD.n4801 0.4505
R7907 DVDD.n4800 DVDD.n4799 0.4505
R7908 DVDD.n465 DVDD.n460 0.4505
R7909 DVDD.n9243 DVDD.n9242 0.4505
R7910 DVDD.n467 DVDD.n466 0.4505
R7911 DVDD.n9238 DVDD.n9237 0.4505
R7912 DVDD.n9236 DVDD.n9235 0.4505
R7913 DVDD.n9234 DVDD.n470 0.4505
R7914 DVDD.n9233 DVDD.n9232 0.4505
R7915 DVDD.n472 DVDD.n471 0.4505
R7916 DVDD.n9228 DVDD.n9227 0.4505
R7917 DVDD.n9226 DVDD.n475 0.4505
R7918 DVDD.n9225 DVDD.n9224 0.4505
R7919 DVDD.n477 DVDD.n476 0.4505
R7920 DVDD.n9220 DVDD.n9219 0.4505
R7921 DVDD.n9218 DVDD.n479 0.4505
R7922 DVDD.n9217 DVDD.n9216 0.4505
R7923 DVDD.n481 DVDD.n480 0.4505
R7924 DVDD.n9212 DVDD.n9211 0.4505
R7925 DVDD.n489 DVDD.n483 0.4505
R7926 DVDD.n504 DVDD.n503 0.4505
R7927 DVDD.n501 DVDD.n499 0.4505
R7928 DVDD.n9207 DVDD.n9206 0.4505
R7929 DVDD.n502 DVDD.n500 0.4505
R7930 DVDD.n9202 DVDD.n9201 0.4505
R7931 DVDD.n9200 DVDD.n508 0.4505
R7932 DVDD.n9199 DVDD.n9198 0.4505
R7933 DVDD.n510 DVDD.n509 0.4505
R7934 DVDD.n9194 DVDD.n9193 0.4505
R7935 DVDD.n9192 DVDD.n512 0.4505
R7936 DVDD.n9191 DVDD.n9190 0.4505
R7937 DVDD.n514 DVDD.n513 0.4505
R7938 DVDD.n9186 DVDD.n9185 0.4505
R7939 DVDD.n9184 DVDD.n516 0.4505
R7940 DVDD.n9183 DVDD.n9182 0.4505
R7941 DVDD.n518 DVDD.n517 0.4505
R7942 DVDD.n9178 DVDD.n9177 0.4505
R7943 DVDD.n9176 DVDD.n520 0.4505
R7944 DVDD.n9129 DVDD.n526 0.4505
R7945 DVDD.n9127 DVDD.n9126 0.4505
R7946 DVDD.n9172 DVDD.n9171 0.4505
R7947 DVDD.n9134 DVDD.n9128 0.4505
R7948 DVDD.n9167 DVDD.n9166 0.4505
R7949 DVDD.n9165 DVDD.n9133 0.4505
R7950 DVDD.n9164 DVDD.n9163 0.4505
R7951 DVDD.n9136 DVDD.n9135 0.4505
R7952 DVDD.n9159 DVDD.n9158 0.4505
R7953 DVDD.n9157 DVDD.n9138 0.4505
R7954 DVDD.n9156 DVDD.n9155 0.4505
R7955 DVDD.n9140 DVDD.n9139 0.4505
R7956 DVDD.n9151 DVDD.n9150 0.4505
R7957 DVDD.n9149 DVDD.n9142 0.4505
R7958 DVDD.n9148 DVDD.n9147 0.4505
R7959 DVDD.n9144 DVDD.n9143 0.4505
R7960 DVDD.n9650 DVDD.n9649 0.4505
R7961 DVDD.n9651 DVDD.n56 0.4505
R7962 DVDD.n9653 DVDD.n9652 0.4505
R7963 DVDD.n54 DVDD.n53 0.4505
R7964 DVDD.n9658 DVDD.n9657 0.4505
R7965 DVDD.n9659 DVDD.n52 0.4505
R7966 DVDD.n9661 DVDD.n9660 0.4505
R7967 DVDD.n50 DVDD.n49 0.4505
R7968 DVDD.n9666 DVDD.n9665 0.4505
R7969 DVDD.n9667 DVDD.n48 0.4505
R7970 DVDD.n9669 DVDD.n9668 0.4505
R7971 DVDD.n23 DVDD.n22 0.4505
R7972 DVDD.n9677 DVDD.n9676 0.4505
R7973 DVDD.n9678 DVDD.n21 0.4505
R7974 DVDD.n9680 DVDD.n9679 0.4505
R7975 DVDD.n19 DVDD.n18 0.4505
R7976 DVDD.n9685 DVDD.n9684 0.4505
R7977 DVDD.n9686 DVDD.n17 0.4505
R7978 DVDD.n9689 DVDD.n9688 0.4505
R7979 DVDD.n9687 DVDD.n2 0.4505
R7980 DVDD.n9695 DVDD.n1 0.4505
R7981 DVDD.n9697 DVDD.n9696 0.4505
R7982 DVDD.n9699 DVDD.n9698 0.4505
R7983 DVDD.n4760 DVDD.n4758 0.4505
R7984 DVDD.n4762 DVDD.n4761 0.4505
R7985 DVDD.n4763 DVDD.n4755 0.4505
R7986 DVDD.n4767 DVDD.n4766 0.4505
R7987 DVDD.n4768 DVDD.n4754 0.4505
R7988 DVDD.n4771 DVDD.n4770 0.4505
R7989 DVDD.n4769 DVDD.n4752 0.4505
R7990 DVDD.n4789 DVDD.n4751 0.4505
R7991 DVDD.n4792 DVDD.n4791 0.4505
R7992 DVDD.n4793 DVDD.n4749 0.4505
R7993 DVDD.n4814 DVDD.n4813 0.4505
R7994 DVDD.n4812 DVDD.n4750 0.4505
R7995 DVDD.n4811 DVDD.n4810 0.4505
R7996 DVDD.n4795 DVDD.n4794 0.4505
R7997 DVDD.n4806 DVDD.n4805 0.4505
R7998 DVDD.n4804 DVDD.n4797 0.4505
R7999 DVDD.n4803 DVDD.n4802 0.4505
R8000 DVDD.n4799 DVDD.n4798 0.4505
R8001 DVDD.n468 DVDD.n465 0.4505
R8002 DVDD.n9242 DVDD.n9241 0.4505
R8003 DVDD.n9240 DVDD.n467 0.4505
R8004 DVDD.n9239 DVDD.n9238 0.4505
R8005 DVDD.n9236 DVDD.n469 0.4505
R8006 DVDD.n473 DVDD.n470 0.4505
R8007 DVDD.n9232 DVDD.n9231 0.4505
R8008 DVDD.n9230 DVDD.n472 0.4505
R8009 DVDD.n9229 DVDD.n9228 0.4505
R8010 DVDD.n475 DVDD.n474 0.4505
R8011 DVDD.n9224 DVDD.n9223 0.4505
R8012 DVDD.n9222 DVDD.n477 0.4505
R8013 DVDD.n9221 DVDD.n9220 0.4505
R8014 DVDD.n479 DVDD.n478 0.4505
R8015 DVDD.n9216 DVDD.n9215 0.4505
R8016 DVDD.n9214 DVDD.n481 0.4505
R8017 DVDD.n9213 DVDD.n9212 0.4505
R8018 DVDD.n483 DVDD.n482 0.4505
R8019 DVDD.n505 DVDD.n504 0.4505
R8020 DVDD.n506 DVDD.n501 0.4505
R8021 DVDD.n9206 DVDD.n9205 0.4505
R8022 DVDD.n9204 DVDD.n502 0.4505
R8023 DVDD.n9203 DVDD.n9202 0.4505
R8024 DVDD.n508 DVDD.n507 0.4505
R8025 DVDD.n9198 DVDD.n9197 0.4505
R8026 DVDD.n9196 DVDD.n510 0.4505
R8027 DVDD.n9195 DVDD.n9194 0.4505
R8028 DVDD.n512 DVDD.n511 0.4505
R8029 DVDD.n9190 DVDD.n9189 0.4505
R8030 DVDD.n9188 DVDD.n514 0.4505
R8031 DVDD.n9187 DVDD.n9186 0.4505
R8032 DVDD.n516 DVDD.n515 0.4505
R8033 DVDD.n9182 DVDD.n9181 0.4505
R8034 DVDD.n9180 DVDD.n518 0.4505
R8035 DVDD.n9179 DVDD.n9178 0.4505
R8036 DVDD.n520 DVDD.n519 0.4505
R8037 DVDD.n9130 DVDD.n9129 0.4505
R8038 DVDD.n9131 DVDD.n9127 0.4505
R8039 DVDD.n9171 DVDD.n9170 0.4505
R8040 DVDD.n9169 DVDD.n9128 0.4505
R8041 DVDD.n9168 DVDD.n9167 0.4505
R8042 DVDD.n9133 DVDD.n9132 0.4505
R8043 DVDD.n9163 DVDD.n9162 0.4505
R8044 DVDD.n9161 DVDD.n9136 0.4505
R8045 DVDD.n9160 DVDD.n9159 0.4505
R8046 DVDD.n9138 DVDD.n9137 0.4505
R8047 DVDD.n9155 DVDD.n9154 0.4505
R8048 DVDD.n9153 DVDD.n9140 0.4505
R8049 DVDD.n9152 DVDD.n9151 0.4505
R8050 DVDD.n9142 DVDD.n9141 0.4505
R8051 DVDD.n9147 DVDD.n9146 0.4505
R8052 DVDD.n9145 DVDD.n9144 0.4505
R8053 DVDD.n58 DVDD.n57 0.4505
R8054 DVDD.n72 DVDD.n58 0.4505
R8055 DVDD.n8421 DVDD.n8420 0.440926
R8056 DVDD.n8438 DVDD.n8435 0.440926
R8057 DVDD.n8507 DVDD.n1415 0.440926
R8058 DVDD.n8498 DVDD.n8497 0.440926
R8059 DVDD.n8513 DVDD.n1409 0.440926
R8060 DVDD.n8597 DVDD.n8596 0.440926
R8061 DVDD.n8632 DVDD.n1317 0.399122
R8062 DVDD.n8637 DVDD.n1309 0.399122
R8063 DVDD.n7429 DVDD.n7363 0.399122
R8064 DVDD.n8371 DVDD.n8370 0.399122
R8065 DVDD.n8647 DVDD.n8646 0.399122
R8066 DVDD.n7486 DVDD.n1502 0.399122
R8067 DVDD.n3500 DVDD.n3490 0.383973
R8068 DVDD.n6457 DVDD.n6456 0.383973
R8069 DVDD.n797 DVDD.n672 0.3821
R8070 DVDD.n8795 DVDD.n8794 0.3821
R8071 DVDD.n8877 DVDD.n8876 0.375556
R8072 DVDD.n3801 DVDD.n3752 0.374243
R8073 DVDD.n7189 DVDD.n7186 0.365885
R8074 DVDD.n7180 DVDD.n7177 0.365885
R8075 DVDD.n8376 DVDD.n1508 0.365885
R8076 DVDD.n8636 DVDD.n8633 0.365885
R8077 DVDD.n5912 DVDD.n5908 0.35585
R8078 DVDD.n228 DVDD.n223 0.355277
R8079 DVDD.n9616 DVDD.n111 0.355277
R8080 DVDD.n9425 DVDD.n187 0.35501
R8081 DVDD.n228 DVDD.n220 0.35405
R8082 DVDD.n5912 DVDD.n5907 0.353477
R8083 DVDD.n9425 DVDD.n188 0.353477
R8084 DVDD.n9616 DVDD.n122 0.353373
R8085 DVDD.n9673 DVDD.n46 0.347744
R8086 DVDD.n9318 DVDD.n432 0.347744
R8087 DVDD.n7507 DVDD.n7506 0.346681
R8088 DVDD.n8119 DVDD.n1747 0.346681
R8089 DVDD.n8289 DVDD.n8288 0.346681
R8090 DVDD.n8322 DVDD.n1620 0.346681
R8091 DVDD.n8360 DVDD.n8359 0.346681
R8092 DVDD.n8662 DVDD.n8661 0.346681
R8093 DVDD.n8650 DVDD.n8649 0.346681
R8094 DVDD.n6770 DVDD.n6769 0.346681
R8095 DVDD.n7287 DVDD.n7286 0.346681
R8096 DVDD.n8416 DVDD.n8415 0.343745
R8097 DVDD.n8441 DVDD.n8440 0.343745
R8098 DVDD.n1485 DVDD.n1382 0.343745
R8099 DVDD.n8494 DVDD.n8493 0.343745
R8100 DVDD.n8557 DVDD.n1393 0.343745
R8101 DVDD.n8602 DVDD.n8601 0.343745
R8102 DVDD.n9579 DVDD.n187 0.339299
R8103 DVDD.n9561 DVDD.n223 0.339029
R8104 DVDD.n9354 DVDD.n111 0.339029
R8105 DVDD.n6082 DVDD.n5908 0.338454
R8106 DVDD.n9354 DVDD.n122 0.338164
R8107 DVDD.n6082 DVDD.n5907 0.337829
R8108 DVDD.n9579 DVDD.n188 0.337829
R8109 DVDD.n9561 DVDD.n220 0.337254
R8110 DVDD.n8550 DVDD.n8549 0.334762
R8111 DVDD.n8531 DVDD.n8530 0.334761
R8112 DVDD.n2368 DVDD.n2335 0.274902
R8113 DVDD.n7743 DVDD.n2335 0.274902
R8114 DVDD.n7726 DVDD.n7702 0.274902
R8115 DVDD.n7726 DVDD.n7725 0.274902
R8116 DVDD.n8430 DVDD.n8428 0.269064
R8117 DVDD.n8433 DVDD.n8430 0.269064
R8118 DVDD.n8504 DVDD.n8503 0.269064
R8119 DVDD.n8503 DVDD.n8501 0.269064
R8120 DVDD.n8591 DVDD.n1370 0.269064
R8121 DVDD.n8592 DVDD.n8591 0.269064
R8122 DVDD.n7192 DVDD.n7191 0.256654
R8123 DVDD.n7175 DVDD.n7172 0.256654
R8124 DVDD.n8379 DVDD.n8378 0.256654
R8125 DVDD.n8631 DVDD.n1296 0.256654
R8126 DVDD.n744 DVDD.n649 0.243741
R8127 DVDD.n7184 DVDD.n7183 0.222038
R8128 DVDD.n7183 DVDD.n7182 0.222038
R8129 DVDD.n8639 DVDD.n1306 0.222038
R8130 DVDD.n8639 DVDD.n8638 0.222038
R8131 DVDD.n4614 DVDD.n4568 0.221946
R8132 DVDD.n9320 DVDD.n9319 0.218099
R8133 DVDD.n4111 DVDD.n3998 0.218099
R8134 DVDD.n9471 DVDD.n289 0.218099
R8135 DVDD.n8788 DVDD.n8787 0.218099
R8136 DVDD.n6777 DVDD.n2957 0.217859
R8137 DVDD.n9547 DVDD.n254 0.217859
R8138 DVDD.n4210 DVDD.n4151 0.217859
R8139 DVDD.n3588 DVDD.n1052 0.217859
R8140 DVDD.n8449 DVDD.n1302 0.21611
R8141 DVDD.n8387 DVDD.n8386 0.21611
R8142 DVDD.n5528 DVDD.n5508 0.214786
R8143 DVDD.n5526 DVDD.n5509 0.214786
R8144 DVDD.n5524 DVDD.n5510 0.214786
R8145 DVDD.n5513 DVDD.n5511 0.214786
R8146 DVDD.n5520 DVDD.n5514 0.214786
R8147 DVDD.n5519 DVDD.n5515 0.214786
R8148 DVDD.n5518 DVDD.n5517 0.214786
R8149 DVDD.n5516 DVDD.n3061 0.214786
R8150 DVDD.n6753 DVDD.n3062 0.214786
R8151 DVDD.n6752 DVDD.n6749 0.214786
R8152 DVDD.n6747 DVDD.n6746 0.214786
R8153 DVDD.n3064 DVDD.n3063 0.214786
R8154 DVDD.n6742 DVDD.n3066 0.214786
R8155 DVDD.n6741 DVDD.n3067 0.214786
R8156 DVDD.n6740 DVDD.n3068 0.214786
R8157 DVDD.n3071 DVDD.n3069 0.214786
R8158 DVDD.n6736 DVDD.n3072 0.214786
R8159 DVDD.n6735 DVDD.n3073 0.214786
R8160 DVDD.n6734 DVDD.n3074 0.214786
R8161 DVDD.n6732 DVDD.n3075 0.214786
R8162 DVDD.n6730 DVDD.n3076 0.214786
R8163 DVDD.n6728 DVDD.n3077 0.214786
R8164 DVDD.n6727 DVDD.n3078 0.214786
R8165 DVDD.n6726 DVDD.n3079 0.214786
R8166 DVDD.n3082 DVDD.n3080 0.214786
R8167 DVDD.n6722 DVDD.n3083 0.214786
R8168 DVDD.n6721 DVDD.n3084 0.214786
R8169 DVDD.n6720 DVDD.n3085 0.214786
R8170 DVDD.n3088 DVDD.n3086 0.214786
R8171 DVDD.n6716 DVDD.n3089 0.214786
R8172 DVDD.n6715 DVDD.n3090 0.214786
R8173 DVDD.n6714 DVDD.n3091 0.214786
R8174 DVDD.n3093 DVDD.n3092 0.214786
R8175 DVDD.n6710 DVDD.n3094 0.214786
R8176 DVDD.n6708 DVDD.n3095 0.214786
R8177 DVDD.n3188 DVDD.n3096 0.214786
R8178 DVDD.n3191 DVDD.n3190 0.214786
R8179 DVDD.n3192 DVDD.n3187 0.214786
R8180 DVDD.n6699 DVDD.n3193 0.214786
R8181 DVDD.n6698 DVDD.n3194 0.214786
R8182 DVDD.n6697 DVDD.n3195 0.214786
R8183 DVDD.n3198 DVDD.n3196 0.214786
R8184 DVDD.n6693 DVDD.n3199 0.214786
R8185 DVDD.n6692 DVDD.n3200 0.214786
R8186 DVDD.n6691 DVDD.n3201 0.214786
R8187 DVDD.n3204 DVDD.n3202 0.214786
R8188 DVDD.n6687 DVDD.n3205 0.214786
R8189 DVDD.n6686 DVDD.n3206 0.214786
R8190 DVDD.n6685 DVDD.n3207 0.214786
R8191 DVDD.n3210 DVDD.n3208 0.214786
R8192 DVDD.n6681 DVDD.n3211 0.214786
R8193 DVDD.n6680 DVDD.n3212 0.214786
R8194 DVDD.n6679 DVDD.n3213 0.214786
R8195 DVDD.n3308 DVDD.n3214 0.214786
R8196 DVDD.n3310 DVDD.n3309 0.214786
R8197 DVDD.n3311 DVDD.n3307 0.214786
R8198 DVDD.n6672 DVDD.n3312 0.214786
R8199 DVDD.n6671 DVDD.n3313 0.214786
R8200 DVDD.n6667 DVDD.n3316 0.214786
R8201 DVDD.n6666 DVDD.n3317 0.214786
R8202 DVDD.n6665 DVDD.n3318 0.214786
R8203 DVDD.n3321 DVDD.n3319 0.214786
R8204 DVDD.n6661 DVDD.n3322 0.214786
R8205 DVDD.n6660 DVDD.n3323 0.214786
R8206 DVDD.n6659 DVDD.n3324 0.214786
R8207 DVDD.n3327 DVDD.n3325 0.214786
R8208 DVDD.n6655 DVDD.n3328 0.214786
R8209 DVDD.n6654 DVDD.n3329 0.214786
R8210 DVDD.n6653 DVDD.n3330 0.214786
R8211 DVDD.n3366 DVDD.n3331 0.214786
R8212 DVDD.n3368 DVDD.n3367 0.214786
R8213 DVDD.n3371 DVDD.n3370 0.214786
R8214 DVDD.n3372 DVDD.n3365 0.214786
R8215 DVDD.n6643 DVDD.n3373 0.214786
R8216 DVDD.n6642 DVDD.n3374 0.214786
R8217 DVDD.n6641 DVDD.n3375 0.214786
R8218 DVDD.n3378 DVDD.n3376 0.214786
R8219 DVDD.n6637 DVDD.n3379 0.214786
R8220 DVDD.n6636 DVDD.n3380 0.214786
R8221 DVDD.n6635 DVDD.n3381 0.214786
R8222 DVDD.n3383 DVDD.n3382 0.214786
R8223 DVDD.n6631 DVDD.n3384 0.214786
R8224 DVDD.n6629 DVDD.n3385 0.214786
R8225 DVDD.n6628 DVDD.n3386 0.214786
R8226 DVDD.n6615 DVDD.n3387 0.214786
R8227 DVDD.n6613 DVDD.n3388 0.214786
R8228 DVDD.n3391 DVDD.n3389 0.214786
R8229 DVDD.n6609 DVDD.n3392 0.214786
R8230 DVDD.n6608 DVDD.n3393 0.214786
R8231 DVDD.n6607 DVDD.n3394 0.214786
R8232 DVDD.n6595 DVDD.n3395 0.214786
R8233 DVDD.n6596 DVDD.n6594 0.214786
R8234 DVDD.n6601 DVDD.n6597 0.214786
R8235 DVDD.n6600 DVDD.n6598 0.214786
R8236 DVDD.n7016 DVDD.n2551 0.214786
R8237 DVDD.n7015 DVDD.n2552 0.214786
R8238 DVDD.n7013 DVDD.n2553 0.214786
R8239 DVDD.n2556 DVDD.n2554 0.214786
R8240 DVDD.n7009 DVDD.n2557 0.214786
R8241 DVDD.n7008 DVDD.n2558 0.214786
R8242 DVDD.n7007 DVDD.n2559 0.214786
R8243 DVDD.n2612 DVDD.n2560 0.214786
R8244 DVDD.n2613 DVDD.n2611 0.214786
R8245 DVDD.n7001 DVDD.n2614 0.214786
R8246 DVDD.n6999 DVDD.n2616 0.214786
R8247 DVDD.n2619 DVDD.n2617 0.214786
R8248 DVDD.n6995 DVDD.n2620 0.214786
R8249 DVDD.n6994 DVDD.n2621 0.214786
R8250 DVDD.n6993 DVDD.n2622 0.214786
R8251 DVDD.n2625 DVDD.n2623 0.214786
R8252 DVDD.n6989 DVDD.n2626 0.214786
R8253 DVDD.n6988 DVDD.n2627 0.214786
R8254 DVDD.n6987 DVDD.n2628 0.214786
R8255 DVDD.n6942 DVDD.n2629 0.214786
R8256 DVDD.n6975 DVDD.n6943 0.214786
R8257 DVDD.n6974 DVDD.n6944 0.214786
R8258 DVDD.n6973 DVDD.n6945 0.214786
R8259 DVDD.n6972 DVDD.n6946 0.214786
R8260 DVDD.n6949 DVDD.n6947 0.214786
R8261 DVDD.n6968 DVDD.n6950 0.214786
R8262 DVDD.n6967 DVDD.n6951 0.214786
R8263 DVDD.n6966 DVDD.n6952 0.214786
R8264 DVDD.n6955 DVDD.n6953 0.214786
R8265 DVDD.n6962 DVDD.n6956 0.214786
R8266 DVDD.n6961 DVDD.n6957 0.214786
R8267 DVDD.n6960 DVDD.n6958 0.214786
R8268 DVDD.n2202 DVDD.n2201 0.214786
R8269 DVDD.n7789 DVDD.n7788 0.214786
R8270 DVDD.n7791 DVDD.n2197 0.214786
R8271 DVDD.n7793 DVDD.n7792 0.214786
R8272 DVDD.n2170 DVDD.n2169 0.214786
R8273 DVDD.n7809 DVDD.n7808 0.214786
R8274 DVDD.n7810 DVDD.n2168 0.214786
R8275 DVDD.n7812 DVDD.n7811 0.214786
R8276 DVDD.n2166 DVDD.n2165 0.214786
R8277 DVDD.n7817 DVDD.n7816 0.214786
R8278 DVDD.n7818 DVDD.n2164 0.214786
R8279 DVDD.n7820 DVDD.n7819 0.214786
R8280 DVDD.n2162 DVDD.n2161 0.214786
R8281 DVDD.n7825 DVDD.n7824 0.214786
R8282 DVDD.n7826 DVDD.n2160 0.214786
R8283 DVDD.n7828 DVDD.n7827 0.214786
R8284 DVDD.n2158 DVDD.n2157 0.214786
R8285 DVDD.n7833 DVDD.n7832 0.214786
R8286 DVDD.n7834 DVDD.n2156 0.214786
R8287 DVDD.n7836 DVDD.n7835 0.214786
R8288 DVDD.n2154 DVDD.n2153 0.214786
R8289 DVDD.n7845 DVDD.n7844 0.214786
R8290 DVDD.n7846 DVDD.n2152 0.214786
R8291 DVDD.n7849 DVDD.n7848 0.214786
R8292 DVDD.n7847 DVDD.n2118 0.214786
R8293 DVDD.n7855 DVDD.n2119 0.214786
R8294 DVDD.n7858 DVDD.n7857 0.214786
R8295 DVDD.n2115 DVDD.n2114 0.214786
R8296 DVDD.n7863 DVDD.n7862 0.214786
R8297 DVDD.n7864 DVDD.n2113 0.214786
R8298 DVDD.n7866 DVDD.n7865 0.214786
R8299 DVDD.n2111 DVDD.n2110 0.214786
R8300 DVDD.n7871 DVDD.n7870 0.214786
R8301 DVDD.n7872 DVDD.n2109 0.214786
R8302 DVDD.n7875 DVDD.n7874 0.214786
R8303 DVDD.n7873 DVDD.n2107 0.214786
R8304 DVDD.n7879 DVDD.n2106 0.214786
R8305 DVDD.n7881 DVDD.n7880 0.214786
R8306 DVDD.n7882 DVDD.n2105 0.214786
R8307 DVDD.n7884 DVDD.n7883 0.214786
R8308 DVDD.n2073 DVDD.n2072 0.214786
R8309 DVDD.n7896 DVDD.n7895 0.214786
R8310 DVDD.n7897 DVDD.n2071 0.214786
R8311 DVDD.n7899 DVDD.n7898 0.214786
R8312 DVDD.n2069 DVDD.n2068 0.214786
R8313 DVDD.n7904 DVDD.n7903 0.214786
R8314 DVDD.n7905 DVDD.n2067 0.214786
R8315 DVDD.n7907 DVDD.n7906 0.214786
R8316 DVDD.n2065 DVDD.n2064 0.214786
R8317 DVDD.n7912 DVDD.n7911 0.214786
R8318 DVDD.n7915 DVDD.n7914 0.214786
R8319 DVDD.n7928 DVDD.n2062 0.214786
R8320 DVDD.n7931 DVDD.n7930 0.214786
R8321 DVDD.n7932 DVDD.n2061 0.214786
R8322 DVDD.n7935 DVDD.n7934 0.214786
R8323 DVDD.n7933 DVDD.n2059 0.214786
R8324 DVDD.n7939 DVDD.n2058 0.214786
R8325 DVDD.n7941 DVDD.n7940 0.214786
R8326 DVDD.n7942 DVDD.n2057 0.214786
R8327 DVDD.n7950 DVDD.n7943 0.214786
R8328 DVDD.n7949 DVDD.n7944 0.214786
R8329 DVDD.n7947 DVDD.n7945 0.214786
R8330 DVDD.n2507 DVDD.n2506 0.214786
R8331 DVDD.n7553 DVDD.n7552 0.214786
R8332 DVDD.n7554 DVDD.n2505 0.214786
R8333 DVDD.n7556 DVDD.n7555 0.214786
R8334 DVDD.n2503 DVDD.n2502 0.214786
R8335 DVDD.n7561 DVDD.n7560 0.214786
R8336 DVDD.n7562 DVDD.n2501 0.214786
R8337 DVDD.n7564 DVDD.n7563 0.214786
R8338 DVDD.n2470 DVDD.n2469 0.214786
R8339 DVDD.n7596 DVDD.n7595 0.214786
R8340 DVDD.n7598 DVDD.n2466 0.214786
R8341 DVDD.n7600 DVDD.n7599 0.214786
R8342 DVDD.n2464 DVDD.n2463 0.214786
R8343 DVDD.n7605 DVDD.n7604 0.214786
R8344 DVDD.n7606 DVDD.n2462 0.214786
R8345 DVDD.n7608 DVDD.n7607 0.214786
R8346 DVDD.n2460 DVDD.n2459 0.214786
R8347 DVDD.n7613 DVDD.n7612 0.214786
R8348 DVDD.n7614 DVDD.n2458 0.214786
R8349 DVDD.n7655 DVDD.n7615 0.214786
R8350 DVDD.n7654 DVDD.n7616 0.214786
R8351 DVDD.n7652 DVDD.n7617 0.214786
R8352 DVDD.n7651 DVDD.n7618 0.214786
R8353 DVDD.n7650 DVDD.n7619 0.214786
R8354 DVDD.n7622 DVDD.n7620 0.214786
R8355 DVDD.n7646 DVDD.n7623 0.214786
R8356 DVDD.n7645 DVDD.n7624 0.214786
R8357 DVDD.n7644 DVDD.n7625 0.214786
R8358 DVDD.n7628 DVDD.n7626 0.214786
R8359 DVDD.n7640 DVDD.n7629 0.214786
R8360 DVDD.n7639 DVDD.n7630 0.214786
R8361 DVDD.n7638 DVDD.n7631 0.214786
R8362 DVDD.n7635 DVDD.n7632 0.214786
R8363 DVDD.n7634 DVDD.n7633 0.214786
R8364 DVDD.n7783 DVDD.n2208 0.214786
R8365 DVDD.n7782 DVDD.n2209 0.214786
R8366 DVDD.n2253 DVDD.n2210 0.214786
R8367 DVDD.n2254 DVDD.n2252 0.214786
R8368 DVDD.n7772 DVDD.n2255 0.214786
R8369 DVDD.n7771 DVDD.n2256 0.214786
R8370 DVDD.n7770 DVDD.n2257 0.214786
R8371 DVDD.n2260 DVDD.n2258 0.214786
R8372 DVDD.n7766 DVDD.n2261 0.214786
R8373 DVDD.n7765 DVDD.n2262 0.214786
R8374 DVDD.n7764 DVDD.n2263 0.214786
R8375 DVDD.n2266 DVDD.n2264 0.214786
R8376 DVDD.n7760 DVDD.n2267 0.214786
R8377 DVDD.n7759 DVDD.n2268 0.214786
R8378 DVDD.n7758 DVDD.n2269 0.214786
R8379 DVDD.n2272 DVDD.n2270 0.214786
R8380 DVDD.n7754 DVDD.n2273 0.214786
R8381 DVDD.n7753 DVDD.n2274 0.214786
R8382 DVDD.n7752 DVDD.n2275 0.214786
R8383 DVDD.n2309 DVDD.n2276 0.214786
R8384 DVDD.n2311 DVDD.n2310 0.214786
R8385 DVDD.n2312 DVDD.n2308 0.214786
R8386 DVDD.n2314 DVDD.n2313 0.214786
R8387 DVDD.n2315 DVDD.n1925 0.214786
R8388 DVDD.n8077 DVDD.n8076 0.214786
R8389 DVDD.n1928 DVDD.n1926 0.214786
R8390 DVDD.n8072 DVDD.n1931 0.214786
R8391 DVDD.n8071 DVDD.n1932 0.214786
R8392 DVDD.n8070 DVDD.n1933 0.214786
R8393 DVDD.n1936 DVDD.n1934 0.214786
R8394 DVDD.n8066 DVDD.n1937 0.214786
R8395 DVDD.n8065 DVDD.n1938 0.214786
R8396 DVDD.n8064 DVDD.n1939 0.214786
R8397 DVDD.n1942 DVDD.n1940 0.214786
R8398 DVDD.n8060 DVDD.n1943 0.214786
R8399 DVDD.n8059 DVDD.n1944 0.214786
R8400 DVDD.n8058 DVDD.n1945 0.214786
R8401 DVDD.n1990 DVDD.n1946 0.214786
R8402 DVDD.n1991 DVDD.n1989 0.214786
R8403 DVDD.n8048 DVDD.n1992 0.214786
R8404 DVDD.n8047 DVDD.n1993 0.214786
R8405 DVDD.n8046 DVDD.n1994 0.214786
R8406 DVDD.n1997 DVDD.n1995 0.214786
R8407 DVDD.n8042 DVDD.n1998 0.214786
R8408 DVDD.n8041 DVDD.n1999 0.214786
R8409 DVDD.n8040 DVDD.n2000 0.214786
R8410 DVDD.n2002 DVDD.n2001 0.214786
R8411 DVDD.n8036 DVDD.n2003 0.214786
R8412 DVDD.n8034 DVDD.n2005 0.214786
R8413 DVDD.n8033 DVDD.n2006 0.214786
R8414 DVDD.n8020 DVDD.n2007 0.214786
R8415 DVDD.n8018 DVDD.n2008 0.214786
R8416 DVDD.n2011 DVDD.n2009 0.214786
R8417 DVDD.n8014 DVDD.n2012 0.214786
R8418 DVDD.n8013 DVDD.n2013 0.214786
R8419 DVDD.n8012 DVDD.n2014 0.214786
R8420 DVDD.n8000 DVDD.n2015 0.214786
R8421 DVDD.n8001 DVDD.n7999 0.214786
R8422 DVDD.n8006 DVDD.n8002 0.214786
R8423 DVDD.n8005 DVDD.n8003 0.214786
R8424 DVDD.n8107 DVDD.n8106 0.214786
R8425 DVDD.n1852 DVDD.n1851 0.214786
R8426 DVDD.n8123 DVDD.n8122 0.214786
R8427 DVDD.n8124 DVDD.n1850 0.214786
R8428 DVDD.n8126 DVDD.n8125 0.214786
R8429 DVDD.n1848 DVDD.n1847 0.214786
R8430 DVDD.n8131 DVDD.n8130 0.214786
R8431 DVDD.n8132 DVDD.n1846 0.214786
R8432 DVDD.n8134 DVDD.n8133 0.214786
R8433 DVDD.n1844 DVDD.n1843 0.214786
R8434 DVDD.n8139 DVDD.n8138 0.214786
R8435 DVDD.n8142 DVDD.n8141 0.214786
R8436 DVDD.n8153 DVDD.n1840 0.214786
R8437 DVDD.n8156 DVDD.n8155 0.214786
R8438 DVDD.n8157 DVDD.n1839 0.214786
R8439 DVDD.n8160 DVDD.n8159 0.214786
R8440 DVDD.n8158 DVDD.n1837 0.214786
R8441 DVDD.n8164 DVDD.n1836 0.214786
R8442 DVDD.n8166 DVDD.n8165 0.214786
R8443 DVDD.n8167 DVDD.n1835 0.214786
R8444 DVDD.n8175 DVDD.n8168 0.214786
R8445 DVDD.n8174 DVDD.n8169 0.214786
R8446 DVDD.n8172 DVDD.n8170 0.214786
R8447 DVDD.n7224 DVDD.n7210 0.214786
R8448 DVDD.n7227 DVDD.n7226 0.214786
R8449 DVDD.n7228 DVDD.n7209 0.214786
R8450 DVDD.n7231 DVDD.n7230 0.214786
R8451 DVDD.n7229 DVDD.n7207 0.214786
R8452 DVDD.n7235 DVDD.n7206 0.214786
R8453 DVDD.n7237 DVDD.n7236 0.214786
R8454 DVDD.n7238 DVDD.n7205 0.214786
R8455 DVDD.n7271 DVDD.n7239 0.214786
R8456 DVDD.n7270 DVDD.n7240 0.214786
R8457 DVDD.n7267 DVDD.n7241 0.214786
R8458 DVDD.n7244 DVDD.n7242 0.214786
R8459 DVDD.n7263 DVDD.n7245 0.214786
R8460 DVDD.n7262 DVDD.n7246 0.214786
R8461 DVDD.n7261 DVDD.n7247 0.214786
R8462 DVDD.n7250 DVDD.n7248 0.214786
R8463 DVDD.n7257 DVDD.n7251 0.214786
R8464 DVDD.n7256 DVDD.n7252 0.214786
R8465 DVDD.n7255 DVDD.n7254 0.214786
R8466 DVDD.n7253 DVDD.n1563 0.214786
R8467 DVDD.n8347 DVDD.n1564 0.214786
R8468 DVDD.n8346 DVDD.n1565 0.214786
R8469 DVDD.n8344 DVDD.n1566 0.214786
R8470 DVDD.n1569 DVDD.n1567 0.214786
R8471 DVDD.n8340 DVDD.n1570 0.214786
R8472 DVDD.n8339 DVDD.n1571 0.214786
R8473 DVDD.n8338 DVDD.n1572 0.214786
R8474 DVDD.n1575 DVDD.n1573 0.214786
R8475 DVDD.n8334 DVDD.n1576 0.214786
R8476 DVDD.n8333 DVDD.n1577 0.214786
R8477 DVDD.n8332 DVDD.n1578 0.214786
R8478 DVDD.n1581 DVDD.n1579 0.214786
R8479 DVDD.n8328 DVDD.n1582 0.214786
R8480 DVDD.n8327 DVDD.n1583 0.214786
R8481 DVDD.n8325 DVDD.n1585 0.214786
R8482 DVDD.n1631 DVDD.n1586 0.214786
R8483 DVDD.n1632 DVDD.n1630 0.214786
R8484 DVDD.n8319 DVDD.n1633 0.214786
R8485 DVDD.n8318 DVDD.n1634 0.214786
R8486 DVDD.n1637 DVDD.n1635 0.214786
R8487 DVDD.n8314 DVDD.n1638 0.214786
R8488 DVDD.n8313 DVDD.n1639 0.214786
R8489 DVDD.n8312 DVDD.n1640 0.214786
R8490 DVDD.n1643 DVDD.n1641 0.214786
R8491 DVDD.n8308 DVDD.n1644 0.214786
R8492 DVDD.n8307 DVDD.n1645 0.214786
R8493 DVDD.n8306 DVDD.n1646 0.214786
R8494 DVDD.n1649 DVDD.n1647 0.214786
R8495 DVDD.n8302 DVDD.n1650 0.214786
R8496 DVDD.n8301 DVDD.n1651 0.214786
R8497 DVDD.n8300 DVDD.n1652 0.214786
R8498 DVDD.n1655 DVDD.n1653 0.214786
R8499 DVDD.n8296 DVDD.n1656 0.214786
R8500 DVDD.n8295 DVDD.n1657 0.214786
R8501 DVDD.n8294 DVDD.n1658 0.214786
R8502 DVDD.n1918 DVDD.n1659 0.214786
R8503 DVDD.n1920 DVDD.n1919 0.214786
R8504 DVDD.n1923 DVDD.n1922 0.214786
R8505 DVDD.n8081 DVDD.n8080 0.214786
R8506 DVDD.n1915 DVDD.n1914 0.214786
R8507 DVDD.n8086 DVDD.n8085 0.214786
R8508 DVDD.n8087 DVDD.n1913 0.214786
R8509 DVDD.n8089 DVDD.n8088 0.214786
R8510 DVDD.n1911 DVDD.n1910 0.214786
R8511 DVDD.n8094 DVDD.n8093 0.214786
R8512 DVDD.n8095 DVDD.n1909 0.214786
R8513 DVDD.n8098 DVDD.n8097 0.214786
R8514 DVDD.n8096 DVDD.n1907 0.214786
R8515 DVDD.n8102 DVDD.n1906 0.214786
R8516 DVDD.n8104 DVDD.n8103 0.214786
R8517 DVDD.n8105 DVDD.n1905 0.214786
R8518 DVDD.n8174 DVDD.n8173 0.214786
R8519 DVDD.n8176 DVDD.n8175 0.214786
R8520 DVDD.n1835 DVDD.n1814 0.214786
R8521 DVDD.n8165 DVDD.n1801 0.214786
R8522 DVDD.n8164 DVDD.n8163 0.214786
R8523 DVDD.n8162 DVDD.n1837 0.214786
R8524 DVDD.n8161 DVDD.n8160 0.214786
R8525 DVDD.n1839 DVDD.n1838 0.214786
R8526 DVDD.n8155 DVDD.n8154 0.214786
R8527 DVDD.n8153 DVDD.n8152 0.214786
R8528 DVDD.n8142 DVDD.n1249 0.214786
R8529 DVDD.n8138 DVDD.n8137 0.214786
R8530 DVDD.n8136 DVDD.n1844 0.214786
R8531 DVDD.n8135 DVDD.n8134 0.214786
R8532 DVDD.n1846 DVDD.n1845 0.214786
R8533 DVDD.n8130 DVDD.n8129 0.214786
R8534 DVDD.n8128 DVDD.n1848 0.214786
R8535 DVDD.n8127 DVDD.n8126 0.214786
R8536 DVDD.n1850 DVDD.n1849 0.214786
R8537 DVDD.n8122 DVDD.n8121 0.214786
R8538 DVDD.n1853 DVDD.n1852 0.214786
R8539 DVDD.n8108 DVDD.n8107 0.214786
R8540 DVDD.n7211 DVDD.n7043 0.214786
R8541 DVDD.n7224 DVDD.n7223 0.214786
R8542 DVDD.n7226 DVDD.n7225 0.214786
R8543 DVDD.n7209 DVDD.n7208 0.214786
R8544 DVDD.n7232 DVDD.n7231 0.214786
R8545 DVDD.n7233 DVDD.n7207 0.214786
R8546 DVDD.n7235 DVDD.n7234 0.214786
R8547 DVDD.n7236 DVDD.n7108 0.214786
R8548 DVDD.n7205 DVDD.n7120 0.214786
R8549 DVDD.n7272 DVDD.n7271 0.214786
R8550 DVDD.n7270 DVDD.n7269 0.214786
R8551 DVDD.n7267 DVDD.n7266 0.214786
R8552 DVDD.n7265 DVDD.n7242 0.214786
R8553 DVDD.n7264 DVDD.n7263 0.214786
R8554 DVDD.n7262 DVDD.n7243 0.214786
R8555 DVDD.n7261 DVDD.n7260 0.214786
R8556 DVDD.n7259 DVDD.n7248 0.214786
R8557 DVDD.n7258 DVDD.n7257 0.214786
R8558 DVDD.n7256 DVDD.n7249 0.214786
R8559 DVDD.n7255 DVDD.n1531 0.214786
R8560 DVDD.n1563 DVDD.n1544 0.214786
R8561 DVDD.n8348 DVDD.n8347 0.214786
R8562 DVDD.n8346 DVDD.n8345 0.214786
R8563 DVDD.n8344 DVDD.n8343 0.214786
R8564 DVDD.n8342 DVDD.n1567 0.214786
R8565 DVDD.n8341 DVDD.n8340 0.214786
R8566 DVDD.n8339 DVDD.n1568 0.214786
R8567 DVDD.n8338 DVDD.n8337 0.214786
R8568 DVDD.n8336 DVDD.n1573 0.214786
R8569 DVDD.n8335 DVDD.n8334 0.214786
R8570 DVDD.n8333 DVDD.n1574 0.214786
R8571 DVDD.n8332 DVDD.n8331 0.214786
R8572 DVDD.n8330 DVDD.n1579 0.214786
R8573 DVDD.n8329 DVDD.n8328 0.214786
R8574 DVDD.n8327 DVDD.n1580 0.214786
R8575 DVDD.n8325 DVDD.n8324 0.214786
R8576 DVDD.n1600 DVDD.n1586 0.214786
R8577 DVDD.n1630 DVDD.n1629 0.214786
R8578 DVDD.n8320 DVDD.n8319 0.214786
R8579 DVDD.n8318 DVDD.n8317 0.214786
R8580 DVDD.n8316 DVDD.n1635 0.214786
R8581 DVDD.n8315 DVDD.n8314 0.214786
R8582 DVDD.n8313 DVDD.n1636 0.214786
R8583 DVDD.n8312 DVDD.n8311 0.214786
R8584 DVDD.n8310 DVDD.n1641 0.214786
R8585 DVDD.n8309 DVDD.n8308 0.214786
R8586 DVDD.n8307 DVDD.n1642 0.214786
R8587 DVDD.n8306 DVDD.n8305 0.214786
R8588 DVDD.n8304 DVDD.n1647 0.214786
R8589 DVDD.n8303 DVDD.n8302 0.214786
R8590 DVDD.n8301 DVDD.n1648 0.214786
R8591 DVDD.n8300 DVDD.n8299 0.214786
R8592 DVDD.n8298 DVDD.n1653 0.214786
R8593 DVDD.n8297 DVDD.n8296 0.214786
R8594 DVDD.n8295 DVDD.n1654 0.214786
R8595 DVDD.n8294 DVDD.n8293 0.214786
R8596 DVDD.n1665 DVDD.n1659 0.214786
R8597 DVDD.n1920 DVDD.n1688 0.214786
R8598 DVDD.n1922 DVDD.n1921 0.214786
R8599 DVDD.n8082 DVDD.n8081 0.214786
R8600 DVDD.n8083 DVDD.n1915 0.214786
R8601 DVDD.n8085 DVDD.n8084 0.214786
R8602 DVDD.n1913 DVDD.n1912 0.214786
R8603 DVDD.n8090 DVDD.n8089 0.214786
R8604 DVDD.n8091 DVDD.n1911 0.214786
R8605 DVDD.n8093 DVDD.n8092 0.214786
R8606 DVDD.n1909 DVDD.n1908 0.214786
R8607 DVDD.n8099 DVDD.n8098 0.214786
R8608 DVDD.n8100 DVDD.n1907 0.214786
R8609 DVDD.n8102 DVDD.n8101 0.214786
R8610 DVDD.n8103 DVDD.n1892 0.214786
R8611 DVDD.n1905 DVDD.n1899 0.214786
R8612 DVDD.n8007 DVDD.n8006 0.214786
R8613 DVDD.n7999 DVDD.n7998 0.214786
R8614 DVDD.n7961 DVDD.n2015 0.214786
R8615 DVDD.n8012 DVDD.n8011 0.214786
R8616 DVDD.n8013 DVDD.n2010 0.214786
R8617 DVDD.n8015 DVDD.n8014 0.214786
R8618 DVDD.n8016 DVDD.n2009 0.214786
R8619 DVDD.n8018 DVDD.n8017 0.214786
R8620 DVDD.n8020 DVDD.n8019 0.214786
R8621 DVDD.n8033 DVDD.n8032 0.214786
R8622 DVDD.n8034 DVDD.n1210 0.214786
R8623 DVDD.n8037 DVDD.n8036 0.214786
R8624 DVDD.n8038 DVDD.n2001 0.214786
R8625 DVDD.n8040 DVDD.n8039 0.214786
R8626 DVDD.n8041 DVDD.n1996 0.214786
R8627 DVDD.n8043 DVDD.n8042 0.214786
R8628 DVDD.n8044 DVDD.n1995 0.214786
R8629 DVDD.n8046 DVDD.n8045 0.214786
R8630 DVDD.n8047 DVDD.n1988 0.214786
R8631 DVDD.n8049 DVDD.n8048 0.214786
R8632 DVDD.n1989 DVDD.n1973 0.214786
R8633 DVDD.n1954 DVDD.n1946 0.214786
R8634 DVDD.n8058 DVDD.n8057 0.214786
R8635 DVDD.n8059 DVDD.n1941 0.214786
R8636 DVDD.n8061 DVDD.n8060 0.214786
R8637 DVDD.n8062 DVDD.n1940 0.214786
R8638 DVDD.n8064 DVDD.n8063 0.214786
R8639 DVDD.n8065 DVDD.n1935 0.214786
R8640 DVDD.n8067 DVDD.n8066 0.214786
R8641 DVDD.n8068 DVDD.n1934 0.214786
R8642 DVDD.n8070 DVDD.n8069 0.214786
R8643 DVDD.n8071 DVDD.n1930 0.214786
R8644 DVDD.n8073 DVDD.n8072 0.214786
R8645 DVDD.n8074 DVDD.n1928 0.214786
R8646 DVDD.n8076 DVDD.n8075 0.214786
R8647 DVDD.n2316 DVDD.n2315 0.214786
R8648 DVDD.n2314 DVDD.n2295 0.214786
R8649 DVDD.n2308 DVDD.n2307 0.214786
R8650 DVDD.n2310 DVDD.n2285 0.214786
R8651 DVDD.n7750 DVDD.n2276 0.214786
R8652 DVDD.n7752 DVDD.n7751 0.214786
R8653 DVDD.n7753 DVDD.n2271 0.214786
R8654 DVDD.n7755 DVDD.n7754 0.214786
R8655 DVDD.n7756 DVDD.n2270 0.214786
R8656 DVDD.n7758 DVDD.n7757 0.214786
R8657 DVDD.n7759 DVDD.n2265 0.214786
R8658 DVDD.n7761 DVDD.n7760 0.214786
R8659 DVDD.n7762 DVDD.n2264 0.214786
R8660 DVDD.n7764 DVDD.n7763 0.214786
R8661 DVDD.n7765 DVDD.n2259 0.214786
R8662 DVDD.n7767 DVDD.n7766 0.214786
R8663 DVDD.n7768 DVDD.n2258 0.214786
R8664 DVDD.n7770 DVDD.n7769 0.214786
R8665 DVDD.n7771 DVDD.n2251 0.214786
R8666 DVDD.n7773 DVDD.n7772 0.214786
R8667 DVDD.n2252 DVDD.n2236 0.214786
R8668 DVDD.n2217 DVDD.n2210 0.214786
R8669 DVDD.n7782 DVDD.n7781 0.214786
R8670 DVDD.n7784 DVDD.n7783 0.214786
R8671 DVDD.n7634 DVDD.n2206 0.214786
R8672 DVDD.n7636 DVDD.n7635 0.214786
R8673 DVDD.n7638 DVDD.n7637 0.214786
R8674 DVDD.n7639 DVDD.n7627 0.214786
R8675 DVDD.n7641 DVDD.n7640 0.214786
R8676 DVDD.n7642 DVDD.n7626 0.214786
R8677 DVDD.n7644 DVDD.n7643 0.214786
R8678 DVDD.n7645 DVDD.n7621 0.214786
R8679 DVDD.n7647 DVDD.n7646 0.214786
R8680 DVDD.n7648 DVDD.n7620 0.214786
R8681 DVDD.n7650 DVDD.n7649 0.214786
R8682 DVDD.n7651 DVDD.n2388 0.214786
R8683 DVDD.n7652 DVDD.n2375 0.214786
R8684 DVDD.n7654 DVDD.n7653 0.214786
R8685 DVDD.n7656 DVDD.n7655 0.214786
R8686 DVDD.n2458 DVDD.n2451 0.214786
R8687 DVDD.n7612 DVDD.n7611 0.214786
R8688 DVDD.n7610 DVDD.n2460 0.214786
R8689 DVDD.n7609 DVDD.n7608 0.214786
R8690 DVDD.n2462 DVDD.n2461 0.214786
R8691 DVDD.n7604 DVDD.n7603 0.214786
R8692 DVDD.n7602 DVDD.n2464 0.214786
R8693 DVDD.n7601 DVDD.n7600 0.214786
R8694 DVDD.n2466 DVDD.n2465 0.214786
R8695 DVDD.n7595 DVDD.n7594 0.214786
R8696 DVDD.n7576 DVDD.n2470 0.214786
R8697 DVDD.n7565 DVDD.n7564 0.214786
R8698 DVDD.n2501 DVDD.n2489 0.214786
R8699 DVDD.n7560 DVDD.n7559 0.214786
R8700 DVDD.n7558 DVDD.n2503 0.214786
R8701 DVDD.n7557 DVDD.n7556 0.214786
R8702 DVDD.n2505 DVDD.n2504 0.214786
R8703 DVDD.n7552 DVDD.n7551 0.214786
R8704 DVDD.n7534 DVDD.n2507 0.214786
R8705 DVDD.n7523 DVDD.n7522 0.214786
R8706 DVDD.n7949 DVDD.n7948 0.214786
R8707 DVDD.n7951 DVDD.n7950 0.214786
R8708 DVDD.n2057 DVDD.n2043 0.214786
R8709 DVDD.n7940 DVDD.n2030 0.214786
R8710 DVDD.n7939 DVDD.n7938 0.214786
R8711 DVDD.n7937 DVDD.n2059 0.214786
R8712 DVDD.n7936 DVDD.n7935 0.214786
R8713 DVDD.n2061 DVDD.n2060 0.214786
R8714 DVDD.n7930 DVDD.n7929 0.214786
R8715 DVDD.n7928 DVDD.n7927 0.214786
R8716 DVDD.n7915 DVDD.n1171 0.214786
R8717 DVDD.n7911 DVDD.n7910 0.214786
R8718 DVDD.n7909 DVDD.n2065 0.214786
R8719 DVDD.n7908 DVDD.n7907 0.214786
R8720 DVDD.n2067 DVDD.n2066 0.214786
R8721 DVDD.n7903 DVDD.n7902 0.214786
R8722 DVDD.n7901 DVDD.n2069 0.214786
R8723 DVDD.n7900 DVDD.n7899 0.214786
R8724 DVDD.n2071 DVDD.n2070 0.214786
R8725 DVDD.n7895 DVDD.n7894 0.214786
R8726 DVDD.n2074 DVDD.n2073 0.214786
R8727 DVDD.n7885 DVDD.n7884 0.214786
R8728 DVDD.n2105 DVDD.n2101 0.214786
R8729 DVDD.n7880 DVDD.n2097 0.214786
R8730 DVDD.n7879 DVDD.n7878 0.214786
R8731 DVDD.n7877 DVDD.n2107 0.214786
R8732 DVDD.n7876 DVDD.n7875 0.214786
R8733 DVDD.n2109 DVDD.n2108 0.214786
R8734 DVDD.n7870 DVDD.n7869 0.214786
R8735 DVDD.n7868 DVDD.n2111 0.214786
R8736 DVDD.n7867 DVDD.n7866 0.214786
R8737 DVDD.n2113 DVDD.n2112 0.214786
R8738 DVDD.n7862 DVDD.n7861 0.214786
R8739 DVDD.n7860 DVDD.n2115 0.214786
R8740 DVDD.n7859 DVDD.n7858 0.214786
R8741 DVDD.n7855 DVDD.n7854 0.214786
R8742 DVDD.n2120 DVDD.n2118 0.214786
R8743 DVDD.n7850 DVDD.n7849 0.214786
R8744 DVDD.n2152 DVDD.n2151 0.214786
R8745 DVDD.n7844 DVDD.n7843 0.214786
R8746 DVDD.n7838 DVDD.n2154 0.214786
R8747 DVDD.n7837 DVDD.n7836 0.214786
R8748 DVDD.n2156 DVDD.n2155 0.214786
R8749 DVDD.n7832 DVDD.n7831 0.214786
R8750 DVDD.n7830 DVDD.n2158 0.214786
R8751 DVDD.n7829 DVDD.n7828 0.214786
R8752 DVDD.n2160 DVDD.n2159 0.214786
R8753 DVDD.n7824 DVDD.n7823 0.214786
R8754 DVDD.n7822 DVDD.n2162 0.214786
R8755 DVDD.n7821 DVDD.n7820 0.214786
R8756 DVDD.n2164 DVDD.n2163 0.214786
R8757 DVDD.n7816 DVDD.n7815 0.214786
R8758 DVDD.n7814 DVDD.n2166 0.214786
R8759 DVDD.n7813 DVDD.n7812 0.214786
R8760 DVDD.n2168 DVDD.n2167 0.214786
R8761 DVDD.n7808 DVDD.n7807 0.214786
R8762 DVDD.n7798 DVDD.n2170 0.214786
R8763 DVDD.n7794 DVDD.n7793 0.214786
R8764 DVDD.n2197 DVDD.n2193 0.214786
R8765 DVDD.n7788 DVDD.n7787 0.214786
R8766 DVDD.n2204 DVDD.n2202 0.214786
R8767 DVDD.n6960 DVDD.n6959 0.214786
R8768 DVDD.n6961 DVDD.n6954 0.214786
R8769 DVDD.n6963 DVDD.n6962 0.214786
R8770 DVDD.n6964 DVDD.n6953 0.214786
R8771 DVDD.n6966 DVDD.n6965 0.214786
R8772 DVDD.n6967 DVDD.n6948 0.214786
R8773 DVDD.n6969 DVDD.n6968 0.214786
R8774 DVDD.n6970 DVDD.n6947 0.214786
R8775 DVDD.n6972 DVDD.n6971 0.214786
R8776 DVDD.n6973 DVDD.n6939 0.214786
R8777 DVDD.n6974 DVDD.n6935 0.214786
R8778 DVDD.n6976 DVDD.n6975 0.214786
R8779 DVDD.n2638 DVDD.n2629 0.214786
R8780 DVDD.n6987 DVDD.n6986 0.214786
R8781 DVDD.n6988 DVDD.n2624 0.214786
R8782 DVDD.n6990 DVDD.n6989 0.214786
R8783 DVDD.n6991 DVDD.n2623 0.214786
R8784 DVDD.n6993 DVDD.n6992 0.214786
R8785 DVDD.n6994 DVDD.n2618 0.214786
R8786 DVDD.n6996 DVDD.n6995 0.214786
R8787 DVDD.n6997 DVDD.n2617 0.214786
R8788 DVDD.n6999 DVDD.n6998 0.214786
R8789 DVDD.n7002 DVDD.n7001 0.214786
R8790 DVDD.n2611 DVDD.n2610 0.214786
R8791 DVDD.n2573 DVDD.n2560 0.214786
R8792 DVDD.n7007 DVDD.n7006 0.214786
R8793 DVDD.n7008 DVDD.n2555 0.214786
R8794 DVDD.n7010 DVDD.n7009 0.214786
R8795 DVDD.n7011 DVDD.n2554 0.214786
R8796 DVDD.n7013 DVDD.n7012 0.214786
R8797 DVDD.n7015 DVDD.n7014 0.214786
R8798 DVDD.n7017 DVDD.n7016 0.214786
R8799 DVDD.n2550 DVDD.n2536 0.214786
R8800 DVDD.n6602 DVDD.n6601 0.214786
R8801 DVDD.n6594 DVDD.n6593 0.214786
R8802 DVDD.n3408 DVDD.n3395 0.214786
R8803 DVDD.n6607 DVDD.n6606 0.214786
R8804 DVDD.n6608 DVDD.n3390 0.214786
R8805 DVDD.n6610 DVDD.n6609 0.214786
R8806 DVDD.n6611 DVDD.n3389 0.214786
R8807 DVDD.n6613 DVDD.n6612 0.214786
R8808 DVDD.n6615 DVDD.n6614 0.214786
R8809 DVDD.n6628 DVDD.n6627 0.214786
R8810 DVDD.n6629 DVDD.n1132 0.214786
R8811 DVDD.n6632 DVDD.n6631 0.214786
R8812 DVDD.n6633 DVDD.n3382 0.214786
R8813 DVDD.n6635 DVDD.n6634 0.214786
R8814 DVDD.n6636 DVDD.n3377 0.214786
R8815 DVDD.n6638 DVDD.n6637 0.214786
R8816 DVDD.n6639 DVDD.n3376 0.214786
R8817 DVDD.n6641 DVDD.n6640 0.214786
R8818 DVDD.n6642 DVDD.n3364 0.214786
R8819 DVDD.n6644 DVDD.n6643 0.214786
R8820 DVDD.n3365 DVDD.n3363 0.214786
R8821 DVDD.n3370 DVDD.n3369 0.214786
R8822 DVDD.n3368 DVDD.n3344 0.214786
R8823 DVDD.n6651 DVDD.n3331 0.214786
R8824 DVDD.n6653 DVDD.n6652 0.214786
R8825 DVDD.n6654 DVDD.n3326 0.214786
R8826 DVDD.n6656 DVDD.n6655 0.214786
R8827 DVDD.n6657 DVDD.n3325 0.214786
R8828 DVDD.n6659 DVDD.n6658 0.214786
R8829 DVDD.n6660 DVDD.n3320 0.214786
R8830 DVDD.n6662 DVDD.n6661 0.214786
R8831 DVDD.n6663 DVDD.n3319 0.214786
R8832 DVDD.n6665 DVDD.n6664 0.214786
R8833 DVDD.n6666 DVDD.n3314 0.214786
R8834 DVDD.n6668 DVDD.n6667 0.214786
R8835 DVDD.n6671 DVDD.n6670 0.214786
R8836 DVDD.n6673 DVDD.n6672 0.214786
R8837 DVDD.n3307 DVDD.n3297 0.214786
R8838 DVDD.n3309 DVDD.n3227 0.214786
R8839 DVDD.n6677 DVDD.n3214 0.214786
R8840 DVDD.n6679 DVDD.n6678 0.214786
R8841 DVDD.n6680 DVDD.n3209 0.214786
R8842 DVDD.n6682 DVDD.n6681 0.214786
R8843 DVDD.n6683 DVDD.n3208 0.214786
R8844 DVDD.n6685 DVDD.n6684 0.214786
R8845 DVDD.n6686 DVDD.n3203 0.214786
R8846 DVDD.n6688 DVDD.n6687 0.214786
R8847 DVDD.n6689 DVDD.n3202 0.214786
R8848 DVDD.n6691 DVDD.n6690 0.214786
R8849 DVDD.n6692 DVDD.n3197 0.214786
R8850 DVDD.n6694 DVDD.n6693 0.214786
R8851 DVDD.n6695 DVDD.n3196 0.214786
R8852 DVDD.n6697 DVDD.n6696 0.214786
R8853 DVDD.n6698 DVDD.n3186 0.214786
R8854 DVDD.n6700 DVDD.n6699 0.214786
R8855 DVDD.n3187 DVDD.n3185 0.214786
R8856 DVDD.n3190 DVDD.n3189 0.214786
R8857 DVDD.n3109 DVDD.n3096 0.214786
R8858 DVDD.n6708 DVDD.n6707 0.214786
R8859 DVDD.n6711 DVDD.n6710 0.214786
R8860 DVDD.n6712 DVDD.n3092 0.214786
R8861 DVDD.n6714 DVDD.n6713 0.214786
R8862 DVDD.n6715 DVDD.n3087 0.214786
R8863 DVDD.n6717 DVDD.n6716 0.214786
R8864 DVDD.n6718 DVDD.n3086 0.214786
R8865 DVDD.n6720 DVDD.n6719 0.214786
R8866 DVDD.n6721 DVDD.n3081 0.214786
R8867 DVDD.n6723 DVDD.n6722 0.214786
R8868 DVDD.n6724 DVDD.n3080 0.214786
R8869 DVDD.n6726 DVDD.n6725 0.214786
R8870 DVDD.n6727 DVDD.n2672 0.214786
R8871 DVDD.n6728 DVDD.n2660 0.214786
R8872 DVDD.n6730 DVDD.n6729 0.214786
R8873 DVDD.n6732 DVDD.n6731 0.214786
R8874 DVDD.n6734 DVDD.n6733 0.214786
R8875 DVDD.n6735 DVDD.n3070 0.214786
R8876 DVDD.n6737 DVDD.n6736 0.214786
R8877 DVDD.n6738 DVDD.n3069 0.214786
R8878 DVDD.n6740 DVDD.n6739 0.214786
R8879 DVDD.n6741 DVDD.n3065 0.214786
R8880 DVDD.n6743 DVDD.n6742 0.214786
R8881 DVDD.n6744 DVDD.n3064 0.214786
R8882 DVDD.n6746 DVDD.n6745 0.214786
R8883 DVDD.n6752 DVDD.n6751 0.214786
R8884 DVDD.n6754 DVDD.n6753 0.214786
R8885 DVDD.n3061 DVDD.n3038 0.214786
R8886 DVDD.n5518 DVDD.n3026 0.214786
R8887 DVDD.n5519 DVDD.n5512 0.214786
R8888 DVDD.n5521 DVDD.n5520 0.214786
R8889 DVDD.n5522 DVDD.n5511 0.214786
R8890 DVDD.n5524 DVDD.n5523 0.214786
R8891 DVDD.n5526 DVDD.n5525 0.214786
R8892 DVDD.n5528 DVDD.n5527 0.214786
R8893 DVDD.n5530 DVDD.n5529 0.214786
R8894 DVDD.n5414 DVDD.n5378 0.214786
R8895 DVDD.n5412 DVDD.n5379 0.214786
R8896 DVDD.n5410 DVDD.n5380 0.214786
R8897 DVDD.n5383 DVDD.n5381 0.214786
R8898 DVDD.n5406 DVDD.n5384 0.214786
R8899 DVDD.n5405 DVDD.n5385 0.214786
R8900 DVDD.n5404 DVDD.n5386 0.214786
R8901 DVDD.n5403 DVDD.n5387 0.214786
R8902 DVDD.n5402 DVDD.n5389 0.214786
R8903 DVDD.n5388 DVDD.n4449 0.214786
R8904 DVDD.n5712 DVDD.n5711 0.214786
R8905 DVDD.n5713 DVDD.n4447 0.214786
R8906 DVDD.n5715 DVDD.n5714 0.214786
R8907 DVDD.n4445 DVDD.n4444 0.214786
R8908 DVDD.n5720 DVDD.n5719 0.214786
R8909 DVDD.n5721 DVDD.n4443 0.214786
R8910 DVDD.n5723 DVDD.n5722 0.214786
R8911 DVDD.n4441 DVDD.n4440 0.214786
R8912 DVDD.n5728 DVDD.n5727 0.214786
R8913 DVDD.n5729 DVDD.n4439 0.214786
R8914 DVDD.n5732 DVDD.n5730 0.214786
R8915 DVDD.n5733 DVDD.n4437 0.214786
R8916 DVDD.n5735 DVDD.n5734 0.214786
R8917 DVDD.n5736 DVDD.n4436 0.214786
R8918 DVDD.n5738 DVDD.n5737 0.214786
R8919 DVDD.n4434 DVDD.n4433 0.214786
R8920 DVDD.n5743 DVDD.n5742 0.214786
R8921 DVDD.n5744 DVDD.n4432 0.214786
R8922 DVDD.n5746 DVDD.n5745 0.214786
R8923 DVDD.n4430 DVDD.n4429 0.214786
R8924 DVDD.n5752 DVDD.n5751 0.214786
R8925 DVDD.n5753 DVDD.n4428 0.214786
R8926 DVDD.n5755 DVDD.n5754 0.214786
R8927 DVDD.n5756 DVDD.n4391 0.214786
R8928 DVDD.n6102 DVDD.n4390 0.214786
R8929 DVDD.n6104 DVDD.n6103 0.214786
R8930 DVDD.n4304 DVDD.n4303 0.214786
R8931 DVDD.n6116 DVDD.n6115 0.214786
R8932 DVDD.n6117 DVDD.n4302 0.214786
R8933 DVDD.n6119 DVDD.n6118 0.214786
R8934 DVDD.n4300 DVDD.n4299 0.214786
R8935 DVDD.n6124 DVDD.n6123 0.214786
R8936 DVDD.n6125 DVDD.n4298 0.214786
R8937 DVDD.n6127 DVDD.n6126 0.214786
R8938 DVDD.n4296 DVDD.n4295 0.214786
R8939 DVDD.n6132 DVDD.n6131 0.214786
R8940 DVDD.n6133 DVDD.n4294 0.214786
R8941 DVDD.n6135 DVDD.n6134 0.214786
R8942 DVDD.n4292 DVDD.n4291 0.214786
R8943 DVDD.n6140 DVDD.n6139 0.214786
R8944 DVDD.n6141 DVDD.n4290 0.214786
R8945 DVDD.n6143 DVDD.n6142 0.214786
R8946 DVDD.n4288 DVDD.n4287 0.214786
R8947 DVDD.n6148 DVDD.n6147 0.214786
R8948 DVDD.n6149 DVDD.n4286 0.214786
R8949 DVDD.n6151 DVDD.n6150 0.214786
R8950 DVDD.n3945 DVDD.n3944 0.214786
R8951 DVDD.n6158 DVDD.n6157 0.214786
R8952 DVDD.n6161 DVDD.n6160 0.214786
R8953 DVDD.n3911 DVDD.n3910 0.214786
R8954 DVDD.n6166 DVDD.n6165 0.214786
R8955 DVDD.n6167 DVDD.n3909 0.214786
R8956 DVDD.n6169 DVDD.n6168 0.214786
R8957 DVDD.n3907 DVDD.n3906 0.214786
R8958 DVDD.n6174 DVDD.n6173 0.214786
R8959 DVDD.n6175 DVDD.n3905 0.214786
R8960 DVDD.n6177 DVDD.n6176 0.214786
R8961 DVDD.n3903 DVDD.n3902 0.214786
R8962 DVDD.n6183 DVDD.n6182 0.214786
R8963 DVDD.n6184 DVDD.n3901 0.214786
R8964 DVDD.n6187 DVDD.n6185 0.214786
R8965 DVDD.n6189 DVDD.n3900 0.214786
R8966 DVDD.n6191 DVDD.n6190 0.214786
R8967 DVDD.n6192 DVDD.n3899 0.214786
R8968 DVDD.n6194 DVDD.n6193 0.214786
R8969 DVDD.n3898 DVDD.n3897 0.214786
R8970 DVDD.n6199 DVDD.n6198 0.214786
R8971 DVDD.n6200 DVDD.n3896 0.214786
R8972 DVDD.n6202 DVDD.n6201 0.214786
R8973 DVDD.n3894 DVDD.n3893 0.214786
R8974 DVDD.n6208 DVDD.n6207 0.214786
R8975 DVDD.n6209 DVDD.n3510 0.214786
R8976 DVDD.n6423 DVDD.n3511 0.214786
R8977 DVDD.n6422 DVDD.n3512 0.214786
R8978 DVDD.n6409 DVDD.n3513 0.214786
R8979 DVDD.n6407 DVDD.n3514 0.214786
R8980 DVDD.n3517 DVDD.n3515 0.214786
R8981 DVDD.n6403 DVDD.n3518 0.214786
R8982 DVDD.n6402 DVDD.n3519 0.214786
R8983 DVDD.n6401 DVDD.n3520 0.214786
R8984 DVDD.n6389 DVDD.n3521 0.214786
R8985 DVDD.n6390 DVDD.n6388 0.214786
R8986 DVDD.n6395 DVDD.n6391 0.214786
R8987 DVDD.n6394 DVDD.n6392 0.214786
R8988 DVDD.n6396 DVDD.n6395 0.214786
R8989 DVDD.n6388 DVDD.n6387 0.214786
R8990 DVDD.n3534 DVDD.n3521 0.214786
R8991 DVDD.n6401 DVDD.n6400 0.214786
R8992 DVDD.n6402 DVDD.n3516 0.214786
R8993 DVDD.n6404 DVDD.n6403 0.214786
R8994 DVDD.n6405 DVDD.n3515 0.214786
R8995 DVDD.n6407 DVDD.n6406 0.214786
R8996 DVDD.n6409 DVDD.n6408 0.214786
R8997 DVDD.n6422 DVDD.n6421 0.214786
R8998 DVDD.n6423 DVDD.n1070 0.214786
R8999 DVDD.n6205 DVDD.n3510 0.214786
R9000 DVDD.n6207 DVDD.n6206 0.214786
R9001 DVDD.n6204 DVDD.n3894 0.214786
R9002 DVDD.n6203 DVDD.n6202 0.214786
R9003 DVDD.n3896 DVDD.n3895 0.214786
R9004 DVDD.n6198 DVDD.n6197 0.214786
R9005 DVDD.n6196 DVDD.n3898 0.214786
R9006 DVDD.n6195 DVDD.n6194 0.214786
R9007 DVDD.n3899 DVDD.n3808 0.214786
R9008 DVDD.n6190 DVDD.n3561 0.214786
R9009 DVDD.n6189 DVDD.n6188 0.214786
R9010 DVDD.n6187 DVDD.n6186 0.214786
R9011 DVDD.n6180 DVDD.n3901 0.214786
R9012 DVDD.n6182 DVDD.n6181 0.214786
R9013 DVDD.n6179 DVDD.n3903 0.214786
R9014 DVDD.n6178 DVDD.n6177 0.214786
R9015 DVDD.n3905 DVDD.n3904 0.214786
R9016 DVDD.n6173 DVDD.n6172 0.214786
R9017 DVDD.n6171 DVDD.n3907 0.214786
R9018 DVDD.n6170 DVDD.n6169 0.214786
R9019 DVDD.n3909 DVDD.n3908 0.214786
R9020 DVDD.n6165 DVDD.n6164 0.214786
R9021 DVDD.n6163 DVDD.n3911 0.214786
R9022 DVDD.n6162 DVDD.n6161 0.214786
R9023 DVDD.n6157 DVDD.n6156 0.214786
R9024 DVDD.n3946 DVDD.n3945 0.214786
R9025 DVDD.n6152 DVDD.n6151 0.214786
R9026 DVDD.n4286 DVDD.n4283 0.214786
R9027 DVDD.n6147 DVDD.n6146 0.214786
R9028 DVDD.n6145 DVDD.n4288 0.214786
R9029 DVDD.n6144 DVDD.n6143 0.214786
R9030 DVDD.n4290 DVDD.n4289 0.214786
R9031 DVDD.n6139 DVDD.n6138 0.214786
R9032 DVDD.n6137 DVDD.n4292 0.214786
R9033 DVDD.n6136 DVDD.n6135 0.214786
R9034 DVDD.n4294 DVDD.n4293 0.214786
R9035 DVDD.n6131 DVDD.n6130 0.214786
R9036 DVDD.n6129 DVDD.n4296 0.214786
R9037 DVDD.n6128 DVDD.n6127 0.214786
R9038 DVDD.n4298 DVDD.n4297 0.214786
R9039 DVDD.n6123 DVDD.n6122 0.214786
R9040 DVDD.n6121 DVDD.n4300 0.214786
R9041 DVDD.n6120 DVDD.n6119 0.214786
R9042 DVDD.n4302 DVDD.n4301 0.214786
R9043 DVDD.n6115 DVDD.n6114 0.214786
R9044 DVDD.n6106 DVDD.n4304 0.214786
R9045 DVDD.n6105 DVDD.n6104 0.214786
R9046 DVDD.n5758 DVDD.n4390 0.214786
R9047 DVDD.n5757 DVDD.n5756 0.214786
R9048 DVDD.n5755 DVDD.n4427 0.214786
R9049 DVDD.n5749 DVDD.n4428 0.214786
R9050 DVDD.n5751 DVDD.n5750 0.214786
R9051 DVDD.n5748 DVDD.n4430 0.214786
R9052 DVDD.n5747 DVDD.n5746 0.214786
R9053 DVDD.n4432 DVDD.n4431 0.214786
R9054 DVDD.n5742 DVDD.n5741 0.214786
R9055 DVDD.n5740 DVDD.n4434 0.214786
R9056 DVDD.n5739 DVDD.n5738 0.214786
R9057 DVDD.n4436 DVDD.n4435 0.214786
R9058 DVDD.n5734 DVDD.n2820 0.214786
R9059 DVDD.n5733 DVDD.n2808 0.214786
R9060 DVDD.n5732 DVDD.n5731 0.214786
R9061 DVDD.n4439 DVDD.n4438 0.214786
R9062 DVDD.n5727 DVDD.n5726 0.214786
R9063 DVDD.n5725 DVDD.n4441 0.214786
R9064 DVDD.n5724 DVDD.n5723 0.214786
R9065 DVDD.n4443 DVDD.n4442 0.214786
R9066 DVDD.n5719 DVDD.n5718 0.214786
R9067 DVDD.n5717 DVDD.n4445 0.214786
R9068 DVDD.n5716 DVDD.n5715 0.214786
R9069 DVDD.n4447 DVDD.n4446 0.214786
R9070 DVDD.n5711 DVDD.n5710 0.214786
R9071 DVDD.n5676 DVDD.n4449 0.214786
R9072 DVDD.n5402 DVDD.n5401 0.214786
R9073 DVDD.n5403 DVDD.n2975 0.214786
R9074 DVDD.n5404 DVDD.n2963 0.214786
R9075 DVDD.n5405 DVDD.n5382 0.214786
R9076 DVDD.n5407 DVDD.n5406 0.214786
R9077 DVDD.n5408 DVDD.n5381 0.214786
R9078 DVDD.n5410 DVDD.n5409 0.214786
R9079 DVDD.n5412 DVDD.n5411 0.214786
R9080 DVDD.n5414 DVDD.n5413 0.214786
R9081 DVDD.n5416 DVDD.n5415 0.214786
R9082 DVDD.n2893 DVDD.n226 0.214786
R9083 DVDD.n9564 DVDD.n212 0.214786
R9084 DVDD.n9565 DVDD.n211 0.214786
R9085 DVDD.n4508 DVDD.n209 0.214786
R9086 DVDD.n9571 DVDD.n206 0.214786
R9087 DVDD.n393 DVDD.n204 0.214786
R9088 DVDD.n9333 DVDD.n358 0.214786
R9089 DVDD.n9334 DVDD.n170 0.214786
R9090 DVDD.n9332 DVDD.n167 0.214786
R9091 DVDD.n9338 DVDD.n166 0.214786
R9092 DVDD.n9340 DVDD.n146 0.214786
R9093 DVDD.n9346 DVDD.n108 0.214786
R9094 DVDD.n9324 DVDD.n106 0.214786
R9095 DVDD.n9323 DVDD.n409 0.214786
R9096 DVDD.n9322 DVDD.n428 0.214786
R9097 DVDD.n430 DVDD.n427 0.214786
R9098 DVDD.n9345 DVDD.n129 0.214786
R9099 DVDD.n9344 DVDD.n9328 0.214786
R9100 DVDD.n9330 DVDD.n9329 0.214786
R9101 DVDD.n9339 DVDD.n151 0.214786
R9102 DVDD.n9577 DVDD.n201 0.214786
R9103 DVDD.n9576 DVDD.n202 0.214786
R9104 DVDD.n9575 DVDD.n203 0.214786
R9105 DVDD.n9570 DVDD.n207 0.214786
R9106 DVDD.n9569 DVDD.n208 0.214786
R9107 DVDD.n5297 DVDD.n2894 0.214786
R9108 DVDD.n5300 DVDD.n2898 0.214786
R9109 DVDD.n5302 DVDD.n5301 0.214786
R9110 DVDD.n5300 DVDD.n5299 0.214786
R9111 DVDD.n5298 DVDD.n5297 0.214786
R9112 DVDD.n237 DVDD.n226 0.214786
R9113 DVDD.n9564 DVDD.n210 0.214786
R9114 DVDD.n9566 DVDD.n9565 0.214786
R9115 DVDD.n9567 DVDD.n209 0.214786
R9116 DVDD.n9569 DVDD.n9568 0.214786
R9117 DVDD.n9570 DVDD.n205 0.214786
R9118 DVDD.n9572 DVDD.n9571 0.214786
R9119 DVDD.n9573 DVDD.n204 0.214786
R9120 DVDD.n9575 DVDD.n9574 0.214786
R9121 DVDD.n9576 DVDD.n199 0.214786
R9122 DVDD.n9578 DVDD.n9577 0.214786
R9123 DVDD.n9333 DVDD.n198 0.214786
R9124 DVDD.n9335 DVDD.n9334 0.214786
R9125 DVDD.n9336 DVDD.n9332 0.214786
R9126 DVDD.n9338 DVDD.n9337 0.214786
R9127 DVDD.n9339 DVDD.n9331 0.214786
R9128 DVDD.n9341 DVDD.n9340 0.214786
R9129 DVDD.n9342 DVDD.n9330 0.214786
R9130 DVDD.n9344 DVDD.n9343 0.214786
R9131 DVDD.n9345 DVDD.n9326 0.214786
R9132 DVDD.n9347 DVDD.n9346 0.214786
R9133 DVDD.n9325 DVDD.n9324 0.214786
R9134 DVDD.n9323 DVDD.n426 0.214786
R9135 DVDD.n9322 DVDD.n9321 0.214786
R9136 DVDD.n241 DVDD.n240 0.214786
R9137 DVDD.n9559 DVDD.n9558 0.214786
R9138 DVDD.n9560 DVDD.n222 0.214786
R9139 DVDD.n239 DVDD.n221 0.214786
R9140 DVDD.n9502 DVDD.n9501 0.214786
R9141 DVDD.n9500 DVDD.n269 0.214786
R9142 DVDD.n9499 DVDD.n9498 0.214786
R9143 DVDD.n271 DVDD.n270 0.214786
R9144 DVDD.n9489 DVDD.n9488 0.214786
R9145 DVDD.n9487 DVDD.n278 0.214786
R9146 DVDD.n9486 DVDD.n9485 0.214786
R9147 DVDD.n280 DVDD.n279 0.214786
R9148 DVDD.n360 DVDD.n195 0.214786
R9149 DVDD.n9429 DVDD.n196 0.214786
R9150 DVDD.n9428 DVDD.n9427 0.214786
R9151 DVDD.n9426 DVDD.n328 0.214786
R9152 DVDD.n9441 DVDD.n327 0.214786
R9153 DVDD.n9442 DVDD.n326 0.214786
R9154 DVDD.n9443 DVDD.n325 0.214786
R9155 DVDD.n324 DVDD.n312 0.214786
R9156 DVDD.n9454 DVDD.n311 0.214786
R9157 DVDD.n9455 DVDD.n310 0.214786
R9158 DVDD.n425 DVDD.n309 0.214786
R9159 DVDD.n418 DVDD.n417 0.214786
R9160 DVDD.n416 DVDD.n292 0.214786
R9161 DVDD.n9468 DVDD.n291 0.214786
R9162 DVDD.n242 DVDD.n222 0.214786
R9163 DVDD.n9504 DVDD.n221 0.214786
R9164 DVDD.n9503 DVDD.n9502 0.214786
R9165 DVDD.n273 DVDD.n269 0.214786
R9166 DVDD.n9490 DVDD.n9489 0.214786
R9167 DVDD.n278 DVDD.n276 0.214786
R9168 DVDD.n9430 DVDD.n9429 0.214786
R9169 DVDD.n9428 DVDD.n347 0.214786
R9170 DVDD.n330 DVDD.n328 0.214786
R9171 DVDD.n9441 DVDD.n9440 0.214786
R9172 DVDD.n9444 DVDD.n9443 0.214786
R9173 DVDD.n309 DVDD.n124 0.214786
R9174 DVDD.n417 DVDD.n123 0.214786
R9175 DVDD.n294 DVDD.n292 0.214786
R9176 DVDD.n9468 DVDD.n9467 0.214786
R9177 DVDD.n9470 DVDD.n9469 0.214786
R9178 DVDD.n9456 DVDD.n9455 0.214786
R9179 DVDD.n9454 DVDD.n9453 0.214786
R9180 DVDD.n313 DVDD.n312 0.214786
R9181 DVDD.n9442 DVDD.n323 0.214786
R9182 DVDD.n361 DVDD.n360 0.214786
R9183 DVDD.n362 DVDD.n280 0.214786
R9184 DVDD.n9485 DVDD.n9484 0.214786
R9185 DVDD.n277 DVDD.n271 0.214786
R9186 DVDD.n9498 DVDD.n9497 0.214786
R9187 DVDD.n9558 DVDD.n9557 0.214786
R9188 DVDD.n244 DVDD.n241 0.214786
R9189 DVDD.n253 DVDD.n252 0.214786
R9190 DVDD.n3590 DVDD.n3587 0.214786
R9191 DVDD.n3586 DVDD.n3585 0.214786
R9192 DVDD.n231 DVDD.n215 0.214786
R9193 DVDD.n232 DVDD.n216 0.214786
R9194 DVDD.n1030 DVDD.n1029 0.214786
R9195 DVDD.n1031 DVDD.n1028 0.214786
R9196 DVDD.n1027 DVDD.n1015 0.214786
R9197 DVDD.n1026 DVDD.n1025 0.214786
R9198 DVDD.n1024 DVDD.n1016 0.214786
R9199 DVDD.n1023 DVDD.n1022 0.214786
R9200 DVDD.n1021 DVDD.n1017 0.214786
R9201 DVDD.n1020 DVDD.n1019 0.214786
R9202 DVDD.n1018 DVDD.n191 0.214786
R9203 DVDD.n972 DVDD.n190 0.214786
R9204 DVDD.n973 DVDD.n971 0.214786
R9205 DVDD.n974 DVDD.n970 0.214786
R9206 DVDD.n975 DVDD.n969 0.214786
R9207 DVDD.n968 DVDD.n957 0.214786
R9208 DVDD.n967 DVDD.n966 0.214786
R9209 DVDD.n964 DVDD.n958 0.214786
R9210 DVDD.n963 DVDD.n962 0.214786
R9211 DVDD.n961 DVDD.n960 0.214786
R9212 DVDD.n959 DVDD.n419 0.214786
R9213 DVDD.n8783 DVDD.n420 0.214786
R9214 DVDD.n8784 DVDD.n8782 0.214786
R9215 DVDD.n8786 DVDD.n8785 0.214786
R9216 DVDD.n4148 DVDD.n218 0.214786
R9217 DVDD.n4144 DVDD.n219 0.214786
R9218 DVDD.n4143 DVDD.n4142 0.214786
R9219 DVDD.n3982 DVDD.n3978 0.214786
R9220 DVDD.n4130 DVDD.n4129 0.214786
R9221 DVDD.n3987 DVDD.n3985 0.214786
R9222 DVDD.n4081 DVDD.n373 0.214786
R9223 DVDD.n4082 DVDD.n4080 0.214786
R9224 DVDD.n4083 DVDD.n4026 0.214786
R9225 DVDD.n4060 DVDD.n4024 0.214786
R9226 DVDD.n4088 DVDD.n4022 0.214786
R9227 DVDD.n4018 DVDD.n120 0.214786
R9228 DVDD.n4104 DVDD.n121 0.214786
R9229 DVDD.n4105 DVDD.n4103 0.214786
R9230 DVDD.n4108 DVDD.n4000 0.214786
R9231 DVDD.n4110 DVDD.n4109 0.214786
R9232 DVDD.n4094 DVDD.n4093 0.214786
R9233 DVDD.n4041 DVDD.n4019 0.214786
R9234 DVDD.n4089 DVDD.n4021 0.214786
R9235 DVDD.n4087 DVDD.n4023 0.214786
R9236 DVDD.n3989 DVDD.n371 0.214786
R9237 DVDD.n4071 DVDD.n3990 0.214786
R9238 DVDD.n4125 DVDD.n4124 0.214786
R9239 DVDD.n3986 DVDD.n3980 0.214786
R9240 DVDD.n4138 DVDD.n4137 0.214786
R9241 DVDD.n4214 DVDD.n4213 0.214786
R9242 DVDD.n4152 DVDD.n4150 0.214786
R9243 DVDD.n4209 DVDD.n4208 0.214786
R9244 DVDD.n4211 DVDD.n4150 0.214786
R9245 DVDD.n4213 DVDD.n4212 0.214786
R9246 DVDD.n234 DVDD.n218 0.214786
R9247 DVDD.n235 DVDD.n219 0.214786
R9248 DVDD.n4142 DVDD.n4141 0.214786
R9249 DVDD.n4140 DVDD.n3978 0.214786
R9250 DVDD.n4139 DVDD.n4138 0.214786
R9251 DVDD.n3980 DVDD.n3979 0.214786
R9252 DVDD.n4129 DVDD.n4128 0.214786
R9253 DVDD.n4127 DVDD.n3987 0.214786
R9254 DVDD.n4126 DVDD.n4125 0.214786
R9255 DVDD.n3990 DVDD.n3988 0.214786
R9256 DVDD.n3989 DVDD.n185 0.214786
R9257 DVDD.n4081 DVDD.n186 0.214786
R9258 DVDD.n4082 DVDD.n4025 0.214786
R9259 DVDD.n4084 DVDD.n4083 0.214786
R9260 DVDD.n4085 DVDD.n4024 0.214786
R9261 DVDD.n4087 DVDD.n4086 0.214786
R9262 DVDD.n4088 DVDD.n4020 0.214786
R9263 DVDD.n4090 DVDD.n4089 0.214786
R9264 DVDD.n4091 DVDD.n4019 0.214786
R9265 DVDD.n4093 DVDD.n4092 0.214786
R9266 DVDD.n4018 DVDD.n423 0.214786
R9267 DVDD.n4104 DVDD.n424 0.214786
R9268 DVDD.n4106 DVDD.n4105 0.214786
R9269 DVDD.n4108 DVDD.n4107 0.214786
R9270 DVDD.n1037 DVDD.n215 0.214786
R9271 DVDD.n1012 DVDD.n216 0.214786
R9272 DVDD.n1030 DVDD.n1011 0.214786
R9273 DVDD.n1032 DVDD.n1031 0.214786
R9274 DVDD.n1024 DVDD.n907 0.214786
R9275 DVDD.n1023 DVDD.n906 0.214786
R9276 DVDD.n972 DVDD.n352 0.214786
R9277 DVDD.n973 DVDD.n883 0.214786
R9278 DVDD.n974 DVDD.n882 0.214786
R9279 DVDD.n976 DVDD.n975 0.214786
R9280 DVDD.n966 DVDD.n965 0.214786
R9281 DVDD.n959 DVDD.n116 0.214786
R9282 DVDD.n8783 DVDD.n117 0.214786
R9283 DVDD.n8784 DVDD.n89 0.214786
R9284 DVDD.n8785 DVDD.n88 0.214786
R9285 DVDD.n8781 DVDD.n84 0.214786
R9286 DVDD.n960 DVDD.n850 0.214786
R9287 DVDD.n963 DVDD.n853 0.214786
R9288 DVDD.n964 DVDD.n866 0.214786
R9289 DVDD.n957 DVDD.n870 0.214786
R9290 DVDD.n1018 DVDD.n349 0.214786
R9291 DVDD.n1019 DVDD.n891 0.214786
R9292 DVDD.n1017 DVDD.n894 0.214786
R9293 DVDD.n1025 DVDD.n911 0.214786
R9294 DVDD.n1015 DVDD.n912 0.214786
R9295 DVDD.n3585 DVDD.n1038 0.214786
R9296 DVDD.n3591 DVDD.n3590 0.214786
R9297 DVDD.n3589 DVDD.n1051 0.214786
R9298 DVDD.n8495 DVDD.n1432 0.210972
R9299 DVDD.n8600 DVDD.n1354 0.210972
R9300 DVDD.n8499 DVDD.n1424 0.210972
R9301 DVDD.n8595 DVDD.n1363 0.210972
R9302 DVDD.n8505 DVDD.n1418 0.210972
R9303 DVDD.n8511 DVDD.n8508 0.210972
R9304 DVDD.n8417 DVDD.n1488 0.210972
R9305 DVDD.n1486 DVDD.n1483 0.210972
R9306 DVDD.n8628 DVDD.n8627 0.210618
R9307 DVDD.n1330 DVDD.n1314 0.210618
R9308 DVDD.n7359 DVDD.n7358 0.210618
R9309 DVDD.n8377 DVDD.n1506 0.210618
R9310 DVDD.n353 DVDD 0.209761
R9311 DVDD.n9425 DVDD.n184 0.207132
R9312 DVDD.n9616 DVDD.n104 0.207064
R9313 DVDD.n228 DVDD.n227 0.207064
R9314 DVDD.n8625 DVDD.n1328 0.206898
R9315 DVDD.n8598 DVDD.n1360 0.206898
R9316 DVDD.n8622 DVDD.n1334 0.206898
R9317 DVDD.n8593 DVDD.n1369 0.206898
R9318 DVDD.n8427 DVDD.n1458 0.206898
R9319 DVDD.n8516 DVDD.n8514 0.206898
R9320 DVDD.n8419 DVDD.n1462 0.206898
R9321 DVDD.n1481 DVDD.n1401 0.206898
R9322 DVDD.n9562 DVDD.n228 0.2068
R9323 DVDD.n5646 DVDD.n5640 0.2067
R9324 DVDD.n5645 DVDD.n5640 0.206533
R9325 DVDD.n9425 DVDD.n183 0.206229
R9326 DVDD.n9616 DVDD.n105 0.205961
R9327 DVDD.n353 DVDD 0.203577
R9328 DVDD.n9579 DVDD.n184 0.199885
R9329 DVDD.n5647 DVDD.n5646 0.19985
R9330 DVDD.n9354 DVDD.n104 0.19948
R9331 DVDD.n9561 DVDD.n227 0.19948
R9332 DVDD.n9354 DVDD.n105 0.199195
R9333 DVDD.n9579 DVDD.n183 0.198923
R9334 DVDD.n5647 DVDD.n5645 0.198626
R9335 DVDD.n9562 DVDD.n9561 0.198351
R9336 DVDD.n3764 DVDD.n3533 0.178448
R9337 DVDD.n228 DVDD.n213 0.174559
R9338 DVDD.n9425 DVDD.n192 0.174559
R9339 DVDD.n9616 DVDD.n119 0.173987
R9340 DVDD.n229 DVDD 0.172062
R9341 DVDD.n422 DVDD 0.172062
R9342 DVDD.n9354 DVDD.n119 0.167884
R9343 DVDD.n9561 DVDD.n213 0.16731
R9344 DVDD.n9579 DVDD.n192 0.16731
R9345 DVDD DVDD.n229 0.165645
R9346 DVDD DVDD.n422 0.165645
R9347 DVDD.n747 DVDD.n746 0.164201
R9348 DVDD.n8836 DVDD.n8835 0.164201
R9349 DVDD.n9634 DVDD.n9633 0.164201
R9350 DVDD.n3703 DVDD.n3702 0.164201
R9351 DVDD.n9070 DVDD.n9018 0.164201
R9352 DVDD.n9106 DVDD.n9074 0.164201
R9353 DVDD.n4114 DVDD.n540 0.164201
R9354 DVDD.n4275 DVDD.n4223 0.164201
R9355 DVDD.n4996 DVDD.n4995 0.164201
R9356 DVDD.n4953 DVDD.n4950 0.164201
R9357 DVDD.n9474 DVDD.n287 0.164201
R9358 DVDD.n4371 DVDD.n265 0.164201
R9359 DVDD.n5215 DVDD.n5161 0.164201
R9360 DVDD.n9298 DVDD.n451 0.164201
R9361 DVDD.n9302 DVDD.n9301 0.164201
R9362 DVDD.n6850 DVDD.n6798 0.164201
R9363 DVDD.n8702 DVDD.n1001 0.15215
R9364 DVDD.n4695 DVDD.n4694 0.150736
R9365 DVDD.n5219 DVDD.n5218 0.150736
R9366 DVDD.n5264 DVDD.n5262 0.150736
R9367 DVDD.n5339 DVDD.n5338 0.150736
R9368 DVDD.n8009 DVDD.n1813 0.13721
R9369 DVDD.n7960 DVDD.n7959 0.13721
R9370 DVDD.n8204 DVDD 0.130618
R9371 DVDD.n8891 DVDD 0.130618
R9372 DVDD.n9700 DVDD 0.13017
R9373 DVDD.n1383 DVDD.n1374 0.119165
R9374 DVDD.n8490 DVDD.n1341 0.119165
R9375 DVDD.n8531 DVDD.n8523 0.114109
R9376 DVDD.n8549 DVDD.n1373 0.114108
R9377 DVDD.n7505 DVDD.n7070 0.113915
R9378 DVDD.n5249 DVDD.n4545 0.113652
R9379 DVDD.n4707 DVDD.n4625 0.113565
R9380 DVDD.n291 DVDD.n289 0.110634
R9381 DVDD.n254 DVDD.n240 0.110634
R9382 DVDD.n9321 DVDD.n9320 0.110634
R9383 DVDD.n5299 DVDD.n2957 0.110634
R9384 DVDD.n4107 DVDD.n3998 0.110634
R9385 DVDD.n4211 DVDD.n4210 0.110634
R9386 DVDD.n8787 DVDD.n8786 0.110634
R9387 DVDD.n3588 DVDD.n3587 0.110634
R9388 DVDD DVDD.n9700 0.101194
R9389 DVDD DVDD.n8204 0.10093
R9390 DVDD DVDD.n8891 0.10093
R9391 DVDD.n7500 DVDD.n7070 0.0901335
R9392 DVDD.n4707 DVDD.n4611 0.0896854
R9393 DVDD.n4760 DVDD.n4545 0.0896255
R9394 DVDD.n3807 DVDD.n3804 0.0842992
R9395 DVDD.n6154 DVDD.n4279 0.0842992
R9396 DVDD.n4376 DVDD.n4375 0.0842992
R9397 DVDD.n6855 DVDD.n6853 0.0842992
R9398 DVDD.n5377 DVDD.n5376 0.0775669
R9399 DVDD.n8707 DVDD.n905 0.0642795
R9400 DVDD.n4133 DVDD.n4132 0.0642795
R9401 DVDD.n9493 DVDD.n9492 0.0642795
R9402 DVDD.n9408 DVDD.n392 0.0642795
R9403 DVDD.n8751 DVDD.n8750 0.0642795
R9404 DVDD.n8705 DVDD.n8704 0.0642795
R9405 DVDD.n9598 DVDD.n9597 0.0642795
R9406 DVDD.n5270 DVDD.n4519 0.0642795
R9407 DVDD.n8004 DVDD 0.0638222
R9408 DVDD.n7946 DVDD 0.0638222
R9409 DVDD.n6599 DVDD 0.0638222
R9410 DVDD.n8171 DVDD 0.0638222
R9411 DVDD.n6393 DVDD 0.0638222
R9412 DVDD.n8665 DVDD.n8664 0.0632165
R9413 DVDD.n6773 DVDD.n6772 0.0632165
R9414 DVDD.n7026 DVDD.n7025 0.0621535
R9415 DVDD.n7549 DVDD.n7509 0.0621535
R9416 DVDD.n8055 DVDD.n1865 0.0621535
R9417 DVDD.n2284 DVDD.n1661 0.0621535
R9418 DVDD.n7779 DVDD.n1599 0.0621535
R9419 DVDD.n2387 DVDD.n1532 0.0621535
R9420 DVDD.n8659 DVDD.n8658 0.0621535
R9421 DVDD.n8656 DVDD.n8655 0.0621535
R9422 DVDD.n8653 DVDD.n8652 0.0621535
R9423 DVDD.n6767 DVDD.n2572 0.0621535
R9424 DVDD.n7004 DVDD.n2486 0.0621535
R9425 DVDD.n7591 DVDD.n2488 0.0621535
R9426 DVDD.n7687 DVDD.n2343 0.0610769
R9427 DVDD.n7729 DVDD.n7728 0.0610769
R9428 DVDD.n5268 DVDD.n5267 0.0602047
R9429 DVDD.n8876 DVDD.n660 0.0563
R9430 DVDD.n8872 DVDD.n660 0.0563
R9431 DVDD.n8872 DVDD.n8871 0.0563
R9432 DVDD.n8871 DVDD.n8870 0.0563
R9433 DVDD.n8870 DVDD.n662 0.0563
R9434 DVDD.n8866 DVDD.n662 0.0563
R9435 DVDD.n8866 DVDD.n8865 0.0563
R9436 DVDD.n8865 DVDD.n8864 0.0563
R9437 DVDD.n8864 DVDD.n664 0.0563
R9438 DVDD.n8860 DVDD.n664 0.0563
R9439 DVDD.n8860 DVDD.n8859 0.0563
R9440 DVDD.n8859 DVDD.n8858 0.0563
R9441 DVDD.n8858 DVDD.n666 0.0563
R9442 DVDD.n8854 DVDD.n666 0.0563
R9443 DVDD.n8854 DVDD.n8853 0.0563
R9444 DVDD.n8853 DVDD.n8852 0.0563
R9445 DVDD.n8852 DVDD.n668 0.0563
R9446 DVDD.n8848 DVDD.n668 0.0563
R9447 DVDD.n8848 DVDD.n8847 0.0563
R9448 DVDD.n8847 DVDD.n8846 0.0563
R9449 DVDD.n8846 DVDD.n670 0.0563
R9450 DVDD.n8842 DVDD.n670 0.0563
R9451 DVDD.n8842 DVDD.n8841 0.0563
R9452 DVDD.n8841 DVDD.n8840 0.0563
R9453 DVDD.n8840 DVDD.n672 0.0563
R9454 DVDD.n799 DVDD.n797 0.0563
R9455 DVDD.n800 DVDD.n799 0.0563
R9456 DVDD.n801 DVDD.n800 0.0563
R9457 DVDD.n801 DVDD.n795 0.0563
R9458 DVDD.n805 DVDD.n795 0.0563
R9459 DVDD.n806 DVDD.n805 0.0563
R9460 DVDD.n807 DVDD.n806 0.0563
R9461 DVDD.n830 DVDD.n15 0.0563
R9462 DVDD.n831 DVDD.n830 0.0563
R9463 DVDD.n832 DVDD.n831 0.0563
R9464 DVDD.n832 DVDD.n792 0.0563
R9465 DVDD.n836 DVDD.n792 0.0563
R9466 DVDD.n837 DVDD.n836 0.0563
R9467 DVDD.n8795 DVDD.n837 0.0563
R9468 DVDD.n8794 DVDD.n838 0.0563
R9469 DVDD.n950 DVDD.n949 0.0563
R9470 DVDD.n951 DVDD.n950 0.0563
R9471 DVDD.n8702 DVDD.n8701 0.0563
R9472 DVDD.n8701 DVDD.n1002 0.0563
R9473 DVDD.n1033 DVDD.n1002 0.0563
R9474 DVDD.n1033 DVDD.n1013 0.0563
R9475 DVDD.n3627 DVDD.n3626 0.0563
R9476 DVDD.n3626 DVDD.n3593 0.0563
R9477 DVDD.n3622 DVDD.n3593 0.0563
R9478 DVDD.n3622 DVDD.n3621 0.0563
R9479 DVDD.n3621 DVDD.n3620 0.0563
R9480 DVDD.n3620 DVDD.n3595 0.0563
R9481 DVDD.n3616 DVDD.n3595 0.0563
R9482 DVDD.n3616 DVDD.n3615 0.0563
R9483 DVDD.n3615 DVDD.n3614 0.0563
R9484 DVDD.n3614 DVDD.n3597 0.0563
R9485 DVDD.n3610 DVDD.n3597 0.0563
R9486 DVDD.n3610 DVDD.n3609 0.0563
R9487 DVDD.n3609 DVDD.n3608 0.0563
R9488 DVDD.n3608 DVDD.n3599 0.0563
R9489 DVDD.n3604 DVDD.n3599 0.0563
R9490 DVDD.n3604 DVDD.n3603 0.0563
R9491 DVDD.n3603 DVDD.n3602 0.0563
R9492 DVDD.n3602 DVDD.n3579 0.0563
R9493 DVDD.n3752 DVDD.n3579 0.0563
R9494 DVDD.n5614 DVDD.n5496 0.055969
R9495 DVDD.n7024 DVDD.n2523 0.055969
R9496 DVDD.n7548 DVDD.n7510 0.055969
R9497 DVDD.n5466 DVDD.n4473 0.055969
R9498 DVDD.n7508 DVDD.n7031 0.0553109
R9499 DVDD.n807 DVDD.n9 0.05315
R9500 DVDD.n809 DVDD.n8 0.05315
R9501 DVDD.n811 DVDD.n10 0.05315
R9502 DVDD.n813 DVDD.n7 0.05315
R9503 DVDD.n815 DVDD.n11 0.05315
R9504 DVDD.n817 DVDD.n6 0.05315
R9505 DVDD.n819 DVDD.n12 0.05315
R9506 DVDD.n821 DVDD.n5 0.05315
R9507 DVDD.n823 DVDD.n13 0.05315
R9508 DVDD.n825 DVDD.n4 0.05315
R9509 DVDD.n9692 DVDD.n14 0.05315
R9510 DVDD.n5910 DVDD.n5908 0.0515891
R9511 DVDD.n9563 DVDD.n223 0.0515849
R9512 DVDD.n111 DVDD.n103 0.0515849
R9513 DVDD.n200 DVDD.n187 0.0515835
R9514 DVDD.n8789 DVDD.n838 0.05135
R9515 DVDD.n8790 DVDD.n86 0.05135
R9516 DVDD.n8779 DVDD.n8778 0.05135
R9517 DVDD.n8777 DVDD.n90 0.05135
R9518 DVDD.n8774 DVDD.n8773 0.05135
R9519 DVDD.n840 DVDD.n115 0.05135
R9520 DVDD.n924 DVDD.n851 0.05135
R9521 DVDD.n926 DVDD.n854 0.05135
R9522 DVDD.n943 DVDD.n929 0.05135
R9523 DVDD.n944 DVDD.n868 0.05135
R9524 DVDD.n946 DVDD.n923 0.05135
R9525 DVDD.n122 DVDD.n103 0.0498479
R9526 DVDD.n2421 DVDD.n2405 0.049839
R9527 DVDD.n2421 DVDD.n2420 0.049839
R9528 DVDD.n2420 DVDD.n2406 0.049839
R9529 DVDD.n2415 DVDD.n2407 0.049839
R9530 DVDD.n2415 DVDD.n2414 0.049839
R9531 DVDD.n2414 DVDD.n2408 0.049839
R9532 DVDD.n2444 DVDD.n2428 0.049839
R9533 DVDD.n2444 DVDD.n2443 0.049839
R9534 DVDD.n2443 DVDD.n2429 0.049839
R9535 DVDD.n2438 DVDD.n2430 0.049839
R9536 DVDD.n2438 DVDD.n2437 0.049839
R9537 DVDD.n2437 DVDD.n2431 0.049839
R9538 DVDD.n7674 DVDD.n7661 0.049839
R9539 DVDD.n7662 DVDD.n7661 0.049839
R9540 DVDD.n7663 DVDD.n7662 0.049839
R9541 DVDD.n7670 DVDD.n7669 0.049839
R9542 DVDD.n7669 DVDD.n7668 0.049839
R9543 DVDD.n7668 DVDD.n7667 0.049839
R9544 DVDD.n1873 DVDD.n1869 0.049839
R9545 DVDD.n1869 DVDD.n1868 0.049839
R9546 DVDD.n1868 DVDD.n1867 0.049839
R9547 DVDD.n1881 DVDD.n1880 0.049839
R9548 DVDD.n9563 DVDD.n220 0.0497891
R9549 DVDD.n5910 DVDD.n5907 0.0497849
R9550 DVDD.n200 DVDD.n188 0.0497849
R9551 DVDD.n3749 DVDD.n3748 0.04955
R9552 DVDD.n3747 DVDD.n1039 0.04955
R9553 DVDD.n3744 DVDD.n3743 0.04955
R9554 DVDD.n3633 DVDD.n3584 0.04955
R9555 DVDD.n3632 DVDD.n1053 0.04955
R9556 DVDD.n3629 DVDD.n3628 0.04955
R9557 DVDD.n1879 DVDD.n1878 0.0491
R9558 DVDD.n8171 DVDD 0.0487259
R9559 DVDD.n8004 DVDD 0.0487259
R9560 DVDD.n7946 DVDD 0.0487259
R9561 DVDD.n6599 DVDD 0.0487259
R9562 DVDD.n6393 DVDD 0.0487259
R9563 DVDD.n4628 DVDD.n4568 0.0480684
R9564 DVDD.n744 DVDD.n743 0.0466307
R9565 DVDD.n951 DVDD.n872 0.04595
R9566 DVDD.n955 DVDD.n954 0.04595
R9567 DVDD.n978 DVDD.n956 0.04595
R9568 DVDD.n979 DVDD.n884 0.04595
R9569 DVDD.n981 DVDD.n886 0.04595
R9570 DVDD.n983 DVDD.n350 0.04595
R9571 DVDD.n985 DVDD.n892 0.04595
R9572 DVDD.n987 DVDD.n895 0.04595
R9573 DVDD.n989 DVDD.n920 0.04595
R9574 DVDD.n994 DVDD.n992 0.04595
R9575 DVDD.n993 DVDD.n908 0.04595
R9576 DVDD.n7348 DVDD.n7347 0.0450718
R9577 DVDD.n7356 DVDD.n7354 0.0450718
R9578 DVDD.n8620 DVDD.n1333 0.0450718
R9579 DVDD.n1327 DVDD.n1323 0.0450718
R9580 DVDD.n1398 DVDD.n1396 0.0450718
R9581 DVDD.n1404 DVDD.n1402 0.0450718
R9582 DVDD.n8519 DVDD.n8517 0.0450718
R9583 DVDD.n8537 DVDD.n8536 0.0450718
R9584 DVDD.n4879 DVDD.n4878 0.0450675
R9585 DVDD.n5159 DVDD.n4569 0.0450675
R9586 DVDD.n9015 DVDD.n547 0.0450675
R9587 DVDD.n725 DVDD.n724 0.0450675
R9588 DVDD.n8454 DVDD.n8446 0.0442838
R9589 DVDD.n8455 DVDD.n8454 0.0442838
R9590 DVDD.n8456 DVDD.n8455 0.0442838
R9591 DVDD.n8456 DVDD.n1338 0.0442838
R9592 DVDD.n8460 DVDD.n1338 0.0442838
R9593 DVDD.n8461 DVDD.n8460 0.0442838
R9594 DVDD.n8462 DVDD.n8461 0.0442838
R9595 DVDD.n8462 DVDD.n1445 0.0442838
R9596 DVDD.n7351 DVDD.n7349 0.0442838
R9597 DVDD.n7352 DVDD.n7351 0.0442838
R9598 DVDD.n7357 DVDD.n7355 0.0442838
R9599 DVDD.n7355 DVDD.n1335 0.0442838
R9600 DVDD.n1332 DVDD.n1329 0.0442838
R9601 DVDD.n8623 DVDD.n1329 0.0442838
R9602 DVDD.n1325 DVDD.n1324 0.0442838
R9603 DVDD.n8626 DVDD.n1325 0.0442838
R9604 DVDD.n8390 DVDD.n1494 0.0442838
R9605 DVDD.n8394 DVDD.n1494 0.0442838
R9606 DVDD.n8395 DVDD.n8394 0.0442838
R9607 DVDD.n8396 DVDD.n8395 0.0442838
R9608 DVDD.n8396 DVDD.n1492 0.0442838
R9609 DVDD.n8400 DVDD.n1492 0.0442838
R9610 DVDD.n8401 DVDD.n8400 0.0442838
R9611 DVDD.n8402 DVDD.n8401 0.0442838
R9612 DVDD.n8412 DVDD.n8411 0.0442838
R9613 DVDD.n8411 DVDD.n8410 0.0442838
R9614 DVDD.n8410 DVDD.n1377 0.0442838
R9615 DVDD.n8585 DVDD.n1377 0.0442838
R9616 DVDD.n8585 DVDD.n1378 0.0442838
R9617 DVDD.n8581 DVDD.n1378 0.0442838
R9618 DVDD.n8581 DVDD.n8580 0.0442838
R9619 DVDD.n8580 DVDD.n8579 0.0442838
R9620 DVDD.n8469 DVDD.n1443 0.0442838
R9621 DVDD.n8473 DVDD.n1443 0.0442838
R9622 DVDD.n8474 DVDD.n8473 0.0442838
R9623 DVDD.n8475 DVDD.n8474 0.0442838
R9624 DVDD.n8475 DVDD.n1441 0.0442838
R9625 DVDD.n8479 DVDD.n1441 0.0442838
R9626 DVDD.n8480 DVDD.n8479 0.0442838
R9627 DVDD.n8481 DVDD.n8480 0.0442838
R9628 DVDD.n8487 DVDD.n8486 0.0442838
R9629 DVDD.n8486 DVDD.n8485 0.0442838
R9630 DVDD.n8485 DVDD.n1344 0.0442838
R9631 DVDD.n8614 DVDD.n1344 0.0442838
R9632 DVDD.n8614 DVDD.n1345 0.0442838
R9633 DVDD.n8610 DVDD.n1345 0.0442838
R9634 DVDD.n8610 DVDD.n8609 0.0442838
R9635 DVDD.n8609 DVDD.n8608 0.0442838
R9636 DVDD.n8571 DVDD.n8570 0.0442838
R9637 DVDD.n8570 DVDD.n8569 0.0442838
R9638 DVDD.n8569 DVDD.n1385 0.0442838
R9639 DVDD.n8565 DVDD.n1385 0.0442838
R9640 DVDD.n8565 DVDD.n8564 0.0442838
R9641 DVDD.n8564 DVDD.n8563 0.0442838
R9642 DVDD.n8563 DVDD.n1387 0.0442838
R9643 DVDD.n8559 DVDD.n1387 0.0442838
R9644 DVDD.n8553 DVDD.n1389 0.0442838
R9645 DVDD.n8553 DVDD.n8552 0.0442838
R9646 DVDD.n8552 DVDD.n8551 0.0442838
R9647 DVDD.n8551 DVDD.n1373 0.0442838
R9648 DVDD.n8527 DVDD.n8525 0.0442838
R9649 DVDD.n8528 DVDD.n8527 0.0442838
R9650 DVDD.n8529 DVDD.n8528 0.0442838
R9651 DVDD.n8529 DVDD.n8523 0.0442838
R9652 DVDD.n1400 DVDD.n1399 0.0442838
R9653 DVDD.n8546 DVDD.n1399 0.0442838
R9654 DVDD.n8515 DVDD.n1405 0.0442838
R9655 DVDD.n8543 DVDD.n1405 0.0442838
R9656 DVDD.n8521 DVDD.n8520 0.0442838
R9657 DVDD.n8539 DVDD.n8521 0.0442838
R9658 DVDD.n8535 DVDD.n8534 0.0442838
R9659 DVDD.n8534 DVDD.n8532 0.0442838
R9660 DVDD.n7210 DVDD.n7031 0.0437872
R9661 DVDD.n7510 DVDD.n2506 0.0433572
R9662 DVDD.n2551 DVDD.n2523 0.0433572
R9663 DVDD.n5508 DVDD.n5496 0.0433572
R9664 DVDD.n5378 DVDD.n4473 0.0433572
R9665 DVDD DVDD.t31 0.0375588
R9666 DVDD DVDD.t37 0.0375588
R9667 DVDD DVDD.t6 0.0375588
R9668 DVDD DVDD.t25 0.0375588
R9669 DVDD.n8888 DVDD.n655 0.0349444
R9670 DVDD.n8884 DVDD.n655 0.0349444
R9671 DVDD.n8884 DVDD.n8883 0.0349444
R9672 DVDD.n8883 DVDD.n8882 0.0349444
R9673 DVDD.n8882 DVDD.n658 0.0349444
R9674 DVDD.n8878 DVDD.n658 0.0349444
R9675 DVDD.n8878 DVDD.n8877 0.0349444
R9676 DVDD.n1500 DVDD.n1305 0.0345541
R9677 DVDD.n8642 DVDD.n8641 0.0345541
R9678 DVDD.n8448 DVDD.n8446 0.0337432
R9679 DVDD.n8468 DVDD.n1445 0.0337432
R9680 DVDD.n8390 DVDD.n8389 0.0337432
R9681 DVDD.n8402 DVDD.n1489 0.0337432
R9682 DVDD.n8412 DVDD.n1489 0.0337432
R9683 DVDD.n8579 DVDD.n1381 0.0337432
R9684 DVDD.n8469 DVDD.n8468 0.0337432
R9685 DVDD.n8481 DVDD.n1438 0.0337432
R9686 DVDD.n8487 DVDD.n1438 0.0337432
R9687 DVDD.n8608 DVDD.n1348 0.0337432
R9688 DVDD.n8571 DVDD.n1381 0.0337432
R9689 DVDD.n8559 DVDD.n8558 0.0337432
R9690 DVDD.n8558 DVDD.n1389 0.0337432
R9691 DVDD.n8525 DVDD.n1348 0.0337432
R9692 DVDD.n2342 DVDD.n2335 0.0329742
R9693 DVDD.n7727 DVDD.n7726 0.0329742
R9694 DVDD.n8695 DVDD.n1007 0.03245
R9695 DVDD.n8695 DVDD.n8690 0.03245
R9696 DVDD.n8690 DVDD.n214 0.03245
R9697 DVDD.n8678 DVDD.n217 0.03245
R9698 DVDD.n8678 DVDD.n1045 0.03245
R9699 DVDD.n8674 DVDD.n1045 0.03245
R9700 DVDD.n6318 DVDD.n3869 0.03245
R9701 DVDD.n6318 DVDD.n6317 0.03245
R9702 DVDD.n6317 DVDD.n3872 0.03245
R9703 DVDD.n6307 DVDD.n3880 0.03245
R9704 DVDD.n6307 DVDD.n6306 0.03245
R9705 DVDD.n6306 DVDD.n6238 0.03245
R9706 DVDD.n6870 DVDD.n2794 0.03245
R9707 DVDD.n6870 DVDD.n2790 0.03245
R9708 DVDD.n6880 DVDD.n2790 0.03245
R9709 DVDD.n6884 DVDD.n2781 0.03245
R9710 DVDD.n6896 DVDD.n2781 0.03245
R9711 DVDD.n6896 DVDD.n2779 0.03245
R9712 DVDD.n180 DVDD.n176 0.03245
R9713 DVDD.n9582 DVDD.n176 0.03245
R9714 DVDD.n9582 DVDD.n177 0.03245
R9715 DVDD.n400 DVDD.n399 0.03245
R9716 DVDD.n9404 DVDD.n400 0.03245
R9717 DVDD.n9404 DVDD.n397 0.03245
R9718 DVDD.n5276 DVDD.n4513 0.03245
R9719 DVDD.n5280 DVDD.n4513 0.03245
R9720 DVDD.n5280 DVDD.n225 0.03245
R9721 DVDD.n2911 DVDD.n224 0.03245
R9722 DVDD.n2914 DVDD.n2911 0.03245
R9723 DVDD.n2914 DVDD.n2908 0.03245
R9724 DVDD.n440 DVDD.n413 0.03245
R9725 DVDD.n9357 DVDD.n413 0.03245
R9726 DVDD.n9357 DVDD.n414 0.03245
R9727 DVDD.n9352 DVDD.n9351 0.03245
R9728 DVDD.n9351 DVDD.n140 0.03245
R9729 DVDD.n9603 DVDD.n140 0.03245
R9730 DVDD.n8727 DVDD.n8724 0.03245
R9731 DVDD.n8731 DVDD.n8727 0.03245
R9732 DVDD.n8731 DVDD.n8728 0.03245
R9733 DVDD.n900 DVDD.n899 0.03245
R9734 DVDD.n8711 DVDD.n900 0.03245
R9735 DVDD.n8711 DVDD.n901 0.03245
R9736 DVDD.n98 DVDD.n95 0.03245
R9737 DVDD.n9619 DVDD.n95 0.03245
R9738 DVDD.n9619 DVDD.n9618 0.03245
R9739 DVDD.n859 DVDD.n858 0.03245
R9740 DVDD.n8758 DVDD.n859 0.03245
R9741 DVDD.n8758 DVDD.n8757 0.03245
R9742 DVDD.n6592 DVDD.n6486 0.0306622
R9743 DVDD.n6588 DVDD.n6486 0.0306622
R9744 DVDD.n3466 DVDD.n3465 0.0306622
R9745 DVDD.n3465 DVDD.n3422 0.0306622
R9746 DVDD.n3461 DVDD.n3422 0.0306622
R9747 DVDD.n3461 DVDD.n3460 0.0306622
R9748 DVDD.n3460 DVDD.n3459 0.0306622
R9749 DVDD.n3459 DVDD.n3424 0.0306622
R9750 DVDD.n3455 DVDD.n3424 0.0306622
R9751 DVDD.n3455 DVDD.n3454 0.0306622
R9752 DVDD.n3454 DVDD.n3453 0.0306622
R9753 DVDD.n3453 DVDD.n3426 0.0306622
R9754 DVDD.n3449 DVDD.n3426 0.0306622
R9755 DVDD.n3449 DVDD.n3448 0.0306622
R9756 DVDD.n3448 DVDD.n3447 0.0306622
R9757 DVDD.n3447 DVDD.n3428 0.0306622
R9758 DVDD.n3443 DVDD.n3428 0.0306622
R9759 DVDD.n6386 DVDD.n3552 0.0306622
R9760 DVDD.n6382 DVDD.n3552 0.0306622
R9761 DVDD.n3801 DVDD.n3800 0.0306622
R9762 DVDD.n3800 DVDD.n3799 0.0306622
R9763 DVDD.n3799 DVDD.n3753 0.0306622
R9764 DVDD.n3795 DVDD.n3753 0.0306622
R9765 DVDD.n3795 DVDD.n3794 0.0306622
R9766 DVDD.n3794 DVDD.n3793 0.0306622
R9767 DVDD.n3793 DVDD.n3755 0.0306622
R9768 DVDD.n3789 DVDD.n3755 0.0306622
R9769 DVDD.n3789 DVDD.n3788 0.0306622
R9770 DVDD.n3788 DVDD.n3787 0.0306622
R9771 DVDD.n3787 DVDD.n3757 0.0306622
R9772 DVDD.n3783 DVDD.n3757 0.0306622
R9773 DVDD.n3783 DVDD.n3782 0.0306622
R9774 DVDD.n3782 DVDD.n3781 0.0306622
R9775 DVDD.n3781 DVDD.n3759 0.0306622
R9776 DVDD.n3777 DVDD.n3759 0.0306622
R9777 DVDD.n3777 DVDD.n3776 0.0306622
R9778 DVDD.n3776 DVDD.n3775 0.0306622
R9779 DVDD.n3775 DVDD.n3761 0.0306622
R9780 DVDD.n3771 DVDD.n3761 0.0306622
R9781 DVDD.n3771 DVDD.n3770 0.0306622
R9782 DVDD.n3770 DVDD.n3769 0.0306622
R9783 DVDD.n3769 DVDD.n3763 0.0306622
R9784 DVDD.n3765 DVDD.n3763 0.0306622
R9785 DVDD.n3765 DVDD.n3764 0.0306622
R9786 DVDD.n8618 DVDD.t0 0.028625
R9787 DVDD.n8619 DVDD.n8618 0.028625
R9788 DVDD.n8542 DVDD.n1372 0.028625
R9789 DVDD.n1372 DVDD.t0 0.028625
R9790 DVDD.n8893 DVDD.n8888 0.0284117
R9791 DVDD.n8698 DVDD.n8697 0.0284
R9792 DVDD.n8672 DVDD.n1046 0.0284
R9793 DVDD.n8747 DVDD.n8746 0.0284
R9794 DVDD.n917 DVDD.n898 0.0284
R9795 DVDD.n6326 DVDD.n6325 0.0284
R9796 DVDD.n6304 DVDD.n6239 0.0284
R9797 DVDD.n6867 DVDD.n2796 0.0284
R9798 DVDD.n6894 DVDD.n2783 0.0284
R9799 DVDD.n178 DVDD.n155 0.0284
R9800 DVDD.n395 DVDD.n388 0.0284
R9801 DVDD.n5274 DVDD.n4515 0.0284
R9802 DVDD.n6780 DVDD.n6779 0.0284
R9803 DVDD.n9314 DVDD.n9313 0.0284
R9804 DVDD.n9601 DVDD.n139 0.0284
R9805 DVDD.n841 DVDD.n83 0.0284
R9806 DVDD.n8755 DVDD.n863 0.0284
R9807 DVDD.n8673 DVDD.n1048 0.027725
R9808 DVDD.n8725 DVDD.n876 0.027725
R9809 DVDD.n6320 DVDD.n3866 0.027725
R9810 DVDD.n2795 DVDD.n2793 0.027725
R9811 DVDD.n179 DVDD.n164 0.027725
R9812 DVDD.n2912 DVDD.n2907 0.027725
R9813 DVDD.n9605 DVDD.n9604 0.027725
R9814 DVDD.n8756 DVDD.n857 0.027725
R9815 DVDD.n8691 DVDD.n1005 0.027275
R9816 DVDD.n8708 DVDD.n903 0.027275
R9817 DVDD.n6244 DVDD.n6242 0.027275
R9818 DVDD.n6899 DVDD.n2778 0.027275
R9819 DVDD.n9407 DVDD.n396 0.027275
R9820 DVDD.n5275 DVDD.n4514 0.027275
R9821 DVDD.n441 DVDD.n438 0.027275
R9822 DVDD.n97 DVDD.n96 0.027275
R9823 DVDD.n7682 DVDD.n7681 0.026913
R9824 DVDD.n7684 DVDD.n2358 0.026913
R9825 DVDD.n2366 DVDD.n2365 0.026913
R9826 DVDD.n2368 DVDD.n2363 0.026913
R9827 DVDD.n7738 DVDD.n7737 0.026913
R9828 DVDD.n7732 DVDD.n7731 0.026913
R9829 DVDD.n7734 DVDD.n2340 0.026913
R9830 DVDD.n8389 DVDD.n8388 0.0268514
R9831 DVDD.n8448 DVDD.n1326 0.0268514
R9832 DVDD.n8418 DVDD.n1465 0.0263511
R9833 DVDD.n8418 DVDD.n1466 0.0263511
R9834 DVDD.n8426 DVDD.n8424 0.0263511
R9835 DVDD.n8426 DVDD.n8425 0.0263511
R9836 DVDD.n8431 DVDD.n1455 0.0263511
R9837 DVDD.n1455 DVDD.n1454 0.0263511
R9838 DVDD.n8436 DVDD.n1450 0.0263511
R9839 DVDD.n1450 DVDD.n1449 0.0263511
R9840 DVDD.n1487 DVDD.n1470 0.0263511
R9841 DVDD.n1487 DVDD.n1472 0.0263511
R9842 DVDD.n1417 DVDD.n1414 0.0263511
R9843 DVDD.n1419 DVDD.n1414 0.0263511
R9844 DVDD.n1426 DVDD.n1423 0.0263511
R9845 DVDD.n1427 DVDD.n1426 0.0263511
R9846 DVDD.n1434 DVDD.n1431 0.0263511
R9847 DVDD.n1435 DVDD.n1434 0.0263511
R9848 DVDD.n1482 DVDD.n1476 0.0263511
R9849 DVDD.n1482 DVDD.n1478 0.0263511
R9850 DVDD.n1411 DVDD.n1408 0.0263511
R9851 DVDD.n8509 DVDD.n1408 0.0263511
R9852 DVDD.n8594 DVDD.n1366 0.0263511
R9853 DVDD.n8594 DVDD.n1367 0.0263511
R9854 DVDD.n8599 DVDD.n1357 0.0263511
R9855 DVDD.n8599 DVDD.n1358 0.0263511
R9856 DVDD.n200 DVDD.n184 0.0257401
R9857 DVDD.n104 DVDD.n103 0.0255962
R9858 DVDD.n9563 DVDD.n227 0.0255962
R9859 DVDD.n5646 DVDD.n5644 0.0255952
R9860 DVDD.n8696 DVDD.n1006 0.025475
R9861 DVDD.n8713 DVDD.n8712 0.025475
R9862 DVDD.n6305 DVDD.n3879 0.025475
R9863 DVDD.n6895 DVDD.n2782 0.025475
R9864 DVDD.n9403 DVDD.n9402 0.025475
R9865 DVDD.n5282 DVDD.n4510 0.025475
R9866 DVDD.n442 DVDD.n412 0.025475
R9867 DVDD.n9621 DVDD.n93 0.025475
R9868 DVDD.n2418 DVDD.n2406 0.0251695
R9869 DVDD.n2412 DVDD.n2408 0.0251695
R9870 DVDD.n2441 DVDD.n2429 0.0251695
R9871 DVDD.n2435 DVDD.n2431 0.0251695
R9872 DVDD.n7672 DVDD.n7663 0.0251695
R9873 DVDD.n7667 DVDD.n7666 0.0251695
R9874 DVDD.n1875 DVDD.n1867 0.0251695
R9875 DVDD.n1878 DVDD.n1877 0.0251695
R9876 DVDD.n1882 DVDD.n1881 0.0251695
R9877 DVDD.n1880 DVDD.n1879 0.0251695
R9878 DVDD.n1877 DVDD.n1876 0.0251695
R9879 DVDD.n7671 DVDD.n7670 0.0251695
R9880 DVDD.n2440 DVDD.n2430 0.0251695
R9881 DVDD.n2417 DVDD.n2407 0.0251695
R9882 DVDD.n1873 DVDD.n1872 0.0251695
R9883 DVDD.n7675 DVDD.n7674 0.0251695
R9884 DVDD.n2446 DVDD.n2428 0.0251695
R9885 DVDD.n2423 DVDD.n2405 0.0251695
R9886 DVDD.n9563 DVDD.n9562 0.0247655
R9887 DVDD.n5645 DVDD.n5644 0.0247646
R9888 DVDD.n200 DVDD.n183 0.0247619
R9889 DVDD.n105 DVDD.n103 0.0247609
R9890 DVDD.n7362 DVDD.n7344 0.0243462
R9891 DVDD.n7344 DVDD.n1306 0.0243462
R9892 DVDD.n1312 DVDD.n1311 0.0243462
R9893 DVDD.n8636 DVDD.n1312 0.0243462
R9894 DVDD.n1320 DVDD.n1319 0.0243462
R9895 DVDD.n8631 DVDD.n1320 0.0243462
R9896 DVDD.n1047 DVDD.n1044 0.023675
R9897 DVDD.n8726 DVDD.n881 0.023675
R9898 DVDD.n6319 DVDD.n3868 0.023675
R9899 DVDD.n6872 DVDD.n6871 0.023675
R9900 DVDD.n9584 DVDD.n174 0.023675
R9901 DVDD.n2913 DVDD.n2900 0.023675
R9902 DVDD.n9349 DVDD.n138 0.023675
R9903 DVDD.n8760 DVDD.n8759 0.023675
R9904 DVDD.n742 DVDD.n649 0.0227991
R9905 DVDD.n740 DVDD.n647 0.0227991
R9906 DVDD.n738 DVDD.n650 0.0227991
R9907 DVDD.n736 DVDD.n646 0.0227991
R9908 DVDD.n734 DVDD.n651 0.0227991
R9909 DVDD.n732 DVDD.n645 0.0227991
R9910 DVDD.n730 DVDD.n652 0.0227991
R9911 DVDD.n728 DVDD.n644 0.0227991
R9912 DVDD.n726 DVDD.n653 0.0227991
R9913 DVDD.n654 DVDD.n643 0.0227991
R9914 DVDD.n8536 DVDD.n8535 0.0227859
R9915 DVDD.n8538 DVDD.n8537 0.0227859
R9916 DVDD.n8624 DVDD.n1323 0.0227859
R9917 DVDD.n1327 DVDD.n1324 0.0227859
R9918 DVDD.n8541 DVDD.n8517 0.0227859
R9919 DVDD.n8520 DVDD.n8519 0.0227859
R9920 DVDD.n8621 DVDD.n8620 0.0227859
R9921 DVDD.n1333 DVDD.n1332 0.0227859
R9922 DVDD.n8545 DVDD.n1402 0.0227859
R9923 DVDD.n8515 DVDD.n1404 0.0227859
R9924 DVDD.n7354 DVDD.n7353 0.0227859
R9925 DVDD.n7357 DVDD.n7356 0.0227859
R9926 DVDD.n8548 DVDD.n1396 0.0227859
R9927 DVDD.n1400 DVDD.n1398 0.0227859
R9928 DVDD.n7347 DVDD.n1497 0.0227859
R9929 DVDD.n7349 DVDD.n7348 0.0227859
R9930 DVDD.n9563 DVDD.n213 0.0227712
R9931 DVDD.n200 DVDD.n192 0.0227712
R9932 DVDD.n119 DVDD.n103 0.0227678
R9933 DVDD.n4706 DVDD.n4626 0.0224685
R9934 DVDD.n4702 DVDD.n4626 0.0224685
R9935 DVDD.n4702 DVDD.n4701 0.0224685
R9936 DVDD.n4701 DVDD.n4700 0.0224685
R9937 DVDD.n4700 DVDD.n4647 0.0224685
R9938 DVDD.n4696 DVDD.n4647 0.0224685
R9939 DVDD.n4696 DVDD.n4695 0.0224685
R9940 DVDD.n4694 DVDD.n4693 0.0224685
R9941 DVDD.n4693 DVDD.n4648 0.0224685
R9942 DVDD.n4689 DVDD.n4648 0.0224685
R9943 DVDD.n4689 DVDD.n4688 0.0224685
R9944 DVDD.n4688 DVDD.n4687 0.0224685
R9945 DVDD.n4687 DVDD.n4650 0.0224685
R9946 DVDD.n4683 DVDD.n4650 0.0224685
R9947 DVDD.n4683 DVDD.n4682 0.0224685
R9948 DVDD.n4682 DVDD.n4681 0.0224685
R9949 DVDD.n4681 DVDD.n4652 0.0224685
R9950 DVDD.n4677 DVDD.n4652 0.0224685
R9951 DVDD.n4677 DVDD.n4676 0.0224685
R9952 DVDD.n4676 DVDD.n4675 0.0224685
R9953 DVDD.n4675 DVDD.n4654 0.0224685
R9954 DVDD.n4671 DVDD.n4654 0.0224685
R9955 DVDD.n4671 DVDD.n4670 0.0224685
R9956 DVDD.n4670 DVDD.n4669 0.0224685
R9957 DVDD.n4669 DVDD.n4656 0.0224685
R9958 DVDD.n4665 DVDD.n4656 0.0224685
R9959 DVDD.n4665 DVDD.n4664 0.0224685
R9960 DVDD.n4664 DVDD.n4663 0.0224685
R9961 DVDD.n4663 DVDD.n4658 0.0224685
R9962 DVDD.n4659 DVDD.n4658 0.0224685
R9963 DVDD.n4659 DVDD.n4560 0.0224685
R9964 DVDD.n5218 DVDD.n4560 0.0224685
R9965 DVDD.n5221 DVDD.n5219 0.0224685
R9966 DVDD.n5222 DVDD.n5221 0.0224685
R9967 DVDD.n5223 DVDD.n5222 0.0224685
R9968 DVDD.n5223 DVDD.n4558 0.0224685
R9969 DVDD.n5227 DVDD.n4558 0.0224685
R9970 DVDD.n5228 DVDD.n5227 0.0224685
R9971 DVDD.n5229 DVDD.n5228 0.0224685
R9972 DVDD.n5251 DVDD.n4539 0.0224685
R9973 DVDD.n5255 DVDD.n4539 0.0224685
R9974 DVDD.n5256 DVDD.n5255 0.0224685
R9975 DVDD.n5257 DVDD.n5256 0.0224685
R9976 DVDD.n5257 DVDD.n4537 0.0224685
R9977 DVDD.n5261 DVDD.n4537 0.0224685
R9978 DVDD.n5262 DVDD.n5261 0.0224685
R9979 DVDD.n5264 DVDD.n5263 0.0224685
R9980 DVDD.n9378 DVDD.n9377 0.0224685
R9981 DVDD.n9379 DVDD.n9378 0.0224685
R9982 DVDD.n5268 DVDD.n4518 0.0224685
R9983 DVDD.n4518 DVDD.n4517 0.0224685
R9984 DVDD.n4517 DVDD.n4506 0.0224685
R9985 DVDD.n5288 DVDD.n4506 0.0224685
R9986 DVDD.n5309 DVDD.n4504 0.0224685
R9987 DVDD.n5313 DVDD.n4504 0.0224685
R9988 DVDD.n5314 DVDD.n5313 0.0224685
R9989 DVDD.n5315 DVDD.n5314 0.0224685
R9990 DVDD.n5315 DVDD.n4502 0.0224685
R9991 DVDD.n5319 DVDD.n4502 0.0224685
R9992 DVDD.n5320 DVDD.n5319 0.0224685
R9993 DVDD.n5321 DVDD.n5320 0.0224685
R9994 DVDD.n5321 DVDD.n4500 0.0224685
R9995 DVDD.n5325 DVDD.n4500 0.0224685
R9996 DVDD.n5326 DVDD.n5325 0.0224685
R9997 DVDD.n5327 DVDD.n5326 0.0224685
R9998 DVDD.n5327 DVDD.n4498 0.0224685
R9999 DVDD.n5331 DVDD.n4498 0.0224685
R10000 DVDD.n5332 DVDD.n5331 0.0224685
R10001 DVDD.n5333 DVDD.n5332 0.0224685
R10002 DVDD.n5333 DVDD.n4496 0.0224685
R10003 DVDD.n5337 DVDD.n4496 0.0224685
R10004 DVDD.n5338 DVDD.n5337 0.0224685
R10005 DVDD.n5340 DVDD.n5339 0.0224685
R10006 DVDD.n5341 DVDD.n5340 0.0224685
R10007 DVDD.n5341 DVDD.n4494 0.0224685
R10008 DVDD.n5345 DVDD.n4494 0.0224685
R10009 DVDD.n5346 DVDD.n5345 0.0224685
R10010 DVDD.n5347 DVDD.n5346 0.0224685
R10011 DVDD.n5347 DVDD.n4492 0.0224685
R10012 DVDD.n5351 DVDD.n4492 0.0224685
R10013 DVDD.n5352 DVDD.n5351 0.0224685
R10014 DVDD.n5353 DVDD.n5352 0.0224685
R10015 DVDD.n5353 DVDD.n4490 0.0224685
R10016 DVDD.n5357 DVDD.n4490 0.0224685
R10017 DVDD.n5358 DVDD.n5357 0.0224685
R10018 DVDD.n5359 DVDD.n5358 0.0224685
R10019 DVDD.n5359 DVDD.n4488 0.0224685
R10020 DVDD.n5363 DVDD.n4488 0.0224685
R10021 DVDD.n5364 DVDD.n5363 0.0224685
R10022 DVDD.n5365 DVDD.n5364 0.0224685
R10023 DVDD.n5365 DVDD.n4486 0.0224685
R10024 DVDD.n5369 DVDD.n4486 0.0224685
R10025 DVDD.n5370 DVDD.n5369 0.0224685
R10026 DVDD.n5371 DVDD.n5370 0.0224685
R10027 DVDD.n5371 DVDD.n4484 0.0224685
R10028 DVDD.n5375 DVDD.n4484 0.0224685
R10029 DVDD.n5376 DVDD.n5375 0.0224685
R10030 DVDD.n5472 DVDD.n5471 0.0224685
R10031 DVDD.n5473 DVDD.n5472 0.0224685
R10032 DVDD.n5639 DVDD.n5484 0.0224685
R10033 DVDD.n5635 DVDD.n5484 0.0224685
R10034 DVDD.n5635 DVDD.n5634 0.0224685
R10035 DVDD.n5634 DVDD.n5633 0.0224685
R10036 DVDD.n5633 DVDD.n5486 0.0224685
R10037 DVDD.n5629 DVDD.n5486 0.0224685
R10038 DVDD.n5629 DVDD.n5628 0.0224685
R10039 DVDD.n5628 DVDD.n5627 0.0224685
R10040 DVDD.n5627 DVDD.n5488 0.0224685
R10041 DVDD.n5623 DVDD.n5488 0.0224685
R10042 DVDD.n5623 DVDD.n5622 0.0224685
R10043 DVDD.n5622 DVDD.n5621 0.0224685
R10044 DVDD.n5621 DVDD.n5490 0.0224685
R10045 DVDD.n5617 DVDD.n5490 0.0224685
R10046 DVDD.n5617 DVDD.n5616 0.0224685
R10047 DVDD.n5612 DVDD.n5566 0.0224685
R10048 DVDD.n5608 DVDD.n5566 0.0224685
R10049 DVDD.n8699 DVDD.n905 0.0224685
R10050 DVDD.n8699 DVDD.n1004 0.0224685
R10051 DVDD.n1009 DVDD.n1004 0.0224685
R10052 DVDD.n8687 DVDD.n1009 0.0224685
R10053 DVDD.n4135 DVDD.n4133 0.0224685
R10054 DVDD.n4135 DVDD.n4134 0.0224685
R10055 DVDD.n4134 DVDD.n3976 0.0224685
R10056 DVDD.n4146 DVDD.n3976 0.0224685
R10057 DVDD.n9495 DVDD.n9493 0.0224685
R10058 DVDD.n9495 DVDD.n9494 0.0224685
R10059 DVDD.n9494 DVDD.n267 0.0224685
R10060 DVDD.n9506 DVDD.n267 0.0224685
R10061 DVDD.n5273 DVDD.n392 0.0224685
R10062 DVDD.n5273 DVDD.n4509 0.0224685
R10063 DVDD.n5283 DVDD.n4509 0.0224685
R10064 DVDD.n5283 DVDD.n2889 0.0224685
R10065 DVDD.n9626 DVDD.n46 0.0224685
R10066 DVDD.n9626 DVDD.n9625 0.0224685
R10067 DVDD.n9625 DVDD.n9624 0.0224685
R10068 DVDD.n9624 DVDD.n87 0.0224685
R10069 DVDD.n113 DVDD.n87 0.0224685
R10070 DVDD.n8764 DVDD.n113 0.0224685
R10071 DVDD.n8764 DVDD.n8763 0.0224685
R10072 DVDD.n8763 DVDD.n852 0.0224685
R10073 DVDD.n8752 DVDD.n852 0.0224685
R10074 DVDD.n8752 DVDD.n8751 0.0224685
R10075 DVDD.n8750 DVDD.n869 0.0224685
R10076 DVDD.n885 DVDD.n869 0.0224685
R10077 DVDD.n8737 DVDD.n885 0.0224685
R10078 DVDD.n8737 DVDD.n8736 0.0224685
R10079 DVDD.n8736 DVDD.n351 0.0224685
R10080 DVDD.n8717 DVDD.n351 0.0224685
R10081 DVDD.n8717 DVDD.n8716 0.0224685
R10082 DVDD.n8716 DVDD.n893 0.0224685
R10083 DVDD.n909 DVDD.n893 0.0224685
R10084 DVDD.n8705 DVDD.n909 0.0224685
R10085 DVDD.n8704 DVDD.n910 0.0224685
R10086 DVDD.n1014 DVDD.n910 0.0224685
R10087 DVDD.n1035 DVDD.n1014 0.0224685
R10088 DVDD.n8685 DVDD.n1035 0.0224685
R10089 DVDD.n8685 DVDD.n8684 0.0224685
R10090 DVDD.n8684 DVDD.n8683 0.0224685
R10091 DVDD.n8683 DVDD.n1036 0.0224685
R10092 DVDD.n1054 DVDD.n1036 0.0224685
R10093 DVDD.n8669 DVDD.n1054 0.0224685
R10094 DVDD.n8669 DVDD.n8668 0.0224685
R10095 DVDD.n8646 DVDD.n1297 0.0224685
R10096 DVDD.n8644 DVDD.n1297 0.0224685
R10097 DVDD.n9318 DVDD.n9317 0.0224685
R10098 DVDD.n9317 DVDD.n433 0.0224685
R10099 DVDD.n4527 DVDD.n433 0.0224685
R10100 DVDD.n4527 DVDD.n127 0.0224685
R10101 DVDD.n9615 DVDD.n127 0.0224685
R10102 DVDD.n9615 DVDD.n9614 0.0224685
R10103 DVDD.n9614 DVDD.n128 0.0224685
R10104 DVDD.n148 DVDD.n128 0.0224685
R10105 DVDD.n149 DVDD.n148 0.0224685
R10106 DVDD.n9598 DVDD.n149 0.0224685
R10107 DVDD.n9597 DVDD.n150 0.0224685
R10108 DVDD.n9588 DVDD.n150 0.0224685
R10109 DVDD.n9588 DVDD.n9587 0.0224685
R10110 DVDD.n9587 DVDD.n169 0.0224685
R10111 DVDD.n359 DVDD.n169 0.0224685
R10112 DVDD.n383 DVDD.n359 0.0224685
R10113 DVDD.n9417 DVDD.n383 0.0224685
R10114 DVDD.n9417 DVDD.n9416 0.0224685
R10115 DVDD.n9416 DVDD.n384 0.0224685
R10116 DVDD.n4519 DVDD.n384 0.0224685
R10117 DVDD.n5271 DVDD.n5270 0.0224685
R10118 DVDD.n5271 DVDD.n4507 0.0224685
R10119 DVDD.n5285 DVDD.n4507 0.0224685
R10120 DVDD.n5286 DVDD.n5285 0.0224685
R10121 DVDD.n5286 DVDD.n2896 0.0224685
R10122 DVDD.n6790 DVDD.n2896 0.0224685
R10123 DVDD.n6790 DVDD.n6789 0.0224685
R10124 DVDD.n6789 DVDD.n2897 0.0224685
R10125 DVDD.n2959 DVDD.n2897 0.0224685
R10126 DVDD.n6776 DVDD.n2959 0.0224685
R10127 DVDD.n8382 DVDD.n1502 0.0224685
R10128 DVDD.n8382 DVDD.n1501 0.0224685
R10129 DVDD.n7183 DVDD.n1304 0.0218559
R10130 DVDD.n8640 DVDD.n8639 0.0218559
R10131 DVDD.n3871 DVDD.n3870 0.0218
R10132 DVDD.n3881 DVDD.n3871 0.0218
R10133 DVDD.n6236 DVDD.n6235 0.0218
R10134 DVDD.n6237 DVDD.n6236 0.0218
R10135 DVDD.n6869 DVDD.n2789 0.0218
R10136 DVDD.n6881 DVDD.n2789 0.0218
R10137 DVDD.n6883 DVDD.n2780 0.0218
R10138 DVDD.n6897 DVDD.n2780 0.0218
R10139 DVDD.n9581 DVDD.n182 0.0218
R10140 DVDD.n9581 DVDD.n9580 0.0218
R10141 DVDD.n398 DVDD.n197 0.0218
R10142 DVDD.n9405 DVDD.n398 0.0218
R10143 DVDD.n8694 DVDD.n8693 0.0218
R10144 DVDD.n8693 DVDD.n230 0.0218
R10145 DVDD.n8677 DVDD.n233 0.0218
R10146 DVDD.n8677 DVDD.n8676 0.0218
R10147 DVDD.n5279 DVDD.n5278 0.0218
R10148 DVDD.n5279 DVDD.n236 0.0218
R10149 DVDD.n2909 DVDD.n238 0.0218
R10150 DVDD.n2915 DVDD.n2909 0.0218
R10151 DVDD.n9356 DVDD.n415 0.0218
R10152 DVDD.n9356 DVDD.n9355 0.0218
R10153 DVDD.n9353 DVDD.n9348 0.0218
R10154 DVDD.n9348 DVDD.n141 0.0218
R10155 DVDD.n8730 DVDD.n8729 0.0218
R10156 DVDD.n8730 DVDD.n194 0.0218
R10157 DVDD.n902 DVDD.n189 0.0218
R10158 DVDD.n8710 DVDD.n902 0.0218
R10159 DVDD.n101 DVDD.n100 0.0218
R10160 DVDD.n102 DVDD.n101 0.0218
R10161 DVDD.n860 DVDD.n421 0.0218
R10162 DVDD.n861 DVDD.n860 0.0218
R10163 DVDD.n8689 DVDD.n8688 0.021425
R10164 DVDD.n897 DVDD.n890 0.021425
R10165 DVDD.n6309 DVDD.n6308 0.021425
R10166 DVDD.n6887 DVDD.n6886 0.021425
R10167 DVDD.n9401 DVDD.n9400 0.021425
R10168 DVDD.n5281 DVDD.n4512 0.021425
R10169 DVDD.n9359 DVDD.n9358 0.021425
R10170 DVDD.n9620 DVDD.n94 0.021425
R10171 DVDD DVDD.n353 0.0213137
R10172 DVDD.n5229 DVDD.n4552 0.0212283
R10173 DVDD.n5231 DVDD.n4550 0.0212283
R10174 DVDD.n5233 DVDD.n4553 0.0212283
R10175 DVDD.n5235 DVDD.n4549 0.0212283
R10176 DVDD.n5237 DVDD.n4554 0.0212283
R10177 DVDD.n5239 DVDD.n4548 0.0212283
R10178 DVDD.n5241 DVDD.n4555 0.0212283
R10179 DVDD.n5243 DVDD.n4547 0.0212283
R10180 DVDD.n5248 DVDD.n4556 0.0212283
R10181 DVDD.n5247 DVDD.n4546 0.0212283
R10182 DVDD.n5250 DVDD.n4541 0.0212283
R10183 DVDD.n8465 DVDD.n8443 0.0205933
R10184 DVDD.n8443 DVDD.n8442 0.0205933
R10185 DVDD.n8492 DVDD.n1439 0.0205933
R10186 DVDD.n1439 DVDD.n1437 0.0205933
R10187 DVDD.n1350 DVDD.n1349 0.0205933
R10188 DVDD.n8603 DVDD.n1350 0.0205933
R10189 DVDD.n8405 DVDD.n1490 0.0205933
R10190 DVDD.n8407 DVDD.n1490 0.0205933
R10191 DVDD.n8576 DVDD.n8575 0.0205933
R10192 DVDD.n8575 DVDD.n8574 0.0205933
R10193 DVDD.n1392 DVDD.n1391 0.0205933
R10194 DVDD.n1394 DVDD.n1392 0.0205933
R10195 DVDD.n5263 DVDD.n429 0.0205197
R10196 DVDD.n4534 DVDD.n435 0.0205197
R10197 DVDD.n4532 DVDD.n4531 0.0205197
R10198 DVDD.n4530 DVDD.n4529 0.0205197
R10199 DVDD.n9362 DVDD.n408 0.0205197
R10200 DVDD.n9363 DVDD.n107 0.0205197
R10201 DVDD.n9365 DVDD.n130 0.0205197
R10202 DVDD.n9367 DVDD.n406 0.0205197
R10203 DVDD.n9371 DVDD.n9370 0.0205197
R10204 DVDD.n9373 DVDD.n9372 0.0205197
R10205 DVDD.n9374 DVDD.n147 0.0205197
R10206 DVDD.n7733 DVDD.n1972 0.0203425
R10207 DVDD.n7746 DVDD.n7745 0.0203425
R10208 DVDD.n2367 DVDD.n2235 0.0203425
R10209 DVDD.n7683 DVDD.n7680 0.0203425
R10210 DVDD.n229 DVDD 0.0202739
R10211 DVDD.n422 DVDD 0.0202739
R10212 DVDD.n4627 DVDD.n4614 0.0201654
R10213 DVDD.n4629 DVDD.n4623 0.0201654
R10214 DVDD.n4631 DVDD.n4615 0.0201654
R10215 DVDD.n4633 DVDD.n4622 0.0201654
R10216 DVDD.n4635 DVDD.n4616 0.0201654
R10217 DVDD.n4637 DVDD.n4621 0.0201654
R10218 DVDD.n4639 DVDD.n4617 0.0201654
R10219 DVDD.n4641 DVDD.n4620 0.0201654
R10220 DVDD.n4643 DVDD.n4618 0.0201654
R10221 DVDD.n4624 DVDD.n4619 0.0201654
R10222 DVDD.n4712 DVDD.n4706 0.0201654
R10223 DVDD.n5290 DVDD.n5289 0.019811
R10224 DVDD.n5291 DVDD.n2895 0.019811
R10225 DVDD.n5293 DVDD.n2899 0.019811
R10226 DVDD.n5304 DVDD.n5296 0.019811
R10227 DVDD.n5306 DVDD.n5305 0.019811
R10228 DVDD.n5307 DVDD.n2958 0.019811
R10229 DVDD.n721 DVDD.n720 0.0196339
R10230 DVDD.n705 DVDD.n704 0.0196339
R10231 DVDD.n699 DVDD.n590 0.0196339
R10232 DVDD.n699 DVDD.n698 0.0196339
R10233 DVDD.n698 DVDD.n697 0.0196339
R10234 DVDD.n697 DVDD.n690 0.0196339
R10235 DVDD.n693 DVDD.n690 0.0196339
R10236 DVDD.n693 DVDD.n692 0.0196339
R10237 DVDD.n692 DVDD.n687 0.0196339
R10238 DVDD.n746 DVDD.n687 0.0196339
R10239 DVDD.n747 DVDD.n686 0.0196339
R10240 DVDD.n751 DVDD.n686 0.0196339
R10241 DVDD.n752 DVDD.n751 0.0196339
R10242 DVDD.n753 DVDD.n752 0.0196339
R10243 DVDD.n753 DVDD.n684 0.0196339
R10244 DVDD.n757 DVDD.n684 0.0196339
R10245 DVDD.n758 DVDD.n757 0.0196339
R10246 DVDD.n759 DVDD.n758 0.0196339
R10247 DVDD.n759 DVDD.n682 0.0196339
R10248 DVDD.n763 DVDD.n682 0.0196339
R10249 DVDD.n764 DVDD.n763 0.0196339
R10250 DVDD.n765 DVDD.n764 0.0196339
R10251 DVDD.n765 DVDD.n680 0.0196339
R10252 DVDD.n769 DVDD.n680 0.0196339
R10253 DVDD.n770 DVDD.n769 0.0196339
R10254 DVDD.n771 DVDD.n770 0.0196339
R10255 DVDD.n771 DVDD.n678 0.0196339
R10256 DVDD.n775 DVDD.n678 0.0196339
R10257 DVDD.n776 DVDD.n775 0.0196339
R10258 DVDD.n777 DVDD.n776 0.0196339
R10259 DVDD.n777 DVDD.n676 0.0196339
R10260 DVDD.n781 DVDD.n676 0.0196339
R10261 DVDD.n782 DVDD.n781 0.0196339
R10262 DVDD.n783 DVDD.n782 0.0196339
R10263 DVDD.n783 DVDD.n674 0.0196339
R10264 DVDD.n787 DVDD.n674 0.0196339
R10265 DVDD.n788 DVDD.n787 0.0196339
R10266 DVDD.n8836 DVDD.n788 0.0196339
R10267 DVDD.n8835 DVDD.n789 0.0196339
R10268 DVDD.n8831 DVDD.n789 0.0196339
R10269 DVDD.n8831 DVDD.n8830 0.0196339
R10270 DVDD.n8830 DVDD.n8829 0.0196339
R10271 DVDD.n8829 DVDD.n8798 0.0196339
R10272 DVDD.n8825 DVDD.n8798 0.0196339
R10273 DVDD.n8825 DVDD.n8824 0.0196339
R10274 DVDD.n8824 DVDD.n8823 0.0196339
R10275 DVDD.n8818 DVDD.n8817 0.0196339
R10276 DVDD.n8802 DVDD.n8801 0.0196339
R10277 DVDD.n9645 DVDD.n74 0.0196339
R10278 DVDD.n9641 DVDD.n74 0.0196339
R10279 DVDD.n9641 DVDD.n9640 0.0196339
R10280 DVDD.n9640 DVDD.n9639 0.0196339
R10281 DVDD.n9639 DVDD.n77 0.0196339
R10282 DVDD.n9635 DVDD.n77 0.0196339
R10283 DVDD.n9635 DVDD.n9634 0.0196339
R10284 DVDD.n9633 DVDD.n79 0.0196339
R10285 DVDD.n843 DVDD.n82 0.0196339
R10286 DVDD.n940 DVDD.n855 0.0196339
R10287 DVDD.n935 DVDD.n934 0.0196339
R10288 DVDD.n934 DVDD.n873 0.0196339
R10289 DVDD.n8741 DVDD.n8740 0.0196339
R10290 DVDD.n997 DVDD.n904 0.0196339
R10291 DVDD.n3740 DVDD.n3636 0.0196339
R10292 DVDD.n3734 DVDD.n3733 0.0196339
R10293 DVDD.n3733 DVDD.n3732 0.0196339
R10294 DVDD.n3732 DVDD.n3641 0.0196339
R10295 DVDD.n3728 DVDD.n3641 0.0196339
R10296 DVDD.n3728 DVDD.n3727 0.0196339
R10297 DVDD.n3727 DVDD.n3726 0.0196339
R10298 DVDD.n3726 DVDD.n3643 0.0196339
R10299 DVDD.n3722 DVDD.n3643 0.0196339
R10300 DVDD.n3722 DVDD.n3721 0.0196339
R10301 DVDD.n3721 DVDD.n3720 0.0196339
R10302 DVDD.n3720 DVDD.n3645 0.0196339
R10303 DVDD.n3716 DVDD.n3645 0.0196339
R10304 DVDD.n3716 DVDD.n3715 0.0196339
R10305 DVDD.n3715 DVDD.n3714 0.0196339
R10306 DVDD.n3714 DVDD.n3647 0.0196339
R10307 DVDD.n3710 DVDD.n3647 0.0196339
R10308 DVDD.n3710 DVDD.n3709 0.0196339
R10309 DVDD.n3709 DVDD.n3708 0.0196339
R10310 DVDD.n3708 DVDD.n3649 0.0196339
R10311 DVDD.n3704 DVDD.n3649 0.0196339
R10312 DVDD.n3704 DVDD.n3703 0.0196339
R10313 DVDD.n3702 DVDD.n3701 0.0196339
R10314 DVDD.n3701 DVDD.n3650 0.0196339
R10315 DVDD.n3697 DVDD.n3650 0.0196339
R10316 DVDD.n3697 DVDD.n3696 0.0196339
R10317 DVDD.n3696 DVDD.n3695 0.0196339
R10318 DVDD.n3695 DVDD.n3652 0.0196339
R10319 DVDD.n3691 DVDD.n3652 0.0196339
R10320 DVDD.n3691 DVDD.n3690 0.0196339
R10321 DVDD.n3690 DVDD.n3689 0.0196339
R10322 DVDD.n3689 DVDD.n3654 0.0196339
R10323 DVDD.n3685 DVDD.n3654 0.0196339
R10324 DVDD.n3685 DVDD.n3684 0.0196339
R10325 DVDD.n3684 DVDD.n3683 0.0196339
R10326 DVDD.n3683 DVDD.n3656 0.0196339
R10327 DVDD.n3679 DVDD.n3656 0.0196339
R10328 DVDD.n3679 DVDD.n3678 0.0196339
R10329 DVDD.n3678 DVDD.n3677 0.0196339
R10330 DVDD.n3677 DVDD.n3658 0.0196339
R10331 DVDD.n3673 DVDD.n3658 0.0196339
R10332 DVDD.n3673 DVDD.n3672 0.0196339
R10333 DVDD.n3672 DVDD.n3671 0.0196339
R10334 DVDD.n3671 DVDD.n3660 0.0196339
R10335 DVDD.n3667 DVDD.n3660 0.0196339
R10336 DVDD.n3667 DVDD.n3666 0.0196339
R10337 DVDD.n3666 DVDD.n3665 0.0196339
R10338 DVDD.n3665 DVDD.n3662 0.0196339
R10339 DVDD.n3662 DVDD.n3574 0.0196339
R10340 DVDD.n3804 DVDD.n3574 0.0196339
R10341 DVDD.n3826 DVDD.n3825 0.0196339
R10342 DVDD.n3842 DVDD.n3841 0.0196339
R10343 DVDD.n3858 DVDD.n3857 0.0196339
R10344 DVDD.n6332 DVDD.n3819 0.0196339
R10345 DVDD.n6328 DVDD.n3819 0.0196339
R10346 DVDD.n6298 DVDD.n6245 0.0196339
R10347 DVDD.n6294 DVDD.n6245 0.0196339
R10348 DVDD.n6294 DVDD.n6293 0.0196339
R10349 DVDD.n6293 DVDD.n6292 0.0196339
R10350 DVDD.n6292 DVDD.n6247 0.0196339
R10351 DVDD.n6288 DVDD.n6247 0.0196339
R10352 DVDD.n6288 DVDD.n6287 0.0196339
R10353 DVDD.n6287 DVDD.n6286 0.0196339
R10354 DVDD.n6286 DVDD.n6249 0.0196339
R10355 DVDD.n6282 DVDD.n6249 0.0196339
R10356 DVDD.n6282 DVDD.n6281 0.0196339
R10357 DVDD.n6281 DVDD.n6280 0.0196339
R10358 DVDD.n6280 DVDD.n6251 0.0196339
R10359 DVDD.n6276 DVDD.n6251 0.0196339
R10360 DVDD.n6276 DVDD.n6275 0.0196339
R10361 DVDD.n6275 DVDD.n6274 0.0196339
R10362 DVDD.n6274 DVDD.n6253 0.0196339
R10363 DVDD.n6264 DVDD.n6263 0.0196339
R10364 DVDD.n6532 DVDD.n6531 0.0196339
R10365 DVDD.n6524 DVDD.n3358 0.0196339
R10366 DVDD.n6524 DVDD.n6523 0.0196339
R10367 DVDD.n6516 DVDD.n6515 0.0196339
R10368 DVDD.n6500 DVDD.n6499 0.0196339
R10369 DVDD.n8979 DVDD.n8978 0.0196339
R10370 DVDD.n9008 DVDD.n9007 0.0196339
R10371 DVDD.n9002 DVDD.n9001 0.0196339
R10372 DVDD.n9001 DVDD.n9000 0.0196339
R10373 DVDD.n9000 DVDD.n8991 0.0196339
R10374 DVDD.n8996 DVDD.n8991 0.0196339
R10375 DVDD.n8996 DVDD.n8995 0.0196339
R10376 DVDD.n8995 DVDD.n8994 0.0196339
R10377 DVDD.n8994 DVDD.n545 0.0196339
R10378 DVDD.n9018 DVDD.n545 0.0196339
R10379 DVDD.n9070 DVDD.n9069 0.0196339
R10380 DVDD.n9069 DVDD.n9068 0.0196339
R10381 DVDD.n9068 DVDD.n9019 0.0196339
R10382 DVDD.n9064 DVDD.n9019 0.0196339
R10383 DVDD.n9064 DVDD.n9063 0.0196339
R10384 DVDD.n9063 DVDD.n9062 0.0196339
R10385 DVDD.n9062 DVDD.n9021 0.0196339
R10386 DVDD.n9058 DVDD.n9021 0.0196339
R10387 DVDD.n9058 DVDD.n9057 0.0196339
R10388 DVDD.n9057 DVDD.n9056 0.0196339
R10389 DVDD.n9056 DVDD.n9023 0.0196339
R10390 DVDD.n9052 DVDD.n9023 0.0196339
R10391 DVDD.n9052 DVDD.n9051 0.0196339
R10392 DVDD.n9051 DVDD.n9050 0.0196339
R10393 DVDD.n9050 DVDD.n9025 0.0196339
R10394 DVDD.n9046 DVDD.n9025 0.0196339
R10395 DVDD.n9046 DVDD.n9045 0.0196339
R10396 DVDD.n9045 DVDD.n9044 0.0196339
R10397 DVDD.n9044 DVDD.n9027 0.0196339
R10398 DVDD.n9040 DVDD.n9027 0.0196339
R10399 DVDD.n9040 DVDD.n9039 0.0196339
R10400 DVDD.n9039 DVDD.n9038 0.0196339
R10401 DVDD.n9038 DVDD.n9029 0.0196339
R10402 DVDD.n9034 DVDD.n9029 0.0196339
R10403 DVDD.n9034 DVDD.n9033 0.0196339
R10404 DVDD.n9033 DVDD.n9032 0.0196339
R10405 DVDD.n9032 DVDD.n542 0.0196339
R10406 DVDD.n9074 DVDD.n542 0.0196339
R10407 DVDD.n9106 DVDD.n9105 0.0196339
R10408 DVDD.n9105 DVDD.n9104 0.0196339
R10409 DVDD.n9104 DVDD.n9075 0.0196339
R10410 DVDD.n9100 DVDD.n9075 0.0196339
R10411 DVDD.n9100 DVDD.n9099 0.0196339
R10412 DVDD.n9099 DVDD.n9098 0.0196339
R10413 DVDD.n9098 DVDD.n9077 0.0196339
R10414 DVDD.n9094 DVDD.n9077 0.0196339
R10415 DVDD.n9090 DVDD.n9089 0.0196339
R10416 DVDD.n9125 DVDD.n535 0.0196339
R10417 DVDD.n9119 DVDD.n9118 0.0196339
R10418 DVDD.n9118 DVDD.n9117 0.0196339
R10419 DVDD.n9117 DVDD.n538 0.0196339
R10420 DVDD.n9113 DVDD.n538 0.0196339
R10421 DVDD.n9113 DVDD.n9112 0.0196339
R10422 DVDD.n9112 DVDD.n9111 0.0196339
R10423 DVDD.n9111 DVDD.n540 0.0196339
R10424 DVDD.n4114 DVDD.n4113 0.0196339
R10425 DVDD.n4008 DVDD.n4007 0.0196339
R10426 DVDD.n4040 DVDD.n4037 0.0196339
R10427 DVDD.n4052 DVDD.n4051 0.0196339
R10428 DVDD.n4053 DVDD.n4052 0.0196339
R10429 DVDD.n4065 DVDD.n4063 0.0196339
R10430 DVDD.n4118 DVDD.n3984 0.0196339
R10431 DVDD.n4161 DVDD.n4159 0.0196339
R10432 DVDD.n4202 DVDD.n4201 0.0196339
R10433 DVDD.n4201 DVDD.n4200 0.0196339
R10434 DVDD.n4200 DVDD.n4165 0.0196339
R10435 DVDD.n4196 DVDD.n4165 0.0196339
R10436 DVDD.n4196 DVDD.n4195 0.0196339
R10437 DVDD.n4195 DVDD.n4194 0.0196339
R10438 DVDD.n4194 DVDD.n4167 0.0196339
R10439 DVDD.n4190 DVDD.n4167 0.0196339
R10440 DVDD.n4190 DVDD.n4189 0.0196339
R10441 DVDD.n4189 DVDD.n4188 0.0196339
R10442 DVDD.n4188 DVDD.n4169 0.0196339
R10443 DVDD.n4184 DVDD.n4169 0.0196339
R10444 DVDD.n4184 DVDD.n4183 0.0196339
R10445 DVDD.n4183 DVDD.n4182 0.0196339
R10446 DVDD.n4182 DVDD.n4171 0.0196339
R10447 DVDD.n4178 DVDD.n4171 0.0196339
R10448 DVDD.n4178 DVDD.n4177 0.0196339
R10449 DVDD.n4177 DVDD.n4176 0.0196339
R10450 DVDD.n4176 DVDD.n4173 0.0196339
R10451 DVDD.n4173 DVDD.n3973 0.0196339
R10452 DVDD.n4223 DVDD.n3973 0.0196339
R10453 DVDD.n4275 DVDD.n4274 0.0196339
R10454 DVDD.n4274 DVDD.n4273 0.0196339
R10455 DVDD.n4273 DVDD.n4224 0.0196339
R10456 DVDD.n4269 DVDD.n4224 0.0196339
R10457 DVDD.n4269 DVDD.n4268 0.0196339
R10458 DVDD.n4268 DVDD.n4267 0.0196339
R10459 DVDD.n4267 DVDD.n4226 0.0196339
R10460 DVDD.n4263 DVDD.n4226 0.0196339
R10461 DVDD.n4263 DVDD.n4262 0.0196339
R10462 DVDD.n4262 DVDD.n4261 0.0196339
R10463 DVDD.n4261 DVDD.n4228 0.0196339
R10464 DVDD.n4257 DVDD.n4228 0.0196339
R10465 DVDD.n4257 DVDD.n4256 0.0196339
R10466 DVDD.n4256 DVDD.n4255 0.0196339
R10467 DVDD.n4255 DVDD.n4230 0.0196339
R10468 DVDD.n4251 DVDD.n4230 0.0196339
R10469 DVDD.n4251 DVDD.n4250 0.0196339
R10470 DVDD.n4250 DVDD.n4249 0.0196339
R10471 DVDD.n4249 DVDD.n4232 0.0196339
R10472 DVDD.n4245 DVDD.n4232 0.0196339
R10473 DVDD.n4245 DVDD.n4244 0.0196339
R10474 DVDD.n4244 DVDD.n4243 0.0196339
R10475 DVDD.n4243 DVDD.n4234 0.0196339
R10476 DVDD.n4239 DVDD.n4234 0.0196339
R10477 DVDD.n4239 DVDD.n4238 0.0196339
R10478 DVDD.n4238 DVDD.n4237 0.0196339
R10479 DVDD.n4237 DVDD.n3970 0.0196339
R10480 DVDD.n4279 DVDD.n3970 0.0196339
R10481 DVDD.n6044 DVDD.n6043 0.0196339
R10482 DVDD.n6028 DVDD.n6027 0.0196339
R10483 DVDD.n6012 DVDD.n6011 0.0196339
R10484 DVDD.n6006 DVDD.n6005 0.0196339
R10485 DVDD.n6005 DVDD.n5931 0.0196339
R10486 DVDD.n5989 DVDD.n5988 0.0196339
R10487 DVDD.n5988 DVDD.n5987 0.0196339
R10488 DVDD.n5987 DVDD.n5935 0.0196339
R10489 DVDD.n5983 DVDD.n5935 0.0196339
R10490 DVDD.n5983 DVDD.n5982 0.0196339
R10491 DVDD.n5982 DVDD.n5981 0.0196339
R10492 DVDD.n5981 DVDD.n5937 0.0196339
R10493 DVDD.n5977 DVDD.n5937 0.0196339
R10494 DVDD.n5977 DVDD.n5976 0.0196339
R10495 DVDD.n5976 DVDD.n5975 0.0196339
R10496 DVDD.n5975 DVDD.n5939 0.0196339
R10497 DVDD.n5971 DVDD.n5939 0.0196339
R10498 DVDD.n5971 DVDD.n5970 0.0196339
R10499 DVDD.n5970 DVDD.n5969 0.0196339
R10500 DVDD.n5969 DVDD.n5941 0.0196339
R10501 DVDD.n5965 DVDD.n5941 0.0196339
R10502 DVDD.n5965 DVDD.n5964 0.0196339
R10503 DVDD.n5955 DVDD.n5954 0.0196339
R10504 DVDD.n3296 DVDD.n3239 0.0196339
R10505 DVDD.n3288 DVDD.n3287 0.0196339
R10506 DVDD.n3287 DVDD.n3286 0.0196339
R10507 DVDD.n3279 DVDD.n3278 0.0196339
R10508 DVDD.n3263 DVDD.n3262 0.0196339
R10509 DVDD.n4875 DVDD.n4868 0.0196339
R10510 DVDD.n5014 DVDD.n5013 0.0196339
R10511 DVDD.n5008 DVDD.n5007 0.0196339
R10512 DVDD.n5007 DVDD.n5006 0.0196339
R10513 DVDD.n5006 DVDD.n4872 0.0196339
R10514 DVDD.n5002 DVDD.n4872 0.0196339
R10515 DVDD.n5002 DVDD.n5001 0.0196339
R10516 DVDD.n5001 DVDD.n5000 0.0196339
R10517 DVDD.n5000 DVDD.n4874 0.0196339
R10518 DVDD.n4996 DVDD.n4874 0.0196339
R10519 DVDD.n4995 DVDD.n4881 0.0196339
R10520 DVDD.n4991 DVDD.n4881 0.0196339
R10521 DVDD.n4991 DVDD.n4990 0.0196339
R10522 DVDD.n4990 DVDD.n4989 0.0196339
R10523 DVDD.n4989 DVDD.n4883 0.0196339
R10524 DVDD.n4985 DVDD.n4883 0.0196339
R10525 DVDD.n4985 DVDD.n4984 0.0196339
R10526 DVDD.n4984 DVDD.n4983 0.0196339
R10527 DVDD.n4983 DVDD.n4885 0.0196339
R10528 DVDD.n4979 DVDD.n4885 0.0196339
R10529 DVDD.n4979 DVDD.n4978 0.0196339
R10530 DVDD.n4978 DVDD.n4977 0.0196339
R10531 DVDD.n4977 DVDD.n4887 0.0196339
R10532 DVDD.n4973 DVDD.n4887 0.0196339
R10533 DVDD.n4973 DVDD.n4972 0.0196339
R10534 DVDD.n4972 DVDD.n4971 0.0196339
R10535 DVDD.n4971 DVDD.n4889 0.0196339
R10536 DVDD.n4967 DVDD.n4889 0.0196339
R10537 DVDD.n4967 DVDD.n4966 0.0196339
R10538 DVDD.n4966 DVDD.n4965 0.0196339
R10539 DVDD.n4965 DVDD.n4891 0.0196339
R10540 DVDD.n4961 DVDD.n4891 0.0196339
R10541 DVDD.n4961 DVDD.n4960 0.0196339
R10542 DVDD.n4960 DVDD.n4959 0.0196339
R10543 DVDD.n4959 DVDD.n4893 0.0196339
R10544 DVDD.n4955 DVDD.n4893 0.0196339
R10545 DVDD.n4955 DVDD.n4954 0.0196339
R10546 DVDD.n4954 DVDD.n4953 0.0196339
R10547 DVDD.n4950 DVDD.n4895 0.0196339
R10548 DVDD.n4946 DVDD.n4895 0.0196339
R10549 DVDD.n4946 DVDD.n4945 0.0196339
R10550 DVDD.n4945 DVDD.n4944 0.0196339
R10551 DVDD.n4944 DVDD.n4897 0.0196339
R10552 DVDD.n4940 DVDD.n4897 0.0196339
R10553 DVDD.n4940 DVDD.n4939 0.0196339
R10554 DVDD.n4939 DVDD.n4938 0.0196339
R10555 DVDD.n4933 DVDD.n4932 0.0196339
R10556 DVDD.n4917 DVDD.n4916 0.0196339
R10557 DVDD.n4911 DVDD.n497 0.0196339
R10558 DVDD.n4911 DVDD.n4910 0.0196339
R10559 DVDD.n4910 DVDD.n4909 0.0196339
R10560 DVDD.n4909 DVDD.n4900 0.0196339
R10561 DVDD.n4905 DVDD.n4900 0.0196339
R10562 DVDD.n4905 DVDD.n4904 0.0196339
R10563 DVDD.n4904 DVDD.n287 0.0196339
R10564 DVDD.n9474 DVDD.n9473 0.0196339
R10565 DVDD.n303 DVDD.n301 0.0196339
R10566 DVDD.n317 DVDD.n314 0.0196339
R10567 DVDD.n335 DVDD.n321 0.0196339
R10568 DVDD.n336 DVDD.n335 0.0196339
R10569 DVDD.n9437 DVDD.n332 0.0196339
R10570 DVDD.n9478 DVDD.n275 0.0196339
R10571 DVDD.n9554 DVDD.n246 0.0196339
R10572 DVDD.n9545 DVDD.n255 0.0196339
R10573 DVDD.n9541 DVDD.n255 0.0196339
R10574 DVDD.n9541 DVDD.n9540 0.0196339
R10575 DVDD.n9540 DVDD.n9539 0.0196339
R10576 DVDD.n9539 DVDD.n257 0.0196339
R10577 DVDD.n9535 DVDD.n257 0.0196339
R10578 DVDD.n9535 DVDD.n9534 0.0196339
R10579 DVDD.n9534 DVDD.n9533 0.0196339
R10580 DVDD.n9533 DVDD.n259 0.0196339
R10581 DVDD.n9529 DVDD.n259 0.0196339
R10582 DVDD.n9529 DVDD.n9528 0.0196339
R10583 DVDD.n9528 DVDD.n9527 0.0196339
R10584 DVDD.n9527 DVDD.n261 0.0196339
R10585 DVDD.n9523 DVDD.n261 0.0196339
R10586 DVDD.n9523 DVDD.n9522 0.0196339
R10587 DVDD.n9522 DVDD.n9521 0.0196339
R10588 DVDD.n9521 DVDD.n263 0.0196339
R10589 DVDD.n9517 DVDD.n263 0.0196339
R10590 DVDD.n9517 DVDD.n9516 0.0196339
R10591 DVDD.n9516 DVDD.n9515 0.0196339
R10592 DVDD.n9515 DVDD.n265 0.0196339
R10593 DVDD.n4371 DVDD.n4370 0.0196339
R10594 DVDD.n4370 DVDD.n4369 0.0196339
R10595 DVDD.n4369 DVDD.n4320 0.0196339
R10596 DVDD.n4365 DVDD.n4320 0.0196339
R10597 DVDD.n4365 DVDD.n4364 0.0196339
R10598 DVDD.n4364 DVDD.n4363 0.0196339
R10599 DVDD.n4363 DVDD.n4322 0.0196339
R10600 DVDD.n4359 DVDD.n4322 0.0196339
R10601 DVDD.n4359 DVDD.n4358 0.0196339
R10602 DVDD.n4358 DVDD.n4357 0.0196339
R10603 DVDD.n4357 DVDD.n4324 0.0196339
R10604 DVDD.n4353 DVDD.n4324 0.0196339
R10605 DVDD.n4353 DVDD.n4352 0.0196339
R10606 DVDD.n4352 DVDD.n4351 0.0196339
R10607 DVDD.n4351 DVDD.n4326 0.0196339
R10608 DVDD.n4347 DVDD.n4326 0.0196339
R10609 DVDD.n4347 DVDD.n4346 0.0196339
R10610 DVDD.n4346 DVDD.n4345 0.0196339
R10611 DVDD.n4345 DVDD.n4328 0.0196339
R10612 DVDD.n4341 DVDD.n4328 0.0196339
R10613 DVDD.n4341 DVDD.n4340 0.0196339
R10614 DVDD.n4340 DVDD.n4339 0.0196339
R10615 DVDD.n4339 DVDD.n4330 0.0196339
R10616 DVDD.n4335 DVDD.n4330 0.0196339
R10617 DVDD.n4335 DVDD.n4334 0.0196339
R10618 DVDD.n4334 DVDD.n4333 0.0196339
R10619 DVDD.n4333 DVDD.n4317 0.0196339
R10620 DVDD.n4375 DVDD.n4317 0.0196339
R10621 DVDD.n5811 DVDD.n5810 0.0196339
R10622 DVDD.n5795 DVDD.n5794 0.0196339
R10623 DVDD.n5779 DVDD.n5778 0.0196339
R10624 DVDD.n5773 DVDD.n4389 0.0196339
R10625 DVDD.n5773 DVDD.n5772 0.0196339
R10626 DVDD.n5887 DVDD.n5830 0.0196339
R10627 DVDD.n5883 DVDD.n5830 0.0196339
R10628 DVDD.n5883 DVDD.n5882 0.0196339
R10629 DVDD.n5882 DVDD.n5881 0.0196339
R10630 DVDD.n5881 DVDD.n5833 0.0196339
R10631 DVDD.n5877 DVDD.n5833 0.0196339
R10632 DVDD.n5877 DVDD.n5876 0.0196339
R10633 DVDD.n5876 DVDD.n5875 0.0196339
R10634 DVDD.n5875 DVDD.n5835 0.0196339
R10635 DVDD.n5871 DVDD.n5835 0.0196339
R10636 DVDD.n5871 DVDD.n5870 0.0196339
R10637 DVDD.n5870 DVDD.n5869 0.0196339
R10638 DVDD.n5869 DVDD.n5837 0.0196339
R10639 DVDD.n5865 DVDD.n5837 0.0196339
R10640 DVDD.n5865 DVDD.n5864 0.0196339
R10641 DVDD.n5864 DVDD.n5863 0.0196339
R10642 DVDD.n5863 DVDD.n5839 0.0196339
R10643 DVDD.n5853 DVDD.n5852 0.0196339
R10644 DVDD.n3129 DVDD.n3128 0.0196339
R10645 DVDD.n3180 DVDD.n3123 0.0196339
R10646 DVDD.n3176 DVDD.n3123 0.0196339
R10647 DVDD.n3170 DVDD.n3169 0.0196339
R10648 DVDD.n3154 DVDD.n3153 0.0196339
R10649 DVDD.n5123 DVDD.n5122 0.0196339
R10650 DVDD.n5152 DVDD.n5151 0.0196339
R10651 DVDD.n5146 DVDD.n5145 0.0196339
R10652 DVDD.n5145 DVDD.n5144 0.0196339
R10653 DVDD.n5144 DVDD.n5135 0.0196339
R10654 DVDD.n5140 DVDD.n5135 0.0196339
R10655 DVDD.n5140 DVDD.n5139 0.0196339
R10656 DVDD.n5139 DVDD.n5138 0.0196339
R10657 DVDD.n5138 DVDD.n4565 0.0196339
R10658 DVDD.n5161 DVDD.n4565 0.0196339
R10659 DVDD.n5215 DVDD.n5214 0.0196339
R10660 DVDD.n5214 DVDD.n5213 0.0196339
R10661 DVDD.n5213 DVDD.n5162 0.0196339
R10662 DVDD.n5209 DVDD.n5162 0.0196339
R10663 DVDD.n5209 DVDD.n5208 0.0196339
R10664 DVDD.n5208 DVDD.n5207 0.0196339
R10665 DVDD.n5207 DVDD.n5164 0.0196339
R10666 DVDD.n5203 DVDD.n5164 0.0196339
R10667 DVDD.n5203 DVDD.n5202 0.0196339
R10668 DVDD.n5202 DVDD.n5201 0.0196339
R10669 DVDD.n5201 DVDD.n5166 0.0196339
R10670 DVDD.n5197 DVDD.n5166 0.0196339
R10671 DVDD.n5197 DVDD.n5196 0.0196339
R10672 DVDD.n5196 DVDD.n5195 0.0196339
R10673 DVDD.n5195 DVDD.n5168 0.0196339
R10674 DVDD.n5191 DVDD.n5168 0.0196339
R10675 DVDD.n5191 DVDD.n5190 0.0196339
R10676 DVDD.n5190 DVDD.n5189 0.0196339
R10677 DVDD.n5189 DVDD.n5170 0.0196339
R10678 DVDD.n5185 DVDD.n5170 0.0196339
R10679 DVDD.n5185 DVDD.n5184 0.0196339
R10680 DVDD.n5184 DVDD.n5183 0.0196339
R10681 DVDD.n5183 DVDD.n5172 0.0196339
R10682 DVDD.n5179 DVDD.n5172 0.0196339
R10683 DVDD.n5179 DVDD.n5178 0.0196339
R10684 DVDD.n5178 DVDD.n5177 0.0196339
R10685 DVDD.n5177 DVDD.n5174 0.0196339
R10686 DVDD.n5174 DVDD.n451 0.0196339
R10687 DVDD.n9298 DVDD.n9297 0.0196339
R10688 DVDD.n9297 DVDD.n9296 0.0196339
R10689 DVDD.n9296 DVDD.n452 0.0196339
R10690 DVDD.n9292 DVDD.n452 0.0196339
R10691 DVDD.n9292 DVDD.n9291 0.0196339
R10692 DVDD.n9291 DVDD.n9290 0.0196339
R10693 DVDD.n9290 DVDD.n454 0.0196339
R10694 DVDD.n9286 DVDD.n454 0.0196339
R10695 DVDD.n9253 DVDD.n9252 0.0196339
R10696 DVDD.n9282 DVDD.n9250 0.0196339
R10697 DVDD.n9276 DVDD.n9275 0.0196339
R10698 DVDD.n9275 DVDD.n9274 0.0196339
R10699 DVDD.n9274 DVDD.n9267 0.0196339
R10700 DVDD.n9270 DVDD.n9267 0.0196339
R10701 DVDD.n9270 DVDD.n9269 0.0196339
R10702 DVDD.n9269 DVDD.n446 0.0196339
R10703 DVDD.n9301 DVDD.n446 0.0196339
R10704 DVDD.n9303 DVDD.n9302 0.0196339
R10705 DVDD.n443 DVDD.n437 0.0196339
R10706 DVDD.n9608 DVDD.n9607 0.0196339
R10707 DVDD.n160 DVDD.n143 0.0196339
R10708 DVDD.n160 DVDD.n154 0.0196339
R10709 DVDD.n172 DVDD.n165 0.0196339
R10710 DVDD.n9410 DVDD.n9409 0.0196339
R10711 DVDD.n6786 DVDD.n2901 0.0196339
R10712 DVDD.n2956 DVDD.n2917 0.0196339
R10713 DVDD.n2952 DVDD.n2917 0.0196339
R10714 DVDD.n2952 DVDD.n2951 0.0196339
R10715 DVDD.n2951 DVDD.n2950 0.0196339
R10716 DVDD.n2950 DVDD.n2919 0.0196339
R10717 DVDD.n2946 DVDD.n2919 0.0196339
R10718 DVDD.n2946 DVDD.n2945 0.0196339
R10719 DVDD.n2945 DVDD.n2944 0.0196339
R10720 DVDD.n2944 DVDD.n2921 0.0196339
R10721 DVDD.n2940 DVDD.n2921 0.0196339
R10722 DVDD.n2940 DVDD.n2939 0.0196339
R10723 DVDD.n2939 DVDD.n2938 0.0196339
R10724 DVDD.n2938 DVDD.n2923 0.0196339
R10725 DVDD.n2934 DVDD.n2923 0.0196339
R10726 DVDD.n2934 DVDD.n2933 0.0196339
R10727 DVDD.n2933 DVDD.n2932 0.0196339
R10728 DVDD.n2932 DVDD.n2925 0.0196339
R10729 DVDD.n2928 DVDD.n2925 0.0196339
R10730 DVDD.n2928 DVDD.n2927 0.0196339
R10731 DVDD.n2927 DVDD.n2884 0.0196339
R10732 DVDD.n6798 DVDD.n2884 0.0196339
R10733 DVDD.n6850 DVDD.n6849 0.0196339
R10734 DVDD.n6849 DVDD.n6848 0.0196339
R10735 DVDD.n6848 DVDD.n6799 0.0196339
R10736 DVDD.n6844 DVDD.n6799 0.0196339
R10737 DVDD.n6844 DVDD.n6843 0.0196339
R10738 DVDD.n6843 DVDD.n6842 0.0196339
R10739 DVDD.n6842 DVDD.n6801 0.0196339
R10740 DVDD.n6838 DVDD.n6801 0.0196339
R10741 DVDD.n6838 DVDD.n6837 0.0196339
R10742 DVDD.n6837 DVDD.n6836 0.0196339
R10743 DVDD.n6836 DVDD.n6803 0.0196339
R10744 DVDD.n6832 DVDD.n6803 0.0196339
R10745 DVDD.n6832 DVDD.n6831 0.0196339
R10746 DVDD.n6831 DVDD.n6830 0.0196339
R10747 DVDD.n6830 DVDD.n6805 0.0196339
R10748 DVDD.n6826 DVDD.n6805 0.0196339
R10749 DVDD.n6826 DVDD.n6825 0.0196339
R10750 DVDD.n6825 DVDD.n6824 0.0196339
R10751 DVDD.n6824 DVDD.n6807 0.0196339
R10752 DVDD.n6820 DVDD.n6807 0.0196339
R10753 DVDD.n6820 DVDD.n6819 0.0196339
R10754 DVDD.n6819 DVDD.n6818 0.0196339
R10755 DVDD.n6818 DVDD.n6809 0.0196339
R10756 DVDD.n6814 DVDD.n6809 0.0196339
R10757 DVDD.n6814 DVDD.n6813 0.0196339
R10758 DVDD.n6813 DVDD.n6812 0.0196339
R10759 DVDD.n6812 DVDD.n2879 0.0196339
R10760 DVDD.n6853 DVDD.n2879 0.0196339
R10761 DVDD.n2871 DVDD.n2870 0.0196339
R10762 DVDD.n2855 DVDD.n2854 0.0196339
R10763 DVDD.n2839 DVDD.n2838 0.0196339
R10764 DVDD.n2833 DVDD.n2832 0.0196339
R10765 DVDD.n2832 DVDD.n2797 0.0196339
R10766 DVDD.n2776 DVDD.n2775 0.0196339
R10767 DVDD.n2775 DVDD.n2744 0.0196339
R10768 DVDD.n2771 DVDD.n2744 0.0196339
R10769 DVDD.n2771 DVDD.n2770 0.0196339
R10770 DVDD.n2770 DVDD.n2769 0.0196339
R10771 DVDD.n2769 DVDD.n2746 0.0196339
R10772 DVDD.n2765 DVDD.n2746 0.0196339
R10773 DVDD.n2765 DVDD.n2764 0.0196339
R10774 DVDD.n2764 DVDD.n2763 0.0196339
R10775 DVDD.n2763 DVDD.n2748 0.0196339
R10776 DVDD.n2759 DVDD.n2748 0.0196339
R10777 DVDD.n2759 DVDD.n2758 0.0196339
R10778 DVDD.n2758 DVDD.n2757 0.0196339
R10779 DVDD.n2757 DVDD.n2750 0.0196339
R10780 DVDD.n2753 DVDD.n2750 0.0196339
R10781 DVDD.n2753 DVDD.n2752 0.0196339
R10782 DVDD.n2752 DVDD.n2737 0.0196339
R10783 DVDD.n6915 DVDD.n6914 0.0196339
R10784 DVDD.n2717 DVDD.n2716 0.0196339
R10785 DVDD.n2709 DVDD.n2708 0.0196339
R10786 DVDD.n2708 DVDD.n2707 0.0196339
R10787 DVDD.n2700 DVDD.n2699 0.0196339
R10788 DVDD.n2684 DVDD.n2683 0.0196339
R10789 DVDD.n8452 DVDD.n8451 0.0196339
R10790 DVDD.n8453 DVDD.n8452 0.0196339
R10791 DVDD.n8453 DVDD.n8445 0.0196339
R10792 DVDD.n8457 DVDD.n8445 0.0196339
R10793 DVDD.n8458 DVDD.n8457 0.0196339
R10794 DVDD.n8459 DVDD.n8458 0.0196339
R10795 DVDD.n8459 DVDD.n8444 0.0196339
R10796 DVDD.n8463 DVDD.n8444 0.0196339
R10797 DVDD.n8464 DVDD.n8463 0.0196339
R10798 DVDD.n8466 DVDD.n8464 0.0196339
R10799 DVDD.n8470 DVDD.n1444 0.0196339
R10800 DVDD.n8471 DVDD.n8470 0.0196339
R10801 DVDD.n8472 DVDD.n8471 0.0196339
R10802 DVDD.n8472 DVDD.n1442 0.0196339
R10803 DVDD.n8476 DVDD.n1442 0.0196339
R10804 DVDD.n8477 DVDD.n8476 0.0196339
R10805 DVDD.n8478 DVDD.n8477 0.0196339
R10806 DVDD.n8478 DVDD.n1440 0.0196339
R10807 DVDD.n8482 DVDD.n1440 0.0196339
R10808 DVDD.n8491 DVDD.n8482 0.0196339
R10809 DVDD.n8489 DVDD.n8488 0.0196339
R10810 DVDD.n8488 DVDD.n8483 0.0196339
R10811 DVDD.n8484 DVDD.n8483 0.0196339
R10812 DVDD.n8484 DVDD.n1346 0.0196339
R10813 DVDD.n8613 DVDD.n1346 0.0196339
R10814 DVDD.n8613 DVDD.n8612 0.0196339
R10815 DVDD.n8612 DVDD.n8611 0.0196339
R10816 DVDD.n8611 DVDD.n1347 0.0196339
R10817 DVDD.n8607 DVDD.n1347 0.0196339
R10818 DVDD.n8607 DVDD.n8606 0.0196339
R10819 DVDD.n8604 DVDD.n1351 0.0196339
R10820 DVDD.n8526 DVDD.n1351 0.0196339
R10821 DVDD.n8526 DVDD.n8524 0.0196339
R10822 DVDD.n8530 DVDD.n8524 0.0196339
R10823 DVDD.n8391 DVDD.n1495 0.0196339
R10824 DVDD.n8392 DVDD.n8391 0.0196339
R10825 DVDD.n8393 DVDD.n8392 0.0196339
R10826 DVDD.n8393 DVDD.n1493 0.0196339
R10827 DVDD.n8397 DVDD.n1493 0.0196339
R10828 DVDD.n8398 DVDD.n8397 0.0196339
R10829 DVDD.n8399 DVDD.n8398 0.0196339
R10830 DVDD.n8399 DVDD.n1491 0.0196339
R10831 DVDD.n8403 DVDD.n1491 0.0196339
R10832 DVDD.n8404 DVDD.n8403 0.0196339
R10833 DVDD.n8414 DVDD.n8413 0.0196339
R10834 DVDD.n8413 DVDD.n8408 0.0196339
R10835 DVDD.n8409 DVDD.n8408 0.0196339
R10836 DVDD.n8409 DVDD.n1379 0.0196339
R10837 DVDD.n8584 DVDD.n1379 0.0196339
R10838 DVDD.n8584 DVDD.n8583 0.0196339
R10839 DVDD.n8583 DVDD.n8582 0.0196339
R10840 DVDD.n8582 DVDD.n1380 0.0196339
R10841 DVDD.n8578 DVDD.n1380 0.0196339
R10842 DVDD.n8578 DVDD.n8577 0.0196339
R10843 DVDD.n8573 DVDD.n8572 0.0196339
R10844 DVDD.n8572 DVDD.n1384 0.0196339
R10845 DVDD.n8568 DVDD.n1384 0.0196339
R10846 DVDD.n8568 DVDD.n8567 0.0196339
R10847 DVDD.n8567 DVDD.n8566 0.0196339
R10848 DVDD.n8566 DVDD.n1386 0.0196339
R10849 DVDD.n8562 DVDD.n1386 0.0196339
R10850 DVDD.n8562 DVDD.n8561 0.0196339
R10851 DVDD.n8561 DVDD.n8560 0.0196339
R10852 DVDD.n8560 DVDD.n1388 0.0196339
R10853 DVDD.n8556 DVDD.n8555 0.0196339
R10854 DVDD.n8555 DVDD.n8554 0.0196339
R10855 DVDD.n8554 DVDD.n1395 0.0196339
R10856 DVDD.n8550 DVDD.n1395 0.0196339
R10857 DVDD.n8680 DVDD.n8679 0.019625
R10858 DVDD.n8733 DVDD.n8732 0.019625
R10859 DVDD.n6316 DVDD.n6315 0.019625
R10860 DVDD.n6878 DVDD.n2791 0.019625
R10861 DVDD.n9583 DVDD.n175 0.019625
R10862 DVDD.n2910 DVDD.n2891 0.019625
R10863 DVDD.n9350 DVDD.n132 0.019625
R10864 DVDD.n856 DVDD.n849 0.019625
R10865 DVDD.n8430 DVDD.n8429 0.0195909
R10866 DVDD.n8503 DVDD.n8502 0.0195909
R10867 DVDD.n8591 DVDD.n8590 0.0195909
R10868 DVDD.n8429 DVDD.t0 0.0195909
R10869 DVDD.n8502 DVDD.t0 0.0195909
R10870 DVDD.n8590 DVDD.t0 0.0195909
R10871 DVDD.n707 DVDD.n581 0.0194567
R10872 DVDD.n9629 DVDD.n9628 0.0194567
R10873 DVDD.n996 DVDD.n916 0.0194567
R10874 DVDD.n3828 DVDD.n3569 0.0194567
R10875 DVDD.n9011 DVDD.n8973 0.0194567
R10876 DVDD.n4004 DVDD.n3997 0.0194567
R10877 DVDD.n4121 DVDD.n3994 0.0194567
R10878 DVDD.n6040 DVDD.n3966 0.0194567
R10879 DVDD.n5016 DVDD.n4859 0.0194567
R10880 DVDD.n300 DVDD.n288 0.0194567
R10881 DVDD.n9481 DVDD.n284 0.0194567
R10882 DVDD.n5807 DVDD.n4313 0.0194567
R10883 DVDD.n5155 DVDD.n5117 0.0194567
R10884 DVDD.n9315 DVDD.n436 0.0194567
R10885 DVDD.n9413 DVDD.n389 0.0194567
R10886 DVDD.n2867 DVDD.n2828 0.0194567
R10887 DVDD.n941 DVDD.n864 0.0191024
R10888 DVDD.n6266 DVDD.n3346 0.0191024
R10889 DVDD.n4044 DVDD.n4043 0.0191024
R10890 DVDD.n5957 DVDD.n3217 0.0191024
R10891 DVDD.n9451 DVDD.n9450 0.0191024
R10892 DVDD.n5855 DVDD.n3111 0.0191024
R10893 DVDD.n9606 DVDD.n136 0.0191024
R10894 DVDD.n6917 DVDD.n2662 0.0191024
R10895 DVDD.n723 DVDD.n586 0.018748
R10896 DVDD.n8804 DVDD.n70 0.018748
R10897 DVDD.n8744 DVDD.n877 0.018748
R10898 DVDD.n3741 DVDD.n1042 0.018748
R10899 DVDD.n3844 DVDD.n3814 0.018748
R10900 DVDD.n3874 DVDD.n3867 0.018748
R10901 DVDD.n6512 DVDD.n2084 0.018748
R10902 DVDD.n554 DVDD.n550 0.018748
R10903 DVDD.n9174 DVDD.n532 0.018748
R10904 DVDD.n4062 DVDD.n4030 0.018748
R10905 DVDD.n4158 DVDD.n4147 0.018748
R10906 DVDD.n6024 DVDD.n3954 0.018748
R10907 DVDD.n6055 DVDD.n5924 0.018748
R10908 DVDD.n3275 DVDD.n2142 0.018748
R10909 DVDD.n4877 DVDD.n4857 0.018748
R10910 DVDD.n4919 DVDD.n494 0.018748
R10911 DVDD.n9438 DVDD.n331 0.018748
R10912 DVDD.n9555 DVDD.n245 0.018748
R10913 DVDD.n5791 DVDD.n4383 0.018748
R10914 DVDD.n5823 DVDD.n5763 0.018748
R10915 DVDD.n3166 DVDD.n2181 0.018748
R10916 DVDD.n4576 DVDD.n4572 0.018748
R10917 DVDD.n9283 DVDD.n9249 0.018748
R10918 DVDD.n9591 DVDD.n9590 0.018748
R10919 DVDD.n6787 DVDD.n2892 0.018748
R10920 DVDD.n2851 DVDD.n2815 0.018748
R10921 DVDD.n6873 DVDD.n2792 0.018748
R10922 DVDD.n2696 DVDD.n2634 0.018748
R10923 DVDD.n9379 DVDD.n153 0.0183937
R10924 DVDD.n9383 DVDD.n9382 0.0183937
R10925 DVDD.n9384 DVDD.n168 0.0183937
R10926 DVDD.n9386 DVDD.n171 0.0183937
R10927 DVDD.n9390 DVDD.n9389 0.0183937
R10928 DVDD.n9424 DVDD.n377 0.0183937
R10929 DVDD.n9423 DVDD.n378 0.0183937
R10930 DVDD.n9420 DVDD.n9419 0.0183937
R10931 DVDD.n386 DVDD.n381 0.0183937
R10932 DVDD.n4523 DVDD.n4522 0.0183937
R10933 DVDD.n4524 DVDD.n4520 0.0183937
R10934 DVDD.n8814 DVDD.n67 0.0183937
R10935 DVDD.n3854 DVDD.n3817 0.0183937
R10936 DVDD.n6534 DVDD.n3333 0.0183937
R10937 DVDD.n6502 DVDD.n2087 0.0183937
R10938 DVDD.n9086 DVDD.n529 0.0183937
R10939 DVDD.n6014 DVDD.n3957 0.0183937
R10940 DVDD.n6675 DVDD.n3236 0.0183937
R10941 DVDD.n3265 DVDD.n2139 0.0183937
R10942 DVDD.n4929 DVDD.n491 0.0183937
R10943 DVDD.n5781 DVDD.n4386 0.0183937
R10944 DVDD.n3131 DVDD.n3098 0.0183937
R10945 DVDD.n3156 DVDD.n2184 0.0183937
R10946 DVDD.n9255 DVDD.n9246 0.0183937
R10947 DVDD.n2841 DVDD.n2818 0.0183937
R10948 DVDD.n2719 DVDD.n2674 0.0183937
R10949 DVDD.n2686 DVDD.n2631 0.0183937
R10950 DVDD.n8820 DVDD.n64 0.0180394
R10951 DVDD.n3818 DVDD.n3562 0.0180394
R10952 DVDD.n6528 DVDD.n3355 0.0180394
R10953 DVDD.n6496 DVDD.n2077 0.0180394
R10954 DVDD.n9092 DVDD.n530 0.0180394
R10955 DVDD.n6008 DVDD.n3959 0.0180394
R10956 DVDD.n3292 DVDD.n3225 0.0180394
R10957 DVDD.n3259 DVDD.n2126 0.0180394
R10958 DVDD.n4935 DVDD.n488 0.0180394
R10959 DVDD.n4387 DVDD.n4306 0.0180394
R10960 DVDD.n3125 DVDD.n3120 0.0180394
R10961 DVDD.n3150 DVDD.n2174 0.0180394
R10962 DVDD.n9247 DVDD.n458 0.0180394
R10963 DVDD.n2835 DVDD.n2821 0.0180394
R10964 DVDD.n2713 DVDD.n2670 0.0180394
R10965 DVDD.n2680 DVDD.n2636 0.0180394
R10966 DVDD.n8450 DVDD.n8448 0.0179324
R10967 DVDD.n7719 DVDD.n1886 0.0178622
R10968 DVDD.n7724 DVDD.n1693 0.0178622
R10969 DVDD.n7701 DVDD.n1604 0.0178622
R10970 DVDD.n7694 DVDD.n1549 0.0178622
R10971 DVDD.n717 DVDD.n585 0.017685
R10972 DVDD.n71 DVDD.n60 0.017685
R10973 DVDD.n8739 DVDD.n880 0.017685
R10974 DVDD.n3635 DVDD.n1049 0.017685
R10975 DVDD.n3838 DVDD.n3566 0.017685
R10976 DVDD.n6518 DVDD.n2081 0.017685
R10977 DVDD.n8981 DVDD.n555 0.017685
R10978 DVDD.n9121 DVDD.n525 0.017685
R10979 DVDD.n4064 DVDD.n4028 0.017685
R10980 DVDD.n4160 DVDD.n4154 0.017685
R10981 DVDD.n6030 DVDD.n3963 0.017685
R10982 DVDD.n3281 DVDD.n2122 0.017685
R10983 DVDD.n5081 DVDD.n5027 0.017685
R10984 DVDD.n495 DVDD.n484 0.017685
R10985 DVDD.n9433 DVDD.n344 0.017685
R10986 DVDD.n9550 DVDD.n249 0.017685
R10987 DVDD.n5797 DVDD.n4310 0.017685
R10988 DVDD.n3172 DVDD.n2178 0.017685
R10989 DVDD.n5125 DVDD.n4577 0.017685
R10990 DVDD.n9278 DVDD.n464 0.017685
R10991 DVDD.n9585 DVDD.n173 0.017685
R10992 DVDD.n6782 DVDD.n2904 0.017685
R10993 DVDD.n2857 DVDD.n2825 0.017685
R10994 DVDD.n2702 DVDD.n2647 0.017685
R10995 DVDD.n9406 DVDD.n397 0.0174342
R10996 DVDD.n9603 DVDD.n9602 0.0174342
R10997 DVDD.n8709 DVDD.n901 0.0174342
R10998 DVDD.n1008 DVDD.n228 0.017375
R10999 DVDD.n9563 DVDD.n214 0.017375
R11000 DVDD.n9425 DVDD.n357 0.017375
R11001 DVDD.n3884 DVDD.n3880 0.017375
R11002 DVDD.n3878 DVDD.n3876 0.017375
R11003 DVDD.n6885 DVDD.n2785 0.017375
R11004 DVDD.n6884 DVDD.n2786 0.017375
R11005 DVDD.n9425 DVDD.n374 0.017375
R11006 DVDD.n399 DVDD.n200 0.017375
R11007 DVDD.n4511 DVDD.n228 0.017375
R11008 DVDD.n9563 DVDD.n225 0.017375
R11009 DVDD.n9616 DVDD.n109 0.017375
R11010 DVDD.n414 DVDD.n103 0.017375
R11011 DVDD.n899 DVDD.n200 0.017375
R11012 DVDD.n9618 DVDD.n103 0.017375
R11013 DVDD.n9617 DVDD.n9616 0.017375
R11014 DVDD.n8761 DVDD.n848 0.0173307
R11015 DVDD.n6260 DVDD.n3341 0.0173307
R11016 DVDD.n2409 DVDD.n1977 0.0173307
R11017 DVDD.n4036 DVDD.n4016 0.0173307
R11018 DVDD.n5951 DVDD.n3219 0.0173307
R11019 DVDD.n2416 DVDD.n2301 0.0173307
R11020 DVDD.n316 DVDD.n307 0.0173307
R11021 DVDD.n5849 DVDD.n3106 0.0173307
R11022 DVDD.n2422 DVDD.n2240 0.0173307
R11023 DVDD.n9611 DVDD.n133 0.0173307
R11024 DVDD.n6911 DVDD.n2735 0.0173307
R11025 DVDD.n2425 DVDD.n2381 0.0173307
R11026 DVDD.n588 DVDD.n583 0.0169764
R11027 DVDD.n842 DVDD.n91 0.0169764
R11028 DVDD.n3822 DVDD.n3810 0.0169764
R11029 DVDD.n3415 DVDD.n3349 0.0169764
R11030 DVDD.n9004 DVDD.n557 0.0169764
R11031 DVDD.n4012 DVDD.n4010 0.0169764
R11032 DVDD.n6046 DVDD.n3950 0.0169764
R11033 DVDD.n5943 DVDD.n3298 0.0169764
R11034 DVDD.n5010 DVDD.n4866 0.0169764
R11035 DVDD.n302 DVDD.n295 0.0169764
R11036 DVDD.n5813 DVDD.n4379 0.0169764
R11037 DVDD.n5841 DVDD.n3114 0.0169764
R11038 DVDD.n5148 DVDD.n4579 0.0169764
R11039 DVDD.n9312 DVDD.n9311 0.0169764
R11040 DVDD.n2874 DVDD.n2811 0.0169764
R11041 DVDD.n6903 DVDD.n2665 0.0169764
R11042 DVDD.n7090 DVDD.n7070 0.0168728
R11043 DVDD.n6243 DVDD.n6238 0.0166964
R11044 DVDD.n3869 DVDD.n3865 0.0166964
R11045 DVDD.n6898 DVDD.n2779 0.0166964
R11046 DVDD.n6868 DVDD.n2794 0.0166964
R11047 DVDD.n181 DVDD.n180 0.0166964
R11048 DVDD.n8675 DVDD.n8674 0.0166964
R11049 DVDD.n8692 DVDD.n1007 0.0166964
R11050 DVDD.n2916 DVDD.n2908 0.0166964
R11051 DVDD.n5277 DVDD.n5276 0.0166964
R11052 DVDD.n440 DVDD.n439 0.0166964
R11053 DVDD.n8724 DVDD.n875 0.0166964
R11054 DVDD.n8757 DVDD.n862 0.0166964
R11055 DVDD.n99 DVDD.n98 0.0166964
R11056 DVDD.n4756 DVDD.n4545 0.0166902
R11057 DVDD.n4708 DVDD.n4707 0.0166877
R11058 DVDD.n709 DVDD.n577 0.016622
R11059 DVDD.n81 DVDD.n79 0.016622
R11060 DVDD.n918 DVDD.n896 0.016622
R11061 DVDD.n3830 DVDD.n3811 0.016622
R11062 DVDD.n2432 DVDD.n1966 0.016622
R11063 DVDD.n9012 DVDD.n8976 0.016622
R11064 DVDD.n4113 DVDD.n4112 0.016622
R11065 DVDD.n4122 DVDD.n3993 0.016622
R11066 DVDD.n6038 DVDD.n3951 0.016622
R11067 DVDD.n2439 DVDD.n2323 0.016622
R11068 DVDD.n5018 DVDD.n4865 0.016622
R11069 DVDD.n9473 DVDD.n9472 0.016622
R11070 DVDD.n9482 DVDD.n283 0.016622
R11071 DVDD.n5805 DVDD.n4380 0.016622
R11072 DVDD.n2445 DVDD.n2229 0.016622
R11073 DVDD.n5156 DVDD.n5120 0.016622
R11074 DVDD.n9303 DVDD.n431 0.016622
R11075 DVDD.n9414 DVDD.n387 0.016622
R11076 DVDD.n2865 DVDD.n2812 0.016622
R11077 DVDD.n2448 DVDD.n2395 0.016622
R11078 DVDD.n6466 DVDD.n6465 0.0165042
R11079 DVDD.n8754 DVDD.n865 0.0162677
R11080 DVDD.n6268 DVDD.n3342 0.0162677
R11081 DVDD.n6488 DVDD.n2090 0.0162677
R11082 DVDD.n4048 DVDD.n4047 0.0162677
R11083 DVDD.n5959 DVDD.n3233 0.0162677
R11084 DVDD.n3251 DVDD.n2136 0.0162677
R11085 DVDD.n9447 DVDD.n315 0.0162677
R11086 DVDD.n5857 DVDD.n3107 0.0162677
R11087 DVDD.n3142 DVDD.n2187 0.0162677
R11088 DVDD.n144 DVDD.n142 0.0162677
R11089 DVDD.n6919 DVDD.n2736 0.0162677
R11090 DVDD.n6928 DVDD.n2642 0.0162677
R11091 DVDD.n6374 DVDD.n3531 0.0161276
R11092 DVDD.n6372 DVDD.n3537 0.0161276
R11093 DVDD.n6370 DVDD.n3530 0.0161276
R11094 DVDD.n6368 DVDD.n3538 0.0161276
R11095 DVDD.n6366 DVDD.n3529 0.0161276
R11096 DVDD.n6364 DVDD.n3539 0.0161276
R11097 DVDD.n6362 DVDD.n3528 0.0161276
R11098 DVDD.n6360 DVDD.n3540 0.0161276
R11099 DVDD.n6358 DVDD.n3527 0.0161276
R11100 DVDD.n6356 DVDD.n3541 0.0161276
R11101 DVDD.n6354 DVDD.n3526 0.0161276
R11102 DVDD.n6352 DVDD.n3542 0.0161276
R11103 DVDD.n6350 DVDD.n3525 0.0161276
R11104 DVDD.n6348 DVDD.n3543 0.0161276
R11105 DVDD.n6346 DVDD.n3524 0.0161276
R11106 DVDD.n6344 DVDD.n3544 0.0161276
R11107 DVDD.n6342 DVDD.n3523 0.0161276
R11108 DVDD.n6340 DVDD.n3545 0.0161276
R11109 DVDD.n6338 DVDD.n3522 0.0161276
R11110 DVDD.n6398 DVDD.n3546 0.0161276
R11111 DVDD.n8415 DVDD.n1489 0.0160585
R11112 DVDD.n8468 DVDD.n8441 0.0160585
R11113 DVDD.n1382 DVDD.n1381 0.0160585
R11114 DVDD.n8493 DVDD.n1438 0.0160585
R11115 DVDD.n8558 DVDD.n8557 0.0160585
R11116 DVDD.n8602 DVDD.n1348 0.0160585
R11117 DVDD.n8806 DVDD.n61 0.0159134
R11118 DVDD.n8745 DVDD.n874 0.0159134
R11119 DVDD.n8681 DVDD.n1041 0.0159134
R11120 DVDD.n3846 DVDD.n3565 0.0159134
R11121 DVDD.n6323 DVDD.n6321 0.0159134
R11122 DVDD.n6542 DVDD.n3352 0.0159134
R11123 DVDD.n6510 DVDD.n2080 0.0159134
R11124 DVDD.n8053 DVDD.n1983 0.0159134
R11125 DVDD.n9078 DVDD.n521 0.0159134
R11126 DVDD.n4058 DVDD.n4057 0.0159134
R11127 DVDD.n4217 DVDD.n4216 0.0159134
R11128 DVDD.n6022 DVDD.n3962 0.0159134
R11129 DVDD.n6057 DVDD.n5930 0.0159134
R11130 DVDD.n3248 DVDD.n3230 0.0159134
R11131 DVDD.n3273 DVDD.n2123 0.0159134
R11132 DVDD.n2306 DVDD.n2293 0.0159134
R11133 DVDD.n4921 DVDD.n485 0.0159134
R11134 DVDD.n340 DVDD.n339 0.0159134
R11135 DVDD.n9508 DVDD.n9507 0.0159134
R11136 DVDD.n5789 DVDD.n4309 0.0159134
R11137 DVDD.n5824 DVDD.n5767 0.0159134
R11138 DVDD.n3139 DVDD.n3117 0.0159134
R11139 DVDD.n3164 DVDD.n2177 0.0159134
R11140 DVDD.n7777 DVDD.n2246 0.0159134
R11141 DVDD.n9263 DVDD.n461 0.0159134
R11142 DVDD.n9594 DVDD.n156 0.0159134
R11143 DVDD.n6793 DVDD.n6792 0.0159134
R11144 DVDD.n2849 DVDD.n2824 0.0159134
R11145 DVDD.n6862 DVDD.n6861 0.0159134
R11146 DVDD.n6926 DVDD.n2655 0.0159134
R11147 DVDD.n2694 DVDD.n2645 0.0159134
R11148 DVDD.n7677 DVDD.n2386 0.0159134
R11149 DVDD.n1043 DVDD.n228 0.015575
R11150 DVDD.n9563 DVDD.n217 0.015575
R11151 DVDD.n9425 DVDD.n348 0.015575
R11152 DVDD.n3884 DVDD.n3872 0.015575
R11153 DVDD.n3876 DVDD.n3873 0.015575
R11154 DVDD.n6879 DVDD.n2785 0.015575
R11155 DVDD.n6880 DVDD.n2786 0.015575
R11156 DVDD.n9425 DVDD.n376 0.015575
R11157 DVDD.n200 DVDD.n177 0.015575
R11158 DVDD.n2890 DVDD.n228 0.015575
R11159 DVDD.n9563 DVDD.n224 0.015575
R11160 DVDD.n9616 DVDD.n110 0.015575
R11161 DVDD.n9352 DVDD.n103 0.015575
R11162 DVDD.n8728 DVDD.n200 0.015575
R11163 DVDD.n858 DVDD.n103 0.015575
R11164 DVDD.n9616 DVDD.n118 0.015575
R11165 DVDD.n5658 DVDD.n5481 0.0155591
R11166 DVDD.n8812 DVDD.n63 0.0155591
R11167 DVDD.n3852 DVDD.n3563 0.0155591
R11168 DVDD.n6536 DVDD.n3354 0.0155591
R11169 DVDD.n6504 DVDD.n2078 0.0155591
R11170 DVDD.n9084 DVDD.n524 0.0155591
R11171 DVDD.n6016 DVDD.n3960 0.0155591
R11172 DVDD.n3242 DVDD.n3215 0.0155591
R11173 DVDD.n3267 DVDD.n2125 0.0155591
R11174 DVDD.n4927 DVDD.n487 0.0155591
R11175 DVDD.n5783 DVDD.n4307 0.0155591
R11176 DVDD.n3133 DVDD.n3119 0.0155591
R11177 DVDD.n3158 DVDD.n2175 0.0155591
R11178 DVDD.n9257 DVDD.n463 0.0155591
R11179 DVDD.n2843 DVDD.n2822 0.0155591
R11180 DVDD.n2722 DVDD.n2669 0.0155591
R11181 DVDD.n2688 DVDD.n2648 0.0155591
R11182 DVDD.n5421 DVDD.n4482 0.0152047
R11183 DVDD.n5431 DVDD.n5423 0.0152047
R11184 DVDD.n5433 DVDD.n4481 0.0152047
R11185 DVDD.n5435 DVDD.n5424 0.0152047
R11186 DVDD.n5437 DVDD.n4480 0.0152047
R11187 DVDD.n5439 DVDD.n5425 0.0152047
R11188 DVDD.n5441 DVDD.n4479 0.0152047
R11189 DVDD.n5443 DVDD.n5426 0.0152047
R11190 DVDD.n5445 DVDD.n4478 0.0152047
R11191 DVDD.n5447 DVDD.n5427 0.0152047
R11192 DVDD.n5449 DVDD.n4477 0.0152047
R11193 DVDD.n5451 DVDD.n5428 0.0152047
R11194 DVDD.n5453 DVDD.n4476 0.0152047
R11195 DVDD.n5455 DVDD.n5429 0.0152047
R11196 DVDD.n5457 DVDD.n4475 0.0152047
R11197 DVDD.n5459 DVDD.n5430 0.0152047
R11198 DVDD.n5461 DVDD.n4474 0.0152047
R11199 DVDD.n5465 DVDD.n5464 0.0152047
R11200 DVDD.n5467 DVDD.n4469 0.0152047
R11201 DVDD.n5468 DVDD.n4467 0.0152047
R11202 DVDD.n8823 DVDD.n66 0.0152047
R11203 DVDD.n6333 DVDD.n6332 0.0152047
R11204 DVDD.n3356 DVDD.n3332 0.0152047
R11205 DVDD.n6494 DVDD.n2088 0.0152047
R11206 DVDD.n9094 DVDD.n523 0.0152047
R11207 DVDD.n6006 DVDD.n3958 0.0152047
R11208 DVDD.n3290 DVDD.n3228 0.0152047
R11209 DVDD.n3257 DVDD.n2138 0.0152047
R11210 DVDD.n4938 DVDD.n490 0.0152047
R11211 DVDD.n6112 DVDD.n4389 0.0152047
R11212 DVDD.n3121 DVDD.n3097 0.0152047
R11213 DVDD.n3148 DVDD.n2185 0.0152047
R11214 DVDD.n9286 DVDD.n9285 0.0152047
R11215 DVDD.n2833 DVDD.n2819 0.0152047
R11216 DVDD.n2711 DVDD.n2673 0.0152047
R11217 DVDD.n2678 DVDD.n2643 0.0152047
R11218 DVDD.n7710 DVDD.n1861 0.0150276
R11219 DVDD.n7703 DVDD.n1664 0.0150276
R11220 DVDD.n7697 DVDD.n1595 0.0150276
R11221 DVDD.n7690 DVDD.n1540 0.0150276
R11222 DVDD.n715 DVDD.n580 0.0148504
R11223 DVDD.n9646 DVDD.n9645 0.0148504
R11224 DVDD.n8734 DVDD.n8723 0.0148504
R11225 DVDD.n8671 DVDD.n1050 0.0148504
R11226 DVDD.n3836 DVDD.n3813 0.0148504
R11227 DVDD.n6520 DVDD.n2083 0.0148504
R11228 DVDD.n1866 DVDD.n1865 0.0148504
R11229 DVDD.n8983 DVDD.n8974 0.0148504
R11230 DVDD.n9119 DVDD.n527 0.0148504
R11231 DVDD.n4078 DVDD.n4077 0.0148504
R11232 DVDD.n4206 DVDD.n4205 0.0148504
R11233 DVDD.n6032 DVDD.n3953 0.0148504
R11234 DVDD.n3283 DVDD.n2143 0.0148504
R11235 DVDD.n1677 DVDD.n1661 0.0148504
R11236 DVDD.n5024 DVDD.n4863 0.0148504
R11237 DVDD.n9209 DVDD.n497 0.0148504
R11238 DVDD.n9432 DVDD.n345 0.0148504
R11239 DVDD.n9549 DVDD.n250 0.0148504
R11240 DVDD.n5799 DVDD.n4382 0.0148504
R11241 DVDD.n3174 DVDD.n2180 0.0148504
R11242 DVDD.n1874 DVDD.n1599 0.0148504
R11243 DVDD.n5127 DVDD.n5118 0.0148504
R11244 DVDD.n9276 DVDD.n9244 0.0148504
R11245 DVDD.n9393 DVDD.n9392 0.0148504
R11246 DVDD.n6781 DVDD.n2905 0.0148504
R11247 DVDD.n2859 DVDD.n2814 0.0148504
R11248 DVDD.n2704 DVDD.n2633 0.0148504
R11249 DVDD.n1561 DVDD.n1532 0.0148504
R11250 DVDD.n6556 DVDD.n3399 0.0146213
R11251 DVDD.n6554 DVDD.n6474 0.0146213
R11252 DVDD.n6552 DVDD.n3398 0.0146213
R11253 DVDD.n6550 DVDD.n6475 0.0146213
R11254 DVDD.n6548 DVDD.n3397 0.0146213
R11255 DVDD.n6546 DVDD.n6476 0.0146213
R11256 DVDD.n6544 DVDD.n3396 0.0146213
R11257 DVDD.n6604 DVDD.n6477 0.0146213
R11258 DVDD.n8767 DVDD.n8766 0.0144961
R11259 DVDD.n6336 DVDD.n3556 0.0144961
R11260 DVDD.n6258 DVDD.n3347 0.0144961
R11261 DVDD.n2410 DVDD.n1953 0.0144961
R11262 DVDD.n4097 DVDD.n4096 0.0144961
R11263 DVDD.n6052 DVDD.n3948 0.0144961
R11264 DVDD.n5949 DVDD.n3231 0.0144961
R11265 DVDD.n2413 DVDD.n2289 0.0144961
R11266 DVDD.n9459 DVDD.n9458 0.0144961
R11267 DVDD.n5819 DVDD.n4377 0.0144961
R11268 DVDD.n5847 DVDD.n3112 0.0144961
R11269 DVDD.n2419 DVDD.n2216 0.0144961
R11270 DVDD.n9612 DVDD.n131 0.0144961
R11271 DVDD.n6858 DVDD.n2803 0.0144961
R11272 DVDD.n6909 DVDD.n2663 0.0144961
R11273 DVDD.n2426 DVDD.n2404 0.0144961
R11274 DVDD.n8891 DVDD.n8889 0.0142903
R11275 DVDD.n8204 DVDD.n8203 0.0142903
R11276 DVDD.n9700 DVDD.n9699 0.0142808
R11277 DVDD.n6586 DVDD.n2042 0.0142448
R11278 DVDD.n6584 DVDD.n2044 0.0142448
R11279 DVDD.n6582 DVDD.n2041 0.0142448
R11280 DVDD.n6580 DVDD.n2045 0.0142448
R11281 DVDD.n6578 DVDD.n2040 0.0142448
R11282 DVDD.n6576 DVDD.n2046 0.0142448
R11283 DVDD.n6574 DVDD.n2039 0.0142448
R11284 DVDD.n6572 DVDD.n2047 0.0142448
R11285 DVDD.n6570 DVDD.n2038 0.0142448
R11286 DVDD.n6568 DVDD.n2048 0.0142448
R11287 DVDD.n6566 DVDD.n2037 0.0142448
R11288 DVDD.n6564 DVDD.n2049 0.0142448
R11289 DVDD.n6562 DVDD.n2036 0.0142448
R11290 DVDD.n6560 DVDD.n2050 0.0142448
R11291 DVDD.n6558 DVDD.n2035 0.0142448
R11292 DVDD.n6382 DVDD.n3474 0.0142224
R11293 DVDD.n7681 DVDD.n2354 0.0141679
R11294 DVDD.n7682 DVDD.n2357 0.0141679
R11295 DVDD.n2365 DVDD.n2360 0.0141679
R11296 DVDD.n2366 DVDD.n2362 0.0141679
R11297 DVDD.n7744 DVDD.n2334 0.0141679
R11298 DVDD.n7741 DVDD.n2334 0.0141679
R11299 DVDD.n7738 DVDD.n2333 0.0141679
R11300 DVDD.n7731 DVDD.n2337 0.0141679
R11301 DVDD.n7732 DVDD.n2339 0.0141679
R11302 DVDD.n7744 DVDD.n7743 0.0141679
R11303 DVDD.n7740 DVDD.n2333 0.0141679
R11304 DVDD.n7736 DVDD.n2337 0.0141679
R11305 DVDD.n7741 DVDD.n7740 0.0141679
R11306 DVDD.n2340 DVDD.n2339 0.0141679
R11307 DVDD.n7688 DVDD.n2352 0.0141679
R11308 DVDD.n7691 DVDD.n2352 0.0141679
R11309 DVDD.n7692 DVDD.n2351 0.0141679
R11310 DVDD.n2351 DVDD.n2349 0.0141679
R11311 DVDD.n2348 DVDD.n2347 0.0141679
R11312 DVDD.n7698 DVDD.n2348 0.0141679
R11313 DVDD.n7699 DVDD.n2346 0.0141679
R11314 DVDD.n2346 DVDD.n2344 0.0141679
R11315 DVDD.n7706 DVDD.n7704 0.0141679
R11316 DVDD.n7707 DVDD.n7706 0.0141679
R11317 DVDD.n7721 DVDD.n7705 0.0141679
R11318 DVDD.n7709 DVDD.n7705 0.0141679
R11319 DVDD.n7714 DVDD.n7711 0.0141679
R11320 DVDD.n7715 DVDD.n7714 0.0141679
R11321 DVDD.n7717 DVDD.n7713 0.0141679
R11322 DVDD.n7713 DVDD.n7712 0.0141679
R11323 DVDD.n7725 DVDD.n7704 0.0141679
R11324 DVDD.n7721 DVDD.n7708 0.0141679
R11325 DVDD.n7720 DVDD.n7711 0.0141679
R11326 DVDD.n7718 DVDD.n7717 0.0141679
R11327 DVDD.n7708 DVDD.n7707 0.0141679
R11328 DVDD.n7723 DVDD.n7709 0.0141679
R11329 DVDD.n7718 DVDD.n7715 0.0141679
R11330 DVDD.n7712 DVDD.n2341 0.0141679
R11331 DVDD.n7700 DVDD.n7699 0.0141679
R11332 DVDD.n7700 DVDD.n7698 0.0141679
R11333 DVDD.n7702 DVDD.n2344 0.0141679
R11334 DVDD.n7696 DVDD.n2347 0.0141679
R11335 DVDD.n2370 DVDD.n2360 0.0141679
R11336 DVDD.n2363 DVDD.n2362 0.0141679
R11337 DVDD.n7689 DVDD.n7688 0.0141679
R11338 DVDD.n7693 DVDD.n7692 0.0141679
R11339 DVDD.n7693 DVDD.n7691 0.0141679
R11340 DVDD.n7695 DVDD.n2349 0.0141679
R11341 DVDD.n7686 DVDD.n2354 0.0141679
R11342 DVDD.n2358 DVDD.n2357 0.0141679
R11343 DVDD.n8937 DVDD.n590 0.0141417
R11344 DVDD.n9622 DVDD.n92 0.0141417
R11345 DVDD.n3820 DVDD.n3570 0.0141417
R11346 DVDD.n6301 DVDD.n6300 0.0141417
R11347 DVDD.n6254 DVDD.n3339 0.0141417
R11348 DVDD.n9002 DVDD.n8972 0.0141417
R11349 DVDD.n4011 DVDD.n4002 0.0141417
R11350 DVDD.n6048 DVDD.n3967 0.0141417
R11351 DVDD.n5993 DVDD.n5992 0.0141417
R11352 DVDD.n5945 DVDD.n3216 0.0141417
R11353 DVDD.n5008 DVDD.n4858 0.0141417
R11354 DVDD.n9465 DVDD.n9464 0.0141417
R11355 DVDD.n5815 DVDD.n4314 0.0141417
R11356 DVDD.n5828 DVDD.n5760 0.0141417
R11357 DVDD.n5843 DVDD.n3104 0.0141417
R11358 DVDD.n5146 DVDD.n5116 0.0141417
R11359 DVDD.n444 DVDD.n410 0.0141417
R11360 DVDD.n2875 DVDD.n2829 0.0141417
R11361 DVDD.n6901 DVDD.n2742 0.0141417
R11362 DVDD.n6905 DVDD.n2733 0.0141417
R11363 DVDD.n3499 DVDD.n3491 0.0141393
R11364 DVDD.n3499 DVDD.n3488 0.0141393
R11365 DVDD.n6447 DVDD.n3488 0.0141393
R11366 DVDD.n6454 DVDD.n3486 0.0141393
R11367 DVDD.n6454 DVDD.n3484 0.0141393
R11368 DVDD.n6458 DVDD.n3484 0.0141393
R11369 DVDD.n1465 DVDD.n1464 0.0138885
R11370 DVDD.n8424 DVDD.n8422 0.0138885
R11371 DVDD.n8432 DVDD.n8431 0.0138885
R11372 DVDD.n8437 DVDD.n8436 0.0138885
R11373 DVDD.n1470 DVDD.n1469 0.0138885
R11374 DVDD.n8506 DVDD.n1417 0.0138885
R11375 DVDD.n8500 DVDD.n1423 0.0138885
R11376 DVDD.n8496 DVDD.n1431 0.0138885
R11377 DVDD.n1476 DVDD.n1475 0.0138885
R11378 DVDD.n8512 DVDD.n1411 0.0138885
R11379 DVDD.n1366 DVDD.n1365 0.0138885
R11380 DVDD.n1357 DVDD.n1356 0.0138885
R11381 DVDD.n8438 DVDD.n8437 0.0138885
R11382 DVDD.n8497 DVDD.n8496 0.0138885
R11383 DVDD.n8597 DVDD.n1356 0.0138885
R11384 DVDD.n8433 DVDD.n8432 0.0138885
R11385 DVDD.n8501 DVDD.n8500 0.0138885
R11386 DVDD.n8592 DVDD.n1365 0.0138885
R11387 DVDD.n8422 DVDD.n8421 0.0138885
R11388 DVDD.n8507 DVDD.n8506 0.0138885
R11389 DVDD.n8513 DVDD.n8512 0.0138885
R11390 DVDD.n8416 DVDD.n1464 0.0138885
R11391 DVDD.n1485 DVDD.n1469 0.0138885
R11392 DVDD.n1475 DVDD.n1393 0.0138885
R11393 DVDD.n8420 DVDD.n1460 0.0138885
R11394 DVDD.n8428 DVDD.n1456 0.0138885
R11395 DVDD.n8435 DVDD.n1451 0.0138885
R11396 DVDD.n8440 DVDD.n1446 0.0138885
R11397 DVDD.n1484 DVDD.n1415 0.0138885
R11398 DVDD.n8504 DVDD.n1413 0.0138885
R11399 DVDD.n8498 DVDD.n1428 0.0138885
R11400 DVDD.n8494 DVDD.n1436 0.0138885
R11401 DVDD.n1480 DVDD.n1409 0.0138885
R11402 DVDD.n1407 DVDD.n1370 0.0138885
R11403 DVDD.n8596 DVDD.n1361 0.0138885
R11404 DVDD.n8601 DVDD.n1352 0.0138885
R11405 DVDD.n1449 DVDD.n1446 0.0138885
R11406 DVDD.n1436 DVDD.n1435 0.0138885
R11407 DVDD.n1358 DVDD.n1352 0.0138885
R11408 DVDD.n1454 DVDD.n1451 0.0138885
R11409 DVDD.n1428 DVDD.n1427 0.0138885
R11410 DVDD.n1367 DVDD.n1361 0.0138885
R11411 DVDD.n8425 DVDD.n1456 0.0138885
R11412 DVDD.n1419 DVDD.n1413 0.0138885
R11413 DVDD.n8509 DVDD.n1407 0.0138885
R11414 DVDD.n1466 DVDD.n1460 0.0138885
R11415 DVDD.n1484 DVDD.n1472 0.0138885
R11416 DVDD.n1480 DVDD.n1478 0.0138885
R11417 DVDD.n5560 DVDD.n5500 0.0137874
R11418 DVDD.n5567 DVDD.n5562 0.0137874
R11419 DVDD.n5569 DVDD.n5499 0.0137874
R11420 DVDD.n5571 DVDD.n5563 0.0137874
R11421 DVDD.n5573 DVDD.n5498 0.0137874
R11422 DVDD.n5575 DVDD.n5564 0.0137874
R11423 DVDD.n5577 DVDD.n5497 0.0137874
R11424 DVDD.n5613 DVDD.n5565 0.0137874
R11425 DVDD.n711 DVDD.n587 0.0137874
R11426 DVDD.n8714 DVDD.n889 0.0137874
R11427 DVDD.n3832 DVDD.n3568 0.0137874
R11428 DVDD.n2433 DVDD.n1958 0.0137874
R11429 DVDD.n8987 DVDD.n553 0.0137874
R11430 DVDD.n4070 DVDD.n4069 0.0137874
R11431 DVDD.n6036 DVDD.n3965 0.0137874
R11432 DVDD.n2436 DVDD.n2290 0.0137874
R11433 DVDD.n5020 DVDD.n4860 0.0137874
R11434 DVDD.n366 DVDD.n365 0.0137874
R11435 DVDD.n5803 DVDD.n4312 0.0137874
R11436 DVDD.n2442 DVDD.n2221 0.0137874
R11437 DVDD.n5131 DVDD.n4575 0.0137874
R11438 DVDD.n9397 DVDD.n382 0.0137874
R11439 DVDD.n2863 DVDD.n2827 0.0137874
R11440 DVDD.n2449 DVDD.n2427 0.0137874
R11441 DVDD.n3441 DVDD.n3407 0.0134916
R11442 DVDD.n3439 DVDD.n3409 0.0134916
R11443 DVDD.n3437 DVDD.n3406 0.0134916
R11444 DVDD.n3435 DVDD.n3410 0.0134916
R11445 DVDD.n3433 DVDD.n3405 0.0134916
R11446 DVDD.n3431 DVDD.n3411 0.0134916
R11447 DVDD.n3429 DVDD.n3404 0.0134916
R11448 DVDD.n3413 DVDD.n3412 0.0134916
R11449 DVDD.n6469 DVDD.n3403 0.0134916
R11450 DVDD.n5606 DVDD.n2535 0.0134331
R11451 DVDD.n5604 DVDD.n2537 0.0134331
R11452 DVDD.n5602 DVDD.n2534 0.0134331
R11453 DVDD.n5600 DVDD.n2538 0.0134331
R11454 DVDD.n5598 DVDD.n2533 0.0134331
R11455 DVDD.n5596 DVDD.n2539 0.0134331
R11456 DVDD.n5594 DVDD.n2532 0.0134331
R11457 DVDD.n5592 DVDD.n2540 0.0134331
R11458 DVDD.n5590 DVDD.n2531 0.0134331
R11459 DVDD.n5588 DVDD.n2541 0.0134331
R11460 DVDD.n5586 DVDD.n2530 0.0134331
R11461 DVDD.n5584 DVDD.n2542 0.0134331
R11462 DVDD.n5582 DVDD.n2529 0.0134331
R11463 DVDD.n5580 DVDD.n2543 0.0134331
R11464 DVDD.n2651 DVDD.n2528 0.0134331
R11465 DVDD.n935 DVDD.n933 0.0134331
R11466 DVDD.n6270 DVDD.n3345 0.0134331
R11467 DVDD.n6490 DVDD.n2075 0.0134331
R11468 DVDD.n4051 DVDD.n4034 0.0134331
R11469 DVDD.n5961 DVDD.n3218 0.0134331
R11470 DVDD.n3253 DVDD.n2128 0.0134331
R11471 DVDD.n9446 DVDD.n321 0.0134331
R11472 DVDD.n5859 DVDD.n3110 0.0134331
R11473 DVDD.n3144 DVDD.n2172 0.0134331
R11474 DVDD.n9600 DVDD.n143 0.0134331
R11475 DVDD.n6922 DVDD.n2661 0.0134331
R11476 DVDD.n6931 DVDD.n2630 0.0134331
R11477 DVDD.n8680 DVDD.n1043 0.013325
R11478 DVDD.n8733 DVDD.n348 0.013325
R11479 DVDD.n6315 DVDD.n3873 0.013325
R11480 DVDD.n6879 DVDD.n6878 0.013325
R11481 DVDD.n376 DVDD.n175 0.013325
R11482 DVDD.n2891 DVDD.n2890 0.013325
R11483 DVDD.n132 DVDD.n110 0.013325
R11484 DVDD.n849 DVDD.n118 0.013325
R11485 DVDD.n8808 DVDD.n69 0.0130787
R11486 DVDD.n8748 DVDD.n873 0.0130787
R11487 DVDD.n1040 DVDD.n1010 0.0130787
R11488 DVDD.n3848 DVDD.n3815 0.0130787
R11489 DVDD.n6324 DVDD.n3863 0.0130787
R11490 DVDD.n6540 DVDD.n3335 0.0130787
R11491 DVDD.n6508 DVDD.n2085 0.0130787
R11492 DVDD.n7664 DVDD.n1949 0.0130787
R11493 DVDD.n9080 DVDD.n531 0.0130787
R11494 DVDD.n4053 DVDD.n4032 0.0130787
R11495 DVDD.n4219 DVDD.n4218 0.0130787
R11496 DVDD.n6020 DVDD.n3955 0.0130787
R11497 DVDD.n6060 DVDD.n5923 0.0130787
R11498 DVDD.n3246 DVDD.n3224 0.0130787
R11499 DVDD.n3271 DVDD.n2141 0.0130787
R11500 DVDD.n7748 DVDD.n2291 0.0130787
R11501 DVDD.n4923 DVDD.n493 0.0130787
R11502 DVDD.n338 DVDD.n336 0.0130787
R11503 DVDD.n9510 DVDD.n9509 0.0130787
R11504 DVDD.n5787 DVDD.n4384 0.0130787
R11505 DVDD.n5769 DVDD.n5764 0.0130787
R11506 DVDD.n3137 DVDD.n3100 0.0130787
R11507 DVDD.n3162 DVDD.n2182 0.0130787
R11508 DVDD.n7673 DVDD.n2212 0.0130787
R11509 DVDD.n9261 DVDD.n9248 0.0130787
R11510 DVDD.n9595 DVDD.n154 0.0130787
R11511 DVDD.n6795 DVDD.n6794 0.0130787
R11512 DVDD.n2847 DVDD.n2816 0.0130787
R11513 DVDD.n6865 DVDD.n2798 0.0130787
R11514 DVDD.n6925 DVDD.n2658 0.0130787
R11515 DVDD.n2692 DVDD.n2635 0.0130787
R11516 DVDD.n7678 DVDD.n2450 0.0130787
R11517 DVDD.n7199 DVDD.n7198 0.0128916
R11518 DVDD.n7195 DVDD.n7193 0.0128916
R11519 DVDD.n7196 DVDD.n7192 0.0128916
R11520 DVDD.n7191 DVDD.n7139 0.0128916
R11521 DVDD.n7141 DVDD.n7140 0.0128916
R11522 DVDD.n7188 DVDD.n7140 0.0128916
R11523 DVDD.n7148 DVDD.n7144 0.0128916
R11524 DVDD.n7147 DVDD.n7146 0.0128916
R11525 DVDD.n7184 DVDD.n7150 0.0128916
R11526 DVDD.n7182 DVDD.n7153 0.0128916
R11527 DVDD.n7155 DVDD.n7154 0.0128916
R11528 DVDD.n7179 DVDD.n7154 0.0128916
R11529 DVDD.n7177 DVDD.n7159 0.0128916
R11530 DVDD.n7161 DVDD.n7160 0.0128916
R11531 DVDD.n7174 DVDD.n7160 0.0128916
R11532 DVDD.n7170 DVDD.n7163 0.0128916
R11533 DVDD.n7169 DVDD.n7168 0.0128916
R11534 DVDD.n7167 DVDD.n1303 0.0128916
R11535 DVDD.n7186 DVDD.n7144 0.0128916
R11536 DVDD.n7150 DVDD.n7146 0.0128916
R11537 DVDD.n7156 DVDD.n7155 0.0128916
R11538 DVDD.n7162 DVDD.n7161 0.0128916
R11539 DVDD.n7148 DVDD.n7147 0.0128916
R11540 DVDD.n7156 DVDD.n7153 0.0128916
R11541 DVDD.n7180 DVDD.n7179 0.0128916
R11542 DVDD.n7162 DVDD.n7159 0.0128916
R11543 DVDD.n7175 DVDD.n7174 0.0128916
R11544 DVDD.n8384 DVDD.n8383 0.0128916
R11545 DVDD.n8380 DVDD.n1499 0.0128916
R11546 DVDD.n8381 DVDD.n8379 0.0128916
R11547 DVDD.n1507 DVDD.n1504 0.0128916
R11548 DVDD.n8374 DVDD.n8373 0.0128916
R11549 DVDD.n8375 DVDD.n8374 0.0128916
R11550 DVDD.n7343 DVDD.n1508 0.0128916
R11551 DVDD.n8638 DVDD.n1307 0.0128916
R11552 DVDD.n8633 DVDD.n1315 0.0128916
R11553 DVDD.n1299 DVDD.n1298 0.0128916
R11554 DVDD.n1301 DVDD.n1295 0.0128916
R11555 DVDD.n8645 DVDD.n1300 0.0128916
R11556 DVDD.n7362 DVDD.n7343 0.0128916
R11557 DVDD.n1311 DVDD.n1307 0.0128916
R11558 DVDD.n1319 DVDD.n1315 0.0128916
R11559 DVDD.n8378 DVDD.n1504 0.0128916
R11560 DVDD.n8373 DVDD.n1507 0.0128916
R11561 DVDD.n8376 DVDD.n8375 0.0128916
R11562 DVDD.n7142 DVDD.n7141 0.0128916
R11563 DVDD.n7142 DVDD.n7139 0.0128916
R11564 DVDD.n7189 DVDD.n7188 0.0128916
R11565 DVDD.n1301 DVDD.n1299 0.0128916
R11566 DVDD.n1298 DVDD.n1296 0.0128916
R11567 DVDD.n1300 DVDD.n1295 0.0128916
R11568 DVDD.n7170 DVDD.n7169 0.0128916
R11569 DVDD.n7172 DVDD.n7163 0.0128916
R11570 DVDD.n7168 DVDD.n7167 0.0128916
R11571 DVDD.n8383 DVDD.n1499 0.0128916
R11572 DVDD.n8381 DVDD.n8380 0.0128916
R11573 DVDD.n7198 DVDD.n7193 0.0128916
R11574 DVDD.n7196 DVDD.n7195 0.0128916
R11575 DVDD.n7200 DVDD.n7199 0.0128916
R11576 DVDD.n8385 DVDD.n8384 0.0128916
R11577 DVDD.n6380 DVDD.n3472 0.0127385
R11578 DVDD.n6378 DVDD.n3475 0.0127385
R11579 DVDD.n6376 DVDD.n3471 0.0127385
R11580 DVDD.n5615 DVDD.n5494 0.0127244
R11581 DVDD.n5536 DVDD.n5531 0.0127244
R11582 DVDD.n5538 DVDD.n5507 0.0127244
R11583 DVDD.n5540 DVDD.n5532 0.0127244
R11584 DVDD.n5542 DVDD.n5506 0.0127244
R11585 DVDD.n5544 DVDD.n5533 0.0127244
R11586 DVDD.n5534 DVDD.n5505 0.0127244
R11587 DVDD.n5549 DVDD.n5548 0.0127244
R11588 DVDD.n5550 DVDD.n5504 0.0127244
R11589 DVDD.n8810 DVDD.n68 0.0127244
R11590 DVDD.n3850 DVDD.n3816 0.0127244
R11591 DVDD.n6538 DVDD.n3334 0.0127244
R11592 DVDD.n6506 DVDD.n2086 0.0127244
R11593 DVDD.n9082 DVDD.n528 0.0127244
R11594 DVDD.n6018 DVDD.n3956 0.0127244
R11595 DVDD.n3244 DVDD.n3235 0.0127244
R11596 DVDD.n3269 DVDD.n2140 0.0127244
R11597 DVDD.n4925 DVDD.n492 0.0127244
R11598 DVDD.n5785 DVDD.n4385 0.0127244
R11599 DVDD.n3135 DVDD.n3099 0.0127244
R11600 DVDD.n3160 DVDD.n2183 0.0127244
R11601 DVDD.n9259 DVDD.n9245 0.0127244
R11602 DVDD.n2845 DVDD.n2817 0.0127244
R11603 DVDD.n2723 DVDD.n2675 0.0127244
R11604 DVDD.n2690 DVDD.n2632 0.0127244
R11605 DVDD.n1796 DVDD.n1789 0.0126434
R11606 DVDD.n8199 DVDD.n8194 0.0126434
R11607 DVDD.n1795 DVDD.n1788 0.0126434
R11608 DVDD.n8198 DVDD.n8195 0.0126434
R11609 DVDD.n1794 DVDD.n1787 0.0126434
R11610 DVDD.n8197 DVDD.n8196 0.0126434
R11611 DVDD.n1793 DVDD.n1786 0.0126434
R11612 DVDD.n8207 DVDD.n8206 0.0126434
R11613 DVDD.n1792 DVDD.n1785 0.0126434
R11614 DVDD.n8209 DVDD.n1791 0.0126434
R11615 DVDD.n8193 DVDD.n1789 0.0126434
R11616 DVDD.n8199 DVDD.n1796 0.0126434
R11617 DVDD.n8194 DVDD.n1788 0.0126434
R11618 DVDD.n8198 DVDD.n1795 0.0126434
R11619 DVDD.n8195 DVDD.n1787 0.0126434
R11620 DVDD.n8197 DVDD.n1794 0.0126434
R11621 DVDD.n8196 DVDD.n1786 0.0126434
R11622 DVDD.n8206 DVDD.n1793 0.0126434
R11623 DVDD.n8207 DVDD.n1785 0.0126434
R11624 DVDD.n1792 DVDD.n1791 0.0126434
R11625 DVDD.n8177 DVDD.n1816 0.0126434
R11626 DVDD.n1815 DVDD.n1812 0.0126434
R11627 DVDD.n8178 DVDD.n1818 0.0126434
R11628 DVDD.n1817 DVDD.n1811 0.0126434
R11629 DVDD.n8179 DVDD.n1820 0.0126434
R11630 DVDD.n1819 DVDD.n1810 0.0126434
R11631 DVDD.n8180 DVDD.n1822 0.0126434
R11632 DVDD.n1821 DVDD.n1809 0.0126434
R11633 DVDD.n8181 DVDD.n1824 0.0126434
R11634 DVDD.n1823 DVDD.n1808 0.0126434
R11635 DVDD.n8182 DVDD.n1826 0.0126434
R11636 DVDD.n1825 DVDD.n1807 0.0126434
R11637 DVDD.n8183 DVDD.n1828 0.0126434
R11638 DVDD.n1827 DVDD.n1806 0.0126434
R11639 DVDD.n8184 DVDD.n1830 0.0126434
R11640 DVDD.n1829 DVDD.n1805 0.0126434
R11641 DVDD.n8185 DVDD.n1832 0.0126434
R11642 DVDD.n1831 DVDD.n1804 0.0126434
R11643 DVDD.n8186 DVDD.n1834 0.0126434
R11644 DVDD.n1833 DVDD.n1803 0.0126434
R11645 DVDD.n8190 DVDD.n8188 0.0126434
R11646 DVDD.n8189 DVDD.n1802 0.0126434
R11647 DVDD.n8192 DVDD.n1798 0.0126434
R11648 DVDD.n8177 DVDD.n1813 0.0126434
R11649 DVDD.n1816 DVDD.n1815 0.0126434
R11650 DVDD.n8178 DVDD.n1812 0.0126434
R11651 DVDD.n1818 DVDD.n1817 0.0126434
R11652 DVDD.n8179 DVDD.n1811 0.0126434
R11653 DVDD.n1820 DVDD.n1819 0.0126434
R11654 DVDD.n8180 DVDD.n1810 0.0126434
R11655 DVDD.n1822 DVDD.n1821 0.0126434
R11656 DVDD.n8181 DVDD.n1809 0.0126434
R11657 DVDD.n1824 DVDD.n1823 0.0126434
R11658 DVDD.n8182 DVDD.n1808 0.0126434
R11659 DVDD.n1826 DVDD.n1825 0.0126434
R11660 DVDD.n8183 DVDD.n1807 0.0126434
R11661 DVDD.n1828 DVDD.n1827 0.0126434
R11662 DVDD.n8184 DVDD.n1806 0.0126434
R11663 DVDD.n1830 DVDD.n1829 0.0126434
R11664 DVDD.n8185 DVDD.n1805 0.0126434
R11665 DVDD.n1832 DVDD.n1831 0.0126434
R11666 DVDD.n8186 DVDD.n1804 0.0126434
R11667 DVDD.n1834 DVDD.n1833 0.0126434
R11668 DVDD.n8188 DVDD.n1803 0.0126434
R11669 DVDD.n8190 DVDD.n8189 0.0126434
R11670 DVDD.n1802 DVDD.n1798 0.0126434
R11671 DVDD.n7986 DVDD.n7962 0.0126434
R11672 DVDD.n7984 DVDD.n2026 0.0126434
R11673 DVDD.n7987 DVDD.n7963 0.0126434
R11674 DVDD.n7983 DVDD.n2025 0.0126434
R11675 DVDD.n7988 DVDD.n7964 0.0126434
R11676 DVDD.n7982 DVDD.n2024 0.0126434
R11677 DVDD.n7989 DVDD.n7965 0.0126434
R11678 DVDD.n7981 DVDD.n2023 0.0126434
R11679 DVDD.n7990 DVDD.n7966 0.0126434
R11680 DVDD.n7980 DVDD.n2022 0.0126434
R11681 DVDD.n7991 DVDD.n7967 0.0126434
R11682 DVDD.n7979 DVDD.n2021 0.0126434
R11683 DVDD.n7992 DVDD.n7968 0.0126434
R11684 DVDD.n7978 DVDD.n2020 0.0126434
R11685 DVDD.n7993 DVDD.n7969 0.0126434
R11686 DVDD.n7977 DVDD.n2019 0.0126434
R11687 DVDD.n7994 DVDD.n7970 0.0126434
R11688 DVDD.n7976 DVDD.n2018 0.0126434
R11689 DVDD.n7995 DVDD.n7971 0.0126434
R11690 DVDD.n7975 DVDD.n2017 0.0126434
R11691 DVDD.n7996 DVDD.n7972 0.0126434
R11692 DVDD.n7974 DVDD.n2016 0.0126434
R11693 DVDD.n8009 DVDD.n7973 0.0126434
R11694 DVDD.n7986 DVDD.n7960 0.0126434
R11695 DVDD.n7984 DVDD.n7962 0.0126434
R11696 DVDD.n7987 DVDD.n2026 0.0126434
R11697 DVDD.n7983 DVDD.n7963 0.0126434
R11698 DVDD.n7988 DVDD.n2025 0.0126434
R11699 DVDD.n7982 DVDD.n7964 0.0126434
R11700 DVDD.n7989 DVDD.n2024 0.0126434
R11701 DVDD.n7981 DVDD.n7965 0.0126434
R11702 DVDD.n7990 DVDD.n2023 0.0126434
R11703 DVDD.n7980 DVDD.n7966 0.0126434
R11704 DVDD.n7991 DVDD.n2022 0.0126434
R11705 DVDD.n7979 DVDD.n7967 0.0126434
R11706 DVDD.n7992 DVDD.n2021 0.0126434
R11707 DVDD.n7978 DVDD.n7968 0.0126434
R11708 DVDD.n7993 DVDD.n2020 0.0126434
R11709 DVDD.n7977 DVDD.n7969 0.0126434
R11710 DVDD.n7994 DVDD.n2019 0.0126434
R11711 DVDD.n7976 DVDD.n7970 0.0126434
R11712 DVDD.n7995 DVDD.n2018 0.0126434
R11713 DVDD.n7975 DVDD.n7971 0.0126434
R11714 DVDD.n7996 DVDD.n2017 0.0126434
R11715 DVDD.n7974 DVDD.n7972 0.0126434
R11716 DVDD.n7973 DVDD.n2016 0.0126434
R11717 DVDD.n2051 DVDD.n2034 0.0126434
R11718 DVDD.n7952 DVDD.n2054 0.0126434
R11719 DVDD.n2053 DVDD.n2033 0.0126434
R11720 DVDD.n7953 DVDD.n2056 0.0126434
R11721 DVDD.n2055 DVDD.n2032 0.0126434
R11722 DVDD.n7957 DVDD.n7955 0.0126434
R11723 DVDD.n7956 DVDD.n2031 0.0126434
R11724 DVDD.n7959 DVDD.n2027 0.0126434
R11725 DVDD.n2052 DVDD.n2051 0.0126434
R11726 DVDD.n7952 DVDD.n2034 0.0126434
R11727 DVDD.n2054 DVDD.n2053 0.0126434
R11728 DVDD.n7953 DVDD.n2033 0.0126434
R11729 DVDD.n2056 DVDD.n2055 0.0126434
R11730 DVDD.n7955 DVDD.n2032 0.0126434
R11731 DVDD.n7957 DVDD.n7956 0.0126434
R11732 DVDD.n2031 DVDD.n2027 0.0126434
R11733 DVDD.n6480 DVDD.n3402 0.0126434
R11734 DVDD.n6482 DVDD.n6471 0.0126434
R11735 DVDD.n6479 DVDD.n3401 0.0126434
R11736 DVDD.n6483 DVDD.n6472 0.0126434
R11737 DVDD.n6478 DVDD.n3400 0.0126434
R11738 DVDD.n6484 DVDD.n6473 0.0126434
R11739 DVDD.n6480 DVDD.n6470 0.0126434
R11740 DVDD.n6482 DVDD.n3402 0.0126434
R11741 DVDD.n6479 DVDD.n6471 0.0126434
R11742 DVDD.n6483 DVDD.n3401 0.0126434
R11743 DVDD.n6478 DVDD.n6472 0.0126434
R11744 DVDD.n6484 DVDD.n3400 0.0126434
R11745 DVDD.n3478 DVDD.n3476 0.0126434
R11746 DVDD.n3478 DVDD.n3477 0.0126434
R11747 DVDD.n3481 DVDD.n3479 0.0126434
R11748 DVDD.n3481 DVDD.n3480 0.0126434
R11749 DVDD.n6463 DVDD.n3482 0.0126434
R11750 DVDD.n6463 DVDD.n6462 0.0126434
R11751 DVDD.n3476 DVDD.n3471 0.0126434
R11752 DVDD.n3477 DVDD.n3470 0.0126434
R11753 DVDD.n3479 DVDD.n3470 0.0126434
R11754 DVDD.n3480 DVDD.n3469 0.0126434
R11755 DVDD.n3482 DVDD.n3469 0.0126434
R11756 DVDD.n6462 DVDD.n3419 0.0126434
R11757 DVDD.n3547 DVDD.n3535 0.0126434
R11758 DVDD.n3550 DVDD.n3532 0.0126434
R11759 DVDD.n3548 DVDD.n3536 0.0126434
R11760 DVDD.n3547 DVDD.n3533 0.0126434
R11761 DVDD.n3550 DVDD.n3535 0.0126434
R11762 DVDD.n3548 DVDD.n3532 0.0126434
R11763 DVDD.n3493 DVDD.n3492 0.0124104
R11764 DVDD.n6461 DVDD.n6460 0.0124104
R11765 DVDD.n6649 DVDD.n3358 0.0123701
R11766 DVDD.n6492 DVDD.n2076 0.0123701
R11767 DVDD.n3288 DVDD.n3226 0.0123701
R11768 DVDD.n3255 DVDD.n2127 0.0123701
R11769 DVDD.n6705 DVDD.n3180 0.0123701
R11770 DVDD.n3146 DVDD.n2173 0.0123701
R11771 DVDD.n2709 DVDD.n2671 0.0123701
R11772 DVDD.n2649 DVDD.n2637 0.0123701
R11773 DVDD.n7716 DVDD.n1887 0.0121929
R11774 DVDD.n7722 DVDD.n1669 0.0121929
R11775 DVDD.n2345 DVDD.n1605 0.0121929
R11776 DVDD.n2350 DVDD.n1550 0.0121929
R11777 DVDD.n3495 DVDD.n3494 0.0121222
R11778 DVDD.n5473 DVDD.n4465 0.0120157
R11779 DVDD.n5475 DVDD.n4464 0.0120157
R11780 DVDD.n5480 DVDD.n5478 0.0120157
R11781 DVDD.n5479 DVDD.n4463 0.0120157
R11782 DVDD.n713 DVDD.n584 0.0120157
R11783 DVDD.n8720 DVDD.n356 0.0120157
R11784 DVDD.n3734 DVDD.n3640 0.0120157
R11785 DVDD.n3834 DVDD.n3567 0.0120157
R11786 DVDD.n6523 DVDD.n2082 0.0120157
R11787 DVDD.n1885 DVDD.n1884 0.0120157
R11788 DVDD.n8985 DVDD.n556 0.0120157
R11789 DVDD.n4074 DVDD.n372 0.0120157
R11790 DVDD.n4202 DVDD.n4155 0.0120157
R11791 DVDD.n6034 DVDD.n3964 0.0120157
R11792 DVDD.n3286 DVDD.n2121 0.0120157
R11793 DVDD.n8291 DVDD.n1679 0.0120157
R11794 DVDD.n5022 DVDD.n4861 0.0120157
R11795 DVDD.n370 DVDD.n369 0.0120157
R11796 DVDD.n9546 DVDD.n9545 0.0120157
R11797 DVDD.n5801 DVDD.n4311 0.0120157
R11798 DVDD.n3176 DVDD.n2179 0.0120157
R11799 DVDD.n1871 DVDD.n1601 0.0120157
R11800 DVDD.n5129 DVDD.n4578 0.0120157
R11801 DVDD.n401 DVDD.n375 0.0120157
R11802 DVDD.n6778 DVDD.n2956 0.0120157
R11803 DVDD.n2861 DVDD.n2826 0.0120157
R11804 DVDD.n2707 DVDD.n2646 0.0120157
R11805 DVDD.n8357 DVDD.n1562 0.0120157
R11806 DVDD.n5419 DVDD.n5417 0.0119575
R11807 DVDD.n5418 DVDD.n4483 0.0119575
R11808 DVDD.n5422 DVDD.n5420 0.0119575
R11809 DVDD.n5652 DVDD.n5651 0.0119575
R11810 DVDD.n5643 DVDD.n4462 0.0119575
R11811 DVDD.n5654 DVDD.n5653 0.0119575
R11812 DVDD.n5642 DVDD.n4461 0.0119575
R11813 DVDD.n5656 DVDD.n5655 0.0119575
R11814 DVDD.n5641 DVDD.n4460 0.0119575
R11815 DVDD.n5551 DVDD.n5503 0.0119575
R11816 DVDD.n5555 DVDD.n5553 0.0119575
R11817 DVDD.n5554 DVDD.n5502 0.0119575
R11818 DVDD.n5558 DVDD.n5556 0.0119575
R11819 DVDD.n5557 DVDD.n5501 0.0119575
R11820 DVDD.n5561 DVDD.n5559 0.0119575
R11821 DVDD.n2544 DVDD.n2527 0.0119575
R11822 DVDD.n7018 DVDD.n2547 0.0119575
R11823 DVDD.n2546 DVDD.n2526 0.0119575
R11824 DVDD.n7019 DVDD.n2549 0.0119575
R11825 DVDD.n2548 DVDD.n2525 0.0119575
R11826 DVDD.n7023 DVDD.n7021 0.0119575
R11827 DVDD.n7022 DVDD.n2524 0.0119575
R11828 DVDD.n7025 DVDD.n2520 0.0119575
R11829 DVDD.n7535 DVDD.n7524 0.0119575
R11830 DVDD.n7521 DVDD.n2519 0.0119575
R11831 DVDD.n7536 DVDD.n7525 0.0119575
R11832 DVDD.n7520 DVDD.n2518 0.0119575
R11833 DVDD.n7537 DVDD.n7526 0.0119575
R11834 DVDD.n7519 DVDD.n2517 0.0119575
R11835 DVDD.n7538 DVDD.n7527 0.0119575
R11836 DVDD.n7518 DVDD.n2516 0.0119575
R11837 DVDD.n7539 DVDD.n7528 0.0119575
R11838 DVDD.n7517 DVDD.n2515 0.0119575
R11839 DVDD.n7540 DVDD.n7529 0.0119575
R11840 DVDD.n7516 DVDD.n2514 0.0119575
R11841 DVDD.n7541 DVDD.n7530 0.0119575
R11842 DVDD.n7515 DVDD.n2513 0.0119575
R11843 DVDD.n7542 DVDD.n7531 0.0119575
R11844 DVDD.n7514 DVDD.n2512 0.0119575
R11845 DVDD.n7543 DVDD.n7532 0.0119575
R11846 DVDD.n7513 DVDD.n2511 0.0119575
R11847 DVDD.n7544 DVDD.n7533 0.0119575
R11848 DVDD.n7512 DVDD.n2510 0.0119575
R11849 DVDD.n7547 DVDD.n7546 0.0119575
R11850 DVDD.n7511 DVDD.n2509 0.0119575
R11851 DVDD.n7549 DVDD.n7027 0.0119575
R11852 DVDD.n7045 DVDD.n7028 0.0119575
R11853 DVDD.n7044 DVDD.n7042 0.0119575
R11854 DVDD.n7212 DVDD.n7047 0.0119575
R11855 DVDD.n7046 DVDD.n7041 0.0119575
R11856 DVDD.n7213 DVDD.n7049 0.0119575
R11857 DVDD.n7048 DVDD.n7040 0.0119575
R11858 DVDD.n7214 DVDD.n7051 0.0119575
R11859 DVDD.n7050 DVDD.n7039 0.0119575
R11860 DVDD.n7215 DVDD.n7053 0.0119575
R11861 DVDD.n7052 DVDD.n7038 0.0119575
R11862 DVDD.n7216 DVDD.n7055 0.0119575
R11863 DVDD.n7054 DVDD.n7037 0.0119575
R11864 DVDD.n7217 DVDD.n7057 0.0119575
R11865 DVDD.n7056 DVDD.n7036 0.0119575
R11866 DVDD.n7218 DVDD.n7059 0.0119575
R11867 DVDD.n7058 DVDD.n7035 0.0119575
R11868 DVDD.n7219 DVDD.n7061 0.0119575
R11869 DVDD.n7060 DVDD.n7034 0.0119575
R11870 DVDD.n7220 DVDD.n7063 0.0119575
R11871 DVDD.n7062 DVDD.n7033 0.0119575
R11872 DVDD.n7221 DVDD.n7065 0.0119575
R11873 DVDD.n7064 DVDD.n7032 0.0119575
R11874 DVDD.n7507 DVDD.n7066 0.0119575
R11875 DVDD.n7075 DVDD.n7067 0.0119575
R11876 DVDD.n7078 DVDD.n7077 0.0119575
R11877 DVDD.n7089 DVDD.n7074 0.0119575
R11878 DVDD.n7080 DVDD.n7079 0.0119575
R11879 DVDD.n7088 DVDD.n7073 0.0119575
R11880 DVDD.n7082 DVDD.n7081 0.0119575
R11881 DVDD.n7087 DVDD.n7072 0.0119575
R11882 DVDD.n7084 DVDD.n7083 0.0119575
R11883 DVDD.n7086 DVDD.n7071 0.0119575
R11884 DVDD.n7504 DVDD.n7085 0.0119575
R11885 DVDD.n5417 DVDD.n5377 0.0119575
R11886 DVDD.n5419 DVDD.n5418 0.0119575
R11887 DVDD.n5420 DVDD.n4483 0.0119575
R11888 DVDD.n5651 DVDD.n4463 0.0119575
R11889 DVDD.n5652 DVDD.n4462 0.0119575
R11890 DVDD.n5653 DVDD.n5643 0.0119575
R11891 DVDD.n5654 DVDD.n4461 0.0119575
R11892 DVDD.n5655 DVDD.n5642 0.0119575
R11893 DVDD.n5656 DVDD.n4460 0.0119575
R11894 DVDD.n5552 DVDD.n5551 0.0119575
R11895 DVDD.n5553 DVDD.n5503 0.0119575
R11896 DVDD.n5555 DVDD.n5554 0.0119575
R11897 DVDD.n5556 DVDD.n5502 0.0119575
R11898 DVDD.n5558 DVDD.n5557 0.0119575
R11899 DVDD.n5559 DVDD.n5501 0.0119575
R11900 DVDD.n2545 DVDD.n2544 0.0119575
R11901 DVDD.n7018 DVDD.n2527 0.0119575
R11902 DVDD.n2547 DVDD.n2546 0.0119575
R11903 DVDD.n7019 DVDD.n2526 0.0119575
R11904 DVDD.n2549 DVDD.n2548 0.0119575
R11905 DVDD.n7021 DVDD.n2525 0.0119575
R11906 DVDD.n7023 DVDD.n7022 0.0119575
R11907 DVDD.n2524 DVDD.n2520 0.0119575
R11908 DVDD.n7535 DVDD.n7026 0.0119575
R11909 DVDD.n7524 DVDD.n2519 0.0119575
R11910 DVDD.n7536 DVDD.n7521 0.0119575
R11911 DVDD.n7525 DVDD.n2518 0.0119575
R11912 DVDD.n7537 DVDD.n7520 0.0119575
R11913 DVDD.n7526 DVDD.n2517 0.0119575
R11914 DVDD.n7538 DVDD.n7519 0.0119575
R11915 DVDD.n7527 DVDD.n2516 0.0119575
R11916 DVDD.n7539 DVDD.n7518 0.0119575
R11917 DVDD.n7528 DVDD.n2515 0.0119575
R11918 DVDD.n7540 DVDD.n7517 0.0119575
R11919 DVDD.n7529 DVDD.n2514 0.0119575
R11920 DVDD.n7541 DVDD.n7516 0.0119575
R11921 DVDD.n7530 DVDD.n2513 0.0119575
R11922 DVDD.n7542 DVDD.n7515 0.0119575
R11923 DVDD.n7531 DVDD.n2512 0.0119575
R11924 DVDD.n7543 DVDD.n7514 0.0119575
R11925 DVDD.n7532 DVDD.n2511 0.0119575
R11926 DVDD.n7544 DVDD.n7513 0.0119575
R11927 DVDD.n7533 DVDD.n2510 0.0119575
R11928 DVDD.n7546 DVDD.n7512 0.0119575
R11929 DVDD.n7547 DVDD.n2509 0.0119575
R11930 DVDD.n7511 DVDD.n7027 0.0119575
R11931 DVDD.n7509 DVDD.n7028 0.0119575
R11932 DVDD.n7045 DVDD.n7044 0.0119575
R11933 DVDD.n7212 DVDD.n7042 0.0119575
R11934 DVDD.n7047 DVDD.n7046 0.0119575
R11935 DVDD.n7213 DVDD.n7041 0.0119575
R11936 DVDD.n7049 DVDD.n7048 0.0119575
R11937 DVDD.n7214 DVDD.n7040 0.0119575
R11938 DVDD.n7051 DVDD.n7050 0.0119575
R11939 DVDD.n7215 DVDD.n7039 0.0119575
R11940 DVDD.n7053 DVDD.n7052 0.0119575
R11941 DVDD.n7216 DVDD.n7038 0.0119575
R11942 DVDD.n7055 DVDD.n7054 0.0119575
R11943 DVDD.n7217 DVDD.n7037 0.0119575
R11944 DVDD.n7057 DVDD.n7056 0.0119575
R11945 DVDD.n7218 DVDD.n7036 0.0119575
R11946 DVDD.n7059 DVDD.n7058 0.0119575
R11947 DVDD.n7219 DVDD.n7035 0.0119575
R11948 DVDD.n7061 DVDD.n7060 0.0119575
R11949 DVDD.n7220 DVDD.n7034 0.0119575
R11950 DVDD.n7063 DVDD.n7062 0.0119575
R11951 DVDD.n7221 DVDD.n7033 0.0119575
R11952 DVDD.n7065 DVDD.n7064 0.0119575
R11953 DVDD.n7066 DVDD.n7032 0.0119575
R11954 DVDD.n3806 DVDD.n3805 0.0119575
R11955 DVDD.n3573 DVDD.n3572 0.0119575
R11956 DVDD.n3571 DVDD.n3556 0.0119575
R11957 DVDD.n6314 DVDD.n3875 0.0119575
R11958 DVDD.n6314 DVDD.n6313 0.0119575
R11959 DVDD.n6311 DVDD.n6310 0.0119575
R11960 DVDD.n6310 DVDD.n3877 0.0119575
R11961 DVDD.n6303 DVDD.n6241 0.0119575
R11962 DVDD.n6303 DVDD.n6302 0.0119575
R11963 DVDD.n3361 DVDD.n3338 0.0119575
R11964 DVDD.n6645 DVDD.n3350 0.0119575
R11965 DVDD.n3360 DVDD.n3337 0.0119575
R11966 DVDD.n6646 DVDD.n3351 0.0119575
R11967 DVDD.n3359 DVDD.n3336 0.0119575
R11968 DVDD.n6647 DVDD.n3352 0.0119575
R11969 DVDD.n2104 DVDD.n2100 0.0119575
R11970 DVDD.n2102 DVDD.n2091 0.0119575
R11971 DVDD.n2103 DVDD.n2099 0.0119575
R11972 DVDD.n7888 DVDD.n2092 0.0119575
R11973 DVDD.n7887 DVDD.n2098 0.0119575
R11974 DVDD.n7889 DVDD.n2093 0.0119575
R11975 DVDD.n7891 DVDD.n2095 0.0119575
R11976 DVDD.n7892 DVDD.n2094 0.0119575
R11977 DVDD.n1974 DVDD.n1955 0.0119575
R11978 DVDD.n1987 DVDD.n1971 0.0119575
R11979 DVDD.n1975 DVDD.n1956 0.0119575
R11980 DVDD.n1986 DVDD.n1970 0.0119575
R11981 DVDD.n1976 DVDD.n1957 0.0119575
R11982 DVDD.n1969 DVDD.n1952 0.0119575
R11983 DVDD.n8050 DVDD.n1978 0.0119575
R11984 DVDD.n1968 DVDD.n1951 0.0119575
R11985 DVDD.n8051 DVDD.n1979 0.0119575
R11986 DVDD.n1967 DVDD.n1950 0.0119575
R11987 DVDD.n1980 DVDD.n1959 0.0119575
R11988 DVDD.n1985 DVDD.n1965 0.0119575
R11989 DVDD.n1981 DVDD.n1960 0.0119575
R11990 DVDD.n1984 DVDD.n1964 0.0119575
R11991 DVDD.n1982 DVDD.n1961 0.0119575
R11992 DVDD.n1963 DVDD.n1948 0.0119575
R11993 DVDD.n8055 DVDD.n1962 0.0119575
R11994 DVDD.n8109 DVDD.n1900 0.0119575
R11995 DVDD.n1898 DVDD.n1863 0.0119575
R11996 DVDD.n8110 DVDD.n1901 0.0119575
R11997 DVDD.n1897 DVDD.n1862 0.0119575
R11998 DVDD.n8111 DVDD.n1886 0.0119575
R11999 DVDD.n8112 DVDD.n1902 0.0119575
R12000 DVDD.n1896 DVDD.n1859 0.0119575
R12001 DVDD.n8113 DVDD.n1903 0.0119575
R12002 DVDD.n1895 DVDD.n1858 0.0119575
R12003 DVDD.n8114 DVDD.n1904 0.0119575
R12004 DVDD.n1894 DVDD.n1855 0.0119575
R12005 DVDD.n8117 DVDD.n8116 0.0119575
R12006 DVDD.n1893 DVDD.n1854 0.0119575
R12007 DVDD.n8119 DVDD.n1890 0.0119575
R12008 DVDD.n1756 DVDD.n1745 0.0119575
R12009 DVDD.n1759 DVDD.n1748 0.0119575
R12010 DVDD.n1755 DVDD.n1744 0.0119575
R12011 DVDD.n1760 DVDD.n1749 0.0119575
R12012 DVDD.n1754 DVDD.n1743 0.0119575
R12013 DVDD.n1761 DVDD.n1750 0.0119575
R12014 DVDD.n1753 DVDD.n1742 0.0119575
R12015 DVDD.n8251 DVDD.n1751 0.0119575
R12016 DVDD.n1752 DVDD.n1741 0.0119575
R12017 DVDD.n1762 DVDD.n1317 0.0119575
R12018 DVDD.n1321 DVDD.n1318 0.0119575
R12019 DVDD.n8630 DVDD.n1316 0.0119575
R12020 DVDD.n8629 DVDD.n8628 0.0119575
R12021 DVDD.n3807 DVDD.n3806 0.0119575
R12022 DVDD.n3805 DVDD.n3573 0.0119575
R12023 DVDD.n3572 DVDD.n3571 0.0119575
R12024 DVDD.n3875 DVDD.n3874 0.0119575
R12025 DVDD.n6312 DVDD.n6311 0.0119575
R12026 DVDD.n6313 DVDD.n6312 0.0119575
R12027 DVDD.n6241 DVDD.n6240 0.0119575
R12028 DVDD.n6240 DVDD.n3877 0.0119575
R12029 DVDD.n6302 DVDD.n6301 0.0119575
R12030 DVDD.n3361 DVDD.n3349 0.0119575
R12031 DVDD.n6645 DVDD.n3338 0.0119575
R12032 DVDD.n3360 DVDD.n3350 0.0119575
R12033 DVDD.n6646 DVDD.n3337 0.0119575
R12034 DVDD.n3359 DVDD.n3351 0.0119575
R12035 DVDD.n6647 DVDD.n3336 0.0119575
R12036 DVDD.n2104 DVDD.n2090 0.0119575
R12037 DVDD.n2100 DVDD.n2091 0.0119575
R12038 DVDD.n2103 DVDD.n2102 0.0119575
R12039 DVDD.n2099 DVDD.n2092 0.0119575
R12040 DVDD.n7888 DVDD.n7887 0.0119575
R12041 DVDD.n2098 DVDD.n2093 0.0119575
R12042 DVDD.n7889 DVDD.n2095 0.0119575
R12043 DVDD.n7892 DVDD.n7891 0.0119575
R12044 DVDD.n1972 DVDD.n1955 0.0119575
R12045 DVDD.n1987 DVDD.n1974 0.0119575
R12046 DVDD.n1971 DVDD.n1956 0.0119575
R12047 DVDD.n1986 DVDD.n1975 0.0119575
R12048 DVDD.n1970 DVDD.n1957 0.0119575
R12049 DVDD.n1977 DVDD.n1952 0.0119575
R12050 DVDD.n8050 DVDD.n1969 0.0119575
R12051 DVDD.n1978 DVDD.n1951 0.0119575
R12052 DVDD.n8051 DVDD.n1968 0.0119575
R12053 DVDD.n1979 DVDD.n1950 0.0119575
R12054 DVDD.n1966 DVDD.n1959 0.0119575
R12055 DVDD.n1985 DVDD.n1980 0.0119575
R12056 DVDD.n1965 DVDD.n1960 0.0119575
R12057 DVDD.n1984 DVDD.n1981 0.0119575
R12058 DVDD.n1964 DVDD.n1961 0.0119575
R12059 DVDD.n8053 DVDD.n1948 0.0119575
R12060 DVDD.n1963 DVDD.n1962 0.0119575
R12061 DVDD.n8109 DVDD.n1864 0.0119575
R12062 DVDD.n1900 DVDD.n1863 0.0119575
R12063 DVDD.n8110 DVDD.n1898 0.0119575
R12064 DVDD.n1901 DVDD.n1862 0.0119575
R12065 DVDD.n8111 DVDD.n1897 0.0119575
R12066 DVDD.n8112 DVDD.n1860 0.0119575
R12067 DVDD.n1902 DVDD.n1859 0.0119575
R12068 DVDD.n8113 DVDD.n1896 0.0119575
R12069 DVDD.n1903 DVDD.n1858 0.0119575
R12070 DVDD.n8114 DVDD.n1856 0.0119575
R12071 DVDD.n1904 DVDD.n1855 0.0119575
R12072 DVDD.n8116 DVDD.n1894 0.0119575
R12073 DVDD.n8117 DVDD.n1854 0.0119575
R12074 DVDD.n1893 DVDD.n1890 0.0119575
R12075 DVDD.n4280 DVDD.n3947 0.0119575
R12076 DVDD.n4281 DVDD.n3969 0.0119575
R12077 DVDD.n4284 DVDD.n3948 0.0119575
R12078 DVDD.n6001 DVDD.n6000 0.0119575
R12079 DVDD.n5932 DVDD.n5925 0.0119575
R12080 DVDD.n5999 DVDD.n5998 0.0119575
R12081 DVDD.n5933 DVDD.n5926 0.0119575
R12082 DVDD.n5997 DVDD.n5996 0.0119575
R12083 DVDD.n5993 DVDD.n5927 0.0119575
R12084 DVDD.n3299 DVDD.n3221 0.0119575
R12085 DVDD.n3301 DVDD.n3300 0.0119575
R12086 DVDD.n3302 DVDD.n3222 0.0119575
R12087 DVDD.n3304 DVDD.n3303 0.0119575
R12088 DVDD.n3305 DVDD.n3223 0.0119575
R12089 DVDD.n3306 DVDD.n3230 0.0119575
R12090 DVDD.n2145 DVDD.n2129 0.0119575
R12091 DVDD.n7841 DVDD.n2135 0.0119575
R12092 DVDD.n2146 DVDD.n2130 0.0119575
R12093 DVDD.n7840 DVDD.n2134 0.0119575
R12094 DVDD.n2147 DVDD.n2131 0.0119575
R12095 DVDD.n7839 DVDD.n2133 0.0119575
R12096 DVDD.n2148 DVDD.n2132 0.0119575
R12097 DVDD.n7852 DVDD.n2144 0.0119575
R12098 DVDD.n2299 DVDD.n2280 0.0119575
R12099 DVDD.n2331 DVDD.n2330 0.0119575
R12100 DVDD.n2300 DVDD.n2281 0.0119575
R12101 DVDD.n2329 DVDD.n2328 0.0119575
R12102 DVDD.n2298 DVDD.n2279 0.0119575
R12103 DVDD.n2327 DVDD.n2288 0.0119575
R12104 DVDD.n2326 DVDD.n2302 0.0119575
R12105 DVDD.n2325 DVDD.n2287 0.0119575
R12106 DVDD.n2324 DVDD.n2303 0.0119575
R12107 DVDD.n2297 DVDD.n2278 0.0119575
R12108 DVDD.n2304 DVDD.n2282 0.0119575
R12109 DVDD.n2322 DVDD.n2321 0.0119575
R12110 DVDD.n2305 DVDD.n2283 0.0119575
R12111 DVDD.n2320 DVDD.n2319 0.0119575
R12112 DVDD.n2296 DVDD.n2277 0.0119575
R12113 DVDD.n2318 DVDD.n2286 0.0119575
R12114 DVDD.n2317 DVDD.n2284 0.0119575
R12115 DVDD.n1690 DVDD.n1666 0.0119575
R12116 DVDD.n1689 DVDD.n1686 0.0119575
R12117 DVDD.n1692 DVDD.n1667 0.0119575
R12118 DVDD.n1691 DVDD.n1685 0.0119575
R12119 DVDD.n1693 DVDD.n1668 0.0119575
R12120 DVDD.n1695 DVDD.n1670 0.0119575
R12121 DVDD.n1694 DVDD.n1683 0.0119575
R12122 DVDD.n1697 DVDD.n1671 0.0119575
R12123 DVDD.n1696 DVDD.n1663 0.0119575
R12124 DVDD.n1699 DVDD.n1674 0.0119575
R12125 DVDD.n1698 DVDD.n1681 0.0119575
R12126 DVDD.n1701 DVDD.n1675 0.0119575
R12127 DVDD.n1700 DVDD.n1680 0.0119575
R12128 DVDD.n8289 DVDD.n1676 0.0119575
R12129 DVDD.n1711 DVDD.n1702 0.0119575
R12130 DVDD.n1714 DVDD.n1713 0.0119575
R12131 DVDD.n1722 DVDD.n1710 0.0119575
R12132 DVDD.n1716 DVDD.n1715 0.0119575
R12133 DVDD.n1721 DVDD.n1709 0.0119575
R12134 DVDD.n1718 DVDD.n1717 0.0119575
R12135 DVDD.n1720 DVDD.n1708 0.0119575
R12136 DVDD.n8286 DVDD.n1719 0.0119575
R12137 DVDD.n8285 DVDD.n1707 0.0119575
R12138 DVDD.n1706 DVDD.n1309 0.0119575
R12139 DVDD.n1313 DVDD.n1310 0.0119575
R12140 DVDD.n8635 DVDD.n1308 0.0119575
R12141 DVDD.n8634 DVDD.n1314 0.0119575
R12142 DVDD.n1687 DVDD.n1666 0.0119575
R12143 DVDD.n1690 DVDD.n1689 0.0119575
R12144 DVDD.n1686 DVDD.n1667 0.0119575
R12145 DVDD.n1692 DVDD.n1691 0.0119575
R12146 DVDD.n1685 DVDD.n1668 0.0119575
R12147 DVDD.n1684 DVDD.n1670 0.0119575
R12148 DVDD.n1695 DVDD.n1694 0.0119575
R12149 DVDD.n1683 DVDD.n1671 0.0119575
R12150 DVDD.n1697 DVDD.n1696 0.0119575
R12151 DVDD.n1682 DVDD.n1674 0.0119575
R12152 DVDD.n1699 DVDD.n1698 0.0119575
R12153 DVDD.n1681 DVDD.n1675 0.0119575
R12154 DVDD.n1701 DVDD.n1700 0.0119575
R12155 DVDD.n1680 DVDD.n1676 0.0119575
R12156 DVDD.n2318 DVDD.n2317 0.0119575
R12157 DVDD.n2306 DVDD.n2286 0.0119575
R12158 DVDD.n2320 DVDD.n2277 0.0119575
R12159 DVDD.n2319 DVDD.n2305 0.0119575
R12160 DVDD.n2322 DVDD.n2283 0.0119575
R12161 DVDD.n2321 DVDD.n2304 0.0119575
R12162 DVDD.n2323 DVDD.n2282 0.0119575
R12163 DVDD.n2303 DVDD.n2278 0.0119575
R12164 DVDD.n2325 DVDD.n2324 0.0119575
R12165 DVDD.n2302 DVDD.n2287 0.0119575
R12166 DVDD.n2327 DVDD.n2326 0.0119575
R12167 DVDD.n2301 DVDD.n2288 0.0119575
R12168 DVDD.n2329 DVDD.n2279 0.0119575
R12169 DVDD.n2328 DVDD.n2300 0.0119575
R12170 DVDD.n2331 DVDD.n2281 0.0119575
R12171 DVDD.n2330 DVDD.n2299 0.0119575
R12172 DVDD.n7746 DVDD.n2280 0.0119575
R12173 DVDD.n2144 DVDD.n2132 0.0119575
R12174 DVDD.n2148 DVDD.n2133 0.0119575
R12175 DVDD.n7839 DVDD.n2131 0.0119575
R12176 DVDD.n2147 DVDD.n2134 0.0119575
R12177 DVDD.n7840 DVDD.n2130 0.0119575
R12178 DVDD.n2146 DVDD.n2135 0.0119575
R12179 DVDD.n7841 DVDD.n2129 0.0119575
R12180 DVDD.n2145 DVDD.n2136 0.0119575
R12181 DVDD.n3306 DVDD.n3305 0.0119575
R12182 DVDD.n3303 DVDD.n3223 0.0119575
R12183 DVDD.n3304 DVDD.n3302 0.0119575
R12184 DVDD.n3300 DVDD.n3222 0.0119575
R12185 DVDD.n3301 DVDD.n3299 0.0119575
R12186 DVDD.n3298 DVDD.n3221 0.0119575
R12187 DVDD.n5997 DVDD.n5927 0.0119575
R12188 DVDD.n5996 DVDD.n5933 0.0119575
R12189 DVDD.n5999 DVDD.n5926 0.0119575
R12190 DVDD.n5998 DVDD.n5932 0.0119575
R12191 DVDD.n6001 DVDD.n5925 0.0119575
R12192 DVDD.n6000 DVDD.n5924 0.0119575
R12193 DVDD.n4284 DVDD.n3969 0.0119575
R12194 DVDD.n4281 DVDD.n3947 0.0119575
R12195 DVDD.n6154 DVDD.n4280 0.0119575
R12196 DVDD.n6108 DVDD.n6107 0.0119575
R12197 DVDD.n6109 DVDD.n4316 0.0119575
R12198 DVDD.n6110 DVDD.n4377 0.0119575
R12199 DVDD.n5888 DVDD.n5825 0.0119575
R12200 DVDD.n5895 DVDD.n5762 0.0119575
R12201 DVDD.n5889 DVDD.n5826 0.0119575
R12202 DVDD.n5894 DVDD.n5761 0.0119575
R12203 DVDD.n5890 DVDD.n5827 0.0119575
R12204 DVDD.n5893 DVDD.n5760 0.0119575
R12205 DVDD.n3183 DVDD.n3103 0.0119575
R12206 DVDD.n6701 DVDD.n3115 0.0119575
R12207 DVDD.n3182 DVDD.n3102 0.0119575
R12208 DVDD.n6702 DVDD.n3116 0.0119575
R12209 DVDD.n3181 DVDD.n3101 0.0119575
R12210 DVDD.n6703 DVDD.n3117 0.0119575
R12211 DVDD.n7797 DVDD.n2196 0.0119575
R12212 DVDD.n7795 DVDD.n2188 0.0119575
R12213 DVDD.n7796 DVDD.n2195 0.0119575
R12214 DVDD.n7801 DVDD.n2189 0.0119575
R12215 DVDD.n7800 DVDD.n2194 0.0119575
R12216 DVDD.n7802 DVDD.n2190 0.0119575
R12217 DVDD.n7804 DVDD.n2192 0.0119575
R12218 DVDD.n7805 DVDD.n2191 0.0119575
R12219 DVDD.n2237 DVDD.n2218 0.0119575
R12220 DVDD.n2250 DVDD.n2234 0.0119575
R12221 DVDD.n2238 DVDD.n2219 0.0119575
R12222 DVDD.n2249 DVDD.n2233 0.0119575
R12223 DVDD.n2239 DVDD.n2220 0.0119575
R12224 DVDD.n2232 DVDD.n2215 0.0119575
R12225 DVDD.n7774 DVDD.n2241 0.0119575
R12226 DVDD.n2231 DVDD.n2214 0.0119575
R12227 DVDD.n7775 DVDD.n2242 0.0119575
R12228 DVDD.n2230 DVDD.n2213 0.0119575
R12229 DVDD.n2243 DVDD.n2222 0.0119575
R12230 DVDD.n2248 DVDD.n2228 0.0119575
R12231 DVDD.n2244 DVDD.n2223 0.0119575
R12232 DVDD.n2247 DVDD.n2227 0.0119575
R12233 DVDD.n2245 DVDD.n2224 0.0119575
R12234 DVDD.n2226 DVDD.n2211 0.0119575
R12235 DVDD.n7779 DVDD.n2225 0.0119575
R12236 DVDD.n1621 DVDD.n1602 0.0119575
R12237 DVDD.n1618 DVDD.n1597 0.0119575
R12238 DVDD.n1622 DVDD.n1603 0.0119575
R12239 DVDD.n1617 DVDD.n1596 0.0119575
R12240 DVDD.n1623 DVDD.n1604 0.0119575
R12241 DVDD.n1624 DVDD.n1606 0.0119575
R12242 DVDD.n1616 DVDD.n1593 0.0119575
R12243 DVDD.n1625 DVDD.n1607 0.0119575
R12244 DVDD.n1615 DVDD.n1592 0.0119575
R12245 DVDD.n1626 DVDD.n1610 0.0119575
R12246 DVDD.n1614 DVDD.n1589 0.0119575
R12247 DVDD.n1627 DVDD.n1611 0.0119575
R12248 DVDD.n1613 DVDD.n1588 0.0119575
R12249 DVDD.n8322 DVDD.n1612 0.0119575
R12250 DVDD.n7368 DVDD.n7338 0.0119575
R12251 DVDD.n7422 DVDD.n7370 0.0119575
R12252 DVDD.n7367 DVDD.n7337 0.0119575
R12253 DVDD.n7423 DVDD.n7371 0.0119575
R12254 DVDD.n7366 DVDD.n7336 0.0119575
R12255 DVDD.n7424 DVDD.n7372 0.0119575
R12256 DVDD.n7365 DVDD.n7335 0.0119575
R12257 DVDD.n7427 DVDD.n7426 0.0119575
R12258 DVDD.n7364 DVDD.n7334 0.0119575
R12259 DVDD.n7429 DVDD.n7340 0.0119575
R12260 DVDD.n7342 DVDD.n7341 0.0119575
R12261 DVDD.n7361 DVDD.n7345 0.0119575
R12262 DVDD.n7360 DVDD.n7359 0.0119575
R12263 DVDD.n6108 DVDD.n4376 0.0119575
R12264 DVDD.n6107 DVDD.n4316 0.0119575
R12265 DVDD.n6110 DVDD.n6109 0.0119575
R12266 DVDD.n5888 DVDD.n5763 0.0119575
R12267 DVDD.n5895 DVDD.n5825 0.0119575
R12268 DVDD.n5889 DVDD.n5762 0.0119575
R12269 DVDD.n5894 DVDD.n5826 0.0119575
R12270 DVDD.n5890 DVDD.n5761 0.0119575
R12271 DVDD.n5893 DVDD.n5827 0.0119575
R12272 DVDD.n3183 DVDD.n3114 0.0119575
R12273 DVDD.n6701 DVDD.n3103 0.0119575
R12274 DVDD.n3182 DVDD.n3115 0.0119575
R12275 DVDD.n6702 DVDD.n3102 0.0119575
R12276 DVDD.n3181 DVDD.n3116 0.0119575
R12277 DVDD.n6703 DVDD.n3101 0.0119575
R12278 DVDD.n7797 DVDD.n2187 0.0119575
R12279 DVDD.n2196 DVDD.n2188 0.0119575
R12280 DVDD.n7796 DVDD.n7795 0.0119575
R12281 DVDD.n2195 DVDD.n2189 0.0119575
R12282 DVDD.n7801 DVDD.n7800 0.0119575
R12283 DVDD.n2194 DVDD.n2190 0.0119575
R12284 DVDD.n7802 DVDD.n2192 0.0119575
R12285 DVDD.n7805 DVDD.n7804 0.0119575
R12286 DVDD.n2235 DVDD.n2218 0.0119575
R12287 DVDD.n2250 DVDD.n2237 0.0119575
R12288 DVDD.n2234 DVDD.n2219 0.0119575
R12289 DVDD.n2249 DVDD.n2238 0.0119575
R12290 DVDD.n2233 DVDD.n2220 0.0119575
R12291 DVDD.n2240 DVDD.n2215 0.0119575
R12292 DVDD.n7774 DVDD.n2232 0.0119575
R12293 DVDD.n2241 DVDD.n2214 0.0119575
R12294 DVDD.n7775 DVDD.n2231 0.0119575
R12295 DVDD.n2242 DVDD.n2213 0.0119575
R12296 DVDD.n2229 DVDD.n2222 0.0119575
R12297 DVDD.n2248 DVDD.n2243 0.0119575
R12298 DVDD.n2228 DVDD.n2223 0.0119575
R12299 DVDD.n2247 DVDD.n2244 0.0119575
R12300 DVDD.n2227 DVDD.n2224 0.0119575
R12301 DVDD.n7777 DVDD.n2211 0.0119575
R12302 DVDD.n2226 DVDD.n2225 0.0119575
R12303 DVDD.n1621 DVDD.n1598 0.0119575
R12304 DVDD.n1618 DVDD.n1602 0.0119575
R12305 DVDD.n1622 DVDD.n1597 0.0119575
R12306 DVDD.n1617 DVDD.n1603 0.0119575
R12307 DVDD.n1623 DVDD.n1596 0.0119575
R12308 DVDD.n1624 DVDD.n1594 0.0119575
R12309 DVDD.n1616 DVDD.n1606 0.0119575
R12310 DVDD.n1625 DVDD.n1593 0.0119575
R12311 DVDD.n1615 DVDD.n1607 0.0119575
R12312 DVDD.n1626 DVDD.n1590 0.0119575
R12313 DVDD.n1614 DVDD.n1610 0.0119575
R12314 DVDD.n1627 DVDD.n1589 0.0119575
R12315 DVDD.n1613 DVDD.n1611 0.0119575
R12316 DVDD.n1612 DVDD.n1588 0.0119575
R12317 DVDD.n7361 DVDD.n7360 0.0119575
R12318 DVDD.n8635 DVDD.n8634 0.0119575
R12319 DVDD.n8630 DVDD.n8629 0.0119575
R12320 DVDD.n7345 DVDD.n7342 0.0119575
R12321 DVDD.n1313 DVDD.n1308 0.0119575
R12322 DVDD.n1321 DVDD.n1316 0.0119575
R12323 DVDD.n7363 DVDD.n7341 0.0119575
R12324 DVDD.n8637 DVDD.n1310 0.0119575
R12325 DVDD.n8632 DVDD.n1318 0.0119575
R12326 DVDD.n6854 DVDD.n2809 0.0119575
R12327 DVDD.n2878 DVDD.n2876 0.0119575
R12328 DVDD.n2877 DVDD.n2803 0.0119575
R12329 DVDD.n6877 DVDD.n6874 0.0119575
R12330 DVDD.n6876 DVDD.n6875 0.0119575
R12331 DVDD.n6888 DVDD.n2784 0.0119575
R12332 DVDD.n6890 DVDD.n6889 0.0119575
R12333 DVDD.n6893 DVDD.n6891 0.0119575
R12334 DVDD.n6892 DVDD.n2742 0.0119575
R12335 DVDD.n2732 DVDD.n2730 0.0119575
R12336 DVDD.n2731 DVDD.n2666 0.0119575
R12337 DVDD.n2729 DVDD.n2727 0.0119575
R12338 DVDD.n2728 DVDD.n2667 0.0119575
R12339 DVDD.n2726 DVDD.n2724 0.0119575
R12340 DVDD.n2725 DVDD.n2655 0.0119575
R12341 DVDD.n6977 DVDD.n6936 0.0119575
R12342 DVDD.n6981 DVDD.n2641 0.0119575
R12343 DVDD.n6980 DVDD.n6937 0.0119575
R12344 DVDD.n6941 DVDD.n2640 0.0119575
R12345 DVDD.n6978 DVDD.n6938 0.0119575
R12346 DVDD.n6940 DVDD.n2639 0.0119575
R12347 DVDD.n6983 DVDD.n6933 0.0119575
R12348 DVDD.n6984 DVDD.n2355 0.0119575
R12349 DVDD.n2379 DVDD.n2373 0.0119575
R12350 DVDD.n2403 DVDD.n2402 0.0119575
R12351 DVDD.n2455 DVDD.n2380 0.0119575
R12352 DVDD.n2401 DVDD.n2400 0.0119575
R12353 DVDD.n2454 DVDD.n2378 0.0119575
R12354 DVDD.n7659 DVDD.n2399 0.0119575
R12355 DVDD.n2398 DVDD.n2382 0.0119575
R12356 DVDD.n7658 DVDD.n2397 0.0119575
R12357 DVDD.n2396 DVDD.n2383 0.0119575
R12358 DVDD.n2453 DVDD.n2377 0.0119575
R12359 DVDD.n2456 DVDD.n2384 0.0119575
R12360 DVDD.n2394 DVDD.n2393 0.0119575
R12361 DVDD.n2457 DVDD.n2385 0.0119575
R12362 DVDD.n2392 DVDD.n2391 0.0119575
R12363 DVDD.n2452 DVDD.n2376 0.0119575
R12364 DVDD.n7657 DVDD.n2390 0.0119575
R12365 DVDD.n2389 DVDD.n2387 0.0119575
R12366 DVDD.n8349 DVDD.n1546 0.0119575
R12367 DVDD.n1545 DVDD.n1542 0.0119575
R12368 DVDD.n8350 DVDD.n1548 0.0119575
R12369 DVDD.n1547 DVDD.n1541 0.0119575
R12370 DVDD.n8351 DVDD.n1549 0.0119575
R12371 DVDD.n8352 DVDD.n1552 0.0119575
R12372 DVDD.n1551 DVDD.n1538 0.0119575
R12373 DVDD.n8353 DVDD.n1554 0.0119575
R12374 DVDD.n1553 DVDD.n1537 0.0119575
R12375 DVDD.n8354 DVDD.n1558 0.0119575
R12376 DVDD.n1557 DVDD.n1534 0.0119575
R12377 DVDD.n8355 DVDD.n1560 0.0119575
R12378 DVDD.n1559 DVDD.n1533 0.0119575
R12379 DVDD.n8359 DVDD.n1528 0.0119575
R12380 DVDD.n8361 DVDD.n1519 0.0119575
R12381 DVDD.n8362 DVDD.n1522 0.0119575
R12382 DVDD.n1521 DVDD.n1518 0.0119575
R12383 DVDD.n8363 DVDD.n1524 0.0119575
R12384 DVDD.n1523 DVDD.n1517 0.0119575
R12385 DVDD.n8364 DVDD.n1526 0.0119575
R12386 DVDD.n1525 DVDD.n1516 0.0119575
R12387 DVDD.n8368 DVDD.n8366 0.0119575
R12388 DVDD.n8367 DVDD.n1515 0.0119575
R12389 DVDD.n8370 DVDD.n1511 0.0119575
R12390 DVDD.n8371 DVDD.n1503 0.0119575
R12391 DVDD.n1510 DVDD.n1509 0.0119575
R12392 DVDD.n8377 DVDD.n1505 0.0119575
R12393 DVDD.n1509 DVDD.n1505 0.0119575
R12394 DVDD.n8372 DVDD.n1503 0.0119575
R12395 DVDD.n8372 DVDD.n1510 0.0119575
R12396 DVDD.n8349 DVDD.n1543 0.0119575
R12397 DVDD.n1546 DVDD.n1545 0.0119575
R12398 DVDD.n8350 DVDD.n1542 0.0119575
R12399 DVDD.n1548 DVDD.n1547 0.0119575
R12400 DVDD.n8351 DVDD.n1541 0.0119575
R12401 DVDD.n8352 DVDD.n1539 0.0119575
R12402 DVDD.n1552 DVDD.n1551 0.0119575
R12403 DVDD.n8353 DVDD.n1538 0.0119575
R12404 DVDD.n1554 DVDD.n1553 0.0119575
R12405 DVDD.n8354 DVDD.n1535 0.0119575
R12406 DVDD.n1558 DVDD.n1557 0.0119575
R12407 DVDD.n8355 DVDD.n1534 0.0119575
R12408 DVDD.n1560 DVDD.n1559 0.0119575
R12409 DVDD.n1533 DVDD.n1528 0.0119575
R12410 DVDD.n2390 DVDD.n2389 0.0119575
R12411 DVDD.n7657 DVDD.n2386 0.0119575
R12412 DVDD.n2452 DVDD.n2392 0.0119575
R12413 DVDD.n2391 DVDD.n2385 0.0119575
R12414 DVDD.n2457 DVDD.n2394 0.0119575
R12415 DVDD.n2393 DVDD.n2384 0.0119575
R12416 DVDD.n2456 DVDD.n2395 0.0119575
R12417 DVDD.n2453 DVDD.n2383 0.0119575
R12418 DVDD.n2397 DVDD.n2396 0.0119575
R12419 DVDD.n7658 DVDD.n2382 0.0119575
R12420 DVDD.n2399 DVDD.n2398 0.0119575
R12421 DVDD.n7659 DVDD.n2381 0.0119575
R12422 DVDD.n2454 DVDD.n2401 0.0119575
R12423 DVDD.n2400 DVDD.n2380 0.0119575
R12424 DVDD.n2455 DVDD.n2403 0.0119575
R12425 DVDD.n2402 DVDD.n2379 0.0119575
R12426 DVDD.n7680 DVDD.n2373 0.0119575
R12427 DVDD.n6984 DVDD.n6983 0.0119575
R12428 DVDD.n6940 DVDD.n6933 0.0119575
R12429 DVDD.n6938 DVDD.n2639 0.0119575
R12430 DVDD.n6978 DVDD.n6941 0.0119575
R12431 DVDD.n6937 DVDD.n2640 0.0119575
R12432 DVDD.n6981 DVDD.n6980 0.0119575
R12433 DVDD.n6936 DVDD.n2641 0.0119575
R12434 DVDD.n6977 DVDD.n2642 0.0119575
R12435 DVDD.n2726 DVDD.n2725 0.0119575
R12436 DVDD.n2724 DVDD.n2667 0.0119575
R12437 DVDD.n2729 DVDD.n2728 0.0119575
R12438 DVDD.n2727 DVDD.n2666 0.0119575
R12439 DVDD.n2732 DVDD.n2731 0.0119575
R12440 DVDD.n2730 DVDD.n2665 0.0119575
R12441 DVDD.n6893 DVDD.n6892 0.0119575
R12442 DVDD.n6891 DVDD.n6890 0.0119575
R12443 DVDD.n6889 DVDD.n6888 0.0119575
R12444 DVDD.n6875 DVDD.n2784 0.0119575
R12445 DVDD.n6877 DVDD.n6876 0.0119575
R12446 DVDD.n6874 DVDD.n6873 0.0119575
R12447 DVDD.n2878 DVDD.n2877 0.0119575
R12448 DVDD.n2876 DVDD.n2809 0.0119575
R12449 DVDD.n6855 DVDD.n6854 0.0119575
R12450 DVDD.n8360 DVDD.n1519 0.0119575
R12451 DVDD.n8362 DVDD.n8361 0.0119575
R12452 DVDD.n1522 DVDD.n1521 0.0119575
R12453 DVDD.n8363 DVDD.n1518 0.0119575
R12454 DVDD.n1524 DVDD.n1523 0.0119575
R12455 DVDD.n8364 DVDD.n1517 0.0119575
R12456 DVDD.n1526 DVDD.n1525 0.0119575
R12457 DVDD.n8366 DVDD.n1516 0.0119575
R12458 DVDD.n8368 DVDD.n8367 0.0119575
R12459 DVDD.n1515 DVDD.n1511 0.0119575
R12460 DVDD.n8288 DVDD.n1702 0.0119575
R12461 DVDD.n1713 DVDD.n1711 0.0119575
R12462 DVDD.n1722 DVDD.n1714 0.0119575
R12463 DVDD.n1715 DVDD.n1710 0.0119575
R12464 DVDD.n1721 DVDD.n1716 0.0119575
R12465 DVDD.n1717 DVDD.n1709 0.0119575
R12466 DVDD.n1720 DVDD.n1718 0.0119575
R12467 DVDD.n1719 DVDD.n1708 0.0119575
R12468 DVDD.n8286 DVDD.n8285 0.0119575
R12469 DVDD.n1707 DVDD.n1706 0.0119575
R12470 DVDD.n7506 DVDD.n7067 0.0119575
R12471 DVDD.n7077 DVDD.n7075 0.0119575
R12472 DVDD.n7089 DVDD.n7078 0.0119575
R12473 DVDD.n7079 DVDD.n7074 0.0119575
R12474 DVDD.n7088 DVDD.n7080 0.0119575
R12475 DVDD.n7081 DVDD.n7073 0.0119575
R12476 DVDD.n7087 DVDD.n7082 0.0119575
R12477 DVDD.n7083 DVDD.n7072 0.0119575
R12478 DVDD.n7086 DVDD.n7084 0.0119575
R12479 DVDD.n7085 DVDD.n7071 0.0119575
R12480 DVDD.n7338 DVDD.n1620 0.0119575
R12481 DVDD.n7422 DVDD.n7368 0.0119575
R12482 DVDD.n7370 DVDD.n7337 0.0119575
R12483 DVDD.n7423 DVDD.n7367 0.0119575
R12484 DVDD.n7371 DVDD.n7336 0.0119575
R12485 DVDD.n7424 DVDD.n7366 0.0119575
R12486 DVDD.n7372 DVDD.n7335 0.0119575
R12487 DVDD.n7426 DVDD.n7365 0.0119575
R12488 DVDD.n7427 DVDD.n7334 0.0119575
R12489 DVDD.n7364 DVDD.n7340 0.0119575
R12490 DVDD.n1756 DVDD.n1747 0.0119575
R12491 DVDD.n1759 DVDD.n1745 0.0119575
R12492 DVDD.n1755 DVDD.n1748 0.0119575
R12493 DVDD.n1760 DVDD.n1744 0.0119575
R12494 DVDD.n1754 DVDD.n1749 0.0119575
R12495 DVDD.n1761 DVDD.n1743 0.0119575
R12496 DVDD.n1753 DVDD.n1750 0.0119575
R12497 DVDD.n1751 DVDD.n1742 0.0119575
R12498 DVDD.n8251 DVDD.n1752 0.0119575
R12499 DVDD.n1762 DVDD.n1741 0.0119575
R12500 DVDD.n618 DVDD.n616 0.0119575
R12501 DVDD.n621 DVDD.n620 0.0119575
R12502 DVDD.n632 DVDD.n615 0.0119575
R12503 DVDD.n623 DVDD.n622 0.0119575
R12504 DVDD.n631 DVDD.n614 0.0119575
R12505 DVDD.n625 DVDD.n624 0.0119575
R12506 DVDD.n630 DVDD.n613 0.0119575
R12507 DVDD.n627 DVDD.n626 0.0119575
R12508 DVDD.n629 DVDD.n612 0.0119575
R12509 DVDD.n8911 DVDD.n628 0.0119575
R12510 DVDD.n31 DVDD.n29 0.0119575
R12511 DVDD.n35 DVDD.n33 0.0119575
R12512 DVDD.n34 DVDD.n28 0.0119575
R12513 DVDD.n38 DVDD.n36 0.0119575
R12514 DVDD.n37 DVDD.n27 0.0119575
R12515 DVDD.n41 DVDD.n39 0.0119575
R12516 DVDD.n40 DVDD.n26 0.0119575
R12517 DVDD.n44 DVDD.n42 0.0119575
R12518 DVDD.n43 DVDD.n25 0.0119575
R12519 DVDD.n9673 DVDD.n45 0.0119575
R12520 DVDD.n1072 DVDD.n1055 0.0119575
R12521 DVDD.n1071 DVDD.n1069 0.0119575
R12522 DVDD.n6410 DVDD.n1074 0.0119575
R12523 DVDD.n1073 DVDD.n1068 0.0119575
R12524 DVDD.n6411 DVDD.n1076 0.0119575
R12525 DVDD.n1075 DVDD.n1067 0.0119575
R12526 DVDD.n6412 DVDD.n1078 0.0119575
R12527 DVDD.n1077 DVDD.n1066 0.0119575
R12528 DVDD.n6413 DVDD.n1080 0.0119575
R12529 DVDD.n1079 DVDD.n1065 0.0119575
R12530 DVDD.n6414 DVDD.n1082 0.0119575
R12531 DVDD.n1081 DVDD.n1064 0.0119575
R12532 DVDD.n6415 DVDD.n1084 0.0119575
R12533 DVDD.n1083 DVDD.n1063 0.0119575
R12534 DVDD.n6416 DVDD.n1086 0.0119575
R12535 DVDD.n1085 DVDD.n1062 0.0119575
R12536 DVDD.n6417 DVDD.n1088 0.0119575
R12537 DVDD.n1087 DVDD.n1061 0.0119575
R12538 DVDD.n6418 DVDD.n1090 0.0119575
R12539 DVDD.n1089 DVDD.n1060 0.0119575
R12540 DVDD.n6419 DVDD.n1092 0.0119575
R12541 DVDD.n1091 DVDD.n1059 0.0119575
R12542 DVDD.n8665 DVDD.n1093 0.0119575
R12543 DVDD.n1101 DVDD.n1094 0.0119575
R12544 DVDD.n1104 DVDD.n1103 0.0119575
R12545 DVDD.n1115 DVDD.n1100 0.0119575
R12546 DVDD.n1106 DVDD.n1105 0.0119575
R12547 DVDD.n1114 DVDD.n1099 0.0119575
R12548 DVDD.n1108 DVDD.n1107 0.0119575
R12549 DVDD.n1113 DVDD.n1098 0.0119575
R12550 DVDD.n1110 DVDD.n1109 0.0119575
R12551 DVDD.n1112 DVDD.n1097 0.0119575
R12552 DVDD.n8662 DVDD.n1111 0.0119575
R12553 DVDD.n1134 DVDD.n1117 0.0119575
R12554 DVDD.n1133 DVDD.n1131 0.0119575
R12555 DVDD.n6616 DVDD.n1136 0.0119575
R12556 DVDD.n1135 DVDD.n1130 0.0119575
R12557 DVDD.n6617 DVDD.n1138 0.0119575
R12558 DVDD.n1137 DVDD.n1129 0.0119575
R12559 DVDD.n6618 DVDD.n1140 0.0119575
R12560 DVDD.n1139 DVDD.n1128 0.0119575
R12561 DVDD.n6619 DVDD.n1142 0.0119575
R12562 DVDD.n1141 DVDD.n1127 0.0119575
R12563 DVDD.n6620 DVDD.n1144 0.0119575
R12564 DVDD.n1143 DVDD.n1126 0.0119575
R12565 DVDD.n6621 DVDD.n1146 0.0119575
R12566 DVDD.n1145 DVDD.n1125 0.0119575
R12567 DVDD.n6622 DVDD.n1148 0.0119575
R12568 DVDD.n1147 DVDD.n1124 0.0119575
R12569 DVDD.n6623 DVDD.n1150 0.0119575
R12570 DVDD.n1149 DVDD.n1123 0.0119575
R12571 DVDD.n6624 DVDD.n1152 0.0119575
R12572 DVDD.n1151 DVDD.n1122 0.0119575
R12573 DVDD.n6625 DVDD.n1154 0.0119575
R12574 DVDD.n1153 DVDD.n1121 0.0119575
R12575 DVDD.n8659 DVDD.n1155 0.0119575
R12576 DVDD.n1173 DVDD.n1156 0.0119575
R12577 DVDD.n1172 DVDD.n1170 0.0119575
R12578 DVDD.n7916 DVDD.n1175 0.0119575
R12579 DVDD.n1174 DVDD.n1169 0.0119575
R12580 DVDD.n7917 DVDD.n1177 0.0119575
R12581 DVDD.n1176 DVDD.n1168 0.0119575
R12582 DVDD.n7918 DVDD.n1179 0.0119575
R12583 DVDD.n1178 DVDD.n1167 0.0119575
R12584 DVDD.n7919 DVDD.n1181 0.0119575
R12585 DVDD.n1180 DVDD.n1166 0.0119575
R12586 DVDD.n7920 DVDD.n1183 0.0119575
R12587 DVDD.n1182 DVDD.n1165 0.0119575
R12588 DVDD.n7921 DVDD.n1185 0.0119575
R12589 DVDD.n1184 DVDD.n1164 0.0119575
R12590 DVDD.n7922 DVDD.n1187 0.0119575
R12591 DVDD.n1186 DVDD.n1163 0.0119575
R12592 DVDD.n7923 DVDD.n1189 0.0119575
R12593 DVDD.n1188 DVDD.n1162 0.0119575
R12594 DVDD.n7924 DVDD.n1191 0.0119575
R12595 DVDD.n1190 DVDD.n1161 0.0119575
R12596 DVDD.n7925 DVDD.n1193 0.0119575
R12597 DVDD.n1192 DVDD.n1160 0.0119575
R12598 DVDD.n8656 DVDD.n1194 0.0119575
R12599 DVDD.n1212 DVDD.n1195 0.0119575
R12600 DVDD.n1211 DVDD.n1209 0.0119575
R12601 DVDD.n8021 DVDD.n1214 0.0119575
R12602 DVDD.n1213 DVDD.n1208 0.0119575
R12603 DVDD.n8022 DVDD.n1216 0.0119575
R12604 DVDD.n1215 DVDD.n1207 0.0119575
R12605 DVDD.n8023 DVDD.n1218 0.0119575
R12606 DVDD.n1217 DVDD.n1206 0.0119575
R12607 DVDD.n8024 DVDD.n1220 0.0119575
R12608 DVDD.n1219 DVDD.n1205 0.0119575
R12609 DVDD.n8025 DVDD.n1222 0.0119575
R12610 DVDD.n1221 DVDD.n1204 0.0119575
R12611 DVDD.n8026 DVDD.n1224 0.0119575
R12612 DVDD.n1223 DVDD.n1203 0.0119575
R12613 DVDD.n8027 DVDD.n1226 0.0119575
R12614 DVDD.n1225 DVDD.n1202 0.0119575
R12615 DVDD.n8028 DVDD.n1228 0.0119575
R12616 DVDD.n1227 DVDD.n1201 0.0119575
R12617 DVDD.n8029 DVDD.n1230 0.0119575
R12618 DVDD.n1229 DVDD.n1200 0.0119575
R12619 DVDD.n8030 DVDD.n1232 0.0119575
R12620 DVDD.n1231 DVDD.n1199 0.0119575
R12621 DVDD.n8653 DVDD.n1233 0.0119575
R12622 DVDD.n1251 DVDD.n1234 0.0119575
R12623 DVDD.n1250 DVDD.n1248 0.0119575
R12624 DVDD.n8143 DVDD.n1253 0.0119575
R12625 DVDD.n1252 DVDD.n1247 0.0119575
R12626 DVDD.n8144 DVDD.n1255 0.0119575
R12627 DVDD.n1254 DVDD.n1246 0.0119575
R12628 DVDD.n8145 DVDD.n1257 0.0119575
R12629 DVDD.n1256 DVDD.n1245 0.0119575
R12630 DVDD.n8146 DVDD.n1259 0.0119575
R12631 DVDD.n1258 DVDD.n1244 0.0119575
R12632 DVDD.n8147 DVDD.n1261 0.0119575
R12633 DVDD.n1260 DVDD.n1243 0.0119575
R12634 DVDD.n8148 DVDD.n1263 0.0119575
R12635 DVDD.n1262 DVDD.n1242 0.0119575
R12636 DVDD.n8149 DVDD.n1267 0.0119575
R12637 DVDD.n1266 DVDD.n1239 0.0119575
R12638 DVDD.n8150 DVDD.n1269 0.0119575
R12639 DVDD.n1268 DVDD.n1238 0.0119575
R12640 DVDD.n8650 DVDD.n1270 0.0119575
R12641 DVDD.n1279 DVDD.n1271 0.0119575
R12642 DVDD.n1282 DVDD.n1281 0.0119575
R12643 DVDD.n1293 DVDD.n1278 0.0119575
R12644 DVDD.n1284 DVDD.n1283 0.0119575
R12645 DVDD.n1292 DVDD.n1277 0.0119575
R12646 DVDD.n1286 DVDD.n1285 0.0119575
R12647 DVDD.n1291 DVDD.n1276 0.0119575
R12648 DVDD.n1288 DVDD.n1287 0.0119575
R12649 DVDD.n1290 DVDD.n1275 0.0119575
R12650 DVDD.n8647 DVDD.n1289 0.0119575
R12651 DVDD.n8643 DVDD.n1302 0.0119575
R12652 DVDD.n8667 DVDD.n1055 0.0119575
R12653 DVDD.n1072 DVDD.n1071 0.0119575
R12654 DVDD.n6410 DVDD.n1069 0.0119575
R12655 DVDD.n1074 DVDD.n1073 0.0119575
R12656 DVDD.n6411 DVDD.n1068 0.0119575
R12657 DVDD.n1076 DVDD.n1075 0.0119575
R12658 DVDD.n6412 DVDD.n1067 0.0119575
R12659 DVDD.n1078 DVDD.n1077 0.0119575
R12660 DVDD.n6413 DVDD.n1066 0.0119575
R12661 DVDD.n1080 DVDD.n1079 0.0119575
R12662 DVDD.n6414 DVDD.n1065 0.0119575
R12663 DVDD.n1082 DVDD.n1081 0.0119575
R12664 DVDD.n6415 DVDD.n1064 0.0119575
R12665 DVDD.n1084 DVDD.n1083 0.0119575
R12666 DVDD.n6416 DVDD.n1063 0.0119575
R12667 DVDD.n1086 DVDD.n1085 0.0119575
R12668 DVDD.n6417 DVDD.n1062 0.0119575
R12669 DVDD.n1088 DVDD.n1087 0.0119575
R12670 DVDD.n6418 DVDD.n1061 0.0119575
R12671 DVDD.n1090 DVDD.n1089 0.0119575
R12672 DVDD.n6419 DVDD.n1060 0.0119575
R12673 DVDD.n1092 DVDD.n1091 0.0119575
R12674 DVDD.n1093 DVDD.n1059 0.0119575
R12675 DVDD.n8664 DVDD.n1094 0.0119575
R12676 DVDD.n1103 DVDD.n1101 0.0119575
R12677 DVDD.n1115 DVDD.n1104 0.0119575
R12678 DVDD.n1105 DVDD.n1100 0.0119575
R12679 DVDD.n1114 DVDD.n1106 0.0119575
R12680 DVDD.n1107 DVDD.n1099 0.0119575
R12681 DVDD.n1113 DVDD.n1108 0.0119575
R12682 DVDD.n1109 DVDD.n1098 0.0119575
R12683 DVDD.n1112 DVDD.n1110 0.0119575
R12684 DVDD.n1111 DVDD.n1097 0.0119575
R12685 DVDD.n8661 DVDD.n1117 0.0119575
R12686 DVDD.n1134 DVDD.n1133 0.0119575
R12687 DVDD.n6616 DVDD.n1131 0.0119575
R12688 DVDD.n1136 DVDD.n1135 0.0119575
R12689 DVDD.n6617 DVDD.n1130 0.0119575
R12690 DVDD.n1138 DVDD.n1137 0.0119575
R12691 DVDD.n6618 DVDD.n1129 0.0119575
R12692 DVDD.n1140 DVDD.n1139 0.0119575
R12693 DVDD.n6619 DVDD.n1128 0.0119575
R12694 DVDD.n1142 DVDD.n1141 0.0119575
R12695 DVDD.n6620 DVDD.n1127 0.0119575
R12696 DVDD.n1144 DVDD.n1143 0.0119575
R12697 DVDD.n6621 DVDD.n1126 0.0119575
R12698 DVDD.n1146 DVDD.n1145 0.0119575
R12699 DVDD.n6622 DVDD.n1125 0.0119575
R12700 DVDD.n1148 DVDD.n1147 0.0119575
R12701 DVDD.n6623 DVDD.n1124 0.0119575
R12702 DVDD.n1150 DVDD.n1149 0.0119575
R12703 DVDD.n6624 DVDD.n1123 0.0119575
R12704 DVDD.n1152 DVDD.n1151 0.0119575
R12705 DVDD.n6625 DVDD.n1122 0.0119575
R12706 DVDD.n1154 DVDD.n1153 0.0119575
R12707 DVDD.n1155 DVDD.n1121 0.0119575
R12708 DVDD.n8658 DVDD.n1156 0.0119575
R12709 DVDD.n1173 DVDD.n1172 0.0119575
R12710 DVDD.n7916 DVDD.n1170 0.0119575
R12711 DVDD.n1175 DVDD.n1174 0.0119575
R12712 DVDD.n7917 DVDD.n1169 0.0119575
R12713 DVDD.n1177 DVDD.n1176 0.0119575
R12714 DVDD.n7918 DVDD.n1168 0.0119575
R12715 DVDD.n1179 DVDD.n1178 0.0119575
R12716 DVDD.n7919 DVDD.n1167 0.0119575
R12717 DVDD.n1181 DVDD.n1180 0.0119575
R12718 DVDD.n7920 DVDD.n1166 0.0119575
R12719 DVDD.n1183 DVDD.n1182 0.0119575
R12720 DVDD.n7921 DVDD.n1165 0.0119575
R12721 DVDD.n1185 DVDD.n1184 0.0119575
R12722 DVDD.n7922 DVDD.n1164 0.0119575
R12723 DVDD.n1187 DVDD.n1186 0.0119575
R12724 DVDD.n7923 DVDD.n1163 0.0119575
R12725 DVDD.n1189 DVDD.n1188 0.0119575
R12726 DVDD.n7924 DVDD.n1162 0.0119575
R12727 DVDD.n1191 DVDD.n1190 0.0119575
R12728 DVDD.n7925 DVDD.n1161 0.0119575
R12729 DVDD.n1193 DVDD.n1192 0.0119575
R12730 DVDD.n1194 DVDD.n1160 0.0119575
R12731 DVDD.n8655 DVDD.n1195 0.0119575
R12732 DVDD.n1212 DVDD.n1211 0.0119575
R12733 DVDD.n8021 DVDD.n1209 0.0119575
R12734 DVDD.n1214 DVDD.n1213 0.0119575
R12735 DVDD.n8022 DVDD.n1208 0.0119575
R12736 DVDD.n1216 DVDD.n1215 0.0119575
R12737 DVDD.n8023 DVDD.n1207 0.0119575
R12738 DVDD.n1218 DVDD.n1217 0.0119575
R12739 DVDD.n8024 DVDD.n1206 0.0119575
R12740 DVDD.n1220 DVDD.n1219 0.0119575
R12741 DVDD.n8025 DVDD.n1205 0.0119575
R12742 DVDD.n1222 DVDD.n1221 0.0119575
R12743 DVDD.n8026 DVDD.n1204 0.0119575
R12744 DVDD.n1224 DVDD.n1223 0.0119575
R12745 DVDD.n8027 DVDD.n1203 0.0119575
R12746 DVDD.n1226 DVDD.n1225 0.0119575
R12747 DVDD.n8028 DVDD.n1202 0.0119575
R12748 DVDD.n1228 DVDD.n1227 0.0119575
R12749 DVDD.n8029 DVDD.n1201 0.0119575
R12750 DVDD.n1230 DVDD.n1229 0.0119575
R12751 DVDD.n8030 DVDD.n1200 0.0119575
R12752 DVDD.n1232 DVDD.n1231 0.0119575
R12753 DVDD.n1233 DVDD.n1199 0.0119575
R12754 DVDD.n8652 DVDD.n1234 0.0119575
R12755 DVDD.n1251 DVDD.n1250 0.0119575
R12756 DVDD.n8143 DVDD.n1248 0.0119575
R12757 DVDD.n1253 DVDD.n1252 0.0119575
R12758 DVDD.n8144 DVDD.n1247 0.0119575
R12759 DVDD.n1255 DVDD.n1254 0.0119575
R12760 DVDD.n8145 DVDD.n1246 0.0119575
R12761 DVDD.n1257 DVDD.n1256 0.0119575
R12762 DVDD.n8146 DVDD.n1245 0.0119575
R12763 DVDD.n1259 DVDD.n1258 0.0119575
R12764 DVDD.n8147 DVDD.n1244 0.0119575
R12765 DVDD.n1261 DVDD.n1260 0.0119575
R12766 DVDD.n8148 DVDD.n1243 0.0119575
R12767 DVDD.n1263 DVDD.n1262 0.0119575
R12768 DVDD.n8149 DVDD.n1240 0.0119575
R12769 DVDD.n1267 DVDD.n1266 0.0119575
R12770 DVDD.n8150 DVDD.n1239 0.0119575
R12771 DVDD.n1269 DVDD.n1268 0.0119575
R12772 DVDD.n1270 DVDD.n1238 0.0119575
R12773 DVDD.n8649 DVDD.n1271 0.0119575
R12774 DVDD.n1281 DVDD.n1279 0.0119575
R12775 DVDD.n1293 DVDD.n1282 0.0119575
R12776 DVDD.n1283 DVDD.n1278 0.0119575
R12777 DVDD.n1292 DVDD.n1284 0.0119575
R12778 DVDD.n1285 DVDD.n1277 0.0119575
R12779 DVDD.n1291 DVDD.n1286 0.0119575
R12780 DVDD.n1287 DVDD.n1276 0.0119575
R12781 DVDD.n1290 DVDD.n1288 0.0119575
R12782 DVDD.n1289 DVDD.n1275 0.0119575
R12783 DVDD.n8644 DVDD.n8643 0.0119575
R12784 DVDD.n619 DVDD.n618 0.0119575
R12785 DVDD.n620 DVDD.n616 0.0119575
R12786 DVDD.n632 DVDD.n621 0.0119575
R12787 DVDD.n622 DVDD.n615 0.0119575
R12788 DVDD.n631 DVDD.n623 0.0119575
R12789 DVDD.n624 DVDD.n614 0.0119575
R12790 DVDD.n630 DVDD.n625 0.0119575
R12791 DVDD.n626 DVDD.n613 0.0119575
R12792 DVDD.n629 DVDD.n627 0.0119575
R12793 DVDD.n628 DVDD.n612 0.0119575
R12794 DVDD.n4605 DVDD.n4599 0.0119575
R12795 DVDD.n4729 DVDD.n4598 0.0119575
R12796 DVDD.n4736 DVDD.n4604 0.0119575
R12797 DVDD.n4730 DVDD.n4597 0.0119575
R12798 DVDD.n4735 DVDD.n4603 0.0119575
R12799 DVDD.n4731 DVDD.n4596 0.0119575
R12800 DVDD.n4734 DVDD.n4602 0.0119575
R12801 DVDD.n4732 DVDD.n4595 0.0119575
R12802 DVDD.n4733 DVDD.n4601 0.0119575
R12803 DVDD.n4818 DVDD.n4594 0.0119575
R12804 DVDD.n4747 DVDD.n4739 0.0119575
R12805 DVDD.n4780 DVDD.n4779 0.0119575
R12806 DVDD.n4778 DVDD.n4746 0.0119575
R12807 DVDD.n4782 DVDD.n4781 0.0119575
R12808 DVDD.n4777 DVDD.n4745 0.0119575
R12809 DVDD.n4784 DVDD.n4783 0.0119575
R12810 DVDD.n4776 DVDD.n4744 0.0119575
R12811 DVDD.n4786 DVDD.n4785 0.0119575
R12812 DVDD.n4775 DVDD.n4743 0.0119575
R12813 DVDD.n4774 DVDD.n432 0.0119575
R12814 DVDD.n2977 DVDD.n2960 0.0119575
R12815 DVDD.n2976 DVDD.n2974 0.0119575
R12816 DVDD.n5390 DVDD.n2979 0.0119575
R12817 DVDD.n2978 DVDD.n2973 0.0119575
R12818 DVDD.n5391 DVDD.n2981 0.0119575
R12819 DVDD.n2980 DVDD.n2972 0.0119575
R12820 DVDD.n5392 DVDD.n2983 0.0119575
R12821 DVDD.n2982 DVDD.n2971 0.0119575
R12822 DVDD.n5393 DVDD.n2985 0.0119575
R12823 DVDD.n2984 DVDD.n2970 0.0119575
R12824 DVDD.n5394 DVDD.n2987 0.0119575
R12825 DVDD.n2986 DVDD.n2969 0.0119575
R12826 DVDD.n5395 DVDD.n2989 0.0119575
R12827 DVDD.n2988 DVDD.n2968 0.0119575
R12828 DVDD.n5396 DVDD.n2991 0.0119575
R12829 DVDD.n2990 DVDD.n2967 0.0119575
R12830 DVDD.n5397 DVDD.n2993 0.0119575
R12831 DVDD.n2992 DVDD.n2966 0.0119575
R12832 DVDD.n5398 DVDD.n2995 0.0119575
R12833 DVDD.n2994 DVDD.n2965 0.0119575
R12834 DVDD.n5399 DVDD.n2997 0.0119575
R12835 DVDD.n2996 DVDD.n2964 0.0119575
R12836 DVDD.n6773 DVDD.n2998 0.0119575
R12837 DVDD.n3007 DVDD.n2999 0.0119575
R12838 DVDD.n3010 DVDD.n3009 0.0119575
R12839 DVDD.n3021 DVDD.n3006 0.0119575
R12840 DVDD.n3012 DVDD.n3011 0.0119575
R12841 DVDD.n3020 DVDD.n3005 0.0119575
R12842 DVDD.n3014 DVDD.n3013 0.0119575
R12843 DVDD.n3019 DVDD.n3004 0.0119575
R12844 DVDD.n3016 DVDD.n3015 0.0119575
R12845 DVDD.n3018 DVDD.n3003 0.0119575
R12846 DVDD.n6770 DVDD.n3017 0.0119575
R12847 DVDD.n3040 DVDD.n3023 0.0119575
R12848 DVDD.n3039 DVDD.n3037 0.0119575
R12849 DVDD.n6755 DVDD.n3042 0.0119575
R12850 DVDD.n3041 DVDD.n3036 0.0119575
R12851 DVDD.n6756 DVDD.n3044 0.0119575
R12852 DVDD.n3043 DVDD.n3035 0.0119575
R12853 DVDD.n6757 DVDD.n3046 0.0119575
R12854 DVDD.n3045 DVDD.n3034 0.0119575
R12855 DVDD.n6758 DVDD.n3048 0.0119575
R12856 DVDD.n3047 DVDD.n3033 0.0119575
R12857 DVDD.n6759 DVDD.n3050 0.0119575
R12858 DVDD.n3049 DVDD.n3032 0.0119575
R12859 DVDD.n6760 DVDD.n3052 0.0119575
R12860 DVDD.n3051 DVDD.n3031 0.0119575
R12861 DVDD.n6761 DVDD.n3054 0.0119575
R12862 DVDD.n3053 DVDD.n3030 0.0119575
R12863 DVDD.n6762 DVDD.n3056 0.0119575
R12864 DVDD.n3055 DVDD.n3029 0.0119575
R12865 DVDD.n6763 DVDD.n3058 0.0119575
R12866 DVDD.n3057 DVDD.n3028 0.0119575
R12867 DVDD.n6764 DVDD.n3060 0.0119575
R12868 DVDD.n3059 DVDD.n3027 0.0119575
R12869 DVDD.n6767 DVDD.n6766 0.0119575
R12870 DVDD.n2598 DVDD.n2574 0.0119575
R12871 DVDD.n2596 DVDD.n2571 0.0119575
R12872 DVDD.n2599 DVDD.n2575 0.0119575
R12873 DVDD.n2595 DVDD.n2570 0.0119575
R12874 DVDD.n2600 DVDD.n2576 0.0119575
R12875 DVDD.n2594 DVDD.n2569 0.0119575
R12876 DVDD.n2601 DVDD.n2577 0.0119575
R12877 DVDD.n2593 DVDD.n2568 0.0119575
R12878 DVDD.n2602 DVDD.n2578 0.0119575
R12879 DVDD.n2592 DVDD.n2567 0.0119575
R12880 DVDD.n2603 DVDD.n2579 0.0119575
R12881 DVDD.n2591 DVDD.n2566 0.0119575
R12882 DVDD.n2604 DVDD.n2580 0.0119575
R12883 DVDD.n2590 DVDD.n2565 0.0119575
R12884 DVDD.n2605 DVDD.n2581 0.0119575
R12885 DVDD.n2589 DVDD.n2564 0.0119575
R12886 DVDD.n2606 DVDD.n2582 0.0119575
R12887 DVDD.n2588 DVDD.n2563 0.0119575
R12888 DVDD.n2607 DVDD.n2583 0.0119575
R12889 DVDD.n2587 DVDD.n2562 0.0119575
R12890 DVDD.n2608 DVDD.n2584 0.0119575
R12891 DVDD.n2586 DVDD.n2561 0.0119575
R12892 DVDD.n7004 DVDD.n2585 0.0119575
R12893 DVDD.n7577 DVDD.n7566 0.0119575
R12894 DVDD.n2500 DVDD.n2485 0.0119575
R12895 DVDD.n7578 DVDD.n7567 0.0119575
R12896 DVDD.n2499 DVDD.n2484 0.0119575
R12897 DVDD.n7579 DVDD.n7568 0.0119575
R12898 DVDD.n2498 DVDD.n2483 0.0119575
R12899 DVDD.n7580 DVDD.n7569 0.0119575
R12900 DVDD.n2497 DVDD.n2482 0.0119575
R12901 DVDD.n7581 DVDD.n7570 0.0119575
R12902 DVDD.n2496 DVDD.n2481 0.0119575
R12903 DVDD.n7582 DVDD.n7571 0.0119575
R12904 DVDD.n2495 DVDD.n2480 0.0119575
R12905 DVDD.n7583 DVDD.n7572 0.0119575
R12906 DVDD.n2494 DVDD.n2479 0.0119575
R12907 DVDD.n7584 DVDD.n7573 0.0119575
R12908 DVDD.n2493 DVDD.n2478 0.0119575
R12909 DVDD.n7585 DVDD.n7574 0.0119575
R12910 DVDD.n2492 DVDD.n2477 0.0119575
R12911 DVDD.n7586 DVDD.n7575 0.0119575
R12912 DVDD.n2491 DVDD.n2476 0.0119575
R12913 DVDD.n7589 DVDD.n7588 0.0119575
R12914 DVDD.n2490 DVDD.n2475 0.0119575
R12915 DVDD.n7591 DVDD.n2487 0.0119575
R12916 DVDD.n7273 DVDD.n7122 0.0119575
R12917 DVDD.n7121 DVDD.n7119 0.0119575
R12918 DVDD.n7274 DVDD.n7124 0.0119575
R12919 DVDD.n7123 DVDD.n7118 0.0119575
R12920 DVDD.n7275 DVDD.n7126 0.0119575
R12921 DVDD.n7125 DVDD.n7117 0.0119575
R12922 DVDD.n7276 DVDD.n7128 0.0119575
R12923 DVDD.n7127 DVDD.n7116 0.0119575
R12924 DVDD.n7277 DVDD.n7130 0.0119575
R12925 DVDD.n7129 DVDD.n7115 0.0119575
R12926 DVDD.n7278 DVDD.n7132 0.0119575
R12927 DVDD.n7131 DVDD.n7114 0.0119575
R12928 DVDD.n7279 DVDD.n7134 0.0119575
R12929 DVDD.n7133 DVDD.n7113 0.0119575
R12930 DVDD.n7280 DVDD.n7204 0.0119575
R12931 DVDD.n7203 DVDD.n7110 0.0119575
R12932 DVDD.n7284 DVDD.n7282 0.0119575
R12933 DVDD.n7283 DVDD.n7109 0.0119575
R12934 DVDD.n7286 DVDD.n7105 0.0119575
R12935 DVDD.n7297 DVDD.n7103 0.0119575
R12936 DVDD.n7300 DVDD.n7288 0.0119575
R12937 DVDD.n7296 DVDD.n7102 0.0119575
R12938 DVDD.n7301 DVDD.n7289 0.0119575
R12939 DVDD.n7295 DVDD.n7101 0.0119575
R12940 DVDD.n7302 DVDD.n7290 0.0119575
R12941 DVDD.n7294 DVDD.n7100 0.0119575
R12942 DVDD.n7303 DVDD.n7291 0.0119575
R12943 DVDD.n7293 DVDD.n7099 0.0119575
R12944 DVDD.n7486 DVDD.n7292 0.0119575
R12945 DVDD.n8386 DVDD.n1498 0.0119575
R12946 DVDD.n4820 DVDD.n4599 0.0119575
R12947 DVDD.n4605 DVDD.n4598 0.0119575
R12948 DVDD.n4736 DVDD.n4729 0.0119575
R12949 DVDD.n4604 DVDD.n4597 0.0119575
R12950 DVDD.n4735 DVDD.n4730 0.0119575
R12951 DVDD.n4603 DVDD.n4596 0.0119575
R12952 DVDD.n4734 DVDD.n4731 0.0119575
R12953 DVDD.n4602 DVDD.n4595 0.0119575
R12954 DVDD.n4733 DVDD.n4732 0.0119575
R12955 DVDD.n4601 DVDD.n4594 0.0119575
R12956 DVDD.n6775 DVDD.n2960 0.0119575
R12957 DVDD.n2977 DVDD.n2976 0.0119575
R12958 DVDD.n5390 DVDD.n2974 0.0119575
R12959 DVDD.n2979 DVDD.n2978 0.0119575
R12960 DVDD.n5391 DVDD.n2973 0.0119575
R12961 DVDD.n2981 DVDD.n2980 0.0119575
R12962 DVDD.n5392 DVDD.n2972 0.0119575
R12963 DVDD.n2983 DVDD.n2982 0.0119575
R12964 DVDD.n5393 DVDD.n2971 0.0119575
R12965 DVDD.n2985 DVDD.n2984 0.0119575
R12966 DVDD.n5394 DVDD.n2970 0.0119575
R12967 DVDD.n2987 DVDD.n2986 0.0119575
R12968 DVDD.n5395 DVDD.n2969 0.0119575
R12969 DVDD.n2989 DVDD.n2988 0.0119575
R12970 DVDD.n5396 DVDD.n2968 0.0119575
R12971 DVDD.n2991 DVDD.n2990 0.0119575
R12972 DVDD.n5397 DVDD.n2967 0.0119575
R12973 DVDD.n2993 DVDD.n2992 0.0119575
R12974 DVDD.n5398 DVDD.n2966 0.0119575
R12975 DVDD.n2995 DVDD.n2994 0.0119575
R12976 DVDD.n5399 DVDD.n2965 0.0119575
R12977 DVDD.n2997 DVDD.n2996 0.0119575
R12978 DVDD.n2998 DVDD.n2964 0.0119575
R12979 DVDD.n6772 DVDD.n2999 0.0119575
R12980 DVDD.n3009 DVDD.n3007 0.0119575
R12981 DVDD.n3021 DVDD.n3010 0.0119575
R12982 DVDD.n3011 DVDD.n3006 0.0119575
R12983 DVDD.n3020 DVDD.n3012 0.0119575
R12984 DVDD.n3013 DVDD.n3005 0.0119575
R12985 DVDD.n3019 DVDD.n3014 0.0119575
R12986 DVDD.n3015 DVDD.n3004 0.0119575
R12987 DVDD.n3018 DVDD.n3016 0.0119575
R12988 DVDD.n3017 DVDD.n3003 0.0119575
R12989 DVDD.n6769 DVDD.n3023 0.0119575
R12990 DVDD.n3040 DVDD.n3039 0.0119575
R12991 DVDD.n6755 DVDD.n3037 0.0119575
R12992 DVDD.n3042 DVDD.n3041 0.0119575
R12993 DVDD.n6756 DVDD.n3036 0.0119575
R12994 DVDD.n3044 DVDD.n3043 0.0119575
R12995 DVDD.n6757 DVDD.n3035 0.0119575
R12996 DVDD.n3046 DVDD.n3045 0.0119575
R12997 DVDD.n6758 DVDD.n3034 0.0119575
R12998 DVDD.n3048 DVDD.n3047 0.0119575
R12999 DVDD.n6759 DVDD.n3033 0.0119575
R13000 DVDD.n3050 DVDD.n3049 0.0119575
R13001 DVDD.n6760 DVDD.n3032 0.0119575
R13002 DVDD.n3052 DVDD.n3051 0.0119575
R13003 DVDD.n6761 DVDD.n3031 0.0119575
R13004 DVDD.n3054 DVDD.n3053 0.0119575
R13005 DVDD.n6762 DVDD.n3030 0.0119575
R13006 DVDD.n3056 DVDD.n3055 0.0119575
R13007 DVDD.n6763 DVDD.n3029 0.0119575
R13008 DVDD.n3058 DVDD.n3057 0.0119575
R13009 DVDD.n6764 DVDD.n3028 0.0119575
R13010 DVDD.n3060 DVDD.n3059 0.0119575
R13011 DVDD.n6766 DVDD.n3027 0.0119575
R13012 DVDD.n2598 DVDD.n2572 0.0119575
R13013 DVDD.n2596 DVDD.n2574 0.0119575
R13014 DVDD.n2599 DVDD.n2571 0.0119575
R13015 DVDD.n2595 DVDD.n2575 0.0119575
R13016 DVDD.n2600 DVDD.n2570 0.0119575
R13017 DVDD.n2594 DVDD.n2576 0.0119575
R13018 DVDD.n2601 DVDD.n2569 0.0119575
R13019 DVDD.n2593 DVDD.n2577 0.0119575
R13020 DVDD.n2602 DVDD.n2568 0.0119575
R13021 DVDD.n2592 DVDD.n2578 0.0119575
R13022 DVDD.n2603 DVDD.n2567 0.0119575
R13023 DVDD.n2591 DVDD.n2579 0.0119575
R13024 DVDD.n2604 DVDD.n2566 0.0119575
R13025 DVDD.n2590 DVDD.n2580 0.0119575
R13026 DVDD.n2605 DVDD.n2565 0.0119575
R13027 DVDD.n2589 DVDD.n2581 0.0119575
R13028 DVDD.n2606 DVDD.n2564 0.0119575
R13029 DVDD.n2588 DVDD.n2582 0.0119575
R13030 DVDD.n2607 DVDD.n2563 0.0119575
R13031 DVDD.n2587 DVDD.n2583 0.0119575
R13032 DVDD.n2608 DVDD.n2562 0.0119575
R13033 DVDD.n2586 DVDD.n2584 0.0119575
R13034 DVDD.n2585 DVDD.n2561 0.0119575
R13035 DVDD.n7577 DVDD.n2486 0.0119575
R13036 DVDD.n7566 DVDD.n2485 0.0119575
R13037 DVDD.n7578 DVDD.n2500 0.0119575
R13038 DVDD.n7567 DVDD.n2484 0.0119575
R13039 DVDD.n7579 DVDD.n2499 0.0119575
R13040 DVDD.n7568 DVDD.n2483 0.0119575
R13041 DVDD.n7580 DVDD.n2498 0.0119575
R13042 DVDD.n7569 DVDD.n2482 0.0119575
R13043 DVDD.n7581 DVDD.n2497 0.0119575
R13044 DVDD.n7570 DVDD.n2481 0.0119575
R13045 DVDD.n7582 DVDD.n2496 0.0119575
R13046 DVDD.n7571 DVDD.n2480 0.0119575
R13047 DVDD.n7583 DVDD.n2495 0.0119575
R13048 DVDD.n7572 DVDD.n2479 0.0119575
R13049 DVDD.n7584 DVDD.n2494 0.0119575
R13050 DVDD.n7573 DVDD.n2478 0.0119575
R13051 DVDD.n7585 DVDD.n2493 0.0119575
R13052 DVDD.n7574 DVDD.n2477 0.0119575
R13053 DVDD.n7586 DVDD.n2492 0.0119575
R13054 DVDD.n7575 DVDD.n2476 0.0119575
R13055 DVDD.n7588 DVDD.n2491 0.0119575
R13056 DVDD.n7589 DVDD.n2475 0.0119575
R13057 DVDD.n2490 DVDD.n2487 0.0119575
R13058 DVDD.n7273 DVDD.n2488 0.0119575
R13059 DVDD.n7122 DVDD.n7121 0.0119575
R13060 DVDD.n7274 DVDD.n7119 0.0119575
R13061 DVDD.n7124 DVDD.n7123 0.0119575
R13062 DVDD.n7275 DVDD.n7118 0.0119575
R13063 DVDD.n7126 DVDD.n7125 0.0119575
R13064 DVDD.n7276 DVDD.n7117 0.0119575
R13065 DVDD.n7128 DVDD.n7127 0.0119575
R13066 DVDD.n7277 DVDD.n7116 0.0119575
R13067 DVDD.n7130 DVDD.n7129 0.0119575
R13068 DVDD.n7278 DVDD.n7115 0.0119575
R13069 DVDD.n7132 DVDD.n7131 0.0119575
R13070 DVDD.n7279 DVDD.n7114 0.0119575
R13071 DVDD.n7134 DVDD.n7133 0.0119575
R13072 DVDD.n7280 DVDD.n7111 0.0119575
R13073 DVDD.n7204 DVDD.n7203 0.0119575
R13074 DVDD.n7282 DVDD.n7110 0.0119575
R13075 DVDD.n7284 DVDD.n7283 0.0119575
R13076 DVDD.n7109 DVDD.n7105 0.0119575
R13077 DVDD.n7297 DVDD.n7287 0.0119575
R13078 DVDD.n7300 DVDD.n7103 0.0119575
R13079 DVDD.n7296 DVDD.n7288 0.0119575
R13080 DVDD.n7301 DVDD.n7102 0.0119575
R13081 DVDD.n7295 DVDD.n7289 0.0119575
R13082 DVDD.n7302 DVDD.n7101 0.0119575
R13083 DVDD.n7294 DVDD.n7290 0.0119575
R13084 DVDD.n7303 DVDD.n7100 0.0119575
R13085 DVDD.n7293 DVDD.n7291 0.0119575
R13086 DVDD.n7292 DVDD.n7099 0.0119575
R13087 DVDD.n1501 DVDD.n1498 0.0119575
R13088 DVDD.n4817 DVDD.n4739 0.0119575
R13089 DVDD.n4779 DVDD.n4747 0.0119575
R13090 DVDD.n4780 DVDD.n4746 0.0119575
R13091 DVDD.n4781 DVDD.n4778 0.0119575
R13092 DVDD.n4782 DVDD.n4745 0.0119575
R13093 DVDD.n4783 DVDD.n4777 0.0119575
R13094 DVDD.n4784 DVDD.n4744 0.0119575
R13095 DVDD.n4785 DVDD.n4776 0.0119575
R13096 DVDD.n4786 DVDD.n4743 0.0119575
R13097 DVDD.n4775 DVDD.n4774 0.0119575
R13098 DVDD.n32 DVDD.n31 0.0119575
R13099 DVDD.n33 DVDD.n29 0.0119575
R13100 DVDD.n35 DVDD.n34 0.0119575
R13101 DVDD.n36 DVDD.n28 0.0119575
R13102 DVDD.n38 DVDD.n37 0.0119575
R13103 DVDD.n39 DVDD.n27 0.0119575
R13104 DVDD.n41 DVDD.n40 0.0119575
R13105 DVDD.n42 DVDD.n26 0.0119575
R13106 DVDD.n44 DVDD.n43 0.0119575
R13107 DVDD.n45 DVDD.n25 0.0119575
R13108 DVDD.n6459 DVDD.n3421 0.0119301
R13109 DVDD.n7176 DVDD.n1888 0.0118386
R13110 DVDD.n7157 DVDD.n1857 0.0118386
R13111 DVDD.n7173 DVDD.n1889 0.0118386
R13112 DVDD.n7158 DVDD.n1856 0.0118386
R13113 DVDD.n7181 DVDD.n1672 0.0118386
R13114 DVDD.n7151 DVDD.n1662 0.0118386
R13115 DVDD.n7178 DVDD.n1673 0.0118386
R13116 DVDD.n7152 DVDD.n1682 0.0118386
R13117 DVDD.n7185 DVDD.n1608 0.0118386
R13118 DVDD.n7143 DVDD.n1591 0.0118386
R13119 DVDD.n7145 DVDD.n1609 0.0118386
R13120 DVDD.n7149 DVDD.n1590 0.0118386
R13121 DVDD.n7190 DVDD.n1555 0.0118386
R13122 DVDD.n7137 DVDD.n1536 0.0118386
R13123 DVDD.n7187 DVDD.n1556 0.0118386
R13124 DVDD.n7138 DVDD.n1535 0.0118386
R13125 DVDD.n7171 DVDD.n1264 0.0118386
R13126 DVDD.n7166 DVDD.n1241 0.0118386
R13127 DVDD.n7165 DVDD.n1265 0.0118386
R13128 DVDD.n7164 DVDD.n1240 0.0118386
R13129 DVDD.n7194 DVDD.n7135 0.0118386
R13130 DVDD.n7197 DVDD.n7112 0.0118386
R13131 DVDD.n7202 DVDD.n7136 0.0118386
R13132 DVDD.n7201 DVDD.n7111 0.0118386
R13133 DVDD.n3443 DVDD.n3407 0.0117899
R13134 DVDD.n6235 DVDD.n6234 0.01175
R13135 DVDD.n6883 DVDD.n6882 0.01175
R13136 DVDD.n9579 DVDD.n197 0.01175
R13137 DVDD.n9561 DVDD.n230 0.01175
R13138 DVDD.n9561 DVDD.n236 0.01175
R13139 DVDD.n9355 DVDD.n9354 0.01175
R13140 DVDD.n9579 DVDD.n189 0.01175
R13141 DVDD.n9354 DVDD.n102 0.01175
R13142 DVDD.n8770 DVDD.n114 0.0116614
R13143 DVDD.n6335 DVDD.n3559 0.0116614
R13144 DVDD.n6256 DVDD.n3340 0.0116614
R13145 DVDD.n4100 DVDD.n112 0.0116614
R13146 DVDD.n6050 DVDD.n3968 0.0116614
R13147 DVDD.n5947 DVDD.n3220 0.0116614
R13148 DVDD.n9461 DVDD.n125 0.0116614
R13149 DVDD.n5817 DVDD.n4315 0.0116614
R13150 DVDD.n5845 DVDD.n3105 0.0116614
R13151 DVDD.n411 DVDD.n126 0.0116614
R13152 DVDD.n6857 DVDD.n2806 0.0116614
R13153 DVDD.n6907 DVDD.n2734 0.0116614
R13154 DVDD.n4630 DVDD.n4628 0.01166
R13155 DVDD.n4632 DVDD.n4630 0.01166
R13156 DVDD.n4634 DVDD.n4632 0.01166
R13157 DVDD.n4636 DVDD.n4634 0.01166
R13158 DVDD.n4638 DVDD.n4636 0.01166
R13159 DVDD.n4640 DVDD.n4638 0.01166
R13160 DVDD.n4642 DVDD.n4640 0.01166
R13161 DVDD.n4644 DVDD.n4642 0.01166
R13162 DVDD.n4645 DVDD.n4644 0.01166
R13163 DVDD.n4705 DVDD.n4645 0.01166
R13164 DVDD.n4705 DVDD.n4704 0.01166
R13165 DVDD.n4704 DVDD.n4703 0.01166
R13166 DVDD.n4703 DVDD.n4646 0.01166
R13167 DVDD.n4699 DVDD.n4646 0.01166
R13168 DVDD.n4699 DVDD.n4698 0.01166
R13169 DVDD.n4698 DVDD.n4697 0.01166
R13170 DVDD.n4697 DVDD.n4567 0.01166
R13171 DVDD.n4692 DVDD.n4563 0.01166
R13172 DVDD.n4692 DVDD.n4691 0.01166
R13173 DVDD.n4691 DVDD.n4690 0.01166
R13174 DVDD.n4690 DVDD.n4649 0.01166
R13175 DVDD.n4686 DVDD.n4649 0.01166
R13176 DVDD.n4686 DVDD.n4685 0.01166
R13177 DVDD.n4685 DVDD.n4684 0.01166
R13178 DVDD.n4684 DVDD.n4651 0.01166
R13179 DVDD.n4680 DVDD.n4651 0.01166
R13180 DVDD.n4680 DVDD.n4679 0.01166
R13181 DVDD.n4679 DVDD.n4678 0.01166
R13182 DVDD.n4678 DVDD.n4653 0.01166
R13183 DVDD.n4674 DVDD.n4653 0.01166
R13184 DVDD.n4674 DVDD.n4673 0.01166
R13185 DVDD.n4673 DVDD.n4672 0.01166
R13186 DVDD.n4672 DVDD.n4655 0.01166
R13187 DVDD.n4668 DVDD.n4655 0.01166
R13188 DVDD.n4668 DVDD.n4667 0.01166
R13189 DVDD.n4667 DVDD.n4666 0.01166
R13190 DVDD.n4666 DVDD.n4657 0.01166
R13191 DVDD.n4662 DVDD.n4657 0.01166
R13192 DVDD.n4662 DVDD.n4661 0.01166
R13193 DVDD.n4661 DVDD.n4660 0.01166
R13194 DVDD.n4660 DVDD.n4561 0.01166
R13195 DVDD.n5217 DVDD.n4561 0.01166
R13196 DVDD.n5220 DVDD.n449 0.01166
R13197 DVDD.n5220 DVDD.n4559 0.01166
R13198 DVDD.n5224 DVDD.n4559 0.01166
R13199 DVDD.n5225 DVDD.n5224 0.01166
R13200 DVDD.n5226 DVDD.n5225 0.01166
R13201 DVDD.n5226 DVDD.n4557 0.01166
R13202 DVDD.n5230 DVDD.n4557 0.01166
R13203 DVDD.n5232 DVDD.n5230 0.01166
R13204 DVDD.n5234 DVDD.n5232 0.01166
R13205 DVDD.n5236 DVDD.n5234 0.01166
R13206 DVDD.n5238 DVDD.n5236 0.01166
R13207 DVDD.n5240 DVDD.n5238 0.01166
R13208 DVDD.n5242 DVDD.n5240 0.01166
R13209 DVDD.n5244 DVDD.n5242 0.01166
R13210 DVDD.n5245 DVDD.n5244 0.01166
R13211 DVDD.n5246 DVDD.n5245 0.01166
R13212 DVDD.n5246 DVDD.n4540 0.01166
R13213 DVDD.n5252 DVDD.n4540 0.01166
R13214 DVDD.n5253 DVDD.n5252 0.01166
R13215 DVDD.n5254 DVDD.n5253 0.01166
R13216 DVDD.n5254 DVDD.n4538 0.01166
R13217 DVDD.n5258 DVDD.n4538 0.01166
R13218 DVDD.n5259 DVDD.n5258 0.01166
R13219 DVDD.n5260 DVDD.n5259 0.01166
R13220 DVDD.n5260 DVDD.n448 0.01166
R13221 DVDD.n5265 DVDD.n4536 0.01166
R13222 DVDD.n4536 DVDD.n4535 0.01166
R13223 DVDD.n4535 DVDD.n4533 0.01166
R13224 DVDD.n4533 DVDD.n4526 0.01166
R13225 DVDD.n4526 DVDD.n407 0.01166
R13226 DVDD.n9364 DVDD.n407 0.01166
R13227 DVDD.n9366 DVDD.n9364 0.01166
R13228 DVDD.n9368 DVDD.n9366 0.01166
R13229 DVDD.n9369 DVDD.n9368 0.01166
R13230 DVDD.n9369 DVDD.n405 0.01166
R13231 DVDD.n9375 DVDD.n405 0.01166
R13232 DVDD.n9376 DVDD.n9375 0.01166
R13233 DVDD.n9376 DVDD.n404 0.01166
R13234 DVDD.n9380 DVDD.n404 0.01166
R13235 DVDD.n9381 DVDD.n9380 0.01166
R13236 DVDD.n9385 DVDD.n9381 0.01166
R13237 DVDD.n9387 DVDD.n9385 0.01166
R13238 DVDD.n9388 DVDD.n9387 0.01166
R13239 DVDD.n9388 DVDD.n379 0.01166
R13240 DVDD.n9422 DVDD.n379 0.01166
R13241 DVDD.n9422 DVDD.n9421 0.01166
R13242 DVDD.n9421 DVDD.n380 0.01166
R13243 DVDD.n4521 DVDD.n380 0.01166
R13244 DVDD.n4525 DVDD.n4521 0.01166
R13245 DVDD.n5266 DVDD.n4525 0.01166
R13246 DVDD.n5292 DVDD.n2887 0.01166
R13247 DVDD.n5294 DVDD.n5292 0.01166
R13248 DVDD.n5295 DVDD.n5294 0.01166
R13249 DVDD.n5295 DVDD.n4505 0.01166
R13250 DVDD.n5308 DVDD.n4505 0.01166
R13251 DVDD.n5310 DVDD.n5308 0.01166
R13252 DVDD.n5311 DVDD.n5310 0.01166
R13253 DVDD.n5312 DVDD.n5311 0.01166
R13254 DVDD.n5312 DVDD.n4503 0.01166
R13255 DVDD.n5316 DVDD.n4503 0.01166
R13256 DVDD.n5317 DVDD.n5316 0.01166
R13257 DVDD.n5318 DVDD.n5317 0.01166
R13258 DVDD.n5318 DVDD.n4501 0.01166
R13259 DVDD.n5322 DVDD.n4501 0.01166
R13260 DVDD.n5323 DVDD.n5322 0.01166
R13261 DVDD.n5324 DVDD.n5323 0.01166
R13262 DVDD.n5324 DVDD.n4499 0.01166
R13263 DVDD.n5328 DVDD.n4499 0.01166
R13264 DVDD.n5329 DVDD.n5328 0.01166
R13265 DVDD.n5330 DVDD.n5329 0.01166
R13266 DVDD.n5330 DVDD.n4497 0.01166
R13267 DVDD.n5334 DVDD.n4497 0.01166
R13268 DVDD.n5335 DVDD.n5334 0.01166
R13269 DVDD.n5336 DVDD.n5335 0.01166
R13270 DVDD.n5336 DVDD.n2886 0.01166
R13271 DVDD.n4495 DVDD.n2882 0.01166
R13272 DVDD.n5342 DVDD.n4495 0.01166
R13273 DVDD.n5343 DVDD.n5342 0.01166
R13274 DVDD.n5344 DVDD.n5343 0.01166
R13275 DVDD.n5344 DVDD.n4493 0.01166
R13276 DVDD.n5348 DVDD.n4493 0.01166
R13277 DVDD.n5349 DVDD.n5348 0.01166
R13278 DVDD.n5350 DVDD.n5349 0.01166
R13279 DVDD.n5350 DVDD.n4491 0.01166
R13280 DVDD.n5354 DVDD.n4491 0.01166
R13281 DVDD.n5355 DVDD.n5354 0.01166
R13282 DVDD.n5356 DVDD.n5355 0.01166
R13283 DVDD.n5356 DVDD.n4489 0.01166
R13284 DVDD.n5360 DVDD.n4489 0.01166
R13285 DVDD.n5361 DVDD.n5360 0.01166
R13286 DVDD.n5362 DVDD.n5361 0.01166
R13287 DVDD.n5362 DVDD.n4487 0.01166
R13288 DVDD.n5366 DVDD.n4487 0.01166
R13289 DVDD.n5367 DVDD.n5366 0.01166
R13290 DVDD.n5368 DVDD.n5367 0.01166
R13291 DVDD.n5368 DVDD.n4485 0.01166
R13292 DVDD.n5372 DVDD.n4485 0.01166
R13293 DVDD.n5373 DVDD.n5372 0.01166
R13294 DVDD.n5374 DVDD.n5373 0.01166
R13295 DVDD.n5374 DVDD.n2881 0.01166
R13296 DVDD.n5432 DVDD.n2801 0.01166
R13297 DVDD.n5434 DVDD.n5432 0.01166
R13298 DVDD.n5436 DVDD.n5434 0.01166
R13299 DVDD.n5438 DVDD.n5436 0.01166
R13300 DVDD.n5440 DVDD.n5438 0.01166
R13301 DVDD.n5442 DVDD.n5440 0.01166
R13302 DVDD.n5444 DVDD.n5442 0.01166
R13303 DVDD.n5446 DVDD.n5444 0.01166
R13304 DVDD.n5448 DVDD.n5446 0.01166
R13305 DVDD.n5450 DVDD.n5448 0.01166
R13306 DVDD.n5452 DVDD.n5450 0.01166
R13307 DVDD.n5454 DVDD.n5452 0.01166
R13308 DVDD.n5456 DVDD.n5454 0.01166
R13309 DVDD.n5458 DVDD.n5456 0.01166
R13310 DVDD.n5460 DVDD.n5458 0.01166
R13311 DVDD.n5462 DVDD.n5460 0.01166
R13312 DVDD.n5463 DVDD.n5462 0.01166
R13313 DVDD.n5463 DVDD.n4468 0.01166
R13314 DVDD.n5469 DVDD.n4468 0.01166
R13315 DVDD.n5470 DVDD.n5469 0.01166
R13316 DVDD.n5470 DVDD.n4466 0.01166
R13317 DVDD.n5474 DVDD.n4466 0.01166
R13318 DVDD.n5476 DVDD.n5474 0.01166
R13319 DVDD.n5477 DVDD.n5476 0.01166
R13320 DVDD.n5477 DVDD.n2800 0.01166
R13321 DVDD.n5638 DVDD.n2740 0.01166
R13322 DVDD.n5638 DVDD.n5637 0.01166
R13323 DVDD.n5637 DVDD.n5636 0.01166
R13324 DVDD.n5636 DVDD.n5485 0.01166
R13325 DVDD.n5632 DVDD.n5485 0.01166
R13326 DVDD.n5632 DVDD.n5631 0.01166
R13327 DVDD.n5631 DVDD.n5630 0.01166
R13328 DVDD.n5630 DVDD.n5487 0.01166
R13329 DVDD.n5626 DVDD.n5487 0.01166
R13330 DVDD.n5626 DVDD.n5625 0.01166
R13331 DVDD.n5625 DVDD.n5624 0.01166
R13332 DVDD.n5624 DVDD.n5489 0.01166
R13333 DVDD.n5620 DVDD.n5489 0.01166
R13334 DVDD.n5620 DVDD.n5619 0.01166
R13335 DVDD.n5619 DVDD.n5618 0.01166
R13336 DVDD.n5618 DVDD.n5491 0.01166
R13337 DVDD.n5535 DVDD.n5491 0.01166
R13338 DVDD.n5537 DVDD.n5535 0.01166
R13339 DVDD.n5539 DVDD.n5537 0.01166
R13340 DVDD.n5541 DVDD.n5539 0.01166
R13341 DVDD.n5543 DVDD.n5541 0.01166
R13342 DVDD.n5545 DVDD.n5543 0.01166
R13343 DVDD.n5546 DVDD.n5545 0.01166
R13344 DVDD.n5547 DVDD.n5546 0.01166
R13345 DVDD.n5547 DVDD.n2739 0.01166
R13346 DVDD.n5568 DVDD.n2653 0.01166
R13347 DVDD.n5570 DVDD.n5568 0.01166
R13348 DVDD.n5572 DVDD.n5570 0.01166
R13349 DVDD.n5574 DVDD.n5572 0.01166
R13350 DVDD.n5576 DVDD.n5574 0.01166
R13351 DVDD.n5578 DVDD.n5576 0.01166
R13352 DVDD.n5579 DVDD.n5578 0.01166
R13353 DVDD.n5611 DVDD.n5579 0.01166
R13354 DVDD.n5611 DVDD.n5610 0.01166
R13355 DVDD.n5610 DVDD.n5609 0.01166
R13356 DVDD.n5609 DVDD.n5607 0.01166
R13357 DVDD.n5607 DVDD.n5605 0.01166
R13358 DVDD.n5605 DVDD.n5603 0.01166
R13359 DVDD.n5603 DVDD.n5601 0.01166
R13360 DVDD.n5601 DVDD.n5599 0.01166
R13361 DVDD.n5599 DVDD.n5597 0.01166
R13362 DVDD.n5597 DVDD.n5595 0.01166
R13363 DVDD.n5595 DVDD.n5593 0.01166
R13364 DVDD.n5593 DVDD.n5591 0.01166
R13365 DVDD.n5591 DVDD.n5589 0.01166
R13366 DVDD.n5589 DVDD.n5587 0.01166
R13367 DVDD.n5587 DVDD.n5585 0.01166
R13368 DVDD.n5585 DVDD.n5583 0.01166
R13369 DVDD.n5583 DVDD.n5581 0.01166
R13370 DVDD.n5581 DVDD.n2652 0.01166
R13371 DVDD.n743 DVDD.n741 0.01166
R13372 DVDD.n741 DVDD.n739 0.01166
R13373 DVDD.n739 DVDD.n737 0.01166
R13374 DVDD.n737 DVDD.n735 0.01166
R13375 DVDD.n735 DVDD.n733 0.01166
R13376 DVDD.n733 DVDD.n731 0.01166
R13377 DVDD.n731 DVDD.n729 0.01166
R13378 DVDD.n729 DVDD.n727 0.01166
R13379 DVDD.n727 DVDD.n656 0.01166
R13380 DVDD.n8887 DVDD.n656 0.01166
R13381 DVDD.n8887 DVDD.n8886 0.01166
R13382 DVDD.n8886 DVDD.n8885 0.01166
R13383 DVDD.n8885 DVDD.n657 0.01166
R13384 DVDD.n8881 DVDD.n657 0.01166
R13385 DVDD.n8881 DVDD.n8880 0.01166
R13386 DVDD.n8880 DVDD.n8879 0.01166
R13387 DVDD.n8879 DVDD.n659 0.01166
R13388 DVDD.n8875 DVDD.n8874 0.01166
R13389 DVDD.n8874 DVDD.n8873 0.01166
R13390 DVDD.n8873 DVDD.n661 0.01166
R13391 DVDD.n8869 DVDD.n661 0.01166
R13392 DVDD.n8869 DVDD.n8868 0.01166
R13393 DVDD.n8868 DVDD.n8867 0.01166
R13394 DVDD.n8867 DVDD.n663 0.01166
R13395 DVDD.n8863 DVDD.n663 0.01166
R13396 DVDD.n8863 DVDD.n8862 0.01166
R13397 DVDD.n8862 DVDD.n8861 0.01166
R13398 DVDD.n8861 DVDD.n665 0.01166
R13399 DVDD.n8857 DVDD.n665 0.01166
R13400 DVDD.n8857 DVDD.n8856 0.01166
R13401 DVDD.n8856 DVDD.n8855 0.01166
R13402 DVDD.n8855 DVDD.n667 0.01166
R13403 DVDD.n8851 DVDD.n667 0.01166
R13404 DVDD.n8851 DVDD.n8850 0.01166
R13405 DVDD.n8850 DVDD.n8849 0.01166
R13406 DVDD.n8849 DVDD.n669 0.01166
R13407 DVDD.n8845 DVDD.n669 0.01166
R13408 DVDD.n8845 DVDD.n8844 0.01166
R13409 DVDD.n8844 DVDD.n8843 0.01166
R13410 DVDD.n8843 DVDD.n671 0.01166
R13411 DVDD.n8839 DVDD.n671 0.01166
R13412 DVDD.n8839 DVDD.n8838 0.01166
R13413 DVDD.n798 DVDD.n790 0.01166
R13414 DVDD.n798 DVDD.n796 0.01166
R13415 DVDD.n802 DVDD.n796 0.01166
R13416 DVDD.n803 DVDD.n802 0.01166
R13417 DVDD.n804 DVDD.n803 0.01166
R13418 DVDD.n804 DVDD.n794 0.01166
R13419 DVDD.n808 DVDD.n794 0.01166
R13420 DVDD.n810 DVDD.n808 0.01166
R13421 DVDD.n812 DVDD.n810 0.01166
R13422 DVDD.n814 DVDD.n812 0.01166
R13423 DVDD.n816 DVDD.n814 0.01166
R13424 DVDD.n818 DVDD.n816 0.01166
R13425 DVDD.n820 DVDD.n818 0.01166
R13426 DVDD.n822 DVDD.n820 0.01166
R13427 DVDD.n824 DVDD.n822 0.01166
R13428 DVDD.n826 DVDD.n824 0.01166
R13429 DVDD.n827 DVDD.n826 0.01166
R13430 DVDD.n828 DVDD.n827 0.01166
R13431 DVDD.n829 DVDD.n828 0.01166
R13432 DVDD.n829 DVDD.n793 0.01166
R13433 DVDD.n833 DVDD.n793 0.01166
R13434 DVDD.n834 DVDD.n833 0.01166
R13435 DVDD.n835 DVDD.n834 0.01166
R13436 DVDD.n835 DVDD.n791 0.01166
R13437 DVDD.n8796 DVDD.n791 0.01166
R13438 DVDD.n8793 DVDD.n8792 0.01166
R13439 DVDD.n8792 DVDD.n8791 0.01166
R13440 DVDD.n8791 DVDD.n8780 0.01166
R13441 DVDD.n8780 DVDD.n8776 0.01166
R13442 DVDD.n8776 DVDD.n8775 0.01166
R13443 DVDD.n8775 DVDD.n839 0.01166
R13444 DVDD.n925 DVDD.n839 0.01166
R13445 DVDD.n927 DVDD.n925 0.01166
R13446 DVDD.n928 DVDD.n927 0.01166
R13447 DVDD.n945 DVDD.n928 0.01166
R13448 DVDD.n947 DVDD.n945 0.01166
R13449 DVDD.n948 DVDD.n947 0.01166
R13450 DVDD.n948 DVDD.n922 0.01166
R13451 DVDD.n952 DVDD.n922 0.01166
R13452 DVDD.n953 DVDD.n952 0.01166
R13453 DVDD.n953 DVDD.n921 0.01166
R13454 DVDD.n980 DVDD.n921 0.01166
R13455 DVDD.n982 DVDD.n980 0.01166
R13456 DVDD.n984 DVDD.n982 0.01166
R13457 DVDD.n986 DVDD.n984 0.01166
R13458 DVDD.n988 DVDD.n986 0.01166
R13459 DVDD.n990 DVDD.n988 0.01166
R13460 DVDD.n991 DVDD.n990 0.01166
R13461 DVDD.n991 DVDD.n913 0.01166
R13462 DVDD.n1000 DVDD.n913 0.01166
R13463 DVDD.n3750 DVDD.n3746 0.01166
R13464 DVDD.n3746 DVDD.n3745 0.01166
R13465 DVDD.n3745 DVDD.n3583 0.01166
R13466 DVDD.n3631 DVDD.n3583 0.01166
R13467 DVDD.n3631 DVDD.n3630 0.01166
R13468 DVDD.n3630 DVDD.n3592 0.01166
R13469 DVDD.n3625 DVDD.n3592 0.01166
R13470 DVDD.n3625 DVDD.n3624 0.01166
R13471 DVDD.n3624 DVDD.n3623 0.01166
R13472 DVDD.n3623 DVDD.n3594 0.01166
R13473 DVDD.n3619 DVDD.n3594 0.01166
R13474 DVDD.n3619 DVDD.n3618 0.01166
R13475 DVDD.n3618 DVDD.n3617 0.01166
R13476 DVDD.n3617 DVDD.n3596 0.01166
R13477 DVDD.n3613 DVDD.n3596 0.01166
R13478 DVDD.n3613 DVDD.n3612 0.01166
R13479 DVDD.n3612 DVDD.n3611 0.01166
R13480 DVDD.n3611 DVDD.n3598 0.01166
R13481 DVDD.n3607 DVDD.n3598 0.01166
R13482 DVDD.n3607 DVDD.n3606 0.01166
R13483 DVDD.n3606 DVDD.n3605 0.01166
R13484 DVDD.n3605 DVDD.n3600 0.01166
R13485 DVDD.n3601 DVDD.n3600 0.01166
R13486 DVDD.n3601 DVDD.n3580 0.01166
R13487 DVDD.n3751 DVDD.n3580 0.01166
R13488 DVDD.n3802 DVDD.n3578 0.01166
R13489 DVDD.n3798 DVDD.n3578 0.01166
R13490 DVDD.n3798 DVDD.n3797 0.01166
R13491 DVDD.n3797 DVDD.n3796 0.01166
R13492 DVDD.n3796 DVDD.n3754 0.01166
R13493 DVDD.n3792 DVDD.n3754 0.01166
R13494 DVDD.n3792 DVDD.n3791 0.01166
R13495 DVDD.n3791 DVDD.n3790 0.01166
R13496 DVDD.n3790 DVDD.n3756 0.01166
R13497 DVDD.n3786 DVDD.n3756 0.01166
R13498 DVDD.n3786 DVDD.n3785 0.01166
R13499 DVDD.n3785 DVDD.n3784 0.01166
R13500 DVDD.n3784 DVDD.n3758 0.01166
R13501 DVDD.n3780 DVDD.n3758 0.01166
R13502 DVDD.n3780 DVDD.n3779 0.01166
R13503 DVDD.n3779 DVDD.n3778 0.01166
R13504 DVDD.n3778 DVDD.n3760 0.01166
R13505 DVDD.n3774 DVDD.n3760 0.01166
R13506 DVDD.n3774 DVDD.n3773 0.01166
R13507 DVDD.n3773 DVDD.n3772 0.01166
R13508 DVDD.n3772 DVDD.n3762 0.01166
R13509 DVDD.n3768 DVDD.n3762 0.01166
R13510 DVDD.n3768 DVDD.n3767 0.01166
R13511 DVDD.n3767 DVDD.n3766 0.01166
R13512 DVDD.n3766 DVDD.n3576 0.01166
R13513 DVDD.n6375 DVDD.n6373 0.01166
R13514 DVDD.n6373 DVDD.n6371 0.01166
R13515 DVDD.n6371 DVDD.n6369 0.01166
R13516 DVDD.n6369 DVDD.n6367 0.01166
R13517 DVDD.n6367 DVDD.n6365 0.01166
R13518 DVDD.n6365 DVDD.n6363 0.01166
R13519 DVDD.n6363 DVDD.n6361 0.01166
R13520 DVDD.n6361 DVDD.n6359 0.01166
R13521 DVDD.n6359 DVDD.n6357 0.01166
R13522 DVDD.n6357 DVDD.n6355 0.01166
R13523 DVDD.n6355 DVDD.n6353 0.01166
R13524 DVDD.n6353 DVDD.n6351 0.01166
R13525 DVDD.n6351 DVDD.n6349 0.01166
R13526 DVDD.n6349 DVDD.n6347 0.01166
R13527 DVDD.n6347 DVDD.n6345 0.01166
R13528 DVDD.n6345 DVDD.n6343 0.01166
R13529 DVDD.n6343 DVDD.n6341 0.01166
R13530 DVDD.n6341 DVDD.n6339 0.01166
R13531 DVDD.n6339 DVDD.n3553 0.01166
R13532 DVDD.n6385 DVDD.n3553 0.01166
R13533 DVDD.n6385 DVDD.n6384 0.01166
R13534 DVDD.n6384 DVDD.n6383 0.01166
R13535 DVDD.n6383 DVDD.n6381 0.01166
R13536 DVDD.n6381 DVDD.n6379 0.01166
R13537 DVDD.n6379 DVDD.n6377 0.01166
R13538 DVDD.n6467 DVDD.n3418 0.01166
R13539 DVDD.n3464 DVDD.n3418 0.01166
R13540 DVDD.n3464 DVDD.n3463 0.01166
R13541 DVDD.n3463 DVDD.n3462 0.01166
R13542 DVDD.n3462 DVDD.n3423 0.01166
R13543 DVDD.n3458 DVDD.n3423 0.01166
R13544 DVDD.n3458 DVDD.n3457 0.01166
R13545 DVDD.n3457 DVDD.n3456 0.01166
R13546 DVDD.n3456 DVDD.n3425 0.01166
R13547 DVDD.n3452 DVDD.n3425 0.01166
R13548 DVDD.n3452 DVDD.n3451 0.01166
R13549 DVDD.n3451 DVDD.n3450 0.01166
R13550 DVDD.n3450 DVDD.n3427 0.01166
R13551 DVDD.n3446 DVDD.n3427 0.01166
R13552 DVDD.n3446 DVDD.n3445 0.01166
R13553 DVDD.n3445 DVDD.n3444 0.01166
R13554 DVDD.n3444 DVDD.n3442 0.01166
R13555 DVDD.n3442 DVDD.n3440 0.01166
R13556 DVDD.n3440 DVDD.n3438 0.01166
R13557 DVDD.n3438 DVDD.n3436 0.01166
R13558 DVDD.n3436 DVDD.n3434 0.01166
R13559 DVDD.n3434 DVDD.n3432 0.01166
R13560 DVDD.n3432 DVDD.n3430 0.01166
R13561 DVDD.n3430 DVDD.n3414 0.01166
R13562 DVDD.n6468 DVDD.n3414 0.01166
R13563 DVDD.n6557 DVDD.n6555 0.01166
R13564 DVDD.n6555 DVDD.n6553 0.01166
R13565 DVDD.n6553 DVDD.n6551 0.01166
R13566 DVDD.n6551 DVDD.n6549 0.01166
R13567 DVDD.n6549 DVDD.n6547 0.01166
R13568 DVDD.n6547 DVDD.n6545 0.01166
R13569 DVDD.n6545 DVDD.n6487 0.01166
R13570 DVDD.n6591 DVDD.n6487 0.01166
R13571 DVDD.n6591 DVDD.n6590 0.01166
R13572 DVDD.n6590 DVDD.n6589 0.01166
R13573 DVDD.n6589 DVDD.n6587 0.01166
R13574 DVDD.n6587 DVDD.n6585 0.01166
R13575 DVDD.n6585 DVDD.n6583 0.01166
R13576 DVDD.n6583 DVDD.n6581 0.01166
R13577 DVDD.n6581 DVDD.n6579 0.01166
R13578 DVDD.n6579 DVDD.n6577 0.01166
R13579 DVDD.n6577 DVDD.n6575 0.01166
R13580 DVDD.n6575 DVDD.n6573 0.01166
R13581 DVDD.n6573 DVDD.n6571 0.01166
R13582 DVDD.n6571 DVDD.n6569 0.01166
R13583 DVDD.n6569 DVDD.n6567 0.01166
R13584 DVDD.n6567 DVDD.n6565 0.01166
R13585 DVDD.n6565 DVDD.n6563 0.01166
R13586 DVDD.n6563 DVDD.n6561 0.01166
R13587 DVDD.n6561 DVDD.n6559 0.01166
R13588 DVDD.n6380 DVDD.n3474 0.0116088
R13589 DVDD.n6378 DVDD.n3472 0.0116088
R13590 DVDD.n6376 DVDD.n3475 0.0116088
R13591 DVDD.n8688 DVDD.n1008 0.011525
R13592 DVDD.n890 DVDD.n357 0.011525
R13593 DVDD.n6309 DVDD.n3878 0.011525
R13594 DVDD.n6887 DVDD.n6885 0.011525
R13595 DVDD.n9400 DVDD.n374 0.011525
R13596 DVDD.n4512 DVDD.n4511 0.011525
R13597 DVDD.n9359 DVDD.n109 0.011525
R13598 DVDD.n9617 DVDD.n94 0.011525
R13599 DVDD.n8771 DVDD.n8770 0.0113071
R13600 DVDD.n3809 DVDD.n3559 0.0113071
R13601 DVDD.n6299 DVDD.n6298 0.0113071
R13602 DVDD.n6256 DVDD.n3348 0.0113071
R13603 DVDD.n4101 DVDD.n4100 0.0113071
R13604 DVDD.n6050 DVDD.n3949 0.0113071
R13605 DVDD.n5989 DVDD.n5929 0.0113071
R13606 DVDD.n5947 DVDD.n3234 0.0113071
R13607 DVDD.n9461 DVDD.n297 0.0113071
R13608 DVDD.n5817 DVDD.n4378 0.0113071
R13609 DVDD.n6096 DVDD.n5887 0.0113071
R13610 DVDD.n5845 DVDD.n3113 0.0113071
R13611 DVDD.n9360 DVDD.n411 0.0113071
R13612 DVDD.n2810 DVDD.n2806 0.0113071
R13613 DVDD.n6900 DVDD.n2776 0.0113071
R13614 DVDD.n6907 DVDD.n2664 0.0113071
R13615 DVDD.n6452 DVDD.n3483 0.0111617
R13616 DVDD.n7176 DVDD.n1895 0.0111299
R13617 DVDD.n7157 DVDD.n1888 0.0111299
R13618 DVDD.n7173 DVDD.n1857 0.0111299
R13619 DVDD.n7158 DVDD.n1889 0.0111299
R13620 DVDD.n7181 DVDD.n1663 0.0111299
R13621 DVDD.n7151 DVDD.n1672 0.0111299
R13622 DVDD.n7178 DVDD.n1662 0.0111299
R13623 DVDD.n7152 DVDD.n1673 0.0111299
R13624 DVDD.n7185 DVDD.n1592 0.0111299
R13625 DVDD.n7143 DVDD.n1608 0.0111299
R13626 DVDD.n7145 DVDD.n1591 0.0111299
R13627 DVDD.n7149 DVDD.n1609 0.0111299
R13628 DVDD.n7190 DVDD.n1537 0.0111299
R13629 DVDD.n7137 DVDD.n1555 0.0111299
R13630 DVDD.n7187 DVDD.n1536 0.0111299
R13631 DVDD.n7138 DVDD.n1556 0.0111299
R13632 DVDD.n7171 DVDD.n1242 0.0111299
R13633 DVDD.n7166 DVDD.n1264 0.0111299
R13634 DVDD.n7165 DVDD.n1241 0.0111299
R13635 DVDD.n7164 DVDD.n1265 0.0111299
R13636 DVDD.n7194 DVDD.n7113 0.0111299
R13637 DVDD.n7197 DVDD.n7135 0.0111299
R13638 DVDD.n7136 DVDD.n7112 0.0111299
R13639 DVDD.n7202 DVDD.n7201 0.0111299
R13640 DVDD.n5475 DVDD.n4465 0.0109528
R13641 DVDD.n5478 DVDD.n4464 0.0109528
R13642 DVDD.n5480 DVDD.n5479 0.0109528
R13643 DVDD.n713 DVDD.n578 0.0109528
R13644 DVDD.n8720 DVDD.n8719 0.0109528
R13645 DVDD.n3834 DVDD.n3812 0.0109528
R13646 DVDD.n1884 DVDD.n1864 0.0109528
R13647 DVDD.n8985 DVDD.n8975 0.0109528
R13648 DVDD.n4074 DVDD.n4073 0.0109528
R13649 DVDD.n6034 DVDD.n3952 0.0109528
R13650 DVDD.n1687 DVDD.n1679 0.0109528
R13651 DVDD.n5022 DVDD.n4864 0.0109528
R13652 DVDD.n369 DVDD.n364 0.0109528
R13653 DVDD.n5801 DVDD.n4381 0.0109528
R13654 DVDD.n1871 DVDD.n1598 0.0109528
R13655 DVDD.n5129 DVDD.n5119 0.0109528
R13656 DVDD.n9399 DVDD.n401 0.0109528
R13657 DVDD.n2861 DVDD.n2813 0.0109528
R13658 DVDD.n1562 DVDD.n1543 0.0109528
R13659 DVDD.n3441 DVDD.n3409 0.0108556
R13660 DVDD.n3439 DVDD.n3406 0.0108556
R13661 DVDD.n3437 DVDD.n3410 0.0108556
R13662 DVDD.n3435 DVDD.n3405 0.0108556
R13663 DVDD.n3433 DVDD.n3411 0.0108556
R13664 DVDD.n3431 DVDD.n3404 0.0108556
R13665 DVDD.n3429 DVDD.n3412 0.0108556
R13666 DVDD.n3413 DVDD.n3403 0.0108556
R13667 DVDD.n6470 DVDD.n6469 0.0108556
R13668 DVDD.n954 DVDD.n872 0.01085
R13669 DVDD.n956 DVDD.n955 0.01085
R13670 DVDD.n979 DVDD.n978 0.01085
R13671 DVDD.n981 DVDD.n884 0.01085
R13672 DVDD.n983 DVDD.n886 0.01085
R13673 DVDD.n985 DVDD.n350 0.01085
R13674 DVDD.n987 DVDD.n892 0.01085
R13675 DVDD.n989 DVDD.n895 0.01085
R13676 DVDD.n992 DVDD.n920 0.01085
R13677 DVDD.n994 DVDD.n993 0.01085
R13678 DVDD.n1001 DVDD.n908 0.01085
R13679 DVDD.n6588 DVDD.n2042 0.010817
R13680 DVDD.n8406 DVDD.n1489 0.0107926
R13681 DVDD.n8468 DVDD.n8467 0.0107926
R13682 DVDD.n1383 DVDD.n1381 0.0107926
R13683 DVDD.n8490 DVDD.n1438 0.0107926
R13684 DVDD.n8558 DVDD.n1390 0.0107926
R13685 DVDD.n8605 DVDD.n1348 0.0107926
R13686 DVDD.n7716 DVDD.n1860 0.0107756
R13687 DVDD.n7722 DVDD.n1684 0.0107756
R13688 DVDD.n2345 DVDD.n1594 0.0107756
R13689 DVDD.n2350 DVDD.n1539 0.0107756
R13690 DVDD.n6253 DVDD.n3343 0.0105984
R13691 DVDD.n6492 DVDD.n2089 0.0105984
R13692 DVDD.n5964 DVDD.n3232 0.0105984
R13693 DVDD.n3255 DVDD.n2137 0.0105984
R13694 DVDD.n5839 DVDD.n3108 0.0105984
R13695 DVDD.n3146 DVDD.n2186 0.0105984
R13696 DVDD.n6923 DVDD.n2737 0.0105984
R13697 DVDD.n6932 DVDD.n2649 0.0105984
R13698 DVDD.n6234 DVDD.n3881 0.01055
R13699 DVDD.n6882 DVDD.n6881 0.01055
R13700 DVDD.n9580 DVDD.n9579 0.01055
R13701 DVDD.n9561 DVDD.n233 0.01055
R13702 DVDD.n9561 DVDD.n238 0.01055
R13703 DVDD.n9354 DVDD.n9353 0.01055
R13704 DVDD.n9579 DVDD.n194 0.01055
R13705 DVDD.n9354 DVDD.n421 0.01055
R13706 DVDD.n2338 DVDD.n2336 0.0105466
R13707 DVDD.n7733 DVDD.n7730 0.0105466
R13708 DVDD.n8625 DVDD.n1322 0.0105466
R13709 DVDD.n8439 DVDD.n1447 0.0105466
R13710 DVDD.n1448 DVDD.n1432 0.0105466
R13711 DVDD.n1433 DVDD.n1429 0.0105466
R13712 DVDD.n1430 DVDD.n1354 0.0105466
R13713 DVDD.n1355 DVDD.n1353 0.0105466
R13714 DVDD.n8598 DVDD.n1359 0.0105466
R13715 DVDD.n8533 DVDD.n8522 0.0105466
R13716 DVDD.n8533 DVDD.n1360 0.0105466
R13717 DVDD.n1447 DVDD.n1328 0.0105466
R13718 DVDD.n8627 DVDD.n1322 0.0105466
R13719 DVDD.n8439 DVDD.n1448 0.0105466
R13720 DVDD.n8495 DVDD.n1433 0.0105466
R13721 DVDD.n1430 DVDD.n1429 0.0105466
R13722 DVDD.n8600 DVDD.n1355 0.0105466
R13723 DVDD.n1359 DVDD.n1353 0.0105466
R13724 DVDD.n7742 DVDD.n7739 0.0105466
R13725 DVDD.n7745 DVDD.n2332 0.0105466
R13726 DVDD.n8622 DVDD.n1331 0.0105466
R13727 DVDD.n8434 DVDD.n1452 0.0105466
R13728 DVDD.n1453 DVDD.n1424 0.0105466
R13729 DVDD.n1425 DVDD.n1421 0.0105466
R13730 DVDD.n1422 DVDD.n1363 0.0105466
R13731 DVDD.n1364 DVDD.n1362 0.0105466
R13732 DVDD.n8593 DVDD.n1368 0.0105466
R13733 DVDD.n8540 DVDD.n8518 0.0105466
R13734 DVDD.n8518 DVDD.n1369 0.0105466
R13735 DVDD.n1452 DVDD.n1334 0.0105466
R13736 DVDD.n1331 DVDD.n1330 0.0105466
R13737 DVDD.n8434 DVDD.n1453 0.0105466
R13738 DVDD.n8499 DVDD.n1425 0.0105466
R13739 DVDD.n1422 DVDD.n1421 0.0105466
R13740 DVDD.n8595 DVDD.n1364 0.0105466
R13741 DVDD.n1368 DVDD.n1362 0.0105466
R13742 DVDD.n7742 DVDD.n2332 0.0105466
R13743 DVDD.n7730 DVDD.n2336 0.0105466
R13744 DVDD.n7739 DVDD.n2150 0.0105466
R13745 DVDD.n7735 DVDD.n2338 0.0105466
R13746 DVDD.n2361 DVDD.n2359 0.0105466
R13747 DVDD.n2367 DVDD.n2364 0.0105466
R13748 DVDD.n7346 DVDD.n1458 0.0105466
R13749 DVDD.n1459 DVDD.n1457 0.0105466
R13750 DVDD.n8423 DVDD.n1418 0.0105466
R13751 DVDD.n1420 DVDD.n1416 0.0105466
R13752 DVDD.n8508 DVDD.n1412 0.0105466
R13753 DVDD.n8510 DVDD.n1410 0.0105466
R13754 DVDD.n8514 DVDD.n1406 0.0105466
R13755 DVDD.n8544 DVDD.n1403 0.0105466
R13756 DVDD.n2364 DVDD.n2359 0.0105466
R13757 DVDD.n2369 DVDD.n2361 0.0105466
R13758 DVDD.n8516 DVDD.n1403 0.0105466
R13759 DVDD.n8427 DVDD.n1459 0.0105466
R13760 DVDD.n7358 DVDD.n7346 0.0105466
R13761 DVDD.n8423 DVDD.n1457 0.0105466
R13762 DVDD.n8505 DVDD.n1420 0.0105466
R13763 DVDD.n1416 DVDD.n1412 0.0105466
R13764 DVDD.n8511 DVDD.n8510 0.0105466
R13765 DVDD.n1410 DVDD.n1406 0.0105466
R13766 DVDD.n2356 DVDD.n2353 0.0105466
R13767 DVDD.n7683 DVDD.n2371 0.0105466
R13768 DVDD.n7350 DVDD.n1462 0.0105466
R13769 DVDD.n1463 DVDD.n1461 0.0105466
R13770 DVDD.n8417 DVDD.n1467 0.0105466
R13771 DVDD.n1471 DVDD.n1468 0.0105466
R13772 DVDD.n1486 DVDD.n1473 0.0105466
R13773 DVDD.n1477 DVDD.n1474 0.0105466
R13774 DVDD.n1481 DVDD.n1479 0.0105466
R13775 DVDD.n8547 DVDD.n1397 0.0105466
R13776 DVDD.n2371 DVDD.n2353 0.0105466
R13777 DVDD.n7685 DVDD.n2356 0.0105466
R13778 DVDD.n1401 DVDD.n1397 0.0105466
R13779 DVDD.n8419 DVDD.n1463 0.0105466
R13780 DVDD.n7350 DVDD.n1506 0.0105466
R13781 DVDD.n1467 DVDD.n1461 0.0105466
R13782 DVDD.n1488 DVDD.n1468 0.0105466
R13783 DVDD.n1473 DVDD.n1471 0.0105466
R13784 DVDD.n1483 DVDD.n1474 0.0105466
R13785 DVDD.n1479 DVDD.n1477 0.0105466
R13786 DVDD.n8451 DVDD.n8447 0.0105466
R13787 DVDD.n8466 DVDD.n8465 0.0105466
R13788 DVDD.n8449 DVDD.n8447 0.0105466
R13789 DVDD.n8492 DVDD.n8491 0.0105466
R13790 DVDD.n8442 DVDD.n1444 0.0105466
R13791 DVDD.n8606 DVDD.n1349 0.0105466
R13792 DVDD.n8489 DVDD.n1437 0.0105466
R13793 DVDD.n8604 DVDD.n8603 0.0105466
R13794 DVDD.n1496 DVDD.n1495 0.0105466
R13795 DVDD.n8414 DVDD.n8407 0.0105466
R13796 DVDD.n8574 DVDD.n8573 0.0105466
R13797 DVDD.n8556 DVDD.n1394 0.0105466
R13798 DVDD.n8387 DVDD.n1496 0.0105466
R13799 DVDD.n1391 DVDD.n1388 0.0105466
R13800 DVDD.n8577 DVDD.n8576 0.0105466
R13801 DVDD.n8405 DVDD.n8404 0.0105466
R13802 DVDD.n151 DVDD.n146 0.0104
R13803 DVDD.n9340 DVDD.n9339 0.0104
R13804 DVDD.n9443 DVDD.n9442 0.0104
R13805 DVDD.n4023 DVDD.n4022 0.0104
R13806 DVDD.n9444 DVDD.n323 0.0104
R13807 DVDD.n966 DVDD.n957 0.0104
R13808 DVDD.n4088 DVDD.n4087 0.0104
R13809 DVDD.n965 DVDD.n870 0.0104
R13810 DVDD.n3498 DVDD.n3497 0.0103933
R13811 DVDD.n6604 DVDD.n6592 0.0103305
R13812 DVDD.n5616 DVDD.n5615 0.0102441
R13813 DVDD.n5531 DVDD.n5494 0.0102441
R13814 DVDD.n5536 DVDD.n5507 0.0102441
R13815 DVDD.n5538 DVDD.n5532 0.0102441
R13816 DVDD.n5540 DVDD.n5506 0.0102441
R13817 DVDD.n5542 DVDD.n5533 0.0102441
R13818 DVDD.n5544 DVDD.n5505 0.0102441
R13819 DVDD.n5549 DVDD.n5534 0.0102441
R13820 DVDD.n5548 DVDD.n5504 0.0102441
R13821 DVDD.n5552 DVDD.n5550 0.0102441
R13822 DVDD.n8810 DVDD.n62 0.0102441
R13823 DVDD.n3850 DVDD.n3564 0.0102441
R13824 DVDD.n6328 DVDD.n6327 0.0102441
R13825 DVDD.n6538 DVDD.n3353 0.0102441
R13826 DVDD.n6506 DVDD.n2079 0.0102441
R13827 DVDD.n9082 DVDD.n522 0.0102441
R13828 DVDD.n6018 DVDD.n3961 0.0102441
R13829 DVDD.n6061 DVDD.n5931 0.0102441
R13830 DVDD.n3244 DVDD.n3229 0.0102441
R13831 DVDD.n3269 DVDD.n2124 0.0102441
R13832 DVDD.n4925 DVDD.n486 0.0102441
R13833 DVDD.n5785 DVDD.n4308 0.0102441
R13834 DVDD.n5772 DVDD.n5766 0.0102441
R13835 DVDD.n3135 DVDD.n3118 0.0102441
R13836 DVDD.n3160 DVDD.n2176 0.0102441
R13837 DVDD.n9259 DVDD.n462 0.0102441
R13838 DVDD.n2845 DVDD.n2823 0.0102441
R13839 DVDD.n6866 DVDD.n2797 0.0102441
R13840 DVDD.n2675 DVDD.n2668 0.0102441
R13841 DVDD.n2690 DVDD.n2644 0.0102441
R13842 DVDD.n4878 DVDD.n4876 0.01022
R13843 DVDD.n4876 DVDD.n4870 0.01022
R13844 DVDD.n5026 DVDD.n4870 0.01022
R13845 DVDD.n5026 DVDD.n5025 0.01022
R13846 DVDD.n5025 DVDD.n5023 0.01022
R13847 DVDD.n5023 DVDD.n5021 0.01022
R13848 DVDD.n5021 DVDD.n5019 0.01022
R13849 DVDD.n5019 DVDD.n5017 0.01022
R13850 DVDD.n5017 DVDD.n5015 0.01022
R13851 DVDD.n5015 DVDD.n5012 0.01022
R13852 DVDD.n5012 DVDD.n5011 0.01022
R13853 DVDD.n5011 DVDD.n5009 0.01022
R13854 DVDD.n5009 DVDD.n4871 0.01022
R13855 DVDD.n5005 DVDD.n4871 0.01022
R13856 DVDD.n5005 DVDD.n5004 0.01022
R13857 DVDD.n5004 DVDD.n5003 0.01022
R13858 DVDD.n5003 DVDD.n4873 0.01022
R13859 DVDD.n4999 DVDD.n4873 0.01022
R13860 DVDD.n4999 DVDD.n4998 0.01022
R13861 DVDD.n4998 DVDD.n4997 0.01022
R13862 DVDD.n4994 DVDD.n4993 0.01022
R13863 DVDD.n4993 DVDD.n4992 0.01022
R13864 DVDD.n4992 DVDD.n4882 0.01022
R13865 DVDD.n4988 DVDD.n4882 0.01022
R13866 DVDD.n4988 DVDD.n4987 0.01022
R13867 DVDD.n4987 DVDD.n4986 0.01022
R13868 DVDD.n4986 DVDD.n4884 0.01022
R13869 DVDD.n4982 DVDD.n4884 0.01022
R13870 DVDD.n4982 DVDD.n4981 0.01022
R13871 DVDD.n4981 DVDD.n4980 0.01022
R13872 DVDD.n4980 DVDD.n4886 0.01022
R13873 DVDD.n4976 DVDD.n4886 0.01022
R13874 DVDD.n4976 DVDD.n4975 0.01022
R13875 DVDD.n4975 DVDD.n4974 0.01022
R13876 DVDD.n4974 DVDD.n4888 0.01022
R13877 DVDD.n4970 DVDD.n4888 0.01022
R13878 DVDD.n4970 DVDD.n4969 0.01022
R13879 DVDD.n4969 DVDD.n4968 0.01022
R13880 DVDD.n4968 DVDD.n4890 0.01022
R13881 DVDD.n4964 DVDD.n4890 0.01022
R13882 DVDD.n4964 DVDD.n4963 0.01022
R13883 DVDD.n4963 DVDD.n4962 0.01022
R13884 DVDD.n4962 DVDD.n4892 0.01022
R13885 DVDD.n4958 DVDD.n4892 0.01022
R13886 DVDD.n4958 DVDD.n4957 0.01022
R13887 DVDD.n4957 DVDD.n4956 0.01022
R13888 DVDD.n4956 DVDD.n4894 0.01022
R13889 DVDD.n4952 DVDD.n4894 0.01022
R13890 DVDD.n4949 DVDD.n4948 0.01022
R13891 DVDD.n4948 DVDD.n4947 0.01022
R13892 DVDD.n4947 DVDD.n4896 0.01022
R13893 DVDD.n4943 DVDD.n4896 0.01022
R13894 DVDD.n4943 DVDD.n4942 0.01022
R13895 DVDD.n4942 DVDD.n4941 0.01022
R13896 DVDD.n4941 DVDD.n4898 0.01022
R13897 DVDD.n4937 DVDD.n4898 0.01022
R13898 DVDD.n4937 DVDD.n4936 0.01022
R13899 DVDD.n4936 DVDD.n4934 0.01022
R13900 DVDD.n4934 DVDD.n4931 0.01022
R13901 DVDD.n4931 DVDD.n4930 0.01022
R13902 DVDD.n4930 DVDD.n4928 0.01022
R13903 DVDD.n4928 DVDD.n4926 0.01022
R13904 DVDD.n4926 DVDD.n4924 0.01022
R13905 DVDD.n4924 DVDD.n4922 0.01022
R13906 DVDD.n4922 DVDD.n4920 0.01022
R13907 DVDD.n4920 DVDD.n4918 0.01022
R13908 DVDD.n4918 DVDD.n4915 0.01022
R13909 DVDD.n4915 DVDD.n4914 0.01022
R13910 DVDD.n4914 DVDD.n4913 0.01022
R13911 DVDD.n4913 DVDD.n4912 0.01022
R13912 DVDD.n4912 DVDD.n4899 0.01022
R13913 DVDD.n4908 DVDD.n4899 0.01022
R13914 DVDD.n4908 DVDD.n4907 0.01022
R13915 DVDD.n4907 DVDD.n4906 0.01022
R13916 DVDD.n4906 DVDD.n4903 0.01022
R13917 DVDD.n4903 DVDD.n4902 0.01022
R13918 DVDD.n9475 DVDD.n286 0.01022
R13919 DVDD.n298 DVDD.n286 0.01022
R13920 DVDD.n299 DVDD.n298 0.01022
R13921 DVDD.n304 DVDD.n299 0.01022
R13922 DVDD.n305 DVDD.n304 0.01022
R13923 DVDD.n9463 DVDD.n305 0.01022
R13924 DVDD.n9463 DVDD.n9462 0.01022
R13925 DVDD.n9462 DVDD.n9460 0.01022
R13926 DVDD.n9460 DVDD.n306 0.01022
R13927 DVDD.n318 DVDD.n306 0.01022
R13928 DVDD.n319 DVDD.n318 0.01022
R13929 DVDD.n9449 DVDD.n319 0.01022
R13930 DVDD.n9449 DVDD.n9448 0.01022
R13931 DVDD.n9448 DVDD.n320 0.01022
R13932 DVDD.n334 DVDD.n320 0.01022
R13933 DVDD.n334 DVDD.n333 0.01022
R13934 DVDD.n341 DVDD.n333 0.01022
R13935 DVDD.n342 DVDD.n341 0.01022
R13936 DVDD.n9436 DVDD.n342 0.01022
R13937 DVDD.n9436 DVDD.n9435 0.01022
R13938 DVDD.n9435 DVDD.n9434 0.01022
R13939 DVDD.n9434 DVDD.n343 0.01022
R13940 DVDD.n368 DVDD.n343 0.01022
R13941 DVDD.n368 DVDD.n367 0.01022
R13942 DVDD.n367 DVDD.n285 0.01022
R13943 DVDD.n9480 DVDD.n285 0.01022
R13944 DVDD.n9480 DVDD.n9479 0.01022
R13945 DVDD.n9479 DVDD.n9477 0.01022
R13946 DVDD.n9511 DVDD.n266 0.01022
R13947 DVDD.n266 DVDD.n247 0.01022
R13948 DVDD.n9553 DVDD.n247 0.01022
R13949 DVDD.n9553 DVDD.n9552 0.01022
R13950 DVDD.n9552 DVDD.n9551 0.01022
R13951 DVDD.n9551 DVDD.n248 0.01022
R13952 DVDD.n9544 DVDD.n248 0.01022
R13953 DVDD.n9544 DVDD.n9543 0.01022
R13954 DVDD.n9543 DVDD.n9542 0.01022
R13955 DVDD.n9542 DVDD.n256 0.01022
R13956 DVDD.n9538 DVDD.n256 0.01022
R13957 DVDD.n9538 DVDD.n9537 0.01022
R13958 DVDD.n9537 DVDD.n9536 0.01022
R13959 DVDD.n9536 DVDD.n258 0.01022
R13960 DVDD.n9532 DVDD.n258 0.01022
R13961 DVDD.n9532 DVDD.n9531 0.01022
R13962 DVDD.n9531 DVDD.n9530 0.01022
R13963 DVDD.n9530 DVDD.n260 0.01022
R13964 DVDD.n9526 DVDD.n260 0.01022
R13965 DVDD.n9526 DVDD.n9525 0.01022
R13966 DVDD.n9525 DVDD.n9524 0.01022
R13967 DVDD.n9524 DVDD.n262 0.01022
R13968 DVDD.n9520 DVDD.n262 0.01022
R13969 DVDD.n9520 DVDD.n9519 0.01022
R13970 DVDD.n9519 DVDD.n9518 0.01022
R13971 DVDD.n9518 DVDD.n264 0.01022
R13972 DVDD.n9514 DVDD.n264 0.01022
R13973 DVDD.n9514 DVDD.n9513 0.01022
R13974 DVDD.n4372 DVDD.n4319 0.01022
R13975 DVDD.n4368 DVDD.n4319 0.01022
R13976 DVDD.n4368 DVDD.n4367 0.01022
R13977 DVDD.n4367 DVDD.n4366 0.01022
R13978 DVDD.n4366 DVDD.n4321 0.01022
R13979 DVDD.n4362 DVDD.n4321 0.01022
R13980 DVDD.n4362 DVDD.n4361 0.01022
R13981 DVDD.n4361 DVDD.n4360 0.01022
R13982 DVDD.n4360 DVDD.n4323 0.01022
R13983 DVDD.n4356 DVDD.n4323 0.01022
R13984 DVDD.n4356 DVDD.n4355 0.01022
R13985 DVDD.n4355 DVDD.n4354 0.01022
R13986 DVDD.n4354 DVDD.n4325 0.01022
R13987 DVDD.n4350 DVDD.n4325 0.01022
R13988 DVDD.n4350 DVDD.n4349 0.01022
R13989 DVDD.n4349 DVDD.n4348 0.01022
R13990 DVDD.n4348 DVDD.n4327 0.01022
R13991 DVDD.n4344 DVDD.n4327 0.01022
R13992 DVDD.n4344 DVDD.n4343 0.01022
R13993 DVDD.n4343 DVDD.n4342 0.01022
R13994 DVDD.n4342 DVDD.n4329 0.01022
R13995 DVDD.n4338 DVDD.n4329 0.01022
R13996 DVDD.n4338 DVDD.n4337 0.01022
R13997 DVDD.n4337 DVDD.n4336 0.01022
R13998 DVDD.n4336 DVDD.n4331 0.01022
R13999 DVDD.n4332 DVDD.n4331 0.01022
R14000 DVDD.n4332 DVDD.n4318 0.01022
R14001 DVDD.n4374 DVDD.n4318 0.01022
R14002 DVDD.n5820 DVDD.n5818 0.01022
R14003 DVDD.n5818 DVDD.n5816 0.01022
R14004 DVDD.n5816 DVDD.n5814 0.01022
R14005 DVDD.n5814 DVDD.n5812 0.01022
R14006 DVDD.n5812 DVDD.n5809 0.01022
R14007 DVDD.n5809 DVDD.n5808 0.01022
R14008 DVDD.n5808 DVDD.n5806 0.01022
R14009 DVDD.n5806 DVDD.n5804 0.01022
R14010 DVDD.n5804 DVDD.n5802 0.01022
R14011 DVDD.n5802 DVDD.n5800 0.01022
R14012 DVDD.n5800 DVDD.n5798 0.01022
R14013 DVDD.n5798 DVDD.n5796 0.01022
R14014 DVDD.n5796 DVDD.n5793 0.01022
R14015 DVDD.n5793 DVDD.n5792 0.01022
R14016 DVDD.n5792 DVDD.n5790 0.01022
R14017 DVDD.n5790 DVDD.n5788 0.01022
R14018 DVDD.n5788 DVDD.n5786 0.01022
R14019 DVDD.n5786 DVDD.n5784 0.01022
R14020 DVDD.n5784 DVDD.n5782 0.01022
R14021 DVDD.n5782 DVDD.n5780 0.01022
R14022 DVDD.n5780 DVDD.n5777 0.01022
R14023 DVDD.n5777 DVDD.n5776 0.01022
R14024 DVDD.n5776 DVDD.n5775 0.01022
R14025 DVDD.n5775 DVDD.n5774 0.01022
R14026 DVDD.n5774 DVDD.n5771 0.01022
R14027 DVDD.n5771 DVDD.n5770 0.01022
R14028 DVDD.n5770 DVDD.n5768 0.01022
R14029 DVDD.n5822 DVDD.n5768 0.01022
R14030 DVDD.n5886 DVDD.n5831 0.01022
R14031 DVDD.n5886 DVDD.n5885 0.01022
R14032 DVDD.n5885 DVDD.n5884 0.01022
R14033 DVDD.n5884 DVDD.n5832 0.01022
R14034 DVDD.n5880 DVDD.n5832 0.01022
R14035 DVDD.n5880 DVDD.n5879 0.01022
R14036 DVDD.n5879 DVDD.n5878 0.01022
R14037 DVDD.n5878 DVDD.n5834 0.01022
R14038 DVDD.n5874 DVDD.n5834 0.01022
R14039 DVDD.n5874 DVDD.n5873 0.01022
R14040 DVDD.n5873 DVDD.n5872 0.01022
R14041 DVDD.n5872 DVDD.n5836 0.01022
R14042 DVDD.n5868 DVDD.n5836 0.01022
R14043 DVDD.n5868 DVDD.n5867 0.01022
R14044 DVDD.n5867 DVDD.n5866 0.01022
R14045 DVDD.n5866 DVDD.n5838 0.01022
R14046 DVDD.n5862 DVDD.n5838 0.01022
R14047 DVDD.n5862 DVDD.n5861 0.01022
R14048 DVDD.n5861 DVDD.n5860 0.01022
R14049 DVDD.n5860 DVDD.n5858 0.01022
R14050 DVDD.n5858 DVDD.n5856 0.01022
R14051 DVDD.n5856 DVDD.n5854 0.01022
R14052 DVDD.n5854 DVDD.n5851 0.01022
R14053 DVDD.n5851 DVDD.n5850 0.01022
R14054 DVDD.n5850 DVDD.n5848 0.01022
R14055 DVDD.n5848 DVDD.n5846 0.01022
R14056 DVDD.n5846 DVDD.n5844 0.01022
R14057 DVDD.n5844 DVDD.n5842 0.01022
R14058 DVDD.n3140 DVDD.n3138 0.01022
R14059 DVDD.n3138 DVDD.n3136 0.01022
R14060 DVDD.n3136 DVDD.n3134 0.01022
R14061 DVDD.n3134 DVDD.n3132 0.01022
R14062 DVDD.n3132 DVDD.n3130 0.01022
R14063 DVDD.n3130 DVDD.n3127 0.01022
R14064 DVDD.n3127 DVDD.n3126 0.01022
R14065 DVDD.n3126 DVDD.n3124 0.01022
R14066 DVDD.n3179 DVDD.n3124 0.01022
R14067 DVDD.n3179 DVDD.n3178 0.01022
R14068 DVDD.n3178 DVDD.n3177 0.01022
R14069 DVDD.n3177 DVDD.n3175 0.01022
R14070 DVDD.n3175 DVDD.n3173 0.01022
R14071 DVDD.n3173 DVDD.n3171 0.01022
R14072 DVDD.n3171 DVDD.n3168 0.01022
R14073 DVDD.n3168 DVDD.n3167 0.01022
R14074 DVDD.n3167 DVDD.n3165 0.01022
R14075 DVDD.n3165 DVDD.n3163 0.01022
R14076 DVDD.n3163 DVDD.n3161 0.01022
R14077 DVDD.n3161 DVDD.n3159 0.01022
R14078 DVDD.n3159 DVDD.n3157 0.01022
R14079 DVDD.n3157 DVDD.n3155 0.01022
R14080 DVDD.n3155 DVDD.n3152 0.01022
R14081 DVDD.n3152 DVDD.n3151 0.01022
R14082 DVDD.n3151 DVDD.n3149 0.01022
R14083 DVDD.n3149 DVDD.n3147 0.01022
R14084 DVDD.n3147 DVDD.n3145 0.01022
R14085 DVDD.n3145 DVDD.n3143 0.01022
R14086 DVDD.n8977 DVDD.n547 0.01022
R14087 DVDD.n8980 DVDD.n8977 0.01022
R14088 DVDD.n8982 DVDD.n8980 0.01022
R14089 DVDD.n8984 DVDD.n8982 0.01022
R14090 DVDD.n8986 DVDD.n8984 0.01022
R14091 DVDD.n8988 DVDD.n8986 0.01022
R14092 DVDD.n8989 DVDD.n8988 0.01022
R14093 DVDD.n9010 DVDD.n8989 0.01022
R14094 DVDD.n9010 DVDD.n9009 0.01022
R14095 DVDD.n9009 DVDD.n9006 0.01022
R14096 DVDD.n9006 DVDD.n9005 0.01022
R14097 DVDD.n9005 DVDD.n9003 0.01022
R14098 DVDD.n9003 DVDD.n8990 0.01022
R14099 DVDD.n8999 DVDD.n8990 0.01022
R14100 DVDD.n8999 DVDD.n8998 0.01022
R14101 DVDD.n8998 DVDD.n8997 0.01022
R14102 DVDD.n8997 DVDD.n8992 0.01022
R14103 DVDD.n8993 DVDD.n8992 0.01022
R14104 DVDD.n8993 DVDD.n546 0.01022
R14105 DVDD.n9017 DVDD.n546 0.01022
R14106 DVDD.n9071 DVDD.n544 0.01022
R14107 DVDD.n9067 DVDD.n544 0.01022
R14108 DVDD.n9067 DVDD.n9066 0.01022
R14109 DVDD.n9066 DVDD.n9065 0.01022
R14110 DVDD.n9065 DVDD.n9020 0.01022
R14111 DVDD.n9061 DVDD.n9020 0.01022
R14112 DVDD.n9061 DVDD.n9060 0.01022
R14113 DVDD.n9060 DVDD.n9059 0.01022
R14114 DVDD.n9059 DVDD.n9022 0.01022
R14115 DVDD.n9055 DVDD.n9022 0.01022
R14116 DVDD.n9055 DVDD.n9054 0.01022
R14117 DVDD.n9054 DVDD.n9053 0.01022
R14118 DVDD.n9053 DVDD.n9024 0.01022
R14119 DVDD.n9049 DVDD.n9024 0.01022
R14120 DVDD.n9049 DVDD.n9048 0.01022
R14121 DVDD.n9048 DVDD.n9047 0.01022
R14122 DVDD.n9047 DVDD.n9026 0.01022
R14123 DVDD.n9043 DVDD.n9026 0.01022
R14124 DVDD.n9043 DVDD.n9042 0.01022
R14125 DVDD.n9042 DVDD.n9041 0.01022
R14126 DVDD.n9041 DVDD.n9028 0.01022
R14127 DVDD.n9037 DVDD.n9028 0.01022
R14128 DVDD.n9037 DVDD.n9036 0.01022
R14129 DVDD.n9036 DVDD.n9035 0.01022
R14130 DVDD.n9035 DVDD.n9030 0.01022
R14131 DVDD.n9031 DVDD.n9030 0.01022
R14132 DVDD.n9031 DVDD.n543 0.01022
R14133 DVDD.n9073 DVDD.n543 0.01022
R14134 DVDD.n9107 DVDD.n541 0.01022
R14135 DVDD.n9103 DVDD.n541 0.01022
R14136 DVDD.n9103 DVDD.n9102 0.01022
R14137 DVDD.n9102 DVDD.n9101 0.01022
R14138 DVDD.n9101 DVDD.n9076 0.01022
R14139 DVDD.n9097 DVDD.n9076 0.01022
R14140 DVDD.n9097 DVDD.n9096 0.01022
R14141 DVDD.n9096 DVDD.n9095 0.01022
R14142 DVDD.n9095 DVDD.n9093 0.01022
R14143 DVDD.n9093 DVDD.n9091 0.01022
R14144 DVDD.n9091 DVDD.n9088 0.01022
R14145 DVDD.n9088 DVDD.n9087 0.01022
R14146 DVDD.n9087 DVDD.n9085 0.01022
R14147 DVDD.n9085 DVDD.n9083 0.01022
R14148 DVDD.n9083 DVDD.n9081 0.01022
R14149 DVDD.n9081 DVDD.n9079 0.01022
R14150 DVDD.n9079 DVDD.n536 0.01022
R14151 DVDD.n9124 DVDD.n536 0.01022
R14152 DVDD.n9124 DVDD.n9123 0.01022
R14153 DVDD.n9123 DVDD.n9122 0.01022
R14154 DVDD.n9122 DVDD.n9120 0.01022
R14155 DVDD.n9120 DVDD.n537 0.01022
R14156 DVDD.n9116 DVDD.n537 0.01022
R14157 DVDD.n9116 DVDD.n9115 0.01022
R14158 DVDD.n9115 DVDD.n9114 0.01022
R14159 DVDD.n9114 DVDD.n539 0.01022
R14160 DVDD.n9110 DVDD.n539 0.01022
R14161 DVDD.n9110 DVDD.n9109 0.01022
R14162 DVDD.n4115 DVDD.n3996 0.01022
R14163 DVDD.n4005 DVDD.n3996 0.01022
R14164 DVDD.n4006 DVDD.n4005 0.01022
R14165 DVDD.n4006 DVDD.n4003 0.01022
R14166 DVDD.n4013 DVDD.n4003 0.01022
R14167 DVDD.n4014 DVDD.n4013 0.01022
R14168 DVDD.n4099 DVDD.n4014 0.01022
R14169 DVDD.n4099 DVDD.n4098 0.01022
R14170 DVDD.n4098 DVDD.n4015 0.01022
R14171 DVDD.n4038 DVDD.n4015 0.01022
R14172 DVDD.n4039 DVDD.n4038 0.01022
R14173 DVDD.n4039 DVDD.n4035 0.01022
R14174 DVDD.n4049 DVDD.n4035 0.01022
R14175 DVDD.n4050 DVDD.n4049 0.01022
R14176 DVDD.n4050 DVDD.n4033 0.01022
R14177 DVDD.n4054 DVDD.n4033 0.01022
R14178 DVDD.n4056 DVDD.n4054 0.01022
R14179 DVDD.n4056 DVDD.n4055 0.01022
R14180 DVDD.n4055 DVDD.n4029 0.01022
R14181 DVDD.n4066 DVDD.n4029 0.01022
R14182 DVDD.n4067 DVDD.n4066 0.01022
R14183 DVDD.n4076 DVDD.n4067 0.01022
R14184 DVDD.n4076 DVDD.n4075 0.01022
R14185 DVDD.n4075 DVDD.n4068 0.01022
R14186 DVDD.n4068 DVDD.n3995 0.01022
R14187 DVDD.n4120 DVDD.n3995 0.01022
R14188 DVDD.n4120 DVDD.n4119 0.01022
R14189 DVDD.n4119 DVDD.n4117 0.01022
R14190 DVDD.n4220 DVDD.n3975 0.01022
R14191 DVDD.n4156 DVDD.n3975 0.01022
R14192 DVDD.n4157 DVDD.n4156 0.01022
R14193 DVDD.n4162 DVDD.n4157 0.01022
R14194 DVDD.n4163 DVDD.n4162 0.01022
R14195 DVDD.n4204 DVDD.n4163 0.01022
R14196 DVDD.n4204 DVDD.n4203 0.01022
R14197 DVDD.n4203 DVDD.n4164 0.01022
R14198 DVDD.n4199 DVDD.n4164 0.01022
R14199 DVDD.n4199 DVDD.n4198 0.01022
R14200 DVDD.n4198 DVDD.n4197 0.01022
R14201 DVDD.n4197 DVDD.n4166 0.01022
R14202 DVDD.n4193 DVDD.n4166 0.01022
R14203 DVDD.n4193 DVDD.n4192 0.01022
R14204 DVDD.n4192 DVDD.n4191 0.01022
R14205 DVDD.n4191 DVDD.n4168 0.01022
R14206 DVDD.n4187 DVDD.n4168 0.01022
R14207 DVDD.n4187 DVDD.n4186 0.01022
R14208 DVDD.n4186 DVDD.n4185 0.01022
R14209 DVDD.n4185 DVDD.n4170 0.01022
R14210 DVDD.n4181 DVDD.n4170 0.01022
R14211 DVDD.n4181 DVDD.n4180 0.01022
R14212 DVDD.n4180 DVDD.n4179 0.01022
R14213 DVDD.n4179 DVDD.n4172 0.01022
R14214 DVDD.n4175 DVDD.n4172 0.01022
R14215 DVDD.n4175 DVDD.n4174 0.01022
R14216 DVDD.n4174 DVDD.n3974 0.01022
R14217 DVDD.n4222 DVDD.n3974 0.01022
R14218 DVDD.n4276 DVDD.n3972 0.01022
R14219 DVDD.n4272 DVDD.n3972 0.01022
R14220 DVDD.n4272 DVDD.n4271 0.01022
R14221 DVDD.n4271 DVDD.n4270 0.01022
R14222 DVDD.n4270 DVDD.n4225 0.01022
R14223 DVDD.n4266 DVDD.n4225 0.01022
R14224 DVDD.n4266 DVDD.n4265 0.01022
R14225 DVDD.n4265 DVDD.n4264 0.01022
R14226 DVDD.n4264 DVDD.n4227 0.01022
R14227 DVDD.n4260 DVDD.n4227 0.01022
R14228 DVDD.n4260 DVDD.n4259 0.01022
R14229 DVDD.n4259 DVDD.n4258 0.01022
R14230 DVDD.n4258 DVDD.n4229 0.01022
R14231 DVDD.n4254 DVDD.n4229 0.01022
R14232 DVDD.n4254 DVDD.n4253 0.01022
R14233 DVDD.n4253 DVDD.n4252 0.01022
R14234 DVDD.n4252 DVDD.n4231 0.01022
R14235 DVDD.n4248 DVDD.n4231 0.01022
R14236 DVDD.n4248 DVDD.n4247 0.01022
R14237 DVDD.n4247 DVDD.n4246 0.01022
R14238 DVDD.n4246 DVDD.n4233 0.01022
R14239 DVDD.n4242 DVDD.n4233 0.01022
R14240 DVDD.n4242 DVDD.n4241 0.01022
R14241 DVDD.n4241 DVDD.n4240 0.01022
R14242 DVDD.n4240 DVDD.n4235 0.01022
R14243 DVDD.n4236 DVDD.n4235 0.01022
R14244 DVDD.n4236 DVDD.n3971 0.01022
R14245 DVDD.n4278 DVDD.n3971 0.01022
R14246 DVDD.n6053 DVDD.n6051 0.01022
R14247 DVDD.n6051 DVDD.n6049 0.01022
R14248 DVDD.n6049 DVDD.n6047 0.01022
R14249 DVDD.n6047 DVDD.n6045 0.01022
R14250 DVDD.n6045 DVDD.n6042 0.01022
R14251 DVDD.n6042 DVDD.n6041 0.01022
R14252 DVDD.n6041 DVDD.n6039 0.01022
R14253 DVDD.n6039 DVDD.n6037 0.01022
R14254 DVDD.n6037 DVDD.n6035 0.01022
R14255 DVDD.n6035 DVDD.n6033 0.01022
R14256 DVDD.n6033 DVDD.n6031 0.01022
R14257 DVDD.n6031 DVDD.n6029 0.01022
R14258 DVDD.n6029 DVDD.n6026 0.01022
R14259 DVDD.n6026 DVDD.n6025 0.01022
R14260 DVDD.n6025 DVDD.n6023 0.01022
R14261 DVDD.n6023 DVDD.n6021 0.01022
R14262 DVDD.n6021 DVDD.n6019 0.01022
R14263 DVDD.n6019 DVDD.n6017 0.01022
R14264 DVDD.n6017 DVDD.n6015 0.01022
R14265 DVDD.n6015 DVDD.n6013 0.01022
R14266 DVDD.n6013 DVDD.n6010 0.01022
R14267 DVDD.n6010 DVDD.n6009 0.01022
R14268 DVDD.n6009 DVDD.n6007 0.01022
R14269 DVDD.n6007 DVDD.n6004 0.01022
R14270 DVDD.n6004 DVDD.n6003 0.01022
R14271 DVDD.n6059 DVDD.n6003 0.01022
R14272 DVDD.n6059 DVDD.n6058 0.01022
R14273 DVDD.n6058 DVDD.n6056 0.01022
R14274 DVDD.n5991 DVDD.n5990 0.01022
R14275 DVDD.n5990 DVDD.n5934 0.01022
R14276 DVDD.n5986 DVDD.n5934 0.01022
R14277 DVDD.n5986 DVDD.n5985 0.01022
R14278 DVDD.n5985 DVDD.n5984 0.01022
R14279 DVDD.n5984 DVDD.n5936 0.01022
R14280 DVDD.n5980 DVDD.n5936 0.01022
R14281 DVDD.n5980 DVDD.n5979 0.01022
R14282 DVDD.n5979 DVDD.n5978 0.01022
R14283 DVDD.n5978 DVDD.n5938 0.01022
R14284 DVDD.n5974 DVDD.n5938 0.01022
R14285 DVDD.n5974 DVDD.n5973 0.01022
R14286 DVDD.n5973 DVDD.n5972 0.01022
R14287 DVDD.n5972 DVDD.n5940 0.01022
R14288 DVDD.n5968 DVDD.n5940 0.01022
R14289 DVDD.n5968 DVDD.n5967 0.01022
R14290 DVDD.n5967 DVDD.n5966 0.01022
R14291 DVDD.n5966 DVDD.n5963 0.01022
R14292 DVDD.n5963 DVDD.n5962 0.01022
R14293 DVDD.n5962 DVDD.n5960 0.01022
R14294 DVDD.n5960 DVDD.n5958 0.01022
R14295 DVDD.n5958 DVDD.n5956 0.01022
R14296 DVDD.n5956 DVDD.n5953 0.01022
R14297 DVDD.n5953 DVDD.n5952 0.01022
R14298 DVDD.n5952 DVDD.n5950 0.01022
R14299 DVDD.n5950 DVDD.n5948 0.01022
R14300 DVDD.n5948 DVDD.n5946 0.01022
R14301 DVDD.n5946 DVDD.n5944 0.01022
R14302 DVDD.n3249 DVDD.n3247 0.01022
R14303 DVDD.n3247 DVDD.n3245 0.01022
R14304 DVDD.n3245 DVDD.n3243 0.01022
R14305 DVDD.n3243 DVDD.n3240 0.01022
R14306 DVDD.n3295 DVDD.n3240 0.01022
R14307 DVDD.n3295 DVDD.n3294 0.01022
R14308 DVDD.n3294 DVDD.n3293 0.01022
R14309 DVDD.n3293 DVDD.n3291 0.01022
R14310 DVDD.n3291 DVDD.n3289 0.01022
R14311 DVDD.n3289 DVDD.n3241 0.01022
R14312 DVDD.n3285 DVDD.n3241 0.01022
R14313 DVDD.n3285 DVDD.n3284 0.01022
R14314 DVDD.n3284 DVDD.n3282 0.01022
R14315 DVDD.n3282 DVDD.n3280 0.01022
R14316 DVDD.n3280 DVDD.n3277 0.01022
R14317 DVDD.n3277 DVDD.n3276 0.01022
R14318 DVDD.n3276 DVDD.n3274 0.01022
R14319 DVDD.n3274 DVDD.n3272 0.01022
R14320 DVDD.n3272 DVDD.n3270 0.01022
R14321 DVDD.n3270 DVDD.n3268 0.01022
R14322 DVDD.n3268 DVDD.n3266 0.01022
R14323 DVDD.n3266 DVDD.n3264 0.01022
R14324 DVDD.n3264 DVDD.n3261 0.01022
R14325 DVDD.n3261 DVDD.n3260 0.01022
R14326 DVDD.n3260 DVDD.n3258 0.01022
R14327 DVDD.n3258 DVDD.n3256 0.01022
R14328 DVDD.n3256 DVDD.n3254 0.01022
R14329 DVDD.n3254 DVDD.n3252 0.01022
R14330 DVDD.n5121 DVDD.n4569 0.01022
R14331 DVDD.n5124 DVDD.n5121 0.01022
R14332 DVDD.n5126 DVDD.n5124 0.01022
R14333 DVDD.n5128 DVDD.n5126 0.01022
R14334 DVDD.n5130 DVDD.n5128 0.01022
R14335 DVDD.n5132 DVDD.n5130 0.01022
R14336 DVDD.n5133 DVDD.n5132 0.01022
R14337 DVDD.n5154 DVDD.n5133 0.01022
R14338 DVDD.n5154 DVDD.n5153 0.01022
R14339 DVDD.n5153 DVDD.n5150 0.01022
R14340 DVDD.n5150 DVDD.n5149 0.01022
R14341 DVDD.n5149 DVDD.n5147 0.01022
R14342 DVDD.n5147 DVDD.n5134 0.01022
R14343 DVDD.n5143 DVDD.n5134 0.01022
R14344 DVDD.n5143 DVDD.n5142 0.01022
R14345 DVDD.n5142 DVDD.n5141 0.01022
R14346 DVDD.n5141 DVDD.n5136 0.01022
R14347 DVDD.n5137 DVDD.n5136 0.01022
R14348 DVDD.n5137 DVDD.n4566 0.01022
R14349 DVDD.n5160 DVDD.n4566 0.01022
R14350 DVDD.n5216 DVDD.n4564 0.01022
R14351 DVDD.n5212 DVDD.n4564 0.01022
R14352 DVDD.n5212 DVDD.n5211 0.01022
R14353 DVDD.n5211 DVDD.n5210 0.01022
R14354 DVDD.n5210 DVDD.n5163 0.01022
R14355 DVDD.n5206 DVDD.n5163 0.01022
R14356 DVDD.n5206 DVDD.n5205 0.01022
R14357 DVDD.n5205 DVDD.n5204 0.01022
R14358 DVDD.n5204 DVDD.n5165 0.01022
R14359 DVDD.n5200 DVDD.n5165 0.01022
R14360 DVDD.n5200 DVDD.n5199 0.01022
R14361 DVDD.n5199 DVDD.n5198 0.01022
R14362 DVDD.n5198 DVDD.n5167 0.01022
R14363 DVDD.n5194 DVDD.n5167 0.01022
R14364 DVDD.n5194 DVDD.n5193 0.01022
R14365 DVDD.n5193 DVDD.n5192 0.01022
R14366 DVDD.n5192 DVDD.n5169 0.01022
R14367 DVDD.n5188 DVDD.n5169 0.01022
R14368 DVDD.n5188 DVDD.n5187 0.01022
R14369 DVDD.n5187 DVDD.n5186 0.01022
R14370 DVDD.n5186 DVDD.n5171 0.01022
R14371 DVDD.n5182 DVDD.n5171 0.01022
R14372 DVDD.n5182 DVDD.n5181 0.01022
R14373 DVDD.n5181 DVDD.n5180 0.01022
R14374 DVDD.n5180 DVDD.n5173 0.01022
R14375 DVDD.n5176 DVDD.n5173 0.01022
R14376 DVDD.n5176 DVDD.n5175 0.01022
R14377 DVDD.n5175 DVDD.n4562 0.01022
R14378 DVDD.n9299 DVDD.n450 0.01022
R14379 DVDD.n9295 DVDD.n450 0.01022
R14380 DVDD.n9295 DVDD.n9294 0.01022
R14381 DVDD.n9294 DVDD.n9293 0.01022
R14382 DVDD.n9293 DVDD.n453 0.01022
R14383 DVDD.n9289 DVDD.n453 0.01022
R14384 DVDD.n9289 DVDD.n9288 0.01022
R14385 DVDD.n9288 DVDD.n9287 0.01022
R14386 DVDD.n9287 DVDD.n455 0.01022
R14387 DVDD.n9251 DVDD.n455 0.01022
R14388 DVDD.n9254 DVDD.n9251 0.01022
R14389 DVDD.n9256 DVDD.n9254 0.01022
R14390 DVDD.n9258 DVDD.n9256 0.01022
R14391 DVDD.n9260 DVDD.n9258 0.01022
R14392 DVDD.n9262 DVDD.n9260 0.01022
R14393 DVDD.n9264 DVDD.n9262 0.01022
R14394 DVDD.n9265 DVDD.n9264 0.01022
R14395 DVDD.n9281 DVDD.n9265 0.01022
R14396 DVDD.n9281 DVDD.n9280 0.01022
R14397 DVDD.n9280 DVDD.n9279 0.01022
R14398 DVDD.n9279 DVDD.n9277 0.01022
R14399 DVDD.n9277 DVDD.n9266 0.01022
R14400 DVDD.n9273 DVDD.n9266 0.01022
R14401 DVDD.n9273 DVDD.n9272 0.01022
R14402 DVDD.n9272 DVDD.n9271 0.01022
R14403 DVDD.n9271 DVDD.n9268 0.01022
R14404 DVDD.n9268 DVDD.n447 0.01022
R14405 DVDD.n9300 DVDD.n447 0.01022
R14406 DVDD.n9304 DVDD.n445 0.01022
R14407 DVDD.n9305 DVDD.n9304 0.01022
R14408 DVDD.n9306 DVDD.n9305 0.01022
R14409 DVDD.n9307 DVDD.n9306 0.01022
R14410 DVDD.n9310 DVDD.n9307 0.01022
R14411 DVDD.n9310 DVDD.n9309 0.01022
R14412 DVDD.n9309 DVDD.n9308 0.01022
R14413 DVDD.n9308 DVDD.n134 0.01022
R14414 DVDD.n9610 DVDD.n134 0.01022
R14415 DVDD.n9610 DVDD.n9609 0.01022
R14416 DVDD.n9609 DVDD.n135 0.01022
R14417 DVDD.n157 DVDD.n135 0.01022
R14418 DVDD.n158 DVDD.n157 0.01022
R14419 DVDD.n159 DVDD.n158 0.01022
R14420 DVDD.n161 DVDD.n159 0.01022
R14421 DVDD.n162 DVDD.n161 0.01022
R14422 DVDD.n9593 DVDD.n162 0.01022
R14423 DVDD.n9593 DVDD.n9592 0.01022
R14424 DVDD.n9592 DVDD.n163 0.01022
R14425 DVDD.n402 DVDD.n163 0.01022
R14426 DVDD.n403 DVDD.n402 0.01022
R14427 DVDD.n9394 DVDD.n403 0.01022
R14428 DVDD.n9395 DVDD.n9394 0.01022
R14429 DVDD.n9396 DVDD.n9395 0.01022
R14430 DVDD.n9396 DVDD.n390 0.01022
R14431 DVDD.n9412 DVDD.n390 0.01022
R14432 DVDD.n9412 DVDD.n9411 0.01022
R14433 DVDD.n9411 DVDD.n391 0.01022
R14434 DVDD.n6796 DVDD.n2888 0.01022
R14435 DVDD.n2902 DVDD.n2888 0.01022
R14436 DVDD.n6785 DVDD.n2902 0.01022
R14437 DVDD.n6785 DVDD.n6784 0.01022
R14438 DVDD.n6784 DVDD.n6783 0.01022
R14439 DVDD.n6783 DVDD.n2903 0.01022
R14440 DVDD.n2955 DVDD.n2903 0.01022
R14441 DVDD.n2955 DVDD.n2954 0.01022
R14442 DVDD.n2954 DVDD.n2953 0.01022
R14443 DVDD.n2953 DVDD.n2918 0.01022
R14444 DVDD.n2949 DVDD.n2918 0.01022
R14445 DVDD.n2949 DVDD.n2948 0.01022
R14446 DVDD.n2948 DVDD.n2947 0.01022
R14447 DVDD.n2947 DVDD.n2920 0.01022
R14448 DVDD.n2943 DVDD.n2920 0.01022
R14449 DVDD.n2943 DVDD.n2942 0.01022
R14450 DVDD.n2942 DVDD.n2941 0.01022
R14451 DVDD.n2941 DVDD.n2922 0.01022
R14452 DVDD.n2937 DVDD.n2922 0.01022
R14453 DVDD.n2937 DVDD.n2936 0.01022
R14454 DVDD.n2936 DVDD.n2935 0.01022
R14455 DVDD.n2935 DVDD.n2924 0.01022
R14456 DVDD.n2931 DVDD.n2924 0.01022
R14457 DVDD.n2931 DVDD.n2930 0.01022
R14458 DVDD.n2930 DVDD.n2929 0.01022
R14459 DVDD.n2929 DVDD.n2926 0.01022
R14460 DVDD.n2926 DVDD.n2885 0.01022
R14461 DVDD.n6797 DVDD.n2885 0.01022
R14462 DVDD.n6851 DVDD.n2883 0.01022
R14463 DVDD.n6847 DVDD.n2883 0.01022
R14464 DVDD.n6847 DVDD.n6846 0.01022
R14465 DVDD.n6846 DVDD.n6845 0.01022
R14466 DVDD.n6845 DVDD.n6800 0.01022
R14467 DVDD.n6841 DVDD.n6800 0.01022
R14468 DVDD.n6841 DVDD.n6840 0.01022
R14469 DVDD.n6840 DVDD.n6839 0.01022
R14470 DVDD.n6839 DVDD.n6802 0.01022
R14471 DVDD.n6835 DVDD.n6802 0.01022
R14472 DVDD.n6835 DVDD.n6834 0.01022
R14473 DVDD.n6834 DVDD.n6833 0.01022
R14474 DVDD.n6833 DVDD.n6804 0.01022
R14475 DVDD.n6829 DVDD.n6804 0.01022
R14476 DVDD.n6829 DVDD.n6828 0.01022
R14477 DVDD.n6828 DVDD.n6827 0.01022
R14478 DVDD.n6827 DVDD.n6806 0.01022
R14479 DVDD.n6823 DVDD.n6806 0.01022
R14480 DVDD.n6823 DVDD.n6822 0.01022
R14481 DVDD.n6822 DVDD.n6821 0.01022
R14482 DVDD.n6821 DVDD.n6808 0.01022
R14483 DVDD.n6817 DVDD.n6808 0.01022
R14484 DVDD.n6817 DVDD.n6816 0.01022
R14485 DVDD.n6816 DVDD.n6815 0.01022
R14486 DVDD.n6815 DVDD.n6810 0.01022
R14487 DVDD.n6811 DVDD.n6810 0.01022
R14488 DVDD.n6811 DVDD.n2880 0.01022
R14489 DVDD.n6852 DVDD.n2880 0.01022
R14490 DVDD.n6859 DVDD.n2802 0.01022
R14491 DVDD.n2830 DVDD.n2802 0.01022
R14492 DVDD.n2873 DVDD.n2830 0.01022
R14493 DVDD.n2873 DVDD.n2872 0.01022
R14494 DVDD.n2872 DVDD.n2869 0.01022
R14495 DVDD.n2869 DVDD.n2868 0.01022
R14496 DVDD.n2868 DVDD.n2866 0.01022
R14497 DVDD.n2866 DVDD.n2864 0.01022
R14498 DVDD.n2864 DVDD.n2862 0.01022
R14499 DVDD.n2862 DVDD.n2860 0.01022
R14500 DVDD.n2860 DVDD.n2858 0.01022
R14501 DVDD.n2858 DVDD.n2856 0.01022
R14502 DVDD.n2856 DVDD.n2853 0.01022
R14503 DVDD.n2853 DVDD.n2852 0.01022
R14504 DVDD.n2852 DVDD.n2850 0.01022
R14505 DVDD.n2850 DVDD.n2848 0.01022
R14506 DVDD.n2848 DVDD.n2846 0.01022
R14507 DVDD.n2846 DVDD.n2844 0.01022
R14508 DVDD.n2844 DVDD.n2842 0.01022
R14509 DVDD.n2842 DVDD.n2840 0.01022
R14510 DVDD.n2840 DVDD.n2837 0.01022
R14511 DVDD.n2837 DVDD.n2836 0.01022
R14512 DVDD.n2836 DVDD.n2834 0.01022
R14513 DVDD.n2834 DVDD.n2831 0.01022
R14514 DVDD.n2831 DVDD.n2799 0.01022
R14515 DVDD.n6864 DVDD.n2799 0.01022
R14516 DVDD.n6864 DVDD.n6863 0.01022
R14517 DVDD.n6863 DVDD.n6860 0.01022
R14518 DVDD.n6902 DVDD.n2741 0.01022
R14519 DVDD.n2774 DVDD.n2741 0.01022
R14520 DVDD.n2774 DVDD.n2773 0.01022
R14521 DVDD.n2773 DVDD.n2772 0.01022
R14522 DVDD.n2772 DVDD.n2745 0.01022
R14523 DVDD.n2768 DVDD.n2745 0.01022
R14524 DVDD.n2768 DVDD.n2767 0.01022
R14525 DVDD.n2767 DVDD.n2766 0.01022
R14526 DVDD.n2766 DVDD.n2747 0.01022
R14527 DVDD.n2762 DVDD.n2747 0.01022
R14528 DVDD.n2762 DVDD.n2761 0.01022
R14529 DVDD.n2761 DVDD.n2760 0.01022
R14530 DVDD.n2760 DVDD.n2749 0.01022
R14531 DVDD.n2756 DVDD.n2749 0.01022
R14532 DVDD.n2756 DVDD.n2755 0.01022
R14533 DVDD.n2755 DVDD.n2754 0.01022
R14534 DVDD.n2754 DVDD.n2751 0.01022
R14535 DVDD.n2751 DVDD.n2738 0.01022
R14536 DVDD.n6921 DVDD.n2738 0.01022
R14537 DVDD.n6921 DVDD.n6920 0.01022
R14538 DVDD.n6920 DVDD.n6918 0.01022
R14539 DVDD.n6918 DVDD.n6916 0.01022
R14540 DVDD.n6916 DVDD.n6913 0.01022
R14541 DVDD.n6913 DVDD.n6912 0.01022
R14542 DVDD.n6912 DVDD.n6910 0.01022
R14543 DVDD.n6910 DVDD.n6908 0.01022
R14544 DVDD.n6908 DVDD.n6906 0.01022
R14545 DVDD.n6906 DVDD.n6904 0.01022
R14546 DVDD.n6927 DVDD.n2654 0.01022
R14547 DVDD.n2676 DVDD.n2654 0.01022
R14548 DVDD.n2721 DVDD.n2676 0.01022
R14549 DVDD.n2721 DVDD.n2720 0.01022
R14550 DVDD.n2720 DVDD.n2718 0.01022
R14551 DVDD.n2718 DVDD.n2715 0.01022
R14552 DVDD.n2715 DVDD.n2714 0.01022
R14553 DVDD.n2714 DVDD.n2712 0.01022
R14554 DVDD.n2712 DVDD.n2710 0.01022
R14555 DVDD.n2710 DVDD.n2677 0.01022
R14556 DVDD.n2706 DVDD.n2677 0.01022
R14557 DVDD.n2706 DVDD.n2705 0.01022
R14558 DVDD.n2705 DVDD.n2703 0.01022
R14559 DVDD.n2703 DVDD.n2701 0.01022
R14560 DVDD.n2701 DVDD.n2698 0.01022
R14561 DVDD.n2698 DVDD.n2697 0.01022
R14562 DVDD.n2697 DVDD.n2695 0.01022
R14563 DVDD.n2695 DVDD.n2693 0.01022
R14564 DVDD.n2693 DVDD.n2691 0.01022
R14565 DVDD.n2691 DVDD.n2689 0.01022
R14566 DVDD.n2689 DVDD.n2687 0.01022
R14567 DVDD.n2687 DVDD.n2685 0.01022
R14568 DVDD.n2685 DVDD.n2682 0.01022
R14569 DVDD.n2682 DVDD.n2681 0.01022
R14570 DVDD.n2681 DVDD.n2679 0.01022
R14571 DVDD.n2679 DVDD.n2650 0.01022
R14572 DVDD.n6930 DVDD.n2650 0.01022
R14573 DVDD.n6930 DVDD.n6929 0.01022
R14574 DVDD.n724 DVDD.n722 0.01022
R14575 DVDD.n722 DVDD.n719 0.01022
R14576 DVDD.n719 DVDD.n718 0.01022
R14577 DVDD.n718 DVDD.n716 0.01022
R14578 DVDD.n716 DVDD.n714 0.01022
R14579 DVDD.n714 DVDD.n712 0.01022
R14580 DVDD.n712 DVDD.n710 0.01022
R14581 DVDD.n710 DVDD.n708 0.01022
R14582 DVDD.n708 DVDD.n706 0.01022
R14583 DVDD.n706 DVDD.n703 0.01022
R14584 DVDD.n703 DVDD.n702 0.01022
R14585 DVDD.n702 DVDD.n701 0.01022
R14586 DVDD.n701 DVDD.n700 0.01022
R14587 DVDD.n700 DVDD.n689 0.01022
R14588 DVDD.n696 DVDD.n689 0.01022
R14589 DVDD.n696 DVDD.n695 0.01022
R14590 DVDD.n695 DVDD.n694 0.01022
R14591 DVDD.n694 DVDD.n691 0.01022
R14592 DVDD.n691 DVDD.n688 0.01022
R14593 DVDD.n745 DVDD.n688 0.01022
R14594 DVDD.n749 DVDD.n748 0.01022
R14595 DVDD.n750 DVDD.n749 0.01022
R14596 DVDD.n750 DVDD.n685 0.01022
R14597 DVDD.n754 DVDD.n685 0.01022
R14598 DVDD.n755 DVDD.n754 0.01022
R14599 DVDD.n756 DVDD.n755 0.01022
R14600 DVDD.n756 DVDD.n683 0.01022
R14601 DVDD.n760 DVDD.n683 0.01022
R14602 DVDD.n761 DVDD.n760 0.01022
R14603 DVDD.n762 DVDD.n761 0.01022
R14604 DVDD.n762 DVDD.n681 0.01022
R14605 DVDD.n766 DVDD.n681 0.01022
R14606 DVDD.n767 DVDD.n766 0.01022
R14607 DVDD.n768 DVDD.n767 0.01022
R14608 DVDD.n768 DVDD.n679 0.01022
R14609 DVDD.n772 DVDD.n679 0.01022
R14610 DVDD.n773 DVDD.n772 0.01022
R14611 DVDD.n774 DVDD.n773 0.01022
R14612 DVDD.n774 DVDD.n677 0.01022
R14613 DVDD.n778 DVDD.n677 0.01022
R14614 DVDD.n779 DVDD.n778 0.01022
R14615 DVDD.n780 DVDD.n779 0.01022
R14616 DVDD.n780 DVDD.n675 0.01022
R14617 DVDD.n784 DVDD.n675 0.01022
R14618 DVDD.n785 DVDD.n784 0.01022
R14619 DVDD.n786 DVDD.n785 0.01022
R14620 DVDD.n786 DVDD.n673 0.01022
R14621 DVDD.n8837 DVDD.n673 0.01022
R14622 DVDD.n8834 DVDD.n8833 0.01022
R14623 DVDD.n8833 DVDD.n8832 0.01022
R14624 DVDD.n8832 DVDD.n8797 0.01022
R14625 DVDD.n8828 DVDD.n8797 0.01022
R14626 DVDD.n8828 DVDD.n8827 0.01022
R14627 DVDD.n8827 DVDD.n8826 0.01022
R14628 DVDD.n8826 DVDD.n8799 0.01022
R14629 DVDD.n8822 DVDD.n8799 0.01022
R14630 DVDD.n8822 DVDD.n8821 0.01022
R14631 DVDD.n8821 DVDD.n8819 0.01022
R14632 DVDD.n8819 DVDD.n8816 0.01022
R14633 DVDD.n8816 DVDD.n8815 0.01022
R14634 DVDD.n8815 DVDD.n8813 0.01022
R14635 DVDD.n8813 DVDD.n8811 0.01022
R14636 DVDD.n8811 DVDD.n8809 0.01022
R14637 DVDD.n8809 DVDD.n8807 0.01022
R14638 DVDD.n8807 DVDD.n8805 0.01022
R14639 DVDD.n8805 DVDD.n8803 0.01022
R14640 DVDD.n8803 DVDD.n8800 0.01022
R14641 DVDD.n8800 DVDD.n75 0.01022
R14642 DVDD.n9644 DVDD.n75 0.01022
R14643 DVDD.n9644 DVDD.n9643 0.01022
R14644 DVDD.n9643 DVDD.n9642 0.01022
R14645 DVDD.n9642 DVDD.n76 0.01022
R14646 DVDD.n9638 DVDD.n76 0.01022
R14647 DVDD.n9638 DVDD.n9637 0.01022
R14648 DVDD.n9637 DVDD.n9636 0.01022
R14649 DVDD.n9636 DVDD.n78 0.01022
R14650 DVDD.n9632 DVDD.n9631 0.01022
R14651 DVDD.n9631 DVDD.n9630 0.01022
R14652 DVDD.n9630 DVDD.n80 0.01022
R14653 DVDD.n844 DVDD.n80 0.01022
R14654 DVDD.n845 DVDD.n844 0.01022
R14655 DVDD.n846 DVDD.n845 0.01022
R14656 DVDD.n8769 DVDD.n846 0.01022
R14657 DVDD.n8769 DVDD.n8768 0.01022
R14658 DVDD.n8768 DVDD.n847 0.01022
R14659 DVDD.n930 DVDD.n847 0.01022
R14660 DVDD.n939 DVDD.n930 0.01022
R14661 DVDD.n939 DVDD.n938 0.01022
R14662 DVDD.n938 DVDD.n937 0.01022
R14663 DVDD.n937 DVDD.n936 0.01022
R14664 DVDD.n936 DVDD.n932 0.01022
R14665 DVDD.n932 DVDD.n931 0.01022
R14666 DVDD.n931 DVDD.n878 0.01022
R14667 DVDD.n8743 DVDD.n878 0.01022
R14668 DVDD.n8743 DVDD.n8742 0.01022
R14669 DVDD.n8742 DVDD.n879 0.01022
R14670 DVDD.n887 DVDD.n879 0.01022
R14671 DVDD.n8722 DVDD.n887 0.01022
R14672 DVDD.n8722 DVDD.n8721 0.01022
R14673 DVDD.n8721 DVDD.n888 0.01022
R14674 DVDD.n914 DVDD.n888 0.01022
R14675 DVDD.n915 DVDD.n914 0.01022
R14676 DVDD.n998 DVDD.n915 0.01022
R14677 DVDD.n999 DVDD.n998 0.01022
R14678 DVDD.n3637 DVDD.n3582 0.01022
R14679 DVDD.n3638 DVDD.n3637 0.01022
R14680 DVDD.n3739 DVDD.n3638 0.01022
R14681 DVDD.n3739 DVDD.n3738 0.01022
R14682 DVDD.n3738 DVDD.n3737 0.01022
R14683 DVDD.n3737 DVDD.n3736 0.01022
R14684 DVDD.n3736 DVDD.n3735 0.01022
R14685 DVDD.n3735 DVDD.n3639 0.01022
R14686 DVDD.n3731 DVDD.n3639 0.01022
R14687 DVDD.n3731 DVDD.n3730 0.01022
R14688 DVDD.n3730 DVDD.n3729 0.01022
R14689 DVDD.n3729 DVDD.n3642 0.01022
R14690 DVDD.n3725 DVDD.n3642 0.01022
R14691 DVDD.n3725 DVDD.n3724 0.01022
R14692 DVDD.n3724 DVDD.n3723 0.01022
R14693 DVDD.n3723 DVDD.n3644 0.01022
R14694 DVDD.n3719 DVDD.n3644 0.01022
R14695 DVDD.n3719 DVDD.n3718 0.01022
R14696 DVDD.n3718 DVDD.n3717 0.01022
R14697 DVDD.n3717 DVDD.n3646 0.01022
R14698 DVDD.n3713 DVDD.n3646 0.01022
R14699 DVDD.n3713 DVDD.n3712 0.01022
R14700 DVDD.n3712 DVDD.n3711 0.01022
R14701 DVDD.n3711 DVDD.n3648 0.01022
R14702 DVDD.n3707 DVDD.n3648 0.01022
R14703 DVDD.n3707 DVDD.n3706 0.01022
R14704 DVDD.n3706 DVDD.n3705 0.01022
R14705 DVDD.n3705 DVDD.n3581 0.01022
R14706 DVDD.n3700 DVDD.n3577 0.01022
R14707 DVDD.n3700 DVDD.n3699 0.01022
R14708 DVDD.n3699 DVDD.n3698 0.01022
R14709 DVDD.n3698 DVDD.n3651 0.01022
R14710 DVDD.n3694 DVDD.n3651 0.01022
R14711 DVDD.n3694 DVDD.n3693 0.01022
R14712 DVDD.n3693 DVDD.n3692 0.01022
R14713 DVDD.n3692 DVDD.n3653 0.01022
R14714 DVDD.n3688 DVDD.n3653 0.01022
R14715 DVDD.n3688 DVDD.n3687 0.01022
R14716 DVDD.n3687 DVDD.n3686 0.01022
R14717 DVDD.n3686 DVDD.n3655 0.01022
R14718 DVDD.n3682 DVDD.n3655 0.01022
R14719 DVDD.n3682 DVDD.n3681 0.01022
R14720 DVDD.n3681 DVDD.n3680 0.01022
R14721 DVDD.n3680 DVDD.n3657 0.01022
R14722 DVDD.n3676 DVDD.n3657 0.01022
R14723 DVDD.n3676 DVDD.n3675 0.01022
R14724 DVDD.n3675 DVDD.n3674 0.01022
R14725 DVDD.n3674 DVDD.n3659 0.01022
R14726 DVDD.n3670 DVDD.n3659 0.01022
R14727 DVDD.n3670 DVDD.n3669 0.01022
R14728 DVDD.n3669 DVDD.n3668 0.01022
R14729 DVDD.n3668 DVDD.n3661 0.01022
R14730 DVDD.n3664 DVDD.n3661 0.01022
R14731 DVDD.n3664 DVDD.n3663 0.01022
R14732 DVDD.n3663 DVDD.n3575 0.01022
R14733 DVDD.n3803 DVDD.n3575 0.01022
R14734 DVDD.n6337 DVDD.n3555 0.01022
R14735 DVDD.n3821 DVDD.n3555 0.01022
R14736 DVDD.n3823 DVDD.n3821 0.01022
R14737 DVDD.n3824 DVDD.n3823 0.01022
R14738 DVDD.n3827 DVDD.n3824 0.01022
R14739 DVDD.n3829 DVDD.n3827 0.01022
R14740 DVDD.n3831 DVDD.n3829 0.01022
R14741 DVDD.n3833 DVDD.n3831 0.01022
R14742 DVDD.n3835 DVDD.n3833 0.01022
R14743 DVDD.n3837 DVDD.n3835 0.01022
R14744 DVDD.n3839 DVDD.n3837 0.01022
R14745 DVDD.n3840 DVDD.n3839 0.01022
R14746 DVDD.n3843 DVDD.n3840 0.01022
R14747 DVDD.n3845 DVDD.n3843 0.01022
R14748 DVDD.n3847 DVDD.n3845 0.01022
R14749 DVDD.n3849 DVDD.n3847 0.01022
R14750 DVDD.n3851 DVDD.n3849 0.01022
R14751 DVDD.n3853 DVDD.n3851 0.01022
R14752 DVDD.n3855 DVDD.n3853 0.01022
R14753 DVDD.n3856 DVDD.n3855 0.01022
R14754 DVDD.n3859 DVDD.n3856 0.01022
R14755 DVDD.n3860 DVDD.n3859 0.01022
R14756 DVDD.n6331 DVDD.n3860 0.01022
R14757 DVDD.n6331 DVDD.n6330 0.01022
R14758 DVDD.n6330 DVDD.n6329 0.01022
R14759 DVDD.n6329 DVDD.n3861 0.01022
R14760 DVDD.n6322 DVDD.n3861 0.01022
R14761 DVDD.n6322 DVDD.n3554 0.01022
R14762 DVDD.n6297 DVDD.n3417 0.01022
R14763 DVDD.n6297 DVDD.n6296 0.01022
R14764 DVDD.n6296 DVDD.n6295 0.01022
R14765 DVDD.n6295 DVDD.n6246 0.01022
R14766 DVDD.n6291 DVDD.n6246 0.01022
R14767 DVDD.n6291 DVDD.n6290 0.01022
R14768 DVDD.n6290 DVDD.n6289 0.01022
R14769 DVDD.n6289 DVDD.n6248 0.01022
R14770 DVDD.n6285 DVDD.n6248 0.01022
R14771 DVDD.n6285 DVDD.n6284 0.01022
R14772 DVDD.n6284 DVDD.n6283 0.01022
R14773 DVDD.n6283 DVDD.n6250 0.01022
R14774 DVDD.n6279 DVDD.n6250 0.01022
R14775 DVDD.n6279 DVDD.n6278 0.01022
R14776 DVDD.n6278 DVDD.n6277 0.01022
R14777 DVDD.n6277 DVDD.n6252 0.01022
R14778 DVDD.n6273 DVDD.n6252 0.01022
R14779 DVDD.n6273 DVDD.n6272 0.01022
R14780 DVDD.n6272 DVDD.n6271 0.01022
R14781 DVDD.n6271 DVDD.n6269 0.01022
R14782 DVDD.n6269 DVDD.n6267 0.01022
R14783 DVDD.n6267 DVDD.n6265 0.01022
R14784 DVDD.n6265 DVDD.n6262 0.01022
R14785 DVDD.n6262 DVDD.n6261 0.01022
R14786 DVDD.n6261 DVDD.n6259 0.01022
R14787 DVDD.n6259 DVDD.n6257 0.01022
R14788 DVDD.n6257 DVDD.n6255 0.01022
R14789 DVDD.n6255 DVDD.n3416 0.01022
R14790 DVDD.n6543 DVDD.n6541 0.01022
R14791 DVDD.n6541 DVDD.n6539 0.01022
R14792 DVDD.n6539 DVDD.n6537 0.01022
R14793 DVDD.n6537 DVDD.n6535 0.01022
R14794 DVDD.n6535 DVDD.n6533 0.01022
R14795 DVDD.n6533 DVDD.n6530 0.01022
R14796 DVDD.n6530 DVDD.n6529 0.01022
R14797 DVDD.n6529 DVDD.n6527 0.01022
R14798 DVDD.n6527 DVDD.n6526 0.01022
R14799 DVDD.n6526 DVDD.n6525 0.01022
R14800 DVDD.n6525 DVDD.n6522 0.01022
R14801 DVDD.n6522 DVDD.n6521 0.01022
R14802 DVDD.n6521 DVDD.n6519 0.01022
R14803 DVDD.n6519 DVDD.n6517 0.01022
R14804 DVDD.n6517 DVDD.n6514 0.01022
R14805 DVDD.n6514 DVDD.n6513 0.01022
R14806 DVDD.n6513 DVDD.n6511 0.01022
R14807 DVDD.n6511 DVDD.n6509 0.01022
R14808 DVDD.n6509 DVDD.n6507 0.01022
R14809 DVDD.n6507 DVDD.n6505 0.01022
R14810 DVDD.n6505 DVDD.n6503 0.01022
R14811 DVDD.n6503 DVDD.n6501 0.01022
R14812 DVDD.n6501 DVDD.n6498 0.01022
R14813 DVDD.n6498 DVDD.n6497 0.01022
R14814 DVDD.n6497 DVDD.n6495 0.01022
R14815 DVDD.n6495 DVDD.n6493 0.01022
R14816 DVDD.n6493 DVDD.n6491 0.01022
R14817 DVDD.n6491 DVDD.n6489 0.01022
R14818 DVDD.n6586 DVDD.n2044 0.0101025
R14819 DVDD.n6584 DVDD.n2041 0.0101025
R14820 DVDD.n6582 DVDD.n2045 0.0101025
R14821 DVDD.n6580 DVDD.n2040 0.0101025
R14822 DVDD.n6578 DVDD.n2046 0.0101025
R14823 DVDD.n6576 DVDD.n2039 0.0101025
R14824 DVDD.n6574 DVDD.n2047 0.0101025
R14825 DVDD.n6572 DVDD.n2038 0.0101025
R14826 DVDD.n6570 DVDD.n2048 0.0101025
R14827 DVDD.n6568 DVDD.n2037 0.0101025
R14828 DVDD.n6566 DVDD.n2049 0.0101025
R14829 DVDD.n6564 DVDD.n2036 0.0101025
R14830 DVDD.n6562 DVDD.n2050 0.0101025
R14831 DVDD.n6560 DVDD.n2035 0.0101025
R14832 DVDD.n6558 DVDD.n2052 0.0101025
R14833 DVDD.n207 DVDD.n206 0.00992
R14834 DVDD.n9571 DVDD.n9570 0.00992
R14835 DVDD.n9489 DVDD.n271 0.00992
R14836 DVDD.n4130 DVDD.n3986 0.00992
R14837 DVDD.n9490 DVDD.n277 0.00992
R14838 DVDD.n1025 DVDD.n1024 0.00992
R14839 DVDD.n4129 DVDD.n3980 0.00992
R14840 DVDD.n911 DVDD.n907 0.00992
R14841 DVDD.n8808 DVDD.n62 0.00988976
R14842 DVDD.n8687 DVDD.n1010 0.00988976
R14843 DVDD.n3848 DVDD.n3564 0.00988976
R14844 DVDD.n6327 DVDD.n3863 0.00988976
R14845 DVDD.n6540 DVDD.n3353 0.00988976
R14846 DVDD.n6508 DVDD.n2079 0.00988976
R14847 DVDD.n7664 DVDD.n1982 0.00988976
R14848 DVDD.n9080 DVDD.n522 0.00988976
R14849 DVDD.n4219 DVDD.n4146 0.00988976
R14850 DVDD.n6020 DVDD.n3961 0.00988976
R14851 DVDD.n6061 DVDD.n6060 0.00988976
R14852 DVDD.n3246 DVDD.n3229 0.00988976
R14853 DVDD.n3271 DVDD.n2124 0.00988976
R14854 DVDD.n2296 DVDD.n2291 0.00988976
R14855 DVDD.n4923 DVDD.n486 0.00988976
R14856 DVDD.n9510 DVDD.n9506 0.00988976
R14857 DVDD.n5787 DVDD.n4308 0.00988976
R14858 DVDD.n5769 DVDD.n5766 0.00988976
R14859 DVDD.n3137 DVDD.n3118 0.00988976
R14860 DVDD.n3162 DVDD.n2176 0.00988976
R14861 DVDD.n7673 DVDD.n2245 0.00988976
R14862 DVDD.n9261 DVDD.n462 0.00988976
R14863 DVDD.n6795 DVDD.n2889 0.00988976
R14864 DVDD.n2847 DVDD.n2823 0.00988976
R14865 DVDD.n6866 DVDD.n6865 0.00988976
R14866 DVDD.n2668 DVDD.n2658 0.00988976
R14867 DVDD.n2692 DVDD.n2644 0.00988976
R14868 DVDD.n2450 DVDD.n2376 0.00988976
R14869 DVDD.n6556 DVDD.n6473 0.00972594
R14870 DVDD.n6554 DVDD.n3399 0.00972594
R14871 DVDD.n6552 DVDD.n6474 0.00972594
R14872 DVDD.n6550 DVDD.n3398 0.00972594
R14873 DVDD.n6548 DVDD.n6475 0.00972594
R14874 DVDD.n6546 DVDD.n3397 0.00972594
R14875 DVDD.n6544 DVDD.n6476 0.00972594
R14876 DVDD.n6477 DVDD.n3396 0.00972594
R14877 DVDD.n4708 DVDD.n4612 0.00962857
R14878 DVDD.n4715 DVDD.n4612 0.00962857
R14879 DVDD.n4715 DVDD.n4610 0.00962857
R14880 DVDD.n4719 DVDD.n4610 0.00962857
R14881 DVDD.n4719 DVDD.n4608 0.00962857
R14882 DVDD.n4723 DVDD.n4608 0.00962857
R14883 DVDD.n4723 DVDD.n4606 0.00962857
R14884 DVDD.n4727 DVDD.n4606 0.00962857
R14885 DVDD.n4727 DVDD.n4592 0.00962857
R14886 DVDD.n4823 DVDD.n4592 0.00962857
R14887 DVDD.n4823 DVDD.n4590 0.00962857
R14888 DVDD.n4827 DVDD.n4590 0.00962857
R14889 DVDD.n4827 DVDD.n4588 0.00962857
R14890 DVDD.n4831 DVDD.n4588 0.00962857
R14891 DVDD.n4831 DVDD.n4586 0.00962857
R14892 DVDD.n4835 DVDD.n4586 0.00962857
R14893 DVDD.n4835 DVDD.n4584 0.00962857
R14894 DVDD.n4839 DVDD.n4584 0.00962857
R14895 DVDD.n4839 DVDD.n4580 0.00962857
R14896 DVDD.n5114 DVDD.n4580 0.00962857
R14897 DVDD.n5114 DVDD.n4582 0.00962857
R14898 DVDD.n5110 DVDD.n4582 0.00962857
R14899 DVDD.n5110 DVDD.n5108 0.00962857
R14900 DVDD.n5108 DVDD.n4843 0.00962857
R14901 DVDD.n5104 DVDD.n4843 0.00962857
R14902 DVDD.n5104 DVDD.n4845 0.00962857
R14903 DVDD.n5100 DVDD.n4845 0.00962857
R14904 DVDD.n5100 DVDD.n4848 0.00962857
R14905 DVDD.n5096 DVDD.n4848 0.00962857
R14906 DVDD.n5096 DVDD.n4850 0.00962857
R14907 DVDD.n5092 DVDD.n4850 0.00962857
R14908 DVDD.n5092 DVDD.n4852 0.00962857
R14909 DVDD.n5088 DVDD.n4852 0.00962857
R14910 DVDD.n5088 DVDD.n4854 0.00962857
R14911 DVDD.n5084 DVDD.n4854 0.00962857
R14912 DVDD.n5084 DVDD.n4856 0.00962857
R14913 DVDD.n5034 DVDD.n4856 0.00962857
R14914 DVDD.n5034 DVDD.n5031 0.00962857
R14915 DVDD.n5078 DVDD.n5031 0.00962857
R14916 DVDD.n5078 DVDD.n5032 0.00962857
R14917 DVDD.n5074 DVDD.n5032 0.00962857
R14918 DVDD.n5074 DVDD.n5038 0.00962857
R14919 DVDD.n5070 DVDD.n5038 0.00962857
R14920 DVDD.n5070 DVDD.n5040 0.00962857
R14921 DVDD.n5066 DVDD.n5040 0.00962857
R14922 DVDD.n5066 DVDD.n5042 0.00962857
R14923 DVDD.n5062 DVDD.n5042 0.00962857
R14924 DVDD.n5062 DVDD.n5044 0.00962857
R14925 DVDD.n5058 DVDD.n5044 0.00962857
R14926 DVDD.n5058 DVDD.n5046 0.00962857
R14927 DVDD.n5054 DVDD.n5046 0.00962857
R14928 DVDD.n5054 DVDD.n5048 0.00962857
R14929 DVDD.n5050 DVDD.n5048 0.00962857
R14930 DVDD.n5050 DVDD.n558 0.00962857
R14931 DVDD.n8970 DVDD.n558 0.00962857
R14932 DVDD.n8970 DVDD.n560 0.00962857
R14933 DVDD.n8966 DVDD.n560 0.00962857
R14934 DVDD.n8966 DVDD.n8964 0.00962857
R14935 DVDD.n8964 DVDD.n563 0.00962857
R14936 DVDD.n8960 DVDD.n563 0.00962857
R14937 DVDD.n8960 DVDD.n565 0.00962857
R14938 DVDD.n8956 DVDD.n565 0.00962857
R14939 DVDD.n8956 DVDD.n568 0.00962857
R14940 DVDD.n8952 DVDD.n568 0.00962857
R14941 DVDD.n8952 DVDD.n570 0.00962857
R14942 DVDD.n8948 DVDD.n570 0.00962857
R14943 DVDD.n8948 DVDD.n572 0.00962857
R14944 DVDD.n8944 DVDD.n572 0.00962857
R14945 DVDD.n8944 DVDD.n574 0.00962857
R14946 DVDD.n8940 DVDD.n574 0.00962857
R14947 DVDD.n8940 DVDD.n576 0.00962857
R14948 DVDD.n597 DVDD.n576 0.00962857
R14949 DVDD.n597 DVDD.n594 0.00962857
R14950 DVDD.n8934 DVDD.n594 0.00962857
R14951 DVDD.n8934 DVDD.n595 0.00962857
R14952 DVDD.n8930 DVDD.n595 0.00962857
R14953 DVDD.n8930 DVDD.n601 0.00962857
R14954 DVDD.n8926 DVDD.n601 0.00962857
R14955 DVDD.n8926 DVDD.n603 0.00962857
R14956 DVDD.n8922 DVDD.n603 0.00962857
R14957 DVDD.n8922 DVDD.n605 0.00962857
R14958 DVDD.n8918 DVDD.n605 0.00962857
R14959 DVDD.n8918 DVDD.n607 0.00962857
R14960 DVDD.n8914 DVDD.n607 0.00962857
R14961 DVDD.n8914 DVDD.n609 0.00962857
R14962 DVDD.n8908 DVDD.n609 0.00962857
R14963 DVDD.n8908 DVDD.n634 0.00962857
R14964 DVDD.n8904 DVDD.n634 0.00962857
R14965 DVDD.n8904 DVDD.n636 0.00962857
R14966 DVDD.n8900 DVDD.n636 0.00962857
R14967 DVDD.n8900 DVDD.n638 0.00962857
R14968 DVDD.n8896 DVDD.n638 0.00962857
R14969 DVDD.n8896 DVDD.n640 0.00962857
R14970 DVDD.n7501 DVDD.n7090 0.00962857
R14971 DVDD.n7501 DVDD.n7092 0.00962857
R14972 DVDD.n7497 DVDD.n7092 0.00962857
R14973 DVDD.n7497 DVDD.n7094 0.00962857
R14974 DVDD.n7493 DVDD.n7094 0.00962857
R14975 DVDD.n7493 DVDD.n7096 0.00962857
R14976 DVDD.n7489 DVDD.n7096 0.00962857
R14977 DVDD.n7489 DVDD.n7098 0.00962857
R14978 DVDD.n7305 DVDD.n7098 0.00962857
R14979 DVDD.n7483 DVDD.n7305 0.00962857
R14980 DVDD.n7483 DVDD.n7306 0.00962857
R14981 DVDD.n7479 DVDD.n7306 0.00962857
R14982 DVDD.n7479 DVDD.n7309 0.00962857
R14983 DVDD.n7475 DVDD.n7309 0.00962857
R14984 DVDD.n7475 DVDD.n7312 0.00962857
R14985 DVDD.n7471 DVDD.n7312 0.00962857
R14986 DVDD.n7471 DVDD.n7314 0.00962857
R14987 DVDD.n7467 DVDD.n7314 0.00962857
R14988 DVDD.n7467 DVDD.n7315 0.00962857
R14989 DVDD.n7463 DVDD.n7315 0.00962857
R14990 DVDD.n7463 DVDD.n7462 0.00962857
R14991 DVDD.n7462 DVDD.n7461 0.00962857
R14992 DVDD.n7461 DVDD.n7317 0.00962857
R14993 DVDD.n7456 DVDD.n7317 0.00962857
R14994 DVDD.n7456 DVDD.n7319 0.00962857
R14995 DVDD.n7452 DVDD.n7319 0.00962857
R14996 DVDD.n7452 DVDD.n7322 0.00962857
R14997 DVDD.n7448 DVDD.n7322 0.00962857
R14998 DVDD.n7448 DVDD.n7324 0.00962857
R14999 DVDD.n7444 DVDD.n7324 0.00962857
R15000 DVDD.n7444 DVDD.n7326 0.00962857
R15001 DVDD.n7440 DVDD.n7326 0.00962857
R15002 DVDD.n7440 DVDD.n7328 0.00962857
R15003 DVDD.n7436 DVDD.n7328 0.00962857
R15004 DVDD.n7436 DVDD.n7330 0.00962857
R15005 DVDD.n7432 DVDD.n7330 0.00962857
R15006 DVDD.n7432 DVDD.n7332 0.00962857
R15007 DVDD.n7374 DVDD.n7332 0.00962857
R15008 DVDD.n7420 DVDD.n7374 0.00962857
R15009 DVDD.n7420 DVDD.n7375 0.00962857
R15010 DVDD.n7416 DVDD.n7375 0.00962857
R15011 DVDD.n7416 DVDD.n7378 0.00962857
R15012 DVDD.n7412 DVDD.n7378 0.00962857
R15013 DVDD.n7412 DVDD.n7380 0.00962857
R15014 DVDD.n7408 DVDD.n7380 0.00962857
R15015 DVDD.n7408 DVDD.n7382 0.00962857
R15016 DVDD.n7404 DVDD.n7382 0.00962857
R15017 DVDD.n7404 DVDD.n7384 0.00962857
R15018 DVDD.n7400 DVDD.n7384 0.00962857
R15019 DVDD.n7400 DVDD.n7386 0.00962857
R15020 DVDD.n7396 DVDD.n7386 0.00962857
R15021 DVDD.n7396 DVDD.n7388 0.00962857
R15022 DVDD.n7392 DVDD.n7388 0.00962857
R15023 DVDD.n7392 DVDD.n7390 0.00962857
R15024 DVDD.n7390 DVDD.n1723 0.00962857
R15025 DVDD.n8282 DVDD.n1723 0.00962857
R15026 DVDD.n8282 DVDD.n1725 0.00962857
R15027 DVDD.n8278 DVDD.n1725 0.00962857
R15028 DVDD.n8278 DVDD.n1728 0.00962857
R15029 DVDD.n8274 DVDD.n1728 0.00962857
R15030 DVDD.n8274 DVDD.n1730 0.00962857
R15031 DVDD.n8270 DVDD.n1730 0.00962857
R15032 DVDD.n8270 DVDD.n1732 0.00962857
R15033 DVDD.n8266 DVDD.n1732 0.00962857
R15034 DVDD.n8266 DVDD.n1734 0.00962857
R15035 DVDD.n8262 DVDD.n1734 0.00962857
R15036 DVDD.n8262 DVDD.n1736 0.00962857
R15037 DVDD.n8258 DVDD.n1736 0.00962857
R15038 DVDD.n8258 DVDD.n1738 0.00962857
R15039 DVDD.n8254 DVDD.n1738 0.00962857
R15040 DVDD.n8254 DVDD.n1740 0.00962857
R15041 DVDD.n1764 DVDD.n1740 0.00962857
R15042 DVDD.n8248 DVDD.n1764 0.00962857
R15043 DVDD.n8248 DVDD.n1765 0.00962857
R15044 DVDD.n8244 DVDD.n1765 0.00962857
R15045 DVDD.n8244 DVDD.n1768 0.00962857
R15046 DVDD.n8240 DVDD.n1768 0.00962857
R15047 DVDD.n8240 DVDD.n1771 0.00962857
R15048 DVDD.n8236 DVDD.n1771 0.00962857
R15049 DVDD.n8236 DVDD.n1773 0.00962857
R15050 DVDD.n8232 DVDD.n1773 0.00962857
R15051 DVDD.n8232 DVDD.n1774 0.00962857
R15052 DVDD.n8228 DVDD.n1774 0.00962857
R15053 DVDD.n8228 DVDD.n8227 0.00962857
R15054 DVDD.n8227 DVDD.n8225 0.00962857
R15055 DVDD.n8225 DVDD.n1776 0.00962857
R15056 DVDD.n8220 DVDD.n1776 0.00962857
R15057 DVDD.n8220 DVDD.n1778 0.00962857
R15058 DVDD.n8216 DVDD.n1778 0.00962857
R15059 DVDD.n8216 DVDD.n1781 0.00962857
R15060 DVDD.n8212 DVDD.n1781 0.00962857
R15061 DVDD.n8212 DVDD.n1783 0.00962857
R15062 DVDD.n8200 DVDD.n1783 0.00962857
R15063 DVDD.n7496 DVDD.n7495 0.00962857
R15064 DVDD.n7495 DVDD.n7494 0.00962857
R15065 DVDD.n7494 DVDD.n7095 0.00962857
R15066 DVDD.n7488 DVDD.n7095 0.00962857
R15067 DVDD.n7478 DVDD.n7310 0.00962857
R15068 DVDD.n7478 DVDD.n7477 0.00962857
R15069 DVDD.n7477 DVDD.n7476 0.00962857
R15070 DVDD.n7476 DVDD.n7311 0.00962857
R15071 DVDD.n7470 DVDD.n7311 0.00962857
R15072 DVDD.n7470 DVDD.n7469 0.00962857
R15073 DVDD.n7469 DVDD.n7468 0.00962857
R15074 DVDD.n7468 DVDD.n1514 0.00962857
R15075 DVDD.n7455 DVDD.n7320 0.00962857
R15076 DVDD.n7455 DVDD.n7454 0.00962857
R15077 DVDD.n7454 DVDD.n7453 0.00962857
R15078 DVDD.n7453 DVDD.n7321 0.00962857
R15079 DVDD.n7447 DVDD.n7321 0.00962857
R15080 DVDD.n7447 DVDD.n7446 0.00962857
R15081 DVDD.n7446 DVDD.n7445 0.00962857
R15082 DVDD.n7445 DVDD.n7325 0.00962857
R15083 DVDD.n7439 DVDD.n7325 0.00962857
R15084 DVDD.n7439 DVDD.n7438 0.00962857
R15085 DVDD.n7438 DVDD.n7437 0.00962857
R15086 DVDD.n7437 DVDD.n7329 0.00962857
R15087 DVDD.n7421 DVDD.n7373 0.00962857
R15088 DVDD.n7415 DVDD.n7373 0.00962857
R15089 DVDD.n7415 DVDD.n7414 0.00962857
R15090 DVDD.n7414 DVDD.n7413 0.00962857
R15091 DVDD.n7413 DVDD.n7379 0.00962857
R15092 DVDD.n7407 DVDD.n7379 0.00962857
R15093 DVDD.n7407 DVDD.n7406 0.00962857
R15094 DVDD.n7406 DVDD.n7405 0.00962857
R15095 DVDD.n7405 DVDD.n7383 0.00962857
R15096 DVDD.n7399 DVDD.n7383 0.00962857
R15097 DVDD.n7399 DVDD.n7398 0.00962857
R15098 DVDD.n7398 DVDD.n7397 0.00962857
R15099 DVDD.n7397 DVDD.n7387 0.00962857
R15100 DVDD.n7391 DVDD.n7387 0.00962857
R15101 DVDD.n7391 DVDD.n1705 0.00962857
R15102 DVDD.n8277 DVDD.n8276 0.00962857
R15103 DVDD.n8276 DVDD.n8275 0.00962857
R15104 DVDD.n8275 DVDD.n1729 0.00962857
R15105 DVDD.n8269 DVDD.n1729 0.00962857
R15106 DVDD.n8269 DVDD.n8268 0.00962857
R15107 DVDD.n8268 DVDD.n8267 0.00962857
R15108 DVDD.n8267 DVDD.n1733 0.00962857
R15109 DVDD.n8261 DVDD.n1733 0.00962857
R15110 DVDD.n8261 DVDD.n8260 0.00962857
R15111 DVDD.n8260 DVDD.n8259 0.00962857
R15112 DVDD.n8259 DVDD.n1737 0.00962857
R15113 DVDD.n8253 DVDD.n1737 0.00962857
R15114 DVDD.n8243 DVDD.n1769 0.00962857
R15115 DVDD.n8243 DVDD.n8242 0.00962857
R15116 DVDD.n8242 DVDD.n8241 0.00962857
R15117 DVDD.n8241 DVDD.n1770 0.00962857
R15118 DVDD.n8235 DVDD.n1770 0.00962857
R15119 DVDD.n8235 DVDD.n8234 0.00962857
R15120 DVDD.n8234 DVDD.n8233 0.00962857
R15121 DVDD.n8233 DVDD.n1274 0.00962857
R15122 DVDD.n8219 DVDD.n1779 0.00962857
R15123 DVDD.n8219 DVDD.n8218 0.00962857
R15124 DVDD.n8218 DVDD.n8217 0.00962857
R15125 DVDD.n8217 DVDD.n1780 0.00962857
R15126 DVDD.n4720 DVDD.n4609 0.00962857
R15127 DVDD.n4721 DVDD.n4720 0.00962857
R15128 DVDD.n4722 DVDD.n4721 0.00962857
R15129 DVDD.n4722 DVDD.n4600 0.00962857
R15130 DVDD.n4828 DVDD.n4589 0.00962857
R15131 DVDD.n4829 DVDD.n4828 0.00962857
R15132 DVDD.n4830 DVDD.n4829 0.00962857
R15133 DVDD.n4830 DVDD.n4585 0.00962857
R15134 DVDD.n4836 DVDD.n4585 0.00962857
R15135 DVDD.n4837 DVDD.n4836 0.00962857
R15136 DVDD.n4838 DVDD.n4837 0.00962857
R15137 DVDD.n4838 DVDD.n4574 0.00962857
R15138 DVDD.n5107 DVDD.n5106 0.00962857
R15139 DVDD.n5106 DVDD.n5105 0.00962857
R15140 DVDD.n5105 DVDD.n4844 0.00962857
R15141 DVDD.n5099 DVDD.n4844 0.00962857
R15142 DVDD.n5099 DVDD.n5098 0.00962857
R15143 DVDD.n5098 DVDD.n5097 0.00962857
R15144 DVDD.n5097 DVDD.n4849 0.00962857
R15145 DVDD.n5091 DVDD.n4849 0.00962857
R15146 DVDD.n5091 DVDD.n5090 0.00962857
R15147 DVDD.n5090 DVDD.n5089 0.00962857
R15148 DVDD.n5089 DVDD.n4853 0.00962857
R15149 DVDD.n5083 DVDD.n4853 0.00962857
R15150 DVDD.n5079 DVDD.n5030 0.00962857
R15151 DVDD.n5073 DVDD.n5030 0.00962857
R15152 DVDD.n5073 DVDD.n5072 0.00962857
R15153 DVDD.n5072 DVDD.n5071 0.00962857
R15154 DVDD.n5071 DVDD.n5039 0.00962857
R15155 DVDD.n5065 DVDD.n5039 0.00962857
R15156 DVDD.n5065 DVDD.n5064 0.00962857
R15157 DVDD.n5064 DVDD.n5063 0.00962857
R15158 DVDD.n5063 DVDD.n5043 0.00962857
R15159 DVDD.n5057 DVDD.n5043 0.00962857
R15160 DVDD.n5057 DVDD.n5056 0.00962857
R15161 DVDD.n5056 DVDD.n5055 0.00962857
R15162 DVDD.n5055 DVDD.n5047 0.00962857
R15163 DVDD.n5049 DVDD.n5047 0.00962857
R15164 DVDD.n5049 DVDD.n552 0.00962857
R15165 DVDD.n8963 DVDD.n8962 0.00962857
R15166 DVDD.n8962 DVDD.n8961 0.00962857
R15167 DVDD.n8961 DVDD.n564 0.00962857
R15168 DVDD.n8955 DVDD.n564 0.00962857
R15169 DVDD.n8955 DVDD.n8954 0.00962857
R15170 DVDD.n8954 DVDD.n8953 0.00962857
R15171 DVDD.n8953 DVDD.n569 0.00962857
R15172 DVDD.n8947 DVDD.n569 0.00962857
R15173 DVDD.n8947 DVDD.n8946 0.00962857
R15174 DVDD.n8946 DVDD.n8945 0.00962857
R15175 DVDD.n8945 DVDD.n573 0.00962857
R15176 DVDD.n8939 DVDD.n573 0.00962857
R15177 DVDD.n8935 DVDD.n593 0.00962857
R15178 DVDD.n8929 DVDD.n593 0.00962857
R15179 DVDD.n8929 DVDD.n8928 0.00962857
R15180 DVDD.n8928 DVDD.n8927 0.00962857
R15181 DVDD.n8927 DVDD.n602 0.00962857
R15182 DVDD.n8921 DVDD.n602 0.00962857
R15183 DVDD.n8921 DVDD.n8920 0.00962857
R15184 DVDD.n8920 DVDD.n8919 0.00962857
R15185 DVDD.n8909 DVDD.n633 0.00962857
R15186 DVDD.n8903 DVDD.n633 0.00962857
R15187 DVDD.n8903 DVDD.n8902 0.00962857
R15188 DVDD.n8902 DVDD.n8901 0.00962857
R15189 DVDD.n4765 DVDD.n4764 0.00962857
R15190 DVDD.n4765 DVDD.n4753 0.00962857
R15191 DVDD.n4772 DVDD.n4753 0.00962857
R15192 DVDD.n4773 DVDD.n4772 0.00962857
R15193 DVDD.n4815 DVDD.n4748 0.00962857
R15194 DVDD.n4809 DVDD.n4748 0.00962857
R15195 DVDD.n4809 DVDD.n4808 0.00962857
R15196 DVDD.n4808 DVDD.n4807 0.00962857
R15197 DVDD.n4807 DVDD.n4796 0.00962857
R15198 DVDD.n4801 DVDD.n4796 0.00962857
R15199 DVDD.n4801 DVDD.n4800 0.00962857
R15200 DVDD.n4800 DVDD.n460 0.00962857
R15201 DVDD.n9235 DVDD.n9234 0.00962857
R15202 DVDD.n9234 DVDD.n9233 0.00962857
R15203 DVDD.n9233 DVDD.n471 0.00962857
R15204 DVDD.n9227 DVDD.n471 0.00962857
R15205 DVDD.n9227 DVDD.n9226 0.00962857
R15206 DVDD.n9226 DVDD.n9225 0.00962857
R15207 DVDD.n9225 DVDD.n476 0.00962857
R15208 DVDD.n9219 DVDD.n476 0.00962857
R15209 DVDD.n9219 DVDD.n9218 0.00962857
R15210 DVDD.n9218 DVDD.n9217 0.00962857
R15211 DVDD.n9217 DVDD.n480 0.00962857
R15212 DVDD.n9211 DVDD.n480 0.00962857
R15213 DVDD.n9207 DVDD.n500 0.00962857
R15214 DVDD.n9201 DVDD.n500 0.00962857
R15215 DVDD.n9201 DVDD.n9200 0.00962857
R15216 DVDD.n9200 DVDD.n9199 0.00962857
R15217 DVDD.n9199 DVDD.n509 0.00962857
R15218 DVDD.n9193 DVDD.n509 0.00962857
R15219 DVDD.n9193 DVDD.n9192 0.00962857
R15220 DVDD.n9192 DVDD.n9191 0.00962857
R15221 DVDD.n9191 DVDD.n513 0.00962857
R15222 DVDD.n9185 DVDD.n513 0.00962857
R15223 DVDD.n9185 DVDD.n9184 0.00962857
R15224 DVDD.n9184 DVDD.n9183 0.00962857
R15225 DVDD.n9183 DVDD.n517 0.00962857
R15226 DVDD.n9177 DVDD.n517 0.00962857
R15227 DVDD.n9177 DVDD.n9176 0.00962857
R15228 DVDD.n9166 DVDD.n9134 0.00962857
R15229 DVDD.n9166 DVDD.n9165 0.00962857
R15230 DVDD.n9165 DVDD.n9164 0.00962857
R15231 DVDD.n9164 DVDD.n9135 0.00962857
R15232 DVDD.n9158 DVDD.n9135 0.00962857
R15233 DVDD.n9158 DVDD.n9157 0.00962857
R15234 DVDD.n9157 DVDD.n9156 0.00962857
R15235 DVDD.n9156 DVDD.n9139 0.00962857
R15236 DVDD.n9150 DVDD.n9139 0.00962857
R15237 DVDD.n9150 DVDD.n9149 0.00962857
R15238 DVDD.n9149 DVDD.n9148 0.00962857
R15239 DVDD.n9148 DVDD.n9143 0.00962857
R15240 DVDD.n9655 DVDD.n9654 0.00962857
R15241 DVDD.n9656 DVDD.n9655 0.00962857
R15242 DVDD.n9656 DVDD.n51 0.00962857
R15243 DVDD.n9662 DVDD.n51 0.00962857
R15244 DVDD.n9663 DVDD.n9662 0.00962857
R15245 DVDD.n9664 DVDD.n9663 0.00962857
R15246 DVDD.n9664 DVDD.n47 0.00962857
R15247 DVDD.n9670 DVDD.n47 0.00962857
R15248 DVDD.n9682 DVDD.n9681 0.00962857
R15249 DVDD.n9683 DVDD.n9682 0.00962857
R15250 DVDD.n9683 DVDD.n16 0.00962857
R15251 DVDD.n9690 DVDD.n16 0.00962857
R15252 DVDD.n9694 DVDD.n0 0.00962857
R15253 DVDD.n4758 DVDD.n4756 0.00962857
R15254 DVDD.n4762 DVDD.n4758 0.00962857
R15255 DVDD.n4763 DVDD.n4762 0.00962857
R15256 DVDD.n4766 DVDD.n4763 0.00962857
R15257 DVDD.n4766 DVDD.n4754 0.00962857
R15258 DVDD.n4771 DVDD.n4754 0.00962857
R15259 DVDD.n4771 DVDD.n4752 0.00962857
R15260 DVDD.n4789 DVDD.n4752 0.00962857
R15261 DVDD.n4791 DVDD.n4789 0.00962857
R15262 DVDD.n4791 DVDD.n4749 0.00962857
R15263 DVDD.n4814 DVDD.n4749 0.00962857
R15264 DVDD.n4814 DVDD.n4750 0.00962857
R15265 DVDD.n4810 DVDD.n4750 0.00962857
R15266 DVDD.n4810 DVDD.n4795 0.00962857
R15267 DVDD.n4806 DVDD.n4795 0.00962857
R15268 DVDD.n4806 DVDD.n4797 0.00962857
R15269 DVDD.n4802 DVDD.n4797 0.00962857
R15270 DVDD.n4802 DVDD.n4799 0.00962857
R15271 DVDD.n4799 DVDD.n465 0.00962857
R15272 DVDD.n9242 DVDD.n465 0.00962857
R15273 DVDD.n9242 DVDD.n467 0.00962857
R15274 DVDD.n9238 DVDD.n467 0.00962857
R15275 DVDD.n9238 DVDD.n9236 0.00962857
R15276 DVDD.n9236 DVDD.n470 0.00962857
R15277 DVDD.n9232 DVDD.n470 0.00962857
R15278 DVDD.n9232 DVDD.n472 0.00962857
R15279 DVDD.n9228 DVDD.n472 0.00962857
R15280 DVDD.n9228 DVDD.n475 0.00962857
R15281 DVDD.n9224 DVDD.n475 0.00962857
R15282 DVDD.n9224 DVDD.n477 0.00962857
R15283 DVDD.n9220 DVDD.n477 0.00962857
R15284 DVDD.n9220 DVDD.n479 0.00962857
R15285 DVDD.n9216 DVDD.n479 0.00962857
R15286 DVDD.n9216 DVDD.n481 0.00962857
R15287 DVDD.n9212 DVDD.n481 0.00962857
R15288 DVDD.n9212 DVDD.n483 0.00962857
R15289 DVDD.n504 DVDD.n483 0.00962857
R15290 DVDD.n504 DVDD.n501 0.00962857
R15291 DVDD.n9206 DVDD.n501 0.00962857
R15292 DVDD.n9206 DVDD.n502 0.00962857
R15293 DVDD.n9202 DVDD.n502 0.00962857
R15294 DVDD.n9202 DVDD.n508 0.00962857
R15295 DVDD.n9198 DVDD.n508 0.00962857
R15296 DVDD.n9198 DVDD.n510 0.00962857
R15297 DVDD.n9194 DVDD.n510 0.00962857
R15298 DVDD.n9194 DVDD.n512 0.00962857
R15299 DVDD.n9190 DVDD.n512 0.00962857
R15300 DVDD.n9190 DVDD.n514 0.00962857
R15301 DVDD.n9186 DVDD.n514 0.00962857
R15302 DVDD.n9186 DVDD.n516 0.00962857
R15303 DVDD.n9182 DVDD.n516 0.00962857
R15304 DVDD.n9182 DVDD.n518 0.00962857
R15305 DVDD.n9178 DVDD.n518 0.00962857
R15306 DVDD.n9178 DVDD.n520 0.00962857
R15307 DVDD.n9129 DVDD.n520 0.00962857
R15308 DVDD.n9129 DVDD.n9127 0.00962857
R15309 DVDD.n9171 DVDD.n9127 0.00962857
R15310 DVDD.n9171 DVDD.n9128 0.00962857
R15311 DVDD.n9167 DVDD.n9128 0.00962857
R15312 DVDD.n9167 DVDD.n9133 0.00962857
R15313 DVDD.n9163 DVDD.n9133 0.00962857
R15314 DVDD.n9163 DVDD.n9136 0.00962857
R15315 DVDD.n9159 DVDD.n9136 0.00962857
R15316 DVDD.n9159 DVDD.n9138 0.00962857
R15317 DVDD.n9155 DVDD.n9138 0.00962857
R15318 DVDD.n9155 DVDD.n9140 0.00962857
R15319 DVDD.n9151 DVDD.n9140 0.00962857
R15320 DVDD.n9151 DVDD.n9142 0.00962857
R15321 DVDD.n9147 DVDD.n9142 0.00962857
R15322 DVDD.n9147 DVDD.n9144 0.00962857
R15323 DVDD.n9144 DVDD.n58 0.00962857
R15324 DVDD.n9649 DVDD.n58 0.00962857
R15325 DVDD.n9649 DVDD.n56 0.00962857
R15326 DVDD.n9653 DVDD.n56 0.00962857
R15327 DVDD.n9653 DVDD.n54 0.00962857
R15328 DVDD.n9657 DVDD.n54 0.00962857
R15329 DVDD.n9657 DVDD.n52 0.00962857
R15330 DVDD.n9661 DVDD.n52 0.00962857
R15331 DVDD.n9661 DVDD.n50 0.00962857
R15332 DVDD.n9665 DVDD.n50 0.00962857
R15333 DVDD.n9665 DVDD.n48 0.00962857
R15334 DVDD.n9669 DVDD.n48 0.00962857
R15335 DVDD.n9669 DVDD.n23 0.00962857
R15336 DVDD.n9676 DVDD.n23 0.00962857
R15337 DVDD.n9676 DVDD.n21 0.00962857
R15338 DVDD.n9680 DVDD.n21 0.00962857
R15339 DVDD.n9680 DVDD.n19 0.00962857
R15340 DVDD.n9684 DVDD.n19 0.00962857
R15341 DVDD.n9684 DVDD.n17 0.00962857
R15342 DVDD.n9689 DVDD.n17 0.00962857
R15343 DVDD.n9689 DVDD.n2 0.00962857
R15344 DVDD.n9695 DVDD.n2 0.00962857
R15345 DVDD.n9696 DVDD.n9695 0.00962857
R15346 DVDD.n3501 DVDD.n3500 0.00959285
R15347 DVDD.n6446 DVDD.n3501 0.00959285
R15348 DVDD.n6455 DVDD.n3485 0.00959285
R15349 DVDD.n6456 DVDD.n6455 0.00959285
R15350 DVDD.n5608 DVDD.n2535 0.00953543
R15351 DVDD.n5606 DVDD.n2537 0.00953543
R15352 DVDD.n5604 DVDD.n2534 0.00953543
R15353 DVDD.n5602 DVDD.n2538 0.00953543
R15354 DVDD.n5600 DVDD.n2533 0.00953543
R15355 DVDD.n5598 DVDD.n2539 0.00953543
R15356 DVDD.n5596 DVDD.n2532 0.00953543
R15357 DVDD.n5594 DVDD.n2540 0.00953543
R15358 DVDD.n5592 DVDD.n2531 0.00953543
R15359 DVDD.n5590 DVDD.n2541 0.00953543
R15360 DVDD.n5588 DVDD.n2530 0.00953543
R15361 DVDD.n5586 DVDD.n2542 0.00953543
R15362 DVDD.n5584 DVDD.n2529 0.00953543
R15363 DVDD.n5582 DVDD.n2543 0.00953543
R15364 DVDD.n5580 DVDD.n2528 0.00953543
R15365 DVDD.n2651 DVDD.n2545 0.00953543
R15366 DVDD.n6270 DVDD.n3343 0.00953543
R15367 DVDD.n6490 DVDD.n2089 0.00953543
R15368 DVDD.n5961 DVDD.n3232 0.00953543
R15369 DVDD.n3253 DVDD.n2137 0.00953543
R15370 DVDD.n5859 DVDD.n3108 0.00953543
R15371 DVDD.n3144 DVDD.n2186 0.00953543
R15372 DVDD.n6923 DVDD.n6922 0.00953543
R15373 DVDD.n6932 DVDD.n6931 0.00953543
R15374 DVDD.n6453 DVDD.n6451 0.00943276
R15375 DVDD.n8679 DVDD.n1044 0.009275
R15376 DVDD.n8732 DVDD.n881 0.009275
R15377 DVDD.n6316 DVDD.n3868 0.009275
R15378 DVDD.n6872 DVDD.n2791 0.009275
R15379 DVDD.n9584 DVDD.n9583 0.009275
R15380 DVDD.n2910 DVDD.n2900 0.009275
R15381 DVDD.n9350 DVDD.n9349 0.009275
R15382 DVDD.n8760 DVDD.n856 0.009275
R15383 DVDD.n5561 DVDD.n5560 0.0091811
R15384 DVDD.n5567 DVDD.n5500 0.0091811
R15385 DVDD.n5569 DVDD.n5562 0.0091811
R15386 DVDD.n5571 DVDD.n5499 0.0091811
R15387 DVDD.n5573 DVDD.n5563 0.0091811
R15388 DVDD.n5575 DVDD.n5498 0.0091811
R15389 DVDD.n5577 DVDD.n5564 0.0091811
R15390 DVDD.n5565 DVDD.n5497 0.0091811
R15391 DVDD.n5613 DVDD.n5612 0.0091811
R15392 DVDD.n711 DVDD.n578 0.0091811
R15393 DVDD.n8719 DVDD.n889 0.0091811
R15394 DVDD.n3832 DVDD.n3812 0.0091811
R15395 DVDD.n2433 DVDD.n1967 0.0091811
R15396 DVDD.n8987 DVDD.n8975 0.0091811
R15397 DVDD.n4073 DVDD.n4070 0.0091811
R15398 DVDD.n6036 DVDD.n3952 0.0091811
R15399 DVDD.n2436 DVDD.n2297 0.0091811
R15400 DVDD.n5020 DVDD.n4864 0.0091811
R15401 DVDD.n366 DVDD.n364 0.0091811
R15402 DVDD.n5803 DVDD.n4381 0.0091811
R15403 DVDD.n2442 DVDD.n2230 0.0091811
R15404 DVDD.n5131 DVDD.n5119 0.0091811
R15405 DVDD.n9399 DVDD.n9397 0.0091811
R15406 DVDD.n2863 DVDD.n2813 0.0091811
R15407 DVDD.n2427 DVDD.n2377 0.0091811
R15408 DVDD.n5529 DVDD.n5496 0.00893735
R15409 DVDD.n2550 DVDD.n2523 0.00893735
R15410 DVDD.n7522 DVDD.n7510 0.00893735
R15411 DVDD.n5415 DVDD.n4473 0.00893735
R15412 DVDD.n7211 DVDD.n7031 0.00891532
R15413 DVDD.n8771 DVDD.n92 0.00882677
R15414 DVDD.n3820 DVDD.n3809 0.00882677
R15415 DVDD.n6300 DVDD.n6299 0.00882677
R15416 DVDD.n6254 DVDD.n3348 0.00882677
R15417 DVDD.n4101 DVDD.n4002 0.00882677
R15418 DVDD.n6048 DVDD.n3949 0.00882677
R15419 DVDD.n5992 DVDD.n5929 0.00882677
R15420 DVDD.n5945 DVDD.n3234 0.00882677
R15421 DVDD.n9464 DVDD.n297 0.00882677
R15422 DVDD.n5815 DVDD.n4378 0.00882677
R15423 DVDD.n6096 DVDD.n5828 0.00882677
R15424 DVDD.n5843 DVDD.n3113 0.00882677
R15425 DVDD.n9360 DVDD.n410 0.00882677
R15426 DVDD.n2829 DVDD.n2810 0.00882677
R15427 DVDD.n6901 DVDD.n6900 0.00882677
R15428 DVDD.n6905 DVDD.n2664 0.00882677
R15429 DVDD.n3496 DVDD.n3487 0.00866435
R15430 DVDD.n3890 DVDD.n3887 0.0084875
R15431 DVDD.n6224 DVDD.n3890 0.0084875
R15432 DVDD.n6224 DVDD.n6223 0.0084875
R15433 DVDD.n6223 DVDD.n6222 0.0084875
R15434 DVDD.n6222 DVDD.n3891 0.0084875
R15435 DVDD.n6216 DVDD.n3891 0.0084875
R15436 DVDD.n6216 DVDD.n6215 0.0084875
R15437 DVDD.n6215 DVDD.n6214 0.0084875
R15438 DVDD.n6433 DVDD.n6432 0.0084875
R15439 DVDD.n6435 DVDD.n6433 0.0084875
R15440 DVDD.n6435 DVDD.n6434 0.0084875
R15441 DVDD.n6434 DVDD.n3468 0.0084875
R15442 DVDD.n6232 DVDD.n6231 0.0084875
R15443 DVDD.n6231 DVDD.n6229 0.0084875
R15444 DVDD.n6229 DVDD.n3886 0.0084875
R15445 DVDD.n6225 DVDD.n3886 0.0084875
R15446 DVDD.n6225 DVDD.n3889 0.0084875
R15447 DVDD.n6221 DVDD.n3889 0.0084875
R15448 DVDD.n6221 DVDD.n3892 0.0084875
R15449 DVDD.n6217 DVDD.n3892 0.0084875
R15450 DVDD.n6217 DVDD.n6213 0.0084875
R15451 DVDD.n6213 DVDD.n3509 0.0084875
R15452 DVDD.n6427 DVDD.n6425 0.0084875
R15453 DVDD.n6427 DVDD.n3507 0.0084875
R15454 DVDD.n6431 DVDD.n3507 0.0084875
R15455 DVDD.n6431 DVDD.n3505 0.0084875
R15456 DVDD.n6436 DVDD.n3505 0.0084875
R15457 DVDD.n6436 DVDD.n3503 0.0084875
R15458 DVDD.n6440 DVDD.n3503 0.0084875
R15459 DVDD.n6441 DVDD.n6440 0.0084875
R15460 DVDD.n6443 DVDD.n6441 0.0084875
R15461 DVDD.n6080 DVDD.n5911 0.0084875
R15462 DVDD.n6076 DVDD.n5911 0.0084875
R15463 DVDD.n6076 DVDD.n5914 0.0084875
R15464 DVDD.n6072 DVDD.n5914 0.0084875
R15465 DVDD.n6072 DVDD.n5916 0.0084875
R15466 DVDD.n6068 DVDD.n5916 0.0084875
R15467 DVDD.n6068 DVDD.n5918 0.0084875
R15468 DVDD.n6064 DVDD.n5918 0.0084875
R15469 DVDD.n6064 DVDD.n5920 0.0084875
R15470 DVDD.n5994 DVDD.n5920 0.0084875
R15471 DVDD.n3942 DVDD.n3916 0.0084875
R15472 DVDD.n3938 DVDD.n3916 0.0084875
R15473 DVDD.n3938 DVDD.n3918 0.0084875
R15474 DVDD.n3934 DVDD.n3918 0.0084875
R15475 DVDD.n3934 DVDD.n3920 0.0084875
R15476 DVDD.n3930 DVDD.n3920 0.0084875
R15477 DVDD.n3930 DVDD.n3922 0.0084875
R15478 DVDD.n3926 DVDD.n3922 0.0084875
R15479 DVDD.n3926 DVDD.n3923 0.0084875
R15480 DVDD.n6079 DVDD.n6078 0.0084875
R15481 DVDD.n6078 DVDD.n6077 0.0084875
R15482 DVDD.n6077 DVDD.n5913 0.0084875
R15483 DVDD.n6071 DVDD.n5913 0.0084875
R15484 DVDD.n6071 DVDD.n6070 0.0084875
R15485 DVDD.n6070 DVDD.n6069 0.0084875
R15486 DVDD.n3941 DVDD.n3940 0.0084875
R15487 DVDD.n3940 DVDD.n3939 0.0084875
R15488 DVDD.n3939 DVDD.n3917 0.0084875
R15489 DVDD.n3933 DVDD.n3917 0.0084875
R15490 DVDD.n3933 DVDD.n3932 0.0084875
R15491 DVDD.n3932 DVDD.n3931 0.0084875
R15492 DVDD.n3931 DVDD.n3921 0.0084875
R15493 DVDD.n3925 DVDD.n3921 0.0084875
R15494 DVDD.n3925 DVDD.n3924 0.0084875
R15495 DVDD.n4408 DVDD.n4404 0.0084875
R15496 DVDD.n4409 DVDD.n4408 0.0084875
R15497 DVDD.n4410 DVDD.n4409 0.0084875
R15498 DVDD.n4410 DVDD.n4400 0.0084875
R15499 DVDD.n4416 DVDD.n4400 0.0084875
R15500 DVDD.n4417 DVDD.n4416 0.0084875
R15501 DVDD.n4419 DVDD.n4417 0.0084875
R15502 DVDD.n4419 DVDD.n4418 0.0084875
R15503 DVDD.n4418 DVDD.n4396 0.0084875
R15504 DVDD.n4426 DVDD.n4396 0.0084875
R15505 DVDD.n6094 DVDD.n5896 0.0084875
R15506 DVDD.n6088 DVDD.n5896 0.0084875
R15507 DVDD.n6088 DVDD.n6087 0.0084875
R15508 DVDD.n6087 DVDD.n6086 0.0084875
R15509 DVDD.n6086 DVDD.n5905 0.0084875
R15510 DVDD.n4407 DVDD.n4405 0.0084875
R15511 DVDD.n4407 DVDD.n4403 0.0084875
R15512 DVDD.n4411 DVDD.n4403 0.0084875
R15513 DVDD.n4411 DVDD.n4401 0.0084875
R15514 DVDD.n4415 DVDD.n4401 0.0084875
R15515 DVDD.n4415 DVDD.n4399 0.0084875
R15516 DVDD.n4420 DVDD.n4399 0.0084875
R15517 DVDD.n4420 DVDD.n4397 0.0084875
R15518 DVDD.n4424 DVDD.n4397 0.0084875
R15519 DVDD.n4425 DVDD.n4424 0.0084875
R15520 DVDD.n6099 DVDD.n4395 0.0084875
R15521 DVDD.n5900 DVDD.n4395 0.0084875
R15522 DVDD.n5900 DVDD.n5897 0.0084875
R15523 DVDD.n6093 DVDD.n5897 0.0084875
R15524 DVDD.n6093 DVDD.n5898 0.0084875
R15525 DVDD.n6089 DVDD.n5898 0.0084875
R15526 DVDD.n6089 DVDD.n5904 0.0084875
R15527 DVDD.n6085 DVDD.n5904 0.0084875
R15528 DVDD.n6085 DVDD.n5906 0.0084875
R15529 DVDD.n5649 DVDD.n4458 0.0084875
R15530 DVDD.n5661 DVDD.n4458 0.0084875
R15531 DVDD.n5661 DVDD.n4456 0.0084875
R15532 DVDD.n5666 DVDD.n4456 0.0084875
R15533 DVDD.n5666 DVDD.n4453 0.0084875
R15534 DVDD.n5670 DVDD.n4453 0.0084875
R15535 DVDD.n5671 DVDD.n5670 0.0084875
R15536 DVDD.n5672 DVDD.n5671 0.0084875
R15537 DVDD.n5672 DVDD.n4451 0.0084875
R15538 DVDD.n5679 DVDD.n4451 0.0084875
R15539 DVDD.n5708 DVDD.n5680 0.0084875
R15540 DVDD.n5704 DVDD.n5680 0.0084875
R15541 DVDD.n5704 DVDD.n5683 0.0084875
R15542 DVDD.n5700 DVDD.n5683 0.0084875
R15543 DVDD.n5700 DVDD.n5686 0.0084875
R15544 DVDD.n5696 DVDD.n5686 0.0084875
R15545 DVDD.n5696 DVDD.n5688 0.0084875
R15546 DVDD.n5692 DVDD.n5688 0.0084875
R15547 DVDD.n5692 DVDD.n5690 0.0084875
R15548 DVDD.n5667 DVDD.n4455 0.0084875
R15549 DVDD.n5668 DVDD.n5667 0.0084875
R15550 DVDD.n5669 DVDD.n5668 0.0084875
R15551 DVDD.n5669 DVDD.n3002 0.0084875
R15552 DVDD.n5707 DVDD.n5706 0.0084875
R15553 DVDD.n5706 DVDD.n5705 0.0084875
R15554 DVDD.n5705 DVDD.n5682 0.0084875
R15555 DVDD.n5699 DVDD.n5682 0.0084875
R15556 DVDD.n5699 DVDD.n5698 0.0084875
R15557 DVDD.n5698 DVDD.n5697 0.0084875
R15558 DVDD.n5697 DVDD.n5687 0.0084875
R15559 DVDD.n5691 DVDD.n5687 0.0084875
R15560 DVDD.n8767 DVDD.n114 0.00847244
R15561 DVDD.n6336 DVDD.n6335 0.00847244
R15562 DVDD.n6258 DVDD.n3340 0.00847244
R15563 DVDD.n2410 DVDD.n1976 0.00847244
R15564 DVDD.n4097 DVDD.n112 0.00847244
R15565 DVDD.n6052 DVDD.n3968 0.00847244
R15566 DVDD.n5949 DVDD.n3220 0.00847244
R15567 DVDD.n2413 DVDD.n2298 0.00847244
R15568 DVDD.n9459 DVDD.n125 0.00847244
R15569 DVDD.n5819 DVDD.n4315 0.00847244
R15570 DVDD.n5847 DVDD.n3105 0.00847244
R15571 DVDD.n2419 DVDD.n2239 0.00847244
R15572 DVDD.n131 DVDD.n126 0.00847244
R15573 DVDD.n6858 DVDD.n6857 0.00847244
R15574 DVDD.n6909 DVDD.n2734 0.00847244
R15575 DVDD.n2404 DVDD.n2378 0.00847244
R15576 DVDD.n6398 DVDD.n6386 0.00838454
R15577 DVDD.n6374 DVDD.n3536 0.00821966
R15578 DVDD.n6372 DVDD.n3531 0.00821966
R15579 DVDD.n6370 DVDD.n3537 0.00821966
R15580 DVDD.n6368 DVDD.n3530 0.00821966
R15581 DVDD.n6366 DVDD.n3538 0.00821966
R15582 DVDD.n6364 DVDD.n3529 0.00821966
R15583 DVDD.n6362 DVDD.n3539 0.00821966
R15584 DVDD.n6360 DVDD.n3528 0.00821966
R15585 DVDD.n6358 DVDD.n3540 0.00821966
R15586 DVDD.n6356 DVDD.n3527 0.00821966
R15587 DVDD.n6354 DVDD.n3541 0.00821966
R15588 DVDD.n6352 DVDD.n3526 0.00821966
R15589 DVDD.n6350 DVDD.n3542 0.00821966
R15590 DVDD.n6348 DVDD.n3525 0.00821966
R15591 DVDD.n6346 DVDD.n3543 0.00821966
R15592 DVDD.n6344 DVDD.n3524 0.00821966
R15593 DVDD.n6342 DVDD.n3544 0.00821966
R15594 DVDD.n6340 DVDD.n3523 0.00821966
R15595 DVDD.n6338 DVDD.n3545 0.00821966
R15596 DVDD.n3546 DVDD.n3522 0.00821966
R15597 DVDD.n715 DVDD.n584 0.00811811
R15598 DVDD.n8723 DVDD.n356 0.00811811
R15599 DVDD.n3640 DVDD.n1050 0.00811811
R15600 DVDD.n3836 DVDD.n3567 0.00811811
R15601 DVDD.n6520 DVDD.n2082 0.00811811
R15602 DVDD.n1885 DVDD.n1866 0.00811811
R15603 DVDD.n8983 DVDD.n556 0.00811811
R15604 DVDD.n4077 DVDD.n372 0.00811811
R15605 DVDD.n4205 DVDD.n4155 0.00811811
R15606 DVDD.n6032 DVDD.n3964 0.00811811
R15607 DVDD.n3283 DVDD.n2121 0.00811811
R15608 DVDD.n8291 DVDD.n1677 0.00811811
R15609 DVDD.n5024 DVDD.n4861 0.00811811
R15610 DVDD.n370 DVDD.n345 0.00811811
R15611 DVDD.n9546 DVDD.n250 0.00811811
R15612 DVDD.n5799 DVDD.n4311 0.00811811
R15613 DVDD.n3174 DVDD.n2179 0.00811811
R15614 DVDD.n1874 DVDD.n1601 0.00811811
R15615 DVDD.n5127 DVDD.n4578 0.00811811
R15616 DVDD.n9393 DVDD.n375 0.00811811
R15617 DVDD.n6778 DVDD.n2905 0.00811811
R15618 DVDD.n2859 DVDD.n2826 0.00811811
R15619 DVDD.n2704 DVDD.n2646 0.00811811
R15620 DVDD.n8357 DVDD.n1561 0.00811811
R15621 DVDD.n7710 DVDD.n1887 0.00794094
R15622 DVDD.n7703 DVDD.n1669 0.00794094
R15623 DVDD.n7697 DVDD.n1605 0.00794094
R15624 DVDD.n7690 DVDD.n1550 0.00794094
R15625 DVDD.n6465 DVDD.n3466 0.00789805
R15626 DVDD.n6466 DVDD.n3419 0.0078431
R15627 DVDD DVDD.n640 0.00782857
R15628 DVDD.n8200 DVDD 0.00782857
R15629 DVDD DVDD.n0 0.00782857
R15630 DVDD.n9696 DVDD 0.00782857
R15631 DVDD.n5422 DVDD.n5421 0.00776378
R15632 DVDD.n5431 DVDD.n4482 0.00776378
R15633 DVDD.n5433 DVDD.n5423 0.00776378
R15634 DVDD.n5435 DVDD.n4481 0.00776378
R15635 DVDD.n5437 DVDD.n5424 0.00776378
R15636 DVDD.n5439 DVDD.n4480 0.00776378
R15637 DVDD.n5441 DVDD.n5425 0.00776378
R15638 DVDD.n5443 DVDD.n4479 0.00776378
R15639 DVDD.n5445 DVDD.n5426 0.00776378
R15640 DVDD.n5447 DVDD.n4478 0.00776378
R15641 DVDD.n5449 DVDD.n5427 0.00776378
R15642 DVDD.n5451 DVDD.n4477 0.00776378
R15643 DVDD.n5453 DVDD.n5428 0.00776378
R15644 DVDD.n5455 DVDD.n4476 0.00776378
R15645 DVDD.n5457 DVDD.n5429 0.00776378
R15646 DVDD.n5459 DVDD.n4475 0.00776378
R15647 DVDD.n5461 DVDD.n5430 0.00776378
R15648 DVDD.n5464 DVDD.n4474 0.00776378
R15649 DVDD.n5465 DVDD.n4469 0.00776378
R15650 DVDD.n5468 DVDD.n5467 0.00776378
R15651 DVDD.n5471 DVDD.n4467 0.00776378
R15652 DVDD.n6649 DVDD.n3356 0.00776378
R15653 DVDD.n6494 DVDD.n2076 0.00776378
R15654 DVDD.n3290 DVDD.n3226 0.00776378
R15655 DVDD.n3257 DVDD.n2127 0.00776378
R15656 DVDD.n6705 DVDD.n3121 0.00776378
R15657 DVDD.n3148 DVDD.n2173 0.00776378
R15658 DVDD.n2711 DVDD.n2671 0.00776378
R15659 DVDD.n2678 DVDD.n2637 0.00776378
R15660 DVDD.n8172 DVDD.n8171 0.00772462
R15661 DVDD.n6600 DVDD.n6599 0.00772462
R15662 DVDD.n7947 DVDD.n7946 0.00772462
R15663 DVDD.n8005 DVDD.n8004 0.00772462
R15664 DVDD.n6394 DVDD.n6393 0.00772462
R15665 DVDD.n6458 DVDD.n6457 0.00771783
R15666 DVDD.n3491 DVDD.n3490 0.00771783
R15667 DVDD.n9425 DVDD.n355 0.00770384
R15668 DVDD.n354 DVDD.n200 0.00770384
R15669 DVDD.n5690 DVDD.n2786 0.0077
R15670 DVDD.n7488 DVDD.n7487 0.00763571
R15671 DVDD.n8369 DVDD.n1514 0.00763571
R15672 DVDD.n7333 DVDD.n7329 0.00763571
R15673 DVDD.n4819 DVDD.n4600 0.00763571
R15674 DVDD.n5157 DVDD.n4574 0.00763571
R15675 DVDD.n5083 DVDD.n5082 0.00763571
R15676 DVDD.n4787 DVDD.n4773 0.00763571
R15677 DVDD.n9284 DVDD.n460 0.00763571
R15678 DVDD.n9211 DVDD.n9210 0.00763571
R15679 DVDD.n8689 DVDD.n1006 0.007475
R15680 DVDD.n8713 DVDD.n897 0.007475
R15681 DVDD.n6308 DVDD.n3879 0.007475
R15682 DVDD.n6886 DVDD.n2782 0.007475
R15683 DVDD.n9402 DVDD.n9401 0.007475
R15684 DVDD.n5282 DVDD.n5281 0.007475
R15685 DVDD.n9358 DVDD.n412 0.007475
R15686 DVDD.n9621 DVDD.n9620 0.007475
R15687 DVDD.n5641 DVDD.n5481 0.00740945
R15688 DVDD.n5658 DVDD.n5639 0.00740945
R15689 DVDD.n8812 DVDD.n68 0.00740945
R15690 DVDD.n3852 DVDD.n3816 0.00740945
R15691 DVDD.n6536 DVDD.n3334 0.00740945
R15692 DVDD.n6504 DVDD.n2086 0.00740945
R15693 DVDD.n9084 DVDD.n528 0.00740945
R15694 DVDD.n6016 DVDD.n3956 0.00740945
R15695 DVDD.n3242 DVDD.n3235 0.00740945
R15696 DVDD.n3267 DVDD.n2140 0.00740945
R15697 DVDD.n4927 DVDD.n492 0.00740945
R15698 DVDD.n5783 DVDD.n4385 0.00740945
R15699 DVDD.n3133 DVDD.n3099 0.00740945
R15700 DVDD.n3158 DVDD.n2183 0.00740945
R15701 DVDD.n9257 DVDD.n9245 0.00740945
R15702 DVDD.n2843 DVDD.n2817 0.00740945
R15703 DVDD.n2723 DVDD.n2722 0.00740945
R15704 DVDD.n2688 DVDD.n2632 0.00740945
R15705 DVDD.n8277 DVDD.n1703 0.00737857
R15706 DVDD.n1769 DVDD.n1763 0.00737857
R15707 DVDD.n1779 DVDD.n1272 0.00737857
R15708 DVDD.n8963 DVDD.n548 0.00737857
R15709 DVDD.n8936 DVDD.n8935 0.00737857
R15710 DVDD.n8910 DVDD.n8909 0.00737857
R15711 DVDD.n9134 DVDD.n533 0.00737857
R15712 DVDD.n9654 DVDD.n55 0.00737857
R15713 DVDD.n9681 DVDD.n20 0.00737857
R15714 DVDD.n5912 DVDD.n5905 0.00725
R15715 DVDD.n5910 DVDD.n5906 0.00725
R15716 DVDD.n3749 DVDD.n1013 0.00725
R15717 DVDD.n3748 DVDD.n3747 0.00725
R15718 DVDD.n3744 DVDD.n1039 0.00725
R15719 DVDD.n3743 DVDD.n3584 0.00725
R15720 DVDD.n3633 DVDD.n3632 0.00725
R15721 DVDD.n3629 DVDD.n1053 0.00725
R15722 DVDD.n3628 DVDD.n3627 0.00725
R15723 DVDD.n6425 DVDD.n6424 0.0071375
R15724 DVDD.n326 DVDD.n325 0.0071
R15725 DVDD.n9341 DVDD.n9331 0.0071
R15726 DVDD.n4086 DVDD.n4020 0.0071
R15727 DVDD.n968 DVDD.n967 0.0071
R15728 DVDD.n8806 DVDD.n69 0.00705512
R15729 DVDD.n8748 DVDD.n874 0.00705512
R15730 DVDD.n1041 DVDD.n1040 0.00705512
R15731 DVDD.n3846 DVDD.n3815 0.00705512
R15732 DVDD.n6324 DVDD.n6323 0.00705512
R15733 DVDD.n6542 DVDD.n3335 0.00705512
R15734 DVDD.n6510 DVDD.n2085 0.00705512
R15735 DVDD.n1983 DVDD.n1949 0.00705512
R15736 DVDD.n9078 DVDD.n531 0.00705512
R15737 DVDD.n4057 DVDD.n4032 0.00705512
R15738 DVDD.n4218 DVDD.n4217 0.00705512
R15739 DVDD.n6022 DVDD.n3955 0.00705512
R15740 DVDD.n6057 DVDD.n5923 0.00705512
R15741 DVDD.n3248 DVDD.n3224 0.00705512
R15742 DVDD.n3273 DVDD.n2141 0.00705512
R15743 DVDD.n7748 DVDD.n2293 0.00705512
R15744 DVDD.n4921 DVDD.n493 0.00705512
R15745 DVDD.n340 DVDD.n338 0.00705512
R15746 DVDD.n9509 DVDD.n9508 0.00705512
R15747 DVDD.n5789 DVDD.n4384 0.00705512
R15748 DVDD.n5767 DVDD.n5764 0.00705512
R15749 DVDD.n3139 DVDD.n3100 0.00705512
R15750 DVDD.n3164 DVDD.n2182 0.00705512
R15751 DVDD.n2246 DVDD.n2212 0.00705512
R15752 DVDD.n9263 DVDD.n9248 0.00705512
R15753 DVDD.n9595 DVDD.n9594 0.00705512
R15754 DVDD.n6794 DVDD.n6793 0.00705512
R15755 DVDD.n2849 DVDD.n2816 0.00705512
R15756 DVDD.n6862 DVDD.n2798 0.00705512
R15757 DVDD.n6926 DVDD.n6925 0.00705512
R15758 DVDD.n2694 DVDD.n2635 0.00705512
R15759 DVDD.n7678 DVDD.n7677 0.00705512
R15760 DVDD.n9694 DVDD.n9693 0.00699286
R15761 DVDD.n6449 DVDD.n6448 0.00693543
R15762 DVDD.n6447 DVDD.n3489 0.00693543
R15763 DVDD.n3923 DVDD.n3884 0.0068
R15764 DVDD.n3924 DVDD.n3876 0.0068
R15765 DVDD.n9488 DVDD.n270 0.00678
R15766 DVDD.n9572 DVDD.n205 0.00678
R15767 DVDD.n4128 DVDD.n3979 0.00678
R15768 DVDD.n1026 DVDD.n1016 0.00678
R15769 DVDD.n6098 DVDD.n6097 0.00674375
R15770 DVDD.n6771 DVDD.n3002 0.00674375
R15771 DVDD.n5691 DVDD.n2743 0.00674375
R15772 DVDD.n933 DVDD.n865 0.00670079
R15773 DVDD.n6268 DVDD.n3345 0.00670079
R15774 DVDD.n6488 DVDD.n2075 0.00670079
R15775 DVDD.n4048 DVDD.n4034 0.00670079
R15776 DVDD.n5959 DVDD.n3218 0.00670079
R15777 DVDD.n3251 DVDD.n2128 0.00670079
R15778 DVDD.n9447 DVDD.n9446 0.00670079
R15779 DVDD.n5857 DVDD.n3110 0.00670079
R15780 DVDD.n3142 DVDD.n2172 0.00670079
R15781 DVDD.n9600 DVDD.n142 0.00670079
R15782 DVDD.n6919 DVDD.n2661 0.00670079
R15783 DVDD.n6928 DVDD.n2630 0.00670079
R15784 DVDD.n3942 DVDD.n3913 0.0066875
R15785 DVDD.n3941 DVDD.n3912 0.0066875
R15786 DVDD.n4761 DVDD.n4760 0.00658571
R15787 DVDD.n4761 DVDD.n4755 0.00658571
R15788 DVDD.n4767 DVDD.n4755 0.00658571
R15789 DVDD.n4768 DVDD.n4767 0.00658571
R15790 DVDD.n4770 DVDD.n4768 0.00658571
R15791 DVDD.n4770 DVDD.n4769 0.00658571
R15792 DVDD.n4769 DVDD.n4751 0.00658571
R15793 DVDD.n4792 DVDD.n4751 0.00658571
R15794 DVDD.n4793 DVDD.n4792 0.00658571
R15795 DVDD.n4813 DVDD.n4793 0.00658571
R15796 DVDD.n4813 DVDD.n4812 0.00658571
R15797 DVDD.n4812 DVDD.n4811 0.00658571
R15798 DVDD.n4811 DVDD.n4794 0.00658571
R15799 DVDD.n4805 DVDD.n4794 0.00658571
R15800 DVDD.n4805 DVDD.n4804 0.00658571
R15801 DVDD.n4804 DVDD.n4803 0.00658571
R15802 DVDD.n4803 DVDD.n4798 0.00658571
R15803 DVDD.n4798 DVDD.n468 0.00658571
R15804 DVDD.n9241 DVDD.n468 0.00658571
R15805 DVDD.n9241 DVDD.n9240 0.00658571
R15806 DVDD.n9240 DVDD.n9239 0.00658571
R15807 DVDD.n9239 DVDD.n469 0.00658571
R15808 DVDD.n473 DVDD.n469 0.00658571
R15809 DVDD.n9231 DVDD.n473 0.00658571
R15810 DVDD.n9231 DVDD.n9230 0.00658571
R15811 DVDD.n9230 DVDD.n9229 0.00658571
R15812 DVDD.n9229 DVDD.n474 0.00658571
R15813 DVDD.n9223 DVDD.n474 0.00658571
R15814 DVDD.n9223 DVDD.n9222 0.00658571
R15815 DVDD.n9222 DVDD.n9221 0.00658571
R15816 DVDD.n9221 DVDD.n478 0.00658571
R15817 DVDD.n9215 DVDD.n478 0.00658571
R15818 DVDD.n9215 DVDD.n9214 0.00658571
R15819 DVDD.n9214 DVDD.n9213 0.00658571
R15820 DVDD.n9213 DVDD.n482 0.00658571
R15821 DVDD.n505 DVDD.n482 0.00658571
R15822 DVDD.n506 DVDD.n505 0.00658571
R15823 DVDD.n9205 DVDD.n506 0.00658571
R15824 DVDD.n9205 DVDD.n9204 0.00658571
R15825 DVDD.n9204 DVDD.n9203 0.00658571
R15826 DVDD.n9203 DVDD.n507 0.00658571
R15827 DVDD.n9197 DVDD.n507 0.00658571
R15828 DVDD.n9197 DVDD.n9196 0.00658571
R15829 DVDD.n9196 DVDD.n9195 0.00658571
R15830 DVDD.n9195 DVDD.n511 0.00658571
R15831 DVDD.n9189 DVDD.n511 0.00658571
R15832 DVDD.n9189 DVDD.n9188 0.00658571
R15833 DVDD.n9188 DVDD.n9187 0.00658571
R15834 DVDD.n9187 DVDD.n515 0.00658571
R15835 DVDD.n9181 DVDD.n515 0.00658571
R15836 DVDD.n9181 DVDD.n9180 0.00658571
R15837 DVDD.n9180 DVDD.n9179 0.00658571
R15838 DVDD.n9179 DVDD.n519 0.00658571
R15839 DVDD.n9130 DVDD.n519 0.00658571
R15840 DVDD.n9131 DVDD.n9130 0.00658571
R15841 DVDD.n9170 DVDD.n9131 0.00658571
R15842 DVDD.n9170 DVDD.n9169 0.00658571
R15843 DVDD.n9169 DVDD.n9168 0.00658571
R15844 DVDD.n9168 DVDD.n9132 0.00658571
R15845 DVDD.n9162 DVDD.n9132 0.00658571
R15846 DVDD.n9162 DVDD.n9161 0.00658571
R15847 DVDD.n9161 DVDD.n9160 0.00658571
R15848 DVDD.n9160 DVDD.n9137 0.00658571
R15849 DVDD.n9154 DVDD.n9137 0.00658571
R15850 DVDD.n9154 DVDD.n9153 0.00658571
R15851 DVDD.n9153 DVDD.n9152 0.00658571
R15852 DVDD.n9152 DVDD.n9141 0.00658571
R15853 DVDD.n9146 DVDD.n9141 0.00658571
R15854 DVDD.n9146 DVDD.n9145 0.00658571
R15855 DVDD.n9145 DVDD.n57 0.00658571
R15856 DVDD.n9650 DVDD.n57 0.00658571
R15857 DVDD.n9651 DVDD.n9650 0.00658571
R15858 DVDD.n9652 DVDD.n9651 0.00658571
R15859 DVDD.n9652 DVDD.n53 0.00658571
R15860 DVDD.n9658 DVDD.n53 0.00658571
R15861 DVDD.n9659 DVDD.n9658 0.00658571
R15862 DVDD.n9660 DVDD.n9659 0.00658571
R15863 DVDD.n9660 DVDD.n49 0.00658571
R15864 DVDD.n9666 DVDD.n49 0.00658571
R15865 DVDD.n9667 DVDD.n9666 0.00658571
R15866 DVDD.n9668 DVDD.n9667 0.00658571
R15867 DVDD.n9668 DVDD.n22 0.00658571
R15868 DVDD.n9677 DVDD.n22 0.00658571
R15869 DVDD.n9678 DVDD.n9677 0.00658571
R15870 DVDD.n9679 DVDD.n9678 0.00658571
R15871 DVDD.n9679 DVDD.n18 0.00658571
R15872 DVDD.n9685 DVDD.n18 0.00658571
R15873 DVDD.n9686 DVDD.n9685 0.00658571
R15874 DVDD.n9688 DVDD.n9686 0.00658571
R15875 DVDD.n9688 DVDD.n9687 0.00658571
R15876 DVDD.n9687 DVDD.n1 0.00658571
R15877 DVDD.n9697 DVDD.n1 0.00658571
R15878 DVDD.n9698 DVDD.n9697 0.00658571
R15879 DVDD.n4716 DVDD.n4611 0.00658571
R15880 DVDD.n4717 DVDD.n4716 0.00658571
R15881 DVDD.n4718 DVDD.n4717 0.00658571
R15882 DVDD.n4718 DVDD.n4607 0.00658571
R15883 DVDD.n4724 DVDD.n4607 0.00658571
R15884 DVDD.n4725 DVDD.n4724 0.00658571
R15885 DVDD.n4726 DVDD.n4725 0.00658571
R15886 DVDD.n4726 DVDD.n4591 0.00658571
R15887 DVDD.n4824 DVDD.n4591 0.00658571
R15888 DVDD.n4825 DVDD.n4824 0.00658571
R15889 DVDD.n4826 DVDD.n4825 0.00658571
R15890 DVDD.n4826 DVDD.n4587 0.00658571
R15891 DVDD.n4832 DVDD.n4587 0.00658571
R15892 DVDD.n4833 DVDD.n4832 0.00658571
R15893 DVDD.n4834 DVDD.n4833 0.00658571
R15894 DVDD.n4834 DVDD.n4583 0.00658571
R15895 DVDD.n4840 DVDD.n4583 0.00658571
R15896 DVDD.n4841 DVDD.n4840 0.00658571
R15897 DVDD.n5113 DVDD.n4841 0.00658571
R15898 DVDD.n5113 DVDD.n5112 0.00658571
R15899 DVDD.n5112 DVDD.n5111 0.00658571
R15900 DVDD.n5111 DVDD.n4842 0.00658571
R15901 DVDD.n4846 DVDD.n4842 0.00658571
R15902 DVDD.n5103 DVDD.n4846 0.00658571
R15903 DVDD.n5103 DVDD.n5102 0.00658571
R15904 DVDD.n5102 DVDD.n5101 0.00658571
R15905 DVDD.n5101 DVDD.n4847 0.00658571
R15906 DVDD.n5095 DVDD.n4847 0.00658571
R15907 DVDD.n5095 DVDD.n5094 0.00658571
R15908 DVDD.n5094 DVDD.n5093 0.00658571
R15909 DVDD.n5093 DVDD.n4851 0.00658571
R15910 DVDD.n5087 DVDD.n4851 0.00658571
R15911 DVDD.n5087 DVDD.n5086 0.00658571
R15912 DVDD.n5086 DVDD.n5085 0.00658571
R15913 DVDD.n5085 DVDD.n4855 0.00658571
R15914 DVDD.n5035 DVDD.n4855 0.00658571
R15915 DVDD.n5036 DVDD.n5035 0.00658571
R15916 DVDD.n5077 DVDD.n5036 0.00658571
R15917 DVDD.n5077 DVDD.n5076 0.00658571
R15918 DVDD.n5076 DVDD.n5075 0.00658571
R15919 DVDD.n5075 DVDD.n5037 0.00658571
R15920 DVDD.n5069 DVDD.n5037 0.00658571
R15921 DVDD.n5069 DVDD.n5068 0.00658571
R15922 DVDD.n5068 DVDD.n5067 0.00658571
R15923 DVDD.n5067 DVDD.n5041 0.00658571
R15924 DVDD.n5061 DVDD.n5041 0.00658571
R15925 DVDD.n5061 DVDD.n5060 0.00658571
R15926 DVDD.n5060 DVDD.n5059 0.00658571
R15927 DVDD.n5059 DVDD.n5045 0.00658571
R15928 DVDD.n5053 DVDD.n5045 0.00658571
R15929 DVDD.n5053 DVDD.n5052 0.00658571
R15930 DVDD.n5052 DVDD.n5051 0.00658571
R15931 DVDD.n5051 DVDD.n561 0.00658571
R15932 DVDD.n8969 DVDD.n561 0.00658571
R15933 DVDD.n8969 DVDD.n8968 0.00658571
R15934 DVDD.n8968 DVDD.n8967 0.00658571
R15935 DVDD.n8967 DVDD.n562 0.00658571
R15936 DVDD.n566 DVDD.n562 0.00658571
R15937 DVDD.n8959 DVDD.n566 0.00658571
R15938 DVDD.n8959 DVDD.n8958 0.00658571
R15939 DVDD.n8958 DVDD.n8957 0.00658571
R15940 DVDD.n8957 DVDD.n567 0.00658571
R15941 DVDD.n8951 DVDD.n567 0.00658571
R15942 DVDD.n8951 DVDD.n8950 0.00658571
R15943 DVDD.n8950 DVDD.n8949 0.00658571
R15944 DVDD.n8949 DVDD.n571 0.00658571
R15945 DVDD.n8943 DVDD.n571 0.00658571
R15946 DVDD.n8943 DVDD.n8942 0.00658571
R15947 DVDD.n8942 DVDD.n8941 0.00658571
R15948 DVDD.n8941 DVDD.n575 0.00658571
R15949 DVDD.n598 DVDD.n575 0.00658571
R15950 DVDD.n599 DVDD.n598 0.00658571
R15951 DVDD.n8933 DVDD.n599 0.00658571
R15952 DVDD.n8933 DVDD.n8932 0.00658571
R15953 DVDD.n8932 DVDD.n8931 0.00658571
R15954 DVDD.n8931 DVDD.n600 0.00658571
R15955 DVDD.n8925 DVDD.n600 0.00658571
R15956 DVDD.n8925 DVDD.n8924 0.00658571
R15957 DVDD.n8924 DVDD.n8923 0.00658571
R15958 DVDD.n8923 DVDD.n604 0.00658571
R15959 DVDD.n8917 DVDD.n604 0.00658571
R15960 DVDD.n8917 DVDD.n8916 0.00658571
R15961 DVDD.n8916 DVDD.n8915 0.00658571
R15962 DVDD.n8915 DVDD.n608 0.00658571
R15963 DVDD.n8907 DVDD.n608 0.00658571
R15964 DVDD.n8907 DVDD.n8906 0.00658571
R15965 DVDD.n8906 DVDD.n8905 0.00658571
R15966 DVDD.n8905 DVDD.n635 0.00658571
R15967 DVDD.n8899 DVDD.n635 0.00658571
R15968 DVDD.n8899 DVDD.n8898 0.00658571
R15969 DVDD.n8898 DVDD.n8897 0.00658571
R15970 DVDD.n8897 DVDD.n639 0.00658571
R15971 DVDD.n8890 DVDD.n639 0.00658571
R15972 DVDD.n7500 DVDD.n7499 0.00658571
R15973 DVDD.n7499 DVDD.n7498 0.00658571
R15974 DVDD.n7498 DVDD.n7093 0.00658571
R15975 DVDD.n7492 DVDD.n7093 0.00658571
R15976 DVDD.n7492 DVDD.n7491 0.00658571
R15977 DVDD.n7491 DVDD.n7490 0.00658571
R15978 DVDD.n7490 DVDD.n7097 0.00658571
R15979 DVDD.n7307 DVDD.n7097 0.00658571
R15980 DVDD.n7482 DVDD.n7307 0.00658571
R15981 DVDD.n7482 DVDD.n7481 0.00658571
R15982 DVDD.n7481 DVDD.n7480 0.00658571
R15983 DVDD.n7480 DVDD.n7308 0.00658571
R15984 DVDD.n7474 DVDD.n7308 0.00658571
R15985 DVDD.n7474 DVDD.n7473 0.00658571
R15986 DVDD.n7473 DVDD.n7472 0.00658571
R15987 DVDD.n7472 DVDD.n7313 0.00658571
R15988 DVDD.n7466 DVDD.n7313 0.00658571
R15989 DVDD.n7466 DVDD.n7465 0.00658571
R15990 DVDD.n7465 DVDD.n7464 0.00658571
R15991 DVDD.n7464 DVDD.n7316 0.00658571
R15992 DVDD.n7459 DVDD.n7316 0.00658571
R15993 DVDD.n7459 DVDD.n7458 0.00658571
R15994 DVDD.n7458 DVDD.n7457 0.00658571
R15995 DVDD.n7457 DVDD.n7318 0.00658571
R15996 DVDD.n7451 DVDD.n7318 0.00658571
R15997 DVDD.n7451 DVDD.n7450 0.00658571
R15998 DVDD.n7450 DVDD.n7449 0.00658571
R15999 DVDD.n7449 DVDD.n7323 0.00658571
R16000 DVDD.n7443 DVDD.n7323 0.00658571
R16001 DVDD.n7443 DVDD.n7442 0.00658571
R16002 DVDD.n7442 DVDD.n7441 0.00658571
R16003 DVDD.n7441 DVDD.n7327 0.00658571
R16004 DVDD.n7435 DVDD.n7327 0.00658571
R16005 DVDD.n7435 DVDD.n7434 0.00658571
R16006 DVDD.n7434 DVDD.n7433 0.00658571
R16007 DVDD.n7433 DVDD.n7331 0.00658571
R16008 DVDD.n7376 DVDD.n7331 0.00658571
R16009 DVDD.n7419 DVDD.n7376 0.00658571
R16010 DVDD.n7419 DVDD.n7418 0.00658571
R16011 DVDD.n7418 DVDD.n7417 0.00658571
R16012 DVDD.n7417 DVDD.n7377 0.00658571
R16013 DVDD.n7411 DVDD.n7377 0.00658571
R16014 DVDD.n7411 DVDD.n7410 0.00658571
R16015 DVDD.n7410 DVDD.n7409 0.00658571
R16016 DVDD.n7409 DVDD.n7381 0.00658571
R16017 DVDD.n7403 DVDD.n7381 0.00658571
R16018 DVDD.n7403 DVDD.n7402 0.00658571
R16019 DVDD.n7402 DVDD.n7401 0.00658571
R16020 DVDD.n7401 DVDD.n7385 0.00658571
R16021 DVDD.n7395 DVDD.n7385 0.00658571
R16022 DVDD.n7395 DVDD.n7394 0.00658571
R16023 DVDD.n7394 DVDD.n7393 0.00658571
R16024 DVDD.n7393 DVDD.n7389 0.00658571
R16025 DVDD.n7389 DVDD.n1726 0.00658571
R16026 DVDD.n8281 DVDD.n1726 0.00658571
R16027 DVDD.n8281 DVDD.n8280 0.00658571
R16028 DVDD.n8280 DVDD.n8279 0.00658571
R16029 DVDD.n8279 DVDD.n1727 0.00658571
R16030 DVDD.n8273 DVDD.n1727 0.00658571
R16031 DVDD.n8273 DVDD.n8272 0.00658571
R16032 DVDD.n8272 DVDD.n8271 0.00658571
R16033 DVDD.n8271 DVDD.n1731 0.00658571
R16034 DVDD.n8265 DVDD.n1731 0.00658571
R16035 DVDD.n8265 DVDD.n8264 0.00658571
R16036 DVDD.n8264 DVDD.n8263 0.00658571
R16037 DVDD.n8263 DVDD.n1735 0.00658571
R16038 DVDD.n8257 DVDD.n1735 0.00658571
R16039 DVDD.n8257 DVDD.n8256 0.00658571
R16040 DVDD.n8256 DVDD.n8255 0.00658571
R16041 DVDD.n8255 DVDD.n1739 0.00658571
R16042 DVDD.n1766 DVDD.n1739 0.00658571
R16043 DVDD.n8247 DVDD.n1766 0.00658571
R16044 DVDD.n8247 DVDD.n8246 0.00658571
R16045 DVDD.n8246 DVDD.n8245 0.00658571
R16046 DVDD.n8245 DVDD.n1767 0.00658571
R16047 DVDD.n8239 DVDD.n1767 0.00658571
R16048 DVDD.n8239 DVDD.n8238 0.00658571
R16049 DVDD.n8238 DVDD.n8237 0.00658571
R16050 DVDD.n8237 DVDD.n1772 0.00658571
R16051 DVDD.n8231 DVDD.n1772 0.00658571
R16052 DVDD.n8231 DVDD.n8230 0.00658571
R16053 DVDD.n8230 DVDD.n8229 0.00658571
R16054 DVDD.n8229 DVDD.n1775 0.00658571
R16055 DVDD.n8223 DVDD.n1775 0.00658571
R16056 DVDD.n8223 DVDD.n8222 0.00658571
R16057 DVDD.n8222 DVDD.n8221 0.00658571
R16058 DVDD.n8221 DVDD.n1777 0.00658571
R16059 DVDD.n8215 DVDD.n1777 0.00658571
R16060 DVDD.n8215 DVDD.n8214 0.00658571
R16061 DVDD.n8214 DVDD.n8213 0.00658571
R16062 DVDD.n8213 DVDD.n1782 0.00658571
R16063 DVDD.n8201 DVDD.n1782 0.00658571
R16064 DVDD.n6450 DVDD 0.00655123
R16065 DVDD DVDD.n3486 0.00655123
R16066 DVDD.n3887 DVDD.n3862 0.00651875
R16067 DVDD.n6432 DVDD.n1095 0.00651875
R16068 DVDD.n6002 DVDD.n5995 0.00651875
R16069 DVDD.n7786 DVDD.n2205 0.0065
R16070 DVDD.n6669 DVDD.n2116 0.0065
R16071 DVDD.n7593 DVDD.n2473 0.0065
R16072 DVDD.n7786 DVDD.n7785 0.0065
R16073 DVDD.n7268 DVDD.n2471 0.0065
R16074 DVDD.n8326 DVDD.n1584 0.0065
R16075 DVDD.n7000 DVDD.n2471 0.0065
R16076 DVDD.n2203 DVDD.n1584 0.0065
R16077 DVDD.n7856 DVDD.n2117 0.0065
R16078 DVDD.n6709 DVDD.n2203 0.0065
R16079 DVDD.n7000 DVDD.n2615 0.0065
R16080 DVDD.n6630 DVDD.n2004 0.0065
R16081 DVDD.n8035 DVDD.n2004 0.0065
R16082 DVDD.n7856 DVDD.n1927 0.0065
R16083 DVDD.n1927 DVDD.n1917 0.0065
R16084 DVDD.n8035 DVDD.n1841 0.0065
R16085 DVDD.n7593 DVDD.n2474 0.0065
R16086 DVDD.n7785 DVDD.n1587 0.0065
R16087 DVDD.n1237 DVDD.n1198 0.0065
R16088 DVDD.n2116 DVDD.n1929 0.0065
R16089 DVDD.n1929 DVDD.n1916 0.0065
R16090 DVDD.n1159 DVDD.n1120 0.0065
R16091 DVDD.n1198 DVDD.n1159 0.0065
R16092 DVDD.n6750 DVDD.n2473 0.0065
R16093 DVDD.n7503 DVDD.n7076 0.00647857
R16094 DVDD.n7298 DVDD.n7104 0.00647857
R16095 DVDD.n8365 DVDD.n1520 0.00647857
R16096 DVDD.n7431 DVDD.n7430 0.00647857
R16097 DVDD.n4711 DVDD.n4709 0.00647857
R16098 DVDD.n4738 DVDD.n4728 0.00647857
R16099 DVDD.n5115 DVDD.n4571 0.00647857
R16100 DVDD.n5028 DVDD.n4862 0.00647857
R16101 DVDD.n4551 DVDD.n4542 0.00647857
R16102 DVDD.n4788 DVDD.n4740 0.00647857
R16103 DVDD.n9243 DVDD.n457 0.00647857
R16104 DVDD.n498 DVDD.n489 0.00647857
R16105 DVDD.n6443 DVDD.n3489 0.00635
R16106 DVDD.n709 DVDD.n587 0.00634646
R16107 DVDD.n8714 DVDD.n896 0.00634646
R16108 DVDD.n3830 DVDD.n3568 0.00634646
R16109 DVDD.n2432 DVDD.n1958 0.00634646
R16110 DVDD.n8976 DVDD.n553 0.00634646
R16111 DVDD.n4069 DVDD.n3993 0.00634646
R16112 DVDD.n6038 DVDD.n3965 0.00634646
R16113 DVDD.n2439 DVDD.n2290 0.00634646
R16114 DVDD.n5018 DVDD.n4860 0.00634646
R16115 DVDD.n365 DVDD.n283 0.00634646
R16116 DVDD.n5805 DVDD.n4312 0.00634646
R16117 DVDD.n2445 DVDD.n2221 0.00634646
R16118 DVDD.n5120 DVDD.n4575 0.00634646
R16119 DVDD.n387 DVDD.n382 0.00634646
R16120 DVDD.n2865 DVDD.n2827 0.00634646
R16121 DVDD.n2449 DVDD.n2448 0.00634646
R16122 DVDD.n6098 DVDD.n5759 0.0062375
R16123 DVDD.n6099 DVDD.n4394 0.0062375
R16124 DVDD.n8287 DVDD.n1705 0.00622143
R16125 DVDD.n1724 DVDD.n1704 0.00622143
R16126 DVDD.n8253 DVDD.n8252 0.00622143
R16127 DVDD.n8250 DVDD.n8249 0.00622143
R16128 DVDD.n8648 DVDD.n1274 0.00622143
R16129 DVDD.n8224 DVDD.n1273 0.00622143
R16130 DVDD.n1784 DVDD.n1780 0.00622143
R16131 DVDD.n8208 DVDD.n1797 0.00622143
R16132 DVDD.n9013 DVDD.n552 0.00622143
R16133 DVDD.n8965 DVDD.n551 0.00622143
R16134 DVDD.n8939 DVDD.n8938 0.00622143
R16135 DVDD.n592 DVDD.n589 0.00622143
R16136 DVDD.n8919 DVDD.n606 0.00622143
R16137 DVDD.n8912 DVDD.n617 0.00622143
R16138 DVDD.n8901 DVDD.n637 0.00622143
R16139 DVDD.n8894 DVDD.n648 0.00622143
R16140 DVDD.n9176 DVDD.n9175 0.00622143
R16141 DVDD.n9173 DVDD.n9172 0.00622143
R16142 DVDD.n9143 DVDD.n73 0.00622143
R16143 DVDD.n9647 DVDD.n65 0.00622143
R16144 DVDD.n9672 DVDD.n9670 0.00622143
R16145 DVDD.n9674 DVDD.n30 0.00622143
R16146 DVDD.n8937 DVDD.n588 0.00599213
R16147 DVDD.n9622 DVDD.n91 0.00599213
R16148 DVDD.n3822 DVDD.n3570 0.00599213
R16149 DVDD.n3415 DVDD.n3339 0.00599213
R16150 DVDD.n9004 DVDD.n8972 0.00599213
R16151 DVDD.n4012 DVDD.n4011 0.00599213
R16152 DVDD.n6046 DVDD.n3967 0.00599213
R16153 DVDD.n5943 DVDD.n3216 0.00599213
R16154 DVDD.n5010 DVDD.n4858 0.00599213
R16155 DVDD.n9465 DVDD.n295 0.00599213
R16156 DVDD.n5813 DVDD.n4314 0.00599213
R16157 DVDD.n5841 DVDD.n3104 0.00599213
R16158 DVDD.n5148 DVDD.n5116 0.00599213
R16159 DVDD.n9311 DVDD.n444 0.00599213
R16160 DVDD.n2875 DVDD.n2874 0.00599213
R16161 DVDD.n6903 DVDD.n2733 0.00599213
R16162 DVDD.n6448 DVDD.n3487 0.00597492
R16163 DVDD.n7496 DVDD.n7068 0.00596429
R16164 DVDD.n7310 DVDD.n7304 0.00596429
R16165 DVDD.n7320 DVDD.n1512 0.00596429
R16166 DVDD.n7425 DVDD.n7421 0.00596429
R16167 DVDD.n4713 DVDD.n4609 0.00596429
R16168 DVDD.n4821 DVDD.n4589 0.00596429
R16169 DVDD.n5107 DVDD.n4570 0.00596429
R16170 DVDD.n5080 DVDD.n5079 0.00596429
R16171 DVDD.n4764 DVDD.n4543 0.00596429
R16172 DVDD.n4816 DVDD.n4815 0.00596429
R16173 DVDD.n9235 DVDD.n456 0.00596429
R16174 DVDD.n9208 DVDD.n9207 0.00596429
R16175 DVDD.n355 DVDD 0.00587887
R16176 DVDD.n354 DVDD 0.00587887
R16177 DVDD.n9691 DVDD.n3 0.00583571
R16178 DVDD.n6233 DVDD.n3883 0.005825
R16179 DVDD.n6228 DVDD.n3883 0.005825
R16180 DVDD.n6228 DVDD.n6227 0.005825
R16181 DVDD.n6227 DVDD.n6226 0.005825
R16182 DVDD.n6226 DVDD.n3888 0.005825
R16183 DVDD.n6220 DVDD.n3888 0.005825
R16184 DVDD.n6220 DVDD.n6219 0.005825
R16185 DVDD.n6219 DVDD.n6218 0.005825
R16186 DVDD.n6218 DVDD.n6212 0.005825
R16187 DVDD.n6212 DVDD.n6211 0.005825
R16188 DVDD.n6428 DVDD.n3508 0.005825
R16189 DVDD.n6429 DVDD.n6428 0.005825
R16190 DVDD.n6430 DVDD.n6429 0.005825
R16191 DVDD.n6430 DVDD.n3504 0.005825
R16192 DVDD.n6437 DVDD.n3504 0.005825
R16193 DVDD.n6438 DVDD.n6437 0.005825
R16194 DVDD.n6439 DVDD.n6438 0.005825
R16195 DVDD.n6439 DVDD.n3502 0.005825
R16196 DVDD.n6444 DVDD.n3502 0.005825
R16197 DVDD.n6081 DVDD.n5909 0.005825
R16198 DVDD.n6075 DVDD.n5909 0.005825
R16199 DVDD.n6075 DVDD.n6074 0.005825
R16200 DVDD.n6074 DVDD.n6073 0.005825
R16201 DVDD.n6073 DVDD.n5915 0.005825
R16202 DVDD.n6067 DVDD.n5915 0.005825
R16203 DVDD.n6067 DVDD.n6066 0.005825
R16204 DVDD.n6066 DVDD.n6065 0.005825
R16205 DVDD.n6065 DVDD.n5919 0.005825
R16206 DVDD.n5919 DVDD.n3914 0.005825
R16207 DVDD.n3943 DVDD.n3915 0.005825
R16208 DVDD.n3937 DVDD.n3915 0.005825
R16209 DVDD.n3937 DVDD.n3936 0.005825
R16210 DVDD.n3936 DVDD.n3935 0.005825
R16211 DVDD.n3935 DVDD.n3919 0.005825
R16212 DVDD.n3929 DVDD.n3919 0.005825
R16213 DVDD.n3929 DVDD.n3928 0.005825
R16214 DVDD.n3928 DVDD.n3927 0.005825
R16215 DVDD.n3927 DVDD.n3882 0.005825
R16216 DVDD.n4406 DVDD.n2787 0.005825
R16217 DVDD.n4406 DVDD.n4402 0.005825
R16218 DVDD.n4412 DVDD.n4402 0.005825
R16219 DVDD.n4413 DVDD.n4412 0.005825
R16220 DVDD.n4414 DVDD.n4413 0.005825
R16221 DVDD.n4414 DVDD.n4398 0.005825
R16222 DVDD.n4421 DVDD.n4398 0.005825
R16223 DVDD.n4422 DVDD.n4421 0.005825
R16224 DVDD.n4423 DVDD.n4422 0.005825
R16225 DVDD.n4423 DVDD.n4392 0.005825
R16226 DVDD.n6100 DVDD.n4393 0.005825
R16227 DVDD.n5901 DVDD.n4393 0.005825
R16228 DVDD.n5902 DVDD.n5901 0.005825
R16229 DVDD.n6092 DVDD.n5902 0.005825
R16230 DVDD.n6092 DVDD.n6091 0.005825
R16231 DVDD.n6091 DVDD.n6090 0.005825
R16232 DVDD.n6090 DVDD.n5903 0.005825
R16233 DVDD.n6084 DVDD.n5903 0.005825
R16234 DVDD.n6084 DVDD.n6083 0.005825
R16235 DVDD.n5648 DVDD.n4457 0.005825
R16236 DVDD.n5662 DVDD.n4457 0.005825
R16237 DVDD.n5663 DVDD.n5662 0.005825
R16238 DVDD.n5665 DVDD.n5663 0.005825
R16239 DVDD.n5665 DVDD.n5664 0.005825
R16240 DVDD.n5664 DVDD.n4454 0.005825
R16241 DVDD.n4454 DVDD.n4452 0.005825
R16242 DVDD.n5673 DVDD.n4452 0.005825
R16243 DVDD.n5674 DVDD.n5673 0.005825
R16244 DVDD.n5675 DVDD.n5674 0.005825
R16245 DVDD.n5684 DVDD.n5681 0.005825
R16246 DVDD.n5703 DVDD.n5684 0.005825
R16247 DVDD.n5703 DVDD.n5702 0.005825
R16248 DVDD.n5702 DVDD.n5701 0.005825
R16249 DVDD.n5701 DVDD.n5685 0.005825
R16250 DVDD.n5695 DVDD.n5685 0.005825
R16251 DVDD.n5695 DVDD.n5694 0.005825
R16252 DVDD.n5694 DVDD.n5693 0.005825
R16253 DVDD.n5693 DVDD.n2788 0.005825
R16254 DVDD.n5709 DVDD.n5708 0.0057875
R16255 DVDD.n5891 DVDD.n5765 0.00573125
R16256 DVDD.n5650 DVDD.n5483 0.00573125
R16257 DVDD.n3022 DVDD.n3008 0.00573125
R16258 DVDD.n5689 DVDD.n2777 0.00573125
R16259 DVDD.n8766 DVDD.n848 0.0056378
R16260 DVDD.n6260 DVDD.n3347 0.0056378
R16261 DVDD.n2409 DVDD.n1953 0.0056378
R16262 DVDD.n4096 DVDD.n4016 0.0056378
R16263 DVDD.n5951 DVDD.n3231 0.0056378
R16264 DVDD.n2416 DVDD.n2289 0.0056378
R16265 DVDD.n9458 DVDD.n307 0.0056378
R16266 DVDD.n5849 DVDD.n3112 0.0056378
R16267 DVDD.n2422 DVDD.n2216 0.0056378
R16268 DVDD.n9612 DVDD.n9611 0.0056378
R16269 DVDD.n6911 DVDD.n2663 0.0056378
R16270 DVDD.n2426 DVDD.n2425 0.0056378
R16271 DVDD.n8205 DVDD 0.00557857
R16272 DVDD.n8892 DVDD 0.00557857
R16273 DVDD.n6230 DVDD.n3864 0.00550625
R16274 DVDD.n3506 DVDD.n1096 0.00550625
R16275 DVDD.n6464 DVDD.n3468 0.00550625
R16276 DVDD.n6069 DVDD.n5917 0.00550625
R16277 DVDD.n6062 DVDD.n5928 0.00550625
R16278 DVDD.n8790 DVDD.n8789 0.00545
R16279 DVDD.n8779 DVDD.n86 0.00545
R16280 DVDD.n8778 DVDD.n8777 0.00545
R16281 DVDD.n8774 DVDD.n90 0.00545
R16282 DVDD.n8773 DVDD.n840 0.00545
R16283 DVDD.n924 DVDD.n115 0.00545
R16284 DVDD.n926 DVDD.n851 0.00545
R16285 DVDD.n929 DVDD.n854 0.00545
R16286 DVDD.n944 DVDD.n943 0.00545
R16287 DVDD.n946 DVDD.n868 0.00545
R16288 DVDD.n949 DVDD.n923 0.00545
R16289 DVDD DVDD.n8201 0.00538571
R16290 DVDD.n7502 DVDD.n7069 0.00532143
R16291 DVDD.n7485 DVDD.n7299 0.00532143
R16292 DVDD.n1527 DVDD.n1513 0.00532143
R16293 DVDD.n7428 DVDD.n7339 0.00532143
R16294 DVDD.n4710 DVDD.n4613 0.00532143
R16295 DVDD.n4737 DVDD.n4593 0.00532143
R16296 DVDD.n4581 DVDD.n4573 0.00532143
R16297 DVDD.n5033 DVDD.n4869 0.00532143
R16298 DVDD.n4757 DVDD.n4544 0.00532143
R16299 DVDD.n4790 DVDD.n4741 0.00532143
R16300 DVDD.n466 DVDD.n459 0.00532143
R16301 DVDD.n503 DVDD.n496 0.00532143
R16302 DVDD.n9579 DVDD.n193 0.00530256
R16303 DVDD.n6882 DVDD.n2788 0.0053
R16304 DVDD.n717 DVDD.n580 0.00528346
R16305 DVDD.n9646 DVDD.n71 0.00528346
R16306 DVDD.n8734 DVDD.n880 0.00528346
R16307 DVDD.n8671 DVDD.n1049 0.00528346
R16308 DVDD.n3838 DVDD.n3813 0.00528346
R16309 DVDD.n6518 DVDD.n2083 0.00528346
R16310 DVDD.n8981 DVDD.n8974 0.00528346
R16311 DVDD.n9121 DVDD.n527 0.00528346
R16312 DVDD.n4078 DVDD.n4028 0.00528346
R16313 DVDD.n4206 DVDD.n4154 0.00528346
R16314 DVDD.n6030 DVDD.n3953 0.00528346
R16315 DVDD.n3281 DVDD.n2143 0.00528346
R16316 DVDD.n5027 DVDD.n4863 0.00528346
R16317 DVDD.n9209 DVDD.n495 0.00528346
R16318 DVDD.n9433 DVDD.n9432 0.00528346
R16319 DVDD.n9550 DVDD.n9549 0.00528346
R16320 DVDD.n5797 DVDD.n4382 0.00528346
R16321 DVDD.n3172 DVDD.n2180 0.00528346
R16322 DVDD.n5125 DVDD.n5118 0.00528346
R16323 DVDD.n9278 DVDD.n9244 0.00528346
R16324 DVDD.n9392 DVDD.n173 0.00528346
R16325 DVDD.n6782 DVDD.n6781 0.00528346
R16326 DVDD.n2857 DVDD.n2814 0.00528346
R16327 DVDD.n2702 DVDD.n2633 0.00528346
R16328 DVDD.n6095 DVDD.n6094 0.00528125
R16329 DVDD.n5659 DVDD.n4455 0.00528125
R16330 DVDD.n5707 DVDD.n3000 0.00528125
R16331 DVDD.n1048 DVDD.n1047 0.005225
R16332 DVDD.n8726 DVDD.n8725 0.005225
R16333 DVDD.n6320 DVDD.n6319 0.005225
R16334 DVDD.n6871 DVDD.n2793 0.005225
R16335 DVDD.n174 DVDD.n164 0.005225
R16336 DVDD.n2913 DVDD.n2912 0.005225
R16337 DVDD.n9605 DVDD.n138 0.005225
R16338 DVDD.n8759 DVDD.n857 0.005225
R16339 DVDD.n6451 DVDD.n6450 0.00520651
R16340 DVDD.n7719 DVDD.n1861 0.0051063
R16341 DVDD.n7724 DVDD.n1664 0.0051063
R16342 DVDD.n7701 DVDD.n1595 0.0051063
R16343 DVDD.n7694 DVDD.n1540 0.0051063
R16344 DVDD.n8284 DVDD.n1712 0.00506429
R16345 DVDD.n8284 DVDD.n8283 0.00506429
R16346 DVDD.n1757 DVDD.n1746 0.00506429
R16347 DVDD.n1758 DVDD.n1757 0.00506429
R16348 DVDD.n1294 DVDD.n1280 0.00506429
R16349 DVDD.n8226 DVDD.n1294 0.00506429
R16350 DVDD.n8211 DVDD.n8210 0.00506429
R16351 DVDD.n8210 DVDD.n1790 0.00506429
R16352 DVDD.n8971 DVDD.n549 0.00506429
R16353 DVDD.n559 DVDD.n549 0.00506429
R16354 DVDD.n591 DVDD.n582 0.00506429
R16355 DVDD.n596 DVDD.n591 0.00506429
R16356 DVDD.n611 DVDD.n610 0.00506429
R16357 DVDD.n8913 DVDD.n611 0.00506429
R16358 DVDD.n642 DVDD.n641 0.00506429
R16359 DVDD.n8895 DVDD.n642 0.00506429
R16360 DVDD.n534 DVDD.n526 0.00506429
R16361 DVDD.n9126 DVDD.n534 0.00506429
R16362 DVDD.n72 DVDD.n59 0.00506429
R16363 DVDD.n9648 DVDD.n59 0.00506429
R16364 DVDD.n9671 DVDD.n24 0.00506429
R16365 DVDD.n9675 DVDD.n24 0.00506429
R16366 DVDD.n6083 DVDD.n6082 0.005
R16367 DVDD.n8820 DVDD.n66 0.00492913
R16368 DVDD.n6333 DVDD.n3818 0.00492913
R16369 DVDD.n6528 DVDD.n3332 0.00492913
R16370 DVDD.n6496 DVDD.n2088 0.00492913
R16371 DVDD.n9092 DVDD.n523 0.00492913
R16372 DVDD.n6008 DVDD.n3958 0.00492913
R16373 DVDD.n3292 DVDD.n3228 0.00492913
R16374 DVDD.n3259 DVDD.n2138 0.00492913
R16375 DVDD.n4935 DVDD.n490 0.00492913
R16376 DVDD.n6112 DVDD.n4387 0.00492913
R16377 DVDD.n3125 DVDD.n3097 0.00492913
R16378 DVDD.n3150 DVDD.n2185 0.00492913
R16379 DVDD.n9285 DVDD.n458 0.00492913
R16380 DVDD.n2835 DVDD.n2819 0.00492913
R16381 DVDD.n2713 DVDD.n2673 0.00492913
R16382 DVDD.n2680 DVDD.n2643 0.00492913
R16383 DVDD.n6210 DVDD.n3508 0.004925
R16384 DVDD.n7091 DVDD.n7069 0.00480714
R16385 DVDD.n7485 DVDD.n7484 0.00480714
R16386 DVDD.n7460 DVDD.n1513 0.00480714
R16387 DVDD.n7428 DVDD.n7369 0.00480714
R16388 DVDD.n4714 DVDD.n4613 0.00480714
R16389 DVDD.n4822 DVDD.n4593 0.00480714
R16390 DVDD.n5109 DVDD.n4573 0.00480714
R16391 DVDD.n5029 DVDD.n4869 0.00480714
R16392 DVDD.n4759 DVDD.n4544 0.00480714
R16393 DVDD.n4742 DVDD.n4741 0.00480714
R16394 DVDD.n9237 DVDD.n459 0.00480714
R16395 DVDD.n499 DVDD.n496 0.00480714
R16396 DVDD.n6446 DVDD.n6445 0.00479029
R16397 DVDD.n5529 DVDD.n5528 0.00476
R16398 DVDD.n5528 DVDD.n5526 0.00476
R16399 DVDD.n5526 DVDD.n5524 0.00476
R16400 DVDD.n5524 DVDD.n5511 0.00476
R16401 DVDD.n5520 DVDD.n5511 0.00476
R16402 DVDD.n5520 DVDD.n5519 0.00476
R16403 DVDD.n5519 DVDD.n5518 0.00476
R16404 DVDD.n5518 DVDD.n3061 0.00476
R16405 DVDD.n6753 DVDD.n3061 0.00476
R16406 DVDD.n6753 DVDD.n6752 0.00476
R16407 DVDD.n6746 DVDD.n3064 0.00476
R16408 DVDD.n6742 DVDD.n3064 0.00476
R16409 DVDD.n6742 DVDD.n6741 0.00476
R16410 DVDD.n6741 DVDD.n6740 0.00476
R16411 DVDD.n6740 DVDD.n3069 0.00476
R16412 DVDD.n6736 DVDD.n3069 0.00476
R16413 DVDD.n6736 DVDD.n6735 0.00476
R16414 DVDD.n6735 DVDD.n6734 0.00476
R16415 DVDD.n6734 DVDD.n6732 0.00476
R16416 DVDD.n6732 DVDD.n6730 0.00476
R16417 DVDD.n6730 DVDD.n6728 0.00476
R16418 DVDD.n6728 DVDD.n6727 0.00476
R16419 DVDD.n6727 DVDD.n6726 0.00476
R16420 DVDD.n6726 DVDD.n3080 0.00476
R16421 DVDD.n6722 DVDD.n3080 0.00476
R16422 DVDD.n6722 DVDD.n6721 0.00476
R16423 DVDD.n6721 DVDD.n6720 0.00476
R16424 DVDD.n6720 DVDD.n3086 0.00476
R16425 DVDD.n6716 DVDD.n3086 0.00476
R16426 DVDD.n6716 DVDD.n6715 0.00476
R16427 DVDD.n6715 DVDD.n6714 0.00476
R16428 DVDD.n6714 DVDD.n3092 0.00476
R16429 DVDD.n6710 DVDD.n3092 0.00476
R16430 DVDD.n6708 DVDD.n3096 0.00476
R16431 DVDD.n3190 DVDD.n3096 0.00476
R16432 DVDD.n3190 DVDD.n3187 0.00476
R16433 DVDD.n6699 DVDD.n3187 0.00476
R16434 DVDD.n6699 DVDD.n6698 0.00476
R16435 DVDD.n6698 DVDD.n6697 0.00476
R16436 DVDD.n6697 DVDD.n3196 0.00476
R16437 DVDD.n6693 DVDD.n3196 0.00476
R16438 DVDD.n6693 DVDD.n6692 0.00476
R16439 DVDD.n6692 DVDD.n6691 0.00476
R16440 DVDD.n6691 DVDD.n3202 0.00476
R16441 DVDD.n6687 DVDD.n3202 0.00476
R16442 DVDD.n6687 DVDD.n6686 0.00476
R16443 DVDD.n6686 DVDD.n6685 0.00476
R16444 DVDD.n6685 DVDD.n3208 0.00476
R16445 DVDD.n6681 DVDD.n3208 0.00476
R16446 DVDD.n6681 DVDD.n6680 0.00476
R16447 DVDD.n6680 DVDD.n6679 0.00476
R16448 DVDD.n6679 DVDD.n3214 0.00476
R16449 DVDD.n3309 DVDD.n3214 0.00476
R16450 DVDD.n3309 DVDD.n3307 0.00476
R16451 DVDD.n6672 DVDD.n3307 0.00476
R16452 DVDD.n6672 DVDD.n6671 0.00476
R16453 DVDD.n6667 DVDD.n6666 0.00476
R16454 DVDD.n6666 DVDD.n6665 0.00476
R16455 DVDD.n6665 DVDD.n3319 0.00476
R16456 DVDD.n6661 DVDD.n3319 0.00476
R16457 DVDD.n6661 DVDD.n6660 0.00476
R16458 DVDD.n6660 DVDD.n6659 0.00476
R16459 DVDD.n6659 DVDD.n3325 0.00476
R16460 DVDD.n6655 DVDD.n3325 0.00476
R16461 DVDD.n6655 DVDD.n6654 0.00476
R16462 DVDD.n6654 DVDD.n6653 0.00476
R16463 DVDD.n6653 DVDD.n3331 0.00476
R16464 DVDD.n3368 DVDD.n3331 0.00476
R16465 DVDD.n3370 DVDD.n3368 0.00476
R16466 DVDD.n3370 DVDD.n3365 0.00476
R16467 DVDD.n6643 DVDD.n3365 0.00476
R16468 DVDD.n6643 DVDD.n6642 0.00476
R16469 DVDD.n6642 DVDD.n6641 0.00476
R16470 DVDD.n6641 DVDD.n3376 0.00476
R16471 DVDD.n6637 DVDD.n3376 0.00476
R16472 DVDD.n6637 DVDD.n6636 0.00476
R16473 DVDD.n6636 DVDD.n6635 0.00476
R16474 DVDD.n6635 DVDD.n3382 0.00476
R16475 DVDD.n6631 DVDD.n3382 0.00476
R16476 DVDD.n6629 DVDD.n6628 0.00476
R16477 DVDD.n6628 DVDD.n6615 0.00476
R16478 DVDD.n6615 DVDD.n6613 0.00476
R16479 DVDD.n6613 DVDD.n3389 0.00476
R16480 DVDD.n6609 DVDD.n3389 0.00476
R16481 DVDD.n6609 DVDD.n6608 0.00476
R16482 DVDD.n6608 DVDD.n6607 0.00476
R16483 DVDD.n6607 DVDD.n3395 0.00476
R16484 DVDD.n6594 DVDD.n3395 0.00476
R16485 DVDD.n6601 DVDD.n6594 0.00476
R16486 DVDD.n7016 DVDD.n2550 0.00476
R16487 DVDD.n7016 DVDD.n7015 0.00476
R16488 DVDD.n7015 DVDD.n7013 0.00476
R16489 DVDD.n7013 DVDD.n2554 0.00476
R16490 DVDD.n7009 DVDD.n2554 0.00476
R16491 DVDD.n7009 DVDD.n7008 0.00476
R16492 DVDD.n7008 DVDD.n7007 0.00476
R16493 DVDD.n7007 DVDD.n2560 0.00476
R16494 DVDD.n2611 DVDD.n2560 0.00476
R16495 DVDD.n7001 DVDD.n2611 0.00476
R16496 DVDD.n6999 DVDD.n2617 0.00476
R16497 DVDD.n6995 DVDD.n2617 0.00476
R16498 DVDD.n6995 DVDD.n6994 0.00476
R16499 DVDD.n6994 DVDD.n6993 0.00476
R16500 DVDD.n6993 DVDD.n2623 0.00476
R16501 DVDD.n6989 DVDD.n2623 0.00476
R16502 DVDD.n6989 DVDD.n6988 0.00476
R16503 DVDD.n6988 DVDD.n6987 0.00476
R16504 DVDD.n6987 DVDD.n2629 0.00476
R16505 DVDD.n6975 DVDD.n2629 0.00476
R16506 DVDD.n6975 DVDD.n6974 0.00476
R16507 DVDD.n6974 DVDD.n6973 0.00476
R16508 DVDD.n6973 DVDD.n6972 0.00476
R16509 DVDD.n6972 DVDD.n6947 0.00476
R16510 DVDD.n6968 DVDD.n6947 0.00476
R16511 DVDD.n6968 DVDD.n6967 0.00476
R16512 DVDD.n6967 DVDD.n6966 0.00476
R16513 DVDD.n6966 DVDD.n6953 0.00476
R16514 DVDD.n6962 DVDD.n6953 0.00476
R16515 DVDD.n6962 DVDD.n6961 0.00476
R16516 DVDD.n6961 DVDD.n6960 0.00476
R16517 DVDD.n6960 DVDD.n2202 0.00476
R16518 DVDD.n7788 DVDD.n2202 0.00476
R16519 DVDD.n7793 DVDD.n2197 0.00476
R16520 DVDD.n7793 DVDD.n2170 0.00476
R16521 DVDD.n7808 DVDD.n2170 0.00476
R16522 DVDD.n7808 DVDD.n2168 0.00476
R16523 DVDD.n7812 DVDD.n2168 0.00476
R16524 DVDD.n7812 DVDD.n2166 0.00476
R16525 DVDD.n7816 DVDD.n2166 0.00476
R16526 DVDD.n7816 DVDD.n2164 0.00476
R16527 DVDD.n7820 DVDD.n2164 0.00476
R16528 DVDD.n7820 DVDD.n2162 0.00476
R16529 DVDD.n7824 DVDD.n2162 0.00476
R16530 DVDD.n7824 DVDD.n2160 0.00476
R16531 DVDD.n7828 DVDD.n2160 0.00476
R16532 DVDD.n7828 DVDD.n2158 0.00476
R16533 DVDD.n7832 DVDD.n2158 0.00476
R16534 DVDD.n7832 DVDD.n2156 0.00476
R16535 DVDD.n7836 DVDD.n2156 0.00476
R16536 DVDD.n7836 DVDD.n2154 0.00476
R16537 DVDD.n7844 DVDD.n2154 0.00476
R16538 DVDD.n7844 DVDD.n2152 0.00476
R16539 DVDD.n7849 DVDD.n2152 0.00476
R16540 DVDD.n7849 DVDD.n2118 0.00476
R16541 DVDD.n7855 DVDD.n2118 0.00476
R16542 DVDD.n7858 DVDD.n2115 0.00476
R16543 DVDD.n7862 DVDD.n2115 0.00476
R16544 DVDD.n7862 DVDD.n2113 0.00476
R16545 DVDD.n7866 DVDD.n2113 0.00476
R16546 DVDD.n7866 DVDD.n2111 0.00476
R16547 DVDD.n7870 DVDD.n2111 0.00476
R16548 DVDD.n7870 DVDD.n2109 0.00476
R16549 DVDD.n7875 DVDD.n2109 0.00476
R16550 DVDD.n7875 DVDD.n2107 0.00476
R16551 DVDD.n7879 DVDD.n2107 0.00476
R16552 DVDD.n7880 DVDD.n7879 0.00476
R16553 DVDD.n7880 DVDD.n2105 0.00476
R16554 DVDD.n7884 DVDD.n2105 0.00476
R16555 DVDD.n7884 DVDD.n2073 0.00476
R16556 DVDD.n7895 DVDD.n2073 0.00476
R16557 DVDD.n7895 DVDD.n2071 0.00476
R16558 DVDD.n7899 DVDD.n2071 0.00476
R16559 DVDD.n7899 DVDD.n2069 0.00476
R16560 DVDD.n7903 DVDD.n2069 0.00476
R16561 DVDD.n7903 DVDD.n2067 0.00476
R16562 DVDD.n7907 DVDD.n2067 0.00476
R16563 DVDD.n7907 DVDD.n2065 0.00476
R16564 DVDD.n7911 DVDD.n2065 0.00476
R16565 DVDD.n7928 DVDD.n7915 0.00476
R16566 DVDD.n7930 DVDD.n7928 0.00476
R16567 DVDD.n7930 DVDD.n2061 0.00476
R16568 DVDD.n7935 DVDD.n2061 0.00476
R16569 DVDD.n7935 DVDD.n2059 0.00476
R16570 DVDD.n7939 DVDD.n2059 0.00476
R16571 DVDD.n7940 DVDD.n7939 0.00476
R16572 DVDD.n7940 DVDD.n2057 0.00476
R16573 DVDD.n7950 DVDD.n2057 0.00476
R16574 DVDD.n7950 DVDD.n7949 0.00476
R16575 DVDD.n7522 DVDD.n2507 0.00476
R16576 DVDD.n7552 DVDD.n2507 0.00476
R16577 DVDD.n7552 DVDD.n2505 0.00476
R16578 DVDD.n7556 DVDD.n2505 0.00476
R16579 DVDD.n7556 DVDD.n2503 0.00476
R16580 DVDD.n7560 DVDD.n2503 0.00476
R16581 DVDD.n7560 DVDD.n2501 0.00476
R16582 DVDD.n7564 DVDD.n2501 0.00476
R16583 DVDD.n7564 DVDD.n2470 0.00476
R16584 DVDD.n7595 DVDD.n2470 0.00476
R16585 DVDD.n7600 DVDD.n2466 0.00476
R16586 DVDD.n7600 DVDD.n2464 0.00476
R16587 DVDD.n7604 DVDD.n2464 0.00476
R16588 DVDD.n7604 DVDD.n2462 0.00476
R16589 DVDD.n7608 DVDD.n2462 0.00476
R16590 DVDD.n7608 DVDD.n2460 0.00476
R16591 DVDD.n7612 DVDD.n2460 0.00476
R16592 DVDD.n7612 DVDD.n2458 0.00476
R16593 DVDD.n7655 DVDD.n2458 0.00476
R16594 DVDD.n7655 DVDD.n7654 0.00476
R16595 DVDD.n7654 DVDD.n7652 0.00476
R16596 DVDD.n7652 DVDD.n7651 0.00476
R16597 DVDD.n7651 DVDD.n7650 0.00476
R16598 DVDD.n7650 DVDD.n7620 0.00476
R16599 DVDD.n7646 DVDD.n7620 0.00476
R16600 DVDD.n7646 DVDD.n7645 0.00476
R16601 DVDD.n7645 DVDD.n7644 0.00476
R16602 DVDD.n7644 DVDD.n7626 0.00476
R16603 DVDD.n7640 DVDD.n7626 0.00476
R16604 DVDD.n7640 DVDD.n7639 0.00476
R16605 DVDD.n7639 DVDD.n7638 0.00476
R16606 DVDD.n7638 DVDD.n7635 0.00476
R16607 DVDD.n7635 DVDD.n7634 0.00476
R16608 DVDD.n7783 DVDD.n7782 0.00476
R16609 DVDD.n7782 DVDD.n2210 0.00476
R16610 DVDD.n2252 DVDD.n2210 0.00476
R16611 DVDD.n7772 DVDD.n2252 0.00476
R16612 DVDD.n7772 DVDD.n7771 0.00476
R16613 DVDD.n7771 DVDD.n7770 0.00476
R16614 DVDD.n7770 DVDD.n2258 0.00476
R16615 DVDD.n7766 DVDD.n2258 0.00476
R16616 DVDD.n7766 DVDD.n7765 0.00476
R16617 DVDD.n7765 DVDD.n7764 0.00476
R16618 DVDD.n7764 DVDD.n2264 0.00476
R16619 DVDD.n7760 DVDD.n2264 0.00476
R16620 DVDD.n7760 DVDD.n7759 0.00476
R16621 DVDD.n7759 DVDD.n7758 0.00476
R16622 DVDD.n7758 DVDD.n2270 0.00476
R16623 DVDD.n7754 DVDD.n2270 0.00476
R16624 DVDD.n7754 DVDD.n7753 0.00476
R16625 DVDD.n7753 DVDD.n7752 0.00476
R16626 DVDD.n7752 DVDD.n2276 0.00476
R16627 DVDD.n2310 DVDD.n2276 0.00476
R16628 DVDD.n2310 DVDD.n2308 0.00476
R16629 DVDD.n2314 DVDD.n2308 0.00476
R16630 DVDD.n2315 DVDD.n2314 0.00476
R16631 DVDD.n8076 DVDD.n1928 0.00476
R16632 DVDD.n8072 DVDD.n1928 0.00476
R16633 DVDD.n8072 DVDD.n8071 0.00476
R16634 DVDD.n8071 DVDD.n8070 0.00476
R16635 DVDD.n8070 DVDD.n1934 0.00476
R16636 DVDD.n8066 DVDD.n1934 0.00476
R16637 DVDD.n8066 DVDD.n8065 0.00476
R16638 DVDD.n8065 DVDD.n8064 0.00476
R16639 DVDD.n8064 DVDD.n1940 0.00476
R16640 DVDD.n8060 DVDD.n1940 0.00476
R16641 DVDD.n8060 DVDD.n8059 0.00476
R16642 DVDD.n8059 DVDD.n8058 0.00476
R16643 DVDD.n8058 DVDD.n1946 0.00476
R16644 DVDD.n1989 DVDD.n1946 0.00476
R16645 DVDD.n8048 DVDD.n1989 0.00476
R16646 DVDD.n8048 DVDD.n8047 0.00476
R16647 DVDD.n8047 DVDD.n8046 0.00476
R16648 DVDD.n8046 DVDD.n1995 0.00476
R16649 DVDD.n8042 DVDD.n1995 0.00476
R16650 DVDD.n8042 DVDD.n8041 0.00476
R16651 DVDD.n8041 DVDD.n8040 0.00476
R16652 DVDD.n8040 DVDD.n2001 0.00476
R16653 DVDD.n8036 DVDD.n2001 0.00476
R16654 DVDD.n8034 DVDD.n8033 0.00476
R16655 DVDD.n8033 DVDD.n8020 0.00476
R16656 DVDD.n8020 DVDD.n8018 0.00476
R16657 DVDD.n8018 DVDD.n2009 0.00476
R16658 DVDD.n8014 DVDD.n2009 0.00476
R16659 DVDD.n8014 DVDD.n8013 0.00476
R16660 DVDD.n8013 DVDD.n8012 0.00476
R16661 DVDD.n8012 DVDD.n2015 0.00476
R16662 DVDD.n7999 DVDD.n2015 0.00476
R16663 DVDD.n8006 DVDD.n7999 0.00476
R16664 DVDD.n7224 DVDD.n7211 0.00476
R16665 DVDD.n7226 DVDD.n7224 0.00476
R16666 DVDD.n7226 DVDD.n7209 0.00476
R16667 DVDD.n7231 DVDD.n7209 0.00476
R16668 DVDD.n7231 DVDD.n7207 0.00476
R16669 DVDD.n7235 DVDD.n7207 0.00476
R16670 DVDD.n7236 DVDD.n7235 0.00476
R16671 DVDD.n7236 DVDD.n7205 0.00476
R16672 DVDD.n7271 DVDD.n7205 0.00476
R16673 DVDD.n7271 DVDD.n7270 0.00476
R16674 DVDD.n7267 DVDD.n7242 0.00476
R16675 DVDD.n7263 DVDD.n7242 0.00476
R16676 DVDD.n7263 DVDD.n7262 0.00476
R16677 DVDD.n7262 DVDD.n7261 0.00476
R16678 DVDD.n7261 DVDD.n7248 0.00476
R16679 DVDD.n7257 DVDD.n7248 0.00476
R16680 DVDD.n7257 DVDD.n7256 0.00476
R16681 DVDD.n7256 DVDD.n7255 0.00476
R16682 DVDD.n7255 DVDD.n1563 0.00476
R16683 DVDD.n8347 DVDD.n1563 0.00476
R16684 DVDD.n8347 DVDD.n8346 0.00476
R16685 DVDD.n8346 DVDD.n8344 0.00476
R16686 DVDD.n8344 DVDD.n1567 0.00476
R16687 DVDD.n8340 DVDD.n1567 0.00476
R16688 DVDD.n8340 DVDD.n8339 0.00476
R16689 DVDD.n8339 DVDD.n8338 0.00476
R16690 DVDD.n8338 DVDD.n1573 0.00476
R16691 DVDD.n8334 DVDD.n1573 0.00476
R16692 DVDD.n8334 DVDD.n8333 0.00476
R16693 DVDD.n8333 DVDD.n8332 0.00476
R16694 DVDD.n8332 DVDD.n1579 0.00476
R16695 DVDD.n8328 DVDD.n1579 0.00476
R16696 DVDD.n8328 DVDD.n8327 0.00476
R16697 DVDD.n8325 DVDD.n1586 0.00476
R16698 DVDD.n1630 DVDD.n1586 0.00476
R16699 DVDD.n8319 DVDD.n1630 0.00476
R16700 DVDD.n8319 DVDD.n8318 0.00476
R16701 DVDD.n8318 DVDD.n1635 0.00476
R16702 DVDD.n8314 DVDD.n1635 0.00476
R16703 DVDD.n8314 DVDD.n8313 0.00476
R16704 DVDD.n8313 DVDD.n8312 0.00476
R16705 DVDD.n8312 DVDD.n1641 0.00476
R16706 DVDD.n8308 DVDD.n1641 0.00476
R16707 DVDD.n8308 DVDD.n8307 0.00476
R16708 DVDD.n8307 DVDD.n8306 0.00476
R16709 DVDD.n8306 DVDD.n1647 0.00476
R16710 DVDD.n8302 DVDD.n1647 0.00476
R16711 DVDD.n8302 DVDD.n8301 0.00476
R16712 DVDD.n8301 DVDD.n8300 0.00476
R16713 DVDD.n8300 DVDD.n1653 0.00476
R16714 DVDD.n8296 DVDD.n1653 0.00476
R16715 DVDD.n8296 DVDD.n8295 0.00476
R16716 DVDD.n8295 DVDD.n8294 0.00476
R16717 DVDD.n8294 DVDD.n1659 0.00476
R16718 DVDD.n1920 DVDD.n1659 0.00476
R16719 DVDD.n1922 DVDD.n1920 0.00476
R16720 DVDD.n8081 DVDD.n1915 0.00476
R16721 DVDD.n8085 DVDD.n1915 0.00476
R16722 DVDD.n8085 DVDD.n1913 0.00476
R16723 DVDD.n8089 DVDD.n1913 0.00476
R16724 DVDD.n8089 DVDD.n1911 0.00476
R16725 DVDD.n8093 DVDD.n1911 0.00476
R16726 DVDD.n8093 DVDD.n1909 0.00476
R16727 DVDD.n8098 DVDD.n1909 0.00476
R16728 DVDD.n8098 DVDD.n1907 0.00476
R16729 DVDD.n8102 DVDD.n1907 0.00476
R16730 DVDD.n8103 DVDD.n8102 0.00476
R16731 DVDD.n8103 DVDD.n1905 0.00476
R16732 DVDD.n8107 DVDD.n1905 0.00476
R16733 DVDD.n8107 DVDD.n1852 0.00476
R16734 DVDD.n8122 DVDD.n1852 0.00476
R16735 DVDD.n8122 DVDD.n1850 0.00476
R16736 DVDD.n8126 DVDD.n1850 0.00476
R16737 DVDD.n8126 DVDD.n1848 0.00476
R16738 DVDD.n8130 DVDD.n1848 0.00476
R16739 DVDD.n8130 DVDD.n1846 0.00476
R16740 DVDD.n8134 DVDD.n1846 0.00476
R16741 DVDD.n8134 DVDD.n1844 0.00476
R16742 DVDD.n8138 DVDD.n1844 0.00476
R16743 DVDD.n8153 DVDD.n8142 0.00476
R16744 DVDD.n8155 DVDD.n8153 0.00476
R16745 DVDD.n8155 DVDD.n1839 0.00476
R16746 DVDD.n8160 DVDD.n1839 0.00476
R16747 DVDD.n8160 DVDD.n1837 0.00476
R16748 DVDD.n8164 DVDD.n1837 0.00476
R16749 DVDD.n8165 DVDD.n8164 0.00476
R16750 DVDD.n8165 DVDD.n1835 0.00476
R16751 DVDD.n8175 DVDD.n1835 0.00476
R16752 DVDD.n8175 DVDD.n8174 0.00476
R16753 DVDD.n7232 DVDD.n7208 0.00476
R16754 DVDD.n7233 DVDD.n7232 0.00476
R16755 DVDD.n7234 DVDD.n7233 0.00476
R16756 DVDD.n7234 DVDD.n7108 0.00476
R16757 DVDD.n7266 DVDD.n7265 0.00476
R16758 DVDD.n7265 DVDD.n7264 0.00476
R16759 DVDD.n7264 DVDD.n7243 0.00476
R16760 DVDD.n7260 DVDD.n7243 0.00476
R16761 DVDD.n7260 DVDD.n7259 0.00476
R16762 DVDD.n7259 DVDD.n7258 0.00476
R16763 DVDD.n7258 DVDD.n7249 0.00476
R16764 DVDD.n7249 DVDD.n1531 0.00476
R16765 DVDD.n8343 DVDD.n8342 0.00476
R16766 DVDD.n8342 DVDD.n8341 0.00476
R16767 DVDD.n8341 DVDD.n1568 0.00476
R16768 DVDD.n8337 DVDD.n1568 0.00476
R16769 DVDD.n8337 DVDD.n8336 0.00476
R16770 DVDD.n8336 DVDD.n8335 0.00476
R16771 DVDD.n8335 DVDD.n1574 0.00476
R16772 DVDD.n8331 DVDD.n1574 0.00476
R16773 DVDD.n8331 DVDD.n8330 0.00476
R16774 DVDD.n8330 DVDD.n8329 0.00476
R16775 DVDD.n8329 DVDD.n1580 0.00476
R16776 DVDD.n8317 DVDD.n8316 0.00476
R16777 DVDD.n8316 DVDD.n8315 0.00476
R16778 DVDD.n8315 DVDD.n1636 0.00476
R16779 DVDD.n8311 DVDD.n1636 0.00476
R16780 DVDD.n8311 DVDD.n8310 0.00476
R16781 DVDD.n8310 DVDD.n8309 0.00476
R16782 DVDD.n8309 DVDD.n1642 0.00476
R16783 DVDD.n8305 DVDD.n1642 0.00476
R16784 DVDD.n8305 DVDD.n8304 0.00476
R16785 DVDD.n8304 DVDD.n8303 0.00476
R16786 DVDD.n8303 DVDD.n1648 0.00476
R16787 DVDD.n8299 DVDD.n1648 0.00476
R16788 DVDD.n8299 DVDD.n8298 0.00476
R16789 DVDD.n8298 DVDD.n8297 0.00476
R16790 DVDD.n8297 DVDD.n1654 0.00476
R16791 DVDD.n8083 DVDD.n8082 0.00476
R16792 DVDD.n8084 DVDD.n8083 0.00476
R16793 DVDD.n8084 DVDD.n1912 0.00476
R16794 DVDD.n8090 DVDD.n1912 0.00476
R16795 DVDD.n8091 DVDD.n8090 0.00476
R16796 DVDD.n8092 DVDD.n8091 0.00476
R16797 DVDD.n8092 DVDD.n1908 0.00476
R16798 DVDD.n8099 DVDD.n1908 0.00476
R16799 DVDD.n8100 DVDD.n8099 0.00476
R16800 DVDD.n8101 DVDD.n8100 0.00476
R16801 DVDD.n8101 DVDD.n1892 0.00476
R16802 DVDD.n8121 DVDD.n1849 0.00476
R16803 DVDD.n8127 DVDD.n1849 0.00476
R16804 DVDD.n8128 DVDD.n8127 0.00476
R16805 DVDD.n8129 DVDD.n8128 0.00476
R16806 DVDD.n8129 DVDD.n1845 0.00476
R16807 DVDD.n8135 DVDD.n1845 0.00476
R16808 DVDD.n8136 DVDD.n8135 0.00476
R16809 DVDD.n8137 DVDD.n8136 0.00476
R16810 DVDD.n8161 DVDD.n1838 0.00476
R16811 DVDD.n8162 DVDD.n8161 0.00476
R16812 DVDD.n8163 DVDD.n8162 0.00476
R16813 DVDD.n8163 DVDD.n1801 0.00476
R16814 DVDD.n7557 DVDD.n2504 0.00476
R16815 DVDD.n7558 DVDD.n7557 0.00476
R16816 DVDD.n7559 DVDD.n7558 0.00476
R16817 DVDD.n7559 DVDD.n2489 0.00476
R16818 DVDD.n7601 DVDD.n2465 0.00476
R16819 DVDD.n7602 DVDD.n7601 0.00476
R16820 DVDD.n7603 DVDD.n7602 0.00476
R16821 DVDD.n7603 DVDD.n2461 0.00476
R16822 DVDD.n7609 DVDD.n2461 0.00476
R16823 DVDD.n7610 DVDD.n7609 0.00476
R16824 DVDD.n7611 DVDD.n7610 0.00476
R16825 DVDD.n7611 DVDD.n2451 0.00476
R16826 DVDD.n7649 DVDD.n2388 0.00476
R16827 DVDD.n7649 DVDD.n7648 0.00476
R16828 DVDD.n7648 DVDD.n7647 0.00476
R16829 DVDD.n7647 DVDD.n7621 0.00476
R16830 DVDD.n7643 DVDD.n7621 0.00476
R16831 DVDD.n7643 DVDD.n7642 0.00476
R16832 DVDD.n7642 DVDD.n7641 0.00476
R16833 DVDD.n7641 DVDD.n7627 0.00476
R16834 DVDD.n7637 DVDD.n7627 0.00476
R16835 DVDD.n7637 DVDD.n7636 0.00476
R16836 DVDD.n7636 DVDD.n2206 0.00476
R16837 DVDD.n7773 DVDD.n2251 0.00476
R16838 DVDD.n7769 DVDD.n2251 0.00476
R16839 DVDD.n7769 DVDD.n7768 0.00476
R16840 DVDD.n7768 DVDD.n7767 0.00476
R16841 DVDD.n7767 DVDD.n2259 0.00476
R16842 DVDD.n7763 DVDD.n2259 0.00476
R16843 DVDD.n7763 DVDD.n7762 0.00476
R16844 DVDD.n7762 DVDD.n7761 0.00476
R16845 DVDD.n7761 DVDD.n2265 0.00476
R16846 DVDD.n7757 DVDD.n2265 0.00476
R16847 DVDD.n7757 DVDD.n7756 0.00476
R16848 DVDD.n7756 DVDD.n7755 0.00476
R16849 DVDD.n7755 DVDD.n2271 0.00476
R16850 DVDD.n7751 DVDD.n2271 0.00476
R16851 DVDD.n7751 DVDD.n7750 0.00476
R16852 DVDD.n8075 DVDD.n8074 0.00476
R16853 DVDD.n8074 DVDD.n8073 0.00476
R16854 DVDD.n8073 DVDD.n1930 0.00476
R16855 DVDD.n8069 DVDD.n1930 0.00476
R16856 DVDD.n8069 DVDD.n8068 0.00476
R16857 DVDD.n8068 DVDD.n8067 0.00476
R16858 DVDD.n8067 DVDD.n1935 0.00476
R16859 DVDD.n8063 DVDD.n1935 0.00476
R16860 DVDD.n8063 DVDD.n8062 0.00476
R16861 DVDD.n8062 DVDD.n8061 0.00476
R16862 DVDD.n8061 DVDD.n1941 0.00476
R16863 DVDD.n8049 DVDD.n1988 0.00476
R16864 DVDD.n8045 DVDD.n1988 0.00476
R16865 DVDD.n8045 DVDD.n8044 0.00476
R16866 DVDD.n8044 DVDD.n8043 0.00476
R16867 DVDD.n8043 DVDD.n1996 0.00476
R16868 DVDD.n8039 DVDD.n1996 0.00476
R16869 DVDD.n8039 DVDD.n8038 0.00476
R16870 DVDD.n8038 DVDD.n8037 0.00476
R16871 DVDD.n8017 DVDD.n8016 0.00476
R16872 DVDD.n8016 DVDD.n8015 0.00476
R16873 DVDD.n8015 DVDD.n2010 0.00476
R16874 DVDD.n8011 DVDD.n2010 0.00476
R16875 DVDD.n7012 DVDD.n7011 0.00476
R16876 DVDD.n7011 DVDD.n7010 0.00476
R16877 DVDD.n7010 DVDD.n2555 0.00476
R16878 DVDD.n7006 DVDD.n2555 0.00476
R16879 DVDD.n6998 DVDD.n6997 0.00476
R16880 DVDD.n6997 DVDD.n6996 0.00476
R16881 DVDD.n6996 DVDD.n2618 0.00476
R16882 DVDD.n6992 DVDD.n2618 0.00476
R16883 DVDD.n6992 DVDD.n6991 0.00476
R16884 DVDD.n6991 DVDD.n6990 0.00476
R16885 DVDD.n6990 DVDD.n2624 0.00476
R16886 DVDD.n6986 DVDD.n2624 0.00476
R16887 DVDD.n6971 DVDD.n6939 0.00476
R16888 DVDD.n6971 DVDD.n6970 0.00476
R16889 DVDD.n6970 DVDD.n6969 0.00476
R16890 DVDD.n6969 DVDD.n6948 0.00476
R16891 DVDD.n6965 DVDD.n6948 0.00476
R16892 DVDD.n6965 DVDD.n6964 0.00476
R16893 DVDD.n6964 DVDD.n6963 0.00476
R16894 DVDD.n6963 DVDD.n6954 0.00476
R16895 DVDD.n6959 DVDD.n6954 0.00476
R16896 DVDD.n6959 DVDD.n2204 0.00476
R16897 DVDD.n7787 DVDD.n2204 0.00476
R16898 DVDD.n7813 DVDD.n2167 0.00476
R16899 DVDD.n7814 DVDD.n7813 0.00476
R16900 DVDD.n7815 DVDD.n7814 0.00476
R16901 DVDD.n7815 DVDD.n2163 0.00476
R16902 DVDD.n7821 DVDD.n2163 0.00476
R16903 DVDD.n7822 DVDD.n7821 0.00476
R16904 DVDD.n7823 DVDD.n7822 0.00476
R16905 DVDD.n7823 DVDD.n2159 0.00476
R16906 DVDD.n7829 DVDD.n2159 0.00476
R16907 DVDD.n7830 DVDD.n7829 0.00476
R16908 DVDD.n7831 DVDD.n7830 0.00476
R16909 DVDD.n7831 DVDD.n2155 0.00476
R16910 DVDD.n7837 DVDD.n2155 0.00476
R16911 DVDD.n7838 DVDD.n7837 0.00476
R16912 DVDD.n7843 DVDD.n7838 0.00476
R16913 DVDD.n7860 DVDD.n7859 0.00476
R16914 DVDD.n7861 DVDD.n7860 0.00476
R16915 DVDD.n7861 DVDD.n2112 0.00476
R16916 DVDD.n7867 DVDD.n2112 0.00476
R16917 DVDD.n7868 DVDD.n7867 0.00476
R16918 DVDD.n7869 DVDD.n7868 0.00476
R16919 DVDD.n7869 DVDD.n2108 0.00476
R16920 DVDD.n7876 DVDD.n2108 0.00476
R16921 DVDD.n7877 DVDD.n7876 0.00476
R16922 DVDD.n7878 DVDD.n7877 0.00476
R16923 DVDD.n7878 DVDD.n2097 0.00476
R16924 DVDD.n7894 DVDD.n2070 0.00476
R16925 DVDD.n7900 DVDD.n2070 0.00476
R16926 DVDD.n7901 DVDD.n7900 0.00476
R16927 DVDD.n7902 DVDD.n7901 0.00476
R16928 DVDD.n7902 DVDD.n2066 0.00476
R16929 DVDD.n7908 DVDD.n2066 0.00476
R16930 DVDD.n7909 DVDD.n7908 0.00476
R16931 DVDD.n7910 DVDD.n7909 0.00476
R16932 DVDD.n7936 DVDD.n2060 0.00476
R16933 DVDD.n7937 DVDD.n7936 0.00476
R16934 DVDD.n7938 DVDD.n7937 0.00476
R16935 DVDD.n7938 DVDD.n2030 0.00476
R16936 DVDD.n5523 DVDD.n5522 0.00476
R16937 DVDD.n5522 DVDD.n5521 0.00476
R16938 DVDD.n5521 DVDD.n5512 0.00476
R16939 DVDD.n5512 DVDD.n3026 0.00476
R16940 DVDD.n6745 DVDD.n6744 0.00476
R16941 DVDD.n6744 DVDD.n6743 0.00476
R16942 DVDD.n6743 DVDD.n3065 0.00476
R16943 DVDD.n6739 DVDD.n3065 0.00476
R16944 DVDD.n6739 DVDD.n6738 0.00476
R16945 DVDD.n6738 DVDD.n6737 0.00476
R16946 DVDD.n6737 DVDD.n3070 0.00476
R16947 DVDD.n6733 DVDD.n3070 0.00476
R16948 DVDD.n6725 DVDD.n2672 0.00476
R16949 DVDD.n6725 DVDD.n6724 0.00476
R16950 DVDD.n6724 DVDD.n6723 0.00476
R16951 DVDD.n6723 DVDD.n3081 0.00476
R16952 DVDD.n6719 DVDD.n3081 0.00476
R16953 DVDD.n6719 DVDD.n6718 0.00476
R16954 DVDD.n6718 DVDD.n6717 0.00476
R16955 DVDD.n6717 DVDD.n3087 0.00476
R16956 DVDD.n6713 DVDD.n3087 0.00476
R16957 DVDD.n6713 DVDD.n6712 0.00476
R16958 DVDD.n6712 DVDD.n6711 0.00476
R16959 DVDD.n6700 DVDD.n3186 0.00476
R16960 DVDD.n6696 DVDD.n3186 0.00476
R16961 DVDD.n6696 DVDD.n6695 0.00476
R16962 DVDD.n6695 DVDD.n6694 0.00476
R16963 DVDD.n6694 DVDD.n3197 0.00476
R16964 DVDD.n6690 DVDD.n3197 0.00476
R16965 DVDD.n6690 DVDD.n6689 0.00476
R16966 DVDD.n6689 DVDD.n6688 0.00476
R16967 DVDD.n6688 DVDD.n3203 0.00476
R16968 DVDD.n6684 DVDD.n3203 0.00476
R16969 DVDD.n6684 DVDD.n6683 0.00476
R16970 DVDD.n6683 DVDD.n6682 0.00476
R16971 DVDD.n6682 DVDD.n3209 0.00476
R16972 DVDD.n6678 DVDD.n3209 0.00476
R16973 DVDD.n6678 DVDD.n6677 0.00476
R16974 DVDD.n6668 DVDD.n3314 0.00476
R16975 DVDD.n6664 DVDD.n3314 0.00476
R16976 DVDD.n6664 DVDD.n6663 0.00476
R16977 DVDD.n6663 DVDD.n6662 0.00476
R16978 DVDD.n6662 DVDD.n3320 0.00476
R16979 DVDD.n6658 DVDD.n3320 0.00476
R16980 DVDD.n6658 DVDD.n6657 0.00476
R16981 DVDD.n6657 DVDD.n6656 0.00476
R16982 DVDD.n6656 DVDD.n3326 0.00476
R16983 DVDD.n6652 DVDD.n3326 0.00476
R16984 DVDD.n6652 DVDD.n6651 0.00476
R16985 DVDD.n6644 DVDD.n3364 0.00476
R16986 DVDD.n6640 DVDD.n3364 0.00476
R16987 DVDD.n6640 DVDD.n6639 0.00476
R16988 DVDD.n6639 DVDD.n6638 0.00476
R16989 DVDD.n6638 DVDD.n3377 0.00476
R16990 DVDD.n6634 DVDD.n3377 0.00476
R16991 DVDD.n6634 DVDD.n6633 0.00476
R16992 DVDD.n6633 DVDD.n6632 0.00476
R16993 DVDD.n6612 DVDD.n6611 0.00476
R16994 DVDD.n6611 DVDD.n6610 0.00476
R16995 DVDD.n6610 DVDD.n3390 0.00476
R16996 DVDD.n6606 DVDD.n3390 0.00476
R16997 DVDD.n5415 DVDD.n5414 0.00476
R16998 DVDD.n5414 DVDD.n5412 0.00476
R16999 DVDD.n5412 DVDD.n5410 0.00476
R17000 DVDD.n5410 DVDD.n5381 0.00476
R17001 DVDD.n5406 DVDD.n5381 0.00476
R17002 DVDD.n5406 DVDD.n5405 0.00476
R17003 DVDD.n5405 DVDD.n5404 0.00476
R17004 DVDD.n5404 DVDD.n5403 0.00476
R17005 DVDD.n5403 DVDD.n5402 0.00476
R17006 DVDD.n5402 DVDD.n4449 0.00476
R17007 DVDD.n5711 DVDD.n4447 0.00476
R17008 DVDD.n5715 DVDD.n4447 0.00476
R17009 DVDD.n5715 DVDD.n4445 0.00476
R17010 DVDD.n5719 DVDD.n4445 0.00476
R17011 DVDD.n5719 DVDD.n4443 0.00476
R17012 DVDD.n5723 DVDD.n4443 0.00476
R17013 DVDD.n5723 DVDD.n4441 0.00476
R17014 DVDD.n5727 DVDD.n4441 0.00476
R17015 DVDD.n5727 DVDD.n4439 0.00476
R17016 DVDD.n5732 DVDD.n4439 0.00476
R17017 DVDD.n5733 DVDD.n5732 0.00476
R17018 DVDD.n5734 DVDD.n5733 0.00476
R17019 DVDD.n5734 DVDD.n4436 0.00476
R17020 DVDD.n5738 DVDD.n4436 0.00476
R17021 DVDD.n5738 DVDD.n4434 0.00476
R17022 DVDD.n5742 DVDD.n4434 0.00476
R17023 DVDD.n5742 DVDD.n4432 0.00476
R17024 DVDD.n5746 DVDD.n4432 0.00476
R17025 DVDD.n5746 DVDD.n4430 0.00476
R17026 DVDD.n5751 DVDD.n4430 0.00476
R17027 DVDD.n5751 DVDD.n4428 0.00476
R17028 DVDD.n5755 DVDD.n4428 0.00476
R17029 DVDD.n5756 DVDD.n5755 0.00476
R17030 DVDD.n6104 DVDD.n4390 0.00476
R17031 DVDD.n6104 DVDD.n4304 0.00476
R17032 DVDD.n6115 DVDD.n4304 0.00476
R17033 DVDD.n6115 DVDD.n4302 0.00476
R17034 DVDD.n6119 DVDD.n4302 0.00476
R17035 DVDD.n6119 DVDD.n4300 0.00476
R17036 DVDD.n6123 DVDD.n4300 0.00476
R17037 DVDD.n6123 DVDD.n4298 0.00476
R17038 DVDD.n6127 DVDD.n4298 0.00476
R17039 DVDD.n6127 DVDD.n4296 0.00476
R17040 DVDD.n6131 DVDD.n4296 0.00476
R17041 DVDD.n6131 DVDD.n4294 0.00476
R17042 DVDD.n6135 DVDD.n4294 0.00476
R17043 DVDD.n6135 DVDD.n4292 0.00476
R17044 DVDD.n6139 DVDD.n4292 0.00476
R17045 DVDD.n6139 DVDD.n4290 0.00476
R17046 DVDD.n6143 DVDD.n4290 0.00476
R17047 DVDD.n6143 DVDD.n4288 0.00476
R17048 DVDD.n6147 DVDD.n4288 0.00476
R17049 DVDD.n6147 DVDD.n4286 0.00476
R17050 DVDD.n6151 DVDD.n4286 0.00476
R17051 DVDD.n6151 DVDD.n3945 0.00476
R17052 DVDD.n6157 DVDD.n3945 0.00476
R17053 DVDD.n6161 DVDD.n3911 0.00476
R17054 DVDD.n6165 DVDD.n3911 0.00476
R17055 DVDD.n6165 DVDD.n3909 0.00476
R17056 DVDD.n6169 DVDD.n3909 0.00476
R17057 DVDD.n6169 DVDD.n3907 0.00476
R17058 DVDD.n6173 DVDD.n3907 0.00476
R17059 DVDD.n6173 DVDD.n3905 0.00476
R17060 DVDD.n6177 DVDD.n3905 0.00476
R17061 DVDD.n6177 DVDD.n3903 0.00476
R17062 DVDD.n6182 DVDD.n3903 0.00476
R17063 DVDD.n6182 DVDD.n3901 0.00476
R17064 DVDD.n6187 DVDD.n3901 0.00476
R17065 DVDD.n6189 DVDD.n6187 0.00476
R17066 DVDD.n6190 DVDD.n6189 0.00476
R17067 DVDD.n6190 DVDD.n3899 0.00476
R17068 DVDD.n6194 DVDD.n3899 0.00476
R17069 DVDD.n6194 DVDD.n3898 0.00476
R17070 DVDD.n6198 DVDD.n3898 0.00476
R17071 DVDD.n6198 DVDD.n3896 0.00476
R17072 DVDD.n6202 DVDD.n3896 0.00476
R17073 DVDD.n6202 DVDD.n3894 0.00476
R17074 DVDD.n6207 DVDD.n3894 0.00476
R17075 DVDD.n6207 DVDD.n3510 0.00476
R17076 DVDD.n6423 DVDD.n6422 0.00476
R17077 DVDD.n6422 DVDD.n6409 0.00476
R17078 DVDD.n6409 DVDD.n6407 0.00476
R17079 DVDD.n6407 DVDD.n3515 0.00476
R17080 DVDD.n6403 DVDD.n3515 0.00476
R17081 DVDD.n6403 DVDD.n6402 0.00476
R17082 DVDD.n6402 DVDD.n6401 0.00476
R17083 DVDD.n6401 DVDD.n3521 0.00476
R17084 DVDD.n6388 DVDD.n3521 0.00476
R17085 DVDD.n6395 DVDD.n6388 0.00476
R17086 DVDD.n5409 DVDD.n5408 0.00476
R17087 DVDD.n5408 DVDD.n5407 0.00476
R17088 DVDD.n5407 DVDD.n5382 0.00476
R17089 DVDD.n5382 DVDD.n2963 0.00476
R17090 DVDD.n5710 DVDD.n4446 0.00476
R17091 DVDD.n5716 DVDD.n4446 0.00476
R17092 DVDD.n5717 DVDD.n5716 0.00476
R17093 DVDD.n5718 DVDD.n5717 0.00476
R17094 DVDD.n5718 DVDD.n4442 0.00476
R17095 DVDD.n5724 DVDD.n4442 0.00476
R17096 DVDD.n5725 DVDD.n5724 0.00476
R17097 DVDD.n5726 DVDD.n5725 0.00476
R17098 DVDD.n4435 DVDD.n2820 0.00476
R17099 DVDD.n5739 DVDD.n4435 0.00476
R17100 DVDD.n5740 DVDD.n5739 0.00476
R17101 DVDD.n5741 DVDD.n5740 0.00476
R17102 DVDD.n5741 DVDD.n4431 0.00476
R17103 DVDD.n5747 DVDD.n4431 0.00476
R17104 DVDD.n5748 DVDD.n5747 0.00476
R17105 DVDD.n5750 DVDD.n5748 0.00476
R17106 DVDD.n5750 DVDD.n5749 0.00476
R17107 DVDD.n5749 DVDD.n4427 0.00476
R17108 DVDD.n5757 DVDD.n4427 0.00476
R17109 DVDD.n6120 DVDD.n4301 0.00476
R17110 DVDD.n6121 DVDD.n6120 0.00476
R17111 DVDD.n6122 DVDD.n6121 0.00476
R17112 DVDD.n6122 DVDD.n4297 0.00476
R17113 DVDD.n6128 DVDD.n4297 0.00476
R17114 DVDD.n6129 DVDD.n6128 0.00476
R17115 DVDD.n6130 DVDD.n6129 0.00476
R17116 DVDD.n6130 DVDD.n4293 0.00476
R17117 DVDD.n6136 DVDD.n4293 0.00476
R17118 DVDD.n6137 DVDD.n6136 0.00476
R17119 DVDD.n6138 DVDD.n6137 0.00476
R17120 DVDD.n6138 DVDD.n4289 0.00476
R17121 DVDD.n6144 DVDD.n4289 0.00476
R17122 DVDD.n6145 DVDD.n6144 0.00476
R17123 DVDD.n6146 DVDD.n6145 0.00476
R17124 DVDD.n6163 DVDD.n6162 0.00476
R17125 DVDD.n6164 DVDD.n6163 0.00476
R17126 DVDD.n6164 DVDD.n3908 0.00476
R17127 DVDD.n6170 DVDD.n3908 0.00476
R17128 DVDD.n6171 DVDD.n6170 0.00476
R17129 DVDD.n6172 DVDD.n6171 0.00476
R17130 DVDD.n6172 DVDD.n3904 0.00476
R17131 DVDD.n6178 DVDD.n3904 0.00476
R17132 DVDD.n6179 DVDD.n6178 0.00476
R17133 DVDD.n6181 DVDD.n6179 0.00476
R17134 DVDD.n6181 DVDD.n6180 0.00476
R17135 DVDD.n6195 DVDD.n3808 0.00476
R17136 DVDD.n6196 DVDD.n6195 0.00476
R17137 DVDD.n6197 DVDD.n6196 0.00476
R17138 DVDD.n6197 DVDD.n3895 0.00476
R17139 DVDD.n6203 DVDD.n3895 0.00476
R17140 DVDD.n6204 DVDD.n6203 0.00476
R17141 DVDD.n6206 DVDD.n6204 0.00476
R17142 DVDD.n6206 DVDD.n6205 0.00476
R17143 DVDD.n6406 DVDD.n6405 0.00476
R17144 DVDD.n6405 DVDD.n6404 0.00476
R17145 DVDD.n6404 DVDD.n3516 0.00476
R17146 DVDD.n6400 DVDD.n3516 0.00476
R17147 DVDD.n9322 DVDD.n427 0.00476
R17148 DVDD.n9323 DVDD.n9322 0.00476
R17149 DVDD.n9324 DVDD.n9323 0.00476
R17150 DVDD.n9346 DVDD.n9345 0.00476
R17151 DVDD.n9345 DVDD.n9344 0.00476
R17152 DVDD.n9344 DVDD.n9330 0.00476
R17153 DVDD.n9340 DVDD.n9330 0.00476
R17154 DVDD.n9339 DVDD.n9338 0.00476
R17155 DVDD.n9338 DVDD.n9332 0.00476
R17156 DVDD.n9334 DVDD.n9332 0.00476
R17157 DVDD.n9334 DVDD.n9333 0.00476
R17158 DVDD.n9577 DVDD.n9576 0.00476
R17159 DVDD.n9576 DVDD.n9575 0.00476
R17160 DVDD.n9575 DVDD.n204 0.00476
R17161 DVDD.n9571 DVDD.n204 0.00476
R17162 DVDD.n9570 DVDD.n9569 0.00476
R17163 DVDD.n9569 DVDD.n209 0.00476
R17164 DVDD.n9565 DVDD.n209 0.00476
R17165 DVDD.n9565 DVDD.n9564 0.00476
R17166 DVDD.n5297 DVDD.n226 0.00476
R17167 DVDD.n5300 DVDD.n5297 0.00476
R17168 DVDD.n5301 DVDD.n5300 0.00476
R17169 DVDD.n9469 DVDD.n9468 0.00476
R17170 DVDD.n9468 DVDD.n292 0.00476
R17171 DVDD.n417 DVDD.n292 0.00476
R17172 DVDD.n9455 DVDD.n309 0.00476
R17173 DVDD.n9455 DVDD.n9454 0.00476
R17174 DVDD.n9454 DVDD.n312 0.00476
R17175 DVDD.n9443 DVDD.n312 0.00476
R17176 DVDD.n9442 DVDD.n9441 0.00476
R17177 DVDD.n9441 DVDD.n328 0.00476
R17178 DVDD.n9428 DVDD.n328 0.00476
R17179 DVDD.n9429 DVDD.n9428 0.00476
R17180 DVDD.n360 DVDD.n280 0.00476
R17181 DVDD.n9485 DVDD.n280 0.00476
R17182 DVDD.n9485 DVDD.n278 0.00476
R17183 DVDD.n9489 DVDD.n278 0.00476
R17184 DVDD.n9498 DVDD.n271 0.00476
R17185 DVDD.n9498 DVDD.n269 0.00476
R17186 DVDD.n9502 DVDD.n269 0.00476
R17187 DVDD.n9502 DVDD.n221 0.00476
R17188 DVDD.n9558 DVDD.n222 0.00476
R17189 DVDD.n9558 DVDD.n241 0.00476
R17190 DVDD.n253 DVDD.n241 0.00476
R17191 DVDD.n8785 DVDD.n8781 0.00476
R17192 DVDD.n8785 DVDD.n8784 0.00476
R17193 DVDD.n8784 DVDD.n8783 0.00476
R17194 DVDD.n960 DVDD.n959 0.00476
R17195 DVDD.n963 DVDD.n960 0.00476
R17196 DVDD.n964 DVDD.n963 0.00476
R17197 DVDD.n966 DVDD.n964 0.00476
R17198 DVDD.n975 DVDD.n957 0.00476
R17199 DVDD.n975 DVDD.n974 0.00476
R17200 DVDD.n974 DVDD.n973 0.00476
R17201 DVDD.n973 DVDD.n972 0.00476
R17202 DVDD.n1019 DVDD.n1018 0.00476
R17203 DVDD.n1019 DVDD.n1017 0.00476
R17204 DVDD.n1023 DVDD.n1017 0.00476
R17205 DVDD.n1024 DVDD.n1023 0.00476
R17206 DVDD.n1025 DVDD.n1015 0.00476
R17207 DVDD.n1031 DVDD.n1015 0.00476
R17208 DVDD.n1031 DVDD.n1030 0.00476
R17209 DVDD.n1030 DVDD.n216 0.00476
R17210 DVDD.n3585 DVDD.n215 0.00476
R17211 DVDD.n3590 DVDD.n3585 0.00476
R17212 DVDD.n3590 DVDD.n3589 0.00476
R17213 DVDD.n4109 DVDD.n4108 0.00476
R17214 DVDD.n4108 DVDD.n4105 0.00476
R17215 DVDD.n4105 DVDD.n4104 0.00476
R17216 DVDD.n4093 DVDD.n4018 0.00476
R17217 DVDD.n4093 DVDD.n4019 0.00476
R17218 DVDD.n4089 DVDD.n4019 0.00476
R17219 DVDD.n4089 DVDD.n4088 0.00476
R17220 DVDD.n4087 DVDD.n4024 0.00476
R17221 DVDD.n4083 DVDD.n4024 0.00476
R17222 DVDD.n4083 DVDD.n4082 0.00476
R17223 DVDD.n4082 DVDD.n4081 0.00476
R17224 DVDD.n3990 DVDD.n3989 0.00476
R17225 DVDD.n4125 DVDD.n3990 0.00476
R17226 DVDD.n4125 DVDD.n3987 0.00476
R17227 DVDD.n4129 DVDD.n3987 0.00476
R17228 DVDD.n4138 DVDD.n3980 0.00476
R17229 DVDD.n4138 DVDD.n3978 0.00476
R17230 DVDD.n4142 DVDD.n3978 0.00476
R17231 DVDD.n4142 DVDD.n219 0.00476
R17232 DVDD.n4213 DVDD.n218 0.00476
R17233 DVDD.n4213 DVDD.n4150 0.00476
R17234 DVDD.n4209 DVDD.n4150 0.00476
R17235 DVDD.n5899 DVDD.n5829 0.00471875
R17236 DVDD.n5482 DVDD.n4459 0.00471875
R17237 DVDD.n4450 DVDD.n3001 0.00471875
R17238 DVDD.n6234 DVDD.n3882 0.0047
R17239 DVDD.n6159 DVDD.n3943 0.004625
R17240 DVDD.n9382 DVDD.n153 0.0045748
R17241 DVDD.n9384 DVDD.n9383 0.0045748
R17242 DVDD.n9386 DVDD.n168 0.0045748
R17243 DVDD.n9389 DVDD.n171 0.0045748
R17244 DVDD.n9390 DVDD.n377 0.0045748
R17245 DVDD.n9424 DVDD.n9423 0.0045748
R17246 DVDD.n9420 DVDD.n378 0.0045748
R17247 DVDD.n9419 DVDD.n381 0.0045748
R17248 DVDD.n4522 DVDD.n386 0.0045748
R17249 DVDD.n4524 DVDD.n4523 0.0045748
R17250 DVDD.n5267 DVDD.n4520 0.0045748
R17251 DVDD.n8814 DVDD.n63 0.0045748
R17252 DVDD.n3854 DVDD.n3563 0.0045748
R17253 DVDD.n6534 DVDD.n3354 0.0045748
R17254 DVDD.n6502 DVDD.n2078 0.0045748
R17255 DVDD.n9086 DVDD.n524 0.0045748
R17256 DVDD.n6014 DVDD.n3960 0.0045748
R17257 DVDD.n3236 DVDD.n3215 0.0045748
R17258 DVDD.n3265 DVDD.n2125 0.0045748
R17259 DVDD.n4929 DVDD.n487 0.0045748
R17260 DVDD.n5781 DVDD.n4307 0.0045748
R17261 DVDD.n3131 DVDD.n3119 0.0045748
R17262 DVDD.n3156 DVDD.n2175 0.0045748
R17263 DVDD.n9255 DVDD.n463 0.0045748
R17264 DVDD.n2841 DVDD.n2822 0.0045748
R17265 DVDD.n2719 DVDD.n2669 0.0045748
R17266 DVDD.n2686 DVDD.n2648 0.0045748
R17267 DVDD DVDD.n3485 0.00453415
R17268 DVDD.n7790 DVDD.n2198 0.0045
R17269 DVDD.n3315 DVDD.n1924 0.0045
R17270 DVDD.n7597 DVDD.n2467 0.0045
R17271 DVDD.n7790 DVDD.n2200 0.0045
R17272 DVDD.n7597 DVDD.n2468 0.0045
R17273 DVDD.n2200 DVDD.n2199 0.0045
R17274 DVDD.n8140 DVDD.n1842 0.0045
R17275 DVDD.n8078 DVDD.n1924 0.0045
R17276 DVDD.n8079 DVDD.n8078 0.0045
R17277 DVDD.n7913 DVDD.n2063 0.0045
R17278 DVDD.n7913 DVDD.n1842 0.0045
R17279 DVDD.n6748 DVDD.n2467 0.0045
R17280 DVDD.n1116 DVDD.n1102 0.00449375
R17281 DVDD.n6426 DVDD.n1116 0.00449375
R17282 DVDD.n3473 DVDD.n3420 0.00449375
R17283 DVDD.n6442 DVDD.n3420 0.00449375
R17284 DVDD.n5922 DVDD.n5921 0.00449375
R17285 DVDD.n6063 DVDD.n5922 0.00449375
R17286 DVDD.n6445 DVDD.n6444 0.0044
R17287 DVDD.n6101 DVDD.n6100 0.004325
R17288 DVDD.n9691 DVDD.n9690 0.00429286
R17289 DVDD.n5892 DVDD.n5829 0.00426875
R17290 DVDD.n5660 DVDD.n4459 0.00426875
R17291 DVDD.n5678 DVDD.n3001 0.00426875
R17292 DVDD.n3497 DVDD.n3496 0.004246
R17293 DVDD.n723 DVDD.n579 0.00422047
R17294 DVDD.n8804 DVDD.n61 0.00422047
R17295 DVDD.n8745 DVDD.n8744 0.00422047
R17296 DVDD.n8681 DVDD.n1042 0.00422047
R17297 DVDD.n3844 DVDD.n3565 0.00422047
R17298 DVDD.n6321 DVDD.n3867 0.00422047
R17299 DVDD.n6512 DVDD.n2080 0.00422047
R17300 DVDD.n9014 DVDD.n550 0.00422047
R17301 DVDD.n532 DVDD.n521 0.00422047
R17302 DVDD.n4058 DVDD.n4030 0.00422047
R17303 DVDD.n4216 DVDD.n4147 0.00422047
R17304 DVDD.n6024 DVDD.n3962 0.00422047
R17305 DVDD.n6055 DVDD.n5930 0.00422047
R17306 DVDD.n3275 DVDD.n2123 0.00422047
R17307 DVDD.n4877 DVDD.n4867 0.00422047
R17308 DVDD.n4919 DVDD.n485 0.00422047
R17309 DVDD.n339 DVDD.n331 0.00422047
R17310 DVDD.n9507 DVDD.n245 0.00422047
R17311 DVDD.n5791 DVDD.n4309 0.00422047
R17312 DVDD.n5824 DVDD.n5823 0.00422047
R17313 DVDD.n3166 DVDD.n2177 0.00422047
R17314 DVDD.n5158 DVDD.n4572 0.00422047
R17315 DVDD.n9249 DVDD.n461 0.00422047
R17316 DVDD.n9591 DVDD.n156 0.00422047
R17317 DVDD.n6792 DVDD.n2892 0.00422047
R17318 DVDD.n2851 DVDD.n2824 0.00422047
R17319 DVDD.n6861 DVDD.n2792 0.00422047
R17320 DVDD.n2696 DVDD.n2645 0.00422047
R17321 DVDD.n9316 DVDD.n434 0.00422
R17322 DVDD.n9599 DVDD.n145 0.00422
R17323 DVDD.n9596 DVDD.n152 0.00422
R17324 DVDD.n9415 DVDD.n385 0.00422
R17325 DVDD.n5272 DVDD.n4516 0.00422
R17326 DVDD.n6777 DVDD.n2906 0.00422
R17327 DVDD.n4009 DVDD.n3999 0.00422
R17328 DVDD.n4046 DVDD.n4045 0.00422
R17329 DVDD.n4059 DVDD.n4031 0.00422
R17330 DVDD.n4123 DVDD.n3992 0.00422
R17331 DVDD.n4136 DVDD.n3983 0.00422
R17332 DVDD.n4207 DVDD.n4151 0.00422
R17333 DVDD.n293 DVDD.n290 0.00422
R17334 DVDD.n9445 DVDD.n322 0.00422
R17335 DVDD.n337 DVDD.n329 0.00422
R17336 DVDD.n9483 DVDD.n282 0.00422
R17337 DVDD.n9496 DVDD.n274 0.00422
R17338 DVDD.n9548 DVDD.n9547 0.00422
R17339 DVDD.n9627 DVDD.n85 0.00422
R17340 DVDD.n8753 DVDD.n867 0.00422
R17341 DVDD.n8749 DVDD.n871 0.00422
R17342 DVDD.n995 DVDD.n919 0.00422
R17343 DVDD.n8700 DVDD.n1003 0.00422
R17344 DVDD.n8670 DVDD.n1052 0.00422
R17345 DVDD.n7091 DVDD.n7068 0.00416429
R17346 DVDD.n7484 DVDD.n7304 0.00416429
R17347 DVDD.n7460 DVDD.n1512 0.00416429
R17348 DVDD.n7425 DVDD.n7369 0.00416429
R17349 DVDD.n4714 DVDD.n4713 0.00416429
R17350 DVDD.n4822 DVDD.n4821 0.00416429
R17351 DVDD.n5109 DVDD.n4570 0.00416429
R17352 DVDD.n5080 DVDD.n5029 0.00416429
R17353 DVDD.n4759 DVDD.n4543 0.00416429
R17354 DVDD.n4816 DVDD.n4742 0.00416429
R17355 DVDD.n9237 DVDD.n456 0.00416429
R17356 DVDD.n9208 DVDD.n499 0.00416429
R17357 DVDD.n8663 DVDD.n1058 0.00415625
R17358 DVDD.n9329 DVDD.n137 0.00413
R17359 DVDD.n9589 DVDD.n166 0.00413
R17360 DVDD.n5303 DVDD.n5302 0.00413
R17361 DVDD.n4042 DVDD.n4021 0.00413
R17362 DVDD.n4061 DVDD.n4060 0.00413
R17363 DVDD.n4208 DVDD.n4153 0.00413
R17364 DVDD.n9452 DVDD.n313 0.00413
R17365 DVDD.n9440 DVDD.n9439 0.00413
R17366 DVDD.n252 DVDD.n251 0.00413
R17367 DVDD.n942 DVDD.n866 0.00413
R17368 DVDD.n977 DVDD.n976 0.00413
R17369 DVDD.n3634 DVDD.n1051 0.00413
R17370 DVDD DVDD.n193 0.00408591
R17371 DVDD.n9319 DVDD.n430 0.00407
R17372 DVDD.n394 DVDD.n393 0.00407
R17373 DVDD.n5269 DVDD.n208 0.00407
R17374 DVDD.n4111 DVDD.n4110 0.00407
R17375 DVDD.n4131 DVDD.n3985 0.00407
R17376 DVDD.n4137 DVDD.n3981 0.00407
R17377 DVDD.n9471 DVDD.n9470 0.00407
R17378 DVDD.n9491 DVDD.n276 0.00407
R17379 DVDD.n9497 DVDD.n272 0.00407
R17380 DVDD.n8788 DVDD.n84 0.00407
R17381 DVDD.n8706 DVDD.n906 0.00407
R17382 DVDD.n8703 DVDD.n912 0.00407
R17383 DVDD.n7735 DVDD.n2094 0.00404331
R17384 DVDD.n7852 DVDD.n2150 0.00404331
R17385 DVDD.n2369 DVDD.n2191 0.00404331
R17386 DVDD.n7685 DVDD.n2355 0.00404331
R17387 DVDD.n6630 DVDD.n6629 0.00404
R17388 DVDD.n7915 DVDD.n2004 0.00404
R17389 DVDD.n8035 DVDD.n8034 0.00404
R17390 DVDD.n8142 DVDD.n1841 0.00404
R17391 DVDD.n6424 DVDD.n6423 0.00404
R17392 DVDD.n5681 DVDD.n4448 0.004025
R17393 DVDD.n6601 DVDD 0.00392
R17394 DVDD.n7949 DVDD 0.00392
R17395 DVDD.n8006 DVDD 0.00392
R17396 DVDD.n8174 DVDD 0.00392
R17397 DVDD.n6395 DVDD 0.00392
R17398 DVDD.n8287 DVDD.n1712 0.00390714
R17399 DVDD.n8283 DVDD.n1704 0.00390714
R17400 DVDD.n8252 DVDD.n1746 0.00390714
R17401 DVDD.n8250 DVDD.n1758 0.00390714
R17402 DVDD.n8648 DVDD.n1280 0.00390714
R17403 DVDD.n8226 DVDD.n1273 0.00390714
R17404 DVDD.n8211 DVDD.n1784 0.00390714
R17405 DVDD.n8208 DVDD.n1790 0.00390714
R17406 DVDD.n9013 DVDD.n8971 0.00390714
R17407 DVDD.n559 DVDD.n551 0.00390714
R17408 DVDD.n8938 DVDD.n582 0.00390714
R17409 DVDD.n596 DVDD.n589 0.00390714
R17410 DVDD.n610 DVDD.n606 0.00390714
R17411 DVDD.n8913 DVDD.n8912 0.00390714
R17412 DVDD.n641 DVDD.n637 0.00390714
R17413 DVDD.n8895 DVDD.n8894 0.00390714
R17414 DVDD.n9175 DVDD.n526 0.00390714
R17415 DVDD.n9173 DVDD.n9126 0.00390714
R17416 DVDD.n73 DVDD.n72 0.00390714
R17417 DVDD.n9648 DVDD.n9647 0.00390714
R17418 DVDD.n9672 DVDD.n9671 0.00390714
R17419 DVDD.n9675 DVDD.n9674 0.00390714
R17420 DVDD.n8754 DVDD.n864 0.00386614
R17421 DVDD.n6266 DVDD.n3342 0.00386614
R17422 DVDD.n4047 DVDD.n4044 0.00386614
R17423 DVDD.n5957 DVDD.n3233 0.00386614
R17424 DVDD.n9450 DVDD.n315 0.00386614
R17425 DVDD.n5855 DVDD.n3107 0.00386614
R17426 DVDD.n144 DVDD.n136 0.00386614
R17427 DVDD.n6917 DVDD.n2736 0.00386614
R17428 DVDD.n7285 DVDD.n7108 0.00383
R17429 DVDD.n8358 DVDD.n1531 0.00383
R17430 DVDD.n8324 DVDD.n8323 0.00383
R17431 DVDD.n7590 DVDD.n2489 0.00383
R17432 DVDD.n7660 DVDD.n2451 0.00383
R17433 DVDD.n7784 DVDD.n2207 0.00383
R17434 DVDD.n7006 DVDD.n7005 0.00383
R17435 DVDD.n6986 DVDD.n6985 0.00383
R17436 DVDD.n7803 DVDD.n2193 0.00383
R17437 DVDD.n6768 DVDD.n3026 0.00383
R17438 DVDD.n6733 DVDD.n2657 0.00383
R17439 DVDD.n6707 DVDD.n6706 0.00383
R17440 DVDD.n6774 DVDD.n2963 0.00383
R17441 DVDD.n5726 DVDD.n2805 0.00383
R17442 DVDD.n5758 DVDD.n4388 0.00383
R17443 DVDD.n4528 DVDD.n428 0.00383
R17444 DVDD.n9418 DVDD.n203 0.00383
R17445 DVDD.n5284 DVDD.n4508 0.00383
R17446 DVDD.n4001 DVDD.n4000 0.00383
R17447 DVDD.n4124 DVDD.n3991 0.00383
R17448 DVDD.n3982 DVDD.n3977 0.00383
R17449 DVDD.n9467 DVDD.n9466 0.00383
R17450 DVDD.n9484 DVDD.n281 0.00383
R17451 DVDD.n273 DVDD.n268 0.00383
R17452 DVDD.n9623 DVDD.n88 0.00383
R17453 DVDD.n8715 DVDD.n894 0.00383
R17454 DVDD.n1034 DVDD.n1032 0.00383
R17455 DVDD.n6667 DVDD.n2117 0.0038
R17456 DVDD.n7858 DVDD.n7856 0.0038
R17457 DVDD.n8076 DVDD.n1927 0.0038
R17458 DVDD.n8081 DVDD.n1917 0.0038
R17459 DVDD.n8082 DVDD.n1916 0.0038
R17460 DVDD.n8075 DVDD.n1929 0.0038
R17461 DVDD.n7859 DVDD.n2116 0.0038
R17462 DVDD.n6669 DVDD.n6668 0.0038
R17463 DVDD.n6161 DVDD.n3913 0.0038
R17464 DVDD.n6162 DVDD.n3912 0.0038
R17465 DVDD DVDD.n228 0.00376574
R17466 DVDD.n9563 DVDD 0.00376574
R17467 DVDD.n9616 DVDD 0.00376574
R17468 DVDD DVDD.n103 0.00376574
R17469 DVDD.n1921 DVDD.n1678 0.00371
R17470 DVDD.n8121 DVDD.n8120 0.00371
R17471 DVDD.n1838 DVDD.n1235 0.00371
R17472 DVDD.n7747 DVDD.n2316 0.00371
R17473 DVDD.n8052 DVDD.n8049 0.00371
R17474 DVDD.n8017 DVDD.n1196 0.00371
R17475 DVDD.n7854 DVDD.n7853 0.00371
R17476 DVDD.n7894 DVDD.n7893 0.00371
R17477 DVDD.n2060 DVDD.n1157 0.00371
R17478 DVDD.n6670 DVDD.n3237 0.00371
R17479 DVDD.n6648 DVDD.n6644 0.00371
R17480 DVDD.n6612 DVDD.n1118 0.00371
R17481 DVDD.n6156 DVDD.n6155 0.00371
R17482 DVDD.n6334 DVDD.n3808 0.00371
R17483 DVDD.n6406 DVDD.n1056 0.00371
R17484 DVDD.n6095 DVDD.n5892 0.00370625
R17485 DVDD.n5660 DVDD.n5659 0.00370625
R17486 DVDD.n3885 DVDD.n3876 0.00365
R17487 DVDD.n6232 DVDD.n3884 0.00365
R17488 DVDD.n7503 DVDD.n7502 0.00365
R17489 DVDD.n7299 DVDD.n7298 0.00365
R17490 DVDD.n8365 DVDD.n1527 0.00365
R17491 DVDD.n7430 DVDD.n7339 0.00365
R17492 DVDD.n809 DVDD.n9 0.00365
R17493 DVDD.n811 DVDD.n8 0.00365
R17494 DVDD.n813 DVDD.n10 0.00365
R17495 DVDD.n815 DVDD.n7 0.00365
R17496 DVDD.n817 DVDD.n11 0.00365
R17497 DVDD.n819 DVDD.n6 0.00365
R17498 DVDD.n821 DVDD.n12 0.00365
R17499 DVDD.n823 DVDD.n5 0.00365
R17500 DVDD.n825 DVDD.n13 0.00365
R17501 DVDD.n14 DVDD.n4 0.00365
R17502 DVDD.n9692 DVDD.n15 0.00365
R17503 DVDD.n4711 DVDD.n4710 0.00365
R17504 DVDD.n4738 DVDD.n4737 0.00365
R17505 DVDD.n4581 DVDD.n4571 0.00365
R17506 DVDD.n5033 DVDD.n5028 0.00365
R17507 DVDD.n4757 DVDD.n4542 0.00365
R17508 DVDD.n4790 DVDD.n4740 0.00365
R17509 DVDD.n466 DVDD.n457 0.00365
R17510 DVDD.n503 DVDD.n498 0.00365
R17511 DVDD.n9328 DVDD.n9327 0.00359
R17512 DVDD.n9586 DVDD.n167 0.00359
R17513 DVDD.n6788 DVDD.n2898 0.00359
R17514 DVDD.n4041 DVDD.n4017 0.00359
R17515 DVDD.n4027 DVDD.n4026 0.00359
R17516 DVDD.n4152 DVDD.n4149 0.00359
R17517 DVDD.n9453 DVDD.n308 0.00359
R17518 DVDD.n346 DVDD.n330 0.00359
R17519 DVDD.n9556 DVDD.n244 0.00359
R17520 DVDD.n8762 DVDD.n853 0.00359
R17521 DVDD.n8738 DVDD.n882 0.00359
R17522 DVDD.n3742 DVDD.n3591 0.00359
R17523 DVDD.n6709 DVDD.n6708 0.00356
R17524 DVDD.n2203 DVDD.n2197 0.00356
R17525 DVDD.n7783 DVDD.n1584 0.00356
R17526 DVDD.n8326 DVDD.n8325 0.00356
R17527 DVDD.n8324 DVDD.n1587 0.00356
R17528 DVDD.n7785 DVDD.n7784 0.00356
R17529 DVDD.n7786 DVDD.n2193 0.00356
R17530 DVDD.n6707 DVDD.n2205 0.00356
R17531 DVDD.n4394 DVDD.n4390 0.00356
R17532 DVDD.n5759 DVDD.n5758 0.00356
R17533 DVDD.n707 DVDD.n577 0.00351181
R17534 DVDD.n9629 DVDD.n81 0.00351181
R17535 DVDD.n918 DVDD.n916 0.00351181
R17536 DVDD.n3828 DVDD.n3811 0.00351181
R17537 DVDD.n9012 DVDD.n9011 0.00351181
R17538 DVDD.n4112 DVDD.n3997 0.00351181
R17539 DVDD.n4122 DVDD.n4121 0.00351181
R17540 DVDD.n6040 DVDD.n3951 0.00351181
R17541 DVDD.n5016 DVDD.n4865 0.00351181
R17542 DVDD.n9472 DVDD.n288 0.00351181
R17543 DVDD.n9482 DVDD.n9481 0.00351181
R17544 DVDD.n5807 DVDD.n4380 0.00351181
R17545 DVDD.n5156 DVDD.n5155 0.00351181
R17546 DVDD.n436 DVDD.n431 0.00351181
R17547 DVDD.n9414 DVDD.n9413 0.00351181
R17548 DVDD.n2867 DVDD.n2812 0.00351181
R17549 DVDD.n3885 DVDD.n3864 0.00348125
R17550 DVDD.n8663 DVDD.n1102 0.00348125
R17551 DVDD.n6426 DVDD.n1096 0.00348125
R17552 DVDD.n6464 DVDD.n3473 0.00348125
R17553 DVDD.n6442 DVDD.n3467 0.00348125
R17554 DVDD.n5921 DVDD.n5917 0.00348125
R17555 DVDD.n6063 DVDD.n6062 0.00348125
R17556 DVDD.n6453 DVDD.n6452 0.00347759
R17557 DVDD.n8697 DVDD.n8696 0.003425
R17558 DVDD.n8712 DVDD.n898 0.003425
R17559 DVDD.n6305 DVDD.n6304 0.003425
R17560 DVDD.n6895 DVDD.n6894 0.003425
R17561 DVDD.n9403 DVDD.n388 0.003425
R17562 DVDD.n4515 DVDD.n4510 0.003425
R17563 DVDD.n9313 DVDD.n442 0.003425
R17564 DVDD.n841 DVDD.n93 0.003425
R17565 DVDD.n6449 DVDD.n3467 0.00336875
R17566 DVDD.n7227 DVDD.n7210 0.00334
R17567 DVDD.n7228 DVDD.n7227 0.00334
R17568 DVDD.n7230 DVDD.n7228 0.00334
R17569 DVDD.n7230 DVDD.n7229 0.00334
R17570 DVDD.n7229 DVDD.n7206 0.00334
R17571 DVDD.n7237 DVDD.n7206 0.00334
R17572 DVDD.n7238 DVDD.n7237 0.00334
R17573 DVDD.n7239 DVDD.n7238 0.00334
R17574 DVDD.n7240 DVDD.n7239 0.00334
R17575 DVDD.n7244 DVDD.n7241 0.00334
R17576 DVDD.n7245 DVDD.n7244 0.00334
R17577 DVDD.n7246 DVDD.n7245 0.00334
R17578 DVDD.n7247 DVDD.n7246 0.00334
R17579 DVDD.n7250 DVDD.n7247 0.00334
R17580 DVDD.n7251 DVDD.n7250 0.00334
R17581 DVDD.n7252 DVDD.n7251 0.00334
R17582 DVDD.n7254 DVDD.n7252 0.00334
R17583 DVDD.n7254 DVDD.n7253 0.00334
R17584 DVDD.n7253 DVDD.n1564 0.00334
R17585 DVDD.n1565 DVDD.n1564 0.00334
R17586 DVDD.n1566 DVDD.n1565 0.00334
R17587 DVDD.n1569 DVDD.n1566 0.00334
R17588 DVDD.n1570 DVDD.n1569 0.00334
R17589 DVDD.n1571 DVDD.n1570 0.00334
R17590 DVDD.n1572 DVDD.n1571 0.00334
R17591 DVDD.n1575 DVDD.n1572 0.00334
R17592 DVDD.n1576 DVDD.n1575 0.00334
R17593 DVDD.n1577 DVDD.n1576 0.00334
R17594 DVDD.n1578 DVDD.n1577 0.00334
R17595 DVDD.n1581 DVDD.n1578 0.00334
R17596 DVDD.n1582 DVDD.n1581 0.00334
R17597 DVDD.n1583 DVDD.n1582 0.00334
R17598 DVDD.n1631 DVDD.n1585 0.00334
R17599 DVDD.n1632 DVDD.n1631 0.00334
R17600 DVDD.n1633 DVDD.n1632 0.00334
R17601 DVDD.n1634 DVDD.n1633 0.00334
R17602 DVDD.n1637 DVDD.n1634 0.00334
R17603 DVDD.n1638 DVDD.n1637 0.00334
R17604 DVDD.n1639 DVDD.n1638 0.00334
R17605 DVDD.n1640 DVDD.n1639 0.00334
R17606 DVDD.n1643 DVDD.n1640 0.00334
R17607 DVDD.n1644 DVDD.n1643 0.00334
R17608 DVDD.n1645 DVDD.n1644 0.00334
R17609 DVDD.n1646 DVDD.n1645 0.00334
R17610 DVDD.n1649 DVDD.n1646 0.00334
R17611 DVDD.n1650 DVDD.n1649 0.00334
R17612 DVDD.n1651 DVDD.n1650 0.00334
R17613 DVDD.n1652 DVDD.n1651 0.00334
R17614 DVDD.n1655 DVDD.n1652 0.00334
R17615 DVDD.n1656 DVDD.n1655 0.00334
R17616 DVDD.n1657 DVDD.n1656 0.00334
R17617 DVDD.n1658 DVDD.n1657 0.00334
R17618 DVDD.n1918 DVDD.n1658 0.00334
R17619 DVDD.n1919 DVDD.n1918 0.00334
R17620 DVDD.n1923 DVDD.n1919 0.00334
R17621 DVDD.n8080 DVDD.n1914 0.00334
R17622 DVDD.n8086 DVDD.n1914 0.00334
R17623 DVDD.n8087 DVDD.n8086 0.00334
R17624 DVDD.n8088 DVDD.n8087 0.00334
R17625 DVDD.n8088 DVDD.n1910 0.00334
R17626 DVDD.n8094 DVDD.n1910 0.00334
R17627 DVDD.n8095 DVDD.n8094 0.00334
R17628 DVDD.n8097 DVDD.n8095 0.00334
R17629 DVDD.n8097 DVDD.n8096 0.00334
R17630 DVDD.n8096 DVDD.n1906 0.00334
R17631 DVDD.n8104 DVDD.n1906 0.00334
R17632 DVDD.n8105 DVDD.n8104 0.00334
R17633 DVDD.n8106 DVDD.n8105 0.00334
R17634 DVDD.n8106 DVDD.n1851 0.00334
R17635 DVDD.n8123 DVDD.n1851 0.00334
R17636 DVDD.n8124 DVDD.n8123 0.00334
R17637 DVDD.n8125 DVDD.n8124 0.00334
R17638 DVDD.n8125 DVDD.n1847 0.00334
R17639 DVDD.n8131 DVDD.n1847 0.00334
R17640 DVDD.n8132 DVDD.n8131 0.00334
R17641 DVDD.n8133 DVDD.n8132 0.00334
R17642 DVDD.n8133 DVDD.n1843 0.00334
R17643 DVDD.n8139 DVDD.n1843 0.00334
R17644 DVDD.n8141 DVDD.n1840 0.00334
R17645 DVDD.n8156 DVDD.n1840 0.00334
R17646 DVDD.n8157 DVDD.n8156 0.00334
R17647 DVDD.n8159 DVDD.n8157 0.00334
R17648 DVDD.n8159 DVDD.n8158 0.00334
R17649 DVDD.n8158 DVDD.n1836 0.00334
R17650 DVDD.n8166 DVDD.n1836 0.00334
R17651 DVDD.n8167 DVDD.n8166 0.00334
R17652 DVDD.n8168 DVDD.n8167 0.00334
R17653 DVDD.n8169 DVDD.n8168 0.00334
R17654 DVDD.n7553 DVDD.n2506 0.00334
R17655 DVDD.n7554 DVDD.n7553 0.00334
R17656 DVDD.n7555 DVDD.n7554 0.00334
R17657 DVDD.n7555 DVDD.n2502 0.00334
R17658 DVDD.n7561 DVDD.n2502 0.00334
R17659 DVDD.n7562 DVDD.n7561 0.00334
R17660 DVDD.n7563 DVDD.n7562 0.00334
R17661 DVDD.n7563 DVDD.n2469 0.00334
R17662 DVDD.n7596 DVDD.n2469 0.00334
R17663 DVDD.n7599 DVDD.n7598 0.00334
R17664 DVDD.n7599 DVDD.n2463 0.00334
R17665 DVDD.n7605 DVDD.n2463 0.00334
R17666 DVDD.n7606 DVDD.n7605 0.00334
R17667 DVDD.n7607 DVDD.n7606 0.00334
R17668 DVDD.n7607 DVDD.n2459 0.00334
R17669 DVDD.n7613 DVDD.n2459 0.00334
R17670 DVDD.n7614 DVDD.n7613 0.00334
R17671 DVDD.n7615 DVDD.n7614 0.00334
R17672 DVDD.n7616 DVDD.n7615 0.00334
R17673 DVDD.n7617 DVDD.n7616 0.00334
R17674 DVDD.n7618 DVDD.n7617 0.00334
R17675 DVDD.n7619 DVDD.n7618 0.00334
R17676 DVDD.n7622 DVDD.n7619 0.00334
R17677 DVDD.n7623 DVDD.n7622 0.00334
R17678 DVDD.n7624 DVDD.n7623 0.00334
R17679 DVDD.n7625 DVDD.n7624 0.00334
R17680 DVDD.n7628 DVDD.n7625 0.00334
R17681 DVDD.n7629 DVDD.n7628 0.00334
R17682 DVDD.n7630 DVDD.n7629 0.00334
R17683 DVDD.n7631 DVDD.n7630 0.00334
R17684 DVDD.n7632 DVDD.n7631 0.00334
R17685 DVDD.n7633 DVDD.n7632 0.00334
R17686 DVDD.n2209 DVDD.n2208 0.00334
R17687 DVDD.n2253 DVDD.n2209 0.00334
R17688 DVDD.n2254 DVDD.n2253 0.00334
R17689 DVDD.n2255 DVDD.n2254 0.00334
R17690 DVDD.n2256 DVDD.n2255 0.00334
R17691 DVDD.n2257 DVDD.n2256 0.00334
R17692 DVDD.n2260 DVDD.n2257 0.00334
R17693 DVDD.n2261 DVDD.n2260 0.00334
R17694 DVDD.n2262 DVDD.n2261 0.00334
R17695 DVDD.n2263 DVDD.n2262 0.00334
R17696 DVDD.n2266 DVDD.n2263 0.00334
R17697 DVDD.n2267 DVDD.n2266 0.00334
R17698 DVDD.n2268 DVDD.n2267 0.00334
R17699 DVDD.n2269 DVDD.n2268 0.00334
R17700 DVDD.n2272 DVDD.n2269 0.00334
R17701 DVDD.n2273 DVDD.n2272 0.00334
R17702 DVDD.n2274 DVDD.n2273 0.00334
R17703 DVDD.n2275 DVDD.n2274 0.00334
R17704 DVDD.n2309 DVDD.n2275 0.00334
R17705 DVDD.n2311 DVDD.n2309 0.00334
R17706 DVDD.n2312 DVDD.n2311 0.00334
R17707 DVDD.n2313 DVDD.n2312 0.00334
R17708 DVDD.n2313 DVDD.n1925 0.00334
R17709 DVDD.n8077 DVDD.n1926 0.00334
R17710 DVDD.n1931 DVDD.n1926 0.00334
R17711 DVDD.n1932 DVDD.n1931 0.00334
R17712 DVDD.n1933 DVDD.n1932 0.00334
R17713 DVDD.n1936 DVDD.n1933 0.00334
R17714 DVDD.n1937 DVDD.n1936 0.00334
R17715 DVDD.n1938 DVDD.n1937 0.00334
R17716 DVDD.n1939 DVDD.n1938 0.00334
R17717 DVDD.n1942 DVDD.n1939 0.00334
R17718 DVDD.n1943 DVDD.n1942 0.00334
R17719 DVDD.n1944 DVDD.n1943 0.00334
R17720 DVDD.n1945 DVDD.n1944 0.00334
R17721 DVDD.n1990 DVDD.n1945 0.00334
R17722 DVDD.n1991 DVDD.n1990 0.00334
R17723 DVDD.n1992 DVDD.n1991 0.00334
R17724 DVDD.n1993 DVDD.n1992 0.00334
R17725 DVDD.n1994 DVDD.n1993 0.00334
R17726 DVDD.n1997 DVDD.n1994 0.00334
R17727 DVDD.n1998 DVDD.n1997 0.00334
R17728 DVDD.n1999 DVDD.n1998 0.00334
R17729 DVDD.n2000 DVDD.n1999 0.00334
R17730 DVDD.n2002 DVDD.n2000 0.00334
R17731 DVDD.n2003 DVDD.n2002 0.00334
R17732 DVDD.n2006 DVDD.n2005 0.00334
R17733 DVDD.n2007 DVDD.n2006 0.00334
R17734 DVDD.n2008 DVDD.n2007 0.00334
R17735 DVDD.n2011 DVDD.n2008 0.00334
R17736 DVDD.n2012 DVDD.n2011 0.00334
R17737 DVDD.n2013 DVDD.n2012 0.00334
R17738 DVDD.n2014 DVDD.n2013 0.00334
R17739 DVDD.n8000 DVDD.n2014 0.00334
R17740 DVDD.n8001 DVDD.n8000 0.00334
R17741 DVDD.n8002 DVDD.n8001 0.00334
R17742 DVDD.n2552 DVDD.n2551 0.00334
R17743 DVDD.n2553 DVDD.n2552 0.00334
R17744 DVDD.n2556 DVDD.n2553 0.00334
R17745 DVDD.n2557 DVDD.n2556 0.00334
R17746 DVDD.n2558 DVDD.n2557 0.00334
R17747 DVDD.n2559 DVDD.n2558 0.00334
R17748 DVDD.n2612 DVDD.n2559 0.00334
R17749 DVDD.n2613 DVDD.n2612 0.00334
R17750 DVDD.n2614 DVDD.n2613 0.00334
R17751 DVDD.n2619 DVDD.n2616 0.00334
R17752 DVDD.n2620 DVDD.n2619 0.00334
R17753 DVDD.n2621 DVDD.n2620 0.00334
R17754 DVDD.n2622 DVDD.n2621 0.00334
R17755 DVDD.n2625 DVDD.n2622 0.00334
R17756 DVDD.n2626 DVDD.n2625 0.00334
R17757 DVDD.n2627 DVDD.n2626 0.00334
R17758 DVDD.n2628 DVDD.n2627 0.00334
R17759 DVDD.n6942 DVDD.n2628 0.00334
R17760 DVDD.n6943 DVDD.n6942 0.00334
R17761 DVDD.n6944 DVDD.n6943 0.00334
R17762 DVDD.n6945 DVDD.n6944 0.00334
R17763 DVDD.n6946 DVDD.n6945 0.00334
R17764 DVDD.n6949 DVDD.n6946 0.00334
R17765 DVDD.n6950 DVDD.n6949 0.00334
R17766 DVDD.n6951 DVDD.n6950 0.00334
R17767 DVDD.n6952 DVDD.n6951 0.00334
R17768 DVDD.n6955 DVDD.n6952 0.00334
R17769 DVDD.n6956 DVDD.n6955 0.00334
R17770 DVDD.n6957 DVDD.n6956 0.00334
R17771 DVDD.n6958 DVDD.n6957 0.00334
R17772 DVDD.n6958 DVDD.n2201 0.00334
R17773 DVDD.n7789 DVDD.n2201 0.00334
R17774 DVDD.n7792 DVDD.n7791 0.00334
R17775 DVDD.n7792 DVDD.n2169 0.00334
R17776 DVDD.n7809 DVDD.n2169 0.00334
R17777 DVDD.n7810 DVDD.n7809 0.00334
R17778 DVDD.n7811 DVDD.n7810 0.00334
R17779 DVDD.n7811 DVDD.n2165 0.00334
R17780 DVDD.n7817 DVDD.n2165 0.00334
R17781 DVDD.n7818 DVDD.n7817 0.00334
R17782 DVDD.n7819 DVDD.n7818 0.00334
R17783 DVDD.n7819 DVDD.n2161 0.00334
R17784 DVDD.n7825 DVDD.n2161 0.00334
R17785 DVDD.n7826 DVDD.n7825 0.00334
R17786 DVDD.n7827 DVDD.n7826 0.00334
R17787 DVDD.n7827 DVDD.n2157 0.00334
R17788 DVDD.n7833 DVDD.n2157 0.00334
R17789 DVDD.n7834 DVDD.n7833 0.00334
R17790 DVDD.n7835 DVDD.n7834 0.00334
R17791 DVDD.n7835 DVDD.n2153 0.00334
R17792 DVDD.n7845 DVDD.n2153 0.00334
R17793 DVDD.n7846 DVDD.n7845 0.00334
R17794 DVDD.n7848 DVDD.n7846 0.00334
R17795 DVDD.n7848 DVDD.n7847 0.00334
R17796 DVDD.n7847 DVDD.n2119 0.00334
R17797 DVDD.n7857 DVDD.n2114 0.00334
R17798 DVDD.n7863 DVDD.n2114 0.00334
R17799 DVDD.n7864 DVDD.n7863 0.00334
R17800 DVDD.n7865 DVDD.n7864 0.00334
R17801 DVDD.n7865 DVDD.n2110 0.00334
R17802 DVDD.n7871 DVDD.n2110 0.00334
R17803 DVDD.n7872 DVDD.n7871 0.00334
R17804 DVDD.n7874 DVDD.n7872 0.00334
R17805 DVDD.n7874 DVDD.n7873 0.00334
R17806 DVDD.n7873 DVDD.n2106 0.00334
R17807 DVDD.n7881 DVDD.n2106 0.00334
R17808 DVDD.n7882 DVDD.n7881 0.00334
R17809 DVDD.n7883 DVDD.n7882 0.00334
R17810 DVDD.n7883 DVDD.n2072 0.00334
R17811 DVDD.n7896 DVDD.n2072 0.00334
R17812 DVDD.n7897 DVDD.n7896 0.00334
R17813 DVDD.n7898 DVDD.n7897 0.00334
R17814 DVDD.n7898 DVDD.n2068 0.00334
R17815 DVDD.n7904 DVDD.n2068 0.00334
R17816 DVDD.n7905 DVDD.n7904 0.00334
R17817 DVDD.n7906 DVDD.n7905 0.00334
R17818 DVDD.n7906 DVDD.n2064 0.00334
R17819 DVDD.n7912 DVDD.n2064 0.00334
R17820 DVDD.n7914 DVDD.n2062 0.00334
R17821 DVDD.n7931 DVDD.n2062 0.00334
R17822 DVDD.n7932 DVDD.n7931 0.00334
R17823 DVDD.n7934 DVDD.n7932 0.00334
R17824 DVDD.n7934 DVDD.n7933 0.00334
R17825 DVDD.n7933 DVDD.n2058 0.00334
R17826 DVDD.n7941 DVDD.n2058 0.00334
R17827 DVDD.n7942 DVDD.n7941 0.00334
R17828 DVDD.n7943 DVDD.n7942 0.00334
R17829 DVDD.n7944 DVDD.n7943 0.00334
R17830 DVDD.n7945 DVDD.n7944 0.00334
R17831 DVDD.n5509 DVDD.n5508 0.00334
R17832 DVDD.n5510 DVDD.n5509 0.00334
R17833 DVDD.n5513 DVDD.n5510 0.00334
R17834 DVDD.n5514 DVDD.n5513 0.00334
R17835 DVDD.n5515 DVDD.n5514 0.00334
R17836 DVDD.n5517 DVDD.n5515 0.00334
R17837 DVDD.n5517 DVDD.n5516 0.00334
R17838 DVDD.n5516 DVDD.n3062 0.00334
R17839 DVDD.n6749 DVDD.n3062 0.00334
R17840 DVDD.n6747 DVDD.n3063 0.00334
R17841 DVDD.n3066 DVDD.n3063 0.00334
R17842 DVDD.n3067 DVDD.n3066 0.00334
R17843 DVDD.n3068 DVDD.n3067 0.00334
R17844 DVDD.n3071 DVDD.n3068 0.00334
R17845 DVDD.n3072 DVDD.n3071 0.00334
R17846 DVDD.n3073 DVDD.n3072 0.00334
R17847 DVDD.n3074 DVDD.n3073 0.00334
R17848 DVDD.n3075 DVDD.n3074 0.00334
R17849 DVDD.n3076 DVDD.n3075 0.00334
R17850 DVDD.n3077 DVDD.n3076 0.00334
R17851 DVDD.n3078 DVDD.n3077 0.00334
R17852 DVDD.n3079 DVDD.n3078 0.00334
R17853 DVDD.n3082 DVDD.n3079 0.00334
R17854 DVDD.n3083 DVDD.n3082 0.00334
R17855 DVDD.n3084 DVDD.n3083 0.00334
R17856 DVDD.n3085 DVDD.n3084 0.00334
R17857 DVDD.n3088 DVDD.n3085 0.00334
R17858 DVDD.n3089 DVDD.n3088 0.00334
R17859 DVDD.n3090 DVDD.n3089 0.00334
R17860 DVDD.n3091 DVDD.n3090 0.00334
R17861 DVDD.n3093 DVDD.n3091 0.00334
R17862 DVDD.n3094 DVDD.n3093 0.00334
R17863 DVDD.n3188 DVDD.n3095 0.00334
R17864 DVDD.n3191 DVDD.n3188 0.00334
R17865 DVDD.n3192 DVDD.n3191 0.00334
R17866 DVDD.n3193 DVDD.n3192 0.00334
R17867 DVDD.n3194 DVDD.n3193 0.00334
R17868 DVDD.n3195 DVDD.n3194 0.00334
R17869 DVDD.n3198 DVDD.n3195 0.00334
R17870 DVDD.n3199 DVDD.n3198 0.00334
R17871 DVDD.n3200 DVDD.n3199 0.00334
R17872 DVDD.n3201 DVDD.n3200 0.00334
R17873 DVDD.n3204 DVDD.n3201 0.00334
R17874 DVDD.n3205 DVDD.n3204 0.00334
R17875 DVDD.n3206 DVDD.n3205 0.00334
R17876 DVDD.n3207 DVDD.n3206 0.00334
R17877 DVDD.n3210 DVDD.n3207 0.00334
R17878 DVDD.n3211 DVDD.n3210 0.00334
R17879 DVDD.n3212 DVDD.n3211 0.00334
R17880 DVDD.n3213 DVDD.n3212 0.00334
R17881 DVDD.n3308 DVDD.n3213 0.00334
R17882 DVDD.n3310 DVDD.n3308 0.00334
R17883 DVDD.n3311 DVDD.n3310 0.00334
R17884 DVDD.n3312 DVDD.n3311 0.00334
R17885 DVDD.n3313 DVDD.n3312 0.00334
R17886 DVDD.n3317 DVDD.n3316 0.00334
R17887 DVDD.n3318 DVDD.n3317 0.00334
R17888 DVDD.n3321 DVDD.n3318 0.00334
R17889 DVDD.n3322 DVDD.n3321 0.00334
R17890 DVDD.n3323 DVDD.n3322 0.00334
R17891 DVDD.n3324 DVDD.n3323 0.00334
R17892 DVDD.n3327 DVDD.n3324 0.00334
R17893 DVDD.n3328 DVDD.n3327 0.00334
R17894 DVDD.n3329 DVDD.n3328 0.00334
R17895 DVDD.n3330 DVDD.n3329 0.00334
R17896 DVDD.n3366 DVDD.n3330 0.00334
R17897 DVDD.n3367 DVDD.n3366 0.00334
R17898 DVDD.n3371 DVDD.n3367 0.00334
R17899 DVDD.n3372 DVDD.n3371 0.00334
R17900 DVDD.n3373 DVDD.n3372 0.00334
R17901 DVDD.n3374 DVDD.n3373 0.00334
R17902 DVDD.n3375 DVDD.n3374 0.00334
R17903 DVDD.n3378 DVDD.n3375 0.00334
R17904 DVDD.n3379 DVDD.n3378 0.00334
R17905 DVDD.n3380 DVDD.n3379 0.00334
R17906 DVDD.n3381 DVDD.n3380 0.00334
R17907 DVDD.n3383 DVDD.n3381 0.00334
R17908 DVDD.n3384 DVDD.n3383 0.00334
R17909 DVDD.n3386 DVDD.n3385 0.00334
R17910 DVDD.n3387 DVDD.n3386 0.00334
R17911 DVDD.n3388 DVDD.n3387 0.00334
R17912 DVDD.n3391 DVDD.n3388 0.00334
R17913 DVDD.n3392 DVDD.n3391 0.00334
R17914 DVDD.n3393 DVDD.n3392 0.00334
R17915 DVDD.n3394 DVDD.n3393 0.00334
R17916 DVDD.n6595 DVDD.n3394 0.00334
R17917 DVDD.n6596 DVDD.n6595 0.00334
R17918 DVDD.n6597 DVDD.n6596 0.00334
R17919 DVDD.n5379 DVDD.n5378 0.00334
R17920 DVDD.n5380 DVDD.n5379 0.00334
R17921 DVDD.n5383 DVDD.n5380 0.00334
R17922 DVDD.n5384 DVDD.n5383 0.00334
R17923 DVDD.n5385 DVDD.n5384 0.00334
R17924 DVDD.n5386 DVDD.n5385 0.00334
R17925 DVDD.n5387 DVDD.n5386 0.00334
R17926 DVDD.n5389 DVDD.n5387 0.00334
R17927 DVDD.n5389 DVDD.n5388 0.00334
R17928 DVDD.n5713 DVDD.n5712 0.00334
R17929 DVDD.n5714 DVDD.n5713 0.00334
R17930 DVDD.n5714 DVDD.n4444 0.00334
R17931 DVDD.n5720 DVDD.n4444 0.00334
R17932 DVDD.n5721 DVDD.n5720 0.00334
R17933 DVDD.n5722 DVDD.n5721 0.00334
R17934 DVDD.n5722 DVDD.n4440 0.00334
R17935 DVDD.n5728 DVDD.n4440 0.00334
R17936 DVDD.n5729 DVDD.n5728 0.00334
R17937 DVDD.n5730 DVDD.n5729 0.00334
R17938 DVDD.n5730 DVDD.n4437 0.00334
R17939 DVDD.n5735 DVDD.n4437 0.00334
R17940 DVDD.n5736 DVDD.n5735 0.00334
R17941 DVDD.n5737 DVDD.n5736 0.00334
R17942 DVDD.n5737 DVDD.n4433 0.00334
R17943 DVDD.n5743 DVDD.n4433 0.00334
R17944 DVDD.n5744 DVDD.n5743 0.00334
R17945 DVDD.n5745 DVDD.n5744 0.00334
R17946 DVDD.n5745 DVDD.n4429 0.00334
R17947 DVDD.n5752 DVDD.n4429 0.00334
R17948 DVDD.n5753 DVDD.n5752 0.00334
R17949 DVDD.n5754 DVDD.n5753 0.00334
R17950 DVDD.n5754 DVDD.n4391 0.00334
R17951 DVDD.n6103 DVDD.n6102 0.00334
R17952 DVDD.n6103 DVDD.n4303 0.00334
R17953 DVDD.n6116 DVDD.n4303 0.00334
R17954 DVDD.n6117 DVDD.n6116 0.00334
R17955 DVDD.n6118 DVDD.n6117 0.00334
R17956 DVDD.n6118 DVDD.n4299 0.00334
R17957 DVDD.n6124 DVDD.n4299 0.00334
R17958 DVDD.n6125 DVDD.n6124 0.00334
R17959 DVDD.n6126 DVDD.n6125 0.00334
R17960 DVDD.n6126 DVDD.n4295 0.00334
R17961 DVDD.n6132 DVDD.n4295 0.00334
R17962 DVDD.n6133 DVDD.n6132 0.00334
R17963 DVDD.n6134 DVDD.n6133 0.00334
R17964 DVDD.n6134 DVDD.n4291 0.00334
R17965 DVDD.n6140 DVDD.n4291 0.00334
R17966 DVDD.n6141 DVDD.n6140 0.00334
R17967 DVDD.n6142 DVDD.n6141 0.00334
R17968 DVDD.n6142 DVDD.n4287 0.00334
R17969 DVDD.n6148 DVDD.n4287 0.00334
R17970 DVDD.n6149 DVDD.n6148 0.00334
R17971 DVDD.n6150 DVDD.n6149 0.00334
R17972 DVDD.n6150 DVDD.n3944 0.00334
R17973 DVDD.n6158 DVDD.n3944 0.00334
R17974 DVDD.n6160 DVDD.n3910 0.00334
R17975 DVDD.n6166 DVDD.n3910 0.00334
R17976 DVDD.n6167 DVDD.n6166 0.00334
R17977 DVDD.n6168 DVDD.n6167 0.00334
R17978 DVDD.n6168 DVDD.n3906 0.00334
R17979 DVDD.n6174 DVDD.n3906 0.00334
R17980 DVDD.n6175 DVDD.n6174 0.00334
R17981 DVDD.n6176 DVDD.n6175 0.00334
R17982 DVDD.n6176 DVDD.n3902 0.00334
R17983 DVDD.n6183 DVDD.n3902 0.00334
R17984 DVDD.n6184 DVDD.n6183 0.00334
R17985 DVDD.n6185 DVDD.n6184 0.00334
R17986 DVDD.n6185 DVDD.n3900 0.00334
R17987 DVDD.n6191 DVDD.n3900 0.00334
R17988 DVDD.n6192 DVDD.n6191 0.00334
R17989 DVDD.n6193 DVDD.n6192 0.00334
R17990 DVDD.n6193 DVDD.n3897 0.00334
R17991 DVDD.n6199 DVDD.n3897 0.00334
R17992 DVDD.n6200 DVDD.n6199 0.00334
R17993 DVDD.n6201 DVDD.n6200 0.00334
R17994 DVDD.n6201 DVDD.n3893 0.00334
R17995 DVDD.n6208 DVDD.n3893 0.00334
R17996 DVDD.n6209 DVDD.n6208 0.00334
R17997 DVDD.n3512 DVDD.n3511 0.00334
R17998 DVDD.n3513 DVDD.n3512 0.00334
R17999 DVDD.n3514 DVDD.n3513 0.00334
R18000 DVDD.n3517 DVDD.n3514 0.00334
R18001 DVDD.n3518 DVDD.n3517 0.00334
R18002 DVDD.n3519 DVDD.n3518 0.00334
R18003 DVDD.n3520 DVDD.n3519 0.00334
R18004 DVDD.n6389 DVDD.n3520 0.00334
R18005 DVDD.n6390 DVDD.n6389 0.00334
R18006 DVDD.n6391 DVDD.n6390 0.00334
R18007 DVDD.n416 DVDD.n291 0.00334
R18008 DVDD.n418 DVDD.n416 0.00334
R18009 DVDD.n425 DVDD.n310 0.00334
R18010 DVDD.n311 DVDD.n310 0.00334
R18011 DVDD.n324 DVDD.n311 0.00334
R18012 DVDD.n325 DVDD.n324 0.00334
R18013 DVDD.n327 DVDD.n326 0.00334
R18014 DVDD.n9426 DVDD.n327 0.00334
R18015 DVDD.n9427 DVDD.n9426 0.00334
R18016 DVDD.n9427 DVDD.n196 0.00334
R18017 DVDD.n279 DVDD.n195 0.00334
R18018 DVDD.n9486 DVDD.n279 0.00334
R18019 DVDD.n9487 DVDD.n9486 0.00334
R18020 DVDD.n9488 DVDD.n9487 0.00334
R18021 DVDD.n9499 DVDD.n270 0.00334
R18022 DVDD.n9500 DVDD.n9499 0.00334
R18023 DVDD.n9501 DVDD.n9500 0.00334
R18024 DVDD.n9501 DVDD.n239 0.00334
R18025 DVDD.n9560 DVDD.n9559 0.00334
R18026 DVDD.n9559 DVDD.n240 0.00334
R18027 DVDD.n9321 DVDD.n426 0.00334
R18028 DVDD.n9325 DVDD.n426 0.00334
R18029 DVDD.n9347 DVDD.n9326 0.00334
R18030 DVDD.n9343 DVDD.n9326 0.00334
R18031 DVDD.n9343 DVDD.n9342 0.00334
R18032 DVDD.n9342 DVDD.n9341 0.00334
R18033 DVDD.n9337 DVDD.n9331 0.00334
R18034 DVDD.n9337 DVDD.n9336 0.00334
R18035 DVDD.n9336 DVDD.n9335 0.00334
R18036 DVDD.n9335 DVDD.n198 0.00334
R18037 DVDD.n9578 DVDD.n199 0.00334
R18038 DVDD.n9574 DVDD.n199 0.00334
R18039 DVDD.n9574 DVDD.n9573 0.00334
R18040 DVDD.n9573 DVDD.n9572 0.00334
R18041 DVDD.n9568 DVDD.n205 0.00334
R18042 DVDD.n9568 DVDD.n9567 0.00334
R18043 DVDD.n9567 DVDD.n9566 0.00334
R18044 DVDD.n9566 DVDD.n210 0.00334
R18045 DVDD.n5298 DVDD.n237 0.00334
R18046 DVDD.n5299 DVDD.n5298 0.00334
R18047 DVDD.n4107 DVDD.n4106 0.00334
R18048 DVDD.n4106 DVDD.n424 0.00334
R18049 DVDD.n4092 DVDD.n423 0.00334
R18050 DVDD.n4092 DVDD.n4091 0.00334
R18051 DVDD.n4091 DVDD.n4090 0.00334
R18052 DVDD.n4090 DVDD.n4020 0.00334
R18053 DVDD.n4086 DVDD.n4085 0.00334
R18054 DVDD.n4085 DVDD.n4084 0.00334
R18055 DVDD.n4084 DVDD.n4025 0.00334
R18056 DVDD.n4025 DVDD.n186 0.00334
R18057 DVDD.n3988 DVDD.n185 0.00334
R18058 DVDD.n4126 DVDD.n3988 0.00334
R18059 DVDD.n4127 DVDD.n4126 0.00334
R18060 DVDD.n4128 DVDD.n4127 0.00334
R18061 DVDD.n4139 DVDD.n3979 0.00334
R18062 DVDD.n4140 DVDD.n4139 0.00334
R18063 DVDD.n4141 DVDD.n4140 0.00334
R18064 DVDD.n4141 DVDD.n235 0.00334
R18065 DVDD.n4212 DVDD.n234 0.00334
R18066 DVDD.n4212 DVDD.n4211 0.00334
R18067 DVDD.n8786 DVDD.n8782 0.00334
R18068 DVDD.n8782 DVDD.n420 0.00334
R18069 DVDD.n961 DVDD.n419 0.00334
R18070 DVDD.n962 DVDD.n961 0.00334
R18071 DVDD.n962 DVDD.n958 0.00334
R18072 DVDD.n967 DVDD.n958 0.00334
R18073 DVDD.n969 DVDD.n968 0.00334
R18074 DVDD.n970 DVDD.n969 0.00334
R18075 DVDD.n971 DVDD.n970 0.00334
R18076 DVDD.n971 DVDD.n190 0.00334
R18077 DVDD.n1020 DVDD.n191 0.00334
R18078 DVDD.n1021 DVDD.n1020 0.00334
R18079 DVDD.n1022 DVDD.n1021 0.00334
R18080 DVDD.n1022 DVDD.n1016 0.00334
R18081 DVDD.n1027 DVDD.n1026 0.00334
R18082 DVDD.n1028 DVDD.n1027 0.00334
R18083 DVDD.n1029 DVDD.n1028 0.00334
R18084 DVDD.n1029 DVDD.n232 0.00334
R18085 DVDD.n3586 DVDD.n231 0.00334
R18086 DVDD.n3587 DVDD.n3586 0.00334
R18087 DVDD.n6746 DVDD.n2615 0.00332
R18088 DVDD.n7000 DVDD.n6999 0.00332
R18089 DVDD.n2471 DVDD.n2466 0.00332
R18090 DVDD.n7268 DVDD.n7267 0.00332
R18091 DVDD.n5711 DVDD.n5709 0.00332
R18092 DVDD.n7222 DVDD.n7043 0.00329
R18093 DVDD.n7281 DVDD.n7120 0.00329
R18094 DVDD.n8356 DVDD.n1544 0.00329
R18095 DVDD.n1628 DVDD.n1600 0.00329
R18096 DVDD.n7545 DVDD.n7523 0.00329
R18097 DVDD.n7587 DVDD.n7565 0.00329
R18098 DVDD.n7656 DVDD.n2374 0.00329
R18099 DVDD.n7781 DVDD.n7780 0.00329
R18100 DVDD.n7020 DVDD.n2536 0.00329
R18101 DVDD.n2609 DVDD.n2573 0.00329
R18102 DVDD.n6934 DVDD.n2638 0.00329
R18103 DVDD.n7799 DVDD.n7794 0.00329
R18104 DVDD.n5530 DVDD.n5492 0.00329
R18105 DVDD.n6765 DVDD.n3038 0.00329
R18106 DVDD.n6731 DVDD.n2659 0.00329
R18107 DVDD.n3184 DVDD.n3109 0.00329
R18108 DVDD.n5416 DVDD.n4470 0.00329
R18109 DVDD.n5400 DVDD.n2975 0.00329
R18110 DVDD.n4438 DVDD.n2807 0.00329
R18111 DVDD.n6111 DVDD.n6105 0.00329
R18112 DVDD.n9361 DVDD.n409 0.00329
R18113 DVDD.n9398 DVDD.n202 0.00329
R18114 DVDD.n5287 DVDD.n211 0.00329
R18115 DVDD.n4103 DVDD.n4102 0.00329
R18116 DVDD.n4072 DVDD.n4071 0.00329
R18117 DVDD.n4145 DVDD.n4143 0.00329
R18118 DVDD.n296 DVDD.n294 0.00329
R18119 DVDD.n363 DVDD.n362 0.00329
R18120 DVDD.n9505 DVDD.n9503 0.00329
R18121 DVDD.n8772 DVDD.n89 0.00329
R18122 DVDD.n8718 DVDD.n891 0.00329
R18123 DVDD.n8686 DVDD.n1011 0.00329
R18124 DVDD.n5899 DVDD.n5891 0.00325625
R18125 DVDD.n5483 DVDD.n5482 0.00325625
R18126 DVDD.n4450 DVDD.n3022 0.00325625
R18127 DVDD.n6080 DVDD.n5910 0.0032
R18128 DVDD.n6079 DVDD.n5912 0.0032
R18129 DVDD.n5709 DVDD.n5679 0.0032
R18130 DVDD.n5678 DVDD.n5677 0.0032
R18131 DVDD.n1660 DVDD.n1654 0.00317
R18132 DVDD.n8290 DVDD.n1688 0.00317
R18133 DVDD.n8118 DVDD.n1892 0.00317
R18134 DVDD.n1891 DVDD.n1853 0.00317
R18135 DVDD.n8154 DVDD.n1236 0.00317
R18136 DVDD.n8191 DVDD.n1801 0.00317
R18137 DVDD.n8173 DVDD.n1800 0.00317
R18138 DVDD.n7750 DVDD.n7749 0.00317
R18139 DVDD.n2295 DVDD.n2292 0.00317
R18140 DVDD.n1947 DVDD.n1941 0.00317
R18141 DVDD.n8054 DVDD.n1973 0.00317
R18142 DVDD.n8019 DVDD.n1197 0.00317
R18143 DVDD.n8011 DVDD.n8010 0.00317
R18144 DVDD.n8008 DVDD.n8007 0.00317
R18145 DVDD.n7843 DVDD.n7842 0.00317
R18146 DVDD.n2149 DVDD.n2120 0.00317
R18147 DVDD.n7890 DVDD.n2097 0.00317
R18148 DVDD.n2096 DVDD.n2074 0.00317
R18149 DVDD.n7929 DVDD.n1158 0.00317
R18150 DVDD.n7958 DVDD.n2030 0.00317
R18151 DVDD.n7948 DVDD.n2029 0.00317
R18152 DVDD.n6677 DVDD.n6676 0.00317
R18153 DVDD.n6674 DVDD.n6673 0.00317
R18154 DVDD.n6651 DVDD.n6650 0.00317
R18155 DVDD.n3363 DVDD.n3357 0.00317
R18156 DVDD.n6614 DVDD.n1119 0.00317
R18157 DVDD.n6606 DVDD.n6605 0.00317
R18158 DVDD.n6603 DVDD.n6602 0.00317
R18159 DVDD.n6146 DVDD.n4282 0.00317
R18160 DVDD.n4285 DVDD.n3946 0.00317
R18161 DVDD.n6180 DVDD.n3557 0.00317
R18162 DVDD.n3561 DVDD.n3558 0.00317
R18163 DVDD.n6408 DVDD.n1057 0.00317
R18164 DVDD.n6400 DVDD.n6399 0.00317
R18165 DVDD.n6397 DVDD.n6396 0.00317
R18166 DVDD.n5289 DVDD.n5288 0.00315748
R18167 DVDD.n5291 DVDD.n5290 0.00315748
R18168 DVDD.n5293 DVDD.n2895 0.00315748
R18169 DVDD.n5296 DVDD.n2899 0.00315748
R18170 DVDD.n5305 DVDD.n5304 0.00315748
R18171 DVDD.n5307 DVDD.n5306 0.00315748
R18172 DVDD.n5309 DVDD.n2958 0.00315748
R18173 DVDD.n704 DVDD.n583 0.00315748
R18174 DVDD.n843 DVDD.n842 0.00315748
R18175 DVDD.n8707 DVDD.n904 0.00315748
R18176 DVDD.n3825 DVDD.n3810 0.00315748
R18177 DVDD.n9007 DVDD.n557 0.00315748
R18178 DVDD.n4010 DVDD.n4008 0.00315748
R18179 DVDD.n4132 DVDD.n3984 0.00315748
R18180 DVDD.n6044 DVDD.n3950 0.00315748
R18181 DVDD.n5013 DVDD.n4866 0.00315748
R18182 DVDD.n303 DVDD.n302 0.00315748
R18183 DVDD.n9492 DVDD.n275 0.00315748
R18184 DVDD.n5811 DVDD.n4379 0.00315748
R18185 DVDD.n5151 DVDD.n4579 0.00315748
R18186 DVDD.n9312 DVDD.n443 0.00315748
R18187 DVDD.n9409 DVDD.n9408 0.00315748
R18188 DVDD.n2871 DVDD.n2811 0.00315748
R18189 DVDD.n9693 DVDD.n3 0.00313571
R18190 DVDD.n742 DVDD.n647 0.00311161
R18191 DVDD.n740 DVDD.n650 0.00311161
R18192 DVDD.n738 DVDD.n646 0.00311161
R18193 DVDD.n736 DVDD.n651 0.00311161
R18194 DVDD.n734 DVDD.n645 0.00311161
R18195 DVDD.n732 DVDD.n652 0.00311161
R18196 DVDD.n730 DVDD.n644 0.00311161
R18197 DVDD.n728 DVDD.n653 0.00311161
R18198 DVDD.n726 DVDD.n643 0.00311161
R18199 DVDD.n8893 DVDD.n654 0.00311161
R18200 DVDD.n5301 DVDD.n2957 0.00309529
R18201 DVDD.n9320 DVDD.n427 0.00309529
R18202 DVDD.n254 DVDD.n253 0.00309529
R18203 DVDD.n9469 DVDD.n289 0.00309529
R18204 DVDD.n3589 DVDD.n3588 0.00309529
R18205 DVDD.n8787 DVDD.n8781 0.00309529
R18206 DVDD.n4210 DVDD.n4209 0.00309529
R18207 DVDD.n4109 DVDD.n3998 0.00309529
R18208 DVDD.n7208 DVDD.n7029 0.00305
R18209 DVDD.n7266 DVDD.n7106 0.00305
R18210 DVDD.n8343 DVDD.n1529 0.00305
R18211 DVDD.n8317 DVDD.n1619 0.00305
R18212 DVDD.n7550 DVDD.n2504 0.00305
R18213 DVDD.n7592 DVDD.n2465 0.00305
R18214 DVDD.n7679 DVDD.n2388 0.00305
R18215 DVDD.n7776 DVDD.n7773 0.00305
R18216 DVDD.n7012 DVDD.n2521 0.00305
R18217 DVDD.n6998 DVDD.n2597 0.00305
R18218 DVDD.n6982 DVDD.n6939 0.00305
R18219 DVDD.n7806 DVDD.n2167 0.00305
R18220 DVDD.n5523 DVDD.n5493 0.00305
R18221 DVDD.n6745 DVDD.n3024 0.00305
R18222 DVDD.n6924 DVDD.n2672 0.00305
R18223 DVDD.n6704 DVDD.n6700 0.00305
R18224 DVDD.n5409 DVDD.n4471 0.00305
R18225 DVDD.n5710 DVDD.n2961 0.00305
R18226 DVDD.n6856 DVDD.n2820 0.00305
R18227 DVDD.n6113 DVDD.n4301 0.00305
R18228 DVDD.n9613 DVDD.n129 0.00305
R18229 DVDD.n9391 DVDD.n170 0.00305
R18230 DVDD.n6791 DVDD.n2894 0.00305
R18231 DVDD.n4095 DVDD.n4094 0.00305
R18232 DVDD.n4080 DVDD.n4079 0.00305
R18233 DVDD.n4215 DVDD.n4214 0.00305
R18234 DVDD.n9457 DVDD.n9456 0.00305
R18235 DVDD.n9431 DVDD.n347 0.00305
R18236 DVDD.n9557 DVDD.n243 0.00305
R18237 DVDD.n8765 DVDD.n850 0.00305
R18238 DVDD.n8735 DVDD.n883 0.00305
R18239 DVDD.n8682 DVDD.n1038 0.00305
R18240 DVDD DVDD.n1799 0.00287
R18241 DVDD DVDD.n7985 0.00287
R18242 DVDD DVDD.n2028 0.00287
R18243 DVDD DVDD.n6485 0.00287
R18244 DVDD DVDD.n3551 0.00287
R18245 DVDD.n8141 DVDD.n8140 0.00286
R18246 DVDD.n2005 DVDD.n1842 0.00286
R18247 DVDD.n7914 DVDD.n7913 0.00286
R18248 DVDD.n3385 DVDD.n2063 0.00286
R18249 DVDD.n6210 DVDD.n3511 0.00286
R18250 DVDD.n4627 DVDD.n4623 0.00280315
R18251 DVDD.n4629 DVDD.n4615 0.00280315
R18252 DVDD.n4631 DVDD.n4622 0.00280315
R18253 DVDD.n4633 DVDD.n4616 0.00280315
R18254 DVDD.n4635 DVDD.n4621 0.00280315
R18255 DVDD.n4637 DVDD.n4617 0.00280315
R18256 DVDD.n4639 DVDD.n4620 0.00280315
R18257 DVDD.n4641 DVDD.n4618 0.00280315
R18258 DVDD.n4643 DVDD.n4619 0.00280315
R18259 DVDD.n4712 DVDD.n4624 0.00280315
R18260 DVDD.n8761 DVDD.n855 0.00280315
R18261 DVDD.n6263 DVDD.n3341 0.00280315
R18262 DVDD.n4037 DVDD.n4036 0.00280315
R18263 DVDD.n5954 DVDD.n3219 0.00280315
R18264 DVDD.n317 DVDD.n316 0.00280315
R18265 DVDD.n5852 DVDD.n3106 0.00280315
R18266 DVDD.n9608 DVDD.n133 0.00280315
R18267 DVDD.n6914 DVDD.n2735 0.00280315
R18268 DVDD DVDD.n8169 0.00278
R18269 DVDD DVDD.n8002 0.00278
R18270 DVDD DVDD.n6597 0.00278
R18271 DVDD DVDD.n6391 0.00278
R18272 DVDD.n7223 DVDD.n7030 0.00275
R18273 DVDD.n7272 DVDD.n7107 0.00275
R18274 DVDD.n8348 DVDD.n1530 0.00275
R18275 DVDD.n8321 DVDD.n1629 0.00275
R18276 DVDD.n7534 DVDD.n2508 0.00275
R18277 DVDD.n7576 DVDD.n2472 0.00275
R18278 DVDD.n7653 DVDD.n2372 0.00275
R18279 DVDD.n7778 DVDD.n2217 0.00275
R18280 DVDD.n7017 DVDD.n2522 0.00275
R18281 DVDD.n7003 DVDD.n2610 0.00275
R18282 DVDD.n6979 DVDD.n6976 0.00275
R18283 DVDD.n7798 DVDD.n2171 0.00275
R18284 DVDD.n5527 DVDD.n5495 0.00275
R18285 DVDD.n6754 DVDD.n3025 0.00275
R18286 DVDD.n6729 DVDD.n2656 0.00275
R18287 DVDD.n3189 DVDD.n3122 0.00275
R18288 DVDD.n4404 DVDD.n2785 0.00275
R18289 DVDD.n5759 DVDD.n4426 0.00275
R18290 DVDD.n4405 DVDD.n2786 0.00275
R18291 DVDD.n4425 DVDD.n4394 0.00275
R18292 DVDD.n5413 DVDD.n4472 0.00275
R18293 DVDD.n5401 DVDD.n2962 0.00275
R18294 DVDD.n5731 DVDD.n2804 0.00275
R18295 DVDD.n6106 DVDD.n4305 0.00275
R18296 DVDD.n9616 DVDD.n106 0.00275
R18297 DVDD.n9425 DVDD.n201 0.00275
R18298 DVDD.n228 DVDD.n212 0.00275
R18299 DVDD.n9324 DVDD.n103 0.00275
R18300 DVDD.n9577 DVDD.n200 0.00275
R18301 DVDD.n9564 DVDD.n9563 0.00275
R18302 DVDD.n417 DVDD.n103 0.00275
R18303 DVDD.n360 DVDD.n200 0.00275
R18304 DVDD.n9563 DVDD.n221 0.00275
R18305 DVDD.n9616 DVDD.n121 0.00275
R18306 DVDD.n9425 DVDD.n371 0.00275
R18307 DVDD.n4144 DVDD.n228 0.00275
R18308 DVDD.n9616 DVDD.n123 0.00275
R18309 DVDD.n9425 DVDD.n361 0.00275
R18310 DVDD.n9504 DVDD.n228 0.00275
R18311 DVDD.n8783 DVDD.n103 0.00275
R18312 DVDD.n1018 DVDD.n200 0.00275
R18313 DVDD.n9563 DVDD.n216 0.00275
R18314 DVDD.n4104 DVDD.n103 0.00275
R18315 DVDD.n3989 DVDD.n200 0.00275
R18316 DVDD.n9563 DVDD.n219 0.00275
R18317 DVDD.n1724 DVDD.n1703 0.00275
R18318 DVDD.n8249 DVDD.n1763 0.00275
R18319 DVDD.n8224 DVDD.n1272 0.00275
R18320 DVDD.n8205 DVDD.n1797 0.00275
R18321 DVDD.n9616 DVDD.n117 0.00275
R18322 DVDD.n9425 DVDD.n349 0.00275
R18323 DVDD.n1012 DVDD.n228 0.00275
R18324 DVDD.n8965 DVDD.n548 0.00275
R18325 DVDD.n8936 DVDD.n592 0.00275
R18326 DVDD.n8910 DVDD.n617 0.00275
R18327 DVDD.n8892 DVDD.n648 0.00275
R18328 DVDD.n9172 DVDD.n533 0.00275
R18329 DVDD.n65 DVDD.n55 0.00275
R18330 DVDD.n30 DVDD.n20 0.00275
R18331 DVDD.n8080 DVDD.n8079 0.0027
R18332 DVDD.n8078 DVDD.n8077 0.0027
R18333 DVDD.n7857 DVDD.n1924 0.0027
R18334 DVDD.n3316 DVDD.n3315 0.0027
R18335 DVDD.n6160 DVDD.n6159 0.0027
R18336 DVDD.n9561 DVDD 0.00267716
R18337 DVDD.n9354 DVDD 0.00267716
R18338 DVDD.n8293 DVDD.n8292 0.00263
R18339 DVDD.n8292 DVDD.n1665 0.00263
R18340 DVDD.n8115 DVDD.n1899 0.00263
R18341 DVDD.n8115 DVDD.n8108 0.00263
R18342 DVDD.n8151 DVDD.n1249 0.00263
R18343 DVDD.n8152 DVDD.n8151 0.00263
R18344 DVDD.n8187 DVDD.n1814 0.00263
R18345 DVDD.n8187 DVDD.n8176 0.00263
R18346 DVDD.n2294 DVDD.n2285 0.00263
R18347 DVDD.n2307 DVDD.n2294 0.00263
R18348 DVDD.n8057 DVDD.n8056 0.00263
R18349 DVDD.n8056 DVDD.n1954 0.00263
R18350 DVDD.n8031 DVDD.n1210 0.00263
R18351 DVDD.n8032 DVDD.n8031 0.00263
R18352 DVDD.n7997 DVDD.n7961 0.00263
R18353 DVDD.n7998 DVDD.n7997 0.00263
R18354 DVDD.n7851 DVDD.n2151 0.00263
R18355 DVDD.n7851 DVDD.n7850 0.00263
R18356 DVDD.n7886 DVDD.n2101 0.00263
R18357 DVDD.n7886 DVDD.n7885 0.00263
R18358 DVDD.n7926 DVDD.n1171 0.00263
R18359 DVDD.n7927 DVDD.n7926 0.00263
R18360 DVDD.n7954 DVDD.n2043 0.00263
R18361 DVDD.n7954 DVDD.n7951 0.00263
R18362 DVDD.n3238 DVDD.n3227 0.00263
R18363 DVDD.n3297 DVDD.n3238 0.00263
R18364 DVDD.n3362 DVDD.n3344 0.00263
R18365 DVDD.n3369 DVDD.n3362 0.00263
R18366 DVDD.n6626 DVDD.n1132 0.00263
R18367 DVDD.n6627 DVDD.n6626 0.00263
R18368 DVDD.n6481 DVDD.n3408 0.00263
R18369 DVDD.n6593 DVDD.n6481 0.00263
R18370 DVDD.n6153 DVDD.n4283 0.00263
R18371 DVDD.n6153 DVDD.n6152 0.00263
R18372 DVDD.n6186 DVDD.n3560 0.00263
R18373 DVDD.n6188 DVDD.n3560 0.00263
R18374 DVDD.n6420 DVDD.n1070 0.00263
R18375 DVDD.n6421 DVDD.n6420 0.00263
R18376 DVDD.n3549 DVDD.n3534 0.00263
R18377 DVDD.n6387 DVDD.n3549 0.00263
R18378 DVDD.n6234 DVDD.n6233 0.0026
R18379 DVDD.n2199 DVDD.n1585 0.00254
R18380 DVDD.n2208 DVDD.n2200 0.00254
R18381 DVDD.n7791 DVDD.n7790 0.00254
R18382 DVDD.n3095 DVDD.n2198 0.00254
R18383 DVDD.n6102 DVDD.n6101 0.00254
R18384 DVDD.n3498 DVDD.n3495 0.00251708
R18385 DVDD.n7225 DVDD.n7030 0.00251
R18386 DVDD.n7269 DVDD.n7107 0.00251
R18387 DVDD.n8345 DVDD.n1530 0.00251
R18388 DVDD.n8321 DVDD.n8320 0.00251
R18389 DVDD.n7551 DVDD.n2508 0.00251
R18390 DVDD.n7594 DVDD.n2472 0.00251
R18391 DVDD.n2375 DVDD.n2372 0.00251
R18392 DVDD.n7778 DVDD.n2236 0.00251
R18393 DVDD.n7014 DVDD.n2522 0.00251
R18394 DVDD.n7003 DVDD.n7002 0.00251
R18395 DVDD.n6979 DVDD.n6935 0.00251
R18396 DVDD.n7807 DVDD.n2171 0.00251
R18397 DVDD.n5525 DVDD.n5495 0.00251
R18398 DVDD.n6751 DVDD.n3025 0.00251
R18399 DVDD.n2660 DVDD.n2656 0.00251
R18400 DVDD.n3185 DVDD.n3122 0.00251
R18401 DVDD.n5411 DVDD.n4472 0.00251
R18402 DVDD.n5676 DVDD.n2962 0.00251
R18403 DVDD.n2808 DVDD.n2804 0.00251
R18404 DVDD.n6114 DVDD.n4305 0.00251
R18405 DVDD.n9616 DVDD.n108 0.00251
R18406 DVDD.n9425 DVDD.n358 0.00251
R18407 DVDD.n2893 DVDD.n228 0.00251
R18408 DVDD.n9346 DVDD.n103 0.00251
R18409 DVDD.n9333 DVDD.n200 0.00251
R18410 DVDD.n9563 DVDD.n226 0.00251
R18411 DVDD.n309 DVDD.n103 0.00251
R18412 DVDD.n9429 DVDD.n200 0.00251
R18413 DVDD.n9563 DVDD.n222 0.00251
R18414 DVDD.n9616 DVDD.n120 0.00251
R18415 DVDD.n9425 DVDD.n373 0.00251
R18416 DVDD.n4148 DVDD.n228 0.00251
R18417 DVDD.n9616 DVDD.n124 0.00251
R18418 DVDD.n9430 DVDD.n9425 0.00251
R18419 DVDD.n242 DVDD.n228 0.00251
R18420 DVDD.n959 DVDD.n103 0.00251
R18421 DVDD.n972 DVDD.n200 0.00251
R18422 DVDD.n9563 DVDD.n215 0.00251
R18423 DVDD.n4018 DVDD.n103 0.00251
R18424 DVDD.n4081 DVDD.n200 0.00251
R18425 DVDD.n9563 DVDD.n218 0.00251
R18426 DVDD.n9616 DVDD.n116 0.00251
R18427 DVDD.n9425 DVDD.n352 0.00251
R18428 DVDD.n1037 DVDD.n228 0.00251
R18429 DVDD.n7505 DVDD.n7076 0.00249286
R18430 DVDD.n7487 DVDD.n7104 0.00249286
R18431 DVDD.n8369 DVDD.n1520 0.00249286
R18432 DVDD.n7431 DVDD.n7333 0.00249286
R18433 DVDD.n4709 DVDD.n4625 0.00249286
R18434 DVDD.n4819 DVDD.n4728 0.00249286
R18435 DVDD.n5157 DVDD.n5115 0.00249286
R18436 DVDD.n5082 DVDD.n4862 0.00249286
R18437 DVDD.n5249 DVDD.n4551 0.00249286
R18438 DVDD.n4788 DVDD.n4787 0.00249286
R18439 DVDD.n9284 DVDD.n9243 0.00249286
R18440 DVDD.n9210 DVDD.n489 0.00249286
R18441 DVDD.n6230 DVDD.n3862 0.00246875
R18442 DVDD.n3506 DVDD.n1095 0.00246875
R18443 DVDD.n6002 DVDD.n5928 0.00246875
R18444 DVDD.n2785 DVDD.n2777 0.00246875
R18445 DVDD.n8651 DVDD.n1237 0.00245
R18446 DVDD.n8654 DVDD.n1198 0.00245
R18447 DVDD.n8657 DVDD.n1159 0.00245
R18448 DVDD.n8660 DVDD.n1120 0.00245
R18449 DVDD.n8666 DVDD.n1058 0.00245
R18450 DVDD.n4534 DVDD.n429 0.00244882
R18451 DVDD.n4532 DVDD.n435 0.00244882
R18452 DVDD.n4531 DVDD.n4530 0.00244882
R18453 DVDD.n4529 DVDD.n408 0.00244882
R18454 DVDD.n9363 DVDD.n9362 0.00244882
R18455 DVDD.n9365 DVDD.n107 0.00244882
R18456 DVDD.n9367 DVDD.n130 0.00244882
R18457 DVDD.n9370 DVDD.n406 0.00244882
R18458 DVDD.n9372 DVDD.n9371 0.00244882
R18459 DVDD.n9374 DVDD.n9373 0.00244882
R18460 DVDD.n9377 DVDD.n147 0.00244882
R18461 DVDD.n720 DVDD.n585 0.00244882
R18462 DVDD.n8801 DVDD.n60 0.00244882
R18463 DVDD.n8740 DVDD.n8739 0.00244882
R18464 DVDD.n3636 DVDD.n3635 0.00244882
R18465 DVDD.n3841 DVDD.n3566 0.00244882
R18466 DVDD.n6516 DVDD.n2081 0.00244882
R18467 DVDD.n8979 DVDD.n555 0.00244882
R18468 DVDD.n535 DVDD.n525 0.00244882
R18469 DVDD.n4065 DVDD.n4064 0.00244882
R18470 DVDD.n4161 DVDD.n4160 0.00244882
R18471 DVDD.n6028 DVDD.n3963 0.00244882
R18472 DVDD.n3279 DVDD.n2122 0.00244882
R18473 DVDD.n5081 DVDD.n4868 0.00244882
R18474 DVDD.n4916 DVDD.n484 0.00244882
R18475 DVDD.n344 DVDD.n332 0.00244882
R18476 DVDD.n249 DVDD.n246 0.00244882
R18477 DVDD.n5795 DVDD.n4310 0.00244882
R18478 DVDD.n3170 DVDD.n2178 0.00244882
R18479 DVDD.n5123 DVDD.n4577 0.00244882
R18480 DVDD.n9250 DVDD.n464 0.00244882
R18481 DVDD.n9585 DVDD.n172 0.00244882
R18482 DVDD.n2904 DVDD.n2901 0.00244882
R18483 DVDD.n2855 DVDD.n2825 0.00244882
R18484 DVDD.n2700 DVDD.n2647 0.00244882
R18485 DVDD.n7241 DVDD.n2468 0.00238
R18486 DVDD.n7598 DVDD.n7597 0.00238
R18487 DVDD.n2616 DVDD.n2467 0.00238
R18488 DVDD.n6748 DVDD.n6747 0.00238
R18489 DVDD.n5712 DVDD.n4448 0.00238
R18490 DVDD.n8889 DVDD 0.0023
R18491 DVDD.n8203 DVDD 0.0023
R18492 DVDD.n5994 DVDD.n3913 0.0023
R18493 DVDD.n5995 DVDD.n3912 0.0023
R18494 DVDD.n6082 DVDD.n6081 0.0023
R18495 DVDD.n5675 DVDD.n4448 0.0023
R18496 DVDD.n5649 DVDD.n5644 0.0023
R18497 DVDD.n9699 DVDD 0.0023
R18498 DVDD.n6097 DVDD.n5765 0.00224375
R18499 DVDD.n5657 DVDD.n5650 0.00224375
R18500 DVDD.n6771 DVDD.n3008 0.00224375
R18501 DVDD.n5689 DVDD.n2743 0.00224375
R18502 DVDD.n7225 DVDD.n7029 0.00221
R18503 DVDD.n8345 DVDD.n1529 0.00221
R18504 DVDD.n8320 DVDD.n1619 0.00221
R18505 DVDD.n7551 DVDD.n7550 0.00221
R18506 DVDD.n7679 DVDD.n2375 0.00221
R18507 DVDD.n7776 DVDD.n2236 0.00221
R18508 DVDD.n7014 DVDD.n2521 0.00221
R18509 DVDD.n6982 DVDD.n6935 0.00221
R18510 DVDD.n7807 DVDD.n7806 0.00221
R18511 DVDD.n5525 DVDD.n5493 0.00221
R18512 DVDD.n6924 DVDD.n2660 0.00221
R18513 DVDD.n6704 DVDD.n3185 0.00221
R18514 DVDD.n5411 DVDD.n4471 0.00221
R18515 DVDD.n6856 DVDD.n2808 0.00221
R18516 DVDD.n6114 DVDD.n6113 0.00221
R18517 DVDD.n9613 DVDD.n108 0.00221
R18518 DVDD.n9391 DVDD.n358 0.00221
R18519 DVDD.n6791 DVDD.n2893 0.00221
R18520 DVDD.n4095 DVDD.n120 0.00221
R18521 DVDD.n4079 DVDD.n373 0.00221
R18522 DVDD.n4215 DVDD.n4148 0.00221
R18523 DVDD.n9457 DVDD.n124 0.00221
R18524 DVDD.n9431 DVDD.n9430 0.00221
R18525 DVDD.n243 DVDD.n242 0.00221
R18526 DVDD.n8765 DVDD.n116 0.00221
R18527 DVDD.n8735 DVDD.n352 0.00221
R18528 DVDD.n8682 DVDD.n1037 0.00221
R18529 DVDD.n8818 DVDD.n64 0.00209449
R18530 DVDD.n3858 DVDD.n3562 0.00209449
R18531 DVDD.n6531 DVDD.n3355 0.00209449
R18532 DVDD.n6499 DVDD.n2077 0.00209449
R18533 DVDD.n9090 DVDD.n530 0.00209449
R18534 DVDD.n6011 DVDD.n3959 0.00209449
R18535 DVDD.n3239 DVDD.n3225 0.00209449
R18536 DVDD.n3262 DVDD.n2126 0.00209449
R18537 DVDD.n4933 DVDD.n488 0.00209449
R18538 DVDD.n5778 DVDD.n4306 0.00209449
R18539 DVDD.n3128 DVDD.n3120 0.00209449
R18540 DVDD.n3153 DVDD.n2174 0.00209449
R18541 DVDD.n9252 DVDD.n9247 0.00209449
R18542 DVDD.n2838 DVDD.n2821 0.00209449
R18543 DVDD.n2716 DVDD.n2670 0.00209449
R18544 DVDD.n2683 DVDD.n2636 0.00209449
R18545 DVDD.n8293 DVDD.n1660 0.00209
R18546 DVDD.n8290 DVDD.n1665 0.00209
R18547 DVDD.n8118 DVDD.n1899 0.00209
R18548 DVDD.n8108 DVDD.n1891 0.00209
R18549 DVDD.n8651 DVDD.n1249 0.00209
R18550 DVDD.n8152 DVDD.n1236 0.00209
R18551 DVDD.n8191 DVDD.n1814 0.00209
R18552 DVDD.n8176 DVDD.n1800 0.00209
R18553 DVDD.n7749 DVDD.n2285 0.00209
R18554 DVDD.n2307 DVDD.n2292 0.00209
R18555 DVDD.n8057 DVDD.n1947 0.00209
R18556 DVDD.n8054 DVDD.n1954 0.00209
R18557 DVDD.n8654 DVDD.n1210 0.00209
R18558 DVDD.n8032 DVDD.n1197 0.00209
R18559 DVDD.n8010 DVDD.n7961 0.00209
R18560 DVDD.n8008 DVDD.n7998 0.00209
R18561 DVDD.n7842 DVDD.n2151 0.00209
R18562 DVDD.n7850 DVDD.n2149 0.00209
R18563 DVDD.n7890 DVDD.n2101 0.00209
R18564 DVDD.n7885 DVDD.n2096 0.00209
R18565 DVDD.n8657 DVDD.n1171 0.00209
R18566 DVDD.n7927 DVDD.n1158 0.00209
R18567 DVDD.n7958 DVDD.n2043 0.00209
R18568 DVDD.n7951 DVDD.n2029 0.00209
R18569 DVDD.n6676 DVDD.n3227 0.00209
R18570 DVDD.n6674 DVDD.n3297 0.00209
R18571 DVDD.n6650 DVDD.n3344 0.00209
R18572 DVDD.n3369 DVDD.n3357 0.00209
R18573 DVDD.n8660 DVDD.n1132 0.00209
R18574 DVDD.n6627 DVDD.n1119 0.00209
R18575 DVDD.n6605 DVDD.n3408 0.00209
R18576 DVDD.n6603 DVDD.n6593 0.00209
R18577 DVDD.n4283 DVDD.n4282 0.00209
R18578 DVDD.n6152 DVDD.n4285 0.00209
R18579 DVDD.n6186 DVDD.n3557 0.00209
R18580 DVDD.n6188 DVDD.n3558 0.00209
R18581 DVDD.n8666 DVDD.n1070 0.00209
R18582 DVDD.n6421 DVDD.n1057 0.00209
R18583 DVDD.n6399 DVDD.n3534 0.00209
R18584 DVDD.n6397 DVDD.n6387 0.00209
R18585 DVDD.n6882 DVDD.n2787 0.002
R18586 DVDD.n6101 DVDD.n4392 0.002
R18587 DVDD.n9354 DVDD.n418 0.002
R18588 DVDD.n9579 DVDD.n195 0.002
R18589 DVDD.n9561 DVDD.n239 0.002
R18590 DVDD.n9354 DVDD.n9325 0.002
R18591 DVDD.n9579 DVDD.n9578 0.002
R18592 DVDD.n9561 DVDD.n210 0.002
R18593 DVDD.n9354 DVDD.n424 0.002
R18594 DVDD.n9579 DVDD.n185 0.002
R18595 DVDD.n9561 DVDD.n235 0.002
R18596 DVDD.n9354 DVDD.n420 0.002
R18597 DVDD.n9579 DVDD.n191 0.002
R18598 DVDD.n9561 DVDD.n232 0.002
R18599 DVDD.n7223 DVDD.n7222 0.00197
R18600 DVDD.n7281 DVDD.n7272 0.00197
R18601 DVDD.n8356 DVDD.n8348 0.00197
R18602 DVDD.n1629 DVDD.n1628 0.00197
R18603 DVDD.n7545 DVDD.n7534 0.00197
R18604 DVDD.n7587 DVDD.n7576 0.00197
R18605 DVDD.n7653 DVDD.n2374 0.00197
R18606 DVDD.n7780 DVDD.n2217 0.00197
R18607 DVDD.n7020 DVDD.n7017 0.00197
R18608 DVDD.n2610 DVDD.n2609 0.00197
R18609 DVDD.n6976 DVDD.n6934 0.00197
R18610 DVDD.n7799 DVDD.n7798 0.00197
R18611 DVDD.n5527 DVDD.n5492 0.00197
R18612 DVDD.n6765 DVDD.n6754 0.00197
R18613 DVDD.n6729 DVDD.n2659 0.00197
R18614 DVDD.n3189 DVDD.n3184 0.00197
R18615 DVDD.n5413 DVDD.n4470 0.00197
R18616 DVDD.n5401 DVDD.n5400 0.00197
R18617 DVDD.n5731 DVDD.n2807 0.00197
R18618 DVDD.n6111 DVDD.n6106 0.00197
R18619 DVDD.n9361 DVDD.n106 0.00197
R18620 DVDD.n9398 DVDD.n201 0.00197
R18621 DVDD.n5287 DVDD.n212 0.00197
R18622 DVDD.n4102 DVDD.n121 0.00197
R18623 DVDD.n4072 DVDD.n371 0.00197
R18624 DVDD.n4145 DVDD.n4144 0.00197
R18625 DVDD.n296 DVDD.n123 0.00197
R18626 DVDD.n363 DVDD.n361 0.00197
R18627 DVDD.n9505 DVDD.n9504 0.00197
R18628 DVDD.n8772 DVDD.n117 0.00197
R18629 DVDD.n8718 DVDD.n349 0.00197
R18630 DVDD.n8686 DVDD.n1012 0.00197
R18631 DVDD.n6752 DVDD.n2615 0.00194
R18632 DVDD.n7001 DVDD.n7000 0.00194
R18633 DVDD.n7595 DVDD.n2471 0.00194
R18634 DVDD.n7270 DVDD.n7268 0.00194
R18635 DVDD.n7269 DVDD.n2474 0.00194
R18636 DVDD.n7594 DVDD.n7593 0.00194
R18637 DVDD.n7002 DVDD.n2473 0.00194
R18638 DVDD.n6751 DVDD.n6750 0.00194
R18639 DVDD.n5709 DVDD.n4449 0.00194
R18640 DVDD.n5677 DVDD.n5676 0.00194
R18641 DVDD.n6214 DVDD.n1058 0.00185
R18642 DVDD.n6424 DVDD.n3509 0.00185
R18643 DVDD.n9354 DVDD.n425 0.00184
R18644 DVDD.n9579 DVDD.n196 0.00184
R18645 DVDD.n9561 DVDD.n9560 0.00184
R18646 DVDD.n9354 DVDD.n9347 0.00184
R18647 DVDD.n9579 DVDD.n198 0.00184
R18648 DVDD.n9561 DVDD.n237 0.00184
R18649 DVDD.n9354 DVDD.n423 0.00184
R18650 DVDD.n9579 DVDD.n186 0.00184
R18651 DVDD.n9561 DVDD.n234 0.00184
R18652 DVDD.n9354 DVDD.n419 0.00184
R18653 DVDD.n9579 DVDD.n190 0.00184
R18654 DVDD.n9561 DVDD.n231 0.00184
R18655 DVDD.n6461 DVDD.n3483 0.00174867
R18656 DVDD.n5231 DVDD.n4552 0.00174016
R18657 DVDD.n5233 DVDD.n4550 0.00174016
R18658 DVDD.n5235 DVDD.n4553 0.00174016
R18659 DVDD.n5237 DVDD.n4549 0.00174016
R18660 DVDD.n5239 DVDD.n4554 0.00174016
R18661 DVDD.n5241 DVDD.n4548 0.00174016
R18662 DVDD.n5243 DVDD.n4555 0.00174016
R18663 DVDD.n4556 DVDD.n4547 0.00174016
R18664 DVDD.n5248 DVDD.n5247 0.00174016
R18665 DVDD.n4546 DVDD.n4541 0.00174016
R18666 DVDD.n5251 DVDD.n5250 0.00174016
R18667 DVDD.n8817 DVDD.n67 0.00174016
R18668 DVDD.n3857 DVDD.n3817 0.00174016
R18669 DVDD.n6532 DVDD.n3333 0.00174016
R18670 DVDD.n6500 DVDD.n2087 0.00174016
R18671 DVDD.n9089 DVDD.n529 0.00174016
R18672 DVDD.n6012 DVDD.n3957 0.00174016
R18673 DVDD.n6675 DVDD.n3296 0.00174016
R18674 DVDD.n3263 DVDD.n2139 0.00174016
R18675 DVDD.n4932 DVDD.n491 0.00174016
R18676 DVDD.n5779 DVDD.n4386 0.00174016
R18677 DVDD.n3129 DVDD.n3098 0.00174016
R18678 DVDD.n3154 DVDD.n2184 0.00174016
R18679 DVDD.n9253 DVDD.n9246 0.00174016
R18680 DVDD.n2839 DVDD.n2818 0.00174016
R18681 DVDD.n2717 DVDD.n2674 0.00174016
R18682 DVDD.n2684 DVDD.n2631 0.00174016
R18683 DVDD.n8202 DVDD 0.0017
R18684 DVDD.n6710 DVDD.n6709 0.0017
R18685 DVDD.n7788 DVDD.n2203 0.0017
R18686 DVDD.n7634 DVDD.n1584 0.0017
R18687 DVDD.n8327 DVDD.n8326 0.0017
R18688 DVDD.n1587 DVDD.n1580 0.0017
R18689 DVDD.n7785 DVDD.n2206 0.0017
R18690 DVDD.n7787 DVDD.n7786 0.0017
R18691 DVDD.n6711 DVDD.n2205 0.0017
R18692 DVDD.n6159 DVDD.n3914 0.0017
R18693 DVDD.n5648 DVDD.n5647 0.0017
R18694 DVDD.n5756 DVDD.n4394 0.0017
R18695 DVDD.n5759 DVDD.n5757 0.0017
R18696 DVDD.n9327 DVDD.n129 0.00167
R18697 DVDD.n9586 DVDD.n170 0.00167
R18698 DVDD.n6788 DVDD.n2894 0.00167
R18699 DVDD.n4094 DVDD.n4017 0.00167
R18700 DVDD.n4080 DVDD.n4027 0.00167
R18701 DVDD.n4214 DVDD.n4149 0.00167
R18702 DVDD.n9456 DVDD.n308 0.00167
R18703 DVDD.n347 DVDD.n346 0.00167
R18704 DVDD.n9557 DVDD.n9556 0.00167
R18705 DVDD.n8762 DVDD.n850 0.00167
R18706 DVDD.n8738 DVDD.n883 0.00167
R18707 DVDD.n3742 DVDD.n1038 0.00167
R18708 DVDD DVDD.n6449 0.00165261
R18709 DVDD.n3489 DVDD 0.00165261
R18710 DVDD.n8698 DVDD.n1005 0.001625
R18711 DVDD.n917 DVDD.n903 0.001625
R18712 DVDD.n6242 DVDD.n6239 0.001625
R18713 DVDD.n2783 DVDD.n2778 0.001625
R18714 DVDD.n396 DVDD.n395 0.001625
R18715 DVDD.n5275 DVDD.n5274 0.001625
R18716 DVDD.n9314 DVDD.n441 0.001625
R18717 DVDD.n97 DVDD.n83 0.001625
R18718 DVDD.n1688 DVDD.n1678 0.00155
R18719 DVDD.n8120 DVDD.n1853 0.00155
R18720 DVDD.n8154 DVDD.n1235 0.00155
R18721 DVDD.n8173 DVDD.n1799 0.00155
R18722 DVDD.n7747 DVDD.n2295 0.00155
R18723 DVDD.n8052 DVDD.n1973 0.00155
R18724 DVDD.n8019 DVDD.n1196 0.00155
R18725 DVDD.n8007 DVDD.n7985 0.00155
R18726 DVDD.n7853 DVDD.n2120 0.00155
R18727 DVDD.n7893 DVDD.n2074 0.00155
R18728 DVDD.n7929 DVDD.n1157 0.00155
R18729 DVDD.n7948 DVDD.n2028 0.00155
R18730 DVDD.n6673 DVDD.n3237 0.00155
R18731 DVDD.n6648 DVDD.n3363 0.00155
R18732 DVDD.n6614 DVDD.n1118 0.00155
R18733 DVDD.n6602 DVDD.n6485 0.00155
R18734 DVDD.n6155 DVDD.n3946 0.00155
R18735 DVDD.n6334 DVDD.n3561 0.00155
R18736 DVDD.n6408 DVDD.n1056 0.00155
R18737 DVDD.n6396 DVDD.n3551 0.00155
R18738 DVDD.n7240 DVDD.n2468 0.00146
R18739 DVDD.n7597 DVDD.n7596 0.00146
R18740 DVDD.n2614 DVDD.n2467 0.00146
R18741 DVDD.n6749 DVDD.n6748 0.00146
R18742 DVDD.n6671 DVDD.n2117 0.00146
R18743 DVDD.n7856 DVDD.n7855 0.00146
R18744 DVDD.n2315 DVDD.n1927 0.00146
R18745 DVDD.n1922 DVDD.n1917 0.00146
R18746 DVDD.n1921 DVDD.n1916 0.00146
R18747 DVDD.n2316 DVDD.n1929 0.00146
R18748 DVDD.n7854 DVDD.n2116 0.00146
R18749 DVDD.n6670 DVDD.n6669 0.00146
R18750 DVDD.n5388 DVDD.n4448 0.00146
R18751 DVDD.n6157 DVDD.n3913 0.00146
R18752 DVDD.n6156 DVDD.n3912 0.00146
R18753 DVDD.n7508 DVDD.n7043 0.00143
R18754 DVDD.n7285 DVDD.n7120 0.00143
R18755 DVDD.n8358 DVDD.n1544 0.00143
R18756 DVDD.n8323 DVDD.n1600 0.00143
R18757 DVDD.n7548 DVDD.n7523 0.00143
R18758 DVDD.n7590 DVDD.n7565 0.00143
R18759 DVDD.n7660 DVDD.n7656 0.00143
R18760 DVDD.n7781 DVDD.n2207 0.00143
R18761 DVDD.n7024 DVDD.n2536 0.00143
R18762 DVDD.n7005 DVDD.n2573 0.00143
R18763 DVDD.n6985 DVDD.n2638 0.00143
R18764 DVDD.n7803 DVDD.n7794 0.00143
R18765 DVDD.n5614 DVDD.n5530 0.00143
R18766 DVDD.n6768 DVDD.n3038 0.00143
R18767 DVDD.n6731 DVDD.n2657 0.00143
R18768 DVDD.n6706 DVDD.n3109 0.00143
R18769 DVDD.n5466 DVDD.n5416 0.00143
R18770 DVDD.n6774 DVDD.n2975 0.00143
R18771 DVDD.n4438 DVDD.n2805 0.00143
R18772 DVDD.n6105 DVDD.n4388 0.00143
R18773 DVDD.n4528 DVDD.n409 0.00143
R18774 DVDD.n9418 DVDD.n202 0.00143
R18775 DVDD.n5284 DVDD.n211 0.00143
R18776 DVDD.n4103 DVDD.n4001 0.00143
R18777 DVDD.n4071 DVDD.n3991 0.00143
R18778 DVDD.n4143 DVDD.n3977 0.00143
R18779 DVDD.n9466 DVDD.n294 0.00143
R18780 DVDD.n362 DVDD.n281 0.00143
R18781 DVDD.n9503 DVDD.n268 0.00143
R18782 DVDD.n9623 DVDD.n89 0.00143
R18783 DVDD.n8715 DVDD.n891 0.00143
R18784 DVDD.n1034 DVDD.n1011 0.00143
R18785 DVDD.n6211 DVDD.n6210 0.0014
R18786 DVDD.n721 DVDD.n586 0.00138583
R18787 DVDD.n8802 DVDD.n70 0.00138583
R18788 DVDD.n8741 DVDD.n877 0.00138583
R18789 DVDD.n3741 DVDD.n3740 0.00138583
R18790 DVDD.n3842 DVDD.n3814 0.00138583
R18791 DVDD.n6515 DVDD.n2084 0.00138583
R18792 DVDD.n8978 DVDD.n554 0.00138583
R18793 DVDD.n9174 DVDD.n9125 0.00138583
R18794 DVDD.n4063 DVDD.n4062 0.00138583
R18795 DVDD.n4159 DVDD.n4158 0.00138583
R18796 DVDD.n6027 DVDD.n3954 0.00138583
R18797 DVDD.n3278 DVDD.n2142 0.00138583
R18798 DVDD.n4875 DVDD.n4857 0.00138583
R18799 DVDD.n4917 DVDD.n494 0.00138583
R18800 DVDD.n9438 DVDD.n9437 0.00138583
R18801 DVDD.n9555 DVDD.n9554 0.00138583
R18802 DVDD.n5794 DVDD.n4383 0.00138583
R18803 DVDD.n3169 DVDD.n2181 0.00138583
R18804 DVDD.n5122 DVDD.n4576 0.00138583
R18805 DVDD.n9283 DVDD.n9282 0.00138583
R18806 DVDD.n9590 DVDD.n165 0.00138583
R18807 DVDD.n6787 DVDD.n6786 0.00138583
R18808 DVDD.n2854 DVDD.n2815 0.00138583
R18809 DVDD.n2699 DVDD.n2634 0.00138583
R18810 DVDD DVDD.n6600 0.00134
R18811 DVDD DVDD.n7947 0.00134
R18812 DVDD DVDD.n8005 0.00134
R18813 DVDD DVDD.n8172 0.00134
R18814 DVDD DVDD.n6394 0.00134
R18815 DVDD.n2199 DVDD.n1583 0.0013
R18816 DVDD.n7633 DVDD.n2200 0.0013
R18817 DVDD.n7790 DVDD.n7789 0.0013
R18818 DVDD.n3094 DVDD.n2198 0.0013
R18819 DVDD.n6101 DVDD.n4391 0.0013
R18820 DVDD.n6445 DVDD 0.00126841
R18821 DVDD.n6631 DVDD.n6630 0.00122
R18822 DVDD.n7911 DVDD.n2004 0.00122
R18823 DVDD.n8036 DVDD.n8035 0.00122
R18824 DVDD.n8138 DVDD.n1841 0.00122
R18825 DVDD.n8137 DVDD.n1237 0.00122
R18826 DVDD.n8037 DVDD.n1198 0.00122
R18827 DVDD.n7910 DVDD.n1159 0.00122
R18828 DVDD.n6632 DVDD.n1120 0.00122
R18829 DVDD.n6424 DVDD.n3510 0.00122
R18830 DVDD.n6205 DVDD.n1058 0.00122
R18831 DVDD.n394 DVDD.n206 0.00119
R18832 DVDD.n5269 DVDD.n207 0.00119
R18833 DVDD.n4131 DVDD.n4130 0.00119
R18834 DVDD.n3986 DVDD.n3981 0.00119
R18835 DVDD.n9491 DVDD.n9490 0.00119
R18836 DVDD.n277 DVDD.n272 0.00119
R18837 DVDD.n8706 DVDD.n907 0.00119
R18838 DVDD.n8703 DVDD.n911 0.00119
R18839 DVDD.n8673 DVDD.n8672 0.001175
R18840 DVDD.n8746 DVDD.n876 0.001175
R18841 DVDD.n6325 DVDD.n3866 0.001175
R18842 DVDD.n2796 DVDD.n2795 0.001175
R18843 DVDD.n179 DVDD.n178 0.001175
R18844 DVDD.n6780 DVDD.n2907 0.001175
R18845 DVDD.n9604 DVDD.n139 0.001175
R18846 DVDD.n8756 DVDD.n8755 0.001175
R18847 DVDD.n8079 DVDD.n1923 0.00114
R18848 DVDD.n8078 DVDD.n1925 0.00114
R18849 DVDD.n2119 DVDD.n1924 0.00114
R18850 DVDD.n3315 DVDD.n3313 0.00114
R18851 DVDD.n6159 DVDD.n6158 0.00114
R18852 DVDD.n9328 DVDD.n137 0.00113
R18853 DVDD.n9589 DVDD.n167 0.00113
R18854 DVDD.n5303 DVDD.n2898 0.00113
R18855 DVDD.n4042 DVDD.n4041 0.00113
R18856 DVDD.n4061 DVDD.n4026 0.00113
R18857 DVDD.n4153 DVDD.n4152 0.00113
R18858 DVDD.n9453 DVDD.n9452 0.00113
R18859 DVDD.n9439 DVDD.n330 0.00113
R18860 DVDD.n251 DVDD.n244 0.00113
R18861 DVDD.n942 DVDD.n853 0.00113
R18862 DVDD.n977 DVDD.n882 0.00113
R18863 DVDD.n3634 DVDD.n3591 0.00113
R18864 DVDD.n8170 DVDD 0.00106
R18865 DVDD.n8003 DVDD 0.00106
R18866 DVDD.n6598 DVDD 0.00106
R18867 DVDD.n6392 DVDD 0.00106
R18868 DVDD.n941 DVDD.n940 0.0010315
R18869 DVDD.n6264 DVDD.n3346 0.0010315
R18870 DVDD.n4043 DVDD.n4040 0.0010315
R18871 DVDD.n5955 DVDD.n3217 0.0010315
R18872 DVDD.n9451 DVDD.n314 0.0010315
R18873 DVDD.n5853 DVDD.n3111 0.0010315
R18874 DVDD.n9607 DVDD.n9606 0.0010315
R18875 DVDD.n6915 DVDD.n2662 0.0010315
R18876 DVDD.n5677 DVDD.n3000 0.00100625
R18877 DVDD.n6460 DVDD.n6459 0.000980256
R18878 DVDD.n8140 DVDD.n8139 0.00098
R18879 DVDD.n2003 DVDD.n1842 0.00098
R18880 DVDD.n7913 DVDD.n7912 0.00098
R18881 DVDD.n3384 DVDD.n2063 0.00098
R18882 DVDD.n6210 DVDD.n6209 0.00098
R18883 DVDD.n9599 DVDD.n146 0.00095
R18884 DVDD.n9596 DVDD.n151 0.00095
R18885 DVDD.n4045 DVDD.n4022 0.00095
R18886 DVDD.n4031 DVDD.n4023 0.00095
R18887 DVDD.n9445 DVDD.n9444 0.00095
R18888 DVDD.n337 DVDD.n323 0.00095
R18889 DVDD.n965 DVDD.n867 0.00095
R18890 DVDD.n8749 DVDD.n870 0.00095
R18891 DVDD.n434 DVDD.n428 0.00089
R18892 DVDD.n9415 DVDD.n203 0.00089
R18893 DVDD.n4516 DVDD.n4508 0.00089
R18894 DVDD.n4009 DVDD.n4000 0.00089
R18895 DVDD.n4124 DVDD.n4123 0.00089
R18896 DVDD.n3983 DVDD.n3982 0.00089
R18897 DVDD.n9467 DVDD.n293 0.00089
R18898 DVDD.n9484 DVDD.n9483 0.00089
R18899 DVDD.n274 DVDD.n273 0.00089
R18900 DVDD.n88 DVDD.n85 0.00089
R18901 DVDD.n919 DVDD.n894 0.00089
R18902 DVDD.n1032 DVDD.n1003 0.00089
R18903 DVDD.n3494 DVDD.n3493 0.000788154
R18904 DVDD.n7106 DVDD.n2474 0.00077
R18905 DVDD.n7593 DVDD.n7592 0.00077
R18906 DVDD.n2597 DVDD.n2473 0.00077
R18907 DVDD.n6750 DVDD.n3024 0.00077
R18908 DVDD.n5677 DVDD.n2961 0.00077
R18909 DVDD.n705 DVDD.n581 0.000677165
R18910 DVDD.n9628 DVDD.n82 0.000677165
R18911 DVDD.n997 DVDD.n996 0.000677165
R18912 DVDD.n3826 DVDD.n3569 0.000677165
R18913 DVDD.n9008 DVDD.n8973 0.000677165
R18914 DVDD.n4007 DVDD.n4004 0.000677165
R18915 DVDD.n4118 DVDD.n3994 0.000677165
R18916 DVDD.n6043 DVDD.n3966 0.000677165
R18917 DVDD.n5014 DVDD.n4859 0.000677165
R18918 DVDD.n301 DVDD.n300 0.000677165
R18919 DVDD.n9478 DVDD.n284 0.000677165
R18920 DVDD.n5810 DVDD.n4313 0.000677165
R18921 DVDD.n5152 DVDD.n5117 0.000677165
R18922 DVDD.n9315 DVDD.n437 0.000677165
R18923 DVDD.n9410 DVDD.n389 0.000677165
R18924 DVDD.n2870 DVDD.n2828 0.000677165
R18925 DVDD.n9698 DVDD 0.000671429
R18926 DVDD DVDD.n8890 0.000671429
R18927 DVDD.n8202 DVDD 0.000671429
R18928 DVDD.n9316 DVDD.n430 0.00065
R18929 DVDD.n393 DVDD.n385 0.00065
R18930 DVDD.n5272 DVDD.n208 0.00065
R18931 DVDD.n4110 DVDD.n3999 0.00065
R18932 DVDD.n3992 DVDD.n3985 0.00065
R18933 DVDD.n4137 DVDD.n4136 0.00065
R18934 DVDD.n9470 DVDD.n290 0.00065
R18935 DVDD.n282 DVDD.n276 0.00065
R18936 DVDD.n9497 DVDD.n9496 0.00065
R18937 DVDD.n9627 DVDD.n84 0.00065
R18938 DVDD.n995 DVDD.n906 0.00065
R18939 DVDD.n8700 DVDD.n912 0.00065
R18940 DVDD.n9329 DVDD.n145 0.00059
R18941 DVDD.n166 DVDD.n152 0.00059
R18942 DVDD.n5302 DVDD.n2906 0.00059
R18943 DVDD.n4046 DVDD.n4021 0.00059
R18944 DVDD.n4060 DVDD.n4059 0.00059
R18945 DVDD.n4208 DVDD.n4207 0.00059
R18946 DVDD.n322 DVDD.n313 0.00059
R18947 DVDD.n9440 DVDD.n329 0.00059
R18948 DVDD.n9548 DVDD.n252 0.00059
R18949 DVDD.n8753 DVDD.n866 0.00059
R18950 DVDD.n976 DVDD.n871 0.00059
R18951 DVDD.n8670 DVDD.n1051 0.00059
R18952 DVDD DVDD.n8170 0.00058
R18953 DVDD DVDD.n8003 0.00058
R18954 DVDD DVDD.n7945 0.00058
R18955 DVDD DVDD.n6598 0.00058
R18956 DVDD DVDD.n6392 0.00058
R18957 DVDD.n5657 DVDD.n5640 0.00055625
R18958 DVSS.n9388 DVSS.n379 20126
R18959 DVSS.n9388 DVSS.n9387 20126
R18960 DVSS.n7255 DVSS.n380 17859.7
R18961 DVSS.n7256 DVSS.n7255 17859.7
R18962 DVSS.n7256 DVSS.n379 6553.98
R18963 DVSS.n9387 DVSS.n380 6553.98
R18964 DVSS.n9386 DVSS.n9385 6266.18
R18965 DVSS.n750 DVSS.n381 6258.6
R18966 DVSS.n750 DVSS.n379 5490.26
R18967 DVSS.n9387 DVSS.n9386 5490.26
R18968 DVSS.n8297 DVSS.t3 3474.96
R18969 DVSS.n8318 DVSS.t3 3474.96
R18970 DVSS.n8462 DVSS.t37 2918.55
R18971 DVSS.n8500 DVSS.t37 2918.55
R18972 DVSS.n7261 DVSS.n6014 2402.48
R18973 DVSS.n7261 DVSS.n6015 2401.2
R18974 DVSS.n6014 DVSS.n2756 2400.01
R18975 DVSS.n6015 DVSS.n2756 2398.73
R18976 DVSS.n6013 DVSS.n2758 851.766
R18977 DVSS.n5005 DVSS.n2758 851.766
R18978 DVSS.n5006 DVSS.n5005 851.766
R18979 DVSS.n5006 DVSS.n2977 851.766
R18980 DVSS.n7264 DVSS.n2755 851.766
R18981 DVSS.n7264 DVSS.n7263 851.766
R18982 DVSS.n7254 DVSS.n2757 851.766
R18983 DVSS.n7262 DVSS.n2757 794.593
R18984 DVSS.n7255 DVSS.n7254 496.031
R18985 DVSS.n5898 DVSS.n2977 425.884
R18986 DVSS.n5898 DVSS.n2755 425.884
R18987 DVSS.n8501 DVSS.n1081 167.197
R18988 DVSS.n1150 DVSS.n1081 167.197
R18989 DVSS.n8461 DVSS.n1093 167.197
R18990 DVSS.n8499 DVSS.n1093 167.197
R18991 DVSS.n8319 DVSS.n1452 130.218
R18992 DVSS.n1477 DVSS.n1452 130.218
R18993 DVSS.n1473 DVSS.n1456 130.218
R18994 DVSS.n8317 DVSS.n1456 130.218
R18995 DVSS.n8297 DVSS.n1476 127.05
R18996 DVSS.n8318 DVSS.n1454 127.05
R18997 DVSS.n6014 DVSS.n6013 96.6714
R18998 DVSS.n1273 DVSS.n1272 93.6563
R18999 DVSS.n1273 DVSS.n1089 93.6563
R19000 DVSS.n8466 DVSS.n8464 93.6563
R19001 DVSS.n8466 DVSS.n8465 93.6563
R19002 DVSS.n8379 DVSS.n1148 93.6563
R19003 DVSS.n8379 DVSS.n1094 93.6563
R19004 DVSS.n8462 DVSS.n1147 85.7351
R19005 DVSS.n8500 DVSS.n1091 85.7351
R19006 DVSS.n8285 DVSS.n1478 75.5231
R19007 DVSS.n8285 DVSS.n1451 75.5231
R19008 DVSS.n8257 DVSS.n1474 75.5231
R19009 DVSS.n8257 DVSS.n8256 75.5231
R19010 DVSS.n8300 DVSS.n8299 75.5231
R19011 DVSS.n8300 DVSS.n1457 75.5231
R19012 DVSS.n7263 DVSS.n7262 57.1732
R19013 DVSS.n8501 DVSS.n1089 14.4308
R19014 DVSS.n8464 DVSS.n1146 14.4308
R19015 DVSS.n1272 DVSS.n1146 14.4308
R19016 DVSS.n1272 DVSS.n1150 14.4308
R19017 DVSS.n1094 DVSS.n1090 14.4308
R19018 DVSS.n8465 DVSS.n1090 14.4308
R19019 DVSS.n8465 DVSS.n1092 14.4308
R19020 DVSS.n1092 DVSS.n1089 14.4308
R19021 DVSS.n8461 DVSS.n1148 14.4308
R19022 DVSS.n8463 DVSS.n1148 14.4308
R19023 DVSS.n8464 DVSS.n8463 14.4308
R19024 DVSS.n8499 DVSS.n1094 14.4308
R19025 DVSS.n5667 DVSS.n2485 12.7299
R19026 DVSS.n6642 DVSS.n6017 10.4832
R19027 DVSS.n6158 DVSS.n6016 10.4832
R19028 DVSS.n6158 DVSS.n6157 7.99992
R19029 DVSS.n6157 DVSS.n6017 7.96398
R19030 DVSS.n9385 DVSS.n381 7.57947
R19031 DVSS.n7257 DVSS.n6643 7.08357
R19032 DVSS.n7260 DVSS.n7259 7.08357
R19033 DVSS.n8319 DVSS.n1451 6.79968
R19034 DVSS.n8296 DVSS.n1474 6.79968
R19035 DVSS.n8296 DVSS.n1478 6.79968
R19036 DVSS.n1478 DVSS.n1477 6.79968
R19037 DVSS.n1457 DVSS.n1453 6.79968
R19038 DVSS.n8256 DVSS.n1453 6.79968
R19039 DVSS.n8256 DVSS.n1455 6.79968
R19040 DVSS.n1455 DVSS.n1451 6.79968
R19041 DVSS.n8299 DVSS.n1473 6.79968
R19042 DVSS.n8299 DVSS.n8298 6.79968
R19043 DVSS.n8298 DVSS.n1474 6.79968
R19044 DVSS.n8317 DVSS.n1457 6.79968
R19045 DVSS.n6346 DVSS.n6345 6.22149
R19046 DVSS.n6643 DVSS.n6642 6.10967
R19047 DVSS.n7260 DVSS.n6016 6.10909
R19048 DVSS.n7259 DVSS.n7258 5.11349
R19049 DVSS.n7258 DVSS.n7257 5.07814
R19050 DVSS.n3412 DVSS.n3401 4.5005
R19051 DVSS.n5307 DVSS.n3412 4.5005
R19052 DVSS.n3412 DVSS.n3405 4.5005
R19053 DVSS.n5305 DVSS.n3412 4.5005
R19054 DVSS.n3410 DVSS.n3401 4.5005
R19055 DVSS.n5307 DVSS.n3410 4.5005
R19056 DVSS.n3410 DVSS.n3405 4.5005
R19057 DVSS.n5305 DVSS.n3410 4.5005
R19058 DVSS.n3413 DVSS.n3401 4.5005
R19059 DVSS.n5307 DVSS.n3413 4.5005
R19060 DVSS.n3413 DVSS.n3405 4.5005
R19061 DVSS.n5305 DVSS.n3413 4.5005
R19062 DVSS.n3409 DVSS.n3401 4.5005
R19063 DVSS.n5307 DVSS.n3409 4.5005
R19064 DVSS.n3409 DVSS.n3405 4.5005
R19065 DVSS.n5305 DVSS.n3409 4.5005
R19066 DVSS.n3415 DVSS.n3401 4.5005
R19067 DVSS.n5307 DVSS.n3415 4.5005
R19068 DVSS.n5305 DVSS.n3415 4.5005
R19069 DVSS.n5307 DVSS.n3408 4.5005
R19070 DVSS.n5305 DVSS.n3408 4.5005
R19071 DVSS.n5307 DVSS.n3418 4.5005
R19072 DVSS.n5305 DVSS.n3418 4.5005
R19073 DVSS.n5307 DVSS.n3407 4.5005
R19074 DVSS.n5305 DVSS.n3407 4.5005
R19075 DVSS.n5307 DVSS.n3421 4.5005
R19076 DVSS.n5305 DVSS.n3421 4.5005
R19077 DVSS.n5307 DVSS.n3406 4.5005
R19078 DVSS.n5305 DVSS.n3406 4.5005
R19079 DVSS.n5307 DVSS.n5306 4.5005
R19080 DVSS.n5306 DVSS.n3405 4.5005
R19081 DVSS.n5306 DVSS.n5305 4.5005
R19082 DVSS.n5073 DVSS.n3423 4.5005
R19083 DVSS.n5130 DVSS.n3423 4.5005
R19084 DVSS.n5065 DVSS.n3423 4.5005
R19085 DVSS.n5080 DVSS.n5073 4.5005
R19086 DVSS.n5080 DVSS.n5065 4.5005
R19087 DVSS.n5078 DVSS.n5073 4.5005
R19088 DVSS.n5078 DVSS.n5065 4.5005
R19089 DVSS.n5077 DVSS.n5073 4.5005
R19090 DVSS.n5077 DVSS.n5065 4.5005
R19091 DVSS.n5075 DVSS.n5073 4.5005
R19092 DVSS.n5075 DVSS.n5065 4.5005
R19093 DVSS.n5073 DVSS.n5067 4.5005
R19094 DVSS.n5130 DVSS.n5067 4.5005
R19095 DVSS.n5067 DVSS.n5065 4.5005
R19096 DVSS.n5065 DVSS.n3355 4.5005
R19097 DVSS.n5130 DVSS.n3355 4.5005
R19098 DVSS.n5073 DVSS.n3355 4.5005
R19099 DVSS.n5128 DVSS.n3355 4.5005
R19100 DVSS.n5065 DVSS.n3357 4.5005
R19101 DVSS.n5130 DVSS.n3357 4.5005
R19102 DVSS.n5073 DVSS.n3357 4.5005
R19103 DVSS.n5128 DVSS.n3357 4.5005
R19104 DVSS.n5072 DVSS.n5065 4.5005
R19105 DVSS.n5130 DVSS.n5072 4.5005
R19106 DVSS.n5073 DVSS.n5072 4.5005
R19107 DVSS.n5128 DVSS.n5072 4.5005
R19108 DVSS.n5066 DVSS.n5065 4.5005
R19109 DVSS.n5130 DVSS.n5066 4.5005
R19110 DVSS.n5073 DVSS.n5066 4.5005
R19111 DVSS.n5128 DVSS.n5066 4.5005
R19112 DVSS.n5129 DVSS.n5065 4.5005
R19113 DVSS.n5130 DVSS.n5129 4.5005
R19114 DVSS.n5129 DVSS.n5073 4.5005
R19115 DVSS.n5129 DVSS.n5128 4.5005
R19116 DVSS.n8123 DVSS.n8122 4.5005
R19117 DVSS.n8122 DVSS.n1808 4.5005
R19118 DVSS.n8122 DVSS.n8121 4.5005
R19119 DVSS.n1821 DVSS.n1808 4.5005
R19120 DVSS.n8121 DVSS.n1821 4.5005
R19121 DVSS.n1823 DVSS.n1808 4.5005
R19122 DVSS.n8121 DVSS.n1823 4.5005
R19123 DVSS.n1820 DVSS.n1808 4.5005
R19124 DVSS.n8121 DVSS.n1820 4.5005
R19125 DVSS.n1824 DVSS.n1808 4.5005
R19126 DVSS.n8121 DVSS.n1824 4.5005
R19127 DVSS.n1819 DVSS.n1808 4.5005
R19128 DVSS.n8121 DVSS.n1819 4.5005
R19129 DVSS.n1825 DVSS.n1808 4.5005
R19130 DVSS.n8121 DVSS.n1825 4.5005
R19131 DVSS.n1818 DVSS.n1808 4.5005
R19132 DVSS.n8121 DVSS.n1818 4.5005
R19133 DVSS.n1826 DVSS.n1808 4.5005
R19134 DVSS.n8121 DVSS.n1826 4.5005
R19135 DVSS.n1817 DVSS.n1808 4.5005
R19136 DVSS.n8121 DVSS.n1817 4.5005
R19137 DVSS.n8120 DVSS.n1808 4.5005
R19138 DVSS.n8120 DVSS.n1832 4.5005
R19139 DVSS.n8121 DVSS.n8120 4.5005
R19140 DVSS.n1116 DVSS.n1106 4.5005
R19141 DVSS.n1116 DVSS.n1107 4.5005
R19142 DVSS.n8489 DVSS.n1116 4.5005
R19143 DVSS.n1113 DVSS.n1107 4.5005
R19144 DVSS.n8489 DVSS.n1113 4.5005
R19145 DVSS.n1119 DVSS.n1107 4.5005
R19146 DVSS.n8489 DVSS.n1119 4.5005
R19147 DVSS.n1112 DVSS.n1107 4.5005
R19148 DVSS.n8489 DVSS.n1112 4.5005
R19149 DVSS.n1121 DVSS.n1107 4.5005
R19150 DVSS.n1121 DVSS.n1105 4.5005
R19151 DVSS.n8489 DVSS.n1121 4.5005
R19152 DVSS.n8490 DVSS.n1106 4.5005
R19153 DVSS.n8490 DVSS.n1107 4.5005
R19154 DVSS.n8490 DVSS.n1105 4.5005
R19155 DVSS.n8490 DVSS.n8489 4.5005
R19156 DVSS.n8489 DVSS.n1101 4.5005
R19157 DVSS.n1105 DVSS.n1101 4.5005
R19158 DVSS.n1106 DVSS.n1101 4.5005
R19159 DVSS.n1111 DVSS.n1105 4.5005
R19160 DVSS.n8489 DVSS.n1111 4.5005
R19161 DVSS.n1124 DVSS.n1107 4.5005
R19162 DVSS.n8489 DVSS.n1124 4.5005
R19163 DVSS.n1109 DVSS.n1107 4.5005
R19164 DVSS.n8489 DVSS.n1109 4.5005
R19165 DVSS.n8488 DVSS.n1107 4.5005
R19166 DVSS.n8488 DVSS.n1105 4.5005
R19167 DVSS.n8489 DVSS.n8488 4.5005
R19168 DVSS.n4888 DVSS.n3620 4.5005
R19169 DVSS.n3620 DVSS.n3614 4.5005
R19170 DVSS.n3625 DVSS.n3620 4.5005
R19171 DVSS.n4888 DVSS.n3619 4.5005
R19172 DVSS.n3619 DVSS.n3614 4.5005
R19173 DVSS.n4883 DVSS.n3614 4.5005
R19174 DVSS.n4886 DVSS.n4883 4.5005
R19175 DVSS.n3630 DVSS.n3614 4.5005
R19176 DVSS.n4886 DVSS.n3630 4.5005
R19177 DVSS.n4885 DVSS.n3614 4.5005
R19178 DVSS.n4886 DVSS.n4885 4.5005
R19179 DVSS.n3629 DVSS.n3614 4.5005
R19180 DVSS.n4886 DVSS.n3629 4.5005
R19181 DVSS.n4888 DVSS.n3621 4.5005
R19182 DVSS.n3621 DVSS.n3614 4.5005
R19183 DVSS.n4886 DVSS.n3621 4.5005
R19184 DVSS.n4888 DVSS.n3616 4.5005
R19185 DVSS.n3616 DVSS.n3614 4.5005
R19186 DVSS.n3625 DVSS.n3616 4.5005
R19187 DVSS.n4886 DVSS.n3616 4.5005
R19188 DVSS.n4888 DVSS.n3622 4.5005
R19189 DVSS.n3622 DVSS.n3614 4.5005
R19190 DVSS.n3625 DVSS.n3622 4.5005
R19191 DVSS.n4886 DVSS.n3622 4.5005
R19192 DVSS.n4888 DVSS.n3615 4.5005
R19193 DVSS.n3615 DVSS.n3614 4.5005
R19194 DVSS.n3625 DVSS.n3615 4.5005
R19195 DVSS.n4886 DVSS.n3615 4.5005
R19196 DVSS.n4888 DVSS.n4887 4.5005
R19197 DVSS.n4887 DVSS.n3614 4.5005
R19198 DVSS.n4887 DVSS.n3625 4.5005
R19199 DVSS.n4887 DVSS.n4886 4.5005
R19200 DVSS.n4850 DVSS.n4849 4.5005
R19201 DVSS.n4849 DVSS.n3647 4.5005
R19202 DVSS.n4849 DVSS.n4848 4.5005
R19203 DVSS.n3659 DVSS.n3647 4.5005
R19204 DVSS.n4848 DVSS.n3659 4.5005
R19205 DVSS.n3661 DVSS.n3647 4.5005
R19206 DVSS.n4848 DVSS.n3661 4.5005
R19207 DVSS.n3658 DVSS.n3647 4.5005
R19208 DVSS.n4848 DVSS.n3658 4.5005
R19209 DVSS.n3662 DVSS.n3647 4.5005
R19210 DVSS.n4848 DVSS.n3662 4.5005
R19211 DVSS.n3657 DVSS.n3647 4.5005
R19212 DVSS.n4848 DVSS.n3657 4.5005
R19213 DVSS.n4847 DVSS.n3647 4.5005
R19214 DVSS.n4847 DVSS.n3666 4.5005
R19215 DVSS.n4848 DVSS.n4847 4.5005
R19216 DVSS.n4850 DVSS.n3651 4.5005
R19217 DVSS.n3651 DVSS.n3647 4.5005
R19218 DVSS.n3666 DVSS.n3651 4.5005
R19219 DVSS.n4848 DVSS.n3651 4.5005
R19220 DVSS.n4850 DVSS.n3650 4.5005
R19221 DVSS.n3650 DVSS.n3647 4.5005
R19222 DVSS.n3666 DVSS.n3650 4.5005
R19223 DVSS.n4848 DVSS.n3650 4.5005
R19224 DVSS.n4850 DVSS.n3649 4.5005
R19225 DVSS.n3649 DVSS.n3647 4.5005
R19226 DVSS.n3666 DVSS.n3649 4.5005
R19227 DVSS.n4848 DVSS.n3649 4.5005
R19228 DVSS.n4850 DVSS.n3648 4.5005
R19229 DVSS.n3648 DVSS.n3647 4.5005
R19230 DVSS.n3666 DVSS.n3648 4.5005
R19231 DVSS.n4848 DVSS.n3648 4.5005
R19232 DVSS.n3447 DVSS.n3436 4.5005
R19233 DVSS.n5272 DVSS.n3447 4.5005
R19234 DVSS.n3447 DVSS.n3440 4.5005
R19235 DVSS.n5270 DVSS.n3447 4.5005
R19236 DVSS.n3445 DVSS.n3436 4.5005
R19237 DVSS.n5272 DVSS.n3445 4.5005
R19238 DVSS.n3445 DVSS.n3440 4.5005
R19239 DVSS.n5270 DVSS.n3445 4.5005
R19240 DVSS.n3448 DVSS.n3436 4.5005
R19241 DVSS.n5272 DVSS.n3448 4.5005
R19242 DVSS.n3448 DVSS.n3440 4.5005
R19243 DVSS.n5270 DVSS.n3448 4.5005
R19244 DVSS.n3444 DVSS.n3436 4.5005
R19245 DVSS.n5272 DVSS.n3444 4.5005
R19246 DVSS.n3444 DVSS.n3440 4.5005
R19247 DVSS.n5270 DVSS.n3444 4.5005
R19248 DVSS.n3450 DVSS.n3436 4.5005
R19249 DVSS.n5272 DVSS.n3450 4.5005
R19250 DVSS.n5270 DVSS.n3450 4.5005
R19251 DVSS.n5272 DVSS.n3443 4.5005
R19252 DVSS.n5270 DVSS.n3443 4.5005
R19253 DVSS.n5272 DVSS.n3453 4.5005
R19254 DVSS.n5270 DVSS.n3453 4.5005
R19255 DVSS.n5272 DVSS.n3442 4.5005
R19256 DVSS.n5270 DVSS.n3442 4.5005
R19257 DVSS.n5272 DVSS.n3456 4.5005
R19258 DVSS.n5270 DVSS.n3456 4.5005
R19259 DVSS.n5272 DVSS.n3441 4.5005
R19260 DVSS.n5270 DVSS.n3441 4.5005
R19261 DVSS.n5272 DVSS.n5271 4.5005
R19262 DVSS.n5271 DVSS.n3440 4.5005
R19263 DVSS.n5271 DVSS.n5270 4.5005
R19264 DVSS.n5393 DVSS.n3333 4.5005
R19265 DVSS.n3333 DVSS.n3325 4.5005
R19266 DVSS.n3333 DVSS.n3326 4.5005
R19267 DVSS.n3335 DVSS.n3325 4.5005
R19268 DVSS.n3335 DVSS.n3326 4.5005
R19269 DVSS.n3339 DVSS.n3325 4.5005
R19270 DVSS.n3339 DVSS.n3326 4.5005
R19271 DVSS.n3341 DVSS.n3325 4.5005
R19272 DVSS.n3341 DVSS.n3326 4.5005
R19273 DVSS.n3338 DVSS.n3325 4.5005
R19274 DVSS.n3338 DVSS.n3326 4.5005
R19275 DVSS.n5393 DVSS.n3331 4.5005
R19276 DVSS.n3331 DVSS.n3325 4.5005
R19277 DVSS.n3331 DVSS.n3326 4.5005
R19278 DVSS.n3343 DVSS.n3326 4.5005
R19279 DVSS.n3343 DVSS.n3327 4.5005
R19280 DVSS.n3343 DVSS.n3325 4.5005
R19281 DVSS.n5393 DVSS.n3343 4.5005
R19282 DVSS.n3330 DVSS.n3326 4.5005
R19283 DVSS.n3330 DVSS.n3327 4.5005
R19284 DVSS.n3330 DVSS.n3325 4.5005
R19285 DVSS.n5393 DVSS.n3330 4.5005
R19286 DVSS.n5392 DVSS.n3326 4.5005
R19287 DVSS.n5392 DVSS.n3327 4.5005
R19288 DVSS.n5392 DVSS.n3325 4.5005
R19289 DVSS.n5393 DVSS.n5392 4.5005
R19290 DVSS.n3329 DVSS.n3326 4.5005
R19291 DVSS.n3329 DVSS.n3327 4.5005
R19292 DVSS.n3329 DVSS.n3325 4.5005
R19293 DVSS.n5393 DVSS.n3329 4.5005
R19294 DVSS.n5394 DVSS.n3326 4.5005
R19295 DVSS.n5394 DVSS.n3327 4.5005
R19296 DVSS.n5394 DVSS.n3325 4.5005
R19297 DVSS.n5394 DVSS.n5393 4.5005
R19298 DVSS.n7847 DVSS.n7729 4.5005
R19299 DVSS.n7847 DVSS.n7730 4.5005
R19300 DVSS.n7847 DVSS.n7846 4.5005
R19301 DVSS.n7736 DVSS.n7730 4.5005
R19302 DVSS.n7846 DVSS.n7736 4.5005
R19303 DVSS.n7739 DVSS.n7730 4.5005
R19304 DVSS.n7846 DVSS.n7739 4.5005
R19305 DVSS.n7735 DVSS.n7730 4.5005
R19306 DVSS.n7846 DVSS.n7735 4.5005
R19307 DVSS.n7741 DVSS.n7730 4.5005
R19308 DVSS.n7846 DVSS.n7741 4.5005
R19309 DVSS.n7734 DVSS.n7730 4.5005
R19310 DVSS.n7846 DVSS.n7734 4.5005
R19311 DVSS.n7743 DVSS.n7730 4.5005
R19312 DVSS.n7846 DVSS.n7743 4.5005
R19313 DVSS.n7733 DVSS.n7730 4.5005
R19314 DVSS.n7846 DVSS.n7733 4.5005
R19315 DVSS.n7745 DVSS.n7730 4.5005
R19316 DVSS.n7846 DVSS.n7745 4.5005
R19317 DVSS.n7732 DVSS.n7730 4.5005
R19318 DVSS.n7846 DVSS.n7732 4.5005
R19319 DVSS.n7845 DVSS.n7730 4.5005
R19320 DVSS.n7845 DVSS.n7844 4.5005
R19321 DVSS.n7846 DVSS.n7845 4.5005
R19322 DVSS.n8341 DVSS.n1426 4.5005
R19323 DVSS.n8341 DVSS.n1427 4.5005
R19324 DVSS.n8348 DVSS.n8341 4.5005
R19325 DVSS.n1435 DVSS.n1427 4.5005
R19326 DVSS.n8348 DVSS.n1435 4.5005
R19327 DVSS.n8344 DVSS.n1427 4.5005
R19328 DVSS.n8348 DVSS.n8344 4.5005
R19329 DVSS.n1434 DVSS.n1427 4.5005
R19330 DVSS.n8348 DVSS.n1434 4.5005
R19331 DVSS.n1427 DVSS.n1424 4.5005
R19332 DVSS.n1425 DVSS.n1424 4.5005
R19333 DVSS.n8348 DVSS.n1424 4.5005
R19334 DVSS.n8349 DVSS.n1426 4.5005
R19335 DVSS.n8349 DVSS.n1427 4.5005
R19336 DVSS.n8349 DVSS.n1425 4.5005
R19337 DVSS.n8349 DVSS.n8348 4.5005
R19338 DVSS.n8348 DVSS.n1422 4.5005
R19339 DVSS.n1425 DVSS.n1422 4.5005
R19340 DVSS.n1426 DVSS.n1422 4.5005
R19341 DVSS.n1432 DVSS.n1426 4.5005
R19342 DVSS.n8348 DVSS.n1432 4.5005
R19343 DVSS.n8347 DVSS.n1427 4.5005
R19344 DVSS.n8348 DVSS.n8347 4.5005
R19345 DVSS.n1430 DVSS.n1427 4.5005
R19346 DVSS.n8348 DVSS.n1430 4.5005
R19347 DVSS.n1426 DVSS.n1135 4.5005
R19348 DVSS.n1427 DVSS.n1135 4.5005
R19349 DVSS.n8348 DVSS.n1135 4.5005
R19350 DVSS.n8333 DVSS.n1443 4.5005
R19351 DVSS.n8333 DVSS.n1441 4.5005
R19352 DVSS.n7095 DVSS.n7093 4.5005
R19353 DVSS.n7095 DVSS.n7094 4.5005
R19354 DVSS.n7096 DVSS.n7095 4.5005
R19355 DVSS.n7097 DVSS.n7096 4.5005
R19356 DVSS.n8098 DVSS.n8097 4.5005
R19357 DVSS.n7865 DVSS.n7864 4.5005
R19358 DVSS.n7863 DVSS.n2074 4.5005
R19359 DVSS.n7869 DVSS.n2075 4.5005
R19360 DVSS.n7872 DVSS.n7870 4.5005
R19361 DVSS.n7875 DVSS.n7873 4.5005
R19362 DVSS.n7878 DVSS.n7876 4.5005
R19363 DVSS.n7881 DVSS.n7879 4.5005
R19364 DVSS.n7883 DVSS.n7882 4.5005
R19365 DVSS.n7887 DVSS.n7884 4.5005
R19366 DVSS.n7890 DVSS.n7888 4.5005
R19367 DVSS.n7893 DVSS.n7891 4.5005
R19368 DVSS.n7895 DVSS.n2073 4.5005
R19369 DVSS.n7899 DVSS.n7898 4.5005
R19370 DVSS.n2059 DVSS.n2058 4.5005
R19371 DVSS.n7933 DVSS.n7903 4.5005
R19372 DVSS.n7932 DVSS.n7904 4.5005
R19373 DVSS.n7931 DVSS.n7905 4.5005
R19374 DVSS.n7908 DVSS.n7906 4.5005
R19375 DVSS.n7927 DVSS.n7909 4.5005
R19376 DVSS.n7926 DVSS.n7910 4.5005
R19377 DVSS.n7925 DVSS.n7911 4.5005
R19378 DVSS.n7914 DVSS.n7912 4.5005
R19379 DVSS.n7921 DVSS.n7915 4.5005
R19380 DVSS.n7920 DVSS.n7916 4.5005
R19381 DVSS.n7919 DVSS.n7917 4.5005
R19382 DVSS.n1872 DVSS.n1871 4.5005
R19383 DVSS.n7862 DVSS.n2077 4.5005
R19384 DVSS.n7328 DVSS.n7327 4.5005
R19385 DVSS.n7275 DVSS.n7274 4.5005
R19386 DVSS.n7276 DVSS.n2649 4.5005
R19387 DVSS.n7278 DVSS.n7277 4.5005
R19388 DVSS.n2647 DVSS.n2646 4.5005
R19389 DVSS.n7283 DVSS.n7282 4.5005
R19390 DVSS.n7284 DVSS.n2645 4.5005
R19391 DVSS.n7286 DVSS.n7285 4.5005
R19392 DVSS.n2643 DVSS.n2642 4.5005
R19393 DVSS.n7291 DVSS.n7290 4.5005
R19394 DVSS.n7292 DVSS.n2641 4.5005
R19395 DVSS.n7294 DVSS.n7293 4.5005
R19396 DVSS.n2638 DVSS.n2637 4.5005
R19397 DVSS.n7299 DVSS.n7298 4.5005
R19398 DVSS.n7300 DVSS.n2636 4.5005
R19399 DVSS.n7302 DVSS.n7301 4.5005
R19400 DVSS.n2634 DVSS.n2633 4.5005
R19401 DVSS.n7307 DVSS.n7306 4.5005
R19402 DVSS.n7308 DVSS.n2632 4.5005
R19403 DVSS.n7310 DVSS.n7309 4.5005
R19404 DVSS.n2630 DVSS.n2629 4.5005
R19405 DVSS.n7315 DVSS.n7314 4.5005
R19406 DVSS.n7316 DVSS.n2628 4.5005
R19407 DVSS.n7318 DVSS.n7317 4.5005
R19408 DVSS.n2626 DVSS.n2625 4.5005
R19409 DVSS.n7323 DVSS.n7322 4.5005
R19410 DVSS.n7324 DVSS.n2623 4.5005
R19411 DVSS.n2651 DVSS.n2650 4.5005
R19412 DVSS.n2701 DVSS.n2700 4.5005
R19413 DVSS.n5550 DVSS.n5549 4.5005
R19414 DVSS.n5625 DVSS.n5551 4.5005
R19415 DVSS.n5624 DVSS.n5552 4.5005
R19416 DVSS.n5622 DVSS.n5553 4.5005
R19417 DVSS.n5620 DVSS.n5554 4.5005
R19418 DVSS.n5618 DVSS.n5555 4.5005
R19419 DVSS.n5616 DVSS.n5556 4.5005
R19420 DVSS.n5614 DVSS.n5557 4.5005
R19421 DVSS.n5611 DVSS.n5558 4.5005
R19422 DVSS.n5610 DVSS.n5559 4.5005
R19423 DVSS.n5608 DVSS.n5560 4.5005
R19424 DVSS.n5606 DVSS.n5561 4.5005
R19425 DVSS.n5604 DVSS.n5562 4.5005
R19426 DVSS.n5601 DVSS.n5563 4.5005
R19427 DVSS.n5599 DVSS.n5564 4.5005
R19428 DVSS.n5596 DVSS.n5565 4.5005
R19429 DVSS.n5595 DVSS.n5566 4.5005
R19430 DVSS.n5593 DVSS.n5567 4.5005
R19431 DVSS.n5591 DVSS.n5568 4.5005
R19432 DVSS.n5589 DVSS.n5569 4.5005
R19433 DVSS.n5587 DVSS.n5570 4.5005
R19434 DVSS.n5585 DVSS.n5571 4.5005
R19435 DVSS.n5583 DVSS.n5572 4.5005
R19436 DVSS.n5580 DVSS.n5573 4.5005
R19437 DVSS.n5579 DVSS.n5574 4.5005
R19438 DVSS.n5577 DVSS.n5575 4.5005
R19439 DVSS.n5630 DVSS.n5629 4.5005
R19440 DVSS.n5640 DVSS.n5639 4.5005
R19441 DVSS.n5407 DVSS.n5406 4.5005
R19442 DVSS.n5479 DVSS.n5409 4.5005
R19443 DVSS.n5478 DVSS.n5410 4.5005
R19444 DVSS.n5477 DVSS.n5411 4.5005
R19445 DVSS.n5414 DVSS.n5412 4.5005
R19446 DVSS.n5473 DVSS.n5415 4.5005
R19447 DVSS.n5472 DVSS.n5416 4.5005
R19448 DVSS.n5471 DVSS.n5417 4.5005
R19449 DVSS.n5420 DVSS.n5418 4.5005
R19450 DVSS.n5467 DVSS.n5421 4.5005
R19451 DVSS.n5466 DVSS.n5422 4.5005
R19452 DVSS.n5465 DVSS.n5423 4.5005
R19453 DVSS.n5427 DVSS.n5424 4.5005
R19454 DVSS.n5461 DVSS.n5428 4.5005
R19455 DVSS.n5460 DVSS.n5429 4.5005
R19456 DVSS.n5459 DVSS.n5430 4.5005
R19457 DVSS.n5433 DVSS.n5431 4.5005
R19458 DVSS.n5455 DVSS.n5434 4.5005
R19459 DVSS.n5454 DVSS.n5435 4.5005
R19460 DVSS.n5453 DVSS.n5436 4.5005
R19461 DVSS.n5439 DVSS.n5437 4.5005
R19462 DVSS.n5449 DVSS.n5440 4.5005
R19463 DVSS.n5448 DVSS.n5441 4.5005
R19464 DVSS.n5447 DVSS.n5442 4.5005
R19465 DVSS.n5444 DVSS.n5443 4.5005
R19466 DVSS.n3285 DVSS.n3283 4.5005
R19467 DVSS.n5484 DVSS.n5483 4.5005
R19468 DVSS.n5487 DVSS.n3229 4.5005
R19469 DVSS.n5737 DVSS.n3191 4.5005
R19470 DVSS.n5736 DVSS.n3192 4.5005
R19471 DVSS.n3195 DVSS.n3193 4.5005
R19472 DVSS.n5732 DVSS.n3196 4.5005
R19473 DVSS.n5731 DVSS.n3197 4.5005
R19474 DVSS.n5730 DVSS.n3198 4.5005
R19475 DVSS.n3201 DVSS.n3199 4.5005
R19476 DVSS.n5726 DVSS.n3202 4.5005
R19477 DVSS.n5725 DVSS.n3203 4.5005
R19478 DVSS.n5724 DVSS.n3204 4.5005
R19479 DVSS.n3207 DVSS.n3205 4.5005
R19480 DVSS.n5720 DVSS.n3208 4.5005
R19481 DVSS.n5719 DVSS.n3209 4.5005
R19482 DVSS.n5717 DVSS.n3210 4.5005
R19483 DVSS.n3213 DVSS.n3211 4.5005
R19484 DVSS.n5713 DVSS.n3214 4.5005
R19485 DVSS.n5712 DVSS.n3215 4.5005
R19486 DVSS.n5711 DVSS.n3216 4.5005
R19487 DVSS.n3219 DVSS.n3217 4.5005
R19488 DVSS.n5707 DVSS.n3220 4.5005
R19489 DVSS.n5706 DVSS.n3221 4.5005
R19490 DVSS.n5705 DVSS.n3222 4.5005
R19491 DVSS.n3225 DVSS.n3223 4.5005
R19492 DVSS.n5701 DVSS.n3226 4.5005
R19493 DVSS.n5700 DVSS.n3227 4.5005
R19494 DVSS.n5699 DVSS.n3228 4.5005
R19495 DVSS.n5738 DVSS.n3190 4.5005
R19496 DVSS.n5199 DVSS.n5198 4.5005
R19497 DVSS.n3990 DVSS.n3984 4.5005
R19498 DVSS.n3988 DVSS.n3985 4.5005
R19499 DVSS.n3987 DVSS.n3986 4.5005
R19500 DVSS.n3487 DVSS.n3485 4.5005
R19501 DVSS.n5235 DVSS.n5234 4.5005
R19502 DVSS.n3488 DVSS.n3486 4.5005
R19503 DVSS.n5230 DVSS.n3491 4.5005
R19504 DVSS.n5229 DVSS.n3492 4.5005
R19505 DVSS.n5228 DVSS.n3493 4.5005
R19506 DVSS.n3496 DVSS.n3494 4.5005
R19507 DVSS.n5224 DVSS.n3497 4.5005
R19508 DVSS.n5223 DVSS.n3498 4.5005
R19509 DVSS.n5222 DVSS.n3499 4.5005
R19510 DVSS.n5219 DVSS.n3502 4.5005
R19511 DVSS.n5218 DVSS.n3503 4.5005
R19512 DVSS.n5217 DVSS.n3504 4.5005
R19513 DVSS.n3507 DVSS.n3505 4.5005
R19514 DVSS.n5213 DVSS.n3508 4.5005
R19515 DVSS.n5212 DVSS.n3509 4.5005
R19516 DVSS.n5211 DVSS.n3510 4.5005
R19517 DVSS.n3513 DVSS.n3511 4.5005
R19518 DVSS.n5207 DVSS.n3514 4.5005
R19519 DVSS.n5206 DVSS.n3515 4.5005
R19520 DVSS.n5205 DVSS.n3516 4.5005
R19521 DVSS.n5203 DVSS.n3517 4.5005
R19522 DVSS.n5201 DVSS.n3518 4.5005
R19523 DVSS.n3991 DVSS.n3983 4.5005
R19524 DVSS.n4089 DVSS.n3561 4.5005
R19525 DVSS.n4040 DVSS.n4039 4.5005
R19526 DVSS.n4041 DVSS.n4035 4.5005
R19527 DVSS.n4043 DVSS.n4042 4.5005
R19528 DVSS.n4033 DVSS.n4032 4.5005
R19529 DVSS.n4048 DVSS.n4047 4.5005
R19530 DVSS.n4049 DVSS.n4031 4.5005
R19531 DVSS.n4051 DVSS.n4050 4.5005
R19532 DVSS.n4029 DVSS.n4028 4.5005
R19533 DVSS.n4056 DVSS.n4055 4.5005
R19534 DVSS.n4057 DVSS.n4027 4.5005
R19535 DVSS.n4059 DVSS.n4058 4.5005
R19536 DVSS.n4025 DVSS.n4024 4.5005
R19537 DVSS.n4064 DVSS.n4063 4.5005
R19538 DVSS.n4066 DVSS.n4065 4.5005
R19539 DVSS.n4067 DVSS.n4021 4.5005
R19540 DVSS.n4071 DVSS.n4070 4.5005
R19541 DVSS.n4072 DVSS.n4020 4.5005
R19542 DVSS.n4074 DVSS.n4073 4.5005
R19543 DVSS.n4018 DVSS.n4017 4.5005
R19544 DVSS.n4079 DVSS.n4078 4.5005
R19545 DVSS.n4080 DVSS.n4016 4.5005
R19546 DVSS.n4082 DVSS.n4081 4.5005
R19547 DVSS.n4014 DVSS.n4013 4.5005
R19548 DVSS.n4087 DVSS.n4086 4.5005
R19549 DVSS.n4088 DVSS.n4012 4.5005
R19550 DVSS.n4091 DVSS.n4090 4.5005
R19551 DVSS.n4037 DVSS.n4036 4.5005
R19552 DVSS.n4813 DVSS.n4812 4.5005
R19553 DVSS.n4700 DVSS.n4625 4.5005
R19554 DVSS.n4698 DVSS.n4626 4.5005
R19555 DVSS.n4696 DVSS.n4627 4.5005
R19556 DVSS.n4694 DVSS.n4628 4.5005
R19557 DVSS.n4631 DVSS.n4629 4.5005
R19558 DVSS.n4690 DVSS.n4632 4.5005
R19559 DVSS.n4689 DVSS.n4633 4.5005
R19560 DVSS.n4688 DVSS.n4634 4.5005
R19561 DVSS.n4637 DVSS.n4635 4.5005
R19562 DVSS.n4684 DVSS.n4638 4.5005
R19563 DVSS.n4683 DVSS.n4639 4.5005
R19564 DVSS.n4682 DVSS.n4640 4.5005
R19565 DVSS.n4644 DVSS.n4641 4.5005
R19566 DVSS.n4678 DVSS.n4645 4.5005
R19567 DVSS.n4677 DVSS.n4646 4.5005
R19568 DVSS.n4676 DVSS.n4647 4.5005
R19569 DVSS.n4650 DVSS.n4648 4.5005
R19570 DVSS.n4672 DVSS.n4651 4.5005
R19571 DVSS.n4671 DVSS.n4652 4.5005
R19572 DVSS.n4670 DVSS.n4653 4.5005
R19573 DVSS.n4655 DVSS.n4654 4.5005
R19574 DVSS.n4666 DVSS.n4656 4.5005
R19575 DVSS.n4665 DVSS.n4657 4.5005
R19576 DVSS.n4663 DVSS.n4658 4.5005
R19577 DVSS.n4661 DVSS.n4659 4.5005
R19578 DVSS.n3687 DVSS.n3686 4.5005
R19579 DVSS.n4703 DVSS.n4702 4.5005
R19580 DVSS.n4817 DVSS.n3684 4.5005
R19581 DVSS.n3684 DVSS.n3677 4.5005
R19582 DVSS.n3684 DVSS.n3678 4.5005
R19583 DVSS.n4817 DVSS.n3682 4.5005
R19584 DVSS.n3682 DVSS.n3677 4.5005
R19585 DVSS.n3682 DVSS.n3678 4.5005
R19586 DVSS.n4817 DVSS.n3685 4.5005
R19587 DVSS.n3685 DVSS.n3677 4.5005
R19588 DVSS.n3685 DVSS.n3678 4.5005
R19589 DVSS.n3681 DVSS.n3678 4.5005
R19590 DVSS.n3681 DVSS.n3677 4.5005
R19591 DVSS.n4817 DVSS.n3681 4.5005
R19592 DVSS.n4814 DVSS.n3678 4.5005
R19593 DVSS.n4814 DVSS.n3677 4.5005
R19594 DVSS.n4817 DVSS.n4814 4.5005
R19595 DVSS.n3680 DVSS.n3678 4.5005
R19596 DVSS.n4817 DVSS.n3680 4.5005
R19597 DVSS.n4816 DVSS.n3678 4.5005
R19598 DVSS.n4817 DVSS.n4816 4.5005
R19599 DVSS.n3678 DVSS.n3672 4.5005
R19600 DVSS.n3677 DVSS.n3672 4.5005
R19601 DVSS.n4817 DVSS.n3672 4.5005
R19602 DVSS.n3678 DVSS.n3674 4.5005
R19603 DVSS.n3677 DVSS.n3674 4.5005
R19604 DVSS.n4817 DVSS.n3674 4.5005
R19605 DVSS.n3678 DVSS.n3676 4.5005
R19606 DVSS.n3677 DVSS.n3676 4.5005
R19607 DVSS.n4817 DVSS.n3676 4.5005
R19608 DVSS.n4818 DVSS.n3678 4.5005
R19609 DVSS.n4818 DVSS.n3677 4.5005
R19610 DVSS.n4818 DVSS.n4817 4.5005
R19611 DVSS.n3481 DVSS.n3470 4.5005
R19612 DVSS.n5237 DVSS.n3481 4.5005
R19613 DVSS.n3481 DVSS.n3474 4.5005
R19614 DVSS.n3479 DVSS.n3470 4.5005
R19615 DVSS.n5237 DVSS.n3479 4.5005
R19616 DVSS.n3479 DVSS.n3474 4.5005
R19617 DVSS.n3482 DVSS.n3470 4.5005
R19618 DVSS.n5237 DVSS.n3482 4.5005
R19619 DVSS.n3482 DVSS.n3474 4.5005
R19620 DVSS.n3478 DVSS.n3470 4.5005
R19621 DVSS.n5237 DVSS.n3478 4.5005
R19622 DVSS.n3478 DVSS.n3474 4.5005
R19623 DVSS.n4999 DVSS.n3470 4.5005
R19624 DVSS.n4999 DVSS.n3474 4.5005
R19625 DVSS.n3982 DVSS.n3470 4.5005
R19626 DVSS.n3982 DVSS.n3474 4.5005
R19627 DVSS.n3483 DVSS.n3474 4.5005
R19628 DVSS.n5237 DVSS.n3483 4.5005
R19629 DVSS.n3483 DVSS.n3470 4.5005
R19630 DVSS.n3476 DVSS.n3474 4.5005
R19631 DVSS.n5237 DVSS.n3476 4.5005
R19632 DVSS.n3476 DVSS.n3470 4.5005
R19633 DVSS.n3484 DVSS.n3470 4.5005
R19634 DVSS.n5237 DVSS.n3484 4.5005
R19635 DVSS.n3484 DVSS.n3474 4.5005
R19636 DVSS.n3475 DVSS.n3470 4.5005
R19637 DVSS.n5237 DVSS.n3475 4.5005
R19638 DVSS.n3475 DVSS.n3474 4.5005
R19639 DVSS.n5236 DVSS.n3470 4.5005
R19640 DVSS.n5237 DVSS.n5236 4.5005
R19641 DVSS.n5236 DVSS.n3474 4.5005
R19642 DVSS.n5196 DVSS.n5017 4.5005
R19643 DVSS.n5194 DVSS.n5017 4.5005
R19644 DVSS.n5017 DVSS.n5010 4.5005
R19645 DVSS.n5196 DVSS.n5015 4.5005
R19646 DVSS.n5194 DVSS.n5015 4.5005
R19647 DVSS.n5015 DVSS.n5010 4.5005
R19648 DVSS.n5196 DVSS.n5018 4.5005
R19649 DVSS.n5194 DVSS.n5018 4.5005
R19650 DVSS.n5018 DVSS.n5010 4.5005
R19651 DVSS.n5010 DVSS.n5008 4.5005
R19652 DVSS.n5194 DVSS.n5008 4.5005
R19653 DVSS.n5196 DVSS.n5008 4.5005
R19654 DVSS.n5197 DVSS.n5010 4.5005
R19655 DVSS.n5197 DVSS.n5196 4.5005
R19656 DVSS.n5014 DVSS.n5010 4.5005
R19657 DVSS.n5196 DVSS.n5014 4.5005
R19658 DVSS.n5196 DVSS.n5019 4.5005
R19659 DVSS.n5194 DVSS.n5019 4.5005
R19660 DVSS.n5019 DVSS.n5010 4.5005
R19661 DVSS.n5196 DVSS.n5013 4.5005
R19662 DVSS.n5194 DVSS.n5013 4.5005
R19663 DVSS.n5013 DVSS.n5010 4.5005
R19664 DVSS.n5196 DVSS.n5020 4.5005
R19665 DVSS.n5194 DVSS.n5020 4.5005
R19666 DVSS.n5020 DVSS.n5010 4.5005
R19667 DVSS.n5196 DVSS.n5012 4.5005
R19668 DVSS.n5194 DVSS.n5012 4.5005
R19669 DVSS.n5012 DVSS.n5010 4.5005
R19670 DVSS.n5196 DVSS.n5195 4.5005
R19671 DVSS.n5195 DVSS.n5194 4.5005
R19672 DVSS.n5195 DVSS.n5010 4.5005
R19673 DVSS.n7901 DVSS.n2069 4.5005
R19674 DVSS.n2069 DVSS.n2060 4.5005
R19675 DVSS.n2069 DVSS.n2061 4.5005
R19676 DVSS.n7901 DVSS.n2067 4.5005
R19677 DVSS.n2067 DVSS.n2060 4.5005
R19678 DVSS.n2067 DVSS.n2061 4.5005
R19679 DVSS.n2070 DVSS.n2061 4.5005
R19680 DVSS.n2070 DVSS.n2060 4.5005
R19681 DVSS.n7901 DVSS.n2070 4.5005
R19682 DVSS.n2066 DVSS.n2061 4.5005
R19683 DVSS.n2066 DVSS.n2060 4.5005
R19684 DVSS.n7901 DVSS.n2066 4.5005
R19685 DVSS.n2071 DVSS.n2061 4.5005
R19686 DVSS.n2071 DVSS.n2060 4.5005
R19687 DVSS.n7901 DVSS.n2071 4.5005
R19688 DVSS.n2065 DVSS.n2061 4.5005
R19689 DVSS.n2065 DVSS.n2060 4.5005
R19690 DVSS.n7901 DVSS.n2065 4.5005
R19691 DVSS.n7901 DVSS.n2072 4.5005
R19692 DVSS.n2072 DVSS.n2060 4.5005
R19693 DVSS.n2072 DVSS.n2061 4.5005
R19694 DVSS.n7901 DVSS.n2064 4.5005
R19695 DVSS.n2064 DVSS.n2060 4.5005
R19696 DVSS.n2064 DVSS.n2061 4.5005
R19697 DVSS.n7901 DVSS.n7900 4.5005
R19698 DVSS.n7900 DVSS.n2060 4.5005
R19699 DVSS.n7900 DVSS.n2061 4.5005
R19700 DVSS.n2063 DVSS.n2061 4.5005
R19701 DVSS.n2063 DVSS.n2060 4.5005
R19702 DVSS.n7901 DVSS.n2063 4.5005
R19703 DVSS.n7902 DVSS.n2061 4.5005
R19704 DVSS.n7902 DVSS.n2060 4.5005
R19705 DVSS.n7902 DVSS.n7901 4.5005
R19706 DVSS.n8388 DVSS.n1415 4.5005
R19707 DVSS.n1415 DVSS.n1398 4.5005
R19708 DVSS.n1412 DVSS.n1398 4.5005
R19709 DVSS.n1411 DVSS.n1398 4.5005
R19710 DVSS.n8389 DVSS.n1398 4.5005
R19711 DVSS.n8392 DVSS.n8391 4.5005
R19712 DVSS.n8391 DVSS.n1398 4.5005
R19713 DVSS.n8388 DVSS.n1401 4.5005
R19714 DVSS.n8392 DVSS.n1401 4.5005
R19715 DVSS.n1401 DVSS.n1398 4.5005
R19716 DVSS.n8387 DVSS.n1398 4.5005
R19717 DVSS.n8388 DVSS.n8387 4.5005
R19718 DVSS.n1409 DVSS.n1398 4.5005
R19719 DVSS.n1408 DVSS.n1398 4.5005
R19720 DVSS.n1406 DVSS.n1398 4.5005
R19721 DVSS.n8392 DVSS.n1143 4.5005
R19722 DVSS.n1398 DVSS.n1143 4.5005
R19723 DVSS.n8273 DVSS.n8263 4.5005
R19724 DVSS.n8266 DVSS.n8263 4.5005
R19725 DVSS.n8271 DVSS.n8263 4.5005
R19726 DVSS.n8261 DVSS.n1471 4.5005
R19727 DVSS.n8266 DVSS.n1465 4.5005
R19728 DVSS.n8271 DVSS.n1465 4.5005
R19729 DVSS.n8279 DVSS.n8278 4.5005
R19730 DVSS.n8273 DVSS.n8272 4.5005
R19731 DVSS.n8272 DVSS.n8271 4.5005
R19732 DVSS.n8282 DVSS.n1501 4.5005
R19733 DVSS.n8282 DVSS.n8281 4.5005
R19734 DVSS.n8326 DVSS.n1446 4.5005
R19735 DVSS.n8326 DVSS.n8325 4.5005
R19736 DVSS.n8327 DVSS.n8326 4.5005
R19737 DVSS.n8281 DVSS.n8280 4.5005
R19738 DVSS.n8325 DVSS.n1449 4.5005
R19739 DVSS.n8327 DVSS.n1449 4.5005
R19740 DVSS.n8281 DVSS.n1499 4.5005
R19741 DVSS.n8328 DVSS.n1446 4.5005
R19742 DVSS.n8328 DVSS.n8327 4.5005
R19743 DVSS.n8304 DVSS.n1469 4.5005
R19744 DVSS.n8307 DVSS.n1469 4.5005
R19745 DVSS.n8308 DVSS.n1463 4.5005
R19746 DVSS.n8311 DVSS.n1463 4.5005
R19747 DVSS.n8314 DVSS.n1463 4.5005
R19748 DVSS.n8307 DVSS.n1467 4.5005
R19749 DVSS.n8311 DVSS.n1461 4.5005
R19750 DVSS.n8314 DVSS.n1461 4.5005
R19751 DVSS.n8307 DVSS.n8306 4.5005
R19752 DVSS.n8313 DVSS.n8308 4.5005
R19753 DVSS.n8314 DVSS.n8313 4.5005
R19754 DVSS.n8218 DVSS.n1528 4.5005
R19755 DVSS.n8214 DVSS.n8212 4.5005
R19756 DVSS.n8212 DVSS.n1458 4.5005
R19757 DVSS.n8216 DVSS.n1458 4.5005
R19758 DVSS.n8217 DVSS.n8216 4.5005
R19759 DVSS.n8219 DVSS.n8218 4.5005
R19760 DVSS.n8219 DVSS.n1526 4.5005
R19761 DVSS.n8220 DVSS.n8219 4.5005
R19762 DVSS.n7143 DVSS.n1523 4.5005
R19763 DVSS.n1523 DVSS.n1522 4.5005
R19764 DVSS.n8222 DVSS.n1523 4.5005
R19765 DVSS.n8223 DVSS.n8222 4.5005
R19766 DVSS.n7084 DVSS.n7083 4.5005
R19767 DVSS.n8288 DVSS.n1494 4.5005
R19768 DVSS.n8288 DVSS.n8287 4.5005
R19769 DVSS.n8287 DVSS.n1497 4.5005
R19770 DVSS.n8252 DVSS.n1509 4.5005
R19771 DVSS.n8255 DVSS.n1509 4.5005
R19772 DVSS.n8255 DVSS.n1507 4.5005
R19773 DVSS.n8229 DVSS.n8228 4.5005
R19774 DVSS.n8229 DVSS.n1472 4.5005
R19775 DVSS.n8224 DVSS.n1472 4.5005
R19776 DVSS.n1518 DVSS.n1472 4.5005
R19777 DVSS.n8255 DVSS.n8254 4.5005
R19778 DVSS.n8287 DVSS.n1492 4.5005
R19779 DVSS.n7110 DVSS.n7084 4.5005
R19780 DVSS.n7110 DVSS.n7081 4.5005
R19781 DVSS.n7111 DVSS.n7110 4.5005
R19782 DVSS.n7248 DVSS.n6648 4.5005
R19783 DVSS.n8097 DVSS.n8096 4.5005
R19784 DVSS.n1873 DVSS.n1872 4.5005
R19785 DVSS.n7919 DVSS.n7918 4.5005
R19786 DVSS.n7920 DVSS.n7913 4.5005
R19787 DVSS.n7922 DVSS.n7921 4.5005
R19788 DVSS.n7923 DVSS.n7912 4.5005
R19789 DVSS.n7925 DVSS.n7924 4.5005
R19790 DVSS.n7926 DVSS.n7907 4.5005
R19791 DVSS.n7928 DVSS.n7927 4.5005
R19792 DVSS.n7929 DVSS.n7906 4.5005
R19793 DVSS.n7931 DVSS.n7930 4.5005
R19794 DVSS.n7932 DVSS.n2057 4.5005
R19795 DVSS.n7934 DVSS.n7933 4.5005
R19796 DVSS.n2058 DVSS.n2056 4.5005
R19797 DVSS.n7898 DVSS.n7897 4.5005
R19798 DVSS.n7895 DVSS.n7894 4.5005
R19799 DVSS.n7893 DVSS.n7892 4.5005
R19800 DVSS.n7890 DVSS.n7889 4.5005
R19801 DVSS.n7887 DVSS.n7886 4.5005
R19802 DVSS.n7885 DVSS.n7882 4.5005
R19803 DVSS.n7881 DVSS.n7880 4.5005
R19804 DVSS.n7878 DVSS.n7877 4.5005
R19805 DVSS.n7875 DVSS.n7874 4.5005
R19806 DVSS.n7872 DVSS.n7871 4.5005
R19807 DVSS.n7869 DVSS.n7868 4.5005
R19808 DVSS.n7867 DVSS.n2074 4.5005
R19809 DVSS.n7866 DVSS.n7865 4.5005
R19810 DVSS.n2077 DVSS.n2076 4.5005
R19811 DVSS.n7329 DVSS.n7328 4.5005
R19812 DVSS.n2623 DVSS.n2622 4.5005
R19813 DVSS.n7322 DVSS.n7321 4.5005
R19814 DVSS.n7320 DVSS.n2626 4.5005
R19815 DVSS.n7319 DVSS.n7318 4.5005
R19816 DVSS.n2628 DVSS.n2627 4.5005
R19817 DVSS.n7314 DVSS.n7313 4.5005
R19818 DVSS.n7312 DVSS.n2630 4.5005
R19819 DVSS.n7311 DVSS.n7310 4.5005
R19820 DVSS.n2632 DVSS.n2631 4.5005
R19821 DVSS.n7306 DVSS.n7305 4.5005
R19822 DVSS.n7304 DVSS.n2634 4.5005
R19823 DVSS.n7303 DVSS.n7302 4.5005
R19824 DVSS.n2636 DVSS.n2635 4.5005
R19825 DVSS.n7298 DVSS.n7297 4.5005
R19826 DVSS.n7296 DVSS.n2638 4.5005
R19827 DVSS.n7295 DVSS.n7294 4.5005
R19828 DVSS.n2641 DVSS.n2640 4.5005
R19829 DVSS.n7290 DVSS.n7289 4.5005
R19830 DVSS.n7288 DVSS.n2643 4.5005
R19831 DVSS.n7287 DVSS.n7286 4.5005
R19832 DVSS.n2645 DVSS.n2644 4.5005
R19833 DVSS.n7282 DVSS.n7281 4.5005
R19834 DVSS.n7280 DVSS.n2647 4.5005
R19835 DVSS.n7279 DVSS.n7278 4.5005
R19836 DVSS.n2649 DVSS.n2648 4.5005
R19837 DVSS.n7274 DVSS.n7273 4.5005
R19838 DVSS.n7272 DVSS.n2651 4.5005
R19839 DVSS.n2701 DVSS.n2699 4.5005
R19840 DVSS.n5577 DVSS.n5576 4.5005
R19841 DVSS.n5579 DVSS.n5578 4.5005
R19842 DVSS.n5581 DVSS.n5580 4.5005
R19843 DVSS.n5583 DVSS.n5582 4.5005
R19844 DVSS.n5585 DVSS.n5584 4.5005
R19845 DVSS.n5587 DVSS.n5586 4.5005
R19846 DVSS.n5589 DVSS.n5588 4.5005
R19847 DVSS.n5591 DVSS.n5590 4.5005
R19848 DVSS.n5593 DVSS.n5592 4.5005
R19849 DVSS.n5595 DVSS.n5594 4.5005
R19850 DVSS.n5597 DVSS.n5596 4.5005
R19851 DVSS.n5599 DVSS.n5598 4.5005
R19852 DVSS.n5601 DVSS.n5600 4.5005
R19853 DVSS.n5604 DVSS.n5603 4.5005
R19854 DVSS.n5606 DVSS.n5605 4.5005
R19855 DVSS.n5608 DVSS.n5607 4.5005
R19856 DVSS.n5610 DVSS.n5609 4.5005
R19857 DVSS.n5612 DVSS.n5611 4.5005
R19858 DVSS.n5614 DVSS.n5613 4.5005
R19859 DVSS.n5616 DVSS.n5615 4.5005
R19860 DVSS.n5618 DVSS.n5617 4.5005
R19861 DVSS.n5620 DVSS.n5619 4.5005
R19862 DVSS.n5622 DVSS.n5621 4.5005
R19863 DVSS.n5624 DVSS.n5623 4.5005
R19864 DVSS.n5626 DVSS.n5625 4.5005
R19865 DVSS.n5627 DVSS.n5550 4.5005
R19866 DVSS.n5629 DVSS.n5628 4.5005
R19867 DVSS.n5641 DVSS.n5640 4.5005
R19868 DVSS.n3283 DVSS.n3282 4.5005
R19869 DVSS.n5445 DVSS.n5444 4.5005
R19870 DVSS.n5447 DVSS.n5446 4.5005
R19871 DVSS.n5448 DVSS.n5438 4.5005
R19872 DVSS.n5450 DVSS.n5449 4.5005
R19873 DVSS.n5451 DVSS.n5437 4.5005
R19874 DVSS.n5453 DVSS.n5452 4.5005
R19875 DVSS.n5454 DVSS.n5432 4.5005
R19876 DVSS.n5456 DVSS.n5455 4.5005
R19877 DVSS.n5457 DVSS.n5431 4.5005
R19878 DVSS.n5459 DVSS.n5458 4.5005
R19879 DVSS.n5460 DVSS.n5425 4.5005
R19880 DVSS.n5462 DVSS.n5461 4.5005
R19881 DVSS.n5463 DVSS.n5424 4.5005
R19882 DVSS.n5465 DVSS.n5464 4.5005
R19883 DVSS.n5466 DVSS.n5419 4.5005
R19884 DVSS.n5468 DVSS.n5467 4.5005
R19885 DVSS.n5469 DVSS.n5418 4.5005
R19886 DVSS.n5471 DVSS.n5470 4.5005
R19887 DVSS.n5472 DVSS.n5413 4.5005
R19888 DVSS.n5474 DVSS.n5473 4.5005
R19889 DVSS.n5475 DVSS.n5412 4.5005
R19890 DVSS.n5477 DVSS.n5476 4.5005
R19891 DVSS.n5478 DVSS.n5408 4.5005
R19892 DVSS.n5480 DVSS.n5479 4.5005
R19893 DVSS.n5481 DVSS.n5407 4.5005
R19894 DVSS.n5483 DVSS.n5482 4.5005
R19895 DVSS.n5697 DVSS.n3229 4.5005
R19896 DVSS.n5699 DVSS.n5698 4.5005
R19897 DVSS.n5700 DVSS.n3224 4.5005
R19898 DVSS.n5702 DVSS.n5701 4.5005
R19899 DVSS.n5703 DVSS.n3223 4.5005
R19900 DVSS.n5705 DVSS.n5704 4.5005
R19901 DVSS.n5706 DVSS.n3218 4.5005
R19902 DVSS.n5708 DVSS.n5707 4.5005
R19903 DVSS.n5709 DVSS.n3217 4.5005
R19904 DVSS.n5711 DVSS.n5710 4.5005
R19905 DVSS.n5712 DVSS.n3212 4.5005
R19906 DVSS.n5714 DVSS.n5713 4.5005
R19907 DVSS.n5715 DVSS.n3211 4.5005
R19908 DVSS.n5717 DVSS.n5716 4.5005
R19909 DVSS.n5719 DVSS.n3206 4.5005
R19910 DVSS.n5721 DVSS.n5720 4.5005
R19911 DVSS.n5722 DVSS.n3205 4.5005
R19912 DVSS.n5724 DVSS.n5723 4.5005
R19913 DVSS.n5725 DVSS.n3200 4.5005
R19914 DVSS.n5727 DVSS.n5726 4.5005
R19915 DVSS.n5728 DVSS.n3199 4.5005
R19916 DVSS.n5730 DVSS.n5729 4.5005
R19917 DVSS.n5731 DVSS.n3194 4.5005
R19918 DVSS.n5733 DVSS.n5732 4.5005
R19919 DVSS.n5734 DVSS.n3193 4.5005
R19920 DVSS.n5736 DVSS.n5735 4.5005
R19921 DVSS.n5737 DVSS.n3189 4.5005
R19922 DVSS.n5739 DVSS.n5738 4.5005
R19923 DVSS.n5199 DVSS.n3519 4.5005
R19924 DVSS.n5201 DVSS.n5200 4.5005
R19925 DVSS.n5203 DVSS.n5202 4.5005
R19926 DVSS.n5205 DVSS.n5204 4.5005
R19927 DVSS.n5206 DVSS.n3512 4.5005
R19928 DVSS.n5208 DVSS.n5207 4.5005
R19929 DVSS.n5209 DVSS.n3511 4.5005
R19930 DVSS.n5211 DVSS.n5210 4.5005
R19931 DVSS.n5212 DVSS.n3506 4.5005
R19932 DVSS.n5214 DVSS.n5213 4.5005
R19933 DVSS.n5215 DVSS.n3505 4.5005
R19934 DVSS.n5217 DVSS.n5216 4.5005
R19935 DVSS.n5218 DVSS.n3501 4.5005
R19936 DVSS.n5220 DVSS.n5219 4.5005
R19937 DVSS.n5222 DVSS.n5221 4.5005
R19938 DVSS.n5223 DVSS.n3495 4.5005
R19939 DVSS.n5225 DVSS.n5224 4.5005
R19940 DVSS.n5226 DVSS.n3494 4.5005
R19941 DVSS.n5228 DVSS.n5227 4.5005
R19942 DVSS.n5229 DVSS.n3490 4.5005
R19943 DVSS.n5231 DVSS.n5230 4.5005
R19944 DVSS.n5232 DVSS.n3488 4.5005
R19945 DVSS.n5234 DVSS.n5233 4.5005
R19946 DVSS.n3970 DVSS.n3487 4.5005
R19947 DVSS.n3987 DVSS.n3981 4.5005
R19948 DVSS.n3988 DVSS.n3980 4.5005
R19949 DVSS.n3990 DVSS.n3989 4.5005
R19950 DVSS.n3992 DVSS.n3991 4.5005
R19951 DVSS.n4093 DVSS.n3561 4.5005
R19952 DVSS.n4092 DVSS.n4091 4.5005
R19953 DVSS.n4012 DVSS.n4011 4.5005
R19954 DVSS.n4086 DVSS.n4085 4.5005
R19955 DVSS.n4084 DVSS.n4014 4.5005
R19956 DVSS.n4083 DVSS.n4082 4.5005
R19957 DVSS.n4016 DVSS.n4015 4.5005
R19958 DVSS.n4078 DVSS.n4077 4.5005
R19959 DVSS.n4076 DVSS.n4018 4.5005
R19960 DVSS.n4075 DVSS.n4074 4.5005
R19961 DVSS.n4020 DVSS.n4019 4.5005
R19962 DVSS.n4070 DVSS.n4069 4.5005
R19963 DVSS.n4068 DVSS.n4067 4.5005
R19964 DVSS.n4066 DVSS.n4022 4.5005
R19965 DVSS.n4063 DVSS.n4062 4.5005
R19966 DVSS.n4061 DVSS.n4025 4.5005
R19967 DVSS.n4060 DVSS.n4059 4.5005
R19968 DVSS.n4027 DVSS.n4026 4.5005
R19969 DVSS.n4055 DVSS.n4054 4.5005
R19970 DVSS.n4053 DVSS.n4029 4.5005
R19971 DVSS.n4052 DVSS.n4051 4.5005
R19972 DVSS.n4031 DVSS.n4030 4.5005
R19973 DVSS.n4047 DVSS.n4046 4.5005
R19974 DVSS.n4045 DVSS.n4033 4.5005
R19975 DVSS.n4044 DVSS.n4043 4.5005
R19976 DVSS.n4035 DVSS.n4034 4.5005
R19977 DVSS.n4039 DVSS.n4038 4.5005
R19978 DVSS.n4037 DVSS.n3705 4.5005
R19979 DVSS.n4812 DVSS.n4811 4.5005
R19980 DVSS.n3694 DVSS.n3687 4.5005
R19981 DVSS.n4661 DVSS.n4660 4.5005
R19982 DVSS.n4663 DVSS.n4662 4.5005
R19983 DVSS.n4665 DVSS.n4664 4.5005
R19984 DVSS.n4667 DVSS.n4666 4.5005
R19985 DVSS.n4668 DVSS.n4654 4.5005
R19986 DVSS.n4670 DVSS.n4669 4.5005
R19987 DVSS.n4671 DVSS.n4649 4.5005
R19988 DVSS.n4673 DVSS.n4672 4.5005
R19989 DVSS.n4674 DVSS.n4648 4.5005
R19990 DVSS.n4676 DVSS.n4675 4.5005
R19991 DVSS.n4677 DVSS.n4642 4.5005
R19992 DVSS.n4679 DVSS.n4678 4.5005
R19993 DVSS.n4680 DVSS.n4641 4.5005
R19994 DVSS.n4682 DVSS.n4681 4.5005
R19995 DVSS.n4683 DVSS.n4636 4.5005
R19996 DVSS.n4685 DVSS.n4684 4.5005
R19997 DVSS.n4686 DVSS.n4635 4.5005
R19998 DVSS.n4688 DVSS.n4687 4.5005
R19999 DVSS.n4689 DVSS.n4630 4.5005
R20000 DVSS.n4691 DVSS.n4690 4.5005
R20001 DVSS.n4692 DVSS.n4629 4.5005
R20002 DVSS.n4694 DVSS.n4693 4.5005
R20003 DVSS.n4696 DVSS.n4695 4.5005
R20004 DVSS.n4698 DVSS.n4697 4.5005
R20005 DVSS.n4700 DVSS.n4699 4.5005
R20006 DVSS.n4702 DVSS.n4701 4.5005
R20007 DVSS.n3698 DVSS.n3690 4.5005
R20008 DVSS.n3703 DVSS.n3698 4.5005
R20009 DVSS.n4809 DVSS.n3698 4.5005
R20010 DVSS.n3696 DVSS.n3690 4.5005
R20011 DVSS.n3703 DVSS.n3696 4.5005
R20012 DVSS.n4809 DVSS.n3696 4.5005
R20013 DVSS.n3699 DVSS.n3690 4.5005
R20014 DVSS.n3703 DVSS.n3699 4.5005
R20015 DVSS.n4809 DVSS.n3699 4.5005
R20016 DVSS.n3695 DVSS.n3690 4.5005
R20017 DVSS.n3703 DVSS.n3695 4.5005
R20018 DVSS.n4809 DVSS.n3695 4.5005
R20019 DVSS.n3690 DVSS.n3688 4.5005
R20020 DVSS.n3703 DVSS.n3688 4.5005
R20021 DVSS.n4809 DVSS.n3688 4.5005
R20022 DVSS.n4810 DVSS.n3690 4.5005
R20023 DVSS.n4810 DVSS.n4809 4.5005
R20024 DVSS.n3700 DVSS.n3690 4.5005
R20025 DVSS.n4809 DVSS.n3700 4.5005
R20026 DVSS.n3693 DVSS.n3690 4.5005
R20027 DVSS.n3703 DVSS.n3693 4.5005
R20028 DVSS.n4809 DVSS.n3693 4.5005
R20029 DVSS.n3701 DVSS.n3690 4.5005
R20030 DVSS.n3703 DVSS.n3701 4.5005
R20031 DVSS.n4809 DVSS.n3701 4.5005
R20032 DVSS.n3692 DVSS.n3690 4.5005
R20033 DVSS.n3703 DVSS.n3692 4.5005
R20034 DVSS.n4809 DVSS.n3692 4.5005
R20035 DVSS.n4808 DVSS.n3690 4.5005
R20036 DVSS.n4808 DVSS.n3703 4.5005
R20037 DVSS.n4809 DVSS.n4808 4.5005
R20038 DVSS.n4103 DVSS.n3977 4.5005
R20039 DVSS.n4105 DVSS.n3977 4.5005
R20040 DVSS.n3977 DVSS.n3969 4.5005
R20041 DVSS.n4103 DVSS.n3975 4.5005
R20042 DVSS.n4105 DVSS.n3975 4.5005
R20043 DVSS.n3975 DVSS.n3969 4.5005
R20044 DVSS.n4103 DVSS.n3978 4.5005
R20045 DVSS.n4105 DVSS.n3978 4.5005
R20046 DVSS.n3978 DVSS.n3969 4.5005
R20047 DVSS.n4103 DVSS.n3974 4.5005
R20048 DVSS.n4105 DVSS.n3974 4.5005
R20049 DVSS.n3974 DVSS.n3969 4.5005
R20050 DVSS.n4103 DVSS.n4102 4.5005
R20051 DVSS.n4102 DVSS.n3969 4.5005
R20052 DVSS.n4103 DVSS.n3993 4.5005
R20053 DVSS.n3993 DVSS.n3969 4.5005
R20054 DVSS.n4103 DVSS.n3979 4.5005
R20055 DVSS.n4105 DVSS.n3979 4.5005
R20056 DVSS.n3979 DVSS.n3969 4.5005
R20057 DVSS.n4103 DVSS.n3972 4.5005
R20058 DVSS.n4105 DVSS.n3972 4.5005
R20059 DVSS.n3972 DVSS.n3969 4.5005
R20060 DVSS.n4104 DVSS.n4103 4.5005
R20061 DVSS.n4105 DVSS.n4104 4.5005
R20062 DVSS.n4104 DVSS.n3969 4.5005
R20063 DVSS.n4103 DVSS.n3971 4.5005
R20064 DVSS.n4105 DVSS.n3971 4.5005
R20065 DVSS.n3971 DVSS.n3969 4.5005
R20066 DVSS.n4103 DVSS.n3489 4.5005
R20067 DVSS.n4105 DVSS.n3489 4.5005
R20068 DVSS.n3969 DVSS.n3489 4.5005
R20069 DVSS.n5741 DVSS.n3182 4.5005
R20070 DVSS.n3182 DVSS.n3175 4.5005
R20071 DVSS.n3182 DVSS.n3170 4.5005
R20072 DVSS.n5741 DVSS.n3180 4.5005
R20073 DVSS.n3180 DVSS.n3175 4.5005
R20074 DVSS.n3180 DVSS.n3170 4.5005
R20075 DVSS.n5741 DVSS.n3183 4.5005
R20076 DVSS.n3183 DVSS.n3175 4.5005
R20077 DVSS.n3183 DVSS.n3170 4.5005
R20078 DVSS.n5741 DVSS.n3179 4.5005
R20079 DVSS.n3179 DVSS.n3175 4.5005
R20080 DVSS.n3179 DVSS.n3170 4.5005
R20081 DVSS.n5741 DVSS.n3185 4.5005
R20082 DVSS.n3185 DVSS.n3170 4.5005
R20083 DVSS.n5741 DVSS.n3178 4.5005
R20084 DVSS.n3178 DVSS.n3170 4.5005
R20085 DVSS.n3186 DVSS.n3170 4.5005
R20086 DVSS.n3186 DVSS.n3175 4.5005
R20087 DVSS.n5741 DVSS.n3186 4.5005
R20088 DVSS.n3177 DVSS.n3170 4.5005
R20089 DVSS.n3177 DVSS.n3175 4.5005
R20090 DVSS.n5741 DVSS.n3177 4.5005
R20091 DVSS.n3187 DVSS.n3170 4.5005
R20092 DVSS.n3187 DVSS.n3175 4.5005
R20093 DVSS.n5741 DVSS.n3187 4.5005
R20094 DVSS.n3176 DVSS.n3170 4.5005
R20095 DVSS.n3176 DVSS.n3175 4.5005
R20096 DVSS.n5741 DVSS.n3176 4.5005
R20097 DVSS.n5740 DVSS.n3170 4.5005
R20098 DVSS.n5740 DVSS.n3175 4.5005
R20099 DVSS.n5741 DVSS.n5740 4.5005
R20100 DVSS.n7936 DVSS.n2051 4.5005
R20101 DVSS.n2051 DVSS.n2044 4.5005
R20102 DVSS.n2051 DVSS.n2039 4.5005
R20103 DVSS.n7936 DVSS.n2049 4.5005
R20104 DVSS.n2049 DVSS.n2044 4.5005
R20105 DVSS.n2049 DVSS.n2039 4.5005
R20106 DVSS.n7936 DVSS.n2052 4.5005
R20107 DVSS.n2052 DVSS.n2044 4.5005
R20108 DVSS.n2052 DVSS.n2039 4.5005
R20109 DVSS.n7936 DVSS.n2048 4.5005
R20110 DVSS.n2048 DVSS.n2044 4.5005
R20111 DVSS.n2048 DVSS.n2039 4.5005
R20112 DVSS.n7936 DVSS.n2053 4.5005
R20113 DVSS.n2053 DVSS.n2044 4.5005
R20114 DVSS.n2053 DVSS.n2039 4.5005
R20115 DVSS.n7936 DVSS.n2047 4.5005
R20116 DVSS.n2047 DVSS.n2044 4.5005
R20117 DVSS.n2047 DVSS.n2039 4.5005
R20118 DVSS.n7936 DVSS.n2054 4.5005
R20119 DVSS.n2054 DVSS.n2044 4.5005
R20120 DVSS.n2054 DVSS.n2039 4.5005
R20121 DVSS.n7936 DVSS.n2046 4.5005
R20122 DVSS.n2046 DVSS.n2044 4.5005
R20123 DVSS.n2046 DVSS.n2039 4.5005
R20124 DVSS.n7936 DVSS.n2055 4.5005
R20125 DVSS.n2055 DVSS.n2044 4.5005
R20126 DVSS.n2055 DVSS.n2039 4.5005
R20127 DVSS.n7936 DVSS.n2045 4.5005
R20128 DVSS.n2045 DVSS.n2044 4.5005
R20129 DVSS.n2045 DVSS.n2039 4.5005
R20130 DVSS.n7936 DVSS.n7935 4.5005
R20131 DVSS.n7935 DVSS.n2044 4.5005
R20132 DVSS.n7935 DVSS.n2039 4.5005
R20133 DVSS.n8400 DVSS.n1368 4.5005
R20134 DVSS.n8403 DVSS.n1368 4.5005
R20135 DVSS.n8403 DVSS.n1366 4.5005
R20136 DVSS.n8403 DVSS.n1369 4.5005
R20137 DVSS.n8403 DVSS.n1365 4.5005
R20138 DVSS.n1377 DVSS.n1370 4.5005
R20139 DVSS.n8403 DVSS.n1370 4.5005
R20140 DVSS.n8400 DVSS.n1364 4.5005
R20141 DVSS.n1377 DVSS.n1364 4.5005
R20142 DVSS.n8403 DVSS.n1364 4.5005
R20143 DVSS.n8403 DVSS.n1371 4.5005
R20144 DVSS.n8400 DVSS.n1371 4.5005
R20145 DVSS.n8403 DVSS.n1363 4.5005
R20146 DVSS.n8403 DVSS.n1372 4.5005
R20147 DVSS.n8403 DVSS.n1362 4.5005
R20148 DVSS.n8402 DVSS.n1377 4.5005
R20149 DVSS.n8403 DVSS.n8402 4.5005
R20150 DVSS.n8519 DVSS.n1082 4.5005
R20151 DVSS.n8515 DVSS.n1082 4.5005
R20152 DVSS.n8510 DVSS.n8509 4.5005
R20153 DVSS.n8504 DVSS.n8503 4.5005
R20154 DVSS.n8508 DVSS.n8507 4.5005
R20155 DVSS.n8514 DVSS.n8513 4.5005
R20156 DVSS.n8525 DVSS.n8521 4.5005
R20157 DVSS.n8526 DVSS.n8525 4.5005
R20158 DVSS.n1215 DVSS.n1076 4.5005
R20159 DVSS.n8529 DVSS.n1076 4.5005
R20160 DVSS.n8527 DVSS.n1076 4.5005
R20161 DVSS.n8532 DVSS.n8531 4.5005
R20162 DVSS.n7150 DVSS.n7141 4.5005
R20163 DVSS.n7150 DVSS.n7149 4.5005
R20164 DVSS.n7149 DVSS.n7148 4.5005
R20165 DVSS.n7148 DVSS.n7147 4.5005
R20166 DVSS.n7114 DVSS.n1484 4.5005
R20167 DVSS.n7112 DVSS.n1484 4.5005
R20168 DVSS.n8293 DVSS.n1482 4.5005
R20169 DVSS.n1489 DVSS.n1482 4.5005
R20170 DVSS.n8291 DVSS.n1482 4.5005
R20171 DVSS.n1490 DVSS.n1489 4.5005
R20172 DVSS.n8291 DVSS.n1490 4.5005
R20173 DVSS.n8243 DVSS.n8241 4.5005
R20174 DVSS.n8246 DVSS.n8241 4.5005
R20175 DVSS.n8249 DVSS.n8241 4.5005
R20176 DVSS.n8246 DVSS.n8239 4.5005
R20177 DVSS.n8249 DVSS.n8239 4.5005
R20178 DVSS.n8236 DVSS.n1513 4.5005
R20179 DVSS.n8236 DVSS.n8235 4.5005
R20180 DVSS.n8237 DVSS.n8236 4.5005
R20181 DVSS.n8235 DVSS.n1516 4.5005
R20182 DVSS.n8237 DVSS.n1516 4.5005
R20183 DVSS.n8238 DVSS.n1513 4.5005
R20184 DVSS.n8238 DVSS.n8237 4.5005
R20185 DVSS.n8248 DVSS.n8243 4.5005
R20186 DVSS.n8249 DVSS.n8248 4.5005
R20187 DVSS.n8293 DVSS.n8292 4.5005
R20188 DVSS.n8292 DVSS.n8291 4.5005
R20189 DVSS.n7118 DVSS.n7112 4.5005
R20190 DVSS.n7118 DVSS.n7117 4.5005
R20191 DVSS.n7153 DVSS.n7135 4.5005
R20192 DVSS.n7153 DVSS.n7152 4.5005
R20193 DVSS.n7154 DVSS.n7153 4.5005
R20194 DVSS.n7152 DVSS.n6650 4.5005
R20195 DVSS.n7154 DVSS.n6650 4.5005
R20196 DVSS.n7152 DVSS.n7151 4.5005
R20197 DVSS.n7151 DVSS.n7135 4.5005
R20198 DVSS.n4787 DVSS.n3720 4.5005
R20199 DVSS.n4787 DVSS.n3721 4.5005
R20200 DVSS.n4796 DVSS.n4787 4.5005
R20201 DVSS.n3725 DVSS.n3721 4.5005
R20202 DVSS.n4796 DVSS.n3725 4.5005
R20203 DVSS.n4790 DVSS.n3721 4.5005
R20204 DVSS.n4796 DVSS.n4790 4.5005
R20205 DVSS.n3724 DVSS.n3721 4.5005
R20206 DVSS.n4796 DVSS.n3724 4.5005
R20207 DVSS.n4793 DVSS.n3721 4.5005
R20208 DVSS.n4796 DVSS.n4793 4.5005
R20209 DVSS.n3723 DVSS.n3721 4.5005
R20210 DVSS.n4796 DVSS.n3723 4.5005
R20211 DVSS.n4795 DVSS.n3721 4.5005
R20212 DVSS.n4795 DVSS.n3719 4.5005
R20213 DVSS.n4796 DVSS.n4795 4.5005
R20214 DVSS.n3720 DVSS.n3714 4.5005
R20215 DVSS.n3721 DVSS.n3714 4.5005
R20216 DVSS.n3719 DVSS.n3714 4.5005
R20217 DVSS.n4796 DVSS.n3714 4.5005
R20218 DVSS.n3720 DVSS.n3717 4.5005
R20219 DVSS.n3721 DVSS.n3717 4.5005
R20220 DVSS.n3719 DVSS.n3717 4.5005
R20221 DVSS.n4796 DVSS.n3717 4.5005
R20222 DVSS.n3720 DVSS.n3718 4.5005
R20223 DVSS.n3721 DVSS.n3718 4.5005
R20224 DVSS.n3719 DVSS.n3718 4.5005
R20225 DVSS.n4796 DVSS.n3718 4.5005
R20226 DVSS.n4797 DVSS.n3720 4.5005
R20227 DVSS.n4797 DVSS.n3721 4.5005
R20228 DVSS.n4797 DVSS.n3719 4.5005
R20229 DVSS.n4797 DVSS.n4796 4.5005
R20230 DVSS.n3950 DVSS.n3937 4.5005
R20231 DVSS.n4137 DVSS.n3937 4.5005
R20232 DVSS.n3946 DVSS.n3937 4.5005
R20233 DVSS.n4139 DVSS.n3937 4.5005
R20234 DVSS.n3950 DVSS.n3935 4.5005
R20235 DVSS.n4137 DVSS.n3935 4.5005
R20236 DVSS.n3946 DVSS.n3935 4.5005
R20237 DVSS.n4139 DVSS.n3935 4.5005
R20238 DVSS.n3950 DVSS.n3938 4.5005
R20239 DVSS.n4137 DVSS.n3938 4.5005
R20240 DVSS.n3946 DVSS.n3938 4.5005
R20241 DVSS.n4139 DVSS.n3938 4.5005
R20242 DVSS.n3950 DVSS.n3934 4.5005
R20243 DVSS.n4137 DVSS.n3934 4.5005
R20244 DVSS.n3946 DVSS.n3934 4.5005
R20245 DVSS.n4139 DVSS.n3934 4.5005
R20246 DVSS.n3950 DVSS.n3939 4.5005
R20247 DVSS.n4137 DVSS.n3939 4.5005
R20248 DVSS.n4139 DVSS.n3939 4.5005
R20249 DVSS.n4137 DVSS.n3933 4.5005
R20250 DVSS.n4139 DVSS.n3933 4.5005
R20251 DVSS.n4137 DVSS.n3940 4.5005
R20252 DVSS.n4139 DVSS.n3940 4.5005
R20253 DVSS.n4137 DVSS.n3932 4.5005
R20254 DVSS.n4139 DVSS.n3932 4.5005
R20255 DVSS.n4137 DVSS.n3941 4.5005
R20256 DVSS.n4139 DVSS.n3941 4.5005
R20257 DVSS.n4137 DVSS.n3931 4.5005
R20258 DVSS.n4139 DVSS.n3931 4.5005
R20259 DVSS.n4138 DVSS.n4137 4.5005
R20260 DVSS.n4138 DVSS.n3946 4.5005
R20261 DVSS.n4139 DVSS.n4138 4.5005
R20262 DVSS.n5775 DVSS.n3149 4.5005
R20263 DVSS.n5777 DVSS.n3149 4.5005
R20264 DVSS.n3149 DVSS.n3136 4.5005
R20265 DVSS.n5777 DVSS.n3146 4.5005
R20266 DVSS.n3146 DVSS.n3136 4.5005
R20267 DVSS.n5777 DVSS.n3151 4.5005
R20268 DVSS.n3151 DVSS.n3136 4.5005
R20269 DVSS.n5777 DVSS.n3145 4.5005
R20270 DVSS.n3145 DVSS.n3136 4.5005
R20271 DVSS.n5777 DVSS.n3153 4.5005
R20272 DVSS.n3153 DVSS.n3136 4.5005
R20273 DVSS.n5775 DVSS.n3144 4.5005
R20274 DVSS.n5777 DVSS.n3144 4.5005
R20275 DVSS.n3144 DVSS.n3136 4.5005
R20276 DVSS.n3154 DVSS.n3136 4.5005
R20277 DVSS.n3154 DVSS.n3141 4.5005
R20278 DVSS.n5777 DVSS.n3154 4.5005
R20279 DVSS.n5775 DVSS.n3154 4.5005
R20280 DVSS.n3143 DVSS.n3136 4.5005
R20281 DVSS.n3143 DVSS.n3141 4.5005
R20282 DVSS.n5777 DVSS.n3143 4.5005
R20283 DVSS.n5775 DVSS.n3143 4.5005
R20284 DVSS.n3155 DVSS.n3136 4.5005
R20285 DVSS.n3155 DVSS.n3141 4.5005
R20286 DVSS.n5777 DVSS.n3155 4.5005
R20287 DVSS.n5775 DVSS.n3155 4.5005
R20288 DVSS.n3142 DVSS.n3136 4.5005
R20289 DVSS.n3142 DVSS.n3141 4.5005
R20290 DVSS.n5777 DVSS.n3142 4.5005
R20291 DVSS.n5775 DVSS.n3142 4.5005
R20292 DVSS.n5776 DVSS.n3136 4.5005
R20293 DVSS.n5776 DVSS.n3141 4.5005
R20294 DVSS.n5777 DVSS.n5776 4.5005
R20295 DVSS.n5776 DVSS.n5775 4.5005
R20296 DVSS.n7972 DVSS.n2018 4.5005
R20297 DVSS.n7975 DVSS.n2018 4.5005
R20298 DVSS.n2018 DVSS.n2005 4.5005
R20299 DVSS.n7975 DVSS.n2015 4.5005
R20300 DVSS.n2015 DVSS.n2005 4.5005
R20301 DVSS.n7975 DVSS.n2020 4.5005
R20302 DVSS.n2020 DVSS.n2005 4.5005
R20303 DVSS.n7975 DVSS.n2014 4.5005
R20304 DVSS.n2014 DVSS.n2005 4.5005
R20305 DVSS.n7975 DVSS.n2022 4.5005
R20306 DVSS.n2022 DVSS.n2005 4.5005
R20307 DVSS.n7975 DVSS.n2013 4.5005
R20308 DVSS.n2013 DVSS.n2005 4.5005
R20309 DVSS.n7975 DVSS.n2024 4.5005
R20310 DVSS.n2024 DVSS.n2005 4.5005
R20311 DVSS.n7975 DVSS.n2012 4.5005
R20312 DVSS.n2012 DVSS.n2005 4.5005
R20313 DVSS.n7975 DVSS.n2026 4.5005
R20314 DVSS.n2026 DVSS.n2005 4.5005
R20315 DVSS.n7975 DVSS.n2011 4.5005
R20316 DVSS.n2011 DVSS.n2005 4.5005
R20317 DVSS.n7975 DVSS.n7974 4.5005
R20318 DVSS.n7974 DVSS.n2010 4.5005
R20319 DVSS.n7974 DVSS.n2005 4.5005
R20320 DVSS.n1335 DVSS.n1326 4.5005
R20321 DVSS.n1335 DVSS.n1327 4.5005
R20322 DVSS.n8439 DVSS.n1335 4.5005
R20323 DVSS.n1333 DVSS.n1327 4.5005
R20324 DVSS.n8439 DVSS.n1333 4.5005
R20325 DVSS.n1337 DVSS.n1327 4.5005
R20326 DVSS.n8439 DVSS.n1337 4.5005
R20327 DVSS.n1332 DVSS.n1327 4.5005
R20328 DVSS.n8439 DVSS.n1332 4.5005
R20329 DVSS.n1339 DVSS.n1327 4.5005
R20330 DVSS.n8435 DVSS.n1339 4.5005
R20331 DVSS.n8439 DVSS.n1339 4.5005
R20332 DVSS.n1331 DVSS.n1326 4.5005
R20333 DVSS.n1331 DVSS.n1327 4.5005
R20334 DVSS.n8435 DVSS.n1331 4.5005
R20335 DVSS.n8439 DVSS.n1331 4.5005
R20336 DVSS.n8439 DVSS.n1341 4.5005
R20337 DVSS.n8435 DVSS.n1341 4.5005
R20338 DVSS.n1341 DVSS.n1326 4.5005
R20339 DVSS.n1330 DVSS.n1326 4.5005
R20340 DVSS.n8439 DVSS.n1330 4.5005
R20341 DVSS.n8438 DVSS.n1327 4.5005
R20342 DVSS.n8439 DVSS.n8438 4.5005
R20343 DVSS.n1329 DVSS.n1327 4.5005
R20344 DVSS.n8439 DVSS.n1329 4.5005
R20345 DVSS.n8440 DVSS.n1326 4.5005
R20346 DVSS.n8440 DVSS.n1327 4.5005
R20347 DVSS.n8440 DVSS.n8439 4.5005
R20348 DVSS.n1387 DVSS.n1145 4.5005
R20349 DVSS.n8475 DVSS.n8474 4.5005
R20350 DVSS.n8479 DVSS.n8478 4.5005
R20351 DVSS.n8480 DVSS.n8479 4.5005
R20352 DVSS.n8487 DVSS.n1128 4.5005
R20353 DVSS.n8487 DVSS.n8486 4.5005
R20354 DVSS.n8486 DVSS.n8483 4.5005
R20355 DVSS.n8483 DVSS.n1128 4.5005
R20356 DVSS.n8483 DVSS.n8482 4.5005
R20357 DVSS.n8480 DVSS.n1134 4.5005
R20358 DVSS.n8478 DVSS.n1134 4.5005
R20359 DVSS.n8476 DVSS.n1134 4.5005
R20360 DVSS.n8475 DVSS.n1142 4.5005
R20361 DVSS.n8468 DVSS.n1142 4.5005
R20362 DVSS.n1383 DVSS.n1145 4.5005
R20363 DVSS.n1383 DVSS.n1379 4.5005
R20364 DVSS.n8444 DVSS.n1324 4.5005
R20365 DVSS.n8481 DVSS.n1128 4.5005
R20366 DVSS.n8482 DVSS.n8481 4.5005
R20367 DVSS.n8478 DVSS.n8477 4.5005
R20368 DVSS.n8477 DVSS.n8476 4.5005
R20369 DVSS.n8470 DVSS.n8468 4.5005
R20370 DVSS.n1382 DVSS.n1379 4.5005
R20371 DVSS.n8447 DVSS.n1324 4.5005
R20372 DVSS.n8447 DVSS.n1323 4.5005
R20373 DVSS.n8447 DVSS.n8446 4.5005
R20374 DVSS.n8448 DVSS.n8447 4.5005
R20375 DVSS.n1283 DVSS.n1282 4.5005
R20376 DVSS.n1282 DVSS.n1281 4.5005
R20377 DVSS.n1277 DVSS.n1276 4.5005
R20378 DVSS.n1268 DVSS.n1267 4.5005
R20379 DVSS.n1263 DVSS.n1262 4.5005
R20380 DVSS.n1262 DVSS.n1261 4.5005
R20381 DVSS.n1258 DVSS.n1257 4.5005
R20382 DVSS.n1257 DVSS.n1256 4.5005
R20383 DVSS.n1256 DVSS.n1249 4.5005
R20384 DVSS.n1260 DVSS.n1249 4.5005
R20385 DVSS.n1261 DVSS.n1242 4.5005
R20386 DVSS.n1265 DVSS.n1242 4.5005
R20387 DVSS.n1268 DVSS.n1238 4.5005
R20388 DVSS.n1240 DVSS.n1238 4.5005
R20389 DVSS.n1271 DVSS.n1238 4.5005
R20390 DVSS.n1277 DVSS.n1234 4.5005
R20391 DVSS.n1236 DVSS.n1234 4.5005
R20392 DVSS.n1280 DVSS.n1234 4.5005
R20393 DVSS.n1281 DVSS.n1227 4.5005
R20394 DVSS.n1285 DVSS.n1227 4.5005
R20395 DVSS.n1259 DVSS.n1258 4.5005
R20396 DVSS.n1259 DVSS.n1251 4.5005
R20397 DVSS.n1260 DVSS.n1259 4.5005
R20398 DVSS.n1264 DVSS.n1263 4.5005
R20399 DVSS.n1264 DVSS.n1244 4.5005
R20400 DVSS.n1265 DVSS.n1264 4.5005
R20401 DVSS.n1270 DVSS.n1240 4.5005
R20402 DVSS.n1271 DVSS.n1270 4.5005
R20403 DVSS.n1279 DVSS.n1236 4.5005
R20404 DVSS.n1280 DVSS.n1279 4.5005
R20405 DVSS.n1284 DVSS.n1283 4.5005
R20406 DVSS.n1284 DVSS.n1229 4.5005
R20407 DVSS.n1285 DVSS.n1284 4.5005
R20408 DVSS.n8372 DVSS.n8362 4.5005
R20409 DVSS.n8376 DVSS.n8358 4.5005
R20410 DVSS.n8378 DVSS.n8358 4.5005
R20411 DVSS.n8385 DVSS.n1405 4.5005
R20412 DVSS.n8355 DVSS.n1405 4.5005
R20413 DVSS.n8350 DVSS.n1104 4.5005
R20414 DVSS.n8496 DVSS.n1098 4.5005
R20415 DVSS.n8491 DVSS.n1103 4.5005
R20416 DVSS.n8494 DVSS.n8491 4.5005
R20417 DVSS.n8352 DVSS.n1417 4.5005
R20418 DVSS.n8354 DVSS.n1417 4.5005
R20419 DVSS.n8385 DVSS.n8382 4.5005
R20420 DVSS.n8376 DVSS.n8373 4.5005
R20421 DVSS.n8367 DVSS.n8366 4.5005
R20422 DVSS.n8370 DVSS.n8367 4.5005
R20423 DVSS.n8496 DVSS.n8495 4.5005
R20424 DVSS.n8495 DVSS.n1100 4.5005
R20425 DVSS.n8495 DVSS.n1103 4.5005
R20426 DVSS.n8495 DVSS.n8494 4.5005
R20427 DVSS.n8353 DVSS.n1104 4.5005
R20428 DVSS.n8353 DVSS.n1421 4.5005
R20429 DVSS.n8353 DVSS.n8352 4.5005
R20430 DVSS.n8354 DVSS.n8353 4.5005
R20431 DVSS.n8386 DVSS.n8355 4.5005
R20432 DVSS.n8386 DVSS.n8356 4.5005
R20433 DVSS.n8386 DVSS.n8385 4.5005
R20434 DVSS.n8378 DVSS.n8377 4.5005
R20435 DVSS.n8377 DVSS.n8360 4.5005
R20436 DVSS.n8377 DVSS.n8376 4.5005
R20437 DVSS.n8372 DVSS.n8371 4.5005
R20438 DVSS.n8371 DVSS.n8364 4.5005
R20439 DVSS.n8371 DVSS.n8366 4.5005
R20440 DVSS.n8371 DVSS.n8370 4.5005
R20441 DVSS.n7121 DVSS.n7119 4.5005
R20442 DVSS.n7119 DVSS.n7077 4.5005
R20443 DVSS.n7109 DVSS.n7108 4.5005
R20444 DVSS.n7098 DVSS.n1440 4.5005
R20445 DVSS.n8336 DVSS.n8335 4.5005
R20446 DVSS.n8336 DVSS.n1438 4.5005
R20447 DVSS.n1550 DVSS.n1549 4.5005
R20448 DVSS.n1550 DVSS.n1095 4.5005
R20449 DVSS.n1546 DVSS.n1095 4.5005
R20450 DVSS.n1546 DVSS.n1545 4.5005
R20451 DVSS.n8339 DVSS.n1438 4.5005
R20452 DVSS.n8339 DVSS.n8338 4.5005
R20453 DVSS.n7102 DVSS.n1440 4.5005
R20454 DVSS.n7102 DVSS.n7101 4.5005
R20455 DVSS.n7103 DVSS.n7102 4.5005
R20456 DVSS.n7108 DVSS.n7107 4.5005
R20457 DVSS.n7107 DVSS.n7105 4.5005
R20458 DVSS.n7107 DVSS.n7106 4.5005
R20459 DVSS.n7123 DVSS.n7077 4.5005
R20460 DVSS.n7124 DVSS.n7123 4.5005
R20461 DVSS.n7129 DVSS.n1151 4.5005
R20462 DVSS.n7129 DVSS.n7128 4.5005
R20463 DVSS.n7128 DVSS.n7127 4.5005
R20464 DVSS.n7127 DVSS.n7126 4.5005
R20465 DVSS.n1216 DVSS.n1214 4.5005
R20466 DVSS.n8454 DVSS.n1158 4.5005
R20467 DVSS.n8456 DVSS.n1152 4.5005
R20468 DVSS.n8458 DVSS.n1152 4.5005
R20469 DVSS.n8457 DVSS.n1158 4.5005
R20470 DVSS.n8457 DVSS.n1155 4.5005
R20471 DVSS.n8457 DVSS.n8456 4.5005
R20472 DVSS.n8458 DVSS.n8457 4.5005
R20473 DVSS.n8450 DVSS.n1183 4.5005
R20474 DVSS.n8450 DVSS.n8449 4.5005
R20475 DVSS.n8449 DVSS.n1319 4.5005
R20476 DVSS.n1319 DVSS.n1183 4.5005
R20477 DVSS.n1319 DVSS.n1318 4.5005
R20478 DVSS.n1317 DVSS.n1183 4.5005
R20479 DVSS.n1318 DVSS.n1317 4.5005
R20480 DVSS.n1288 DVSS.n1287 4.5005
R20481 DVSS.n1287 DVSS.n1286 4.5005
R20482 DVSS.n1286 DVSS.n1220 4.5005
R20483 DVSS.n1290 DVSS.n1220 4.5005
R20484 DVSS.n1289 DVSS.n1288 4.5005
R20485 DVSS.n1289 DVSS.n1222 4.5005
R20486 DVSS.n1290 DVSS.n1289 4.5005
R20487 DVSS.n1296 DVSS.n1295 4.5005
R20488 DVSS.n4420 DVSS.n4200 4.5005
R20489 DVSS.n4420 DVSS.n4201 4.5005
R20490 DVSS.n4429 DVSS.n4420 4.5005
R20491 DVSS.n4205 DVSS.n4201 4.5005
R20492 DVSS.n4429 DVSS.n4205 4.5005
R20493 DVSS.n4423 DVSS.n4201 4.5005
R20494 DVSS.n4429 DVSS.n4423 4.5005
R20495 DVSS.n4204 DVSS.n4201 4.5005
R20496 DVSS.n4429 DVSS.n4204 4.5005
R20497 DVSS.n4426 DVSS.n4201 4.5005
R20498 DVSS.n4429 DVSS.n4426 4.5005
R20499 DVSS.n4203 DVSS.n4201 4.5005
R20500 DVSS.n4429 DVSS.n4203 4.5005
R20501 DVSS.n4428 DVSS.n4201 4.5005
R20502 DVSS.n4428 DVSS.n4199 4.5005
R20503 DVSS.n4429 DVSS.n4428 4.5005
R20504 DVSS.n4200 DVSS.n4193 4.5005
R20505 DVSS.n4201 DVSS.n4193 4.5005
R20506 DVSS.n4199 DVSS.n4193 4.5005
R20507 DVSS.n4429 DVSS.n4193 4.5005
R20508 DVSS.n4200 DVSS.n4195 4.5005
R20509 DVSS.n4201 DVSS.n4195 4.5005
R20510 DVSS.n4199 DVSS.n4195 4.5005
R20511 DVSS.n4429 DVSS.n4195 4.5005
R20512 DVSS.n4200 DVSS.n4198 4.5005
R20513 DVSS.n4201 DVSS.n4198 4.5005
R20514 DVSS.n4199 DVSS.n4198 4.5005
R20515 DVSS.n4429 DVSS.n4198 4.5005
R20516 DVSS.n4430 DVSS.n4200 4.5005
R20517 DVSS.n4430 DVSS.n4201 4.5005
R20518 DVSS.n4430 DVSS.n4199 4.5005
R20519 DVSS.n4430 DVSS.n4429 4.5005
R20520 DVSS.n3888 DVSS.n3879 4.5005
R20521 DVSS.n3889 DVSS.n3879 4.5005
R20522 DVSS.n3887 DVSS.n3879 4.5005
R20523 DVSS.n4186 DVSS.n3879 4.5005
R20524 DVSS.n4187 DVSS.n3888 4.5005
R20525 DVSS.n4187 DVSS.n3889 4.5005
R20526 DVSS.n4187 DVSS.n3887 4.5005
R20527 DVSS.n4187 DVSS.n4186 4.5005
R20528 DVSS.n4175 DVSS.n3888 4.5005
R20529 DVSS.n4175 DVSS.n3889 4.5005
R20530 DVSS.n4175 DVSS.n3887 4.5005
R20531 DVSS.n4186 DVSS.n4175 4.5005
R20532 DVSS.n3894 DVSS.n3888 4.5005
R20533 DVSS.n3894 DVSS.n3889 4.5005
R20534 DVSS.n3894 DVSS.n3887 4.5005
R20535 DVSS.n4186 DVSS.n3894 4.5005
R20536 DVSS.n4177 DVSS.n3888 4.5005
R20537 DVSS.n4177 DVSS.n3889 4.5005
R20538 DVSS.n4186 DVSS.n4177 4.5005
R20539 DVSS.n3893 DVSS.n3889 4.5005
R20540 DVSS.n4186 DVSS.n3893 4.5005
R20541 DVSS.n4180 DVSS.n3889 4.5005
R20542 DVSS.n4186 DVSS.n4180 4.5005
R20543 DVSS.n3892 DVSS.n3889 4.5005
R20544 DVSS.n4186 DVSS.n3892 4.5005
R20545 DVSS.n4183 DVSS.n3889 4.5005
R20546 DVSS.n4186 DVSS.n4183 4.5005
R20547 DVSS.n3891 DVSS.n3889 4.5005
R20548 DVSS.n4186 DVSS.n3891 4.5005
R20549 DVSS.n4185 DVSS.n3889 4.5005
R20550 DVSS.n4185 DVSS.n3887 4.5005
R20551 DVSS.n4186 DVSS.n4185 4.5005
R20552 DVSS.n5811 DVSS.n3106 4.5005
R20553 DVSS.n3112 DVSS.n3106 4.5005
R20554 DVSS.n5813 DVSS.n3106 4.5005
R20555 DVSS.n3112 DVSS.n3104 4.5005
R20556 DVSS.n5813 DVSS.n3104 4.5005
R20557 DVSS.n3112 DVSS.n3107 4.5005
R20558 DVSS.n5813 DVSS.n3107 4.5005
R20559 DVSS.n3112 DVSS.n3103 4.5005
R20560 DVSS.n5813 DVSS.n3103 4.5005
R20561 DVSS.n3112 DVSS.n3108 4.5005
R20562 DVSS.n5813 DVSS.n3108 4.5005
R20563 DVSS.n5811 DVSS.n3102 4.5005
R20564 DVSS.n3112 DVSS.n3102 4.5005
R20565 DVSS.n5813 DVSS.n3102 4.5005
R20566 DVSS.n5813 DVSS.n3109 4.5005
R20567 DVSS.n3117 DVSS.n3109 4.5005
R20568 DVSS.n3112 DVSS.n3109 4.5005
R20569 DVSS.n5811 DVSS.n3109 4.5005
R20570 DVSS.n5813 DVSS.n3101 4.5005
R20571 DVSS.n3117 DVSS.n3101 4.5005
R20572 DVSS.n3112 DVSS.n3101 4.5005
R20573 DVSS.n5811 DVSS.n3101 4.5005
R20574 DVSS.n5813 DVSS.n3110 4.5005
R20575 DVSS.n3117 DVSS.n3110 4.5005
R20576 DVSS.n3112 DVSS.n3110 4.5005
R20577 DVSS.n5811 DVSS.n3110 4.5005
R20578 DVSS.n5813 DVSS.n3100 4.5005
R20579 DVSS.n3117 DVSS.n3100 4.5005
R20580 DVSS.n3112 DVSS.n3100 4.5005
R20581 DVSS.n5811 DVSS.n3100 4.5005
R20582 DVSS.n5813 DVSS.n5812 4.5005
R20583 DVSS.n5812 DVSS.n3117 4.5005
R20584 DVSS.n5812 DVSS.n3112 4.5005
R20585 DVSS.n5812 DVSS.n5811 4.5005
R20586 DVSS.n8011 DVSS.n1984 4.5005
R20587 DVSS.n8014 DVSS.n1984 4.5005
R20588 DVSS.n1984 DVSS.n1971 4.5005
R20589 DVSS.n8014 DVSS.n1981 4.5005
R20590 DVSS.n1981 DVSS.n1971 4.5005
R20591 DVSS.n8014 DVSS.n1986 4.5005
R20592 DVSS.n1986 DVSS.n1971 4.5005
R20593 DVSS.n8014 DVSS.n1980 4.5005
R20594 DVSS.n1980 DVSS.n1971 4.5005
R20595 DVSS.n8014 DVSS.n1988 4.5005
R20596 DVSS.n1988 DVSS.n1971 4.5005
R20597 DVSS.n8014 DVSS.n1979 4.5005
R20598 DVSS.n1979 DVSS.n1971 4.5005
R20599 DVSS.n8014 DVSS.n1990 4.5005
R20600 DVSS.n1990 DVSS.n1971 4.5005
R20601 DVSS.n8014 DVSS.n1978 4.5005
R20602 DVSS.n1978 DVSS.n1971 4.5005
R20603 DVSS.n8014 DVSS.n1992 4.5005
R20604 DVSS.n1992 DVSS.n1971 4.5005
R20605 DVSS.n8014 DVSS.n1977 4.5005
R20606 DVSS.n1977 DVSS.n1971 4.5005
R20607 DVSS.n8014 DVSS.n8013 4.5005
R20608 DVSS.n8013 DVSS.n1976 4.5005
R20609 DVSS.n8013 DVSS.n1971 4.5005
R20610 DVSS.n1173 DVSS.n1162 4.5005
R20611 DVSS.n1173 DVSS.n1163 4.5005
R20612 DVSS.n8452 DVSS.n1173 4.5005
R20613 DVSS.n1170 DVSS.n1163 4.5005
R20614 DVSS.n8452 DVSS.n1170 4.5005
R20615 DVSS.n1176 DVSS.n1163 4.5005
R20616 DVSS.n8452 DVSS.n1176 4.5005
R20617 DVSS.n1169 DVSS.n1163 4.5005
R20618 DVSS.n8452 DVSS.n1169 4.5005
R20619 DVSS.n1163 DVSS.n1160 4.5005
R20620 DVSS.n1161 DVSS.n1160 4.5005
R20621 DVSS.n8452 DVSS.n1160 4.5005
R20622 DVSS.n8453 DVSS.n1162 4.5005
R20623 DVSS.n8453 DVSS.n1163 4.5005
R20624 DVSS.n8453 DVSS.n1161 4.5005
R20625 DVSS.n8453 DVSS.n8452 4.5005
R20626 DVSS.n8452 DVSS.n1156 4.5005
R20627 DVSS.n1161 DVSS.n1156 4.5005
R20628 DVSS.n1162 DVSS.n1156 4.5005
R20629 DVSS.n1167 DVSS.n1162 4.5005
R20630 DVSS.n8452 DVSS.n1167 4.5005
R20631 DVSS.n1179 DVSS.n1163 4.5005
R20632 DVSS.n8452 DVSS.n1179 4.5005
R20633 DVSS.n1165 DVSS.n1163 4.5005
R20634 DVSS.n8452 DVSS.n1165 4.5005
R20635 DVSS.n8451 DVSS.n1162 4.5005
R20636 DVSS.n8451 DVSS.n1163 4.5005
R20637 DVSS.n8452 DVSS.n8451 4.5005
R20638 DVSS.n2429 DVSS.n2413 4.5005
R20639 DVSS.n7419 DVSS.n2429 4.5005
R20640 DVSS.n2429 DVSS.n2417 4.5005
R20641 DVSS.n2432 DVSS.n2413 4.5005
R20642 DVSS.n7419 DVSS.n2432 4.5005
R20643 DVSS.n7419 DVSS.n2428 4.5005
R20644 DVSS.n7417 DVSS.n2428 4.5005
R20645 DVSS.n7419 DVSS.n2435 4.5005
R20646 DVSS.n7417 DVSS.n2435 4.5005
R20647 DVSS.n7419 DVSS.n2427 4.5005
R20648 DVSS.n7417 DVSS.n2427 4.5005
R20649 DVSS.n7419 DVSS.n2438 4.5005
R20650 DVSS.n7417 DVSS.n2438 4.5005
R20651 DVSS.n7419 DVSS.n2426 4.5005
R20652 DVSS.n7417 DVSS.n2426 4.5005
R20653 DVSS.n7419 DVSS.n2441 4.5005
R20654 DVSS.n7417 DVSS.n2441 4.5005
R20655 DVSS.n7419 DVSS.n2425 4.5005
R20656 DVSS.n7417 DVSS.n2425 4.5005
R20657 DVSS.n7419 DVSS.n2444 4.5005
R20658 DVSS.n7417 DVSS.n2444 4.5005
R20659 DVSS.n7419 DVSS.n2424 4.5005
R20660 DVSS.n7417 DVSS.n2424 4.5005
R20661 DVSS.n7419 DVSS.n2447 4.5005
R20662 DVSS.n7417 DVSS.n2447 4.5005
R20663 DVSS.n7419 DVSS.n2423 4.5005
R20664 DVSS.n7417 DVSS.n2423 4.5005
R20665 DVSS.n7419 DVSS.n2450 4.5005
R20666 DVSS.n7417 DVSS.n2450 4.5005
R20667 DVSS.n7419 DVSS.n2422 4.5005
R20668 DVSS.n7417 DVSS.n2422 4.5005
R20669 DVSS.n7419 DVSS.n2453 4.5005
R20670 DVSS.n7417 DVSS.n2453 4.5005
R20671 DVSS.n7419 DVSS.n2421 4.5005
R20672 DVSS.n7417 DVSS.n2421 4.5005
R20673 DVSS.n7419 DVSS.n2456 4.5005
R20674 DVSS.n7417 DVSS.n2456 4.5005
R20675 DVSS.n7419 DVSS.n2420 4.5005
R20676 DVSS.n7417 DVSS.n2420 4.5005
R20677 DVSS.n7419 DVSS.n2459 4.5005
R20678 DVSS.n7417 DVSS.n2459 4.5005
R20679 DVSS.n7419 DVSS.n2419 4.5005
R20680 DVSS.n7417 DVSS.n2419 4.5005
R20681 DVSS.n7419 DVSS.n2462 4.5005
R20682 DVSS.n7417 DVSS.n2462 4.5005
R20683 DVSS.n7419 DVSS.n2418 4.5005
R20684 DVSS.n7417 DVSS.n2418 4.5005
R20685 DVSS.n7419 DVSS.n7418 4.5005
R20686 DVSS.n7418 DVSS.n2417 4.5005
R20687 DVSS.n7418 DVSS.n7417 4.5005
R20688 DVSS.n2364 DVSS.n2348 4.5005
R20689 DVSS.n7454 DVSS.n2364 4.5005
R20690 DVSS.n7452 DVSS.n2364 4.5005
R20691 DVSS.n7454 DVSS.n2368 4.5005
R20692 DVSS.n7452 DVSS.n2368 4.5005
R20693 DVSS.n7454 DVSS.n2363 4.5005
R20694 DVSS.n7452 DVSS.n2363 4.5005
R20695 DVSS.n7454 DVSS.n2371 4.5005
R20696 DVSS.n7452 DVSS.n2371 4.5005
R20697 DVSS.n7454 DVSS.n2362 4.5005
R20698 DVSS.n7452 DVSS.n2362 4.5005
R20699 DVSS.n7454 DVSS.n2374 4.5005
R20700 DVSS.n7452 DVSS.n2374 4.5005
R20701 DVSS.n7454 DVSS.n2361 4.5005
R20702 DVSS.n7452 DVSS.n2361 4.5005
R20703 DVSS.n7454 DVSS.n2377 4.5005
R20704 DVSS.n7452 DVSS.n2377 4.5005
R20705 DVSS.n7454 DVSS.n2360 4.5005
R20706 DVSS.n7452 DVSS.n2360 4.5005
R20707 DVSS.n7454 DVSS.n2380 4.5005
R20708 DVSS.n7452 DVSS.n2380 4.5005
R20709 DVSS.n7454 DVSS.n2359 4.5005
R20710 DVSS.n7452 DVSS.n2359 4.5005
R20711 DVSS.n7454 DVSS.n2383 4.5005
R20712 DVSS.n7452 DVSS.n2383 4.5005
R20713 DVSS.n7454 DVSS.n2358 4.5005
R20714 DVSS.n7452 DVSS.n2358 4.5005
R20715 DVSS.n7454 DVSS.n2386 4.5005
R20716 DVSS.n7452 DVSS.n2386 4.5005
R20717 DVSS.n7454 DVSS.n2357 4.5005
R20718 DVSS.n7452 DVSS.n2357 4.5005
R20719 DVSS.n7454 DVSS.n2389 4.5005
R20720 DVSS.n7452 DVSS.n2389 4.5005
R20721 DVSS.n7454 DVSS.n2356 4.5005
R20722 DVSS.n7452 DVSS.n2356 4.5005
R20723 DVSS.n7454 DVSS.n2392 4.5005
R20724 DVSS.n7452 DVSS.n2392 4.5005
R20725 DVSS.n7454 DVSS.n2355 4.5005
R20726 DVSS.n7452 DVSS.n2355 4.5005
R20727 DVSS.n7454 DVSS.n2395 4.5005
R20728 DVSS.n7452 DVSS.n2395 4.5005
R20729 DVSS.n7454 DVSS.n2354 4.5005
R20730 DVSS.n7452 DVSS.n2354 4.5005
R20731 DVSS.n7454 DVSS.n2398 4.5005
R20732 DVSS.n7452 DVSS.n2398 4.5005
R20733 DVSS.n7454 DVSS.n2353 4.5005
R20734 DVSS.n7452 DVSS.n2353 4.5005
R20735 DVSS.n7453 DVSS.n2348 4.5005
R20736 DVSS.n7454 DVSS.n7453 4.5005
R20737 DVSS.n7453 DVSS.n7452 4.5005
R20738 DVSS.n7489 DVSS.n2322 4.5005
R20739 DVSS.n2322 DVSS.n2310 4.5005
R20740 DVSS.n7487 DVSS.n2322 4.5005
R20741 DVSS.n7489 DVSS.n2323 4.5005
R20742 DVSS.n2323 DVSS.n2310 4.5005
R20743 DVSS.n7487 DVSS.n2323 4.5005
R20744 DVSS.n7489 DVSS.n2321 4.5005
R20745 DVSS.n2321 DVSS.n2310 4.5005
R20746 DVSS.n7487 DVSS.n2321 4.5005
R20747 DVSS.n7489 DVSS.n2324 4.5005
R20748 DVSS.n2324 DVSS.n2310 4.5005
R20749 DVSS.n7487 DVSS.n2324 4.5005
R20750 DVSS.n7489 DVSS.n2320 4.5005
R20751 DVSS.n2320 DVSS.n2310 4.5005
R20752 DVSS.n7487 DVSS.n2320 4.5005
R20753 DVSS.n7489 DVSS.n2325 4.5005
R20754 DVSS.n2325 DVSS.n2310 4.5005
R20755 DVSS.n7487 DVSS.n2325 4.5005
R20756 DVSS.n7489 DVSS.n2319 4.5005
R20757 DVSS.n2319 DVSS.n2310 4.5005
R20758 DVSS.n7487 DVSS.n2319 4.5005
R20759 DVSS.n7489 DVSS.n2326 4.5005
R20760 DVSS.n2326 DVSS.n2310 4.5005
R20761 DVSS.n7487 DVSS.n2326 4.5005
R20762 DVSS.n7489 DVSS.n2318 4.5005
R20763 DVSS.n2318 DVSS.n2310 4.5005
R20764 DVSS.n7487 DVSS.n2318 4.5005
R20765 DVSS.n7489 DVSS.n2327 4.5005
R20766 DVSS.n2327 DVSS.n2310 4.5005
R20767 DVSS.n7487 DVSS.n2327 4.5005
R20768 DVSS.n7489 DVSS.n2317 4.5005
R20769 DVSS.n2317 DVSS.n2310 4.5005
R20770 DVSS.n7487 DVSS.n2317 4.5005
R20771 DVSS.n7489 DVSS.n2328 4.5005
R20772 DVSS.n2328 DVSS.n2310 4.5005
R20773 DVSS.n7487 DVSS.n2328 4.5005
R20774 DVSS.n7489 DVSS.n2316 4.5005
R20775 DVSS.n2316 DVSS.n2310 4.5005
R20776 DVSS.n7487 DVSS.n2316 4.5005
R20777 DVSS.n7489 DVSS.n2329 4.5005
R20778 DVSS.n2329 DVSS.n2310 4.5005
R20779 DVSS.n7487 DVSS.n2329 4.5005
R20780 DVSS.n7489 DVSS.n2315 4.5005
R20781 DVSS.n2315 DVSS.n2310 4.5005
R20782 DVSS.n7487 DVSS.n2315 4.5005
R20783 DVSS.n7489 DVSS.n2330 4.5005
R20784 DVSS.n2330 DVSS.n2310 4.5005
R20785 DVSS.n7487 DVSS.n2330 4.5005
R20786 DVSS.n7489 DVSS.n2314 4.5005
R20787 DVSS.n2314 DVSS.n2310 4.5005
R20788 DVSS.n7487 DVSS.n2314 4.5005
R20789 DVSS.n7489 DVSS.n2331 4.5005
R20790 DVSS.n2331 DVSS.n2310 4.5005
R20791 DVSS.n7487 DVSS.n2331 4.5005
R20792 DVSS.n7489 DVSS.n2313 4.5005
R20793 DVSS.n2313 DVSS.n2310 4.5005
R20794 DVSS.n7487 DVSS.n2313 4.5005
R20795 DVSS.n7489 DVSS.n2332 4.5005
R20796 DVSS.n2332 DVSS.n2310 4.5005
R20797 DVSS.n7487 DVSS.n2332 4.5005
R20798 DVSS.n7489 DVSS.n2312 4.5005
R20799 DVSS.n2312 DVSS.n2310 4.5005
R20800 DVSS.n7487 DVSS.n2312 4.5005
R20801 DVSS.n7489 DVSS.n2333 4.5005
R20802 DVSS.n2333 DVSS.n2310 4.5005
R20803 DVSS.n7487 DVSS.n2333 4.5005
R20804 DVSS.n7489 DVSS.n2311 4.5005
R20805 DVSS.n7487 DVSS.n2311 4.5005
R20806 DVSS.n7489 DVSS.n7488 4.5005
R20807 DVSS.n7488 DVSS.n7487 4.5005
R20808 DVSS.n7498 DVSS.n2292 4.5005
R20809 DVSS.n2292 DVSS.n2280 4.5005
R20810 DVSS.n7500 DVSS.n2292 4.5005
R20811 DVSS.n7498 DVSS.n2293 4.5005
R20812 DVSS.n2293 DVSS.n2280 4.5005
R20813 DVSS.n7500 DVSS.n2293 4.5005
R20814 DVSS.n7500 DVSS.n2291 4.5005
R20815 DVSS.n2291 DVSS.n2280 4.5005
R20816 DVSS.n7498 DVSS.n2291 4.5005
R20817 DVSS.n7500 DVSS.n2294 4.5005
R20818 DVSS.n2294 DVSS.n2280 4.5005
R20819 DVSS.n7498 DVSS.n2294 4.5005
R20820 DVSS.n7500 DVSS.n2290 4.5005
R20821 DVSS.n2290 DVSS.n2280 4.5005
R20822 DVSS.n7498 DVSS.n2290 4.5005
R20823 DVSS.n7500 DVSS.n2295 4.5005
R20824 DVSS.n2295 DVSS.n2280 4.5005
R20825 DVSS.n7498 DVSS.n2295 4.5005
R20826 DVSS.n7498 DVSS.n2289 4.5005
R20827 DVSS.n2289 DVSS.n2280 4.5005
R20828 DVSS.n7500 DVSS.n2289 4.5005
R20829 DVSS.n7498 DVSS.n2296 4.5005
R20830 DVSS.n2296 DVSS.n2280 4.5005
R20831 DVSS.n7500 DVSS.n2296 4.5005
R20832 DVSS.n7498 DVSS.n2288 4.5005
R20833 DVSS.n2288 DVSS.n2280 4.5005
R20834 DVSS.n7500 DVSS.n2288 4.5005
R20835 DVSS.n7500 DVSS.n2297 4.5005
R20836 DVSS.n2297 DVSS.n2280 4.5005
R20837 DVSS.n7498 DVSS.n2297 4.5005
R20838 DVSS.n7500 DVSS.n2287 4.5005
R20839 DVSS.n2287 DVSS.n2280 4.5005
R20840 DVSS.n7498 DVSS.n2287 4.5005
R20841 DVSS.n7500 DVSS.n2298 4.5005
R20842 DVSS.n2298 DVSS.n2280 4.5005
R20843 DVSS.n7498 DVSS.n2298 4.5005
R20844 DVSS.n7498 DVSS.n2286 4.5005
R20845 DVSS.n2286 DVSS.n2280 4.5005
R20846 DVSS.n7500 DVSS.n2286 4.5005
R20847 DVSS.n7498 DVSS.n2299 4.5005
R20848 DVSS.n2299 DVSS.n2280 4.5005
R20849 DVSS.n7500 DVSS.n2299 4.5005
R20850 DVSS.n7498 DVSS.n2285 4.5005
R20851 DVSS.n2285 DVSS.n2280 4.5005
R20852 DVSS.n7500 DVSS.n2285 4.5005
R20853 DVSS.n7498 DVSS.n2300 4.5005
R20854 DVSS.n2300 DVSS.n2280 4.5005
R20855 DVSS.n7500 DVSS.n2300 4.5005
R20856 DVSS.n7500 DVSS.n2284 4.5005
R20857 DVSS.n2284 DVSS.n2280 4.5005
R20858 DVSS.n7498 DVSS.n2284 4.5005
R20859 DVSS.n7500 DVSS.n2301 4.5005
R20860 DVSS.n2301 DVSS.n2280 4.5005
R20861 DVSS.n7498 DVSS.n2301 4.5005
R20862 DVSS.n7500 DVSS.n2283 4.5005
R20863 DVSS.n2283 DVSS.n2280 4.5005
R20864 DVSS.n7498 DVSS.n2283 4.5005
R20865 DVSS.n7498 DVSS.n2302 4.5005
R20866 DVSS.n2302 DVSS.n2280 4.5005
R20867 DVSS.n7500 DVSS.n2302 4.5005
R20868 DVSS.n7498 DVSS.n2282 4.5005
R20869 DVSS.n2282 DVSS.n2280 4.5005
R20870 DVSS.n7500 DVSS.n2282 4.5005
R20871 DVSS.n7498 DVSS.n2303 4.5005
R20872 DVSS.n2303 DVSS.n2280 4.5005
R20873 DVSS.n7500 DVSS.n2303 4.5005
R20874 DVSS.n7500 DVSS.n2281 4.5005
R20875 DVSS.n7498 DVSS.n2281 4.5005
R20876 DVSS.n7500 DVSS.n7499 4.5005
R20877 DVSS.n7499 DVSS.n7498 4.5005
R20878 DVSS.n7558 DVSS.n2250 4.5005
R20879 DVSS.n2250 DVSS.n2238 4.5005
R20880 DVSS.n7556 DVSS.n2250 4.5005
R20881 DVSS.n7532 DVSS.n2238 4.5005
R20882 DVSS.n7556 DVSS.n7532 4.5005
R20883 DVSS.n2264 DVSS.n2238 4.5005
R20884 DVSS.n7556 DVSS.n2264 4.5005
R20885 DVSS.n7533 DVSS.n2238 4.5005
R20886 DVSS.n7556 DVSS.n7533 4.5005
R20887 DVSS.n2263 DVSS.n2238 4.5005
R20888 DVSS.n7556 DVSS.n2263 4.5005
R20889 DVSS.n7534 DVSS.n2238 4.5005
R20890 DVSS.n7556 DVSS.n7534 4.5005
R20891 DVSS.n2262 DVSS.n2238 4.5005
R20892 DVSS.n7556 DVSS.n2262 4.5005
R20893 DVSS.n7535 DVSS.n2238 4.5005
R20894 DVSS.n7556 DVSS.n7535 4.5005
R20895 DVSS.n2261 DVSS.n2238 4.5005
R20896 DVSS.n7556 DVSS.n2261 4.5005
R20897 DVSS.n7536 DVSS.n2238 4.5005
R20898 DVSS.n7556 DVSS.n7536 4.5005
R20899 DVSS.n2260 DVSS.n2238 4.5005
R20900 DVSS.n7556 DVSS.n2260 4.5005
R20901 DVSS.n7537 DVSS.n2238 4.5005
R20902 DVSS.n7556 DVSS.n7537 4.5005
R20903 DVSS.n2259 DVSS.n2238 4.5005
R20904 DVSS.n7556 DVSS.n2259 4.5005
R20905 DVSS.n7538 DVSS.n2238 4.5005
R20906 DVSS.n7556 DVSS.n7538 4.5005
R20907 DVSS.n2258 DVSS.n2238 4.5005
R20908 DVSS.n7556 DVSS.n2258 4.5005
R20909 DVSS.n7539 DVSS.n2238 4.5005
R20910 DVSS.n7556 DVSS.n7539 4.5005
R20911 DVSS.n2257 DVSS.n2238 4.5005
R20912 DVSS.n7556 DVSS.n2257 4.5005
R20913 DVSS.n7540 DVSS.n2238 4.5005
R20914 DVSS.n7556 DVSS.n7540 4.5005
R20915 DVSS.n2256 DVSS.n2238 4.5005
R20916 DVSS.n7556 DVSS.n2256 4.5005
R20917 DVSS.n7541 DVSS.n2238 4.5005
R20918 DVSS.n7556 DVSS.n7541 4.5005
R20919 DVSS.n2255 DVSS.n2238 4.5005
R20920 DVSS.n7556 DVSS.n2255 4.5005
R20921 DVSS.n7555 DVSS.n2238 4.5005
R20922 DVSS.n7556 DVSS.n7555 4.5005
R20923 DVSS.n2254 DVSS.n2238 4.5005
R20924 DVSS.n7556 DVSS.n2254 4.5005
R20925 DVSS.n7558 DVSS.n7557 4.5005
R20926 DVSS.n7557 DVSS.n2238 4.5005
R20927 DVSS.n7557 DVSS.n7556 4.5005
R20928 DVSS.n7616 DVSS.n2208 4.5005
R20929 DVSS.n2208 DVSS.n2196 4.5005
R20930 DVSS.n7614 DVSS.n2208 4.5005
R20931 DVSS.n7590 DVSS.n2196 4.5005
R20932 DVSS.n7614 DVSS.n7590 4.5005
R20933 DVSS.n2222 DVSS.n2196 4.5005
R20934 DVSS.n7614 DVSS.n2222 4.5005
R20935 DVSS.n7591 DVSS.n2196 4.5005
R20936 DVSS.n7614 DVSS.n7591 4.5005
R20937 DVSS.n2221 DVSS.n2196 4.5005
R20938 DVSS.n7614 DVSS.n2221 4.5005
R20939 DVSS.n7592 DVSS.n2196 4.5005
R20940 DVSS.n7614 DVSS.n7592 4.5005
R20941 DVSS.n2220 DVSS.n2196 4.5005
R20942 DVSS.n7614 DVSS.n2220 4.5005
R20943 DVSS.n7593 DVSS.n2196 4.5005
R20944 DVSS.n7614 DVSS.n7593 4.5005
R20945 DVSS.n2219 DVSS.n2196 4.5005
R20946 DVSS.n7614 DVSS.n2219 4.5005
R20947 DVSS.n7594 DVSS.n2196 4.5005
R20948 DVSS.n7614 DVSS.n7594 4.5005
R20949 DVSS.n2218 DVSS.n2196 4.5005
R20950 DVSS.n7614 DVSS.n2218 4.5005
R20951 DVSS.n7595 DVSS.n2196 4.5005
R20952 DVSS.n7614 DVSS.n7595 4.5005
R20953 DVSS.n2217 DVSS.n2196 4.5005
R20954 DVSS.n7614 DVSS.n2217 4.5005
R20955 DVSS.n7596 DVSS.n2196 4.5005
R20956 DVSS.n7614 DVSS.n7596 4.5005
R20957 DVSS.n2216 DVSS.n2196 4.5005
R20958 DVSS.n7614 DVSS.n2216 4.5005
R20959 DVSS.n7597 DVSS.n2196 4.5005
R20960 DVSS.n7614 DVSS.n7597 4.5005
R20961 DVSS.n2215 DVSS.n2196 4.5005
R20962 DVSS.n7614 DVSS.n2215 4.5005
R20963 DVSS.n7598 DVSS.n2196 4.5005
R20964 DVSS.n7614 DVSS.n7598 4.5005
R20965 DVSS.n2214 DVSS.n2196 4.5005
R20966 DVSS.n7614 DVSS.n2214 4.5005
R20967 DVSS.n7599 DVSS.n2196 4.5005
R20968 DVSS.n7614 DVSS.n7599 4.5005
R20969 DVSS.n2213 DVSS.n2196 4.5005
R20970 DVSS.n7614 DVSS.n2213 4.5005
R20971 DVSS.n7613 DVSS.n2196 4.5005
R20972 DVSS.n7614 DVSS.n7613 4.5005
R20973 DVSS.n2212 DVSS.n2196 4.5005
R20974 DVSS.n7614 DVSS.n2212 4.5005
R20975 DVSS.n7616 DVSS.n7615 4.5005
R20976 DVSS.n7615 DVSS.n2196 4.5005
R20977 DVSS.n7615 DVSS.n7614 4.5005
R20978 DVSS.n7399 DVSS.n2485 4.5005
R20979 DVSS.n2485 DVSS.n2473 4.5005
R20980 DVSS.n7397 DVSS.n2485 4.5005
R20981 DVSS.n7399 DVSS.n2489 4.5005
R20982 DVSS.n7397 DVSS.n2489 4.5005
R20983 DVSS.n7399 DVSS.n2484 4.5005
R20984 DVSS.n7397 DVSS.n2484 4.5005
R20985 DVSS.n7399 DVSS.n2492 4.5005
R20986 DVSS.n7397 DVSS.n2492 4.5005
R20987 DVSS.n7399 DVSS.n2483 4.5005
R20988 DVSS.n7397 DVSS.n2483 4.5005
R20989 DVSS.n7399 DVSS.n2495 4.5005
R20990 DVSS.n7397 DVSS.n2495 4.5005
R20991 DVSS.n7399 DVSS.n2482 4.5005
R20992 DVSS.n7397 DVSS.n2482 4.5005
R20993 DVSS.n7399 DVSS.n2498 4.5005
R20994 DVSS.n7397 DVSS.n2498 4.5005
R20995 DVSS.n7399 DVSS.n2481 4.5005
R20996 DVSS.n7397 DVSS.n2481 4.5005
R20997 DVSS.n7399 DVSS.n2501 4.5005
R20998 DVSS.n7397 DVSS.n2501 4.5005
R20999 DVSS.n7399 DVSS.n2480 4.5005
R21000 DVSS.n7397 DVSS.n2480 4.5005
R21001 DVSS.n7399 DVSS.n2504 4.5005
R21002 DVSS.n7397 DVSS.n2504 4.5005
R21003 DVSS.n7399 DVSS.n2479 4.5005
R21004 DVSS.n7397 DVSS.n2479 4.5005
R21005 DVSS.n7399 DVSS.n2507 4.5005
R21006 DVSS.n7397 DVSS.n2507 4.5005
R21007 DVSS.n7399 DVSS.n2478 4.5005
R21008 DVSS.n7397 DVSS.n2478 4.5005
R21009 DVSS.n7399 DVSS.n2510 4.5005
R21010 DVSS.n7397 DVSS.n2510 4.5005
R21011 DVSS.n7399 DVSS.n2477 4.5005
R21012 DVSS.n7397 DVSS.n2477 4.5005
R21013 DVSS.n7399 DVSS.n2513 4.5005
R21014 DVSS.n7397 DVSS.n2513 4.5005
R21015 DVSS.n7399 DVSS.n2476 4.5005
R21016 DVSS.n7397 DVSS.n2476 4.5005
R21017 DVSS.n7399 DVSS.n2516 4.5005
R21018 DVSS.n7397 DVSS.n2516 4.5005
R21019 DVSS.n7399 DVSS.n2475 4.5005
R21020 DVSS.n7397 DVSS.n2475 4.5005
R21021 DVSS.n7399 DVSS.n2519 4.5005
R21022 DVSS.n7397 DVSS.n2519 4.5005
R21023 DVSS.n7399 DVSS.n2474 4.5005
R21024 DVSS.n7397 DVSS.n2474 4.5005
R21025 DVSS.n7399 DVSS.n7398 4.5005
R21026 DVSS.n7398 DVSS.n2473 4.5005
R21027 DVSS.n7398 DVSS.n7397 4.5005
R21028 DVSS.n8034 DVSS.n1958 4.5005
R21029 DVSS.n8037 DVSS.n1958 4.5005
R21030 DVSS.n1958 DVSS.n1945 4.5005
R21031 DVSS.n8037 DVSS.n1955 4.5005
R21032 DVSS.n1955 DVSS.n1945 4.5005
R21033 DVSS.n8037 DVSS.n1960 4.5005
R21034 DVSS.n1960 DVSS.n1945 4.5005
R21035 DVSS.n8037 DVSS.n1954 4.5005
R21036 DVSS.n1954 DVSS.n1945 4.5005
R21037 DVSS.n8037 DVSS.n1962 4.5005
R21038 DVSS.n1962 DVSS.n1945 4.5005
R21039 DVSS.n8037 DVSS.n1953 4.5005
R21040 DVSS.n1953 DVSS.n1945 4.5005
R21041 DVSS.n8037 DVSS.n1964 4.5005
R21042 DVSS.n1964 DVSS.n1945 4.5005
R21043 DVSS.n8037 DVSS.n1952 4.5005
R21044 DVSS.n1952 DVSS.n1945 4.5005
R21045 DVSS.n8037 DVSS.n1966 4.5005
R21046 DVSS.n1966 DVSS.n1945 4.5005
R21047 DVSS.n8037 DVSS.n1951 4.5005
R21048 DVSS.n1951 DVSS.n1945 4.5005
R21049 DVSS.n8037 DVSS.n8036 4.5005
R21050 DVSS.n8036 DVSS.n1950 4.5005
R21051 DVSS.n8036 DVSS.n1945 4.5005
R21052 DVSS.n7063 DVSS.n6667 4.5005
R21053 DVSS.n7063 DVSS.n6668 4.5005
R21054 DVSS.n7063 DVSS.n7062 4.5005
R21055 DVSS.n6674 DVSS.n6668 4.5005
R21056 DVSS.n7062 DVSS.n6674 4.5005
R21057 DVSS.n6677 DVSS.n6668 4.5005
R21058 DVSS.n7062 DVSS.n6677 4.5005
R21059 DVSS.n6673 DVSS.n6668 4.5005
R21060 DVSS.n7062 DVSS.n6673 4.5005
R21061 DVSS.n6679 DVSS.n6668 4.5005
R21062 DVSS.n7062 DVSS.n6679 4.5005
R21063 DVSS.n6672 DVSS.n6668 4.5005
R21064 DVSS.n7062 DVSS.n6672 4.5005
R21065 DVSS.n6681 DVSS.n6668 4.5005
R21066 DVSS.n7062 DVSS.n6681 4.5005
R21067 DVSS.n6671 DVSS.n6668 4.5005
R21068 DVSS.n7062 DVSS.n6671 4.5005
R21069 DVSS.n6683 DVSS.n6668 4.5005
R21070 DVSS.n7062 DVSS.n6683 4.5005
R21071 DVSS.n6670 DVSS.n6668 4.5005
R21072 DVSS.n7062 DVSS.n6670 4.5005
R21073 DVSS.n7061 DVSS.n6668 4.5005
R21074 DVSS.n7061 DVSS.n6689 4.5005
R21075 DVSS.n7062 DVSS.n7061 4.5005
R21076 DVSS.n5834 DVSS.n3049 4.5005
R21077 DVSS.n5837 DVSS.n3049 4.5005
R21078 DVSS.n5834 DVSS.n3047 4.5005
R21079 DVSS.n5837 DVSS.n3047 4.5005
R21080 DVSS.n5834 DVSS.n3050 4.5005
R21081 DVSS.n5837 DVSS.n3050 4.5005
R21082 DVSS.n5834 DVSS.n3046 4.5005
R21083 DVSS.n5837 DVSS.n3046 4.5005
R21084 DVSS.n5837 DVSS.n5836 4.5005
R21085 DVSS.n5834 DVSS.n5833 4.5005
R21086 DVSS.n5832 DVSS.n5831 4.5005
R21087 DVSS.n5831 DVSS.n3059 4.5005
R21088 DVSS.n5831 DVSS.n3063 4.5005
R21089 DVSS.n5829 DVSS.n3063 4.5005
R21090 DVSS.n5831 DVSS.n3058 4.5005
R21091 DVSS.n5829 DVSS.n3058 4.5005
R21092 DVSS.n5831 DVSS.n3064 4.5005
R21093 DVSS.n5829 DVSS.n3064 4.5005
R21094 DVSS.n5831 DVSS.n3057 4.5005
R21095 DVSS.n5829 DVSS.n3057 4.5005
R21096 DVSS.n5831 DVSS.n5830 4.5005
R21097 DVSS.n5830 DVSS.n5829 4.5005
R21098 DVSS.n4260 DVSS.n4217 4.5005
R21099 DVSS.n4217 DVSS.n4215 4.5005
R21100 DVSS.n4258 DVSS.n4217 4.5005
R21101 DVSS.n4228 DVSS.n4215 4.5005
R21102 DVSS.n4258 DVSS.n4228 4.5005
R21103 DVSS.n4254 DVSS.n4215 4.5005
R21104 DVSS.n4258 DVSS.n4254 4.5005
R21105 DVSS.n4226 DVSS.n4215 4.5005
R21106 DVSS.n4258 DVSS.n4226 4.5005
R21107 DVSS.n4256 DVSS.n4215 4.5005
R21108 DVSS.n4258 DVSS.n4256 4.5005
R21109 DVSS.n4225 DVSS.n4215 4.5005
R21110 DVSS.n4258 DVSS.n4225 4.5005
R21111 DVSS.n4257 DVSS.n4215 4.5005
R21112 DVSS.n4257 DVSS.n4223 4.5005
R21113 DVSS.n4258 DVSS.n4257 4.5005
R21114 DVSS.n4260 DVSS.n3862 4.5005
R21115 DVSS.n4215 DVSS.n3862 4.5005
R21116 DVSS.n4223 DVSS.n3862 4.5005
R21117 DVSS.n4258 DVSS.n3862 4.5005
R21118 DVSS.n4260 DVSS.n3864 4.5005
R21119 DVSS.n4215 DVSS.n3864 4.5005
R21120 DVSS.n4223 DVSS.n3864 4.5005
R21121 DVSS.n4258 DVSS.n3864 4.5005
R21122 DVSS.n4260 DVSS.n4216 4.5005
R21123 DVSS.n4216 DVSS.n4215 4.5005
R21124 DVSS.n4223 DVSS.n4216 4.5005
R21125 DVSS.n4258 DVSS.n4216 4.5005
R21126 DVSS.n4260 DVSS.n4259 4.5005
R21127 DVSS.n4259 DVSS.n4215 4.5005
R21128 DVSS.n4259 DVSS.n4223 4.5005
R21129 DVSS.n4259 DVSS.n4258 4.5005
R21130 DVSS.n4519 DVSS.n3818 4.5005
R21131 DVSS.n3818 DVSS.n3815 4.5005
R21132 DVSS.n4517 DVSS.n3818 4.5005
R21133 DVSS.n3825 DVSS.n3818 4.5005
R21134 DVSS.n4519 DVSS.n3819 4.5005
R21135 DVSS.n3819 DVSS.n3815 4.5005
R21136 DVSS.n3825 DVSS.n3819 4.5005
R21137 DVSS.n4514 DVSS.n3815 4.5005
R21138 DVSS.n4514 DVSS.n3825 4.5005
R21139 DVSS.n4512 DVSS.n3815 4.5005
R21140 DVSS.n4512 DVSS.n3825 4.5005
R21141 DVSS.n4511 DVSS.n3815 4.5005
R21142 DVSS.n4511 DVSS.n3825 4.5005
R21143 DVSS.n4509 DVSS.n3815 4.5005
R21144 DVSS.n4509 DVSS.n3825 4.5005
R21145 DVSS.n4519 DVSS.n3817 4.5005
R21146 DVSS.n3817 DVSS.n3815 4.5005
R21147 DVSS.n3825 DVSS.n3817 4.5005
R21148 DVSS.n3825 DVSS.n3823 4.5005
R21149 DVSS.n4517 DVSS.n3823 4.5005
R21150 DVSS.n4519 DVSS.n3823 4.5005
R21151 DVSS.n3825 DVSS.n3816 4.5005
R21152 DVSS.n4517 DVSS.n3816 4.5005
R21153 DVSS.n4519 DVSS.n3816 4.5005
R21154 DVSS.n4519 DVSS.n4518 4.5005
R21155 DVSS.n4518 DVSS.n3815 4.5005
R21156 DVSS.n4518 DVSS.n3825 4.5005
R21157 DVSS.n4518 DVSS.n4517 4.5005
R21158 DVSS.n4589 DVSS.n3800 4.5005
R21159 DVSS.n4589 DVSS.n3801 4.5005
R21160 DVSS.n4589 DVSS.n3799 4.5005
R21161 DVSS.n4589 DVSS.n4588 4.5005
R21162 DVSS.n4581 DVSS.n3800 4.5005
R21163 DVSS.n4581 DVSS.n3801 4.5005
R21164 DVSS.n4588 DVSS.n4581 4.5005
R21165 DVSS.n3807 DVSS.n3801 4.5005
R21166 DVSS.n4588 DVSS.n3807 4.5005
R21167 DVSS.n4584 DVSS.n3801 4.5005
R21168 DVSS.n4588 DVSS.n4584 4.5005
R21169 DVSS.n3806 DVSS.n3801 4.5005
R21170 DVSS.n4588 DVSS.n3806 4.5005
R21171 DVSS.n4587 DVSS.n3801 4.5005
R21172 DVSS.n4588 DVSS.n4587 4.5005
R21173 DVSS.n3805 DVSS.n3800 4.5005
R21174 DVSS.n3805 DVSS.n3801 4.5005
R21175 DVSS.n4588 DVSS.n3805 4.5005
R21176 DVSS.n4588 DVSS.n3793 4.5005
R21177 DVSS.n3799 DVSS.n3793 4.5005
R21178 DVSS.n3800 DVSS.n3793 4.5005
R21179 DVSS.n4588 DVSS.n3804 4.5005
R21180 DVSS.n3804 DVSS.n3799 4.5005
R21181 DVSS.n3804 DVSS.n3800 4.5005
R21182 DVSS.n3800 DVSS.n3796 4.5005
R21183 DVSS.n3801 DVSS.n3796 4.5005
R21184 DVSS.n4588 DVSS.n3796 4.5005
R21185 DVSS.n3799 DVSS.n3796 4.5005
R21186 DVSS.n3734 DVSS.n3728 4.5005
R21187 DVSS.n3734 DVSS.n3729 4.5005
R21188 DVSS.n4782 DVSS.n3734 4.5005
R21189 DVSS.n4784 DVSS.n3734 4.5005
R21190 DVSS.n3736 DVSS.n3728 4.5005
R21191 DVSS.n3736 DVSS.n3729 4.5005
R21192 DVSS.n4784 DVSS.n3736 4.5005
R21193 DVSS.n3733 DVSS.n3729 4.5005
R21194 DVSS.n4784 DVSS.n3733 4.5005
R21195 DVSS.n3738 DVSS.n3729 4.5005
R21196 DVSS.n4784 DVSS.n3738 4.5005
R21197 DVSS.n3732 DVSS.n3729 4.5005
R21198 DVSS.n4784 DVSS.n3732 4.5005
R21199 DVSS.n3740 DVSS.n3729 4.5005
R21200 DVSS.n4784 DVSS.n3740 4.5005
R21201 DVSS.n4785 DVSS.n3728 4.5005
R21202 DVSS.n4785 DVSS.n3729 4.5005
R21203 DVSS.n4785 DVSS.n4784 4.5005
R21204 DVSS.n4784 DVSS.n3742 4.5005
R21205 DVSS.n4782 DVSS.n3742 4.5005
R21206 DVSS.n3742 DVSS.n3728 4.5005
R21207 DVSS.n4784 DVSS.n3731 4.5005
R21208 DVSS.n4782 DVSS.n3731 4.5005
R21209 DVSS.n3731 DVSS.n3728 4.5005
R21210 DVSS.n4783 DVSS.n3728 4.5005
R21211 DVSS.n4783 DVSS.n3729 4.5005
R21212 DVSS.n4784 DVSS.n4783 4.5005
R21213 DVSS.n4783 DVSS.n4782 4.5005
R21214 DVSS.n4755 DVSS.n3774 4.5005
R21215 DVSS.n3783 DVSS.n3774 4.5005
R21216 DVSS.n4757 DVSS.n3774 4.5005
R21217 DVSS.n4755 DVSS.n3776 4.5005
R21218 DVSS.n4757 DVSS.n3776 4.5005
R21219 DVSS.n4755 DVSS.n3773 4.5005
R21220 DVSS.n4757 DVSS.n3773 4.5005
R21221 DVSS.n4755 DVSS.n3777 4.5005
R21222 DVSS.n3783 DVSS.n3777 4.5005
R21223 DVSS.n4757 DVSS.n3777 4.5005
R21224 DVSS.n4755 DVSS.n3772 4.5005
R21225 DVSS.n3783 DVSS.n3772 4.5005
R21226 DVSS.n4757 DVSS.n3772 4.5005
R21227 DVSS.n4755 DVSS.n3778 4.5005
R21228 DVSS.n3783 DVSS.n3778 4.5005
R21229 DVSS.n4757 DVSS.n3778 4.5005
R21230 DVSS.n4755 DVSS.n3771 4.5005
R21231 DVSS.n3783 DVSS.n3771 4.5005
R21232 DVSS.n4757 DVSS.n3771 4.5005
R21233 DVSS.n4757 DVSS.n3779 4.5005
R21234 DVSS.n4755 DVSS.n3779 4.5005
R21235 DVSS.n4757 DVSS.n3770 4.5005
R21236 DVSS.n4755 DVSS.n3770 4.5005
R21237 DVSS.n4756 DVSS.n4755 4.5005
R21238 DVSS.n4756 DVSS.n3783 4.5005
R21239 DVSS.n4757 DVSS.n4756 4.5005
R21240 DVSS.n4746 DVSS.n4621 4.5005
R21241 DVSS.n4749 DVSS.n4621 4.5005
R21242 DVSS.n4621 DVSS.n4616 4.5005
R21243 DVSS.n4746 DVSS.n4745 4.5005
R21244 DVSS.n4745 DVSS.n4616 4.5005
R21245 DVSS.n4746 DVSS.n4704 4.5005
R21246 DVSS.n4704 DVSS.n4616 4.5005
R21247 DVSS.n4746 DVSS.n4623 4.5005
R21248 DVSS.n4749 DVSS.n4623 4.5005
R21249 DVSS.n4623 DVSS.n4616 4.5005
R21250 DVSS.n4746 DVSS.n4618 4.5005
R21251 DVSS.n4749 DVSS.n4618 4.5005
R21252 DVSS.n4618 DVSS.n4616 4.5005
R21253 DVSS.n4746 DVSS.n4624 4.5005
R21254 DVSS.n4749 DVSS.n4624 4.5005
R21255 DVSS.n4624 DVSS.n4616 4.5005
R21256 DVSS.n4746 DVSS.n4617 4.5005
R21257 DVSS.n4749 DVSS.n4617 4.5005
R21258 DVSS.n4617 DVSS.n4616 4.5005
R21259 DVSS.n4616 DVSS.n2762 4.5005
R21260 DVSS.n4746 DVSS.n2762 4.5005
R21261 DVSS.n4747 DVSS.n4616 4.5005
R21262 DVSS.n4747 DVSS.n4746 4.5005
R21263 DVSS.n4746 DVSS.n2764 4.5005
R21264 DVSS.n4749 DVSS.n2764 4.5005
R21265 DVSS.n4616 DVSS.n2764 4.5005
R21266 DVSS.n2781 DVSS.n2778 4.5005
R21267 DVSS.n2782 DVSS.n2778 4.5005
R21268 DVSS.n6000 DVSS.n2778 4.5005
R21269 DVSS.n6003 DVSS.n2778 4.5005
R21270 DVSS.n6004 DVSS.n2781 4.5005
R21271 DVSS.n6004 DVSS.n2782 4.5005
R21272 DVSS.n6004 DVSS.n6003 4.5005
R21273 DVSS.n2788 DVSS.n2782 4.5005
R21274 DVSS.n6003 DVSS.n2788 4.5005
R21275 DVSS.n2791 DVSS.n2782 4.5005
R21276 DVSS.n6003 DVSS.n2791 4.5005
R21277 DVSS.n2787 DVSS.n2782 4.5005
R21278 DVSS.n6003 DVSS.n2787 4.5005
R21279 DVSS.n6002 DVSS.n2782 4.5005
R21280 DVSS.n6003 DVSS.n6002 4.5005
R21281 DVSS.n2786 DVSS.n2781 4.5005
R21282 DVSS.n2786 DVSS.n2782 4.5005
R21283 DVSS.n6003 DVSS.n2786 4.5005
R21284 DVSS.n6003 DVSS.n2770 4.5005
R21285 DVSS.n6000 DVSS.n2770 4.5005
R21286 DVSS.n2781 DVSS.n2770 4.5005
R21287 DVSS.n6003 DVSS.n2785 4.5005
R21288 DVSS.n6000 DVSS.n2785 4.5005
R21289 DVSS.n2785 DVSS.n2781 4.5005
R21290 DVSS.n2781 DVSS.n2773 4.5005
R21291 DVSS.n2782 DVSS.n2773 4.5005
R21292 DVSS.n6003 DVSS.n2773 4.5005
R21293 DVSS.n6000 DVSS.n2773 4.5005
R21294 DVSS.n2830 DVSS.n2821 4.5005
R21295 DVSS.n2833 DVSS.n2821 4.5005
R21296 DVSS.n5973 DVSS.n2821 4.5005
R21297 DVSS.n5975 DVSS.n2821 4.5005
R21298 DVSS.n2830 DVSS.n2823 4.5005
R21299 DVSS.n2833 DVSS.n2823 4.5005
R21300 DVSS.n5975 DVSS.n2823 4.5005
R21301 DVSS.n2833 DVSS.n2820 4.5005
R21302 DVSS.n5975 DVSS.n2820 4.5005
R21303 DVSS.n2833 DVSS.n2824 4.5005
R21304 DVSS.n5975 DVSS.n2824 4.5005
R21305 DVSS.n2833 DVSS.n2819 4.5005
R21306 DVSS.n5975 DVSS.n2819 4.5005
R21307 DVSS.n2833 DVSS.n2825 4.5005
R21308 DVSS.n5975 DVSS.n2825 4.5005
R21309 DVSS.n2830 DVSS.n2818 4.5005
R21310 DVSS.n2833 DVSS.n2818 4.5005
R21311 DVSS.n5975 DVSS.n2818 4.5005
R21312 DVSS.n5975 DVSS.n2826 4.5005
R21313 DVSS.n5973 DVSS.n2826 4.5005
R21314 DVSS.n2830 DVSS.n2826 4.5005
R21315 DVSS.n5975 DVSS.n2817 4.5005
R21316 DVSS.n5973 DVSS.n2817 4.5005
R21317 DVSS.n2830 DVSS.n2817 4.5005
R21318 DVSS.n5974 DVSS.n2830 4.5005
R21319 DVSS.n5974 DVSS.n2833 4.5005
R21320 DVSS.n5975 DVSS.n5974 4.5005
R21321 DVSS.n5974 DVSS.n5973 4.5005
R21322 DVSS.n2863 DVSS.n2852 4.5005
R21323 DVSS.n2865 DVSS.n2852 4.5005
R21324 DVSS.n5958 DVSS.n2852 4.5005
R21325 DVSS.n5960 DVSS.n2852 4.5005
R21326 DVSS.n2865 DVSS.n2854 4.5005
R21327 DVSS.n5958 DVSS.n2854 4.5005
R21328 DVSS.n5960 DVSS.n2854 4.5005
R21329 DVSS.n2865 DVSS.n2851 4.5005
R21330 DVSS.n5960 DVSS.n2851 4.5005
R21331 DVSS.n2865 DVSS.n2855 4.5005
R21332 DVSS.n5960 DVSS.n2855 4.5005
R21333 DVSS.n2865 DVSS.n2850 4.5005
R21334 DVSS.n5960 DVSS.n2850 4.5005
R21335 DVSS.n2865 DVSS.n2856 4.5005
R21336 DVSS.n5960 DVSS.n2856 4.5005
R21337 DVSS.n2865 DVSS.n2849 4.5005
R21338 DVSS.n5958 DVSS.n2849 4.5005
R21339 DVSS.n5960 DVSS.n2849 4.5005
R21340 DVSS.n4963 DVSS.n3599 4.5005
R21341 DVSS.n4963 DVSS.n3600 4.5005
R21342 DVSS.n4972 DVSS.n4963 4.5005
R21343 DVSS.n3604 DVSS.n3600 4.5005
R21344 DVSS.n4972 DVSS.n3604 4.5005
R21345 DVSS.n4966 DVSS.n3600 4.5005
R21346 DVSS.n4972 DVSS.n4966 4.5005
R21347 DVSS.n3603 DVSS.n3600 4.5005
R21348 DVSS.n4972 DVSS.n3603 4.5005
R21349 DVSS.n4969 DVSS.n3600 4.5005
R21350 DVSS.n4972 DVSS.n4969 4.5005
R21351 DVSS.n3602 DVSS.n3600 4.5005
R21352 DVSS.n4972 DVSS.n3602 4.5005
R21353 DVSS.n4971 DVSS.n3600 4.5005
R21354 DVSS.n4971 DVSS.n3598 4.5005
R21355 DVSS.n4972 DVSS.n4971 4.5005
R21356 DVSS.n3599 DVSS.n3595 4.5005
R21357 DVSS.n3600 DVSS.n3595 4.5005
R21358 DVSS.n3598 DVSS.n3595 4.5005
R21359 DVSS.n4972 DVSS.n3595 4.5005
R21360 DVSS.n3599 DVSS.n3597 4.5005
R21361 DVSS.n3600 DVSS.n3597 4.5005
R21362 DVSS.n3598 DVSS.n3597 4.5005
R21363 DVSS.n4972 DVSS.n3597 4.5005
R21364 DVSS.n4973 DVSS.n3599 4.5005
R21365 DVSS.n4973 DVSS.n3600 4.5005
R21366 DVSS.n4973 DVSS.n3598 4.5005
R21367 DVSS.n4973 DVSS.n4972 4.5005
R21368 DVSS.n3599 DVSS.n3588 4.5005
R21369 DVSS.n3600 DVSS.n3588 4.5005
R21370 DVSS.n3598 DVSS.n3588 4.5005
R21371 DVSS.n4972 DVSS.n3588 4.5005
R21372 DVSS.n5349 DVSS.n3387 4.5005
R21373 DVSS.n3387 DVSS.n3379 4.5005
R21374 DVSS.n3387 DVSS.n3378 4.5005
R21375 DVSS.n5353 DVSS.n3387 4.5005
R21376 DVSS.n5349 DVSS.n3385 4.5005
R21377 DVSS.n3385 DVSS.n3379 4.5005
R21378 DVSS.n3385 DVSS.n3378 4.5005
R21379 DVSS.n5353 DVSS.n3385 4.5005
R21380 DVSS.n5349 DVSS.n3388 4.5005
R21381 DVSS.n3388 DVSS.n3379 4.5005
R21382 DVSS.n3388 DVSS.n3378 4.5005
R21383 DVSS.n5353 DVSS.n3388 4.5005
R21384 DVSS.n5349 DVSS.n3384 4.5005
R21385 DVSS.n3384 DVSS.n3379 4.5005
R21386 DVSS.n3384 DVSS.n3378 4.5005
R21387 DVSS.n5353 DVSS.n3384 4.5005
R21388 DVSS.n5349 DVSS.n3390 4.5005
R21389 DVSS.n3390 DVSS.n3379 4.5005
R21390 DVSS.n5353 DVSS.n3390 4.5005
R21391 DVSS.n3383 DVSS.n3379 4.5005
R21392 DVSS.n5353 DVSS.n3383 4.5005
R21393 DVSS.n3392 DVSS.n3379 4.5005
R21394 DVSS.n5353 DVSS.n3392 4.5005
R21395 DVSS.n3382 DVSS.n3379 4.5005
R21396 DVSS.n5353 DVSS.n3382 4.5005
R21397 DVSS.n5352 DVSS.n3379 4.5005
R21398 DVSS.n5353 DVSS.n5352 4.5005
R21399 DVSS.n3381 DVSS.n3379 4.5005
R21400 DVSS.n5353 DVSS.n3381 4.5005
R21401 DVSS.n5354 DVSS.n3379 4.5005
R21402 DVSS.n5354 DVSS.n3378 4.5005
R21403 DVSS.n5354 DVSS.n5353 4.5005
R21404 DVSS.n5366 DVSS.n5355 4.5005
R21405 DVSS.n5355 DVSS.n3371 4.5005
R21406 DVSS.n5355 DVSS.n3372 4.5005
R21407 DVSS.n5357 DVSS.n3371 4.5005
R21408 DVSS.n5357 DVSS.n3372 4.5005
R21409 DVSS.n5361 DVSS.n3371 4.5005
R21410 DVSS.n5361 DVSS.n3372 4.5005
R21411 DVSS.n5363 DVSS.n3371 4.5005
R21412 DVSS.n5363 DVSS.n3372 4.5005
R21413 DVSS.n5360 DVSS.n3371 4.5005
R21414 DVSS.n5360 DVSS.n3372 4.5005
R21415 DVSS.n5366 DVSS.n3375 4.5005
R21416 DVSS.n3375 DVSS.n3371 4.5005
R21417 DVSS.n3375 DVSS.n3372 4.5005
R21418 DVSS.n3372 DVSS.n3365 4.5005
R21419 DVSS.n3373 DVSS.n3365 4.5005
R21420 DVSS.n3371 DVSS.n3365 4.5005
R21421 DVSS.n5366 DVSS.n3365 4.5005
R21422 DVSS.n3372 DVSS.n3367 4.5005
R21423 DVSS.n3373 DVSS.n3367 4.5005
R21424 DVSS.n3371 DVSS.n3367 4.5005
R21425 DVSS.n5366 DVSS.n3367 4.5005
R21426 DVSS.n3372 DVSS.n3370 4.5005
R21427 DVSS.n3373 DVSS.n3370 4.5005
R21428 DVSS.n3371 DVSS.n3370 4.5005
R21429 DVSS.n5366 DVSS.n3370 4.5005
R21430 DVSS.n5367 DVSS.n3372 4.5005
R21431 DVSS.n5367 DVSS.n3373 4.5005
R21432 DVSS.n5367 DVSS.n3371 4.5005
R21433 DVSS.n5367 DVSS.n5366 4.5005
R21434 DVSS.n5365 DVSS.n3372 4.5005
R21435 DVSS.n5365 DVSS.n3373 4.5005
R21436 DVSS.n5365 DVSS.n3371 4.5005
R21437 DVSS.n5366 DVSS.n5365 4.5005
R21438 DVSS.n7658 DVSS.n2174 4.5005
R21439 DVSS.n2174 DVSS.n2162 4.5005
R21440 DVSS.n7656 DVSS.n2174 4.5005
R21441 DVSS.n7632 DVSS.n2162 4.5005
R21442 DVSS.n7656 DVSS.n7632 4.5005
R21443 DVSS.n2188 DVSS.n2162 4.5005
R21444 DVSS.n7656 DVSS.n2188 4.5005
R21445 DVSS.n7633 DVSS.n2162 4.5005
R21446 DVSS.n7656 DVSS.n7633 4.5005
R21447 DVSS.n2187 DVSS.n2162 4.5005
R21448 DVSS.n7656 DVSS.n2187 4.5005
R21449 DVSS.n7634 DVSS.n2162 4.5005
R21450 DVSS.n7656 DVSS.n7634 4.5005
R21451 DVSS.n2186 DVSS.n2162 4.5005
R21452 DVSS.n7656 DVSS.n2186 4.5005
R21453 DVSS.n7635 DVSS.n2162 4.5005
R21454 DVSS.n7656 DVSS.n7635 4.5005
R21455 DVSS.n2185 DVSS.n2162 4.5005
R21456 DVSS.n7656 DVSS.n2185 4.5005
R21457 DVSS.n7636 DVSS.n2162 4.5005
R21458 DVSS.n7656 DVSS.n7636 4.5005
R21459 DVSS.n2184 DVSS.n2162 4.5005
R21460 DVSS.n7656 DVSS.n2184 4.5005
R21461 DVSS.n7637 DVSS.n2162 4.5005
R21462 DVSS.n7656 DVSS.n7637 4.5005
R21463 DVSS.n2183 DVSS.n2162 4.5005
R21464 DVSS.n7656 DVSS.n2183 4.5005
R21465 DVSS.n7638 DVSS.n2162 4.5005
R21466 DVSS.n7656 DVSS.n7638 4.5005
R21467 DVSS.n2182 DVSS.n2162 4.5005
R21468 DVSS.n7656 DVSS.n2182 4.5005
R21469 DVSS.n7639 DVSS.n2162 4.5005
R21470 DVSS.n7656 DVSS.n7639 4.5005
R21471 DVSS.n2181 DVSS.n2162 4.5005
R21472 DVSS.n7656 DVSS.n2181 4.5005
R21473 DVSS.n7640 DVSS.n2162 4.5005
R21474 DVSS.n7656 DVSS.n7640 4.5005
R21475 DVSS.n2180 DVSS.n2162 4.5005
R21476 DVSS.n7656 DVSS.n2180 4.5005
R21477 DVSS.n7641 DVSS.n2162 4.5005
R21478 DVSS.n7656 DVSS.n7641 4.5005
R21479 DVSS.n2179 DVSS.n2162 4.5005
R21480 DVSS.n7656 DVSS.n2179 4.5005
R21481 DVSS.n7655 DVSS.n2162 4.5005
R21482 DVSS.n7656 DVSS.n7655 4.5005
R21483 DVSS.n2178 DVSS.n2162 4.5005
R21484 DVSS.n7656 DVSS.n2178 4.5005
R21485 DVSS.n7658 DVSS.n7657 4.5005
R21486 DVSS.n7657 DVSS.n2162 4.5005
R21487 DVSS.n7657 DVSS.n7656 4.5005
R21488 DVSS.n8152 DVSS.n1789 4.5005
R21489 DVSS.n1789 DVSS.n1788 4.5005
R21490 DVSS.n8149 DVSS.n1789 4.5005
R21491 DVSS.n1800 DVSS.n1788 4.5005
R21492 DVSS.n8149 DVSS.n1800 4.5005
R21493 DVSS.n8139 DVSS.n1788 4.5005
R21494 DVSS.n8149 DVSS.n8139 4.5005
R21495 DVSS.n1799 DVSS.n1788 4.5005
R21496 DVSS.n8149 DVSS.n1799 4.5005
R21497 DVSS.n8140 DVSS.n1788 4.5005
R21498 DVSS.n8149 DVSS.n8140 4.5005
R21499 DVSS.n1798 DVSS.n1788 4.5005
R21500 DVSS.n8149 DVSS.n1798 4.5005
R21501 DVSS.n8147 DVSS.n1788 4.5005
R21502 DVSS.n8149 DVSS.n8147 4.5005
R21503 DVSS.n1797 DVSS.n1788 4.5005
R21504 DVSS.n8149 DVSS.n1797 4.5005
R21505 DVSS.n8148 DVSS.n1788 4.5005
R21506 DVSS.n8149 DVSS.n8148 4.5005
R21507 DVSS.n8150 DVSS.n1788 4.5005
R21508 DVSS.n8150 DVSS.n8149 4.5005
R21509 DVSS.n1794 DVSS.n1788 4.5005
R21510 DVSS.n8145 DVSS.n1794 4.5005
R21511 DVSS.n8149 DVSS.n1794 4.5005
R21512 DVSS.n1727 DVSS.n1557 4.5005
R21513 DVSS.n1594 DVSS.n1557 4.5005
R21514 DVSS.n1724 DVSS.n1557 4.5005
R21515 DVSS.n1605 DVSS.n1594 4.5005
R21516 DVSS.n1724 DVSS.n1605 4.5005
R21517 DVSS.n1714 DVSS.n1594 4.5005
R21518 DVSS.n1724 DVSS.n1714 4.5005
R21519 DVSS.n1604 DVSS.n1594 4.5005
R21520 DVSS.n1724 DVSS.n1604 4.5005
R21521 DVSS.n1715 DVSS.n1594 4.5005
R21522 DVSS.n1724 DVSS.n1715 4.5005
R21523 DVSS.n1603 DVSS.n1594 4.5005
R21524 DVSS.n1724 DVSS.n1603 4.5005
R21525 DVSS.n1722 DVSS.n1594 4.5005
R21526 DVSS.n1724 DVSS.n1722 4.5005
R21527 DVSS.n1602 DVSS.n1594 4.5005
R21528 DVSS.n1724 DVSS.n1602 4.5005
R21529 DVSS.n1723 DVSS.n1594 4.5005
R21530 DVSS.n1724 DVSS.n1723 4.5005
R21531 DVSS.n1725 DVSS.n1594 4.5005
R21532 DVSS.n1725 DVSS.n1724 4.5005
R21533 DVSS.n1599 DVSS.n1594 4.5005
R21534 DVSS.n1720 DVSS.n1599 4.5005
R21535 DVSS.n1724 DVSS.n1599 4.5005
R21536 DVSS.n5960 DVSS.n2857 4.5005
R21537 DVSS.n5958 DVSS.n2857 4.5005
R21538 DVSS.n2865 DVSS.n2857 4.5005
R21539 DVSS.n5960 DVSS.n2848 4.5005
R21540 DVSS.n5958 DVSS.n2848 4.5005
R21541 DVSS.n2865 DVSS.n2848 4.5005
R21542 DVSS.n5959 DVSS.n2863 4.5005
R21543 DVSS.n5959 DVSS.n2865 4.5005
R21544 DVSS.n5960 DVSS.n5959 4.5005
R21545 DVSS.n5959 DVSS.n5958 4.5005
R21546 DVSS.n9002 DVSS.n716 4.5005
R21547 DVSS.n9004 DVSS.n716 4.5005
R21548 DVSS.n9004 DVSS.n718 4.5005
R21549 DVSS.n9004 DVSS.n715 4.5005
R21550 DVSS.n9003 DVSS.n9002 4.5005
R21551 DVSS.n9004 DVSS.n9003 4.5005
R21552 DVSS.n9010 DVSS.n709 4.5005
R21553 DVSS.n9016 DVSS.n702 4.5005
R21554 DVSS.n9023 DVSS.n9017 4.5005
R21555 DVSS.n9017 DVSS.n382 4.5005
R21556 DVSS.n9383 DVSS.n383 4.5005
R21557 DVSS.n9381 DVSS.n383 4.5005
R21558 DVSS.n9376 DVSS.n9373 4.5005
R21559 DVSS.n9541 DVSS.n330 4.5005
R21560 DVSS.n9008 DVSS.n711 4.5005
R21561 DVSS.n9010 DVSS.n711 4.5005
R21562 DVSS.n9014 DVSS.n704 4.5005
R21563 DVSS.n9016 DVSS.n704 4.5005
R21564 DVSS.n9021 DVSS.n382 4.5005
R21565 DVSS.n9381 DVSS.n9380 4.5005
R21566 DVSS.n9375 DVSS.n9370 4.5005
R21567 DVSS.n9376 DVSS.n9375 4.5005
R21568 DVSS.n9540 DVSS.n326 4.5005
R21569 DVSS.n9541 DVSS.n9540 4.5005
R21570 DVSS.n9008 DVSS.n708 4.5005
R21571 DVSS.n9010 DVSS.n708 4.5005
R21572 DVSS.n9014 DVSS.n701 4.5005
R21573 DVSS.n9016 DVSS.n701 4.5005
R21574 DVSS.n9019 DVSS.n382 4.5005
R21575 DVSS.n9381 DVSS.n388 4.5005
R21576 DVSS.n9372 DVSS.n9370 4.5005
R21577 DVSS.n9376 DVSS.n9372 4.5005
R21578 DVSS.n328 DVSS.n326 4.5005
R21579 DVSS.n9541 DVSS.n328 4.5005
R21580 DVSS.n9009 DVSS.n9006 4.5005
R21581 DVSS.n9009 DVSS.n9008 4.5005
R21582 DVSS.n9010 DVSS.n9009 4.5005
R21583 DVSS.n9015 DVSS.n9012 4.5005
R21584 DVSS.n9015 DVSS.n9014 4.5005
R21585 DVSS.n9016 DVSS.n9015 4.5005
R21586 DVSS.n9024 DVSS.n9023 4.5005
R21587 DVSS.n9024 DVSS.n382 4.5005
R21588 DVSS.n9383 DVSS.n9382 4.5005
R21589 DVSS.n9382 DVSS.n9381 4.5005
R21590 DVSS.n9378 DVSS.n9377 4.5005
R21591 DVSS.n9377 DVSS.n9370 4.5005
R21592 DVSS.n9377 DVSS.n9376 4.5005
R21593 DVSS.n9542 DVSS.n325 4.5005
R21594 DVSS.n9542 DVSS.n326 4.5005
R21595 DVSS.n9542 DVSS.n9541 4.5005
R21596 DVSS.n9537 DVSS.n331 4.5005
R21597 DVSS.n9534 DVSS.n331 4.5005
R21598 DVSS.n9535 DVSS.n9534 4.5005
R21599 DVSS.n9534 DVSS.n334 4.5005
R21600 DVSS.n9537 DVSS.n51 4.5005
R21601 DVSS.n9534 DVSS.n51 4.5005
R21602 DVSS.n786 DVSS.n781 4.5005
R21603 DVSS.n8883 DVSS.n786 4.5005
R21604 DVSS.n8883 DVSS.n8882 4.5005
R21605 DVSS.n8884 DVSS.n781 4.5005
R21606 DVSS.n8885 DVSS.n8884 4.5005
R21607 DVSS.n8884 DVSS.n8883 4.5005
R21608 DVSS.n8875 DVSS.n796 4.5005
R21609 DVSS.n8870 DVSS.n8861 4.5005
R21610 DVSS.n8869 DVSS.n8862 4.5005
R21611 DVSS.n8862 DVSS.n378 4.5005
R21612 DVSS.n9392 DVSS.n372 4.5005
R21613 DVSS.n9395 DVSS.n372 4.5005
R21614 DVSS.n9404 DVSS.n369 4.5005
R21615 DVSS.n9413 DVSS.n367 4.5005
R21616 DVSS.n8877 DVSS.n8876 4.5005
R21617 DVSS.n8876 DVSS.n8875 4.5005
R21618 DVSS.n8872 DVSS.n8871 4.5005
R21619 DVSS.n8871 DVSS.n8870 4.5005
R21620 DVSS.n8867 DVSS.n378 4.5005
R21621 DVSS.n9395 DVSS.n373 4.5005
R21622 DVSS.n9399 DVSS.n370 4.5005
R21623 DVSS.n9404 DVSS.n370 4.5005
R21624 DVSS.n9408 DVSS.n368 4.5005
R21625 DVSS.n9413 DVSS.n368 4.5005
R21626 DVSS.n8875 DVSS.n795 4.5005
R21627 DVSS.n8870 DVSS.n805 4.5005
R21628 DVSS.n9404 DVSS.n224 4.5005
R21629 DVSS.n9413 DVSS.n185 4.5005
R21630 DVSS.n8879 DVSS.n8878 4.5005
R21631 DVSS.n8878 DVSS.n8877 4.5005
R21632 DVSS.n8874 DVSS.n8873 4.5005
R21633 DVSS.n8873 DVSS.n8872 4.5005
R21634 DVSS.n603 DVSS.n378 4.5005
R21635 DVSS.n9395 DVSS.n9394 4.5005
R21636 DVSS.n9397 DVSS.n220 4.5005
R21637 DVSS.n9399 DVSS.n220 4.5005
R21638 DVSS.n9406 DVSS.n181 4.5005
R21639 DVSS.n9408 DVSS.n181 4.5005
R21640 DVSS.n9415 DVSS.n366 4.5005
R21641 DVSS.n9419 DVSS.n366 4.5005
R21642 DVSS.n9419 DVSS.n9418 4.5005
R21643 DVSS.n365 DVSS.n158 4.5005
R21644 DVSS.n9419 DVSS.n158 4.5005
R21645 DVSS.n9419 DVSS.n156 4.5005
R21646 DVSS.n7156 DVSS.n7155 4.5005
R21647 DVSS.n7239 DVSS.n7156 4.5005
R21648 DVSS.n7186 DVSS.n7185 4.5005
R21649 DVSS.n7181 DVSS.n7180 4.5005
R21650 DVSS.n7191 DVSS.n7190 4.5005
R21651 DVSS.n7192 DVSS.n7179 4.5005
R21652 DVSS.n7194 DVSS.n7193 4.5005
R21653 DVSS.n7177 DVSS.n7176 4.5005
R21654 DVSS.n7199 DVSS.n7198 4.5005
R21655 DVSS.n7200 DVSS.n7175 4.5005
R21656 DVSS.n7202 DVSS.n7201 4.5005
R21657 DVSS.n7173 DVSS.n7172 4.5005
R21658 DVSS.n7207 DVSS.n7206 4.5005
R21659 DVSS.n7208 DVSS.n7171 4.5005
R21660 DVSS.n7210 DVSS.n7209 4.5005
R21661 DVSS.n7213 DVSS.n7168 4.5005
R21662 DVSS.n7215 DVSS.n7214 4.5005
R21663 DVSS.n7217 DVSS.n7216 4.5005
R21664 DVSS.n7166 DVSS.n7165 4.5005
R21665 DVSS.n7222 DVSS.n7221 4.5005
R21666 DVSS.n7223 DVSS.n7164 4.5005
R21667 DVSS.n7225 DVSS.n7224 4.5005
R21668 DVSS.n7162 DVSS.n7161 4.5005
R21669 DVSS.n7230 DVSS.n7229 4.5005
R21670 DVSS.n7231 DVSS.n7160 4.5005
R21671 DVSS.n7233 DVSS.n7232 4.5005
R21672 DVSS.n7158 DVSS.n7157 4.5005
R21673 DVSS.n7238 DVSS.n7237 4.5005
R21674 DVSS.n7237 DVSS.n7236 4.5005
R21675 DVSS.n7235 DVSS.n7158 4.5005
R21676 DVSS.n7234 DVSS.n7233 4.5005
R21677 DVSS.n7160 DVSS.n7159 4.5005
R21678 DVSS.n7229 DVSS.n7228 4.5005
R21679 DVSS.n7227 DVSS.n7162 4.5005
R21680 DVSS.n7226 DVSS.n7225 4.5005
R21681 DVSS.n7164 DVSS.n7163 4.5005
R21682 DVSS.n7221 DVSS.n7220 4.5005
R21683 DVSS.n7219 DVSS.n7166 4.5005
R21684 DVSS.n7218 DVSS.n7217 4.5005
R21685 DVSS.n7214 DVSS.n7167 4.5005
R21686 DVSS.n7213 DVSS.n7212 4.5005
R21687 DVSS.n7211 DVSS.n7210 4.5005
R21688 DVSS.n7171 DVSS.n7170 4.5005
R21689 DVSS.n7206 DVSS.n7205 4.5005
R21690 DVSS.n7204 DVSS.n7173 4.5005
R21691 DVSS.n7203 DVSS.n7202 4.5005
R21692 DVSS.n7175 DVSS.n7174 4.5005
R21693 DVSS.n7198 DVSS.n7197 4.5005
R21694 DVSS.n7196 DVSS.n7177 4.5005
R21695 DVSS.n7195 DVSS.n7194 4.5005
R21696 DVSS.n7179 DVSS.n7178 4.5005
R21697 DVSS.n7190 DVSS.n7189 4.5005
R21698 DVSS.n7188 DVSS.n7181 4.5005
R21699 DVSS.n7187 DVSS.n7186 4.5005
R21700 DVSS.n7183 DVSS.n7182 4.5005
R21701 DVSS.n7184 DVSS.n7183 4.5005
R21702 DVSS.n8210 DVSS.n8209 4.5005
R21703 DVSS.n8209 DVSS.n1533 4.5005
R21704 DVSS.n8209 DVSS.n8208 4.5005
R21705 DVSS.n7246 DVSS.n7240 4.5005
R21706 DVSS.n1538 DVSS.n1533 4.5005
R21707 DVSS.n8208 DVSS.n1538 4.5005
R21708 DVSS.n8211 DVSS.n1533 4.5005
R21709 DVSS.n8211 DVSS.n8210 4.5005
R21710 DVSS.n8206 DVSS.n1541 4.5005
R21711 DVSS.n8204 DVSS.n1541 4.5005
R21712 DVSS.n8200 DVSS.n1541 4.5005
R21713 DVSS.n8199 DVSS.n1555 4.5005
R21714 DVSS.n8197 DVSS.n1555 4.5005
R21715 DVSS.n8193 DVSS.n1555 4.5005
R21716 DVSS.n8204 DVSS.n8201 4.5005
R21717 DVSS.n8201 DVSS.n8200 4.5005
R21718 DVSS.n8197 DVSS.n8194 4.5005
R21719 DVSS.n8194 DVSS.n8193 4.5005
R21720 DVSS.n8198 DVSS.n8197 4.5005
R21721 DVSS.n8199 DVSS.n8198 4.5005
R21722 DVSS.n8205 DVSS.n8204 4.5005
R21723 DVSS.n8206 DVSS.n8205 4.5005
R21724 DVSS.n8187 DVSS.n1750 4.5005
R21725 DVSS.n8186 DVSS.n1751 4.5005
R21726 DVSS.n8186 DVSS.n1750 4.5005
R21727 DVSS.n2890 DVSS.n2881 4.5005
R21728 DVSS.n5930 DVSS.n2881 4.5005
R21729 DVSS.n5941 DVSS.n2881 4.5005
R21730 DVSS.n5943 DVSS.n2881 4.5005
R21731 DVSS.n2890 DVSS.n2883 4.5005
R21732 DVSS.n5930 DVSS.n2883 4.5005
R21733 DVSS.n5943 DVSS.n2883 4.5005
R21734 DVSS.n5930 DVSS.n2880 4.5005
R21735 DVSS.n5943 DVSS.n2880 4.5005
R21736 DVSS.n5930 DVSS.n2884 4.5005
R21737 DVSS.n5943 DVSS.n2884 4.5005
R21738 DVSS.n5930 DVSS.n2879 4.5005
R21739 DVSS.n5943 DVSS.n2879 4.5005
R21740 DVSS.n5930 DVSS.n2885 4.5005
R21741 DVSS.n5943 DVSS.n2885 4.5005
R21742 DVSS.n2890 DVSS.n2878 4.5005
R21743 DVSS.n5930 DVSS.n2878 4.5005
R21744 DVSS.n5943 DVSS.n2878 4.5005
R21745 DVSS.n4926 DVSS.n4913 4.5005
R21746 DVSS.n4942 DVSS.n4913 4.5005
R21747 DVSS.n4944 DVSS.n4913 4.5005
R21748 DVSS.n4942 DVSS.n4911 4.5005
R21749 DVSS.n4944 DVSS.n4911 4.5005
R21750 DVSS.n4942 DVSS.n4914 4.5005
R21751 DVSS.n4944 DVSS.n4914 4.5005
R21752 DVSS.n4942 DVSS.n4910 4.5005
R21753 DVSS.n4944 DVSS.n4910 4.5005
R21754 DVSS.n4942 DVSS.n4915 4.5005
R21755 DVSS.n4944 DVSS.n4915 4.5005
R21756 DVSS.n4942 DVSS.n4909 4.5005
R21757 DVSS.n4944 DVSS.n4909 4.5005
R21758 DVSS.n4942 DVSS.n4916 4.5005
R21759 DVSS.n4922 DVSS.n4916 4.5005
R21760 DVSS.n4944 DVSS.n4916 4.5005
R21761 DVSS.n4944 DVSS.n4908 4.5005
R21762 DVSS.n4922 DVSS.n4908 4.5005
R21763 DVSS.n4942 DVSS.n4908 4.5005
R21764 DVSS.n4926 DVSS.n4908 4.5005
R21765 DVSS.n4926 DVSS.n4917 4.5005
R21766 DVSS.n4942 DVSS.n4917 4.5005
R21767 DVSS.n4922 DVSS.n4917 4.5005
R21768 DVSS.n4944 DVSS.n4917 4.5005
R21769 DVSS.n4926 DVSS.n4907 4.5005
R21770 DVSS.n4942 DVSS.n4907 4.5005
R21771 DVSS.n4922 DVSS.n4907 4.5005
R21772 DVSS.n4944 DVSS.n4907 4.5005
R21773 DVSS.n4943 DVSS.n4926 4.5005
R21774 DVSS.n4943 DVSS.n4942 4.5005
R21775 DVSS.n4943 DVSS.n4922 4.5005
R21776 DVSS.n4944 DVSS.n4943 4.5005
R21777 DVSS.n5915 DVSS.n2932 4.5005
R21778 DVSS.n2932 DVSS.n2922 4.5005
R21779 DVSS.n2932 DVSS.n2924 4.5005
R21780 DVSS.n2932 DVSS.n2923 4.5005
R21781 DVSS.n5915 DVSS.n2930 4.5005
R21782 DVSS.n2930 DVSS.n2922 4.5005
R21783 DVSS.n2930 DVSS.n2924 4.5005
R21784 DVSS.n2930 DVSS.n2923 4.5005
R21785 DVSS.n5916 DVSS.n2923 4.5005
R21786 DVSS.n5916 DVSS.n2924 4.5005
R21787 DVSS.n5916 DVSS.n2922 4.5005
R21788 DVSS.n5916 DVSS.n5915 4.5005
R21789 DVSS.n2923 DVSS.n2917 4.5005
R21790 DVSS.n2924 DVSS.n2917 4.5005
R21791 DVSS.n2922 DVSS.n2917 4.5005
R21792 DVSS.n5915 DVSS.n2917 4.5005
R21793 DVSS.n2923 DVSS.n2919 4.5005
R21794 DVSS.n2924 DVSS.n2919 4.5005
R21795 DVSS.n5915 DVSS.n2919 4.5005
R21796 DVSS.n2929 DVSS.n2924 4.5005
R21797 DVSS.n5915 DVSS.n2929 4.5005
R21798 DVSS.n2935 DVSS.n2924 4.5005
R21799 DVSS.n5915 DVSS.n2935 4.5005
R21800 DVSS.n2927 DVSS.n2924 4.5005
R21801 DVSS.n5915 DVSS.n2927 4.5005
R21802 DVSS.n2938 DVSS.n2924 4.5005
R21803 DVSS.n5915 DVSS.n2938 4.5005
R21804 DVSS.n2926 DVSS.n2924 4.5005
R21805 DVSS.n5915 DVSS.n2926 4.5005
R21806 DVSS.n5914 DVSS.n2924 4.5005
R21807 DVSS.n5914 DVSS.n2922 4.5005
R21808 DVSS.n5915 DVSS.n5914 4.5005
R21809 DVSS.n5913 DVSS.n2941 4.5005
R21810 DVSS.n5913 DVSS.n2942 4.5005
R21811 DVSS.n5913 DVSS.n5912 4.5005
R21812 DVSS.n2948 DVSS.n2942 4.5005
R21813 DVSS.n5912 DVSS.n2948 4.5005
R21814 DVSS.n2951 DVSS.n2942 4.5005
R21815 DVSS.n5912 DVSS.n2951 4.5005
R21816 DVSS.n2947 DVSS.n2942 4.5005
R21817 DVSS.n5912 DVSS.n2947 4.5005
R21818 DVSS.n2953 DVSS.n2942 4.5005
R21819 DVSS.n5912 DVSS.n2953 4.5005
R21820 DVSS.n2946 DVSS.n2941 4.5005
R21821 DVSS.n2946 DVSS.n2942 4.5005
R21822 DVSS.n5912 DVSS.n2946 4.5005
R21823 DVSS.n5912 DVSS.n2954 4.5005
R21824 DVSS.n2959 DVSS.n2954 4.5005
R21825 DVSS.n2954 DVSS.n2942 4.5005
R21826 DVSS.n2954 DVSS.n2941 4.5005
R21827 DVSS.n5912 DVSS.n2945 4.5005
R21828 DVSS.n2959 DVSS.n2945 4.5005
R21829 DVSS.n2945 DVSS.n2942 4.5005
R21830 DVSS.n2945 DVSS.n2941 4.5005
R21831 DVSS.n5912 DVSS.n2955 4.5005
R21832 DVSS.n2959 DVSS.n2955 4.5005
R21833 DVSS.n2955 DVSS.n2942 4.5005
R21834 DVSS.n2955 DVSS.n2941 4.5005
R21835 DVSS.n2944 DVSS.n2941 4.5005
R21836 DVSS.n2944 DVSS.n2942 4.5005
R21837 DVSS.n2959 DVSS.n2944 4.5005
R21838 DVSS.n5912 DVSS.n2944 4.5005
R21839 DVSS.n5911 DVSS.n2941 4.5005
R21840 DVSS.n5911 DVSS.n2942 4.5005
R21841 DVSS.n5911 DVSS.n2959 4.5005
R21842 DVSS.n5912 DVSS.n5911 4.5005
R21843 DVSS.n2133 DVSS.n2119 4.5005
R21844 DVSS.n2133 DVSS.n2120 4.5005
R21845 DVSS.n7693 DVSS.n2133 4.5005
R21846 DVSS.n2136 DVSS.n2120 4.5005
R21847 DVSS.n7693 DVSS.n2136 4.5005
R21848 DVSS.n2132 DVSS.n2120 4.5005
R21849 DVSS.n7693 DVSS.n2132 4.5005
R21850 DVSS.n2138 DVSS.n2120 4.5005
R21851 DVSS.n7693 DVSS.n2138 4.5005
R21852 DVSS.n2131 DVSS.n2120 4.5005
R21853 DVSS.n7693 DVSS.n2131 4.5005
R21854 DVSS.n2140 DVSS.n2120 4.5005
R21855 DVSS.n7693 DVSS.n2140 4.5005
R21856 DVSS.n2130 DVSS.n2120 4.5005
R21857 DVSS.n7693 DVSS.n2130 4.5005
R21858 DVSS.n2142 DVSS.n2120 4.5005
R21859 DVSS.n7693 DVSS.n2142 4.5005
R21860 DVSS.n2129 DVSS.n2120 4.5005
R21861 DVSS.n7693 DVSS.n2129 4.5005
R21862 DVSS.n2144 DVSS.n2120 4.5005
R21863 DVSS.n7693 DVSS.n2144 4.5005
R21864 DVSS.n2128 DVSS.n2120 4.5005
R21865 DVSS.n7693 DVSS.n2128 4.5005
R21866 DVSS.n2146 DVSS.n2120 4.5005
R21867 DVSS.n7693 DVSS.n2146 4.5005
R21868 DVSS.n2127 DVSS.n2120 4.5005
R21869 DVSS.n7693 DVSS.n2127 4.5005
R21870 DVSS.n2148 DVSS.n2120 4.5005
R21871 DVSS.n7693 DVSS.n2148 4.5005
R21872 DVSS.n2126 DVSS.n2120 4.5005
R21873 DVSS.n7693 DVSS.n2126 4.5005
R21874 DVSS.n2150 DVSS.n2120 4.5005
R21875 DVSS.n7693 DVSS.n2150 4.5005
R21876 DVSS.n2125 DVSS.n2120 4.5005
R21877 DVSS.n7693 DVSS.n2125 4.5005
R21878 DVSS.n2152 DVSS.n2120 4.5005
R21879 DVSS.n7693 DVSS.n2152 4.5005
R21880 DVSS.n2124 DVSS.n2120 4.5005
R21881 DVSS.n7693 DVSS.n2124 4.5005
R21882 DVSS.n2154 DVSS.n2120 4.5005
R21883 DVSS.n7693 DVSS.n2154 4.5005
R21884 DVSS.n2123 DVSS.n2120 4.5005
R21885 DVSS.n7693 DVSS.n2123 4.5005
R21886 DVSS.n7692 DVSS.n2120 4.5005
R21887 DVSS.n7693 DVSS.n7692 4.5005
R21888 DVSS.n2122 DVSS.n2120 4.5005
R21889 DVSS.n7693 DVSS.n2122 4.5005
R21890 DVSS.n7694 DVSS.n2119 4.5005
R21891 DVSS.n7694 DVSS.n2120 4.5005
R21892 DVSS.n7694 DVSS.n7693 4.5005
R21893 DVSS.n8174 DVSS.n1772 4.5005
R21894 DVSS.n1772 DVSS.n1763 4.5005
R21895 DVSS.n8178 DVSS.n1772 4.5005
R21896 DVSS.n1769 DVSS.n1763 4.5005
R21897 DVSS.n8178 DVSS.n1769 4.5005
R21898 DVSS.n1774 DVSS.n1763 4.5005
R21899 DVSS.n8178 DVSS.n1774 4.5005
R21900 DVSS.n1768 DVSS.n1763 4.5005
R21901 DVSS.n8178 DVSS.n1768 4.5005
R21902 DVSS.n1776 DVSS.n1763 4.5005
R21903 DVSS.n8178 DVSS.n1776 4.5005
R21904 DVSS.n1767 DVSS.n1763 4.5005
R21905 DVSS.n8178 DVSS.n1767 4.5005
R21906 DVSS.n1778 DVSS.n1763 4.5005
R21907 DVSS.n8178 DVSS.n1778 4.5005
R21908 DVSS.n1766 DVSS.n1763 4.5005
R21909 DVSS.n8178 DVSS.n1766 4.5005
R21910 DVSS.n8177 DVSS.n1763 4.5005
R21911 DVSS.n8178 DVSS.n8177 4.5005
R21912 DVSS.n1765 DVSS.n1763 4.5005
R21913 DVSS.n8178 DVSS.n1765 4.5005
R21914 DVSS.n8179 DVSS.n1763 4.5005
R21915 DVSS.n8179 DVSS.n1762 4.5005
R21916 DVSS.n8179 DVSS.n8178 4.5005
R21917 DVSS.n1749 DVSS.n1563 4.5005
R21918 DVSS.n1749 DVSS.n1564 4.5005
R21919 DVSS.n1749 DVSS.n1748 4.5005
R21920 DVSS.n1570 DVSS.n1564 4.5005
R21921 DVSS.n1748 DVSS.n1570 4.5005
R21922 DVSS.n1573 DVSS.n1564 4.5005
R21923 DVSS.n1748 DVSS.n1573 4.5005
R21924 DVSS.n1569 DVSS.n1564 4.5005
R21925 DVSS.n1748 DVSS.n1569 4.5005
R21926 DVSS.n1575 DVSS.n1564 4.5005
R21927 DVSS.n1748 DVSS.n1575 4.5005
R21928 DVSS.n1568 DVSS.n1564 4.5005
R21929 DVSS.n1748 DVSS.n1568 4.5005
R21930 DVSS.n1577 DVSS.n1564 4.5005
R21931 DVSS.n1748 DVSS.n1577 4.5005
R21932 DVSS.n1567 DVSS.n1564 4.5005
R21933 DVSS.n1748 DVSS.n1567 4.5005
R21934 DVSS.n1579 DVSS.n1564 4.5005
R21935 DVSS.n1748 DVSS.n1579 4.5005
R21936 DVSS.n1566 DVSS.n1564 4.5005
R21937 DVSS.n1748 DVSS.n1566 4.5005
R21938 DVSS.n1747 DVSS.n1564 4.5005
R21939 DVSS.n1747 DVSS.n1746 4.5005
R21940 DVSS.n1748 DVSS.n1747 4.5005
R21941 DVSS.n5943 DVSS.n2886 4.5005
R21942 DVSS.n5941 DVSS.n2886 4.5005
R21943 DVSS.n2890 DVSS.n2886 4.5005
R21944 DVSS.n5943 DVSS.n2877 4.5005
R21945 DVSS.n5941 DVSS.n2877 4.5005
R21946 DVSS.n2890 DVSS.n2877 4.5005
R21947 DVSS.n5942 DVSS.n2890 4.5005
R21948 DVSS.n5942 DVSS.n5930 4.5005
R21949 DVSS.n5943 DVSS.n5942 4.5005
R21950 DVSS.n5942 DVSS.n5941 4.5005
R21951 DVSS.n5923 DVSS.n2887 4.5005
R21952 DVSS.n4471 DVSS.n4470 4.5005
R21953 DVSS.n4595 DVSS.n3792 4.5005
R21954 DVSS.n4599 DVSS.n4598 4.5005
R21955 DVSS.n4602 DVSS.n4600 4.5005
R21956 DVSS.n4602 DVSS.n2759 4.5005
R21957 DVSS.n6011 DVSS.n2761 4.5005
R21958 DVSS.n6009 DVSS.n2761 4.5005
R21959 DVSS.n6006 DVSS.n6005 4.5005
R21960 DVSS.n2906 DVSS.n2905 4.5005
R21961 DVSS.n2910 DVSS.n2909 4.5005
R21962 DVSS.n5927 DVSS.n5924 4.5005
R21963 DVSS.n5925 DVSS.n5924 4.5005
R21964 DVSS.n4473 DVSS.n3826 4.5005
R21965 DVSS.n4590 DVSS.n3798 4.5005
R21966 DVSS.n4596 DVSS.n3744 4.5005
R21967 DVSS.n6008 DVSS.n2768 4.5005
R21968 DVSS.n2831 DVSS.n2777 4.5005
R21969 DVSS.n2907 DVSS.n2864 4.5005
R21970 DVSS.n5928 DVSS.n5927 4.5005
R21971 DVSS.n5924 DVSS.n5923 4.5005
R21972 DVSS.n4473 DVSS.n3824 4.5005
R21973 DVSS.n4464 DVSS.n3824 4.5005
R21974 DVSS.n4466 DVSS.n3824 4.5005
R21975 DVSS.n4468 DVSS.n3824 4.5005
R21976 DVSS.n4470 DVSS.n3824 4.5005
R21977 DVSS.n4594 DVSS.n3798 4.5005
R21978 DVSS.n4594 DVSS.n3795 4.5005
R21979 DVSS.n4594 DVSS.n4593 4.5005
R21980 DVSS.n4594 DVSS.n3794 4.5005
R21981 DVSS.n4595 DVSS.n4594 4.5005
R21982 DVSS.n4596 DVSS.n3743 4.5005
R21983 DVSS.n3790 DVSS.n3743 4.5005
R21984 DVSS.n3788 DVSS.n3743 4.5005
R21985 DVSS.n3786 DVSS.n3743 4.5005
R21986 DVSS.n4599 DVSS.n3743 4.5005
R21987 DVSS.n4600 DVSS.n3780 4.5005
R21988 DVSS.n4604 DVSS.n3780 4.5005
R21989 DVSS.n4601 DVSS.n3780 4.5005
R21990 DVSS.n3780 DVSS.n2759 4.5005
R21991 DVSS.n6011 DVSS.n6010 4.5005
R21992 DVSS.n6010 DVSS.n2766 4.5005
R21993 DVSS.n6010 DVSS.n2763 4.5005
R21994 DVSS.n6010 DVSS.n6009 4.5005
R21995 DVSS.n6008 DVSS.n6007 4.5005
R21996 DVSS.n6007 DVSS.n2772 4.5005
R21997 DVSS.n6007 DVSS.n2775 4.5005
R21998 DVSS.n6007 DVSS.n2771 4.5005
R21999 DVSS.n6007 DVSS.n6006 4.5005
R22000 DVSS.n2827 DVSS.n2777 4.5005
R22001 DVSS.n2903 DVSS.n2827 4.5005
R22002 DVSS.n2901 DVSS.n2827 4.5005
R22003 DVSS.n2899 DVSS.n2827 4.5005
R22004 DVSS.n2906 DVSS.n2827 4.5005
R22005 DVSS.n2907 DVSS.n2858 4.5005
R22006 DVSS.n2897 DVSS.n2858 4.5005
R22007 DVSS.n2895 DVSS.n2858 4.5005
R22008 DVSS.n2893 DVSS.n2858 4.5005
R22009 DVSS.n2910 DVSS.n2858 4.5005
R22010 DVSS.n4440 DVSS.n3860 4.5005
R22011 DVSS.n4438 DVSS.n3860 4.5005
R22012 DVSS.n4437 DVSS.n4191 4.5005
R22013 DVSS.n4435 DVSS.n4191 4.5005
R22014 DVSS.n3716 DVSS.n3712 4.5005
R22015 DVSS.n4803 DVSS.n3712 4.5005
R22016 DVSS.n4807 DVSS.n4806 4.5005
R22017 DVSS.n4823 DVSS.n3670 4.5005
R22018 DVSS.n4842 DVSS.n4824 4.5005
R22019 DVSS.n4845 DVSS.n4842 4.5005
R22020 DVSS.n4839 DVSS.n3626 4.5005
R22021 DVSS.n4837 DVSS.n3626 4.5005
R22022 DVSS.n4979 DVSS.n3590 4.5005
R22023 DVSS.n4979 DVSS.n4978 4.5005
R22024 DVSS.n4934 DVSS.n4933 4.5005
R22025 DVSS.n4934 DVSS.n4928 4.5005
R22026 DVSS.n4804 DVSS.n3702 4.5005
R22027 DVSS.n4821 DVSS.n4819 4.5005
R22028 DVSS.n4933 DVSS.n4918 4.5005
R22029 DVSS.n4440 DVSS.n3861 4.5005
R22030 DVSS.n3866 DVSS.n3861 4.5005
R22031 DVSS.n3863 DVSS.n3861 4.5005
R22032 DVSS.n4438 DVSS.n3861 4.5005
R22033 DVSS.n4437 DVSS.n4192 4.5005
R22034 DVSS.n4197 DVSS.n4192 4.5005
R22035 DVSS.n4194 DVSS.n4192 4.5005
R22036 DVSS.n4435 DVSS.n4192 4.5005
R22037 DVSS.n3716 DVSS.n3713 4.5005
R22038 DVSS.n4801 DVSS.n3713 4.5005
R22039 DVSS.n3715 DVSS.n3713 4.5005
R22040 DVSS.n4803 DVSS.n3713 4.5005
R22041 DVSS.n4804 DVSS.n3708 4.5005
R22042 DVSS.n3709 DVSS.n3708 4.5005
R22043 DVSS.n4806 DVSS.n3708 4.5005
R22044 DVSS.n4821 DVSS.n3671 4.5005
R22045 DVSS.n3673 DVSS.n3671 4.5005
R22046 DVSS.n4823 DVSS.n3671 4.5005
R22047 DVSS.n4843 DVSS.n4824 4.5005
R22048 DVSS.n4843 DVSS.n4825 4.5005
R22049 DVSS.n4843 DVSS.n3667 4.5005
R22050 DVSS.n4845 DVSS.n4843 4.5005
R22051 DVSS.n4839 DVSS.n4832 4.5005
R22052 DVSS.n4835 DVSS.n4832 4.5005
R22053 DVSS.n4833 DVSS.n4832 4.5005
R22054 DVSS.n4837 DVSS.n4832 4.5005
R22055 DVSS.n3594 DVSS.n3590 4.5005
R22056 DVSS.n4976 DVSS.n3594 4.5005
R22057 DVSS.n3596 DVSS.n3594 4.5005
R22058 DVSS.n4978 DVSS.n3594 4.5005
R22059 DVSS.n4933 DVSS.n4931 4.5005
R22060 DVSS.n4931 DVSS.n4928 4.5005
R22061 DVSS.n4933 DVSS.n4932 4.5005
R22062 DVSS.n4932 DVSS.n4928 4.5005
R22063 DVSS.n4440 DVSS.n3858 4.5005
R22064 DVSS.n3866 DVSS.n3858 4.5005
R22065 DVSS.n3863 DVSS.n3858 4.5005
R22066 DVSS.n4438 DVSS.n3858 4.5005
R22067 DVSS.n4437 DVSS.n3868 4.5005
R22068 DVSS.n4197 DVSS.n3868 4.5005
R22069 DVSS.n4194 DVSS.n3868 4.5005
R22070 DVSS.n4435 DVSS.n3868 4.5005
R22071 DVSS.n3716 DVSS.n3710 4.5005
R22072 DVSS.n4801 DVSS.n3710 4.5005
R22073 DVSS.n3715 DVSS.n3710 4.5005
R22074 DVSS.n4803 DVSS.n3710 4.5005
R22075 DVSS.n4804 DVSS.n3706 4.5005
R22076 DVSS.n3709 DVSS.n3706 4.5005
R22077 DVSS.n4806 DVSS.n3706 4.5005
R22078 DVSS.n4821 DVSS.n3668 4.5005
R22079 DVSS.n3673 DVSS.n3668 4.5005
R22080 DVSS.n4823 DVSS.n3668 4.5005
R22081 DVSS.n4846 DVSS.n4824 4.5005
R22082 DVSS.n4846 DVSS.n4825 4.5005
R22083 DVSS.n4846 DVSS.n3667 4.5005
R22084 DVSS.n4846 DVSS.n4845 4.5005
R22085 DVSS.n4839 DVSS.n4830 4.5005
R22086 DVSS.n4835 DVSS.n4830 4.5005
R22087 DVSS.n4833 DVSS.n4830 4.5005
R22088 DVSS.n4837 DVSS.n4830 4.5005
R22089 DVSS.n3591 DVSS.n3590 4.5005
R22090 DVSS.n4976 DVSS.n3591 4.5005
R22091 DVSS.n3596 DVSS.n3591 4.5005
R22092 DVSS.n4978 DVSS.n3591 4.5005
R22093 DVSS.n4932 DVSS.n2911 4.5005
R22094 DVSS.n4440 DVSS.n4439 4.5005
R22095 DVSS.n4439 DVSS.n3866 4.5005
R22096 DVSS.n4439 DVSS.n3863 4.5005
R22097 DVSS.n4439 DVSS.n4438 4.5005
R22098 DVSS.n4437 DVSS.n4436 4.5005
R22099 DVSS.n4436 DVSS.n4197 4.5005
R22100 DVSS.n4436 DVSS.n4194 4.5005
R22101 DVSS.n4436 DVSS.n4435 4.5005
R22102 DVSS.n4802 DVSS.n3716 4.5005
R22103 DVSS.n4802 DVSS.n4801 4.5005
R22104 DVSS.n4802 DVSS.n3715 4.5005
R22105 DVSS.n4803 DVSS.n4802 4.5005
R22106 DVSS.n4805 DVSS.n4804 4.5005
R22107 DVSS.n4805 DVSS.n3709 4.5005
R22108 DVSS.n4806 DVSS.n4805 4.5005
R22109 DVSS.n4822 DVSS.n4821 4.5005
R22110 DVSS.n4822 DVSS.n3673 4.5005
R22111 DVSS.n4823 DVSS.n4822 4.5005
R22112 DVSS.n4844 DVSS.n4824 4.5005
R22113 DVSS.n4844 DVSS.n4825 4.5005
R22114 DVSS.n4844 DVSS.n3667 4.5005
R22115 DVSS.n4845 DVSS.n4844 4.5005
R22116 DVSS.n4839 DVSS.n4838 4.5005
R22117 DVSS.n4838 DVSS.n4835 4.5005
R22118 DVSS.n4838 DVSS.n4833 4.5005
R22119 DVSS.n4838 DVSS.n4837 4.5005
R22120 DVSS.n4977 DVSS.n3590 4.5005
R22121 DVSS.n4977 DVSS.n4976 4.5005
R22122 DVSS.n4977 DVSS.n3596 4.5005
R22123 DVSS.n4978 DVSS.n4977 4.5005
R22124 DVSS.n4929 DVSS.n2911 4.5005
R22125 DVSS.n4931 DVSS.n2911 4.5005
R22126 DVSS.n4934 DVSS.n2911 4.5005
R22127 DVSS.n3885 DVSS.n3878 4.5005
R22128 DVSS.n4189 DVSS.n3885 4.5005
R22129 DVSS.n4004 DVSS.n4001 4.5005
R22130 DVSS.n4010 DVSS.n4001 4.5005
R22131 DVSS.n4101 DVSS.n3562 4.5005
R22132 DVSS.n5001 DVSS.n5000 4.5005
R22133 DVSS.n4998 DVSS.n3571 4.5005
R22134 DVSS.n4996 DVSS.n3571 4.5005
R22135 DVSS.n4994 DVSS.n3581 4.5005
R22136 DVSS.n4992 DVSS.n3581 4.5005
R22137 DVSS.n4991 DVSS.n4982 4.5005
R22138 DVSS.n4989 DVSS.n4982 4.5005
R22139 DVSS.n5919 DVSS.n5918 4.5005
R22140 DVSS.n5919 DVSS.n2918 4.5005
R22141 DVSS.n3875 DVSS.n3872 4.5005
R22142 DVSS.n3877 DVSS.n3872 4.5005
R22143 DVSS.n4099 DVSS.n4096 4.5005
R22144 DVSS.n5003 DVSS.n3564 4.5005
R22145 DVSS.n5918 DVSS.n5917 4.5005
R22146 DVSS.n3875 DVSS.n3874 4.5005
R22147 DVSS.n3877 DVSS.n3874 4.5005
R22148 DVSS.n3886 DVSS.n3878 4.5005
R22149 DVSS.n3886 DVSS.n3880 4.5005
R22150 DVSS.n3886 DVSS.n3870 4.5005
R22151 DVSS.n4189 DVSS.n3886 4.5005
R22152 DVSS.n4004 DVSS.n4002 4.5005
R22153 DVSS.n4008 DVSS.n4002 4.5005
R22154 DVSS.n4003 DVSS.n4002 4.5005
R22155 DVSS.n4010 DVSS.n4002 4.5005
R22156 DVSS.n4099 DVSS.n4097 4.5005
R22157 DVSS.n4097 DVSS.n3998 4.5005
R22158 DVSS.n4097 DVSS.n3562 4.5005
R22159 DVSS.n5003 DVSS.n3566 4.5005
R22160 DVSS.n3567 DVSS.n3566 4.5005
R22161 DVSS.n5001 DVSS.n3566 4.5005
R22162 DVSS.n4998 DVSS.n3572 4.5005
R22163 DVSS.n3575 DVSS.n3572 4.5005
R22164 DVSS.n3573 DVSS.n3572 4.5005
R22165 DVSS.n4996 DVSS.n3572 4.5005
R22166 DVSS.n4994 DVSS.n3582 4.5005
R22167 DVSS.n3585 DVSS.n3582 4.5005
R22168 DVSS.n3583 DVSS.n3582 4.5005
R22169 DVSS.n4992 DVSS.n3582 4.5005
R22170 DVSS.n4991 DVSS.n4983 4.5005
R22171 DVSS.n4986 DVSS.n4983 4.5005
R22172 DVSS.n4984 DVSS.n4983 4.5005
R22173 DVSS.n4989 DVSS.n4983 4.5005
R22174 DVSS.n5918 DVSS.n2916 4.5005
R22175 DVSS.n2918 DVSS.n2916 4.5005
R22176 DVSS.n5918 DVSS.n2915 4.5005
R22177 DVSS.n2918 DVSS.n2915 4.5005
R22178 DVSS.n3875 DVSS.n3871 4.5005
R22179 DVSS.n3877 DVSS.n3871 4.5005
R22180 DVSS.n4190 DVSS.n3878 4.5005
R22181 DVSS.n4190 DVSS.n3880 4.5005
R22182 DVSS.n4190 DVSS.n3870 4.5005
R22183 DVSS.n4190 DVSS.n4189 4.5005
R22184 DVSS.n4004 DVSS.n3999 4.5005
R22185 DVSS.n4008 DVSS.n3999 4.5005
R22186 DVSS.n4003 DVSS.n3999 4.5005
R22187 DVSS.n4010 DVSS.n3999 4.5005
R22188 DVSS.n4099 DVSS.n4094 4.5005
R22189 DVSS.n4094 DVSS.n3998 4.5005
R22190 DVSS.n4094 DVSS.n3562 4.5005
R22191 DVSS.n5003 DVSS.n3563 4.5005
R22192 DVSS.n3567 DVSS.n3563 4.5005
R22193 DVSS.n5001 DVSS.n3563 4.5005
R22194 DVSS.n4998 DVSS.n3569 4.5005
R22195 DVSS.n3575 DVSS.n3569 4.5005
R22196 DVSS.n3573 DVSS.n3569 4.5005
R22197 DVSS.n4996 DVSS.n3569 4.5005
R22198 DVSS.n4994 DVSS.n3579 4.5005
R22199 DVSS.n3585 DVSS.n3579 4.5005
R22200 DVSS.n3583 DVSS.n3579 4.5005
R22201 DVSS.n4992 DVSS.n3579 4.5005
R22202 DVSS.n4991 DVSS.n4980 4.5005
R22203 DVSS.n4986 DVSS.n4980 4.5005
R22204 DVSS.n4984 DVSS.n4980 4.5005
R22205 DVSS.n4989 DVSS.n4980 4.5005
R22206 DVSS.n5920 DVSS.n2915 4.5005
R22207 DVSS.n3876 DVSS.n3875 4.5005
R22208 DVSS.n3877 DVSS.n3876 4.5005
R22209 DVSS.n4188 DVSS.n3878 4.5005
R22210 DVSS.n4188 DVSS.n3880 4.5005
R22211 DVSS.n4188 DVSS.n3870 4.5005
R22212 DVSS.n4189 DVSS.n4188 4.5005
R22213 DVSS.n4009 DVSS.n4004 4.5005
R22214 DVSS.n4009 DVSS.n4008 4.5005
R22215 DVSS.n4009 DVSS.n4003 4.5005
R22216 DVSS.n4010 DVSS.n4009 4.5005
R22217 DVSS.n4099 DVSS.n4098 4.5005
R22218 DVSS.n4098 DVSS.n3998 4.5005
R22219 DVSS.n4098 DVSS.n3562 4.5005
R22220 DVSS.n5003 DVSS.n5002 4.5005
R22221 DVSS.n5002 DVSS.n3567 4.5005
R22222 DVSS.n5002 DVSS.n5001 4.5005
R22223 DVSS.n4998 DVSS.n4997 4.5005
R22224 DVSS.n4997 DVSS.n3575 4.5005
R22225 DVSS.n4997 DVSS.n3573 4.5005
R22226 DVSS.n4997 DVSS.n4996 4.5005
R22227 DVSS.n4994 DVSS.n4993 4.5005
R22228 DVSS.n4993 DVSS.n3585 4.5005
R22229 DVSS.n4993 DVSS.n3583 4.5005
R22230 DVSS.n4993 DVSS.n4992 4.5005
R22231 DVSS.n4991 DVSS.n4990 4.5005
R22232 DVSS.n4990 DVSS.n4986 4.5005
R22233 DVSS.n4990 DVSS.n4984 4.5005
R22234 DVSS.n4990 DVSS.n4989 4.5005
R22235 DVSS.n5920 DVSS.n2914 4.5005
R22236 DVSS.n5920 DVSS.n2916 4.5005
R22237 DVSS.n5920 DVSS.n5919 4.5005
R22238 DVSS.n3541 DVSS.n3111 4.5005
R22239 DVSS.n3547 DVSS.n3111 4.5005
R22240 DVSS.n3549 DVSS.n3156 4.5005
R22241 DVSS.n3555 DVSS.n3156 4.5005
R22242 DVSS.n3560 DVSS.n3188 4.5005
R22243 DVSS.n5030 DVSS.n5029 4.5005
R22244 DVSS.n3346 DVSS.n3324 4.5005
R22245 DVSS.n5387 DVSS.n3324 4.5005
R22246 DVSS.n5385 DVSS.n3353 4.5005
R22247 DVSS.n5383 DVSS.n3353 4.5005
R22248 DVSS.n5382 DVSS.n3363 4.5005
R22249 DVSS.n5380 DVSS.n3363 4.5005
R22250 DVSS.n5378 DVSS.n2956 4.5005
R22251 DVSS.n5373 DVSS.n2956 4.5005
R22252 DVSS.n3538 DVSS.n3534 4.5005
R22253 DVSS.n3540 DVSS.n3534 4.5005
R22254 DVSS.n3558 DVSS.n3556 4.5005
R22255 DVSS.n5027 DVSS.n5026 4.5005
R22256 DVSS.n5378 DVSS.n5371 4.5005
R22257 DVSS.n3538 DVSS.n3536 4.5005
R22258 DVSS.n3540 DVSS.n3536 4.5005
R22259 DVSS.n3541 DVSS.n3531 4.5005
R22260 DVSS.n3545 DVSS.n3531 4.5005
R22261 DVSS.n3532 DVSS.n3531 4.5005
R22262 DVSS.n3547 DVSS.n3531 4.5005
R22263 DVSS.n3549 DVSS.n3526 4.5005
R22264 DVSS.n3553 DVSS.n3526 4.5005
R22265 DVSS.n3527 DVSS.n3526 4.5005
R22266 DVSS.n3555 DVSS.n3526 4.5005
R22267 DVSS.n3558 DVSS.n3522 4.5005
R22268 DVSS.n3523 DVSS.n3522 4.5005
R22269 DVSS.n3560 DVSS.n3522 4.5005
R22270 DVSS.n5027 DVSS.n5024 4.5005
R22271 DVSS.n5025 DVSS.n5024 4.5005
R22272 DVSS.n5029 DVSS.n5024 4.5005
R22273 DVSS.n3346 DVSS.n3344 4.5005
R22274 DVSS.n5389 DVSS.n3344 4.5005
R22275 DVSS.n3349 DVSS.n3344 4.5005
R22276 DVSS.n5387 DVSS.n3344 4.5005
R22277 DVSS.n5385 DVSS.n3354 4.5005
R22278 DVSS.n3359 DVSS.n3354 4.5005
R22279 DVSS.n3356 DVSS.n3354 4.5005
R22280 DVSS.n5383 DVSS.n3354 4.5005
R22281 DVSS.n5382 DVSS.n3364 4.5005
R22282 DVSS.n3369 DVSS.n3364 4.5005
R22283 DVSS.n3366 DVSS.n3364 4.5005
R22284 DVSS.n5380 DVSS.n3364 4.5005
R22285 DVSS.n5378 DVSS.n5372 4.5005
R22286 DVSS.n5373 DVSS.n5372 4.5005
R22287 DVSS.n5378 DVSS.n5377 4.5005
R22288 DVSS.n5377 DVSS.n5373 4.5005
R22289 DVSS.n3538 DVSS.n3533 4.5005
R22290 DVSS.n3540 DVSS.n3533 4.5005
R22291 DVSS.n3541 DVSS.n3529 4.5005
R22292 DVSS.n3545 DVSS.n3529 4.5005
R22293 DVSS.n3532 DVSS.n3529 4.5005
R22294 DVSS.n3547 DVSS.n3529 4.5005
R22295 DVSS.n3549 DVSS.n3524 4.5005
R22296 DVSS.n3553 DVSS.n3524 4.5005
R22297 DVSS.n3527 DVSS.n3524 4.5005
R22298 DVSS.n3555 DVSS.n3524 4.5005
R22299 DVSS.n3558 DVSS.n3520 4.5005
R22300 DVSS.n3523 DVSS.n3520 4.5005
R22301 DVSS.n3560 DVSS.n3520 4.5005
R22302 DVSS.n5027 DVSS.n5022 4.5005
R22303 DVSS.n5025 DVSS.n5022 4.5005
R22304 DVSS.n5029 DVSS.n5022 4.5005
R22305 DVSS.n3347 DVSS.n3346 4.5005
R22306 DVSS.n5389 DVSS.n3347 4.5005
R22307 DVSS.n3349 DVSS.n3347 4.5005
R22308 DVSS.n5387 DVSS.n3347 4.5005
R22309 DVSS.n5385 DVSS.n3351 4.5005
R22310 DVSS.n3359 DVSS.n3351 4.5005
R22311 DVSS.n3356 DVSS.n3351 4.5005
R22312 DVSS.n5383 DVSS.n3351 4.5005
R22313 DVSS.n5382 DVSS.n3361 4.5005
R22314 DVSS.n3369 DVSS.n3361 4.5005
R22315 DVSS.n3366 DVSS.n3361 4.5005
R22316 DVSS.n5380 DVSS.n3361 4.5005
R22317 DVSS.n5377 DVSS.n5376 4.5005
R22318 DVSS.n3539 DVSS.n3538 4.5005
R22319 DVSS.n3540 DVSS.n3539 4.5005
R22320 DVSS.n3546 DVSS.n3541 4.5005
R22321 DVSS.n3546 DVSS.n3545 4.5005
R22322 DVSS.n3546 DVSS.n3532 4.5005
R22323 DVSS.n3547 DVSS.n3546 4.5005
R22324 DVSS.n3554 DVSS.n3549 4.5005
R22325 DVSS.n3554 DVSS.n3553 4.5005
R22326 DVSS.n3554 DVSS.n3527 4.5005
R22327 DVSS.n3555 DVSS.n3554 4.5005
R22328 DVSS.n3559 DVSS.n3558 4.5005
R22329 DVSS.n3559 DVSS.n3523 4.5005
R22330 DVSS.n3560 DVSS.n3559 4.5005
R22331 DVSS.n5028 DVSS.n5027 4.5005
R22332 DVSS.n5028 DVSS.n5025 4.5005
R22333 DVSS.n5029 DVSS.n5028 4.5005
R22334 DVSS.n5388 DVSS.n3346 4.5005
R22335 DVSS.n5389 DVSS.n5388 4.5005
R22336 DVSS.n5388 DVSS.n3349 4.5005
R22337 DVSS.n5388 DVSS.n5387 4.5005
R22338 DVSS.n5385 DVSS.n5384 4.5005
R22339 DVSS.n5384 DVSS.n3359 4.5005
R22340 DVSS.n5384 DVSS.n3356 4.5005
R22341 DVSS.n5384 DVSS.n5383 4.5005
R22342 DVSS.n5382 DVSS.n5381 4.5005
R22343 DVSS.n5381 DVSS.n3369 4.5005
R22344 DVSS.n5381 DVSS.n3366 4.5005
R22345 DVSS.n5381 DVSS.n5380 4.5005
R22346 DVSS.n5376 DVSS.n5375 4.5005
R22347 DVSS.n5376 DVSS.n5372 4.5005
R22348 DVSS.n5376 DVSS.n2956 4.5005
R22349 DVSS.n5677 DVSS.n5671 4.5005
R22350 DVSS.n5683 DVSS.n3250 4.5005
R22351 DVSS.n5690 DVSS.n3241 4.5005
R22352 DVSS.n5691 DVSS.n3236 4.5005
R22353 DVSS.n5694 DVSS.n3236 4.5005
R22354 DVSS.n5491 DVSS.n5485 4.5005
R22355 DVSS.n5494 DVSS.n5485 4.5005
R22356 DVSS.n5500 DVSS.n3293 4.5005
R22357 DVSS.n5507 DVSS.n3301 4.5005
R22358 DVSS.n5516 DVSS.n5515 4.5005
R22359 DVSS.n5906 DVSS.n2960 4.5005
R22360 DVSS.n5681 DVSS.n3248 4.5005
R22361 DVSS.n5683 DVSS.n3248 4.5005
R22362 DVSS.n5688 DVSS.n3239 4.5005
R22363 DVSS.n5690 DVSS.n3239 4.5005
R22364 DVSS.n5694 DVSS.n3233 4.5005
R22365 DVSS.n5494 DVSS.n5404 4.5005
R22366 DVSS.n5498 DVSS.n5397 4.5005
R22367 DVSS.n5500 DVSS.n5397 4.5005
R22368 DVSS.n5505 DVSS.n3317 4.5005
R22369 DVSS.n5507 DVSS.n3317 4.5005
R22370 DVSS.n5513 DVSS.n3312 4.5005
R22371 DVSS.n5515 DVSS.n3312 4.5005
R22372 DVSS.n5681 DVSS.n3251 4.5005
R22373 DVSS.n5683 DVSS.n3251 4.5005
R22374 DVSS.n5688 DVSS.n3242 4.5005
R22375 DVSS.n5690 DVSS.n3242 4.5005
R22376 DVSS.n5694 DVSS.n5693 4.5005
R22377 DVSS.n5494 DVSS.n5493 4.5005
R22378 DVSS.n5498 DVSS.n5398 4.5005
R22379 DVSS.n5500 DVSS.n5398 4.5005
R22380 DVSS.n5505 DVSS.n3318 4.5005
R22381 DVSS.n5507 DVSS.n3318 4.5005
R22382 DVSS.n5513 DVSS.n3313 4.5005
R22383 DVSS.n5515 DVSS.n3313 4.5005
R22384 DVSS.n5909 DVSS.n5908 4.5005
R22385 DVSS.n5908 DVSS.n2960 4.5005
R22386 DVSS.n5910 DVSS.n5909 4.5005
R22387 DVSS.n5910 DVSS.n2960 4.5005
R22388 DVSS.n5683 DVSS.n3113 4.5005
R22389 DVSS.n5690 DVSS.n3157 4.5005
R22390 DVSS.n5500 DVSS.n5395 4.5005
R22391 DVSS.n5507 DVSS.n3315 4.5005
R22392 DVSS.n5515 DVSS.n3311 4.5005
R22393 DVSS.n5677 DVSS.n5676 4.5005
R22394 DVSS.n5682 DVSS.n5681 4.5005
R22395 DVSS.n5683 DVSS.n5682 4.5005
R22396 DVSS.n5689 DVSS.n5688 4.5005
R22397 DVSS.n5690 DVSS.n5689 4.5005
R22398 DVSS.n5691 DVSS.n3231 4.5005
R22399 DVSS.n5491 DVSS.n5490 4.5005
R22400 DVSS.n5499 DVSS.n5498 4.5005
R22401 DVSS.n5500 DVSS.n5499 4.5005
R22402 DVSS.n5506 DVSS.n5505 4.5005
R22403 DVSS.n5507 DVSS.n5506 4.5005
R22404 DVSS.n5514 DVSS.n5513 4.5005
R22405 DVSS.n5515 DVSS.n5514 4.5005
R22406 DVSS.n5908 DVSS.n5907 4.5005
R22407 DVSS.n5907 DVSS.n5906 4.5005
R22408 DVSS.n5668 DVSS.n5667 4.5005
R22409 DVSS.n5661 DVSS.n5657 4.5005
R22410 DVSS.n5651 DVSS.n5647 4.5005
R22411 DVSS.n5645 DVSS.n3275 4.5005
R22412 DVSS.n3281 DVSS.n3275 4.5005
R22413 DVSS.n5633 DVSS.n5631 4.5005
R22414 DVSS.n5636 DVSS.n5631 4.5005
R22415 DVSS.n5544 DVSS.n5540 4.5005
R22416 DVSS.n5534 DVSS.n5530 4.5005
R22417 DVSS.n5525 DVSS.n5521 4.5005
R22418 DVSS.n5901 DVSS.n2969 4.5005
R22419 DVSS.n5659 DVSS.n3265 4.5005
R22420 DVSS.n5661 DVSS.n3265 4.5005
R22421 DVSS.n5649 DVSS.n3272 4.5005
R22422 DVSS.n5651 DVSS.n3272 4.5005
R22423 DVSS.n3281 DVSS.n3279 4.5005
R22424 DVSS.n5636 DVSS.n3289 4.5005
R22425 DVSS.n5542 DVSS.n3296 4.5005
R22426 DVSS.n5544 DVSS.n3296 4.5005
R22427 DVSS.n5532 DVSS.n3304 4.5005
R22428 DVSS.n5534 DVSS.n3304 4.5005
R22429 DVSS.n5523 DVSS.n5519 4.5005
R22430 DVSS.n5525 DVSS.n5519 4.5005
R22431 DVSS.n5660 DVSS.n5659 4.5005
R22432 DVSS.n5661 DVSS.n5660 4.5005
R22433 DVSS.n5650 DVSS.n5649 4.5005
R22434 DVSS.n5651 DVSS.n5650 4.5005
R22435 DVSS.n3281 DVSS.n3280 4.5005
R22436 DVSS.n5636 DVSS.n5635 4.5005
R22437 DVSS.n5543 DVSS.n5542 4.5005
R22438 DVSS.n5544 DVSS.n5543 4.5005
R22439 DVSS.n5533 DVSS.n5532 4.5005
R22440 DVSS.n5534 DVSS.n5533 4.5005
R22441 DVSS.n5524 DVSS.n5523 4.5005
R22442 DVSS.n5525 DVSS.n5524 4.5005
R22443 DVSS.n5904 DVSS.n5903 4.5005
R22444 DVSS.n5903 DVSS.n2969 4.5005
R22445 DVSS.n5905 DVSS.n5904 4.5005
R22446 DVSS.n5905 DVSS.n2969 4.5005
R22447 DVSS.n5662 DVSS.n5661 4.5005
R22448 DVSS.n5652 DVSS.n5651 4.5005
R22449 DVSS.n5545 DVSS.n5544 4.5005
R22450 DVSS.n5535 DVSS.n5534 4.5005
R22451 DVSS.n5526 DVSS.n5525 4.5005
R22452 DVSS.n5669 DVSS.n5668 4.5005
R22453 DVSS.n5659 DVSS.n3262 4.5005
R22454 DVSS.n5661 DVSS.n3262 4.5005
R22455 DVSS.n5649 DVSS.n3269 4.5005
R22456 DVSS.n5651 DVSS.n3269 4.5005
R22457 DVSS.n5645 DVSS.n5644 4.5005
R22458 DVSS.n5633 DVSS.n3287 4.5005
R22459 DVSS.n5542 DVSS.n3292 4.5005
R22460 DVSS.n5544 DVSS.n3292 4.5005
R22461 DVSS.n5532 DVSS.n3300 4.5005
R22462 DVSS.n5534 DVSS.n3300 4.5005
R22463 DVSS.n5523 DVSS.n3307 4.5005
R22464 DVSS.n5525 DVSS.n3307 4.5005
R22465 DVSS.n5903 DVSS.n5902 4.5005
R22466 DVSS.n5902 DVSS.n5901 4.5005
R22467 DVSS.n2680 DVSS.n2594 4.5005
R22468 DVSS.n2686 DVSS.n2601 4.5005
R22469 DVSS.n2693 DVSS.n2609 4.5005
R22470 DVSS.n7271 DVSS.n2694 4.5005
R22471 DVSS.n7271 DVSS.n7270 4.5005
R22472 DVSS.n2754 DVSS.n2704 4.5005
R22473 DVSS.n2751 DVSS.n2704 4.5005
R22474 DVSS.n2746 DVSS.n2086 4.5005
R22475 DVSS.n2740 DVSS.n2094 4.5005
R22476 DVSS.n2735 DVSS.n2102 4.5005
R22477 DVSS.n7699 DVSS.n2109 4.5005
R22478 DVSS.n2678 DVSS.n2670 4.5005
R22479 DVSS.n2680 DVSS.n2670 4.5005
R22480 DVSS.n2684 DVSS.n2663 4.5005
R22481 DVSS.n2686 DVSS.n2663 4.5005
R22482 DVSS.n2691 DVSS.n2655 4.5005
R22483 DVSS.n2693 DVSS.n2655 4.5005
R22484 DVSS.n7270 DVSS.n2698 4.5005
R22485 DVSS.n2751 DVSS.n2708 4.5005
R22486 DVSS.n2716 DVSS.n2712 4.5005
R22487 DVSS.n2746 DVSS.n2716 4.5005
R22488 DVSS.n2725 DVSS.n2721 4.5005
R22489 DVSS.n2740 DVSS.n2725 4.5005
R22490 DVSS.n2733 DVSS.n2729 4.5005
R22491 DVSS.n2735 DVSS.n2733 4.5005
R22492 DVSS.n2678 DVSS.n2671 4.5005
R22493 DVSS.n2680 DVSS.n2671 4.5005
R22494 DVSS.n2684 DVSS.n2664 4.5005
R22495 DVSS.n2686 DVSS.n2664 4.5005
R22496 DVSS.n2691 DVSS.n2656 4.5005
R22497 DVSS.n2693 DVSS.n2656 4.5005
R22498 DVSS.n7270 DVSS.n7269 4.5005
R22499 DVSS.n2751 DVSS.n2750 4.5005
R22500 DVSS.n2745 DVSS.n2712 4.5005
R22501 DVSS.n2746 DVSS.n2745 4.5005
R22502 DVSS.n2739 DVSS.n2721 4.5005
R22503 DVSS.n2740 DVSS.n2739 4.5005
R22504 DVSS.n2734 DVSS.n2729 4.5005
R22505 DVSS.n2735 DVSS.n2734 4.5005
R22506 DVSS.n7697 DVSS.n7696 4.5005
R22507 DVSS.n7697 DVSS.n2109 4.5005
R22508 DVSS.n7696 DVSS.n7695 4.5005
R22509 DVSS.n7695 DVSS.n2109 4.5005
R22510 DVSS.n2680 DVSS.n2521 4.5005
R22511 DVSS.n2686 DVSS.n2464 4.5005
R22512 DVSS.n2693 DVSS.n2400 4.5005
R22513 DVSS.n2746 DVSS.n2252 4.5005
R22514 DVSS.n2740 DVSS.n2210 4.5005
R22515 DVSS.n2735 DVSS.n2176 4.5005
R22516 DVSS.n2679 DVSS.n2678 4.5005
R22517 DVSS.n2680 DVSS.n2679 4.5005
R22518 DVSS.n2685 DVSS.n2684 4.5005
R22519 DVSS.n2686 DVSS.n2685 4.5005
R22520 DVSS.n2692 DVSS.n2691 4.5005
R22521 DVSS.n2693 DVSS.n2692 4.5005
R22522 DVSS.n7266 DVSS.n2694 4.5005
R22523 DVSS.n2754 DVSS.n2753 4.5005
R22524 DVSS.n2747 DVSS.n2712 4.5005
R22525 DVSS.n2747 DVSS.n2746 4.5005
R22526 DVSS.n2741 DVSS.n2721 4.5005
R22527 DVSS.n2741 DVSS.n2740 4.5005
R22528 DVSS.n2736 DVSS.n2729 4.5005
R22529 DVSS.n2736 DVSS.n2735 4.5005
R22530 DVSS.n7698 DVSS.n7697 4.5005
R22531 DVSS.n7699 DVSS.n7698 4.5005
R22532 DVSS.n7358 DVSS.n7354 4.5005
R22533 DVSS.n7349 DVSS.n7345 4.5005
R22534 DVSS.n7339 DVSS.n7335 4.5005
R22535 DVSS.n7333 DVSS.n2615 4.5005
R22536 DVSS.n2621 DVSS.n2615 4.5005
R22537 DVSS.n7861 DVSS.n2079 4.5005
R22538 DVSS.n7861 DVSS.n7860 4.5005
R22539 DVSS.n7852 DVSS.n7848 4.5005
R22540 DVSS.n7722 DVSS.n1814 4.5005
R22541 DVSS.n7715 DVSS.n7711 4.5005
R22542 DVSS.n7704 DVSS.n7700 4.5005
R22543 DVSS.n7356 DVSS.n2597 4.5005
R22544 DVSS.n7358 DVSS.n2597 4.5005
R22545 DVSS.n7347 DVSS.n2604 4.5005
R22546 DVSS.n7349 DVSS.n2604 4.5005
R22547 DVSS.n7337 DVSS.n2612 4.5005
R22548 DVSS.n7339 DVSS.n2612 4.5005
R22549 DVSS.n2621 DVSS.n2619 4.5005
R22550 DVSS.n7860 DVSS.n2082 4.5005
R22551 DVSS.n7850 DVSS.n2089 4.5005
R22552 DVSS.n7852 DVSS.n2089 4.5005
R22553 DVSS.n7720 DVSS.n2098 4.5005
R22554 DVSS.n7722 DVSS.n2098 4.5005
R22555 DVSS.n7713 DVSS.n2105 4.5005
R22556 DVSS.n7715 DVSS.n2105 4.5005
R22557 DVSS.n7357 DVSS.n7356 4.5005
R22558 DVSS.n7358 DVSS.n7357 4.5005
R22559 DVSS.n7348 DVSS.n7347 4.5005
R22560 DVSS.n7349 DVSS.n7348 4.5005
R22561 DVSS.n7338 DVSS.n7337 4.5005
R22562 DVSS.n7339 DVSS.n7338 4.5005
R22563 DVSS.n2621 DVSS.n2620 4.5005
R22564 DVSS.n7860 DVSS.n7859 4.5005
R22565 DVSS.n7851 DVSS.n7850 4.5005
R22566 DVSS.n7852 DVSS.n7851 4.5005
R22567 DVSS.n7721 DVSS.n7720 4.5005
R22568 DVSS.n7722 DVSS.n7721 4.5005
R22569 DVSS.n7714 DVSS.n7713 4.5005
R22570 DVSS.n7715 DVSS.n7714 4.5005
R22571 DVSS.n7708 DVSS.n2108 4.5005
R22572 DVSS.n7700 DVSS.n2108 4.5005
R22573 DVSS.n7708 DVSS.n7707 4.5005
R22574 DVSS.n7707 DVSS.n7700 4.5005
R22575 DVSS.n7359 DVSS.n7358 4.5005
R22576 DVSS.n7350 DVSS.n7349 4.5005
R22577 DVSS.n7340 DVSS.n7339 4.5005
R22578 DVSS.n7853 DVSS.n7852 4.5005
R22579 DVSS.n7723 DVSS.n7722 4.5005
R22580 DVSS.n7716 DVSS.n7715 4.5005
R22581 DVSS.n7356 DVSS.n2593 4.5005
R22582 DVSS.n7358 DVSS.n2593 4.5005
R22583 DVSS.n7347 DVSS.n2600 4.5005
R22584 DVSS.n7349 DVSS.n2600 4.5005
R22585 DVSS.n7337 DVSS.n2608 4.5005
R22586 DVSS.n7339 DVSS.n2608 4.5005
R22587 DVSS.n7333 DVSS.n7332 4.5005
R22588 DVSS.n7856 DVSS.n2079 4.5005
R22589 DVSS.n7850 DVSS.n2085 4.5005
R22590 DVSS.n7852 DVSS.n2085 4.5005
R22591 DVSS.n7720 DVSS.n2093 4.5005
R22592 DVSS.n7722 DVSS.n2093 4.5005
R22593 DVSS.n7713 DVSS.n2101 4.5005
R22594 DVSS.n7715 DVSS.n2101 4.5005
R22595 DVSS.n7705 DVSS.n2108 4.5005
R22596 DVSS.n7705 DVSS.n7704 4.5005
R22597 DVSS.n8076 DVSS.n1904 4.5005
R22598 DVSS.n8082 DVSS.n1895 4.5005
R22599 DVSS.n8089 DVSS.n1885 4.5005
R22600 DVSS.n8090 DVSS.n1879 4.5005
R22601 DVSS.n8093 DVSS.n1879 4.5005
R22602 DVSS.n8102 DVSS.n1868 4.5005
R22603 DVSS.n8105 DVSS.n1868 4.5005
R22604 DVSS.n8111 DVSS.n1859 4.5005
R22605 DVSS.n8118 DVSS.n1553 4.5005
R22606 DVSS.n1848 DVSS.n1560 4.5005
R22607 DVSS.n8183 DVSS.n1756 4.5005
R22608 DVSS.n8074 DVSS.n1902 4.5005
R22609 DVSS.n8076 DVSS.n1902 4.5005
R22610 DVSS.n8080 DVSS.n1893 4.5005
R22611 DVSS.n8082 DVSS.n1893 4.5005
R22612 DVSS.n8087 DVSS.n1883 4.5005
R22613 DVSS.n8089 DVSS.n1883 4.5005
R22614 DVSS.n8093 DVSS.n1877 4.5005
R22615 DVSS.n8105 DVSS.n1866 4.5005
R22616 DVSS.n8109 DVSS.n1857 4.5005
R22617 DVSS.n8111 DVSS.n1857 4.5005
R22618 DVSS.n8116 DVSS.n1837 4.5005
R22619 DVSS.n8118 DVSS.n1837 4.5005
R22620 DVSS.n1846 DVSS.n1844 4.5005
R22621 DVSS.n1848 DVSS.n1844 4.5005
R22622 DVSS.n8074 DVSS.n1905 4.5005
R22623 DVSS.n8076 DVSS.n1905 4.5005
R22624 DVSS.n8080 DVSS.n1896 4.5005
R22625 DVSS.n8082 DVSS.n1896 4.5005
R22626 DVSS.n8087 DVSS.n1886 4.5005
R22627 DVSS.n8089 DVSS.n1886 4.5005
R22628 DVSS.n8093 DVSS.n8092 4.5005
R22629 DVSS.n8105 DVSS.n8104 4.5005
R22630 DVSS.n8109 DVSS.n1860 4.5005
R22631 DVSS.n8111 DVSS.n1860 4.5005
R22632 DVSS.n8116 DVSS.n1852 4.5005
R22633 DVSS.n8118 DVSS.n1852 4.5005
R22634 DVSS.n1847 DVSS.n1846 4.5005
R22635 DVSS.n1848 DVSS.n1847 4.5005
R22636 DVSS.n8181 DVSS.n1755 4.5005
R22637 DVSS.n1756 DVSS.n1755 4.5005
R22638 DVSS.n8181 DVSS.n8180 4.5005
R22639 DVSS.n8180 DVSS.n1756 4.5005
R22640 DVSS.n8076 DVSS.n1901 4.5005
R22641 DVSS.n8082 DVSS.n1892 4.5005
R22642 DVSS.n8089 DVSS.n1882 4.5005
R22643 DVSS.n8111 DVSS.n1856 4.5005
R22644 DVSS.n8119 DVSS.n8118 4.5005
R22645 DVSS.n1849 DVSS.n1848 4.5005
R22646 DVSS.n8075 DVSS.n8074 4.5005
R22647 DVSS.n8076 DVSS.n8075 4.5005
R22648 DVSS.n8081 DVSS.n8080 4.5005
R22649 DVSS.n8082 DVSS.n8081 4.5005
R22650 DVSS.n8088 DVSS.n8087 4.5005
R22651 DVSS.n8089 DVSS.n8088 4.5005
R22652 DVSS.n8090 DVSS.n1875 4.5005
R22653 DVSS.n8102 DVSS.n8101 4.5005
R22654 DVSS.n8110 DVSS.n8109 4.5005
R22655 DVSS.n8111 DVSS.n8110 4.5005
R22656 DVSS.n8117 DVSS.n8116 4.5005
R22657 DVSS.n8118 DVSS.n8117 4.5005
R22658 DVSS.n1846 DVSS.n1840 4.5005
R22659 DVSS.n1848 DVSS.n1840 4.5005
R22660 DVSS.n8184 DVSS.n1755 4.5005
R22661 DVSS.n8184 DVSS.n8183 4.5005
R22662 DVSS.n7066 DVSS.n6662 4.5005
R22663 DVSS.n7066 DVSS.n7065 4.5005
R22664 DVSS.n7067 DVSS.n7066 4.5005
R22665 DVSS.n7132 DVSS.n7068 4.5005
R22666 DVSS.n7132 DVSS.n7131 4.5005
R22667 DVSS.n7133 DVSS.n7132 4.5005
R22668 DVSS.n7065 DVSS.n6659 4.5005
R22669 DVSS.n7067 DVSS.n6659 4.5005
R22670 DVSS.n7131 DVSS.n6655 4.5005
R22671 DVSS.n7133 DVSS.n6655 4.5005
R22672 DVSS.n7131 DVSS.n7130 4.5005
R22673 DVSS.n7130 DVSS.n7068 4.5005
R22674 DVSS.n7065 DVSS.n7064 4.5005
R22675 DVSS.n7064 DVSS.n6662 4.5005
R22676 DVSS.n6750 DVSS.n1914 4.5005
R22677 DVSS.n6752 DVSS.n1914 4.5005
R22678 DVSS.n8069 DVSS.n1911 4.5005
R22679 DVSS.n8069 DVSS.n1910 4.5005
R22680 DVSS.n7368 DVSS.n7364 4.5005
R22681 DVSS.n7369 DVSS.n7368 4.5005
R22682 DVSS.n7373 DVSS.n2584 4.5005
R22683 DVSS.n7374 DVSS.n7373 4.5005
R22684 DVSS.n5893 DVSS.n2989 4.5005
R22685 DVSS.n5893 DVSS.n2986 4.5005
R22686 DVSS.n5887 DVSS.n2991 4.5005
R22687 DVSS.n5885 DVSS.n2991 4.5005
R22688 DVSS.n3015 DVSS.n3013 4.5005
R22689 DVSS.n5876 DVSS.n5873 4.5005
R22690 DVSS.n5876 DVSS.n5875 4.5005
R22691 DVSS.n5875 DVSS.n3014 4.5005
R22692 DVSS.n5875 DVSS.n3015 4.5005
R22693 DVSS.n5867 DVSS.n5866 4.5005
R22694 DVSS.n5869 DVSS.n3018 4.5005
R22695 DVSS.n5869 DVSS.n3020 4.5005
R22696 DVSS.n3022 DVSS.n3020 4.5005
R22697 DVSS.n5867 DVSS.n3020 4.5005
R22698 DVSS.n4445 DVSS.n4442 4.5005
R22699 DVSS.n4448 DVSS.n4444 4.5005
R22700 DVSS.n4448 DVSS.n4447 4.5005
R22701 DVSS.n4447 DVSS.n3857 4.5005
R22702 DVSS.n4447 DVSS.n4442 4.5005
R22703 DVSS.n4475 DVSS.n4474 4.5005
R22704 DVSS.n4478 DVSS.n4477 4.5005
R22705 DVSS.n4442 DVSS.n3853 4.5005
R22706 DVSS.n3857 DVSS.n3853 4.5005
R22707 DVSS.n4448 DVSS.n3853 4.5005
R22708 DVSS.n4449 DVSS.n4442 4.5005
R22709 DVSS.n4449 DVSS.n3857 4.5005
R22710 DVSS.n4449 DVSS.n4448 4.5005
R22711 DVSS.n5867 DVSS.n3017 4.5005
R22712 DVSS.n3022 DVSS.n3017 4.5005
R22713 DVSS.n5869 DVSS.n3017 4.5005
R22714 DVSS.n5868 DVSS.n5867 4.5005
R22715 DVSS.n5868 DVSS.n3022 4.5005
R22716 DVSS.n5869 DVSS.n5868 4.5005
R22717 DVSS.n5877 DVSS.n3015 4.5005
R22718 DVSS.n5877 DVSS.n3014 4.5005
R22719 DVSS.n5877 DVSS.n5876 4.5005
R22720 DVSS.n3015 DVSS.n2993 4.5005
R22721 DVSS.n3014 DVSS.n2993 4.5005
R22722 DVSS.n5876 DVSS.n2993 4.5005
R22723 DVSS.n5884 DVSS.n2991 4.5005
R22724 DVSS.n5890 DVSS.n2991 4.5005
R22725 DVSS.n5890 DVSS.n5889 4.5005
R22726 DVSS.n5893 DVSS.n2985 4.5005
R22727 DVSS.n5894 DVSS.n5893 4.5005
R22728 DVSS.n5895 DVSS.n5894 4.5005
R22729 DVSS.n7373 DVSS.n2581 4.5005
R22730 DVSS.n7373 DVSS.n7372 4.5005
R22731 DVSS.n7372 DVSS.n2579 4.5005
R22732 DVSS.n7368 DVSS.n2590 4.5005
R22733 DVSS.n7368 DVSS.n7367 4.5005
R22734 DVSS.n7367 DVSS.n2588 4.5005
R22735 DVSS.n8069 DVSS.n1909 4.5005
R22736 DVSS.n8069 DVSS.n8068 4.5005
R22737 DVSS.n8068 DVSS.n8067 4.5005
R22738 DVSS.n6753 DVSS.n6752 4.5005
R22739 DVSS.n4477 DVSS.n4460 4.5005
R22740 DVSS.n4463 DVSS.n4460 4.5005
R22741 DVSS.n4492 DVSS.n4454 4.5005
R22742 DVSS.n4454 DVSS.n3834 4.5005
R22743 DVSS.n4490 DVSS.n4454 4.5005
R22744 DVSS.n4461 DVSS.n4454 4.5005
R22745 DVSS.n4492 DVSS.n4455 4.5005
R22746 DVSS.n4455 DVSS.n3834 4.5005
R22747 DVSS.n4461 DVSS.n4455 4.5005
R22748 DVSS.n4487 DVSS.n3834 4.5005
R22749 DVSS.n4487 DVSS.n4461 4.5005
R22750 DVSS.n4485 DVSS.n3834 4.5005
R22751 DVSS.n4485 DVSS.n4461 4.5005
R22752 DVSS.n4484 DVSS.n3834 4.5005
R22753 DVSS.n4484 DVSS.n4461 4.5005
R22754 DVSS.n4482 DVSS.n3834 4.5005
R22755 DVSS.n4482 DVSS.n4461 4.5005
R22756 DVSS.n4492 DVSS.n4453 4.5005
R22757 DVSS.n4453 DVSS.n3834 4.5005
R22758 DVSS.n4461 DVSS.n4453 4.5005
R22759 DVSS.n4452 DVSS.n3837 4.5005
R22760 DVSS.n4452 DVSS.n3838 4.5005
R22761 DVSS.n4452 DVSS.n4451 4.5005
R22762 DVSS.n3844 DVSS.n3838 4.5005
R22763 DVSS.n4451 DVSS.n3844 4.5005
R22764 DVSS.n3847 DVSS.n3838 4.5005
R22765 DVSS.n4451 DVSS.n3847 4.5005
R22766 DVSS.n3843 DVSS.n3838 4.5005
R22767 DVSS.n4451 DVSS.n3843 4.5005
R22768 DVSS.n3849 DVSS.n3838 4.5005
R22769 DVSS.n4451 DVSS.n3849 4.5005
R22770 DVSS.n3842 DVSS.n3838 4.5005
R22771 DVSS.n4451 DVSS.n3842 4.5005
R22772 DVSS.n3851 DVSS.n3838 4.5005
R22773 DVSS.n3856 DVSS.n3851 4.5005
R22774 DVSS.n4451 DVSS.n3851 4.5005
R22775 DVSS.n3856 DVSS.n3841 4.5005
R22776 DVSS.n4451 DVSS.n3841 4.5005
R22777 DVSS.n3841 DVSS.n3838 4.5005
R22778 DVSS.n3841 DVSS.n3837 4.5005
R22779 DVSS.n3852 DVSS.n3837 4.5005
R22780 DVSS.n3852 DVSS.n3838 4.5005
R22781 DVSS.n3856 DVSS.n3852 4.5005
R22782 DVSS.n4451 DVSS.n3852 4.5005
R22783 DVSS.n3840 DVSS.n3837 4.5005
R22784 DVSS.n3840 DVSS.n3838 4.5005
R22785 DVSS.n3856 DVSS.n3840 4.5005
R22786 DVSS.n4451 DVSS.n3840 4.5005
R22787 DVSS.n4450 DVSS.n3837 4.5005
R22788 DVSS.n4450 DVSS.n3838 4.5005
R22789 DVSS.n4450 DVSS.n3856 4.5005
R22790 DVSS.n4451 DVSS.n4450 4.5005
R22791 DVSS.n5855 DVSS.n3027 4.5005
R22792 DVSS.n5864 DVSS.n5855 4.5005
R22793 DVSS.n5855 DVSS.n3029 4.5005
R22794 DVSS.n5855 DVSS.n3028 4.5005
R22795 DVSS.n3027 DVSS.n3026 4.5005
R22796 DVSS.n5864 DVSS.n3026 4.5005
R22797 DVSS.n3029 DVSS.n3026 4.5005
R22798 DVSS.n3028 DVSS.n3026 4.5005
R22799 DVSS.n5865 DVSS.n3028 4.5005
R22800 DVSS.n5865 DVSS.n3029 4.5005
R22801 DVSS.n5865 DVSS.n3027 4.5005
R22802 DVSS.n5865 DVSS.n5864 4.5005
R22803 DVSS.n3028 DVSS.n3021 4.5005
R22804 DVSS.n3029 DVSS.n3021 4.5005
R22805 DVSS.n3027 DVSS.n3021 4.5005
R22806 DVSS.n5864 DVSS.n3021 4.5005
R22807 DVSS.n3028 DVSS.n3023 4.5005
R22808 DVSS.n3029 DVSS.n3023 4.5005
R22809 DVSS.n5864 DVSS.n3023 4.5005
R22810 DVSS.n3034 DVSS.n3029 4.5005
R22811 DVSS.n5864 DVSS.n3034 4.5005
R22812 DVSS.n5858 DVSS.n3029 4.5005
R22813 DVSS.n5864 DVSS.n5858 4.5005
R22814 DVSS.n3032 DVSS.n3029 4.5005
R22815 DVSS.n5864 DVSS.n3032 4.5005
R22816 DVSS.n5861 DVSS.n3029 4.5005
R22817 DVSS.n5864 DVSS.n5861 4.5005
R22818 DVSS.n3031 DVSS.n3029 4.5005
R22819 DVSS.n5864 DVSS.n3031 4.5005
R22820 DVSS.n5863 DVSS.n3029 4.5005
R22821 DVSS.n5863 DVSS.n3027 4.5005
R22822 DVSS.n5864 DVSS.n5863 4.5005
R22823 DVSS.n3005 DVSS.n2995 4.5005
R22824 DVSS.n3005 DVSS.n2996 4.5005
R22825 DVSS.n5879 DVSS.n3005 4.5005
R22826 DVSS.n3002 DVSS.n2996 4.5005
R22827 DVSS.n5879 DVSS.n3002 4.5005
R22828 DVSS.n3008 DVSS.n2996 4.5005
R22829 DVSS.n5879 DVSS.n3008 4.5005
R22830 DVSS.n3001 DVSS.n2996 4.5005
R22831 DVSS.n5879 DVSS.n3001 4.5005
R22832 DVSS.n3011 DVSS.n2996 4.5005
R22833 DVSS.n5879 DVSS.n3011 4.5005
R22834 DVSS.n3000 DVSS.n2995 4.5005
R22835 DVSS.n3000 DVSS.n2996 4.5005
R22836 DVSS.n5879 DVSS.n3000 4.5005
R22837 DVSS.n3012 DVSS.n2994 4.5005
R22838 DVSS.n5879 DVSS.n3012 4.5005
R22839 DVSS.n3012 DVSS.n2996 4.5005
R22840 DVSS.n3012 DVSS.n2995 4.5005
R22841 DVSS.n2999 DVSS.n2994 4.5005
R22842 DVSS.n5879 DVSS.n2999 4.5005
R22843 DVSS.n2999 DVSS.n2996 4.5005
R22844 DVSS.n2999 DVSS.n2995 4.5005
R22845 DVSS.n5878 DVSS.n2994 4.5005
R22846 DVSS.n5879 DVSS.n5878 4.5005
R22847 DVSS.n5878 DVSS.n2996 4.5005
R22848 DVSS.n5878 DVSS.n2995 4.5005
R22849 DVSS.n2998 DVSS.n2995 4.5005
R22850 DVSS.n2998 DVSS.n2996 4.5005
R22851 DVSS.n2998 DVSS.n2994 4.5005
R22852 DVSS.n5879 DVSS.n2998 4.5005
R22853 DVSS.n5880 DVSS.n2995 4.5005
R22854 DVSS.n5880 DVSS.n2996 4.5005
R22855 DVSS.n5880 DVSS.n2994 4.5005
R22856 DVSS.n5880 DVSS.n5879 4.5005
R22857 DVSS.n2542 DVSS.n2526 4.5005
R22858 DVSS.n7380 DVSS.n2542 4.5005
R22859 DVSS.n7378 DVSS.n2542 4.5005
R22860 DVSS.n7380 DVSS.n2546 4.5005
R22861 DVSS.n7378 DVSS.n2546 4.5005
R22862 DVSS.n7380 DVSS.n2541 4.5005
R22863 DVSS.n7378 DVSS.n2541 4.5005
R22864 DVSS.n7380 DVSS.n2549 4.5005
R22865 DVSS.n7378 DVSS.n2549 4.5005
R22866 DVSS.n7380 DVSS.n2540 4.5005
R22867 DVSS.n7378 DVSS.n2540 4.5005
R22868 DVSS.n7380 DVSS.n2552 4.5005
R22869 DVSS.n7378 DVSS.n2552 4.5005
R22870 DVSS.n7380 DVSS.n2539 4.5005
R22871 DVSS.n7378 DVSS.n2539 4.5005
R22872 DVSS.n7380 DVSS.n2555 4.5005
R22873 DVSS.n7378 DVSS.n2555 4.5005
R22874 DVSS.n7380 DVSS.n2538 4.5005
R22875 DVSS.n7378 DVSS.n2538 4.5005
R22876 DVSS.n7380 DVSS.n2558 4.5005
R22877 DVSS.n7378 DVSS.n2558 4.5005
R22878 DVSS.n7380 DVSS.n2537 4.5005
R22879 DVSS.n7378 DVSS.n2537 4.5005
R22880 DVSS.n7380 DVSS.n2561 4.5005
R22881 DVSS.n7378 DVSS.n2561 4.5005
R22882 DVSS.n7380 DVSS.n2536 4.5005
R22883 DVSS.n7378 DVSS.n2536 4.5005
R22884 DVSS.n7380 DVSS.n2564 4.5005
R22885 DVSS.n7378 DVSS.n2564 4.5005
R22886 DVSS.n7380 DVSS.n2535 4.5005
R22887 DVSS.n7378 DVSS.n2535 4.5005
R22888 DVSS.n7380 DVSS.n2567 4.5005
R22889 DVSS.n7378 DVSS.n2567 4.5005
R22890 DVSS.n7380 DVSS.n2534 4.5005
R22891 DVSS.n7378 DVSS.n2534 4.5005
R22892 DVSS.n7380 DVSS.n2570 4.5005
R22893 DVSS.n7378 DVSS.n2570 4.5005
R22894 DVSS.n7380 DVSS.n2533 4.5005
R22895 DVSS.n7378 DVSS.n2533 4.5005
R22896 DVSS.n7380 DVSS.n2573 4.5005
R22897 DVSS.n7378 DVSS.n2573 4.5005
R22898 DVSS.n7380 DVSS.n2532 4.5005
R22899 DVSS.n7378 DVSS.n2532 4.5005
R22900 DVSS.n7380 DVSS.n2576 4.5005
R22901 DVSS.n7378 DVSS.n2576 4.5005
R22902 DVSS.n7380 DVSS.n2531 4.5005
R22903 DVSS.n7378 DVSS.n2531 4.5005
R22904 DVSS.n7379 DVSS.n2526 4.5005
R22905 DVSS.n7380 DVSS.n7379 4.5005
R22906 DVSS.n7379 DVSS.n7378 4.5005
R22907 DVSS.n8056 DVSS.n1927 4.5005
R22908 DVSS.n1927 DVSS.n1918 4.5005
R22909 DVSS.n8060 DVSS.n1927 4.5005
R22910 DVSS.n1924 DVSS.n1918 4.5005
R22911 DVSS.n8060 DVSS.n1924 4.5005
R22912 DVSS.n1929 DVSS.n1918 4.5005
R22913 DVSS.n8060 DVSS.n1929 4.5005
R22914 DVSS.n1923 DVSS.n1918 4.5005
R22915 DVSS.n8060 DVSS.n1923 4.5005
R22916 DVSS.n1931 DVSS.n1918 4.5005
R22917 DVSS.n8060 DVSS.n1931 4.5005
R22918 DVSS.n1922 DVSS.n1918 4.5005
R22919 DVSS.n8060 DVSS.n1922 4.5005
R22920 DVSS.n1933 DVSS.n1918 4.5005
R22921 DVSS.n8060 DVSS.n1933 4.5005
R22922 DVSS.n1921 DVSS.n1918 4.5005
R22923 DVSS.n8060 DVSS.n1921 4.5005
R22924 DVSS.n8059 DVSS.n1918 4.5005
R22925 DVSS.n8060 DVSS.n8059 4.5005
R22926 DVSS.n1920 DVSS.n1918 4.5005
R22927 DVSS.n8060 DVSS.n1920 4.5005
R22928 DVSS.n8061 DVSS.n1918 4.5005
R22929 DVSS.n8061 DVSS.n1917 4.5005
R22930 DVSS.n8061 DVSS.n8060 4.5005
R22931 DVSS.n6854 DVSS.n6755 4.5005
R22932 DVSS.n6755 DVSS.n6737 4.5005
R22933 DVSS.n6858 DVSS.n6755 4.5005
R22934 DVSS.n6743 DVSS.n6737 4.5005
R22935 DVSS.n6858 DVSS.n6743 4.5005
R22936 DVSS.n6757 DVSS.n6737 4.5005
R22937 DVSS.n6858 DVSS.n6757 4.5005
R22938 DVSS.n6742 DVSS.n6737 4.5005
R22939 DVSS.n6858 DVSS.n6742 4.5005
R22940 DVSS.n6759 DVSS.n6737 4.5005
R22941 DVSS.n6858 DVSS.n6759 4.5005
R22942 DVSS.n6741 DVSS.n6737 4.5005
R22943 DVSS.n6858 DVSS.n6741 4.5005
R22944 DVSS.n6761 DVSS.n6737 4.5005
R22945 DVSS.n6858 DVSS.n6761 4.5005
R22946 DVSS.n6740 DVSS.n6737 4.5005
R22947 DVSS.n6858 DVSS.n6740 4.5005
R22948 DVSS.n6857 DVSS.n6737 4.5005
R22949 DVSS.n6858 DVSS.n6857 4.5005
R22950 DVSS.n6739 DVSS.n6737 4.5005
R22951 DVSS.n6858 DVSS.n6739 4.5005
R22952 DVSS.n6859 DVSS.n6737 4.5005
R22953 DVSS.n6859 DVSS.n6736 4.5005
R22954 DVSS.n6859 DVSS.n6858 4.5005
R22955 DVSS.n4461 DVSS.n4459 4.5005
R22956 DVSS.n4490 DVSS.n4459 4.5005
R22957 DVSS.n4492 DVSS.n4459 4.5005
R22958 DVSS.n4461 DVSS.n3835 4.5005
R22959 DVSS.n4490 DVSS.n3835 4.5005
R22960 DVSS.n4492 DVSS.n3835 4.5005
R22961 DVSS.n4491 DVSS.n4461 4.5005
R22962 DVSS.n4491 DVSS.n4490 4.5005
R22963 DVSS.n4491 DVSS.n3834 4.5005
R22964 DVSS.n4492 DVSS.n4491 4.5005
R22965 DVSS.n4474 DVSS.n4460 4.5005
R22966 DVSS.n6913 DVSS.n6860 4.5005
R22967 DVSS.n6860 DVSS.n6734 4.5005
R22968 DVSS.n6906 DVSS.n6860 4.5005
R22969 DVSS.n6913 DVSS.n6861 4.5005
R22970 DVSS.n6861 DVSS.n6734 4.5005
R22971 DVSS.n6884 DVSS.n6734 4.5005
R22972 DVSS.n6910 DVSS.n6884 4.5005
R22973 DVSS.n6888 DVSS.n6734 4.5005
R22974 DVSS.n6910 DVSS.n6888 4.5005
R22975 DVSS.n6883 DVSS.n6734 4.5005
R22976 DVSS.n6910 DVSS.n6883 4.5005
R22977 DVSS.n6889 DVSS.n6734 4.5005
R22978 DVSS.n6910 DVSS.n6889 4.5005
R22979 DVSS.n6882 DVSS.n6734 4.5005
R22980 DVSS.n6910 DVSS.n6882 4.5005
R22981 DVSS.n6890 DVSS.n6734 4.5005
R22982 DVSS.n6910 DVSS.n6890 4.5005
R22983 DVSS.n6881 DVSS.n6734 4.5005
R22984 DVSS.n6910 DVSS.n6881 4.5005
R22985 DVSS.n6891 DVSS.n6734 4.5005
R22986 DVSS.n6910 DVSS.n6891 4.5005
R22987 DVSS.n6880 DVSS.n6734 4.5005
R22988 DVSS.n6910 DVSS.n6880 4.5005
R22989 DVSS.n6892 DVSS.n6734 4.5005
R22990 DVSS.n6910 DVSS.n6892 4.5005
R22991 DVSS.n6879 DVSS.n6734 4.5005
R22992 DVSS.n6910 DVSS.n6879 4.5005
R22993 DVSS.n6893 DVSS.n6734 4.5005
R22994 DVSS.n6910 DVSS.n6893 4.5005
R22995 DVSS.n6878 DVSS.n6734 4.5005
R22996 DVSS.n6910 DVSS.n6878 4.5005
R22997 DVSS.n6894 DVSS.n6734 4.5005
R22998 DVSS.n6910 DVSS.n6894 4.5005
R22999 DVSS.n6877 DVSS.n6734 4.5005
R23000 DVSS.n6910 DVSS.n6877 4.5005
R23001 DVSS.n6895 DVSS.n6734 4.5005
R23002 DVSS.n6910 DVSS.n6895 4.5005
R23003 DVSS.n6876 DVSS.n6734 4.5005
R23004 DVSS.n6910 DVSS.n6876 4.5005
R23005 DVSS.n6908 DVSS.n6734 4.5005
R23006 DVSS.n6910 DVSS.n6908 4.5005
R23007 DVSS.n6875 DVSS.n6734 4.5005
R23008 DVSS.n6910 DVSS.n6875 4.5005
R23009 DVSS.n6909 DVSS.n6734 4.5005
R23010 DVSS.n6910 DVSS.n6909 4.5005
R23011 DVSS.n6911 DVSS.n6734 4.5005
R23012 DVSS.n6911 DVSS.n6910 4.5005
R23013 DVSS.n6872 DVSS.n6734 4.5005
R23014 DVSS.n6906 DVSS.n6872 4.5005
R23015 DVSS.n6910 DVSS.n6872 4.5005
R23016 DVSS.n7060 DVSS.n6691 4.5005
R23017 DVSS.n7060 DVSS.n6692 4.5005
R23018 DVSS.n7060 DVSS.n7059 4.5005
R23019 DVSS.n6706 DVSS.n6692 4.5005
R23020 DVSS.n7059 DVSS.n6706 4.5005
R23021 DVSS.n6703 DVSS.n6692 4.5005
R23022 DVSS.n7059 DVSS.n6703 4.5005
R23023 DVSS.n6708 DVSS.n6692 4.5005
R23024 DVSS.n7059 DVSS.n6708 4.5005
R23025 DVSS.n6702 DVSS.n6692 4.5005
R23026 DVSS.n7059 DVSS.n6702 4.5005
R23027 DVSS.n6710 DVSS.n6692 4.5005
R23028 DVSS.n7059 DVSS.n6710 4.5005
R23029 DVSS.n6701 DVSS.n6692 4.5005
R23030 DVSS.n7059 DVSS.n6701 4.5005
R23031 DVSS.n6712 DVSS.n6692 4.5005
R23032 DVSS.n7059 DVSS.n6712 4.5005
R23033 DVSS.n6700 DVSS.n6692 4.5005
R23034 DVSS.n7059 DVSS.n6700 4.5005
R23035 DVSS.n6714 DVSS.n6692 4.5005
R23036 DVSS.n7059 DVSS.n6714 4.5005
R23037 DVSS.n6699 DVSS.n6692 4.5005
R23038 DVSS.n7059 DVSS.n6699 4.5005
R23039 DVSS.n6716 DVSS.n6692 4.5005
R23040 DVSS.n7059 DVSS.n6716 4.5005
R23041 DVSS.n6698 DVSS.n6692 4.5005
R23042 DVSS.n7059 DVSS.n6698 4.5005
R23043 DVSS.n6718 DVSS.n6692 4.5005
R23044 DVSS.n7059 DVSS.n6718 4.5005
R23045 DVSS.n6697 DVSS.n6692 4.5005
R23046 DVSS.n7059 DVSS.n6697 4.5005
R23047 DVSS.n6720 DVSS.n6692 4.5005
R23048 DVSS.n7059 DVSS.n6720 4.5005
R23049 DVSS.n6696 DVSS.n6692 4.5005
R23050 DVSS.n7059 DVSS.n6696 4.5005
R23051 DVSS.n6722 DVSS.n6692 4.5005
R23052 DVSS.n7059 DVSS.n6722 4.5005
R23053 DVSS.n6695 DVSS.n6692 4.5005
R23054 DVSS.n7059 DVSS.n6695 4.5005
R23055 DVSS.n6724 DVSS.n6692 4.5005
R23056 DVSS.n7059 DVSS.n6724 4.5005
R23057 DVSS.n6694 DVSS.n6692 4.5005
R23058 DVSS.n7059 DVSS.n6694 4.5005
R23059 DVSS.n7058 DVSS.n6692 4.5005
R23060 DVSS.n7059 DVSS.n7058 4.5005
R23061 DVSS.n6692 DVSS.n784 4.5005
R23062 DVSS.n7055 DVSS.n784 4.5005
R23063 DVSS.n7059 DVSS.n784 4.5005
R23064 DVSS.n7055 DVSS.n785 4.5005
R23065 DVSS.n7059 DVSS.n785 4.5005
R23066 DVSS.n6692 DVSS.n785 4.5005
R23067 DVSS.n6691 DVSS.n785 4.5005
R23068 DVSS.n1316 DVSS.n1190 4.5005
R23069 DVSS.n1316 DVSS.n1191 4.5005
R23070 DVSS.n1316 DVSS.n1315 4.5005
R23071 DVSS.n1203 DVSS.n1190 4.5005
R23072 DVSS.n1203 DVSS.n1191 4.5005
R23073 DVSS.n1315 DVSS.n1203 4.5005
R23074 DVSS.n1315 DVSS.n1201 4.5005
R23075 DVSS.n1311 DVSS.n1201 4.5005
R23076 DVSS.n1201 DVSS.n1191 4.5005
R23077 DVSS.n1201 DVSS.n1190 4.5005
R23078 DVSS.n1315 DVSS.n1205 4.5005
R23079 DVSS.n1311 DVSS.n1205 4.5005
R23080 DVSS.n1205 DVSS.n1190 4.5005
R23081 DVSS.n1200 DVSS.n1190 4.5005
R23082 DVSS.n1315 DVSS.n1200 4.5005
R23083 DVSS.n1207 DVSS.n1191 4.5005
R23084 DVSS.n1315 DVSS.n1207 4.5005
R23085 DVSS.n1199 DVSS.n1191 4.5005
R23086 DVSS.n1315 DVSS.n1199 4.5005
R23087 DVSS.n1209 DVSS.n1191 4.5005
R23088 DVSS.n1315 DVSS.n1209 4.5005
R23089 DVSS.n1198 DVSS.n1191 4.5005
R23090 DVSS.n1315 DVSS.n1198 4.5005
R23091 DVSS.n1211 DVSS.n1191 4.5005
R23092 DVSS.n1315 DVSS.n1211 4.5005
R23093 DVSS.n1197 DVSS.n1191 4.5005
R23094 DVSS.n1315 DVSS.n1197 4.5005
R23095 DVSS.n1213 DVSS.n1191 4.5005
R23096 DVSS.n1315 DVSS.n1213 4.5005
R23097 DVSS.n1196 DVSS.n1191 4.5005
R23098 DVSS.n1311 DVSS.n1196 4.5005
R23099 DVSS.n1315 DVSS.n1196 4.5005
R23100 DVSS.n1297 DVSS.n1190 4.5005
R23101 DVSS.n1297 DVSS.n1191 4.5005
R23102 DVSS.n1311 DVSS.n1297 4.5005
R23103 DVSS.n1315 DVSS.n1297 4.5005
R23104 DVSS.n1195 DVSS.n1190 4.5005
R23105 DVSS.n1195 DVSS.n1191 4.5005
R23106 DVSS.n1315 DVSS.n1195 4.5005
R23107 DVSS.n1299 DVSS.n1191 4.5005
R23108 DVSS.n1315 DVSS.n1299 4.5005
R23109 DVSS.n1194 DVSS.n1191 4.5005
R23110 DVSS.n1315 DVSS.n1194 4.5005
R23111 DVSS.n1301 DVSS.n1191 4.5005
R23112 DVSS.n1315 DVSS.n1301 4.5005
R23113 DVSS.n1193 DVSS.n1191 4.5005
R23114 DVSS.n1315 DVSS.n1193 4.5005
R23115 DVSS.n1303 DVSS.n1191 4.5005
R23116 DVSS.n1315 DVSS.n1303 4.5005
R23117 DVSS.n1192 DVSS.n1191 4.5005
R23118 DVSS.n1315 DVSS.n1192 4.5005
R23119 DVSS.n1314 DVSS.n1191 4.5005
R23120 DVSS.n1315 DVSS.n1314 4.5005
R23121 DVSS.n1191 DVSS.n789 4.5005
R23122 DVSS.n1311 DVSS.n789 4.5005
R23123 DVSS.n1315 DVSS.n789 4.5005
R23124 DVSS.n1315 DVSS.n791 4.5005
R23125 DVSS.n1311 DVSS.n791 4.5005
R23126 DVSS.n1191 DVSS.n791 4.5005
R23127 DVSS.n1190 DVSS.n791 4.5005
R23128 DVSS.n8561 DVSS.n1073 4.5005
R23129 DVSS.n8534 DVSS.n1073 4.5005
R23130 DVSS.n8559 DVSS.n1073 4.5005
R23131 DVSS.n8561 DVSS.n1074 4.5005
R23132 DVSS.n8534 DVSS.n1074 4.5005
R23133 DVSS.n8559 DVSS.n1074 4.5005
R23134 DVSS.n8559 DVSS.n1072 4.5005
R23135 DVSS.n1078 DVSS.n1072 4.5005
R23136 DVSS.n8534 DVSS.n1072 4.5005
R23137 DVSS.n8561 DVSS.n1072 4.5005
R23138 DVSS.n8559 DVSS.n1075 4.5005
R23139 DVSS.n1078 DVSS.n1075 4.5005
R23140 DVSS.n8561 DVSS.n1075 4.5005
R23141 DVSS.n8561 DVSS.n1071 4.5005
R23142 DVSS.n8559 DVSS.n1071 4.5005
R23143 DVSS.n8544 DVSS.n8534 4.5005
R23144 DVSS.n8559 DVSS.n8544 4.5005
R23145 DVSS.n8541 DVSS.n8534 4.5005
R23146 DVSS.n8559 DVSS.n8541 4.5005
R23147 DVSS.n8546 DVSS.n8534 4.5005
R23148 DVSS.n8559 DVSS.n8546 4.5005
R23149 DVSS.n8540 DVSS.n8534 4.5005
R23150 DVSS.n8559 DVSS.n8540 4.5005
R23151 DVSS.n8548 DVSS.n8534 4.5005
R23152 DVSS.n8559 DVSS.n8548 4.5005
R23153 DVSS.n8539 DVSS.n8534 4.5005
R23154 DVSS.n8559 DVSS.n8539 4.5005
R23155 DVSS.n8550 DVSS.n8534 4.5005
R23156 DVSS.n8559 DVSS.n8550 4.5005
R23157 DVSS.n8538 DVSS.n8534 4.5005
R23158 DVSS.n8538 DVSS.n1078 4.5005
R23159 DVSS.n8559 DVSS.n8538 4.5005
R23160 DVSS.n8561 DVSS.n8560 4.5005
R23161 DVSS.n8560 DVSS.n8534 4.5005
R23162 DVSS.n8560 DVSS.n1078 4.5005
R23163 DVSS.n8560 DVSS.n8559 4.5005
R23164 DVSS.n8561 DVSS.n1066 4.5005
R23165 DVSS.n8534 DVSS.n1066 4.5005
R23166 DVSS.n8559 DVSS.n1066 4.5005
R23167 DVSS.n8552 DVSS.n8534 4.5005
R23168 DVSS.n8559 DVSS.n8552 4.5005
R23169 DVSS.n8537 DVSS.n8534 4.5005
R23170 DVSS.n8559 DVSS.n8537 4.5005
R23171 DVSS.n8554 DVSS.n8534 4.5005
R23172 DVSS.n8559 DVSS.n8554 4.5005
R23173 DVSS.n8536 DVSS.n8534 4.5005
R23174 DVSS.n8559 DVSS.n8536 4.5005
R23175 DVSS.n8556 DVSS.n8534 4.5005
R23176 DVSS.n8559 DVSS.n8556 4.5005
R23177 DVSS.n8535 DVSS.n8534 4.5005
R23178 DVSS.n8559 DVSS.n8535 4.5005
R23179 DVSS.n8558 DVSS.n8534 4.5005
R23180 DVSS.n8559 DVSS.n8558 4.5005
R23181 DVSS.n8534 DVSS.n799 4.5005
R23182 DVSS.n1078 DVSS.n799 4.5005
R23183 DVSS.n8559 DVSS.n799 4.5005
R23184 DVSS.n8559 DVSS.n801 4.5005
R23185 DVSS.n1078 DVSS.n801 4.5005
R23186 DVSS.n8534 DVSS.n801 4.5005
R23187 DVSS.n8561 DVSS.n801 4.5005
R23188 DVSS.n9130 DVSS.n595 4.5005
R23189 DVSS.n9128 DVSS.n595 4.5005
R23190 DVSS.n9130 DVSS.n596 4.5005
R23191 DVSS.n9128 DVSS.n596 4.5005
R23192 DVSS.n9128 DVSS.n594 4.5005
R23193 DVSS.n605 DVSS.n594 4.5005
R23194 DVSS.n9130 DVSS.n594 4.5005
R23195 DVSS.n9128 DVSS.n597 4.5005
R23196 DVSS.n9130 DVSS.n597 4.5005
R23197 DVSS.n9128 DVSS.n616 4.5005
R23198 DVSS.n9128 DVSS.n9113 4.5005
R23199 DVSS.n9128 DVSS.n614 4.5005
R23200 DVSS.n9128 DVSS.n9115 4.5005
R23201 DVSS.n9128 DVSS.n613 4.5005
R23202 DVSS.n9128 DVSS.n9117 4.5005
R23203 DVSS.n9128 DVSS.n612 4.5005
R23204 DVSS.n9128 DVSS.n9119 4.5005
R23205 DVSS.n9130 DVSS.n589 4.5005
R23206 DVSS.n9128 DVSS.n589 4.5005
R23207 DVSS.n9130 DVSS.n598 4.5005
R23208 DVSS.n605 DVSS.n598 4.5005
R23209 DVSS.n9128 DVSS.n598 4.5005
R23210 DVSS.n9130 DVSS.n588 4.5005
R23211 DVSS.n9128 DVSS.n588 4.5005
R23212 DVSS.n9128 DVSS.n9121 4.5005
R23213 DVSS.n9128 DVSS.n611 4.5005
R23214 DVSS.n9128 DVSS.n9123 4.5005
R23215 DVSS.n9128 DVSS.n610 4.5005
R23216 DVSS.n9128 DVSS.n9125 4.5005
R23217 DVSS.n9128 DVSS.n609 4.5005
R23218 DVSS.n9128 DVSS.n9127 4.5005
R23219 DVSS.n608 DVSS.n605 4.5005
R23220 DVSS.n9128 DVSS.n608 4.5005
R23221 DVSS.n9129 DVSS.n9128 4.5005
R23222 DVSS.n9129 DVSS.n605 4.5005
R23223 DVSS.n9130 DVSS.n9129 4.5005
R23224 DVSS.n9159 DVSS.n567 4.5005
R23225 DVSS.n9156 DVSS.n567 4.5005
R23226 DVSS.n9159 DVSS.n568 4.5005
R23227 DVSS.n9156 DVSS.n568 4.5005
R23228 DVSS.n9156 DVSS.n566 4.5005
R23229 DVSS.n9153 DVSS.n566 4.5005
R23230 DVSS.n9159 DVSS.n566 4.5005
R23231 DVSS.n9156 DVSS.n569 4.5005
R23232 DVSS.n9159 DVSS.n569 4.5005
R23233 DVSS.n9156 DVSS.n582 4.5005
R23234 DVSS.n9156 DVSS.n9139 4.5005
R23235 DVSS.n9156 DVSS.n581 4.5005
R23236 DVSS.n9156 DVSS.n9140 4.5005
R23237 DVSS.n9156 DVSS.n580 4.5005
R23238 DVSS.n9156 DVSS.n9141 4.5005
R23239 DVSS.n9156 DVSS.n579 4.5005
R23240 DVSS.n9156 DVSS.n9142 4.5005
R23241 DVSS.n9159 DVSS.n561 4.5005
R23242 DVSS.n9156 DVSS.n561 4.5005
R23243 DVSS.n9159 DVSS.n570 4.5005
R23244 DVSS.n9153 DVSS.n570 4.5005
R23245 DVSS.n9156 DVSS.n570 4.5005
R23246 DVSS.n9159 DVSS.n560 4.5005
R23247 DVSS.n9156 DVSS.n560 4.5005
R23248 DVSS.n9156 DVSS.n9143 4.5005
R23249 DVSS.n9156 DVSS.n578 4.5005
R23250 DVSS.n9156 DVSS.n9144 4.5005
R23251 DVSS.n9156 DVSS.n577 4.5005
R23252 DVSS.n9156 DVSS.n9155 4.5005
R23253 DVSS.n9156 DVSS.n576 4.5005
R23254 DVSS.n9157 DVSS.n9156 4.5005
R23255 DVSS.n9153 DVSS.n374 4.5005
R23256 DVSS.n9156 DVSS.n374 4.5005
R23257 DVSS.n9156 DVSS.n375 4.5005
R23258 DVSS.n9153 DVSS.n375 4.5005
R23259 DVSS.n9159 DVSS.n375 4.5005
R23260 DVSS.n9660 DVSS.n216 4.5005
R23261 DVSS.n222 DVSS.n216 4.5005
R23262 DVSS.n223 DVSS.n216 4.5005
R23263 DVSS.n9660 DVSS.n217 4.5005
R23264 DVSS.n222 DVSS.n217 4.5005
R23265 DVSS.n223 DVSS.n217 4.5005
R23266 DVSS.n223 DVSS.n215 4.5005
R23267 DVSS.n9658 DVSS.n215 4.5005
R23268 DVSS.n222 DVSS.n215 4.5005
R23269 DVSS.n9660 DVSS.n215 4.5005
R23270 DVSS.n223 DVSS.n218 4.5005
R23271 DVSS.n9658 DVSS.n218 4.5005
R23272 DVSS.n9660 DVSS.n218 4.5005
R23273 DVSS.n9660 DVSS.n214 4.5005
R23274 DVSS.n223 DVSS.n214 4.5005
R23275 DVSS.n9636 DVSS.n222 4.5005
R23276 DVSS.n9636 DVSS.n223 4.5005
R23277 DVSS.n9639 DVSS.n222 4.5005
R23278 DVSS.n9639 DVSS.n223 4.5005
R23279 DVSS.n9638 DVSS.n222 4.5005
R23280 DVSS.n9638 DVSS.n223 4.5005
R23281 DVSS.n9642 DVSS.n222 4.5005
R23282 DVSS.n9642 DVSS.n223 4.5005
R23283 DVSS.n9641 DVSS.n222 4.5005
R23284 DVSS.n9641 DVSS.n223 4.5005
R23285 DVSS.n9645 DVSS.n222 4.5005
R23286 DVSS.n9645 DVSS.n223 4.5005
R23287 DVSS.n9644 DVSS.n222 4.5005
R23288 DVSS.n9644 DVSS.n223 4.5005
R23289 DVSS.n227 DVSS.n222 4.5005
R23290 DVSS.n9658 DVSS.n227 4.5005
R23291 DVSS.n227 DVSS.n223 4.5005
R23292 DVSS.n9660 DVSS.n219 4.5005
R23293 DVSS.n222 DVSS.n219 4.5005
R23294 DVSS.n9658 DVSS.n219 4.5005
R23295 DVSS.n223 DVSS.n219 4.5005
R23296 DVSS.n9660 DVSS.n209 4.5005
R23297 DVSS.n222 DVSS.n209 4.5005
R23298 DVSS.n223 DVSS.n209 4.5005
R23299 DVSS.n9647 DVSS.n222 4.5005
R23300 DVSS.n9647 DVSS.n223 4.5005
R23301 DVSS.n9650 DVSS.n222 4.5005
R23302 DVSS.n9650 DVSS.n223 4.5005
R23303 DVSS.n9649 DVSS.n222 4.5005
R23304 DVSS.n9649 DVSS.n223 4.5005
R23305 DVSS.n9653 DVSS.n222 4.5005
R23306 DVSS.n9653 DVSS.n223 4.5005
R23307 DVSS.n9652 DVSS.n222 4.5005
R23308 DVSS.n9652 DVSS.n223 4.5005
R23309 DVSS.n9656 DVSS.n222 4.5005
R23310 DVSS.n9656 DVSS.n223 4.5005
R23311 DVSS.n9655 DVSS.n222 4.5005
R23312 DVSS.n9655 DVSS.n223 4.5005
R23313 DVSS.n226 DVSS.n222 4.5005
R23314 DVSS.n9658 DVSS.n226 4.5005
R23315 DVSS.n226 DVSS.n223 4.5005
R23316 DVSS.n9659 DVSS.n223 4.5005
R23317 DVSS.n9659 DVSS.n9658 4.5005
R23318 DVSS.n9659 DVSS.n222 4.5005
R23319 DVSS.n9660 DVSS.n9659 4.5005
R23320 DVSS.n9717 DVSS.n177 4.5005
R23321 DVSS.n183 DVSS.n177 4.5005
R23322 DVSS.n184 DVSS.n177 4.5005
R23323 DVSS.n9717 DVSS.n178 4.5005
R23324 DVSS.n183 DVSS.n178 4.5005
R23325 DVSS.n184 DVSS.n178 4.5005
R23326 DVSS.n184 DVSS.n176 4.5005
R23327 DVSS.n9715 DVSS.n176 4.5005
R23328 DVSS.n183 DVSS.n176 4.5005
R23329 DVSS.n9717 DVSS.n176 4.5005
R23330 DVSS.n184 DVSS.n179 4.5005
R23331 DVSS.n9715 DVSS.n179 4.5005
R23332 DVSS.n9717 DVSS.n179 4.5005
R23333 DVSS.n9717 DVSS.n175 4.5005
R23334 DVSS.n184 DVSS.n175 4.5005
R23335 DVSS.n9693 DVSS.n183 4.5005
R23336 DVSS.n9693 DVSS.n184 4.5005
R23337 DVSS.n9696 DVSS.n183 4.5005
R23338 DVSS.n9696 DVSS.n184 4.5005
R23339 DVSS.n9695 DVSS.n183 4.5005
R23340 DVSS.n9695 DVSS.n184 4.5005
R23341 DVSS.n9699 DVSS.n183 4.5005
R23342 DVSS.n9699 DVSS.n184 4.5005
R23343 DVSS.n9698 DVSS.n183 4.5005
R23344 DVSS.n9698 DVSS.n184 4.5005
R23345 DVSS.n9702 DVSS.n183 4.5005
R23346 DVSS.n9702 DVSS.n184 4.5005
R23347 DVSS.n9701 DVSS.n183 4.5005
R23348 DVSS.n9701 DVSS.n184 4.5005
R23349 DVSS.n188 DVSS.n183 4.5005
R23350 DVSS.n9715 DVSS.n188 4.5005
R23351 DVSS.n188 DVSS.n184 4.5005
R23352 DVSS.n9717 DVSS.n180 4.5005
R23353 DVSS.n183 DVSS.n180 4.5005
R23354 DVSS.n9715 DVSS.n180 4.5005
R23355 DVSS.n184 DVSS.n180 4.5005
R23356 DVSS.n9717 DVSS.n170 4.5005
R23357 DVSS.n183 DVSS.n170 4.5005
R23358 DVSS.n184 DVSS.n170 4.5005
R23359 DVSS.n9704 DVSS.n183 4.5005
R23360 DVSS.n9704 DVSS.n184 4.5005
R23361 DVSS.n9707 DVSS.n183 4.5005
R23362 DVSS.n9707 DVSS.n184 4.5005
R23363 DVSS.n9706 DVSS.n183 4.5005
R23364 DVSS.n9706 DVSS.n184 4.5005
R23365 DVSS.n9710 DVSS.n183 4.5005
R23366 DVSS.n9710 DVSS.n184 4.5005
R23367 DVSS.n9709 DVSS.n183 4.5005
R23368 DVSS.n9709 DVSS.n184 4.5005
R23369 DVSS.n9713 DVSS.n183 4.5005
R23370 DVSS.n9713 DVSS.n184 4.5005
R23371 DVSS.n9712 DVSS.n183 4.5005
R23372 DVSS.n9712 DVSS.n184 4.5005
R23373 DVSS.n187 DVSS.n183 4.5005
R23374 DVSS.n9715 DVSS.n187 4.5005
R23375 DVSS.n187 DVSS.n184 4.5005
R23376 DVSS.n9716 DVSS.n184 4.5005
R23377 DVSS.n9716 DVSS.n9715 4.5005
R23378 DVSS.n9716 DVSS.n183 4.5005
R23379 DVSS.n9717 DVSS.n9716 4.5005
R23380 DVSS.n9770 DVSS.n155 4.5005
R23381 DVSS.n155 DVSS.n143 4.5005
R23382 DVSS.n157 DVSS.n155 4.5005
R23383 DVSS.n9736 DVSS.n143 4.5005
R23384 DVSS.n9736 DVSS.n157 4.5005
R23385 DVSS.n9739 DVSS.n143 4.5005
R23386 DVSS.n9739 DVSS.n157 4.5005
R23387 DVSS.n9738 DVSS.n143 4.5005
R23388 DVSS.n9738 DVSS.n157 4.5005
R23389 DVSS.n9742 DVSS.n143 4.5005
R23390 DVSS.n9742 DVSS.n157 4.5005
R23391 DVSS.n9741 DVSS.n143 4.5005
R23392 DVSS.n9741 DVSS.n157 4.5005
R23393 DVSS.n9745 DVSS.n143 4.5005
R23394 DVSS.n9745 DVSS.n157 4.5005
R23395 DVSS.n9744 DVSS.n143 4.5005
R23396 DVSS.n9744 DVSS.n157 4.5005
R23397 DVSS.n9748 DVSS.n143 4.5005
R23398 DVSS.n9748 DVSS.n157 4.5005
R23399 DVSS.n9747 DVSS.n143 4.5005
R23400 DVSS.n9747 DVSS.n157 4.5005
R23401 DVSS.n9751 DVSS.n143 4.5005
R23402 DVSS.n9751 DVSS.n157 4.5005
R23403 DVSS.n9750 DVSS.n143 4.5005
R23404 DVSS.n9750 DVSS.n157 4.5005
R23405 DVSS.n9754 DVSS.n143 4.5005
R23406 DVSS.n9754 DVSS.n157 4.5005
R23407 DVSS.n9753 DVSS.n143 4.5005
R23408 DVSS.n9753 DVSS.n157 4.5005
R23409 DVSS.n9757 DVSS.n143 4.5005
R23410 DVSS.n9757 DVSS.n157 4.5005
R23411 DVSS.n9756 DVSS.n143 4.5005
R23412 DVSS.n9756 DVSS.n157 4.5005
R23413 DVSS.n9760 DVSS.n143 4.5005
R23414 DVSS.n9760 DVSS.n157 4.5005
R23415 DVSS.n9759 DVSS.n143 4.5005
R23416 DVSS.n9759 DVSS.n157 4.5005
R23417 DVSS.n9763 DVSS.n143 4.5005
R23418 DVSS.n9763 DVSS.n157 4.5005
R23419 DVSS.n9762 DVSS.n143 4.5005
R23420 DVSS.n9762 DVSS.n157 4.5005
R23421 DVSS.n9766 DVSS.n143 4.5005
R23422 DVSS.n9766 DVSS.n157 4.5005
R23423 DVSS.n9765 DVSS.n143 4.5005
R23424 DVSS.n9765 DVSS.n157 4.5005
R23425 DVSS.n9734 DVSS.n143 4.5005
R23426 DVSS.n9768 DVSS.n9734 4.5005
R23427 DVSS.n9734 DVSS.n157 4.5005
R23428 DVSS.n9769 DVSS.n157 4.5005
R23429 DVSS.n9769 DVSS.n9768 4.5005
R23430 DVSS.n9769 DVSS.n143 4.5005
R23431 DVSS.n9770 DVSS.n9769 4.5005
R23432 DVSS.n112 DVSS.n98 4.5005
R23433 DVSS.n112 DVSS.n99 4.5005
R23434 DVSS.n9803 DVSS.n112 4.5005
R23435 DVSS.n115 DVSS.n99 4.5005
R23436 DVSS.n9803 DVSS.n115 4.5005
R23437 DVSS.n111 DVSS.n99 4.5005
R23438 DVSS.n9803 DVSS.n111 4.5005
R23439 DVSS.n117 DVSS.n99 4.5005
R23440 DVSS.n9803 DVSS.n117 4.5005
R23441 DVSS.n110 DVSS.n99 4.5005
R23442 DVSS.n9803 DVSS.n110 4.5005
R23443 DVSS.n119 DVSS.n99 4.5005
R23444 DVSS.n9803 DVSS.n119 4.5005
R23445 DVSS.n109 DVSS.n99 4.5005
R23446 DVSS.n9803 DVSS.n109 4.5005
R23447 DVSS.n121 DVSS.n99 4.5005
R23448 DVSS.n9803 DVSS.n121 4.5005
R23449 DVSS.n108 DVSS.n99 4.5005
R23450 DVSS.n9803 DVSS.n108 4.5005
R23451 DVSS.n123 DVSS.n99 4.5005
R23452 DVSS.n9803 DVSS.n123 4.5005
R23453 DVSS.n107 DVSS.n99 4.5005
R23454 DVSS.n9803 DVSS.n107 4.5005
R23455 DVSS.n125 DVSS.n99 4.5005
R23456 DVSS.n9803 DVSS.n125 4.5005
R23457 DVSS.n106 DVSS.n99 4.5005
R23458 DVSS.n9803 DVSS.n106 4.5005
R23459 DVSS.n127 DVSS.n99 4.5005
R23460 DVSS.n9803 DVSS.n127 4.5005
R23461 DVSS.n105 DVSS.n99 4.5005
R23462 DVSS.n9803 DVSS.n105 4.5005
R23463 DVSS.n129 DVSS.n99 4.5005
R23464 DVSS.n9803 DVSS.n129 4.5005
R23465 DVSS.n104 DVSS.n99 4.5005
R23466 DVSS.n9803 DVSS.n104 4.5005
R23467 DVSS.n131 DVSS.n99 4.5005
R23468 DVSS.n9803 DVSS.n131 4.5005
R23469 DVSS.n103 DVSS.n99 4.5005
R23470 DVSS.n9803 DVSS.n103 4.5005
R23471 DVSS.n133 DVSS.n99 4.5005
R23472 DVSS.n9803 DVSS.n133 4.5005
R23473 DVSS.n102 DVSS.n99 4.5005
R23474 DVSS.n9803 DVSS.n102 4.5005
R23475 DVSS.n9802 DVSS.n99 4.5005
R23476 DVSS.n9803 DVSS.n9802 4.5005
R23477 DVSS.n101 DVSS.n99 4.5005
R23478 DVSS.n9803 DVSS.n101 4.5005
R23479 DVSS.n9804 DVSS.n98 4.5005
R23480 DVSS.n9804 DVSS.n99 4.5005
R23481 DVSS.n9804 DVSS.n9803 4.5005
R23482 DVSS.n991 DVSS.n977 4.5005
R23483 DVSS.n991 DVSS.n978 4.5005
R23484 DVSS.n8638 DVSS.n991 4.5005
R23485 DVSS.n994 DVSS.n978 4.5005
R23486 DVSS.n8638 DVSS.n994 4.5005
R23487 DVSS.n990 DVSS.n978 4.5005
R23488 DVSS.n8638 DVSS.n990 4.5005
R23489 DVSS.n996 DVSS.n978 4.5005
R23490 DVSS.n8638 DVSS.n996 4.5005
R23491 DVSS.n989 DVSS.n978 4.5005
R23492 DVSS.n8638 DVSS.n989 4.5005
R23493 DVSS.n998 DVSS.n978 4.5005
R23494 DVSS.n8638 DVSS.n998 4.5005
R23495 DVSS.n988 DVSS.n978 4.5005
R23496 DVSS.n8638 DVSS.n988 4.5005
R23497 DVSS.n1000 DVSS.n978 4.5005
R23498 DVSS.n8638 DVSS.n1000 4.5005
R23499 DVSS.n987 DVSS.n978 4.5005
R23500 DVSS.n8638 DVSS.n987 4.5005
R23501 DVSS.n1002 DVSS.n978 4.5005
R23502 DVSS.n8638 DVSS.n1002 4.5005
R23503 DVSS.n986 DVSS.n978 4.5005
R23504 DVSS.n8638 DVSS.n986 4.5005
R23505 DVSS.n1004 DVSS.n978 4.5005
R23506 DVSS.n8638 DVSS.n1004 4.5005
R23507 DVSS.n985 DVSS.n978 4.5005
R23508 DVSS.n8638 DVSS.n985 4.5005
R23509 DVSS.n1006 DVSS.n978 4.5005
R23510 DVSS.n8638 DVSS.n1006 4.5005
R23511 DVSS.n984 DVSS.n978 4.5005
R23512 DVSS.n8638 DVSS.n984 4.5005
R23513 DVSS.n1008 DVSS.n978 4.5005
R23514 DVSS.n8638 DVSS.n1008 4.5005
R23515 DVSS.n983 DVSS.n978 4.5005
R23516 DVSS.n8638 DVSS.n983 4.5005
R23517 DVSS.n1010 DVSS.n978 4.5005
R23518 DVSS.n8638 DVSS.n1010 4.5005
R23519 DVSS.n982 DVSS.n978 4.5005
R23520 DVSS.n8638 DVSS.n982 4.5005
R23521 DVSS.n1012 DVSS.n978 4.5005
R23522 DVSS.n8638 DVSS.n1012 4.5005
R23523 DVSS.n981 DVSS.n978 4.5005
R23524 DVSS.n8638 DVSS.n981 4.5005
R23525 DVSS.n8637 DVSS.n978 4.5005
R23526 DVSS.n8638 DVSS.n8637 4.5005
R23527 DVSS.n980 DVSS.n978 4.5005
R23528 DVSS.n8638 DVSS.n980 4.5005
R23529 DVSS.n8639 DVSS.n977 4.5005
R23530 DVSS.n8639 DVSS.n978 4.5005
R23531 DVSS.n8639 DVSS.n8638 4.5005
R23532 DVSS.n769 DVSS.n755 4.5005
R23533 DVSS.n8937 DVSS.n769 4.5005
R23534 DVSS.n769 DVSS.n757 4.5005
R23535 DVSS.n769 DVSS.n756 4.5005
R23536 DVSS.n771 DVSS.n756 4.5005
R23537 DVSS.n771 DVSS.n757 4.5005
R23538 DVSS.n771 DVSS.n755 4.5005
R23539 DVSS.n8937 DVSS.n771 4.5005
R23540 DVSS.n768 DVSS.n756 4.5005
R23541 DVSS.n768 DVSS.n757 4.5005
R23542 DVSS.n768 DVSS.n755 4.5005
R23543 DVSS.n8937 DVSS.n768 4.5005
R23544 DVSS.n772 DVSS.n756 4.5005
R23545 DVSS.n772 DVSS.n757 4.5005
R23546 DVSS.n772 DVSS.n755 4.5005
R23547 DVSS.n8937 DVSS.n772 4.5005
R23548 DVSS.n767 DVSS.n756 4.5005
R23549 DVSS.n767 DVSS.n757 4.5005
R23550 DVSS.n767 DVSS.n755 4.5005
R23551 DVSS.n8937 DVSS.n767 4.5005
R23552 DVSS.n773 DVSS.n755 4.5005
R23553 DVSS.n8937 DVSS.n773 4.5005
R23554 DVSS.n773 DVSS.n757 4.5005
R23555 DVSS.n773 DVSS.n756 4.5005
R23556 DVSS.n766 DVSS.n755 4.5005
R23557 DVSS.n8937 DVSS.n766 4.5005
R23558 DVSS.n766 DVSS.n757 4.5005
R23559 DVSS.n766 DVSS.n756 4.5005
R23560 DVSS.n774 DVSS.n755 4.5005
R23561 DVSS.n8937 DVSS.n774 4.5005
R23562 DVSS.n774 DVSS.n757 4.5005
R23563 DVSS.n774 DVSS.n756 4.5005
R23564 DVSS.n765 DVSS.n756 4.5005
R23565 DVSS.n765 DVSS.n757 4.5005
R23566 DVSS.n765 DVSS.n755 4.5005
R23567 DVSS.n8937 DVSS.n765 4.5005
R23568 DVSS.n775 DVSS.n756 4.5005
R23569 DVSS.n775 DVSS.n757 4.5005
R23570 DVSS.n775 DVSS.n755 4.5005
R23571 DVSS.n8937 DVSS.n775 4.5005
R23572 DVSS.n764 DVSS.n756 4.5005
R23573 DVSS.n764 DVSS.n757 4.5005
R23574 DVSS.n764 DVSS.n755 4.5005
R23575 DVSS.n8937 DVSS.n764 4.5005
R23576 DVSS.n776 DVSS.n756 4.5005
R23577 DVSS.n776 DVSS.n757 4.5005
R23578 DVSS.n776 DVSS.n755 4.5005
R23579 DVSS.n8937 DVSS.n776 4.5005
R23580 DVSS.n763 DVSS.n755 4.5005
R23581 DVSS.n8937 DVSS.n763 4.5005
R23582 DVSS.n763 DVSS.n757 4.5005
R23583 DVSS.n763 DVSS.n756 4.5005
R23584 DVSS.n777 DVSS.n755 4.5005
R23585 DVSS.n8937 DVSS.n777 4.5005
R23586 DVSS.n777 DVSS.n757 4.5005
R23587 DVSS.n777 DVSS.n756 4.5005
R23588 DVSS.n762 DVSS.n755 4.5005
R23589 DVSS.n8937 DVSS.n762 4.5005
R23590 DVSS.n762 DVSS.n757 4.5005
R23591 DVSS.n762 DVSS.n756 4.5005
R23592 DVSS.n778 DVSS.n756 4.5005
R23593 DVSS.n778 DVSS.n757 4.5005
R23594 DVSS.n778 DVSS.n755 4.5005
R23595 DVSS.n8937 DVSS.n778 4.5005
R23596 DVSS.n761 DVSS.n756 4.5005
R23597 DVSS.n761 DVSS.n757 4.5005
R23598 DVSS.n761 DVSS.n755 4.5005
R23599 DVSS.n8937 DVSS.n761 4.5005
R23600 DVSS.n779 DVSS.n756 4.5005
R23601 DVSS.n779 DVSS.n757 4.5005
R23602 DVSS.n779 DVSS.n755 4.5005
R23603 DVSS.n8937 DVSS.n779 4.5005
R23604 DVSS.n760 DVSS.n755 4.5005
R23605 DVSS.n8937 DVSS.n760 4.5005
R23606 DVSS.n760 DVSS.n757 4.5005
R23607 DVSS.n760 DVSS.n756 4.5005
R23608 DVSS.n780 DVSS.n755 4.5005
R23609 DVSS.n8937 DVSS.n780 4.5005
R23610 DVSS.n780 DVSS.n757 4.5005
R23611 DVSS.n780 DVSS.n756 4.5005
R23612 DVSS.n759 DVSS.n755 4.5005
R23613 DVSS.n8937 DVSS.n759 4.5005
R23614 DVSS.n759 DVSS.n757 4.5005
R23615 DVSS.n759 DVSS.n756 4.5005
R23616 DVSS.n8936 DVSS.n755 4.5005
R23617 DVSS.n8937 DVSS.n8936 4.5005
R23618 DVSS.n8936 DVSS.n757 4.5005
R23619 DVSS.n8936 DVSS.n756 4.5005
R23620 DVSS.n756 DVSS.n754 4.5005
R23621 DVSS.n757 DVSS.n754 4.5005
R23622 DVSS.n755 DVSS.n754 4.5005
R23623 DVSS.n8937 DVSS.n754 4.5005
R23624 DVSS.n8938 DVSS.n756 4.5005
R23625 DVSS.n8938 DVSS.n757 4.5005
R23626 DVSS.n8938 DVSS.n755 4.5005
R23627 DVSS.n8938 DVSS.n8937 4.5005
R23628 DVSS.n7030 DVSS.n6942 4.5005
R23629 DVSS.n6967 DVSS.n6942 4.5005
R23630 DVSS.n6979 DVSS.n6942 4.5005
R23631 DVSS.n6979 DVSS.n6944 4.5005
R23632 DVSS.n7030 DVSS.n6944 4.5005
R23633 DVSS.n7028 DVSS.n6941 4.5005
R23634 DVSS.n7030 DVSS.n6941 4.5005
R23635 DVSS.n7028 DVSS.n6945 4.5005
R23636 DVSS.n7030 DVSS.n6945 4.5005
R23637 DVSS.n7028 DVSS.n6940 4.5005
R23638 DVSS.n7030 DVSS.n6940 4.5005
R23639 DVSS.n7028 DVSS.n6946 4.5005
R23640 DVSS.n7030 DVSS.n6946 4.5005
R23641 DVSS.n7028 DVSS.n6939 4.5005
R23642 DVSS.n7030 DVSS.n6939 4.5005
R23643 DVSS.n7028 DVSS.n6947 4.5005
R23644 DVSS.n7030 DVSS.n6947 4.5005
R23645 DVSS.n7028 DVSS.n6938 4.5005
R23646 DVSS.n7030 DVSS.n6938 4.5005
R23647 DVSS.n7028 DVSS.n6948 4.5005
R23648 DVSS.n7030 DVSS.n6948 4.5005
R23649 DVSS.n7028 DVSS.n6937 4.5005
R23650 DVSS.n7030 DVSS.n6937 4.5005
R23651 DVSS.n7028 DVSS.n6949 4.5005
R23652 DVSS.n7030 DVSS.n6949 4.5005
R23653 DVSS.n7028 DVSS.n6936 4.5005
R23654 DVSS.n7030 DVSS.n6936 4.5005
R23655 DVSS.n7028 DVSS.n6950 4.5005
R23656 DVSS.n7030 DVSS.n6950 4.5005
R23657 DVSS.n7028 DVSS.n6935 4.5005
R23658 DVSS.n7030 DVSS.n6935 4.5005
R23659 DVSS.n7028 DVSS.n6951 4.5005
R23660 DVSS.n7030 DVSS.n6951 4.5005
R23661 DVSS.n7028 DVSS.n6934 4.5005
R23662 DVSS.n7030 DVSS.n6934 4.5005
R23663 DVSS.n7028 DVSS.n6952 4.5005
R23664 DVSS.n7030 DVSS.n6952 4.5005
R23665 DVSS.n7028 DVSS.n6933 4.5005
R23666 DVSS.n7030 DVSS.n6933 4.5005
R23667 DVSS.n7028 DVSS.n6953 4.5005
R23668 DVSS.n7030 DVSS.n6953 4.5005
R23669 DVSS.n7028 DVSS.n6932 4.5005
R23670 DVSS.n7030 DVSS.n6932 4.5005
R23671 DVSS.n7028 DVSS.n6954 4.5005
R23672 DVSS.n7030 DVSS.n6954 4.5005
R23673 DVSS.n7028 DVSS.n6931 4.5005
R23674 DVSS.n7030 DVSS.n6931 4.5005
R23675 DVSS.n7029 DVSS.n7028 4.5005
R23676 DVSS.n7029 DVSS.n6967 4.5005
R23677 DVSS.n7030 DVSS.n7029 4.5005
R23678 DVSS.n8860 DVSS.n807 4.5005
R23679 DVSS.n8860 DVSS.n808 4.5005
R23680 DVSS.n8860 DVSS.n8859 4.5005
R23681 DVSS.n8859 DVSS.n811 4.5005
R23682 DVSS.n811 DVSS.n807 4.5005
R23683 DVSS.n8856 DVSS.n8836 4.5005
R23684 DVSS.n8836 DVSS.n807 4.5005
R23685 DVSS.n8856 DVSS.n8838 4.5005
R23686 DVSS.n8838 DVSS.n807 4.5005
R23687 DVSS.n8856 DVSS.n8834 4.5005
R23688 DVSS.n8834 DVSS.n807 4.5005
R23689 DVSS.n8856 DVSS.n8840 4.5005
R23690 DVSS.n8840 DVSS.n807 4.5005
R23691 DVSS.n8856 DVSS.n8833 4.5005
R23692 DVSS.n8833 DVSS.n807 4.5005
R23693 DVSS.n8856 DVSS.n8842 4.5005
R23694 DVSS.n8842 DVSS.n807 4.5005
R23695 DVSS.n8856 DVSS.n8832 4.5005
R23696 DVSS.n8832 DVSS.n807 4.5005
R23697 DVSS.n8856 DVSS.n8844 4.5005
R23698 DVSS.n8844 DVSS.n807 4.5005
R23699 DVSS.n8856 DVSS.n8831 4.5005
R23700 DVSS.n8831 DVSS.n807 4.5005
R23701 DVSS.n8856 DVSS.n8846 4.5005
R23702 DVSS.n8846 DVSS.n807 4.5005
R23703 DVSS.n8856 DVSS.n8830 4.5005
R23704 DVSS.n8830 DVSS.n807 4.5005
R23705 DVSS.n8856 DVSS.n8848 4.5005
R23706 DVSS.n8848 DVSS.n807 4.5005
R23707 DVSS.n8856 DVSS.n8829 4.5005
R23708 DVSS.n8829 DVSS.n807 4.5005
R23709 DVSS.n8856 DVSS.n8850 4.5005
R23710 DVSS.n8850 DVSS.n807 4.5005
R23711 DVSS.n8856 DVSS.n8828 4.5005
R23712 DVSS.n8828 DVSS.n807 4.5005
R23713 DVSS.n8856 DVSS.n8852 4.5005
R23714 DVSS.n8852 DVSS.n807 4.5005
R23715 DVSS.n8856 DVSS.n8827 4.5005
R23716 DVSS.n8827 DVSS.n807 4.5005
R23717 DVSS.n8856 DVSS.n8854 4.5005
R23718 DVSS.n8854 DVSS.n807 4.5005
R23719 DVSS.n8856 DVSS.n8826 4.5005
R23720 DVSS.n8826 DVSS.n807 4.5005
R23721 DVSS.n8856 DVSS.n8855 4.5005
R23722 DVSS.n8855 DVSS.n807 4.5005
R23723 DVSS.n8857 DVSS.n8856 4.5005
R23724 DVSS.n8857 DVSS.n807 4.5005
R23725 DVSS.n8856 DVSS.n822 4.5005
R23726 DVSS.n822 DVSS.n808 4.5005
R23727 DVSS.n822 DVSS.n807 4.5005
R23728 DVSS.n9063 DVSS.n648 4.5005
R23729 DVSS.n9065 DVSS.n648 4.5005
R23730 DVSS.n9063 DVSS.n9040 4.5005
R23731 DVSS.n9063 DVSS.n9038 4.5005
R23732 DVSS.n9063 DVSS.n9041 4.5005
R23733 DVSS.n9063 DVSS.n9037 4.5005
R23734 DVSS.n9063 DVSS.n9042 4.5005
R23735 DVSS.n9063 DVSS.n9036 4.5005
R23736 DVSS.n9063 DVSS.n9043 4.5005
R23737 DVSS.n9063 DVSS.n9035 4.5005
R23738 DVSS.n9063 DVSS.n9044 4.5005
R23739 DVSS.n9063 DVSS.n9034 4.5005
R23740 DVSS.n9063 DVSS.n9045 4.5005
R23741 DVSS.n9063 DVSS.n9033 4.5005
R23742 DVSS.n9063 DVSS.n9046 4.5005
R23743 DVSS.n9063 DVSS.n9032 4.5005
R23744 DVSS.n9063 DVSS.n9047 4.5005
R23745 DVSS.n9063 DVSS.n9031 4.5005
R23746 DVSS.n9063 DVSS.n9048 4.5005
R23747 DVSS.n9063 DVSS.n9030 4.5005
R23748 DVSS.n9063 DVSS.n9049 4.5005
R23749 DVSS.n9063 DVSS.n9029 4.5005
R23750 DVSS.n9063 DVSS.n9062 4.5005
R23751 DVSS.n9063 DVSS.n9028 4.5005
R23752 DVSS.n9065 DVSS.n9064 4.5005
R23753 DVSS.n9064 DVSS.n9063 4.5005
R23754 DVSS.n9212 DVSS.n515 4.5005
R23755 DVSS.n515 DVSS.n502 4.5005
R23756 DVSS.n9212 DVSS.n518 4.5005
R23757 DVSS.n9212 DVSS.n514 4.5005
R23758 DVSS.n9212 DVSS.n520 4.5005
R23759 DVSS.n9212 DVSS.n513 4.5005
R23760 DVSS.n9212 DVSS.n522 4.5005
R23761 DVSS.n9212 DVSS.n512 4.5005
R23762 DVSS.n9212 DVSS.n524 4.5005
R23763 DVSS.n9212 DVSS.n511 4.5005
R23764 DVSS.n9212 DVSS.n526 4.5005
R23765 DVSS.n9212 DVSS.n510 4.5005
R23766 DVSS.n9212 DVSS.n528 4.5005
R23767 DVSS.n9212 DVSS.n509 4.5005
R23768 DVSS.n9212 DVSS.n530 4.5005
R23769 DVSS.n9212 DVSS.n508 4.5005
R23770 DVSS.n9212 DVSS.n532 4.5005
R23771 DVSS.n9212 DVSS.n507 4.5005
R23772 DVSS.n9212 DVSS.n534 4.5005
R23773 DVSS.n9212 DVSS.n506 4.5005
R23774 DVSS.n9212 DVSS.n536 4.5005
R23775 DVSS.n9212 DVSS.n505 4.5005
R23776 DVSS.n9212 DVSS.n9211 4.5005
R23777 DVSS.n9212 DVSS.n504 4.5005
R23778 DVSS.n9213 DVSS.n502 4.5005
R23779 DVSS.n9213 DVSS.n9212 4.5005
R23780 DVSS.n457 DVSS.n421 4.5005
R23781 DVSS.n421 DVSS.n407 4.5005
R23782 DVSS.n453 DVSS.n421 4.5005
R23783 DVSS.n453 DVSS.n424 4.5005
R23784 DVSS.n457 DVSS.n424 4.5005
R23785 DVSS.n420 DVSS.n408 4.5005
R23786 DVSS.n457 DVSS.n420 4.5005
R23787 DVSS.n426 DVSS.n408 4.5005
R23788 DVSS.n457 DVSS.n426 4.5005
R23789 DVSS.n419 DVSS.n408 4.5005
R23790 DVSS.n457 DVSS.n419 4.5005
R23791 DVSS.n428 DVSS.n408 4.5005
R23792 DVSS.n457 DVSS.n428 4.5005
R23793 DVSS.n418 DVSS.n408 4.5005
R23794 DVSS.n457 DVSS.n418 4.5005
R23795 DVSS.n430 DVSS.n408 4.5005
R23796 DVSS.n457 DVSS.n430 4.5005
R23797 DVSS.n417 DVSS.n408 4.5005
R23798 DVSS.n457 DVSS.n417 4.5005
R23799 DVSS.n432 DVSS.n408 4.5005
R23800 DVSS.n457 DVSS.n432 4.5005
R23801 DVSS.n416 DVSS.n408 4.5005
R23802 DVSS.n457 DVSS.n416 4.5005
R23803 DVSS.n434 DVSS.n408 4.5005
R23804 DVSS.n457 DVSS.n434 4.5005
R23805 DVSS.n415 DVSS.n408 4.5005
R23806 DVSS.n457 DVSS.n415 4.5005
R23807 DVSS.n436 DVSS.n408 4.5005
R23808 DVSS.n457 DVSS.n436 4.5005
R23809 DVSS.n414 DVSS.n408 4.5005
R23810 DVSS.n457 DVSS.n414 4.5005
R23811 DVSS.n438 DVSS.n408 4.5005
R23812 DVSS.n457 DVSS.n438 4.5005
R23813 DVSS.n413 DVSS.n408 4.5005
R23814 DVSS.n457 DVSS.n413 4.5005
R23815 DVSS.n440 DVSS.n408 4.5005
R23816 DVSS.n457 DVSS.n440 4.5005
R23817 DVSS.n412 DVSS.n408 4.5005
R23818 DVSS.n457 DVSS.n412 4.5005
R23819 DVSS.n442 DVSS.n408 4.5005
R23820 DVSS.n457 DVSS.n442 4.5005
R23821 DVSS.n411 DVSS.n408 4.5005
R23822 DVSS.n457 DVSS.n411 4.5005
R23823 DVSS.n456 DVSS.n408 4.5005
R23824 DVSS.n457 DVSS.n456 4.5005
R23825 DVSS.n410 DVSS.n408 4.5005
R23826 DVSS.n457 DVSS.n410 4.5005
R23827 DVSS.n458 DVSS.n408 4.5005
R23828 DVSS.n458 DVSS.n407 4.5005
R23829 DVSS.n458 DVSS.n457 4.5005
R23830 DVSS.n9580 DVSS.n268 4.5005
R23831 DVSS.n9576 DVSS.n268 4.5005
R23832 DVSS.n9583 DVSS.n268 4.5005
R23833 DVSS.n9583 DVSS.n273 4.5005
R23834 DVSS.n9580 DVSS.n273 4.5005
R23835 DVSS.n9558 DVSS.n267 4.5005
R23836 DVSS.n9580 DVSS.n9558 4.5005
R23837 DVSS.n9559 DVSS.n267 4.5005
R23838 DVSS.n9580 DVSS.n9559 4.5005
R23839 DVSS.n9557 DVSS.n267 4.5005
R23840 DVSS.n9580 DVSS.n9557 4.5005
R23841 DVSS.n9560 DVSS.n267 4.5005
R23842 DVSS.n9580 DVSS.n9560 4.5005
R23843 DVSS.n9556 DVSS.n267 4.5005
R23844 DVSS.n9580 DVSS.n9556 4.5005
R23845 DVSS.n9561 DVSS.n267 4.5005
R23846 DVSS.n9580 DVSS.n9561 4.5005
R23847 DVSS.n9555 DVSS.n267 4.5005
R23848 DVSS.n9580 DVSS.n9555 4.5005
R23849 DVSS.n9562 DVSS.n267 4.5005
R23850 DVSS.n9580 DVSS.n9562 4.5005
R23851 DVSS.n9554 DVSS.n267 4.5005
R23852 DVSS.n9580 DVSS.n9554 4.5005
R23853 DVSS.n9563 DVSS.n267 4.5005
R23854 DVSS.n9580 DVSS.n9563 4.5005
R23855 DVSS.n9553 DVSS.n267 4.5005
R23856 DVSS.n9580 DVSS.n9553 4.5005
R23857 DVSS.n9564 DVSS.n267 4.5005
R23858 DVSS.n9580 DVSS.n9564 4.5005
R23859 DVSS.n9552 DVSS.n267 4.5005
R23860 DVSS.n9580 DVSS.n9552 4.5005
R23861 DVSS.n9565 DVSS.n267 4.5005
R23862 DVSS.n9580 DVSS.n9565 4.5005
R23863 DVSS.n9551 DVSS.n267 4.5005
R23864 DVSS.n9580 DVSS.n9551 4.5005
R23865 DVSS.n9566 DVSS.n267 4.5005
R23866 DVSS.n9580 DVSS.n9566 4.5005
R23867 DVSS.n9550 DVSS.n267 4.5005
R23868 DVSS.n9580 DVSS.n9550 4.5005
R23869 DVSS.n9578 DVSS.n267 4.5005
R23870 DVSS.n9580 DVSS.n9578 4.5005
R23871 DVSS.n9549 DVSS.n267 4.5005
R23872 DVSS.n9580 DVSS.n9549 4.5005
R23873 DVSS.n9579 DVSS.n267 4.5005
R23874 DVSS.n9580 DVSS.n9579 4.5005
R23875 DVSS.n9581 DVSS.n267 4.5005
R23876 DVSS.n9581 DVSS.n9580 4.5005
R23877 DVSS.n9546 DVSS.n267 4.5005
R23878 DVSS.n9576 DVSS.n9546 4.5005
R23879 DVSS.n9580 DVSS.n9546 4.5005
R23880 DVSS.n9471 DVSS.n354 4.5005
R23881 DVSS.n354 DVSS.n340 4.5005
R23882 DVSS.n354 DVSS.n343 4.5005
R23883 DVSS.n354 DVSS.n341 4.5005
R23884 DVSS.n355 DVSS.n341 4.5005
R23885 DVSS.n355 DVSS.n343 4.5005
R23886 DVSS.n355 DVSS.n340 4.5005
R23887 DVSS.n9471 DVSS.n355 4.5005
R23888 DVSS.n353 DVSS.n341 4.5005
R23889 DVSS.n353 DVSS.n343 4.5005
R23890 DVSS.n353 DVSS.n340 4.5005
R23891 DVSS.n9471 DVSS.n353 4.5005
R23892 DVSS.n356 DVSS.n341 4.5005
R23893 DVSS.n356 DVSS.n343 4.5005
R23894 DVSS.n356 DVSS.n340 4.5005
R23895 DVSS.n9471 DVSS.n356 4.5005
R23896 DVSS.n352 DVSS.n341 4.5005
R23897 DVSS.n352 DVSS.n343 4.5005
R23898 DVSS.n352 DVSS.n340 4.5005
R23899 DVSS.n9471 DVSS.n352 4.5005
R23900 DVSS.n9471 DVSS.n357 4.5005
R23901 DVSS.n357 DVSS.n340 4.5005
R23902 DVSS.n357 DVSS.n343 4.5005
R23903 DVSS.n357 DVSS.n341 4.5005
R23904 DVSS.n9471 DVSS.n351 4.5005
R23905 DVSS.n351 DVSS.n340 4.5005
R23906 DVSS.n351 DVSS.n343 4.5005
R23907 DVSS.n351 DVSS.n341 4.5005
R23908 DVSS.n9471 DVSS.n358 4.5005
R23909 DVSS.n358 DVSS.n340 4.5005
R23910 DVSS.n358 DVSS.n343 4.5005
R23911 DVSS.n358 DVSS.n341 4.5005
R23912 DVSS.n350 DVSS.n341 4.5005
R23913 DVSS.n350 DVSS.n343 4.5005
R23914 DVSS.n350 DVSS.n340 4.5005
R23915 DVSS.n9471 DVSS.n350 4.5005
R23916 DVSS.n359 DVSS.n341 4.5005
R23917 DVSS.n359 DVSS.n343 4.5005
R23918 DVSS.n359 DVSS.n340 4.5005
R23919 DVSS.n9471 DVSS.n359 4.5005
R23920 DVSS.n349 DVSS.n341 4.5005
R23921 DVSS.n349 DVSS.n343 4.5005
R23922 DVSS.n349 DVSS.n340 4.5005
R23923 DVSS.n9471 DVSS.n349 4.5005
R23924 DVSS.n360 DVSS.n341 4.5005
R23925 DVSS.n360 DVSS.n343 4.5005
R23926 DVSS.n360 DVSS.n340 4.5005
R23927 DVSS.n9471 DVSS.n360 4.5005
R23928 DVSS.n9471 DVSS.n348 4.5005
R23929 DVSS.n348 DVSS.n340 4.5005
R23930 DVSS.n348 DVSS.n343 4.5005
R23931 DVSS.n348 DVSS.n341 4.5005
R23932 DVSS.n9471 DVSS.n361 4.5005
R23933 DVSS.n361 DVSS.n340 4.5005
R23934 DVSS.n361 DVSS.n343 4.5005
R23935 DVSS.n361 DVSS.n341 4.5005
R23936 DVSS.n9471 DVSS.n347 4.5005
R23937 DVSS.n347 DVSS.n340 4.5005
R23938 DVSS.n347 DVSS.n343 4.5005
R23939 DVSS.n347 DVSS.n341 4.5005
R23940 DVSS.n362 DVSS.n341 4.5005
R23941 DVSS.n362 DVSS.n343 4.5005
R23942 DVSS.n362 DVSS.n340 4.5005
R23943 DVSS.n9471 DVSS.n362 4.5005
R23944 DVSS.n346 DVSS.n341 4.5005
R23945 DVSS.n346 DVSS.n343 4.5005
R23946 DVSS.n346 DVSS.n340 4.5005
R23947 DVSS.n9471 DVSS.n346 4.5005
R23948 DVSS.n363 DVSS.n341 4.5005
R23949 DVSS.n363 DVSS.n343 4.5005
R23950 DVSS.n363 DVSS.n340 4.5005
R23951 DVSS.n9471 DVSS.n363 4.5005
R23952 DVSS.n9471 DVSS.n345 4.5005
R23953 DVSS.n345 DVSS.n340 4.5005
R23954 DVSS.n345 DVSS.n343 4.5005
R23955 DVSS.n345 DVSS.n341 4.5005
R23956 DVSS.n9471 DVSS.n364 4.5005
R23957 DVSS.n364 DVSS.n340 4.5005
R23958 DVSS.n364 DVSS.n343 4.5005
R23959 DVSS.n364 DVSS.n341 4.5005
R23960 DVSS.n9471 DVSS.n344 4.5005
R23961 DVSS.n344 DVSS.n340 4.5005
R23962 DVSS.n344 DVSS.n343 4.5005
R23963 DVSS.n344 DVSS.n341 4.5005
R23964 DVSS.n9471 DVSS.n9470 4.5005
R23965 DVSS.n9470 DVSS.n340 4.5005
R23966 DVSS.n9470 DVSS.n343 4.5005
R23967 DVSS.n9470 DVSS.n341 4.5005
R23968 DVSS.n341 DVSS.n339 4.5005
R23969 DVSS.n343 DVSS.n339 4.5005
R23970 DVSS.n340 DVSS.n339 4.5005
R23971 DVSS.n9471 DVSS.n339 4.5005
R23972 DVSS.n9472 DVSS.n341 4.5005
R23973 DVSS.n9472 DVSS.n343 4.5005
R23974 DVSS.n9472 DVSS.n340 4.5005
R23975 DVSS.n9472 DVSS.n9471 4.5005
R23976 DVSS.n9805 DVSS.n84 4.5005
R23977 DVSS.n9843 DVSS.n9805 4.5005
R23978 DVSS.n9841 DVSS.n9805 4.5005
R23979 DVSS.n9843 DVSS.n9807 4.5005
R23980 DVSS.n9841 DVSS.n9807 4.5005
R23981 DVSS.n9843 DVSS.n96 4.5005
R23982 DVSS.n9841 DVSS.n96 4.5005
R23983 DVSS.n9843 DVSS.n9809 4.5005
R23984 DVSS.n9841 DVSS.n9809 4.5005
R23985 DVSS.n9843 DVSS.n95 4.5005
R23986 DVSS.n9841 DVSS.n95 4.5005
R23987 DVSS.n9843 DVSS.n9811 4.5005
R23988 DVSS.n9841 DVSS.n9811 4.5005
R23989 DVSS.n9843 DVSS.n94 4.5005
R23990 DVSS.n9841 DVSS.n94 4.5005
R23991 DVSS.n9843 DVSS.n9813 4.5005
R23992 DVSS.n9841 DVSS.n9813 4.5005
R23993 DVSS.n9843 DVSS.n93 4.5005
R23994 DVSS.n9841 DVSS.n93 4.5005
R23995 DVSS.n9843 DVSS.n9815 4.5005
R23996 DVSS.n9841 DVSS.n9815 4.5005
R23997 DVSS.n9843 DVSS.n92 4.5005
R23998 DVSS.n9841 DVSS.n92 4.5005
R23999 DVSS.n9843 DVSS.n9817 4.5005
R24000 DVSS.n9841 DVSS.n9817 4.5005
R24001 DVSS.n9843 DVSS.n91 4.5005
R24002 DVSS.n9841 DVSS.n91 4.5005
R24003 DVSS.n9843 DVSS.n9819 4.5005
R24004 DVSS.n9841 DVSS.n9819 4.5005
R24005 DVSS.n9843 DVSS.n90 4.5005
R24006 DVSS.n9841 DVSS.n90 4.5005
R24007 DVSS.n9843 DVSS.n9821 4.5005
R24008 DVSS.n9841 DVSS.n9821 4.5005
R24009 DVSS.n9843 DVSS.n89 4.5005
R24010 DVSS.n9841 DVSS.n89 4.5005
R24011 DVSS.n9843 DVSS.n9823 4.5005
R24012 DVSS.n9841 DVSS.n9823 4.5005
R24013 DVSS.n9843 DVSS.n88 4.5005
R24014 DVSS.n9841 DVSS.n88 4.5005
R24015 DVSS.n9843 DVSS.n9825 4.5005
R24016 DVSS.n9841 DVSS.n9825 4.5005
R24017 DVSS.n9843 DVSS.n87 4.5005
R24018 DVSS.n9841 DVSS.n87 4.5005
R24019 DVSS.n9843 DVSS.n9827 4.5005
R24020 DVSS.n9841 DVSS.n9827 4.5005
R24021 DVSS.n9843 DVSS.n86 4.5005
R24022 DVSS.n9841 DVSS.n86 4.5005
R24023 DVSS.n9842 DVSS.n84 4.5005
R24024 DVSS.n9843 DVSS.n9842 4.5005
R24025 DVSS.n9842 DVSS.n9841 4.5005
R24026 DVSS.n8682 DVSS.n8640 4.5005
R24027 DVSS.n8640 DVSS.n964 4.5005
R24028 DVSS.n8680 DVSS.n8640 4.5005
R24029 DVSS.n8656 DVSS.n964 4.5005
R24030 DVSS.n8680 DVSS.n8656 4.5005
R24031 DVSS.n8653 DVSS.n964 4.5005
R24032 DVSS.n8680 DVSS.n8653 4.5005
R24033 DVSS.n8657 DVSS.n964 4.5005
R24034 DVSS.n8680 DVSS.n8657 4.5005
R24035 DVSS.n8652 DVSS.n964 4.5005
R24036 DVSS.n8680 DVSS.n8652 4.5005
R24037 DVSS.n8658 DVSS.n964 4.5005
R24038 DVSS.n8680 DVSS.n8658 4.5005
R24039 DVSS.n8651 DVSS.n964 4.5005
R24040 DVSS.n8680 DVSS.n8651 4.5005
R24041 DVSS.n8659 DVSS.n964 4.5005
R24042 DVSS.n8680 DVSS.n8659 4.5005
R24043 DVSS.n8650 DVSS.n964 4.5005
R24044 DVSS.n8680 DVSS.n8650 4.5005
R24045 DVSS.n8660 DVSS.n964 4.5005
R24046 DVSS.n8680 DVSS.n8660 4.5005
R24047 DVSS.n8649 DVSS.n964 4.5005
R24048 DVSS.n8680 DVSS.n8649 4.5005
R24049 DVSS.n8661 DVSS.n964 4.5005
R24050 DVSS.n8680 DVSS.n8661 4.5005
R24051 DVSS.n8648 DVSS.n964 4.5005
R24052 DVSS.n8680 DVSS.n8648 4.5005
R24053 DVSS.n8662 DVSS.n964 4.5005
R24054 DVSS.n8680 DVSS.n8662 4.5005
R24055 DVSS.n8647 DVSS.n964 4.5005
R24056 DVSS.n8680 DVSS.n8647 4.5005
R24057 DVSS.n8663 DVSS.n964 4.5005
R24058 DVSS.n8680 DVSS.n8663 4.5005
R24059 DVSS.n8646 DVSS.n964 4.5005
R24060 DVSS.n8680 DVSS.n8646 4.5005
R24061 DVSS.n8664 DVSS.n964 4.5005
R24062 DVSS.n8680 DVSS.n8664 4.5005
R24063 DVSS.n8645 DVSS.n964 4.5005
R24064 DVSS.n8680 DVSS.n8645 4.5005
R24065 DVSS.n8665 DVSS.n964 4.5005
R24066 DVSS.n8680 DVSS.n8665 4.5005
R24067 DVSS.n8644 DVSS.n964 4.5005
R24068 DVSS.n8680 DVSS.n8644 4.5005
R24069 DVSS.n8679 DVSS.n964 4.5005
R24070 DVSS.n8680 DVSS.n8679 4.5005
R24071 DVSS.n8643 DVSS.n964 4.5005
R24072 DVSS.n8680 DVSS.n8643 4.5005
R24073 DVSS.n8682 DVSS.n8681 4.5005
R24074 DVSS.n8681 DVSS.n964 4.5005
R24075 DVSS.n8681 DVSS.n8680 4.5005
R24076 DVSS.n8996 DVSS.n737 4.5005
R24077 DVSS.n737 DVSS.n723 4.5005
R24078 DVSS.n737 DVSS.n724 4.5005
R24079 DVSS.n737 DVSS.n725 4.5005
R24080 DVSS.n739 DVSS.n724 4.5005
R24081 DVSS.n739 DVSS.n725 4.5005
R24082 DVSS.n739 DVSS.n723 4.5005
R24083 DVSS.n8996 DVSS.n739 4.5005
R24084 DVSS.n736 DVSS.n724 4.5005
R24085 DVSS.n736 DVSS.n725 4.5005
R24086 DVSS.n736 DVSS.n723 4.5005
R24087 DVSS.n8996 DVSS.n736 4.5005
R24088 DVSS.n740 DVSS.n724 4.5005
R24089 DVSS.n740 DVSS.n725 4.5005
R24090 DVSS.n740 DVSS.n723 4.5005
R24091 DVSS.n8996 DVSS.n740 4.5005
R24092 DVSS.n8996 DVSS.n735 4.5005
R24093 DVSS.n735 DVSS.n723 4.5005
R24094 DVSS.n735 DVSS.n724 4.5005
R24095 DVSS.n735 DVSS.n725 4.5005
R24096 DVSS.n8996 DVSS.n741 4.5005
R24097 DVSS.n741 DVSS.n723 4.5005
R24098 DVSS.n741 DVSS.n724 4.5005
R24099 DVSS.n741 DVSS.n725 4.5005
R24100 DVSS.n8996 DVSS.n734 4.5005
R24101 DVSS.n734 DVSS.n723 4.5005
R24102 DVSS.n734 DVSS.n724 4.5005
R24103 DVSS.n734 DVSS.n725 4.5005
R24104 DVSS.n742 DVSS.n724 4.5005
R24105 DVSS.n742 DVSS.n725 4.5005
R24106 DVSS.n742 DVSS.n723 4.5005
R24107 DVSS.n8996 DVSS.n742 4.5005
R24108 DVSS.n733 DVSS.n724 4.5005
R24109 DVSS.n733 DVSS.n725 4.5005
R24110 DVSS.n733 DVSS.n723 4.5005
R24111 DVSS.n8996 DVSS.n733 4.5005
R24112 DVSS.n743 DVSS.n724 4.5005
R24113 DVSS.n743 DVSS.n725 4.5005
R24114 DVSS.n743 DVSS.n723 4.5005
R24115 DVSS.n8996 DVSS.n743 4.5005
R24116 DVSS.n732 DVSS.n724 4.5005
R24117 DVSS.n732 DVSS.n725 4.5005
R24118 DVSS.n732 DVSS.n723 4.5005
R24119 DVSS.n8996 DVSS.n732 4.5005
R24120 DVSS.n8996 DVSS.n744 4.5005
R24121 DVSS.n744 DVSS.n723 4.5005
R24122 DVSS.n744 DVSS.n724 4.5005
R24123 DVSS.n744 DVSS.n725 4.5005
R24124 DVSS.n8996 DVSS.n731 4.5005
R24125 DVSS.n731 DVSS.n723 4.5005
R24126 DVSS.n731 DVSS.n724 4.5005
R24127 DVSS.n731 DVSS.n725 4.5005
R24128 DVSS.n8996 DVSS.n745 4.5005
R24129 DVSS.n745 DVSS.n723 4.5005
R24130 DVSS.n745 DVSS.n724 4.5005
R24131 DVSS.n745 DVSS.n725 4.5005
R24132 DVSS.n730 DVSS.n724 4.5005
R24133 DVSS.n730 DVSS.n725 4.5005
R24134 DVSS.n730 DVSS.n723 4.5005
R24135 DVSS.n8996 DVSS.n730 4.5005
R24136 DVSS.n746 DVSS.n724 4.5005
R24137 DVSS.n746 DVSS.n725 4.5005
R24138 DVSS.n746 DVSS.n723 4.5005
R24139 DVSS.n8996 DVSS.n746 4.5005
R24140 DVSS.n729 DVSS.n724 4.5005
R24141 DVSS.n729 DVSS.n725 4.5005
R24142 DVSS.n729 DVSS.n723 4.5005
R24143 DVSS.n8996 DVSS.n729 4.5005
R24144 DVSS.n8996 DVSS.n747 4.5005
R24145 DVSS.n747 DVSS.n723 4.5005
R24146 DVSS.n747 DVSS.n724 4.5005
R24147 DVSS.n747 DVSS.n725 4.5005
R24148 DVSS.n8996 DVSS.n728 4.5005
R24149 DVSS.n728 DVSS.n723 4.5005
R24150 DVSS.n728 DVSS.n724 4.5005
R24151 DVSS.n728 DVSS.n725 4.5005
R24152 DVSS.n8996 DVSS.n748 4.5005
R24153 DVSS.n748 DVSS.n723 4.5005
R24154 DVSS.n748 DVSS.n724 4.5005
R24155 DVSS.n748 DVSS.n725 4.5005
R24156 DVSS.n8996 DVSS.n727 4.5005
R24157 DVSS.n727 DVSS.n723 4.5005
R24158 DVSS.n727 DVSS.n724 4.5005
R24159 DVSS.n727 DVSS.n725 4.5005
R24160 DVSS.n8995 DVSS.n724 4.5005
R24161 DVSS.n8995 DVSS.n725 4.5005
R24162 DVSS.n8995 DVSS.n723 4.5005
R24163 DVSS.n8996 DVSS.n8995 4.5005
R24164 DVSS.n8997 DVSS.n724 4.5005
R24165 DVSS.n8997 DVSS.n725 4.5005
R24166 DVSS.n8997 DVSS.n723 4.5005
R24167 DVSS.n8997 DVSS.n8996 4.5005
R24168 DVSS.n724 DVSS.n719 4.5005
R24169 DVSS.n725 DVSS.n719 4.5005
R24170 DVSS.n723 DVSS.n719 4.5005
R24171 DVSS.n8996 DVSS.n719 4.5005
R24172 DVSS.n915 DVSS.n898 4.5005
R24173 DVSS.n8717 DVSS.n915 4.5005
R24174 DVSS.n8715 DVSS.n915 4.5005
R24175 DVSS.n8717 DVSS.n919 4.5005
R24176 DVSS.n8715 DVSS.n919 4.5005
R24177 DVSS.n8717 DVSS.n914 4.5005
R24178 DVSS.n8715 DVSS.n914 4.5005
R24179 DVSS.n8717 DVSS.n922 4.5005
R24180 DVSS.n8715 DVSS.n922 4.5005
R24181 DVSS.n8717 DVSS.n913 4.5005
R24182 DVSS.n8715 DVSS.n913 4.5005
R24183 DVSS.n8717 DVSS.n925 4.5005
R24184 DVSS.n8715 DVSS.n925 4.5005
R24185 DVSS.n8717 DVSS.n912 4.5005
R24186 DVSS.n8715 DVSS.n912 4.5005
R24187 DVSS.n8717 DVSS.n928 4.5005
R24188 DVSS.n8715 DVSS.n928 4.5005
R24189 DVSS.n8717 DVSS.n911 4.5005
R24190 DVSS.n8715 DVSS.n911 4.5005
R24191 DVSS.n8717 DVSS.n931 4.5005
R24192 DVSS.n8715 DVSS.n931 4.5005
R24193 DVSS.n8717 DVSS.n910 4.5005
R24194 DVSS.n8715 DVSS.n910 4.5005
R24195 DVSS.n8717 DVSS.n934 4.5005
R24196 DVSS.n8715 DVSS.n934 4.5005
R24197 DVSS.n8717 DVSS.n909 4.5005
R24198 DVSS.n8715 DVSS.n909 4.5005
R24199 DVSS.n8717 DVSS.n937 4.5005
R24200 DVSS.n8715 DVSS.n937 4.5005
R24201 DVSS.n8717 DVSS.n908 4.5005
R24202 DVSS.n8715 DVSS.n908 4.5005
R24203 DVSS.n8717 DVSS.n940 4.5005
R24204 DVSS.n8715 DVSS.n940 4.5005
R24205 DVSS.n8717 DVSS.n907 4.5005
R24206 DVSS.n8715 DVSS.n907 4.5005
R24207 DVSS.n8717 DVSS.n943 4.5005
R24208 DVSS.n8715 DVSS.n943 4.5005
R24209 DVSS.n8717 DVSS.n906 4.5005
R24210 DVSS.n8715 DVSS.n906 4.5005
R24211 DVSS.n8717 DVSS.n946 4.5005
R24212 DVSS.n8715 DVSS.n946 4.5005
R24213 DVSS.n8717 DVSS.n905 4.5005
R24214 DVSS.n8715 DVSS.n905 4.5005
R24215 DVSS.n8717 DVSS.n8716 4.5005
R24216 DVSS.n8716 DVSS.n8715 4.5005
R24217 DVSS.n8717 DVSS.n904 4.5005
R24218 DVSS.n8715 DVSS.n904 4.5005
R24219 DVSS.n898 DVSS.n712 4.5005
R24220 DVSS.n8717 DVSS.n712 4.5005
R24221 DVSS.n8715 DVSS.n712 4.5005
R24222 DVSS.n852 DVSS.n835 4.5005
R24223 DVSS.n8752 DVSS.n852 4.5005
R24224 DVSS.n8750 DVSS.n852 4.5005
R24225 DVSS.n8752 DVSS.n856 4.5005
R24226 DVSS.n8750 DVSS.n856 4.5005
R24227 DVSS.n8752 DVSS.n851 4.5005
R24228 DVSS.n8750 DVSS.n851 4.5005
R24229 DVSS.n8752 DVSS.n859 4.5005
R24230 DVSS.n8750 DVSS.n859 4.5005
R24231 DVSS.n8752 DVSS.n850 4.5005
R24232 DVSS.n8750 DVSS.n850 4.5005
R24233 DVSS.n8752 DVSS.n862 4.5005
R24234 DVSS.n8750 DVSS.n862 4.5005
R24235 DVSS.n8752 DVSS.n849 4.5005
R24236 DVSS.n8750 DVSS.n849 4.5005
R24237 DVSS.n8752 DVSS.n865 4.5005
R24238 DVSS.n8750 DVSS.n865 4.5005
R24239 DVSS.n8752 DVSS.n848 4.5005
R24240 DVSS.n8750 DVSS.n848 4.5005
R24241 DVSS.n8752 DVSS.n868 4.5005
R24242 DVSS.n8750 DVSS.n868 4.5005
R24243 DVSS.n8752 DVSS.n847 4.5005
R24244 DVSS.n8750 DVSS.n847 4.5005
R24245 DVSS.n8752 DVSS.n871 4.5005
R24246 DVSS.n8750 DVSS.n871 4.5005
R24247 DVSS.n8752 DVSS.n846 4.5005
R24248 DVSS.n8750 DVSS.n846 4.5005
R24249 DVSS.n8752 DVSS.n874 4.5005
R24250 DVSS.n8750 DVSS.n874 4.5005
R24251 DVSS.n8752 DVSS.n845 4.5005
R24252 DVSS.n8750 DVSS.n845 4.5005
R24253 DVSS.n8752 DVSS.n877 4.5005
R24254 DVSS.n8750 DVSS.n877 4.5005
R24255 DVSS.n8752 DVSS.n844 4.5005
R24256 DVSS.n8750 DVSS.n844 4.5005
R24257 DVSS.n8752 DVSS.n880 4.5005
R24258 DVSS.n8750 DVSS.n880 4.5005
R24259 DVSS.n8752 DVSS.n843 4.5005
R24260 DVSS.n8750 DVSS.n843 4.5005
R24261 DVSS.n8752 DVSS.n883 4.5005
R24262 DVSS.n8750 DVSS.n883 4.5005
R24263 DVSS.n8752 DVSS.n842 4.5005
R24264 DVSS.n8750 DVSS.n842 4.5005
R24265 DVSS.n8752 DVSS.n8751 4.5005
R24266 DVSS.n8751 DVSS.n8750 4.5005
R24267 DVSS.n8752 DVSS.n841 4.5005
R24268 DVSS.n8750 DVSS.n841 4.5005
R24269 DVSS.n835 DVSS.n705 4.5005
R24270 DVSS.n8752 DVSS.n705 4.5005
R24271 DVSS.n8750 DVSS.n705 4.5005
R24272 DVSS.n9027 DVSS.n662 4.5005
R24273 DVSS.n9027 DVSS.n9026 4.5005
R24274 DVSS.n9026 DVSS.n677 4.5005
R24275 DVSS.n9026 DVSS.n674 4.5005
R24276 DVSS.n9026 DVSS.n679 4.5005
R24277 DVSS.n9026 DVSS.n673 4.5005
R24278 DVSS.n9026 DVSS.n681 4.5005
R24279 DVSS.n9026 DVSS.n672 4.5005
R24280 DVSS.n9026 DVSS.n683 4.5005
R24281 DVSS.n9026 DVSS.n671 4.5005
R24282 DVSS.n9026 DVSS.n685 4.5005
R24283 DVSS.n9026 DVSS.n670 4.5005
R24284 DVSS.n9026 DVSS.n687 4.5005
R24285 DVSS.n9026 DVSS.n669 4.5005
R24286 DVSS.n9026 DVSS.n689 4.5005
R24287 DVSS.n9026 DVSS.n668 4.5005
R24288 DVSS.n9026 DVSS.n691 4.5005
R24289 DVSS.n9026 DVSS.n667 4.5005
R24290 DVSS.n9026 DVSS.n693 4.5005
R24291 DVSS.n9026 DVSS.n666 4.5005
R24292 DVSS.n9026 DVSS.n695 4.5005
R24293 DVSS.n9026 DVSS.n665 4.5005
R24294 DVSS.n9026 DVSS.n697 4.5005
R24295 DVSS.n9026 DVSS.n664 4.5005
R24296 DVSS.n9025 DVSS.n662 4.5005
R24297 DVSS.n9026 DVSS.n9025 4.5005
R24298 DVSS.n9214 DVSS.n495 4.5005
R24299 DVSS.n9214 DVSS.n499 4.5005
R24300 DVSS.n9216 DVSS.n499 4.5005
R24301 DVSS.n9218 DVSS.n499 4.5005
R24302 DVSS.n9220 DVSS.n499 4.5005
R24303 DVSS.n9222 DVSS.n499 4.5005
R24304 DVSS.n9224 DVSS.n499 4.5005
R24305 DVSS.n9226 DVSS.n499 4.5005
R24306 DVSS.n9228 DVSS.n499 4.5005
R24307 DVSS.n9230 DVSS.n499 4.5005
R24308 DVSS.n9232 DVSS.n499 4.5005
R24309 DVSS.n9234 DVSS.n499 4.5005
R24310 DVSS.n9236 DVSS.n499 4.5005
R24311 DVSS.n9238 DVSS.n499 4.5005
R24312 DVSS.n9240 DVSS.n499 4.5005
R24313 DVSS.n9242 DVSS.n499 4.5005
R24314 DVSS.n9244 DVSS.n499 4.5005
R24315 DVSS.n9246 DVSS.n499 4.5005
R24316 DVSS.n9248 DVSS.n499 4.5005
R24317 DVSS.n9250 DVSS.n499 4.5005
R24318 DVSS.n9252 DVSS.n499 4.5005
R24319 DVSS.n9254 DVSS.n499 4.5005
R24320 DVSS.n9256 DVSS.n499 4.5005
R24321 DVSS.n9258 DVSS.n499 4.5005
R24322 DVSS.n495 DVSS.n386 4.5005
R24323 DVSS.n499 DVSS.n386 4.5005
R24324 DVSS.n459 DVSS.n392 4.5005
R24325 DVSS.n459 DVSS.n393 4.5005
R24326 DVSS.n9367 DVSS.n459 4.5005
R24327 DVSS.n462 DVSS.n393 4.5005
R24328 DVSS.n9367 DVSS.n462 4.5005
R24329 DVSS.n405 DVSS.n393 4.5005
R24330 DVSS.n9367 DVSS.n405 4.5005
R24331 DVSS.n464 DVSS.n393 4.5005
R24332 DVSS.n9367 DVSS.n464 4.5005
R24333 DVSS.n404 DVSS.n393 4.5005
R24334 DVSS.n9367 DVSS.n404 4.5005
R24335 DVSS.n466 DVSS.n393 4.5005
R24336 DVSS.n9367 DVSS.n466 4.5005
R24337 DVSS.n403 DVSS.n393 4.5005
R24338 DVSS.n9367 DVSS.n403 4.5005
R24339 DVSS.n468 DVSS.n393 4.5005
R24340 DVSS.n9367 DVSS.n468 4.5005
R24341 DVSS.n402 DVSS.n393 4.5005
R24342 DVSS.n9367 DVSS.n402 4.5005
R24343 DVSS.n470 DVSS.n393 4.5005
R24344 DVSS.n9367 DVSS.n470 4.5005
R24345 DVSS.n401 DVSS.n393 4.5005
R24346 DVSS.n9367 DVSS.n401 4.5005
R24347 DVSS.n472 DVSS.n393 4.5005
R24348 DVSS.n9367 DVSS.n472 4.5005
R24349 DVSS.n400 DVSS.n393 4.5005
R24350 DVSS.n9367 DVSS.n400 4.5005
R24351 DVSS.n474 DVSS.n393 4.5005
R24352 DVSS.n9367 DVSS.n474 4.5005
R24353 DVSS.n399 DVSS.n393 4.5005
R24354 DVSS.n9367 DVSS.n399 4.5005
R24355 DVSS.n476 DVSS.n393 4.5005
R24356 DVSS.n9367 DVSS.n476 4.5005
R24357 DVSS.n398 DVSS.n393 4.5005
R24358 DVSS.n9367 DVSS.n398 4.5005
R24359 DVSS.n478 DVSS.n393 4.5005
R24360 DVSS.n9367 DVSS.n478 4.5005
R24361 DVSS.n397 DVSS.n393 4.5005
R24362 DVSS.n9367 DVSS.n397 4.5005
R24363 DVSS.n480 DVSS.n393 4.5005
R24364 DVSS.n9367 DVSS.n480 4.5005
R24365 DVSS.n396 DVSS.n393 4.5005
R24366 DVSS.n9367 DVSS.n396 4.5005
R24367 DVSS.n9366 DVSS.n393 4.5005
R24368 DVSS.n9367 DVSS.n9366 4.5005
R24369 DVSS.n395 DVSS.n393 4.5005
R24370 DVSS.n9367 DVSS.n395 4.5005
R24371 DVSS.n9368 DVSS.n392 4.5005
R24372 DVSS.n9368 DVSS.n393 4.5005
R24373 DVSS.n9368 DVSS.n9367 4.5005
R24374 DVSS.n9545 DVSS.n285 4.5005
R24375 DVSS.n9545 DVSS.n287 4.5005
R24376 DVSS.n9545 DVSS.n9544 4.5005
R24377 DVSS.n302 DVSS.n287 4.5005
R24378 DVSS.n9544 DVSS.n302 4.5005
R24379 DVSS.n299 DVSS.n287 4.5005
R24380 DVSS.n9544 DVSS.n299 4.5005
R24381 DVSS.n304 DVSS.n287 4.5005
R24382 DVSS.n9544 DVSS.n304 4.5005
R24383 DVSS.n298 DVSS.n287 4.5005
R24384 DVSS.n9544 DVSS.n298 4.5005
R24385 DVSS.n306 DVSS.n287 4.5005
R24386 DVSS.n9544 DVSS.n306 4.5005
R24387 DVSS.n297 DVSS.n287 4.5005
R24388 DVSS.n9544 DVSS.n297 4.5005
R24389 DVSS.n308 DVSS.n287 4.5005
R24390 DVSS.n9544 DVSS.n308 4.5005
R24391 DVSS.n296 DVSS.n287 4.5005
R24392 DVSS.n9544 DVSS.n296 4.5005
R24393 DVSS.n310 DVSS.n287 4.5005
R24394 DVSS.n9544 DVSS.n310 4.5005
R24395 DVSS.n295 DVSS.n287 4.5005
R24396 DVSS.n9544 DVSS.n295 4.5005
R24397 DVSS.n312 DVSS.n287 4.5005
R24398 DVSS.n9544 DVSS.n312 4.5005
R24399 DVSS.n294 DVSS.n287 4.5005
R24400 DVSS.n9544 DVSS.n294 4.5005
R24401 DVSS.n314 DVSS.n287 4.5005
R24402 DVSS.n9544 DVSS.n314 4.5005
R24403 DVSS.n293 DVSS.n287 4.5005
R24404 DVSS.n9544 DVSS.n293 4.5005
R24405 DVSS.n316 DVSS.n287 4.5005
R24406 DVSS.n9544 DVSS.n316 4.5005
R24407 DVSS.n292 DVSS.n287 4.5005
R24408 DVSS.n9544 DVSS.n292 4.5005
R24409 DVSS.n318 DVSS.n287 4.5005
R24410 DVSS.n9544 DVSS.n318 4.5005
R24411 DVSS.n291 DVSS.n287 4.5005
R24412 DVSS.n9544 DVSS.n291 4.5005
R24413 DVSS.n320 DVSS.n287 4.5005
R24414 DVSS.n9544 DVSS.n320 4.5005
R24415 DVSS.n290 DVSS.n287 4.5005
R24416 DVSS.n9544 DVSS.n290 4.5005
R24417 DVSS.n322 DVSS.n287 4.5005
R24418 DVSS.n9544 DVSS.n322 4.5005
R24419 DVSS.n289 DVSS.n287 4.5005
R24420 DVSS.n9544 DVSS.n289 4.5005
R24421 DVSS.n9543 DVSS.n285 4.5005
R24422 DVSS.n9543 DVSS.n287 4.5005
R24423 DVSS.n9544 DVSS.n9543 4.5005
R24424 DVSS.n9888 DVSS.n36 4.5005
R24425 DVSS.n49 DVSS.n36 4.5005
R24426 DVSS.n9886 DVSS.n36 4.5005
R24427 DVSS.n50 DVSS.n36 4.5005
R24428 DVSS.n50 DVSS.n37 4.5005
R24429 DVSS.n9886 DVSS.n37 4.5005
R24430 DVSS.n49 DVSS.n37 4.5005
R24431 DVSS.n9888 DVSS.n37 4.5005
R24432 DVSS.n50 DVSS.n35 4.5005
R24433 DVSS.n9886 DVSS.n35 4.5005
R24434 DVSS.n49 DVSS.n35 4.5005
R24435 DVSS.n9888 DVSS.n35 4.5005
R24436 DVSS.n50 DVSS.n38 4.5005
R24437 DVSS.n9886 DVSS.n38 4.5005
R24438 DVSS.n49 DVSS.n38 4.5005
R24439 DVSS.n9888 DVSS.n38 4.5005
R24440 DVSS.n9888 DVSS.n34 4.5005
R24441 DVSS.n49 DVSS.n34 4.5005
R24442 DVSS.n9886 DVSS.n34 4.5005
R24443 DVSS.n50 DVSS.n34 4.5005
R24444 DVSS.n9888 DVSS.n39 4.5005
R24445 DVSS.n49 DVSS.n39 4.5005
R24446 DVSS.n9886 DVSS.n39 4.5005
R24447 DVSS.n50 DVSS.n39 4.5005
R24448 DVSS.n9888 DVSS.n33 4.5005
R24449 DVSS.n49 DVSS.n33 4.5005
R24450 DVSS.n9886 DVSS.n33 4.5005
R24451 DVSS.n50 DVSS.n33 4.5005
R24452 DVSS.n50 DVSS.n40 4.5005
R24453 DVSS.n9886 DVSS.n40 4.5005
R24454 DVSS.n49 DVSS.n40 4.5005
R24455 DVSS.n9888 DVSS.n40 4.5005
R24456 DVSS.n50 DVSS.n32 4.5005
R24457 DVSS.n9886 DVSS.n32 4.5005
R24458 DVSS.n49 DVSS.n32 4.5005
R24459 DVSS.n9888 DVSS.n32 4.5005
R24460 DVSS.n50 DVSS.n41 4.5005
R24461 DVSS.n9886 DVSS.n41 4.5005
R24462 DVSS.n49 DVSS.n41 4.5005
R24463 DVSS.n9888 DVSS.n41 4.5005
R24464 DVSS.n50 DVSS.n31 4.5005
R24465 DVSS.n9886 DVSS.n31 4.5005
R24466 DVSS.n49 DVSS.n31 4.5005
R24467 DVSS.n9888 DVSS.n31 4.5005
R24468 DVSS.n9888 DVSS.n42 4.5005
R24469 DVSS.n49 DVSS.n42 4.5005
R24470 DVSS.n9886 DVSS.n42 4.5005
R24471 DVSS.n50 DVSS.n42 4.5005
R24472 DVSS.n9888 DVSS.n30 4.5005
R24473 DVSS.n49 DVSS.n30 4.5005
R24474 DVSS.n9886 DVSS.n30 4.5005
R24475 DVSS.n50 DVSS.n30 4.5005
R24476 DVSS.n9888 DVSS.n43 4.5005
R24477 DVSS.n49 DVSS.n43 4.5005
R24478 DVSS.n9886 DVSS.n43 4.5005
R24479 DVSS.n50 DVSS.n43 4.5005
R24480 DVSS.n50 DVSS.n29 4.5005
R24481 DVSS.n9886 DVSS.n29 4.5005
R24482 DVSS.n49 DVSS.n29 4.5005
R24483 DVSS.n9888 DVSS.n29 4.5005
R24484 DVSS.n50 DVSS.n44 4.5005
R24485 DVSS.n9886 DVSS.n44 4.5005
R24486 DVSS.n49 DVSS.n44 4.5005
R24487 DVSS.n9888 DVSS.n44 4.5005
R24488 DVSS.n50 DVSS.n28 4.5005
R24489 DVSS.n9886 DVSS.n28 4.5005
R24490 DVSS.n49 DVSS.n28 4.5005
R24491 DVSS.n9888 DVSS.n28 4.5005
R24492 DVSS.n9888 DVSS.n45 4.5005
R24493 DVSS.n49 DVSS.n45 4.5005
R24494 DVSS.n9886 DVSS.n45 4.5005
R24495 DVSS.n50 DVSS.n45 4.5005
R24496 DVSS.n9888 DVSS.n27 4.5005
R24497 DVSS.n49 DVSS.n27 4.5005
R24498 DVSS.n9886 DVSS.n27 4.5005
R24499 DVSS.n50 DVSS.n27 4.5005
R24500 DVSS.n9888 DVSS.n46 4.5005
R24501 DVSS.n49 DVSS.n46 4.5005
R24502 DVSS.n9886 DVSS.n46 4.5005
R24503 DVSS.n50 DVSS.n46 4.5005
R24504 DVSS.n9888 DVSS.n26 4.5005
R24505 DVSS.n49 DVSS.n26 4.5005
R24506 DVSS.n9886 DVSS.n26 4.5005
R24507 DVSS.n50 DVSS.n26 4.5005
R24508 DVSS.n50 DVSS.n47 4.5005
R24509 DVSS.n9886 DVSS.n47 4.5005
R24510 DVSS.n49 DVSS.n47 4.5005
R24511 DVSS.n9888 DVSS.n47 4.5005
R24512 DVSS.n50 DVSS.n25 4.5005
R24513 DVSS.n9886 DVSS.n25 4.5005
R24514 DVSS.n49 DVSS.n25 4.5005
R24515 DVSS.n9888 DVSS.n25 4.5005
R24516 DVSS.n9887 DVSS.n50 4.5005
R24517 DVSS.n9887 DVSS.n9886 4.5005
R24518 DVSS.n9887 DVSS.n49 4.5005
R24519 DVSS.n9888 DVSS.n9887 4.5005
R24520 DVSS.n9934 DVSS.n17 4.5005
R24521 DVSS.n19 DVSS.n17 4.5005
R24522 DVSS.n9932 DVSS.n17 4.5005
R24523 DVSS.n9909 DVSS.n19 4.5005
R24524 DVSS.n9932 DVSS.n9909 4.5005
R24525 DVSS.n9908 DVSS.n19 4.5005
R24526 DVSS.n9932 DVSS.n9908 4.5005
R24527 DVSS.n9910 DVSS.n19 4.5005
R24528 DVSS.n9932 DVSS.n9910 4.5005
R24529 DVSS.n9907 DVSS.n19 4.5005
R24530 DVSS.n9932 DVSS.n9907 4.5005
R24531 DVSS.n9911 DVSS.n19 4.5005
R24532 DVSS.n9932 DVSS.n9911 4.5005
R24533 DVSS.n9906 DVSS.n19 4.5005
R24534 DVSS.n9932 DVSS.n9906 4.5005
R24535 DVSS.n9912 DVSS.n19 4.5005
R24536 DVSS.n9932 DVSS.n9912 4.5005
R24537 DVSS.n9905 DVSS.n19 4.5005
R24538 DVSS.n9932 DVSS.n9905 4.5005
R24539 DVSS.n9913 DVSS.n19 4.5005
R24540 DVSS.n9932 DVSS.n9913 4.5005
R24541 DVSS.n9904 DVSS.n19 4.5005
R24542 DVSS.n9932 DVSS.n9904 4.5005
R24543 DVSS.n9914 DVSS.n19 4.5005
R24544 DVSS.n9932 DVSS.n9914 4.5005
R24545 DVSS.n9903 DVSS.n19 4.5005
R24546 DVSS.n9932 DVSS.n9903 4.5005
R24547 DVSS.n9915 DVSS.n19 4.5005
R24548 DVSS.n9932 DVSS.n9915 4.5005
R24549 DVSS.n9902 DVSS.n19 4.5005
R24550 DVSS.n9932 DVSS.n9902 4.5005
R24551 DVSS.n9916 DVSS.n19 4.5005
R24552 DVSS.n9932 DVSS.n9916 4.5005
R24553 DVSS.n9901 DVSS.n19 4.5005
R24554 DVSS.n9932 DVSS.n9901 4.5005
R24555 DVSS.n9917 DVSS.n19 4.5005
R24556 DVSS.n9932 DVSS.n9917 4.5005
R24557 DVSS.n9900 DVSS.n19 4.5005
R24558 DVSS.n9932 DVSS.n9900 4.5005
R24559 DVSS.n9918 DVSS.n19 4.5005
R24560 DVSS.n9932 DVSS.n9918 4.5005
R24561 DVSS.n9899 DVSS.n19 4.5005
R24562 DVSS.n9932 DVSS.n9899 4.5005
R24563 DVSS.n9931 DVSS.n19 4.5005
R24564 DVSS.n9932 DVSS.n9931 4.5005
R24565 DVSS.n9898 DVSS.n19 4.5005
R24566 DVSS.n9932 DVSS.n9898 4.5005
R24567 DVSS.n9934 DVSS.n9933 4.5005
R24568 DVSS.n9933 DVSS.n19 4.5005
R24569 DVSS.n9933 DVSS.n9932 4.5005
R24570 DVSS.n8186 DVSS.n8185 4.38021
R24571 DVSS.n5923 DVSS.n5922 4.38021
R24572 DVSS.n4477 DVSS.n3016 4.38021
R24573 DVSS.n6747 DVSS.n1915 4.38021
R24574 DVSS.n5870 DVSS.n3016 4.36815
R24575 DVSS.n5922 DVSS.n5921 4.36815
R24576 DVSS.n5921 DVSS.n2912 4.36815
R24577 DVSS.n5871 DVSS.n5870 4.36815
R24578 DVSS.n5871 DVSS.n2978 4.36815
R24579 DVSS.n2968 DVSS.n2912 4.36815
R24580 DVSS.n5896 DVSS.n2980 4.36815
R24581 DVSS.n5900 DVSS.n2112 4.36815
R24582 DVSS.n2112 DVSS.n1752 4.36815
R24583 DVSS.n2980 DVSS.n2979 4.36815
R24584 DVSS.n2979 DVSS.n1915 4.36815
R24585 DVSS.n8185 DVSS.n1752 4.36815
R24586 DVSS.n7248 DVSS.n7247 2.2505
R24587 DVSS.n7247 DVSS.n7246 2.2505
R24588 DVSS.n7253 DVSS.n6645 2.2505
R24589 DVSS.n7253 DVSS.n7252 2.2505
R24590 DVSS.n4930 DVSS.n4929 2.24726
R24591 DVSS.n4927 DVSS.n4918 2.24726
R24592 DVSS.n2921 DVSS.n2914 2.24726
R24593 DVSS.n5917 DVSS.n2913 2.24726
R24594 DVSS.n5375 DVSS.n5370 2.24726
R24595 DVSS.n5374 DVSS.n5371 2.24726
R24596 DVSS.n2965 DVSS.n2963 2.24726
R24597 DVSS.n2967 DVSS.n2966 2.24726
R24598 DVSS.n2974 DVSS.n2972 2.24726
R24599 DVSS.n2976 DVSS.n2975 2.24726
R24600 DVSS.n2117 DVSS.n2114 2.24726
R24601 DVSS.n2115 DVSS.n2111 2.24726
R24602 DVSS.n7701 DVSS.n2106 2.24726
R24603 DVSS.n7703 DVSS.n7702 2.24726
R24604 DVSS.n1760 DVSS.n1759 2.24726
R24605 DVSS.n1757 DVSS.n1753 2.24726
R24606 DVSS.n8062 DVSS.n1912 2.24726
R24607 DVSS.n7371 DVSS.n2587 2.24726
R24608 DVSS.n7376 DVSS.n2578 2.24726
R24609 DVSS.n5892 DVSS.n5891 2.24726
R24610 DVSS.n5882 DVSS.n5881 2.24726
R24611 DVSS.n5874 DVSS.n3013 2.24726
R24612 DVSS.n5873 DVSS.n5872 2.24726
R24613 DVSS.n5866 DVSS.n3019 2.24726
R24614 DVSS.n3024 DVSS.n3018 2.24726
R24615 DVSS.n4446 DVSS.n4445 2.24726
R24616 DVSS.n4444 DVSS.n4443 2.24726
R24617 DVSS.n3865 DVSS.n3860 2.2467
R24618 DVSS.n4196 DVSS.n4191 2.2467
R24619 DVSS.n4800 DVSS.n3712 2.2467
R24620 DVSS.n4807 DVSS.n3704 2.2467
R24621 DVSS.n4820 DVSS.n3670 2.2467
R24622 DVSS.n4842 DVSS.n4841 2.2467
R24623 DVSS.n4834 DVSS.n3626 2.2467
R24624 DVSS.n4979 DVSS.n3589 2.2467
R24625 DVSS.n4221 DVSS.n3859 2.2467
R24626 DVSS.n4221 DVSS.n3867 2.2467
R24627 DVSS.n4431 DVSS.n3869 2.2467
R24628 DVSS.n4432 DVSS.n4431 2.2467
R24629 DVSS.n4799 DVSS.n4798 2.2467
R24630 DVSS.n4798 DVSS.n3711 2.2467
R24631 DVSS.n3707 DVSS.n3702 2.2467
R24632 DVSS.n4819 DVSS.n3669 2.2467
R24633 DVSS.n4827 DVSS.n4826 2.2467
R24634 DVSS.n4828 DVSS.n4827 2.2467
R24635 DVSS.n4831 DVSS.n3623 2.2467
R24636 DVSS.n4836 DVSS.n3623 2.2467
R24637 DVSS.n4975 DVSS.n4974 2.2467
R24638 DVSS.n4974 DVSS.n3592 2.2467
R24639 DVSS.n3873 DVSS.n3051 2.2467
R24640 DVSS.n3885 DVSS.n3884 2.2467
R24641 DVSS.n4007 DVSS.n4001 2.2467
R24642 DVSS.n4101 DVSS.n4100 2.2467
R24643 DVSS.n5000 DVSS.n3565 2.2467
R24644 DVSS.n3574 DVSS.n3571 2.2467
R24645 DVSS.n3584 DVSS.n3581 2.2467
R24646 DVSS.n4985 DVSS.n4982 2.2467
R24647 DVSS.n4174 DVSS.n4173 2.2467
R24648 DVSS.n4174 DVSS.n3881 2.2467
R24649 DVSS.n4006 DVSS.n4005 2.2467
R24650 DVSS.n4005 DVSS.n4000 2.2467
R24651 DVSS.n4096 DVSS.n4095 2.2467
R24652 DVSS.n3568 DVSS.n3564 2.2467
R24653 DVSS.n3576 DVSS.n3570 2.2467
R24654 DVSS.n3577 DVSS.n3576 2.2467
R24655 DVSS.n3586 DVSS.n3580 2.2467
R24656 DVSS.n3587 DVSS.n3586 2.2467
R24657 DVSS.n4987 DVSS.n4981 2.2467
R24658 DVSS.n4988 DVSS.n4987 2.2467
R24659 DVSS.n3535 DVSS.n3065 2.2467
R24660 DVSS.n3544 DVSS.n3111 2.2467
R24661 DVSS.n3552 DVSS.n3156 2.2467
R24662 DVSS.n3557 DVSS.n3188 2.2467
R24663 DVSS.n5030 DVSS.n5021 2.2467
R24664 DVSS.n3348 DVSS.n3324 2.2467
R24665 DVSS.n3358 DVSS.n3353 2.2467
R24666 DVSS.n3368 DVSS.n3363 2.2467
R24667 DVSS.n3543 DVSS.n3542 2.2467
R24668 DVSS.n3542 DVSS.n3530 2.2467
R24669 DVSS.n3551 DVSS.n3550 2.2467
R24670 DVSS.n3550 DVSS.n3525 2.2467
R24671 DVSS.n3556 DVSS.n3521 2.2467
R24672 DVSS.n5026 DVSS.n5023 2.2467
R24673 DVSS.n5391 DVSS.n5390 2.2467
R24674 DVSS.n5391 DVSS.n3345 2.2467
R24675 DVSS.n5071 DVSS.n3352 2.2467
R24676 DVSS.n5071 DVSS.n3360 2.2467
R24677 DVSS.n5368 DVSS.n3362 2.2467
R24678 DVSS.n5369 DVSS.n5368 2.2467
R24679 DVSS.n5680 DVSS.n3250 2.2467
R24680 DVSS.n5687 DVSS.n3241 2.2467
R24681 DVSS.n5497 DVSS.n3293 2.2467
R24682 DVSS.n5504 DVSS.n3301 2.2467
R24683 DVSS.n5516 DVSS.n3309 2.2467
R24684 DVSS.n3255 DVSS.n3066 2.2467
R24685 DVSS.n3254 DVSS.n3113 2.2467
R24686 DVSS.n3245 DVSS.n3157 2.2467
R24687 DVSS.n5696 DVSS.n3230 2.2467
R24688 DVSS.n5489 DVSS.n5488 2.2467
R24689 DVSS.n5401 DVSS.n5395 2.2467
R24690 DVSS.n3321 DVSS.n3315 2.2467
R24691 DVSS.n5512 DVSS.n3311 2.2467
R24692 DVSS.n5657 DVSS.n3261 2.2467
R24693 DVSS.n5647 DVSS.n3268 2.2467
R24694 DVSS.n5540 DVSS.n3291 2.2467
R24695 DVSS.n5530 DVSS.n3299 2.2467
R24696 DVSS.n5521 DVSS.n3306 2.2467
R24697 DVSS.n5670 DVSS.n3257 2.2467
R24698 DVSS.n5662 DVSS.n3263 2.2467
R24699 DVSS.n5652 DVSS.n3270 2.2467
R24700 DVSS.n5642 DVSS.n3273 2.2467
R24701 DVSS.n5638 DVSS.n3286 2.2467
R24702 DVSS.n5545 DVSS.n3294 2.2467
R24703 DVSS.n5535 DVSS.n3302 2.2467
R24704 DVSS.n5526 DVSS.n5517 2.2467
R24705 DVSS.n2677 DVSS.n2594 2.2467
R24706 DVSS.n2683 DVSS.n2601 2.2467
R24707 DVSS.n2690 DVSS.n2609 2.2467
R24708 DVSS.n2710 DVSS.n2086 2.2467
R24709 DVSS.n2719 DVSS.n2094 2.2467
R24710 DVSS.n2727 DVSS.n2102 2.2467
R24711 DVSS.n2674 DVSS.n2521 2.2467
R24712 DVSS.n2667 DVSS.n2464 2.2467
R24713 DVSS.n2659 DVSS.n2400 2.2467
R24714 DVSS.n2695 DVSS.n2335 2.2467
R24715 DVSS.n2702 DVSS.n2305 2.2467
R24716 DVSS.n2713 DVSS.n2252 2.2467
R24717 DVSS.n2722 DVSS.n2210 2.2467
R24718 DVSS.n2730 DVSS.n2176 2.2467
R24719 DVSS.n7354 DVSS.n2592 2.2467
R24720 DVSS.n7345 DVSS.n2599 2.2467
R24721 DVSS.n7335 DVSS.n2607 2.2467
R24722 DVSS.n7848 DVSS.n2084 2.2467
R24723 DVSS.n2092 DVSS.n1814 2.2467
R24724 DVSS.n7711 DVSS.n2100 2.2467
R24725 DVSS.n7359 DVSS.n2595 2.2467
R24726 DVSS.n7350 DVSS.n2602 2.2467
R24727 DVSS.n7340 DVSS.n2610 2.2467
R24728 DVSS.n7330 DVSS.n2613 2.2467
R24729 DVSS.n7326 DVSS.n7325 2.2467
R24730 DVSS.n7853 DVSS.n2087 2.2467
R24731 DVSS.n7723 DVSS.n2095 2.2467
R24732 DVSS.n7716 DVSS.n2103 2.2467
R24733 DVSS.n8073 DVSS.n1904 2.2467
R24734 DVSS.n8079 DVSS.n1895 2.2467
R24735 DVSS.n8086 DVSS.n1885 2.2467
R24736 DVSS.n8108 DVSS.n1859 2.2467
R24737 DVSS.n8115 DVSS.n1553 2.2467
R24738 DVSS.n1839 DVSS.n1560 2.2467
R24739 DVSS.n1908 DVSS.n1901 2.2467
R24740 DVSS.n1899 DVSS.n1892 2.2467
R24741 DVSS.n1889 DVSS.n1882 2.2467
R24742 DVSS.n8095 DVSS.n1874 2.2467
R24743 DVSS.n8100 DVSS.n8099 2.2467
R24744 DVSS.n1863 DVSS.n1856 2.2467
R24745 DVSS.n8119 DVSS.n1833 2.2467
R24746 DVSS.n1849 DVSS.n1841 2.2467
R24747 DVSS.n8332 DVSS.n1444 2.24623
R24748 DVSS.n8269 DVSS.n8268 2.24623
R24749 DVSS.n8265 DVSS.n8264 2.24623
R24750 DVSS.n8322 DVSS.n1448 2.24623
R24751 DVSS.n8324 DVSS.n1445 2.24623
R24752 DVSS.n1462 DVSS.n1460 2.24623
R24753 DVSS.n8310 DVSS.n1464 2.24623
R24754 DVSS.n8213 DVSS.n1530 2.24623
R24755 DVSS.n7142 DVSS.n7139 2.24623
R24756 DVSS.n1487 DVSS.n1486 2.24623
R24757 DVSS.n8240 DVSS.n1511 2.24623
R24758 DVSS.n8232 DVSS.n1515 2.24623
R24759 DVSS.n8234 DVSS.n1512 2.24623
R24760 DVSS.n8245 DVSS.n8242 2.24623
R24761 DVSS.n1488 DVSS.n1483 2.24623
R24762 DVSS.n7113 DVSS.n7078 2.24623
R24763 DVSS.n7138 DVSS.n6651 2.24623
R24764 DVSS.n7137 DVSS.n6652 2.24623
R24765 DVSS.n8448 DVSS.n1321 2.24623
R24766 DVSS.n1129 DVSS.n1126 2.24623
R24767 DVSS.n1139 DVSS.n1136 2.24623
R24768 DVSS.n1132 DVSS.n1131 2.24623
R24769 DVSS.n1140 DVSS.n1138 2.24623
R24770 DVSS.n1322 DVSS.n1320 2.24623
R24771 DVSS.n1255 DVSS.n1254 2.24623
R24772 DVSS.n1248 DVSS.n1247 2.24623
R24773 DVSS.n1233 DVSS.n1232 2.24623
R24774 DVSS.n8492 DVSS.n1099 2.24623
R24775 DVSS.n1423 DVSS.n1419 2.24623
R24776 DVSS.n8368 DVSS.n8363 2.24623
R24777 DVSS.n1548 DVSS.n1543 2.24623
R24778 DVSS.n8334 DVSS.n1437 2.24623
R24779 DVSS.n7120 DVSS.n7076 2.24623
R24780 DVSS.n7074 DVSS.n7072 2.24623
R24781 DVSS.n1159 DVSS.n1154 2.24623
R24782 DVSS.n1184 DVSS.n1181 2.24623
R24783 DVSS.n1187 DVSS.n1186 2.24623
R24784 DVSS.n1226 DVSS.n1225 2.24623
R24785 DVSS.n717 DVSS.n714 2.24623
R24786 DVSS.n9002 DVSS.n9001 2.24623
R24787 DVSS.n720 DVSS.n714 2.24623
R24788 DVSS.n335 DVSS.n332 2.24623
R24789 DVSS.n9537 DVSS.n9536 2.24623
R24790 DVSS.n333 DVSS.n332 2.24623
R24791 DVSS.n8885 DVSS.n782 2.24623
R24792 DVSS.n8881 DVSS.n781 2.24623
R24793 DVSS.n9417 DVSS.n365 2.24623
R24794 DVSS.n9416 DVSS.n9415 2.24623
R24795 DVSS.n1537 DVSS.n1536 2.24623
R24796 DVSS.n1534 DVSS.n1531 2.24623
R24797 DVSS.n8203 DVSS.n8202 2.24623
R24798 DVSS.n8196 DVSS.n8195 2.24623
R24799 DVSS.n1559 DVSS.n1556 2.24623
R24800 DVSS.n1552 DVSS.n1542 2.24623
R24801 DVSS.n8191 DVSS.n8190 2.24623
R24802 DVSS.n5909 DVSS.n2964 2.24623
R24803 DVSS.n5907 DVSS.n2961 2.24623
R24804 DVSS.n5904 DVSS.n2973 2.24623
R24805 DVSS.n5902 DVSS.n2970 2.24623
R24806 DVSS.n7696 DVSS.n2110 2.24623
R24807 DVSS.n7698 DVSS.n2113 2.24623
R24808 DVSS.n7708 DVSS.n2107 2.24623
R24809 DVSS.n7706 DVSS.n7705 2.24623
R24810 DVSS.n8182 DVSS.n8181 2.24623
R24811 DVSS.n8184 DVSS.n1754 2.24623
R24812 DVSS.n6665 DVSS.n6660 2.24623
R24813 DVSS.n7071 DVSS.n6656 2.24623
R24814 DVSS.n7070 DVSS.n6657 2.24623
R24815 DVSS.n6664 DVSS.n6661 2.24623
R24816 DVSS.n6747 DVSS.n6746 2.24623
R24817 DVSS.n8067 DVSS.n8066 2.24623
R24818 DVSS.n8065 DVSS.n8064 2.24623
R24819 DVSS.n8067 DVSS.n8063 2.24623
R24820 DVSS.n7363 DVSS.n2588 2.24623
R24821 DVSS.n7365 DVSS.n2589 2.24623
R24822 DVSS.n7370 DVSS.n2588 2.24623
R24823 DVSS.n2583 DVSS.n2579 2.24623
R24824 DVSS.n2585 DVSS.n2580 2.24623
R24825 DVSS.n7375 DVSS.n2579 2.24623
R24826 DVSS.n5895 DVSS.n2983 2.24623
R24827 DVSS.n2988 DVSS.n2982 2.24623
R24828 DVSS.n5895 DVSS.n2981 2.24623
R24829 DVSS.n5889 DVSS.n5888 2.24623
R24830 DVSS.n5886 DVSS.n5883 2.24623
R24831 DVSS.n5889 DVSS.n2992 2.24623
R24832 DVSS.n5883 DVSS.n2990 2.24623
R24833 DVSS.n2984 DVSS.n2982 2.24623
R24834 DVSS.n2586 DVSS.n2585 2.24623
R24835 DVSS.n7366 DVSS.n7365 2.24623
R24836 DVSS.n8065 DVSS.n1913 2.24623
R24837 DVSS.n8880 DVSS.n783 2.24582
R24838 DVSS.n9414 DVSS.n156 2.24582
R24839 DVSS.n3414 DVSS.n3405 2.24552
R24840 DVSS.n3416 DVSS.n3401 2.24552
R24841 DVSS.n3417 DVSS.n3405 2.24552
R24842 DVSS.n3419 DVSS.n3401 2.24552
R24843 DVSS.n3420 DVSS.n3405 2.24552
R24844 DVSS.n3422 DVSS.n3401 2.24552
R24845 DVSS.n5128 DVSS.n5081 2.24552
R24846 DVSS.n5130 DVSS.n5069 2.24552
R24847 DVSS.n5128 DVSS.n5079 2.24552
R24848 DVSS.n5130 DVSS.n5070 2.24552
R24849 DVSS.n5128 DVSS.n5076 2.24552
R24850 DVSS.n1832 DVSS.n1815 2.24552
R24851 DVSS.n8123 DVSS.n1813 2.24552
R24852 DVSS.n1832 DVSS.n1830 2.24552
R24853 DVSS.n8123 DVSS.n1812 2.24552
R24854 DVSS.n1832 DVSS.n1829 2.24552
R24855 DVSS.n8123 DVSS.n1811 2.24552
R24856 DVSS.n1832 DVSS.n1828 2.24552
R24857 DVSS.n8123 DVSS.n1810 2.24552
R24858 DVSS.n1832 DVSS.n1827 2.24552
R24859 DVSS.n8123 DVSS.n1809 2.24552
R24860 DVSS.n1115 DVSS.n1105 2.24552
R24861 DVSS.n1117 DVSS.n1106 2.24552
R24862 DVSS.n1118 DVSS.n1105 2.24552
R24863 DVSS.n1120 DVSS.n1106 2.24552
R24864 DVSS.n1110 DVSS.n1107 2.24552
R24865 DVSS.n1122 DVSS.n1106 2.24552
R24866 DVSS.n1123 DVSS.n1105 2.24552
R24867 DVSS.n1125 DVSS.n1106 2.24552
R24868 DVSS.n4886 DVSS.n3631 2.24552
R24869 DVSS.n4882 DVSS.n3625 2.24552
R24870 DVSS.n4888 DVSS.n3618 2.24552
R24871 DVSS.n4884 DVSS.n3625 2.24552
R24872 DVSS.n4888 DVSS.n3617 2.24552
R24873 DVSS.n3628 DVSS.n3625 2.24552
R24874 DVSS.n3666 DVSS.n3655 2.24552
R24875 DVSS.n4850 DVSS.n3654 2.24552
R24876 DVSS.n3666 DVSS.n3664 2.24552
R24877 DVSS.n4850 DVSS.n3653 2.24552
R24878 DVSS.n3666 DVSS.n3663 2.24552
R24879 DVSS.n4850 DVSS.n3652 2.24552
R24880 DVSS.n3449 DVSS.n3440 2.24552
R24881 DVSS.n3451 DVSS.n3436 2.24552
R24882 DVSS.n3452 DVSS.n3440 2.24552
R24883 DVSS.n3454 DVSS.n3436 2.24552
R24884 DVSS.n3455 DVSS.n3440 2.24552
R24885 DVSS.n3457 DVSS.n3436 2.24552
R24886 DVSS.n3334 DVSS.n3327 2.24552
R24887 DVSS.n5393 DVSS.n3336 2.24552
R24888 DVSS.n3340 DVSS.n3327 2.24552
R24889 DVSS.n5393 DVSS.n3342 2.24552
R24890 DVSS.n3337 DVSS.n3327 2.24552
R24891 DVSS.n7844 DVSS.n7728 2.24552
R24892 DVSS.n7738 DVSS.n7729 2.24552
R24893 DVSS.n7844 DVSS.n7750 2.24552
R24894 DVSS.n7740 DVSS.n7729 2.24552
R24895 DVSS.n7844 DVSS.n7749 2.24552
R24896 DVSS.n7742 DVSS.n7729 2.24552
R24897 DVSS.n7844 DVSS.n7748 2.24552
R24898 DVSS.n7744 DVSS.n7729 2.24552
R24899 DVSS.n7844 DVSS.n7747 2.24552
R24900 DVSS.n7746 DVSS.n7729 2.24552
R24901 DVSS.n8340 DVSS.n1425 2.24552
R24902 DVSS.n8342 DVSS.n1426 2.24552
R24903 DVSS.n8343 DVSS.n1425 2.24552
R24904 DVSS.n1433 DVSS.n1426 2.24552
R24905 DVSS.n1431 DVSS.n1427 2.24552
R24906 DVSS.n8345 DVSS.n1425 2.24552
R24907 DVSS.n8346 DVSS.n1426 2.24552
R24908 DVSS.n1429 DVSS.n1425 2.24552
R24909 DVSS.n4786 DVSS.n3719 2.24552
R24910 DVSS.n4788 DVSS.n3720 2.24552
R24911 DVSS.n4789 DVSS.n3719 2.24552
R24912 DVSS.n4791 DVSS.n3720 2.24552
R24913 DVSS.n4792 DVSS.n3719 2.24552
R24914 DVSS.n4794 DVSS.n3720 2.24552
R24915 DVSS.n3946 DVSS.n3945 2.24552
R24916 DVSS.n3950 DVSS.n3948 2.24552
R24917 DVSS.n3946 DVSS.n3944 2.24552
R24918 DVSS.n3950 DVSS.n3949 2.24552
R24919 DVSS.n3946 DVSS.n3943 2.24552
R24920 DVSS.n3950 DVSS.n3942 2.24552
R24921 DVSS.n3148 DVSS.n3141 2.24552
R24922 DVSS.n5775 DVSS.n5773 2.24552
R24923 DVSS.n3150 DVSS.n3141 2.24552
R24924 DVSS.n5775 DVSS.n5774 2.24552
R24925 DVSS.n3152 DVSS.n3141 2.24552
R24926 DVSS.n2017 DVSS.n2010 2.24552
R24927 DVSS.n7972 DVSS.n7968 2.24552
R24928 DVSS.n2019 DVSS.n2010 2.24552
R24929 DVSS.n7972 DVSS.n7969 2.24552
R24930 DVSS.n2021 DVSS.n2010 2.24552
R24931 DVSS.n7972 DVSS.n7970 2.24552
R24932 DVSS.n2023 DVSS.n2010 2.24552
R24933 DVSS.n7972 DVSS.n7971 2.24552
R24934 DVSS.n2025 DVSS.n2010 2.24552
R24935 DVSS.n7973 DVSS.n7972 2.24552
R24936 DVSS.n8435 DVSS.n1343 2.24552
R24937 DVSS.n1336 DVSS.n1326 2.24552
R24938 DVSS.n8435 DVSS.n1342 2.24552
R24939 DVSS.n1338 DVSS.n1326 2.24552
R24940 DVSS.n1340 DVSS.n1327 2.24552
R24941 DVSS.n8436 DVSS.n8435 2.24552
R24942 DVSS.n8437 DVSS.n1326 2.24552
R24943 DVSS.n8435 DVSS.n1325 2.24552
R24944 DVSS.n4419 DVSS.n4199 2.24552
R24945 DVSS.n4421 DVSS.n4200 2.24552
R24946 DVSS.n4422 DVSS.n4199 2.24552
R24947 DVSS.n4424 DVSS.n4200 2.24552
R24948 DVSS.n4425 DVSS.n4199 2.24552
R24949 DVSS.n4427 DVSS.n4200 2.24552
R24950 DVSS.n4176 DVSS.n3887 2.24552
R24951 DVSS.n4178 DVSS.n3888 2.24552
R24952 DVSS.n4179 DVSS.n3887 2.24552
R24953 DVSS.n4181 DVSS.n3888 2.24552
R24954 DVSS.n4182 DVSS.n3887 2.24552
R24955 DVSS.n4184 DVSS.n3888 2.24552
R24956 DVSS.n3117 DVSS.n3116 2.24552
R24957 DVSS.n5811 DVSS.n5809 2.24552
R24958 DVSS.n3117 DVSS.n3115 2.24552
R24959 DVSS.n5811 DVSS.n5810 2.24552
R24960 DVSS.n3117 DVSS.n3114 2.24552
R24961 DVSS.n1983 DVSS.n1976 2.24552
R24962 DVSS.n8011 DVSS.n8007 2.24552
R24963 DVSS.n1985 DVSS.n1976 2.24552
R24964 DVSS.n8011 DVSS.n8008 2.24552
R24965 DVSS.n1987 DVSS.n1976 2.24552
R24966 DVSS.n8011 DVSS.n8009 2.24552
R24967 DVSS.n1989 DVSS.n1976 2.24552
R24968 DVSS.n8011 DVSS.n8010 2.24552
R24969 DVSS.n1991 DVSS.n1976 2.24552
R24970 DVSS.n8012 DVSS.n8011 2.24552
R24971 DVSS.n1172 DVSS.n1161 2.24552
R24972 DVSS.n1174 DVSS.n1162 2.24552
R24973 DVSS.n1175 DVSS.n1161 2.24552
R24974 DVSS.n1168 DVSS.n1162 2.24552
R24975 DVSS.n1166 DVSS.n1163 2.24552
R24976 DVSS.n1177 DVSS.n1161 2.24552
R24977 DVSS.n1178 DVSS.n1162 2.24552
R24978 DVSS.n1180 DVSS.n1161 2.24552
R24979 DVSS.n7417 DVSS.n7416 2.24552
R24980 DVSS.n2431 DVSS.n2417 2.24552
R24981 DVSS.n2433 DVSS.n2413 2.24552
R24982 DVSS.n2434 DVSS.n2417 2.24552
R24983 DVSS.n2436 DVSS.n2413 2.24552
R24984 DVSS.n2437 DVSS.n2417 2.24552
R24985 DVSS.n2439 DVSS.n2413 2.24552
R24986 DVSS.n2440 DVSS.n2417 2.24552
R24987 DVSS.n2442 DVSS.n2413 2.24552
R24988 DVSS.n2443 DVSS.n2417 2.24552
R24989 DVSS.n2445 DVSS.n2413 2.24552
R24990 DVSS.n2446 DVSS.n2417 2.24552
R24991 DVSS.n2448 DVSS.n2413 2.24552
R24992 DVSS.n2449 DVSS.n2417 2.24552
R24993 DVSS.n2451 DVSS.n2413 2.24552
R24994 DVSS.n2452 DVSS.n2417 2.24552
R24995 DVSS.n2454 DVSS.n2413 2.24552
R24996 DVSS.n2455 DVSS.n2417 2.24552
R24997 DVSS.n2457 DVSS.n2413 2.24552
R24998 DVSS.n2458 DVSS.n2417 2.24552
R24999 DVSS.n2460 DVSS.n2413 2.24552
R25000 DVSS.n2461 DVSS.n2417 2.24552
R25001 DVSS.n2463 DVSS.n2413 2.24552
R25002 DVSS.n2366 DVSS.n2352 2.24552
R25003 DVSS.n2367 DVSS.n2348 2.24552
R25004 DVSS.n2369 DVSS.n2352 2.24552
R25005 DVSS.n2370 DVSS.n2348 2.24552
R25006 DVSS.n2372 DVSS.n2352 2.24552
R25007 DVSS.n2373 DVSS.n2348 2.24552
R25008 DVSS.n2375 DVSS.n2352 2.24552
R25009 DVSS.n2376 DVSS.n2348 2.24552
R25010 DVSS.n2378 DVSS.n2352 2.24552
R25011 DVSS.n2379 DVSS.n2348 2.24552
R25012 DVSS.n2381 DVSS.n2352 2.24552
R25013 DVSS.n2382 DVSS.n2348 2.24552
R25014 DVSS.n2384 DVSS.n2352 2.24552
R25015 DVSS.n2385 DVSS.n2348 2.24552
R25016 DVSS.n2387 DVSS.n2352 2.24552
R25017 DVSS.n2388 DVSS.n2348 2.24552
R25018 DVSS.n2390 DVSS.n2352 2.24552
R25019 DVSS.n2391 DVSS.n2348 2.24552
R25020 DVSS.n2393 DVSS.n2352 2.24552
R25021 DVSS.n2394 DVSS.n2348 2.24552
R25022 DVSS.n2396 DVSS.n2352 2.24552
R25023 DVSS.n2397 DVSS.n2348 2.24552
R25024 DVSS.n2399 DVSS.n2352 2.24552
R25025 DVSS.n7553 DVSS.n7543 2.24552
R25026 DVSS.n7558 DVSS.n2249 2.24552
R25027 DVSS.n7553 DVSS.n7544 2.24552
R25028 DVSS.n7558 DVSS.n2248 2.24552
R25029 DVSS.n7553 DVSS.n7545 2.24552
R25030 DVSS.n7558 DVSS.n2247 2.24552
R25031 DVSS.n7553 DVSS.n7546 2.24552
R25032 DVSS.n7558 DVSS.n2246 2.24552
R25033 DVSS.n7553 DVSS.n7547 2.24552
R25034 DVSS.n7558 DVSS.n2245 2.24552
R25035 DVSS.n7553 DVSS.n7548 2.24552
R25036 DVSS.n7558 DVSS.n2244 2.24552
R25037 DVSS.n7553 DVSS.n7549 2.24552
R25038 DVSS.n7558 DVSS.n2243 2.24552
R25039 DVSS.n7553 DVSS.n7550 2.24552
R25040 DVSS.n7558 DVSS.n2242 2.24552
R25041 DVSS.n7553 DVSS.n7551 2.24552
R25042 DVSS.n7558 DVSS.n2241 2.24552
R25043 DVSS.n7553 DVSS.n7552 2.24552
R25044 DVSS.n7558 DVSS.n2240 2.24552
R25045 DVSS.n7554 DVSS.n7553 2.24552
R25046 DVSS.n7558 DVSS.n2239 2.24552
R25047 DVSS.n7553 DVSS.n2251 2.24552
R25048 DVSS.n7611 DVSS.n7601 2.24552
R25049 DVSS.n7616 DVSS.n2207 2.24552
R25050 DVSS.n7611 DVSS.n7602 2.24552
R25051 DVSS.n7616 DVSS.n2206 2.24552
R25052 DVSS.n7611 DVSS.n7603 2.24552
R25053 DVSS.n7616 DVSS.n2205 2.24552
R25054 DVSS.n7611 DVSS.n7604 2.24552
R25055 DVSS.n7616 DVSS.n2204 2.24552
R25056 DVSS.n7611 DVSS.n7605 2.24552
R25057 DVSS.n7616 DVSS.n2203 2.24552
R25058 DVSS.n7611 DVSS.n7606 2.24552
R25059 DVSS.n7616 DVSS.n2202 2.24552
R25060 DVSS.n7611 DVSS.n7607 2.24552
R25061 DVSS.n7616 DVSS.n2201 2.24552
R25062 DVSS.n7611 DVSS.n7608 2.24552
R25063 DVSS.n7616 DVSS.n2200 2.24552
R25064 DVSS.n7611 DVSS.n7609 2.24552
R25065 DVSS.n7616 DVSS.n2199 2.24552
R25066 DVSS.n7611 DVSS.n7610 2.24552
R25067 DVSS.n7616 DVSS.n2198 2.24552
R25068 DVSS.n7612 DVSS.n7611 2.24552
R25069 DVSS.n7616 DVSS.n2197 2.24552
R25070 DVSS.n7611 DVSS.n2209 2.24552
R25071 DVSS.n2487 DVSS.n2469 2.24552
R25072 DVSS.n2488 DVSS.n2473 2.24552
R25073 DVSS.n2490 DVSS.n2469 2.24552
R25074 DVSS.n2491 DVSS.n2473 2.24552
R25075 DVSS.n2493 DVSS.n2469 2.24552
R25076 DVSS.n2494 DVSS.n2473 2.24552
R25077 DVSS.n2496 DVSS.n2469 2.24552
R25078 DVSS.n2497 DVSS.n2473 2.24552
R25079 DVSS.n2499 DVSS.n2469 2.24552
R25080 DVSS.n2500 DVSS.n2473 2.24552
R25081 DVSS.n2502 DVSS.n2469 2.24552
R25082 DVSS.n2503 DVSS.n2473 2.24552
R25083 DVSS.n2505 DVSS.n2469 2.24552
R25084 DVSS.n2506 DVSS.n2473 2.24552
R25085 DVSS.n2508 DVSS.n2469 2.24552
R25086 DVSS.n2509 DVSS.n2473 2.24552
R25087 DVSS.n2511 DVSS.n2469 2.24552
R25088 DVSS.n2512 DVSS.n2473 2.24552
R25089 DVSS.n2514 DVSS.n2469 2.24552
R25090 DVSS.n2515 DVSS.n2473 2.24552
R25091 DVSS.n2517 DVSS.n2469 2.24552
R25092 DVSS.n2518 DVSS.n2473 2.24552
R25093 DVSS.n2520 DVSS.n2469 2.24552
R25094 DVSS.n1957 DVSS.n1950 2.24552
R25095 DVSS.n8034 DVSS.n8030 2.24552
R25096 DVSS.n1959 DVSS.n1950 2.24552
R25097 DVSS.n8034 DVSS.n8031 2.24552
R25098 DVSS.n1961 DVSS.n1950 2.24552
R25099 DVSS.n8034 DVSS.n8032 2.24552
R25100 DVSS.n1963 DVSS.n1950 2.24552
R25101 DVSS.n8034 DVSS.n8033 2.24552
R25102 DVSS.n1965 DVSS.n1950 2.24552
R25103 DVSS.n8035 DVSS.n8034 2.24552
R25104 DVSS.n6689 DVSS.n6666 2.24552
R25105 DVSS.n6676 DVSS.n6667 2.24552
R25106 DVSS.n6689 DVSS.n6688 2.24552
R25107 DVSS.n6678 DVSS.n6667 2.24552
R25108 DVSS.n6689 DVSS.n6687 2.24552
R25109 DVSS.n6680 DVSS.n6667 2.24552
R25110 DVSS.n6689 DVSS.n6686 2.24552
R25111 DVSS.n6682 DVSS.n6667 2.24552
R25112 DVSS.n6689 DVSS.n6685 2.24552
R25113 DVSS.n6684 DVSS.n6667 2.24552
R25114 DVSS.n4227 DVSS.n4223 2.24552
R25115 DVSS.n4260 DVSS.n4218 2.24552
R25116 DVSS.n4253 DVSS.n4223 2.24552
R25117 DVSS.n4260 DVSS.n4219 2.24552
R25118 DVSS.n4255 DVSS.n4223 2.24552
R25119 DVSS.n4260 DVSS.n4220 2.24552
R25120 DVSS.n4517 DVSS.n4515 2.24552
R25121 DVSS.n4519 DVSS.n3820 2.24552
R25122 DVSS.n4517 DVSS.n4513 2.24552
R25123 DVSS.n4519 DVSS.n3821 2.24552
R25124 DVSS.n4517 DVSS.n4510 2.24552
R25125 DVSS.n3822 DVSS.n3815 2.24552
R25126 DVSS.n4580 DVSS.n3799 2.24552
R25127 DVSS.n4582 DVSS.n3800 2.24552
R25128 DVSS.n4583 DVSS.n3799 2.24552
R25129 DVSS.n4585 DVSS.n3800 2.24552
R25130 DVSS.n4586 DVSS.n3799 2.24552
R25131 DVSS.n3803 DVSS.n3801 2.24552
R25132 DVSS.n4782 DVSS.n3746 2.24552
R25133 DVSS.n3737 DVSS.n3728 2.24552
R25134 DVSS.n4782 DVSS.n3745 2.24552
R25135 DVSS.n3739 DVSS.n3728 2.24552
R25136 DVSS.n4782 DVSS.n3727 2.24552
R25137 DVSS.n3741 DVSS.n3729 2.24552
R25138 DVSS.n6000 DVSS.n2780 2.24552
R25139 DVSS.n2790 DVSS.n2781 2.24552
R25140 DVSS.n6000 DVSS.n2793 2.24552
R25141 DVSS.n2792 DVSS.n2781 2.24552
R25142 DVSS.n6001 DVSS.n6000 2.24552
R25143 DVSS.n2784 DVSS.n2782 2.24552
R25144 DVSS.n5973 DVSS.n2836 2.24552
R25145 DVSS.n2830 DVSS.n2828 2.24552
R25146 DVSS.n5973 DVSS.n2835 2.24552
R25147 DVSS.n2830 DVSS.n2829 2.24552
R25148 DVSS.n5973 DVSS.n2834 2.24552
R25149 DVSS.n2833 DVSS.n2832 2.24552
R25150 DVSS.n2863 DVSS.n2862 2.24552
R25151 DVSS.n5958 DVSS.n5956 2.24552
R25152 DVSS.n2863 DVSS.n2861 2.24552
R25153 DVSS.n5958 DVSS.n5957 2.24552
R25154 DVSS.n2863 DVSS.n2860 2.24552
R25155 DVSS.n4962 DVSS.n3598 2.24552
R25156 DVSS.n4964 DVSS.n3599 2.24552
R25157 DVSS.n4965 DVSS.n3598 2.24552
R25158 DVSS.n4967 DVSS.n3599 2.24552
R25159 DVSS.n4968 DVSS.n3598 2.24552
R25160 DVSS.n4970 DVSS.n3599 2.24552
R25161 DVSS.n3389 DVSS.n3378 2.24552
R25162 DVSS.n5349 DVSS.n5348 2.24552
R25163 DVSS.n3391 DVSS.n3378 2.24552
R25164 DVSS.n5350 DVSS.n5349 2.24552
R25165 DVSS.n5351 DVSS.n3378 2.24552
R25166 DVSS.n5349 DVSS.n3377 2.24552
R25167 DVSS.n5356 DVSS.n3373 2.24552
R25168 DVSS.n5366 DVSS.n5358 2.24552
R25169 DVSS.n5362 DVSS.n3373 2.24552
R25170 DVSS.n5366 DVSS.n5364 2.24552
R25171 DVSS.n5359 DVSS.n3373 2.24552
R25172 DVSS.n7653 DVSS.n7643 2.24552
R25173 DVSS.n7658 DVSS.n2173 2.24552
R25174 DVSS.n7653 DVSS.n7644 2.24552
R25175 DVSS.n7658 DVSS.n2172 2.24552
R25176 DVSS.n7653 DVSS.n7645 2.24552
R25177 DVSS.n7658 DVSS.n2171 2.24552
R25178 DVSS.n7653 DVSS.n7646 2.24552
R25179 DVSS.n7658 DVSS.n2170 2.24552
R25180 DVSS.n7653 DVSS.n7647 2.24552
R25181 DVSS.n7658 DVSS.n2169 2.24552
R25182 DVSS.n7653 DVSS.n7648 2.24552
R25183 DVSS.n7658 DVSS.n2168 2.24552
R25184 DVSS.n7653 DVSS.n7649 2.24552
R25185 DVSS.n7658 DVSS.n2167 2.24552
R25186 DVSS.n7653 DVSS.n7650 2.24552
R25187 DVSS.n7658 DVSS.n2166 2.24552
R25188 DVSS.n7653 DVSS.n7651 2.24552
R25189 DVSS.n7658 DVSS.n2165 2.24552
R25190 DVSS.n7653 DVSS.n7652 2.24552
R25191 DVSS.n7658 DVSS.n2164 2.24552
R25192 DVSS.n7654 DVSS.n7653 2.24552
R25193 DVSS.n7658 DVSS.n2163 2.24552
R25194 DVSS.n7653 DVSS.n2175 2.24552
R25195 DVSS.n8145 DVSS.n8143 2.24552
R25196 DVSS.n8152 DVSS.n1790 2.24552
R25197 DVSS.n8145 DVSS.n8142 2.24552
R25198 DVSS.n8152 DVSS.n1791 2.24552
R25199 DVSS.n8145 DVSS.n8141 2.24552
R25200 DVSS.n8152 DVSS.n1792 2.24552
R25201 DVSS.n8146 DVSS.n8145 2.24552
R25202 DVSS.n8152 DVSS.n1793 2.24552
R25203 DVSS.n8145 DVSS.n1795 2.24552
R25204 DVSS.n8152 DVSS.n8151 2.24552
R25205 DVSS.n1720 DVSS.n1718 2.24552
R25206 DVSS.n1727 DVSS.n1595 2.24552
R25207 DVSS.n1720 DVSS.n1717 2.24552
R25208 DVSS.n1727 DVSS.n1596 2.24552
R25209 DVSS.n1720 DVSS.n1716 2.24552
R25210 DVSS.n1727 DVSS.n1597 2.24552
R25211 DVSS.n1721 DVSS.n1720 2.24552
R25212 DVSS.n1727 DVSS.n1598 2.24552
R25213 DVSS.n1720 DVSS.n1600 2.24552
R25214 DVSS.n1727 DVSS.n1726 2.24552
R25215 DVSS.n2863 DVSS.n2859 2.24552
R25216 DVSS.n710 DVSS.n707 2.24552
R25217 DVSS.n703 DVSS.n700 2.24552
R25218 DVSS.n9374 DVSS.n9371 2.24552
R25219 DVSS.n9539 DVSS.n327 2.24552
R25220 DVSS.n9006 DVSS.n9005 2.24552
R25221 DVSS.n9012 DVSS.n9011 2.24552
R25222 DVSS.n9378 DVSS.n390 2.24552
R25223 DVSS.n9538 DVSS.n325 2.24552
R25224 DVSS.n713 DVSS.n707 2.24552
R25225 DVSS.n706 DVSS.n700 2.24552
R25226 DVSS.n9371 DVSS.n9369 2.24552
R25227 DVSS.n327 DVSS.n324 2.24552
R25228 DVSS.n794 DVSS.n793 2.24552
R25229 DVSS.n804 DVSS.n803 2.24552
R25230 DVSS.n9402 DVSS.n9401 2.24552
R25231 DVSS.n9411 DVSS.n9410 2.24552
R25232 DVSS.n8879 DVSS.n788 2.24552
R25233 DVSS.n8874 DVSS.n798 2.24552
R25234 DVSS.n9397 DVSS.n9396 2.24552
R25235 DVSS.n9406 DVSS.n9405 2.24552
R25236 DVSS.n5941 DVSS.n5933 2.24552
R25237 DVSS.n2890 DVSS.n2888 2.24552
R25238 DVSS.n5941 DVSS.n5932 2.24552
R25239 DVSS.n2890 DVSS.n2889 2.24552
R25240 DVSS.n5941 DVSS.n5931 2.24552
R25241 DVSS.n4922 DVSS.n4921 2.24552
R25242 DVSS.n4926 DVSS.n4923 2.24552
R25243 DVSS.n4922 DVSS.n4920 2.24552
R25244 DVSS.n4926 DVSS.n4924 2.24552
R25245 DVSS.n4922 DVSS.n4919 2.24552
R25246 DVSS.n4926 DVSS.n4925 2.24552
R25247 DVSS.n2928 DVSS.n2922 2.24552
R25248 DVSS.n2933 DVSS.n2923 2.24552
R25249 DVSS.n2934 DVSS.n2922 2.24552
R25250 DVSS.n2936 DVSS.n2923 2.24552
R25251 DVSS.n2937 DVSS.n2922 2.24552
R25252 DVSS.n2939 DVSS.n2923 2.24552
R25253 DVSS.n2959 DVSS.n2940 2.24552
R25254 DVSS.n2950 DVSS.n2941 2.24552
R25255 DVSS.n2959 DVSS.n2958 2.24552
R25256 DVSS.n2952 DVSS.n2941 2.24552
R25257 DVSS.n2959 DVSS.n2957 2.24552
R25258 DVSS.n7689 DVSS.n7679 2.24552
R25259 DVSS.n2135 DVSS.n2119 2.24552
R25260 DVSS.n7689 DVSS.n7680 2.24552
R25261 DVSS.n2137 DVSS.n2119 2.24552
R25262 DVSS.n7689 DVSS.n7681 2.24552
R25263 DVSS.n2139 DVSS.n2119 2.24552
R25264 DVSS.n7689 DVSS.n7682 2.24552
R25265 DVSS.n2141 DVSS.n2119 2.24552
R25266 DVSS.n7689 DVSS.n7683 2.24552
R25267 DVSS.n2143 DVSS.n2119 2.24552
R25268 DVSS.n7689 DVSS.n7684 2.24552
R25269 DVSS.n2145 DVSS.n2119 2.24552
R25270 DVSS.n7689 DVSS.n7685 2.24552
R25271 DVSS.n2147 DVSS.n2119 2.24552
R25272 DVSS.n7689 DVSS.n7686 2.24552
R25273 DVSS.n2149 DVSS.n2119 2.24552
R25274 DVSS.n7689 DVSS.n7687 2.24552
R25275 DVSS.n2151 DVSS.n2119 2.24552
R25276 DVSS.n7689 DVSS.n7688 2.24552
R25277 DVSS.n2153 DVSS.n2119 2.24552
R25278 DVSS.n7690 DVSS.n7689 2.24552
R25279 DVSS.n7691 DVSS.n2119 2.24552
R25280 DVSS.n7689 DVSS.n2118 2.24552
R25281 DVSS.n1771 DVSS.n1762 2.24552
R25282 DVSS.n8174 DVSS.n8171 2.24552
R25283 DVSS.n1773 DVSS.n1762 2.24552
R25284 DVSS.n8174 DVSS.n8172 2.24552
R25285 DVSS.n1775 DVSS.n1762 2.24552
R25286 DVSS.n8174 DVSS.n8173 2.24552
R25287 DVSS.n1777 DVSS.n1762 2.24552
R25288 DVSS.n8175 DVSS.n8174 2.24552
R25289 DVSS.n8176 DVSS.n1762 2.24552
R25290 DVSS.n8174 DVSS.n1761 2.24552
R25291 DVSS.n1746 DVSS.n1562 2.24552
R25292 DVSS.n1572 DVSS.n1563 2.24552
R25293 DVSS.n1746 DVSS.n1584 2.24552
R25294 DVSS.n1574 DVSS.n1563 2.24552
R25295 DVSS.n1746 DVSS.n1583 2.24552
R25296 DVSS.n1576 DVSS.n1563 2.24552
R25297 DVSS.n1746 DVSS.n1582 2.24552
R25298 DVSS.n1578 DVSS.n1563 2.24552
R25299 DVSS.n1746 DVSS.n1581 2.24552
R25300 DVSS.n1580 DVSS.n1563 2.24552
R25301 DVSS.n5930 DVSS.n5929 2.24552
R25302 DVSS.n3249 DVSS.n3247 2.24552
R25303 DVSS.n3240 DVSS.n3238 2.24552
R25304 DVSS.n5396 DVSS.n3323 2.24552
R25305 DVSS.n3316 DVSS.n3314 2.24552
R25306 DVSS.n3310 DVSS.n3308 2.24552
R25307 DVSS.n5679 DVSS.n5678 2.24552
R25308 DVSS.n5686 DVSS.n5685 2.24552
R25309 DVSS.n5496 DVSS.n5495 2.24552
R25310 DVSS.n5503 DVSS.n5502 2.24552
R25311 DVSS.n5509 DVSS.n5508 2.24552
R25312 DVSS.n3253 DVSS.n3247 2.24552
R25313 DVSS.n3244 DVSS.n3238 2.24552
R25314 DVSS.n5400 DVSS.n3323 2.24552
R25315 DVSS.n3320 DVSS.n3314 2.24552
R25316 DVSS.n5511 DVSS.n3310 2.24552
R25317 DVSS.n5679 DVSS.n3252 2.24552
R25318 DVSS.n5686 DVSS.n3243 2.24552
R25319 DVSS.n5496 DVSS.n5399 2.24552
R25320 DVSS.n5503 DVSS.n3319 2.24552
R25321 DVSS.n5510 DVSS.n5509 2.24552
R25322 DVSS.n5656 DVSS.n3264 2.24552
R25323 DVSS.n5646 DVSS.n3271 2.24552
R25324 DVSS.n5539 DVSS.n3295 2.24552
R25325 DVSS.n5529 DVSS.n3303 2.24552
R25326 DVSS.n5520 DVSS.n5518 2.24552
R25327 DVSS.n5664 DVSS.n3260 2.24552
R25328 DVSS.n5654 DVSS.n3267 2.24552
R25329 DVSS.n5547 DVSS.n3290 2.24552
R25330 DVSS.n5537 DVSS.n3298 2.24552
R25331 DVSS.n5528 DVSS.n3305 2.24552
R25332 DVSS.n5658 DVSS.n3264 2.24552
R25333 DVSS.n5648 DVSS.n3271 2.24552
R25334 DVSS.n5541 DVSS.n3295 2.24552
R25335 DVSS.n5531 DVSS.n3303 2.24552
R25336 DVSS.n5522 DVSS.n5518 2.24552
R25337 DVSS.n5664 DVSS.n5663 2.24552
R25338 DVSS.n5654 DVSS.n5653 2.24552
R25339 DVSS.n5547 DVSS.n5546 2.24552
R25340 DVSS.n5537 DVSS.n5536 2.24552
R25341 DVSS.n5528 DVSS.n5527 2.24552
R25342 DVSS.n2669 DVSS.n2668 2.24552
R25343 DVSS.n2662 DVSS.n2661 2.24552
R25344 DVSS.n2654 DVSS.n2653 2.24552
R25345 DVSS.n2715 DVSS.n2714 2.24552
R25346 DVSS.n2724 DVSS.n2723 2.24552
R25347 DVSS.n2732 DVSS.n2731 2.24552
R25348 DVSS.n2676 DVSS.n2675 2.24552
R25349 DVSS.n2682 DVSS.n2681 2.24552
R25350 DVSS.n2689 DVSS.n2688 2.24552
R25351 DVSS.n2749 DVSS.n2709 2.24552
R25352 DVSS.n2743 DVSS.n2718 2.24552
R25353 DVSS.n2738 DVSS.n2726 2.24552
R25354 DVSS.n2673 DVSS.n2668 2.24552
R25355 DVSS.n2666 DVSS.n2661 2.24552
R25356 DVSS.n2658 DVSS.n2653 2.24552
R25357 DVSS.n2714 DVSS.n2711 2.24552
R25358 DVSS.n2723 DVSS.n2720 2.24552
R25359 DVSS.n2731 DVSS.n2728 2.24552
R25360 DVSS.n2676 DVSS.n2672 2.24552
R25361 DVSS.n2682 DVSS.n2665 2.24552
R25362 DVSS.n2689 DVSS.n2657 2.24552
R25363 DVSS.n2749 DVSS.n2748 2.24552
R25364 DVSS.n2743 DVSS.n2742 2.24552
R25365 DVSS.n2738 DVSS.n2737 2.24552
R25366 DVSS.n7353 DVSS.n2596 2.24552
R25367 DVSS.n7344 DVSS.n2603 2.24552
R25368 DVSS.n7334 DVSS.n2611 2.24552
R25369 DVSS.n7727 DVSS.n2088 2.24552
R25370 DVSS.n2097 DVSS.n2096 2.24552
R25371 DVSS.n7710 DVSS.n2104 2.24552
R25372 DVSS.n7361 DVSS.n2591 2.24552
R25373 DVSS.n7352 DVSS.n2598 2.24552
R25374 DVSS.n7342 DVSS.n2606 2.24552
R25375 DVSS.n7855 DVSS.n2083 2.24552
R25376 DVSS.n7725 DVSS.n2091 2.24552
R25377 DVSS.n7718 DVSS.n2099 2.24552
R25378 DVSS.n7355 DVSS.n2596 2.24552
R25379 DVSS.n7346 DVSS.n2603 2.24552
R25380 DVSS.n7336 DVSS.n2611 2.24552
R25381 DVSS.n7849 DVSS.n2088 2.24552
R25382 DVSS.n7719 DVSS.n2096 2.24552
R25383 DVSS.n7712 DVSS.n2104 2.24552
R25384 DVSS.n7361 DVSS.n7360 2.24552
R25385 DVSS.n7352 DVSS.n7351 2.24552
R25386 DVSS.n7342 DVSS.n7341 2.24552
R25387 DVSS.n7855 DVSS.n7854 2.24552
R25388 DVSS.n7725 DVSS.n7724 2.24552
R25389 DVSS.n7718 DVSS.n7717 2.24552
R25390 DVSS.n1903 DVSS.n1900 2.24552
R25391 DVSS.n1894 DVSS.n1891 2.24552
R25392 DVSS.n1884 DVSS.n1881 2.24552
R25393 DVSS.n1858 DVSS.n1855 2.24552
R25394 DVSS.n1836 DVSS.n1835 2.24552
R25395 DVSS.n1843 DVSS.n1842 2.24552
R25396 DVSS.n8072 DVSS.n8071 2.24552
R25397 DVSS.n8078 DVSS.n8077 2.24552
R25398 DVSS.n8085 DVSS.n8084 2.24552
R25399 DVSS.n8107 DVSS.n8106 2.24552
R25400 DVSS.n8114 DVSS.n8113 2.24552
R25401 DVSS.n1851 DVSS.n1838 2.24552
R25402 DVSS.n1907 DVSS.n1900 2.24552
R25403 DVSS.n1898 DVSS.n1891 2.24552
R25404 DVSS.n1888 DVSS.n1881 2.24552
R25405 DVSS.n1862 DVSS.n1855 2.24552
R25406 DVSS.n1853 DVSS.n1835 2.24552
R25407 DVSS.n1845 DVSS.n1842 2.24552
R25408 DVSS.n8072 DVSS.n1906 2.24552
R25409 DVSS.n8078 DVSS.n1897 2.24552
R25410 DVSS.n8085 DVSS.n1887 2.24552
R25411 DVSS.n8107 DVSS.n1861 2.24552
R25412 DVSS.n8114 DVSS.n1834 2.24552
R25413 DVSS.n1851 DVSS.n1850 2.24552
R25414 DVSS.n4490 DVSS.n4488 2.24552
R25415 DVSS.n4492 DVSS.n4456 2.24552
R25416 DVSS.n4490 DVSS.n4486 2.24552
R25417 DVSS.n4492 DVSS.n4457 2.24552
R25418 DVSS.n4490 DVSS.n4483 2.24552
R25419 DVSS.n3856 DVSS.n3836 2.24552
R25420 DVSS.n3846 DVSS.n3837 2.24552
R25421 DVSS.n3856 DVSS.n3855 2.24552
R25422 DVSS.n3848 DVSS.n3837 2.24552
R25423 DVSS.n3856 DVSS.n3854 2.24552
R25424 DVSS.n3850 DVSS.n3837 2.24552
R25425 DVSS.n3033 DVSS.n3027 2.24552
R25426 DVSS.n5856 DVSS.n3028 2.24552
R25427 DVSS.n5857 DVSS.n3027 2.24552
R25428 DVSS.n5859 DVSS.n3028 2.24552
R25429 DVSS.n5860 DVSS.n3027 2.24552
R25430 DVSS.n5862 DVSS.n3028 2.24552
R25431 DVSS.n3004 DVSS.n2994 2.24552
R25432 DVSS.n3006 DVSS.n2995 2.24552
R25433 DVSS.n3007 DVSS.n2994 2.24552
R25434 DVSS.n3009 DVSS.n2995 2.24552
R25435 DVSS.n3010 DVSS.n2994 2.24552
R25436 DVSS.n2544 DVSS.n2530 2.24552
R25437 DVSS.n2545 DVSS.n2526 2.24552
R25438 DVSS.n2547 DVSS.n2530 2.24552
R25439 DVSS.n2548 DVSS.n2526 2.24552
R25440 DVSS.n2550 DVSS.n2530 2.24552
R25441 DVSS.n2551 DVSS.n2526 2.24552
R25442 DVSS.n2553 DVSS.n2530 2.24552
R25443 DVSS.n2554 DVSS.n2526 2.24552
R25444 DVSS.n2556 DVSS.n2530 2.24552
R25445 DVSS.n2557 DVSS.n2526 2.24552
R25446 DVSS.n2559 DVSS.n2530 2.24552
R25447 DVSS.n2560 DVSS.n2526 2.24552
R25448 DVSS.n2562 DVSS.n2530 2.24552
R25449 DVSS.n2563 DVSS.n2526 2.24552
R25450 DVSS.n2565 DVSS.n2530 2.24552
R25451 DVSS.n2566 DVSS.n2526 2.24552
R25452 DVSS.n2568 DVSS.n2530 2.24552
R25453 DVSS.n2569 DVSS.n2526 2.24552
R25454 DVSS.n2571 DVSS.n2530 2.24552
R25455 DVSS.n2572 DVSS.n2526 2.24552
R25456 DVSS.n2574 DVSS.n2530 2.24552
R25457 DVSS.n2575 DVSS.n2526 2.24552
R25458 DVSS.n2577 DVSS.n2530 2.24552
R25459 DVSS.n1926 DVSS.n1917 2.24552
R25460 DVSS.n8056 DVSS.n8053 2.24552
R25461 DVSS.n1928 DVSS.n1917 2.24552
R25462 DVSS.n8056 DVSS.n8054 2.24552
R25463 DVSS.n1930 DVSS.n1917 2.24552
R25464 DVSS.n8056 DVSS.n8055 2.24552
R25465 DVSS.n1932 DVSS.n1917 2.24552
R25466 DVSS.n8057 DVSS.n8056 2.24552
R25467 DVSS.n8058 DVSS.n1917 2.24552
R25468 DVSS.n8056 DVSS.n1916 2.24552
R25469 DVSS.n6754 DVSS.n6736 2.24552
R25470 DVSS.n6854 DVSS.n6851 2.24552
R25471 DVSS.n6756 DVSS.n6736 2.24552
R25472 DVSS.n6854 DVSS.n6852 2.24552
R25473 DVSS.n6758 DVSS.n6736 2.24552
R25474 DVSS.n6854 DVSS.n6853 2.24552
R25475 DVSS.n6760 DVSS.n6736 2.24552
R25476 DVSS.n6855 DVSS.n6854 2.24552
R25477 DVSS.n6856 DVSS.n6736 2.24552
R25478 DVSS.n6854 DVSS.n6735 2.24552
R25479 DVSS.n4458 DVSS.n3834 2.24552
R25480 DVSS.n6910 DVSS.n6887 2.24552
R25481 DVSS.n6906 DVSS.n6904 2.24552
R25482 DVSS.n6913 DVSS.n6862 2.24552
R25483 DVSS.n6906 DVSS.n6903 2.24552
R25484 DVSS.n6913 DVSS.n6863 2.24552
R25485 DVSS.n6906 DVSS.n6902 2.24552
R25486 DVSS.n6913 DVSS.n6864 2.24552
R25487 DVSS.n6906 DVSS.n6901 2.24552
R25488 DVSS.n6913 DVSS.n6865 2.24552
R25489 DVSS.n6906 DVSS.n6900 2.24552
R25490 DVSS.n6913 DVSS.n6866 2.24552
R25491 DVSS.n6906 DVSS.n6899 2.24552
R25492 DVSS.n6913 DVSS.n6867 2.24552
R25493 DVSS.n6906 DVSS.n6898 2.24552
R25494 DVSS.n6913 DVSS.n6868 2.24552
R25495 DVSS.n6906 DVSS.n6897 2.24552
R25496 DVSS.n6913 DVSS.n6869 2.24552
R25497 DVSS.n6906 DVSS.n6896 2.24552
R25498 DVSS.n6913 DVSS.n6870 2.24552
R25499 DVSS.n6907 DVSS.n6906 2.24552
R25500 DVSS.n6913 DVSS.n6871 2.24552
R25501 DVSS.n6906 DVSS.n6873 2.24552
R25502 DVSS.n6913 DVSS.n6912 2.24552
R25503 DVSS.n7055 DVSS.n6690 2.24552
R25504 DVSS.n6705 DVSS.n6691 2.24552
R25505 DVSS.n7055 DVSS.n7046 2.24552
R25506 DVSS.n6707 DVSS.n6691 2.24552
R25507 DVSS.n7055 DVSS.n7047 2.24552
R25508 DVSS.n6709 DVSS.n6691 2.24552
R25509 DVSS.n7055 DVSS.n7048 2.24552
R25510 DVSS.n6711 DVSS.n6691 2.24552
R25511 DVSS.n7055 DVSS.n7049 2.24552
R25512 DVSS.n6713 DVSS.n6691 2.24552
R25513 DVSS.n7055 DVSS.n7050 2.24552
R25514 DVSS.n6715 DVSS.n6691 2.24552
R25515 DVSS.n7055 DVSS.n7051 2.24552
R25516 DVSS.n6717 DVSS.n6691 2.24552
R25517 DVSS.n7055 DVSS.n7052 2.24552
R25518 DVSS.n6719 DVSS.n6691 2.24552
R25519 DVSS.n7055 DVSS.n7053 2.24552
R25520 DVSS.n6721 DVSS.n6691 2.24552
R25521 DVSS.n7055 DVSS.n7054 2.24552
R25522 DVSS.n6723 DVSS.n6691 2.24552
R25523 DVSS.n7056 DVSS.n7055 2.24552
R25524 DVSS.n7057 DVSS.n6691 2.24552
R25525 DVSS.n1311 DVSS.n1189 2.24552
R25526 DVSS.n1204 DVSS.n1191 2.24552
R25527 DVSS.n1311 DVSS.n1304 2.24552
R25528 DVSS.n1206 DVSS.n1190 2.24552
R25529 DVSS.n1311 DVSS.n1305 2.24552
R25530 DVSS.n1208 DVSS.n1190 2.24552
R25531 DVSS.n1311 DVSS.n1306 2.24552
R25532 DVSS.n1210 DVSS.n1190 2.24552
R25533 DVSS.n1311 DVSS.n1307 2.24552
R25534 DVSS.n1212 DVSS.n1190 2.24552
R25535 DVSS.n1311 DVSS.n1308 2.24552
R25536 DVSS.n1298 DVSS.n1190 2.24552
R25537 DVSS.n1311 DVSS.n1309 2.24552
R25538 DVSS.n1300 DVSS.n1190 2.24552
R25539 DVSS.n1311 DVSS.n1310 2.24552
R25540 DVSS.n1302 DVSS.n1190 2.24552
R25541 DVSS.n1312 DVSS.n1311 2.24552
R25542 DVSS.n1313 DVSS.n1190 2.24552
R25543 DVSS.n1078 DVSS.n1077 2.24552
R25544 DVSS.n8534 DVSS.n8533 2.24552
R25545 DVSS.n8543 DVSS.n1078 2.24552
R25546 DVSS.n8561 DVSS.n1070 2.24552
R25547 DVSS.n8545 DVSS.n1078 2.24552
R25548 DVSS.n8561 DVSS.n1069 2.24552
R25549 DVSS.n8547 DVSS.n1078 2.24552
R25550 DVSS.n8561 DVSS.n1068 2.24552
R25551 DVSS.n8549 DVSS.n1078 2.24552
R25552 DVSS.n8561 DVSS.n1067 2.24552
R25553 DVSS.n8551 DVSS.n1078 2.24552
R25554 DVSS.n8561 DVSS.n1065 2.24552
R25555 DVSS.n8553 DVSS.n1078 2.24552
R25556 DVSS.n8561 DVSS.n1064 2.24552
R25557 DVSS.n8555 DVSS.n1078 2.24552
R25558 DVSS.n8561 DVSS.n1063 2.24552
R25559 DVSS.n8557 DVSS.n1078 2.24552
R25560 DVSS.n8561 DVSS.n1062 2.24552
R25561 DVSS.n9658 DVSS.n9635 2.24552
R25562 DVSS.n222 DVSS.n221 2.24552
R25563 DVSS.n9658 DVSS.n9637 2.24552
R25564 DVSS.n9660 DVSS.n213 2.24552
R25565 DVSS.n9658 DVSS.n9640 2.24552
R25566 DVSS.n9660 DVSS.n212 2.24552
R25567 DVSS.n9658 DVSS.n9643 2.24552
R25568 DVSS.n9660 DVSS.n211 2.24552
R25569 DVSS.n9658 DVSS.n9646 2.24552
R25570 DVSS.n9660 DVSS.n210 2.24552
R25571 DVSS.n9658 DVSS.n9648 2.24552
R25572 DVSS.n9660 DVSS.n208 2.24552
R25573 DVSS.n9658 DVSS.n9651 2.24552
R25574 DVSS.n9660 DVSS.n207 2.24552
R25575 DVSS.n9658 DVSS.n9654 2.24552
R25576 DVSS.n9660 DVSS.n206 2.24552
R25577 DVSS.n9658 DVSS.n9657 2.24552
R25578 DVSS.n9660 DVSS.n205 2.24552
R25579 DVSS.n9715 DVSS.n9692 2.24552
R25580 DVSS.n183 DVSS.n182 2.24552
R25581 DVSS.n9715 DVSS.n9694 2.24552
R25582 DVSS.n9717 DVSS.n174 2.24552
R25583 DVSS.n9715 DVSS.n9697 2.24552
R25584 DVSS.n9717 DVSS.n173 2.24552
R25585 DVSS.n9715 DVSS.n9700 2.24552
R25586 DVSS.n9717 DVSS.n172 2.24552
R25587 DVSS.n9715 DVSS.n9703 2.24552
R25588 DVSS.n9717 DVSS.n171 2.24552
R25589 DVSS.n9715 DVSS.n9705 2.24552
R25590 DVSS.n9717 DVSS.n169 2.24552
R25591 DVSS.n9715 DVSS.n9708 2.24552
R25592 DVSS.n9717 DVSS.n168 2.24552
R25593 DVSS.n9715 DVSS.n9711 2.24552
R25594 DVSS.n9717 DVSS.n167 2.24552
R25595 DVSS.n9715 DVSS.n9714 2.24552
R25596 DVSS.n9717 DVSS.n166 2.24552
R25597 DVSS.n9768 DVSS.n9737 2.24552
R25598 DVSS.n9770 DVSS.n154 2.24552
R25599 DVSS.n9768 DVSS.n9740 2.24552
R25600 DVSS.n9770 DVSS.n153 2.24552
R25601 DVSS.n9768 DVSS.n9743 2.24552
R25602 DVSS.n9770 DVSS.n152 2.24552
R25603 DVSS.n9768 DVSS.n9746 2.24552
R25604 DVSS.n9770 DVSS.n151 2.24552
R25605 DVSS.n9768 DVSS.n9749 2.24552
R25606 DVSS.n9770 DVSS.n150 2.24552
R25607 DVSS.n9768 DVSS.n9752 2.24552
R25608 DVSS.n9770 DVSS.n149 2.24552
R25609 DVSS.n9768 DVSS.n9755 2.24552
R25610 DVSS.n9770 DVSS.n148 2.24552
R25611 DVSS.n9768 DVSS.n9758 2.24552
R25612 DVSS.n9770 DVSS.n147 2.24552
R25613 DVSS.n9768 DVSS.n9761 2.24552
R25614 DVSS.n9770 DVSS.n146 2.24552
R25615 DVSS.n9768 DVSS.n9764 2.24552
R25616 DVSS.n9770 DVSS.n145 2.24552
R25617 DVSS.n9768 DVSS.n9767 2.24552
R25618 DVSS.n9770 DVSS.n144 2.24552
R25619 DVSS.n9799 DVSS.n9789 2.24552
R25620 DVSS.n114 DVSS.n98 2.24552
R25621 DVSS.n9799 DVSS.n9790 2.24552
R25622 DVSS.n116 DVSS.n98 2.24552
R25623 DVSS.n9799 DVSS.n9791 2.24552
R25624 DVSS.n118 DVSS.n98 2.24552
R25625 DVSS.n9799 DVSS.n9792 2.24552
R25626 DVSS.n120 DVSS.n98 2.24552
R25627 DVSS.n9799 DVSS.n9793 2.24552
R25628 DVSS.n122 DVSS.n98 2.24552
R25629 DVSS.n9799 DVSS.n9794 2.24552
R25630 DVSS.n124 DVSS.n98 2.24552
R25631 DVSS.n9799 DVSS.n9795 2.24552
R25632 DVSS.n126 DVSS.n98 2.24552
R25633 DVSS.n9799 DVSS.n9796 2.24552
R25634 DVSS.n128 DVSS.n98 2.24552
R25635 DVSS.n9799 DVSS.n9797 2.24552
R25636 DVSS.n130 DVSS.n98 2.24552
R25637 DVSS.n9799 DVSS.n9798 2.24552
R25638 DVSS.n132 DVSS.n98 2.24552
R25639 DVSS.n9800 DVSS.n9799 2.24552
R25640 DVSS.n9801 DVSS.n98 2.24552
R25641 DVSS.n9799 DVSS.n97 2.24552
R25642 DVSS.n8634 DVSS.n8624 2.24552
R25643 DVSS.n993 DVSS.n977 2.24552
R25644 DVSS.n8634 DVSS.n8625 2.24552
R25645 DVSS.n995 DVSS.n977 2.24552
R25646 DVSS.n8634 DVSS.n8626 2.24552
R25647 DVSS.n997 DVSS.n977 2.24552
R25648 DVSS.n8634 DVSS.n8627 2.24552
R25649 DVSS.n999 DVSS.n977 2.24552
R25650 DVSS.n8634 DVSS.n8628 2.24552
R25651 DVSS.n1001 DVSS.n977 2.24552
R25652 DVSS.n8634 DVSS.n8629 2.24552
R25653 DVSS.n1003 DVSS.n977 2.24552
R25654 DVSS.n8634 DVSS.n8630 2.24552
R25655 DVSS.n1005 DVSS.n977 2.24552
R25656 DVSS.n8634 DVSS.n8631 2.24552
R25657 DVSS.n1007 DVSS.n977 2.24552
R25658 DVSS.n8634 DVSS.n8632 2.24552
R25659 DVSS.n1009 DVSS.n977 2.24552
R25660 DVSS.n8634 DVSS.n8633 2.24552
R25661 DVSS.n1011 DVSS.n977 2.24552
R25662 DVSS.n8635 DVSS.n8634 2.24552
R25663 DVSS.n8636 DVSS.n977 2.24552
R25664 DVSS.n8634 DVSS.n976 2.24552
R25665 DVSS.n7028 DVSS.n7027 2.24552
R25666 DVSS.n6967 DVSS.n6966 2.24552
R25667 DVSS.n6979 DVSS.n6969 2.24552
R25668 DVSS.n6967 DVSS.n6965 2.24552
R25669 DVSS.n6979 DVSS.n6970 2.24552
R25670 DVSS.n6967 DVSS.n6964 2.24552
R25671 DVSS.n6979 DVSS.n6971 2.24552
R25672 DVSS.n6967 DVSS.n6963 2.24552
R25673 DVSS.n6979 DVSS.n6972 2.24552
R25674 DVSS.n6967 DVSS.n6962 2.24552
R25675 DVSS.n6979 DVSS.n6973 2.24552
R25676 DVSS.n6967 DVSS.n6961 2.24552
R25677 DVSS.n6979 DVSS.n6974 2.24552
R25678 DVSS.n6967 DVSS.n6960 2.24552
R25679 DVSS.n6979 DVSS.n6975 2.24552
R25680 DVSS.n6967 DVSS.n6959 2.24552
R25681 DVSS.n6979 DVSS.n6976 2.24552
R25682 DVSS.n6967 DVSS.n6958 2.24552
R25683 DVSS.n6979 DVSS.n6977 2.24552
R25684 DVSS.n6967 DVSS.n6957 2.24552
R25685 DVSS.n6979 DVSS.n6978 2.24552
R25686 DVSS.n6967 DVSS.n6956 2.24552
R25687 DVSS.n6979 DVSS.n6955 2.24552
R25688 DVSS.n8856 DVSS.n806 2.24552
R25689 DVSS.n8835 DVSS.n808 2.24552
R25690 DVSS.n8859 DVSS.n812 2.24552
R25691 DVSS.n8837 DVSS.n808 2.24552
R25692 DVSS.n8859 DVSS.n813 2.24552
R25693 DVSS.n8839 DVSS.n808 2.24552
R25694 DVSS.n8859 DVSS.n814 2.24552
R25695 DVSS.n8841 DVSS.n808 2.24552
R25696 DVSS.n8859 DVSS.n815 2.24552
R25697 DVSS.n8843 DVSS.n808 2.24552
R25698 DVSS.n8859 DVSS.n816 2.24552
R25699 DVSS.n8845 DVSS.n808 2.24552
R25700 DVSS.n8859 DVSS.n817 2.24552
R25701 DVSS.n8847 DVSS.n808 2.24552
R25702 DVSS.n8859 DVSS.n818 2.24552
R25703 DVSS.n8849 DVSS.n808 2.24552
R25704 DVSS.n8859 DVSS.n819 2.24552
R25705 DVSS.n8851 DVSS.n808 2.24552
R25706 DVSS.n8859 DVSS.n820 2.24552
R25707 DVSS.n8853 DVSS.n808 2.24552
R25708 DVSS.n8859 DVSS.n821 2.24552
R25709 DVSS.n823 DVSS.n808 2.24552
R25710 DVSS.n8859 DVSS.n8858 2.24552
R25711 DVSS.n422 DVSS.n408 2.24552
R25712 DVSS.n423 DVSS.n407 2.24552
R25713 DVSS.n453 DVSS.n444 2.24552
R25714 DVSS.n425 DVSS.n407 2.24552
R25715 DVSS.n453 DVSS.n445 2.24552
R25716 DVSS.n427 DVSS.n407 2.24552
R25717 DVSS.n453 DVSS.n446 2.24552
R25718 DVSS.n429 DVSS.n407 2.24552
R25719 DVSS.n453 DVSS.n447 2.24552
R25720 DVSS.n431 DVSS.n407 2.24552
R25721 DVSS.n453 DVSS.n448 2.24552
R25722 DVSS.n433 DVSS.n407 2.24552
R25723 DVSS.n453 DVSS.n449 2.24552
R25724 DVSS.n435 DVSS.n407 2.24552
R25725 DVSS.n453 DVSS.n450 2.24552
R25726 DVSS.n437 DVSS.n407 2.24552
R25727 DVSS.n453 DVSS.n451 2.24552
R25728 DVSS.n439 DVSS.n407 2.24552
R25729 DVSS.n453 DVSS.n452 2.24552
R25730 DVSS.n441 DVSS.n407 2.24552
R25731 DVSS.n454 DVSS.n453 2.24552
R25732 DVSS.n455 DVSS.n407 2.24552
R25733 DVSS.n453 DVSS.n406 2.24552
R25734 DVSS.n272 DVSS.n267 2.24552
R25735 DVSS.n9576 DVSS.n9575 2.24552
R25736 DVSS.n9583 DVSS.n274 2.24552
R25737 DVSS.n9576 DVSS.n9574 2.24552
R25738 DVSS.n9583 DVSS.n275 2.24552
R25739 DVSS.n9576 DVSS.n9573 2.24552
R25740 DVSS.n9583 DVSS.n276 2.24552
R25741 DVSS.n9576 DVSS.n9572 2.24552
R25742 DVSS.n9583 DVSS.n277 2.24552
R25743 DVSS.n9576 DVSS.n9571 2.24552
R25744 DVSS.n9583 DVSS.n278 2.24552
R25745 DVSS.n9576 DVSS.n9570 2.24552
R25746 DVSS.n9583 DVSS.n279 2.24552
R25747 DVSS.n9576 DVSS.n9569 2.24552
R25748 DVSS.n9583 DVSS.n280 2.24552
R25749 DVSS.n9576 DVSS.n9568 2.24552
R25750 DVSS.n9583 DVSS.n281 2.24552
R25751 DVSS.n9576 DVSS.n9567 2.24552
R25752 DVSS.n9583 DVSS.n282 2.24552
R25753 DVSS.n9577 DVSS.n9576 2.24552
R25754 DVSS.n9583 DVSS.n283 2.24552
R25755 DVSS.n9576 DVSS.n9547 2.24552
R25756 DVSS.n9583 DVSS.n9582 2.24552
R25757 DVSS.n9839 DVSS.n9828 2.24552
R25758 DVSS.n9806 DVSS.n84 2.24552
R25759 DVSS.n9839 DVSS.n9829 2.24552
R25760 DVSS.n9808 DVSS.n84 2.24552
R25761 DVSS.n9839 DVSS.n9830 2.24552
R25762 DVSS.n9810 DVSS.n84 2.24552
R25763 DVSS.n9839 DVSS.n9831 2.24552
R25764 DVSS.n9812 DVSS.n84 2.24552
R25765 DVSS.n9839 DVSS.n9832 2.24552
R25766 DVSS.n9814 DVSS.n84 2.24552
R25767 DVSS.n9839 DVSS.n9833 2.24552
R25768 DVSS.n9816 DVSS.n84 2.24552
R25769 DVSS.n9839 DVSS.n9834 2.24552
R25770 DVSS.n9818 DVSS.n84 2.24552
R25771 DVSS.n9839 DVSS.n9835 2.24552
R25772 DVSS.n9820 DVSS.n84 2.24552
R25773 DVSS.n9839 DVSS.n9836 2.24552
R25774 DVSS.n9822 DVSS.n84 2.24552
R25775 DVSS.n9839 DVSS.n9837 2.24552
R25776 DVSS.n9824 DVSS.n84 2.24552
R25777 DVSS.n9839 DVSS.n9838 2.24552
R25778 DVSS.n9826 DVSS.n84 2.24552
R25779 DVSS.n9840 DVSS.n9839 2.24552
R25780 DVSS.n8677 DVSS.n8667 2.24552
R25781 DVSS.n8682 DVSS.n975 2.24552
R25782 DVSS.n8677 DVSS.n8668 2.24552
R25783 DVSS.n8682 DVSS.n974 2.24552
R25784 DVSS.n8677 DVSS.n8669 2.24552
R25785 DVSS.n8682 DVSS.n973 2.24552
R25786 DVSS.n8677 DVSS.n8670 2.24552
R25787 DVSS.n8682 DVSS.n972 2.24552
R25788 DVSS.n8677 DVSS.n8671 2.24552
R25789 DVSS.n8682 DVSS.n971 2.24552
R25790 DVSS.n8677 DVSS.n8672 2.24552
R25791 DVSS.n8682 DVSS.n970 2.24552
R25792 DVSS.n8677 DVSS.n8673 2.24552
R25793 DVSS.n8682 DVSS.n969 2.24552
R25794 DVSS.n8677 DVSS.n8674 2.24552
R25795 DVSS.n8682 DVSS.n968 2.24552
R25796 DVSS.n8677 DVSS.n8675 2.24552
R25797 DVSS.n8682 DVSS.n967 2.24552
R25798 DVSS.n8677 DVSS.n8676 2.24552
R25799 DVSS.n8682 DVSS.n966 2.24552
R25800 DVSS.n8678 DVSS.n8677 2.24552
R25801 DVSS.n8682 DVSS.n965 2.24552
R25802 DVSS.n8677 DVSS.n8641 2.24552
R25803 DVSS.n917 DVSS.n902 2.24552
R25804 DVSS.n918 DVSS.n898 2.24552
R25805 DVSS.n920 DVSS.n902 2.24552
R25806 DVSS.n921 DVSS.n898 2.24552
R25807 DVSS.n923 DVSS.n902 2.24552
R25808 DVSS.n924 DVSS.n898 2.24552
R25809 DVSS.n926 DVSS.n902 2.24552
R25810 DVSS.n927 DVSS.n898 2.24552
R25811 DVSS.n929 DVSS.n902 2.24552
R25812 DVSS.n930 DVSS.n898 2.24552
R25813 DVSS.n932 DVSS.n902 2.24552
R25814 DVSS.n933 DVSS.n898 2.24552
R25815 DVSS.n935 DVSS.n902 2.24552
R25816 DVSS.n936 DVSS.n898 2.24552
R25817 DVSS.n938 DVSS.n902 2.24552
R25818 DVSS.n939 DVSS.n898 2.24552
R25819 DVSS.n941 DVSS.n902 2.24552
R25820 DVSS.n942 DVSS.n898 2.24552
R25821 DVSS.n944 DVSS.n902 2.24552
R25822 DVSS.n945 DVSS.n898 2.24552
R25823 DVSS.n947 DVSS.n902 2.24552
R25824 DVSS.n948 DVSS.n898 2.24552
R25825 DVSS.n903 DVSS.n902 2.24552
R25826 DVSS.n854 DVSS.n839 2.24552
R25827 DVSS.n855 DVSS.n835 2.24552
R25828 DVSS.n857 DVSS.n839 2.24552
R25829 DVSS.n858 DVSS.n835 2.24552
R25830 DVSS.n860 DVSS.n839 2.24552
R25831 DVSS.n861 DVSS.n835 2.24552
R25832 DVSS.n863 DVSS.n839 2.24552
R25833 DVSS.n864 DVSS.n835 2.24552
R25834 DVSS.n866 DVSS.n839 2.24552
R25835 DVSS.n867 DVSS.n835 2.24552
R25836 DVSS.n869 DVSS.n839 2.24552
R25837 DVSS.n870 DVSS.n835 2.24552
R25838 DVSS.n872 DVSS.n839 2.24552
R25839 DVSS.n873 DVSS.n835 2.24552
R25840 DVSS.n875 DVSS.n839 2.24552
R25841 DVSS.n876 DVSS.n835 2.24552
R25842 DVSS.n878 DVSS.n839 2.24552
R25843 DVSS.n879 DVSS.n835 2.24552
R25844 DVSS.n881 DVSS.n839 2.24552
R25845 DVSS.n882 DVSS.n835 2.24552
R25846 DVSS.n884 DVSS.n839 2.24552
R25847 DVSS.n885 DVSS.n835 2.24552
R25848 DVSS.n840 DVSS.n839 2.24552
R25849 DVSS.n9363 DVSS.n9353 2.24552
R25850 DVSS.n461 DVSS.n392 2.24552
R25851 DVSS.n9363 DVSS.n9354 2.24552
R25852 DVSS.n463 DVSS.n392 2.24552
R25853 DVSS.n9363 DVSS.n9355 2.24552
R25854 DVSS.n465 DVSS.n392 2.24552
R25855 DVSS.n9363 DVSS.n9356 2.24552
R25856 DVSS.n467 DVSS.n392 2.24552
R25857 DVSS.n9363 DVSS.n9357 2.24552
R25858 DVSS.n469 DVSS.n392 2.24552
R25859 DVSS.n9363 DVSS.n9358 2.24552
R25860 DVSS.n471 DVSS.n392 2.24552
R25861 DVSS.n9363 DVSS.n9359 2.24552
R25862 DVSS.n473 DVSS.n392 2.24552
R25863 DVSS.n9363 DVSS.n9360 2.24552
R25864 DVSS.n475 DVSS.n392 2.24552
R25865 DVSS.n9363 DVSS.n9361 2.24552
R25866 DVSS.n477 DVSS.n392 2.24552
R25867 DVSS.n9363 DVSS.n9362 2.24552
R25868 DVSS.n479 DVSS.n392 2.24552
R25869 DVSS.n9364 DVSS.n9363 2.24552
R25870 DVSS.n9365 DVSS.n392 2.24552
R25871 DVSS.n9363 DVSS.n391 2.24552
R25872 DVSS.n9324 DVSS.n284 2.24552
R25873 DVSS.n301 DVSS.n285 2.24552
R25874 DVSS.n9324 DVSS.n9314 2.24552
R25875 DVSS.n303 DVSS.n285 2.24552
R25876 DVSS.n9324 DVSS.n9315 2.24552
R25877 DVSS.n305 DVSS.n285 2.24552
R25878 DVSS.n9324 DVSS.n9316 2.24552
R25879 DVSS.n307 DVSS.n285 2.24552
R25880 DVSS.n9324 DVSS.n9317 2.24552
R25881 DVSS.n309 DVSS.n285 2.24552
R25882 DVSS.n9324 DVSS.n9318 2.24552
R25883 DVSS.n311 DVSS.n285 2.24552
R25884 DVSS.n9324 DVSS.n9319 2.24552
R25885 DVSS.n313 DVSS.n285 2.24552
R25886 DVSS.n9324 DVSS.n9320 2.24552
R25887 DVSS.n315 DVSS.n285 2.24552
R25888 DVSS.n9324 DVSS.n9321 2.24552
R25889 DVSS.n317 DVSS.n285 2.24552
R25890 DVSS.n9324 DVSS.n9322 2.24552
R25891 DVSS.n319 DVSS.n285 2.24552
R25892 DVSS.n9324 DVSS.n9323 2.24552
R25893 DVSS.n321 DVSS.n285 2.24552
R25894 DVSS.n9324 DVSS.n323 2.24552
R25895 DVSS.n9929 DVSS.n9919 2.24552
R25896 DVSS.n9934 DVSS.n16 2.24552
R25897 DVSS.n9929 DVSS.n9920 2.24552
R25898 DVSS.n9934 DVSS.n15 2.24552
R25899 DVSS.n9929 DVSS.n9921 2.24552
R25900 DVSS.n9934 DVSS.n14 2.24552
R25901 DVSS.n9929 DVSS.n9922 2.24552
R25902 DVSS.n9934 DVSS.n13 2.24552
R25903 DVSS.n9929 DVSS.n9923 2.24552
R25904 DVSS.n9934 DVSS.n12 2.24552
R25905 DVSS.n9929 DVSS.n9924 2.24552
R25906 DVSS.n9934 DVSS.n11 2.24552
R25907 DVSS.n9929 DVSS.n9925 2.24552
R25908 DVSS.n9934 DVSS.n10 2.24552
R25909 DVSS.n9929 DVSS.n9926 2.24552
R25910 DVSS.n9934 DVSS.n9 2.24552
R25911 DVSS.n9929 DVSS.n9927 2.24552
R25912 DVSS.n9934 DVSS.n8 2.24552
R25913 DVSS.n9929 DVSS.n9928 2.24552
R25914 DVSS.n9934 DVSS.n7 2.24552
R25915 DVSS.n9930 DVSS.n9929 2.24552
R25916 DVSS.n9934 DVSS.n6 2.24552
R25917 DVSS.n9929 DVSS.n18 2.24552
R25918 DVSS.n7091 DVSS.n7089 2.24531
R25919 DVSS.n8259 DVSS.n1505 2.24531
R25920 DVSS.n8275 DVSS.n8274 2.24531
R25921 DVSS.n1503 DVSS.n1500 2.24531
R25922 DVSS.n8284 DVSS.n8283 2.24531
R25923 DVSS.n1468 DVSS.n1466 2.24531
R25924 DVSS.n8302 DVSS.n1470 2.24531
R25925 DVSS.n1527 DVSS.n1525 2.24531
R25926 DVSS.n1521 DVSS.n1519 2.24531
R25927 DVSS.n1496 DVSS.n1493 2.24531
R25928 DVSS.n1508 DVSS.n1506 2.24531
R25929 DVSS.n8226 DVSS.n8225 2.24531
R25930 DVSS.n8231 DVSS.n8230 2.24531
R25931 DVSS.n8250 DVSS.n1510 2.24531
R25932 DVSS.n8290 DVSS.n8289 2.24531
R25933 DVSS.n7082 DVSS.n7080 2.24531
R25934 DVSS.n8469 DVSS.n1144 2.24531
R25935 DVSS.n1380 DVSS.n1378 2.24531
R25936 DVSS.n8472 DVSS.n8471 2.24531
R25937 DVSS.n1385 DVSS.n1384 2.24531
R25938 DVSS.n1266 DVSS.n1241 2.24531
R25939 DVSS.n1275 DVSS.n1237 2.24531
R25940 DVSS.n8384 DVSS.n1416 2.24531
R25941 DVSS.n8375 DVSS.n8359 2.24531
R25942 DVSS.n7100 DVSS.n7099 2.24531
R25943 DVSS.n7087 DVSS.n7085 2.24531
R25944 DVSS.n7245 DVSS.n7242 2.24531
R25945 DVSS.n7250 DVSS.n7249 2.24531
R25946 DVSS.n9007 DVSS.n709 2.24505
R25947 DVSS.n9013 DVSS.n702 2.24505
R25948 DVSS.n9373 DVSS.n389 2.24505
R25949 DVSS.n330 DVSS.n329 2.24505
R25950 DVSS.n796 DVSS.n787 2.24505
R25951 DVSS.n8861 DVSS.n797 2.24505
R25952 DVSS.n9398 DVSS.n369 2.24505
R25953 DVSS.n9407 DVSS.n367 2.24505
R25954 DVSS.n795 DVSS.n792 2.24505
R25955 DVSS.n805 DVSS.n802 2.24505
R25956 DVSS.n8864 DVSS.n606 2.24505
R25957 DVSS.n9390 DVSS.n371 2.24505
R25958 DVSS.n9400 DVSS.n224 2.24505
R25959 DVSS.n9409 DVSS.n185 2.24505
R25960 DVSS.n8878 DVSS.n790 2.24505
R25961 DVSS.n8873 DVSS.n800 2.24505
R25962 DVSS.n8863 DVSS.n603 2.24505
R25963 DVSS.n9394 DVSS.n9393 2.24505
R25964 DVSS.n9403 DVSS.n220 2.24505
R25965 DVSS.n9412 DVSS.n181 2.24505
R25966 DVSS.n8277 DVSS.n8276 2.24456
R25967 DVSS.n8260 DVSS.n1471 2.24456
R25968 DVSS.n8262 DVSS.n1465 2.24456
R25969 DVSS.n8280 DVSS.n1498 2.24456
R25970 DVSS.n8323 DVSS.n1449 2.24456
R25971 DVSS.n8303 DVSS.n1467 2.24456
R25972 DVSS.n8309 DVSS.n1461 2.24456
R25973 DVSS.n1497 DVSS.n1491 2.24456
R25974 DVSS.n8251 DVSS.n1507 2.24456
R25975 DVSS.n8224 DVSS.n1517 2.24456
R25976 DVSS.n1490 DVSS.n1481 2.24456
R25977 DVSS.n8244 DVSS.n8239 2.24456
R25978 DVSS.n8233 DVSS.n1516 2.24456
R25979 DVSS.n8443 DVSS.n8442 2.24456
R25980 DVSS.n8442 DVSS.n8441 2.24456
R25981 DVSS.n1387 DVSS.n1386 2.24456
R25982 DVSS.n8474 DVSS.n8473 2.24456
R25983 DVSS.n8479 DVSS.n1137 2.24456
R25984 DVSS.n8487 DVSS.n1127 2.24456
R25985 DVSS.n8445 DVSS.n8444 2.24456
R25986 DVSS.n1282 DVSS.n1228 2.24456
R25987 DVSS.n1276 DVSS.n1235 2.24456
R25988 DVSS.n1267 DVSS.n1239 2.24456
R25989 DVSS.n1262 DVSS.n1243 2.24456
R25990 DVSS.n1257 DVSS.n1250 2.24456
R25991 DVSS.n1253 DVSS.n1249 2.24456
R25992 DVSS.n1246 DVSS.n1242 2.24456
R25993 DVSS.n1231 DVSS.n1227 2.24456
R25994 DVSS.n8369 DVSS.n8362 2.24456
R25995 DVSS.n8365 DVSS.n8362 2.24456
R25996 DVSS.n8374 DVSS.n8358 2.24456
R25997 DVSS.n8383 DVSS.n1405 2.24456
R25998 DVSS.n8350 DVSS.n1418 2.24456
R25999 DVSS.n8351 DVSS.n8350 2.24456
R26000 DVSS.n8493 DVSS.n1098 2.24456
R26001 DVSS.n1102 DVSS.n1098 2.24456
R26002 DVSS.n8491 DVSS.n1097 2.24456
R26003 DVSS.n1420 DVSS.n1417 2.24456
R26004 DVSS.n8382 DVSS.n8381 2.24456
R26005 DVSS.n8373 DVSS.n8357 2.24456
R26006 DVSS.n8367 DVSS.n8361 2.24456
R26007 DVSS.n8454 DVSS.n1153 2.24456
R26008 DVSS.n8455 DVSS.n8454 2.24456
R26009 DVSS.n1157 DVSS.n1152 2.24456
R26010 DVSS.n8450 DVSS.n1182 2.24456
R26011 DVSS.n1287 DVSS.n1221 2.24456
R26012 DVSS.n1224 DVSS.n1220 2.24456
R26013 DVSS.n8279 DVSS.n1504 2.24456
R26014 DVSS.n8272 DVSS.n8267 2.24456
R26015 DVSS.n1502 DVSS.n1499 2.24456
R26016 DVSS.n8328 DVSS.n1447 2.24456
R26017 DVSS.n8306 DVSS.n8305 2.24456
R26018 DVSS.n8313 DVSS.n8312 2.24456
R26019 DVSS.n8227 DVSS.n1518 2.24456
R26020 DVSS.n8254 DVSS.n8253 2.24456
R26021 DVSS.n1495 DVSS.n1492 2.24456
R26022 DVSS.n8238 DVSS.n1514 2.24456
R26023 DVSS.n8248 DVSS.n8247 2.24456
R26024 DVSS.n8292 DVSS.n1485 2.24456
R26025 DVSS.n8481 DVSS.n1130 2.24456
R26026 DVSS.n8477 DVSS.n1133 2.24456
R26027 DVSS.n8470 DVSS.n1141 2.24456
R26028 DVSS.n1382 DVSS.n1381 2.24456
R26029 DVSS.n1259 DVSS.n1252 2.24456
R26030 DVSS.n1264 DVSS.n1245 2.24456
R26031 DVSS.n1270 DVSS.n1269 2.24456
R26032 DVSS.n1279 DVSS.n1278 2.24456
R26033 DVSS.n1284 DVSS.n1230 2.24456
R26034 DVSS.n1317 DVSS.n1185 2.24456
R26035 DVSS.n1289 DVSS.n1223 2.24456
R26036 DVSS.n4815 DVSS.n3677 2.24447
R26037 DVSS.n5237 DVSS.n3477 2.24447
R26038 DVSS.n5194 DVSS.n5009 2.24447
R26039 DVSS.n8388 DVSS.n1413 2.24447
R26040 DVSS.n8392 DVSS.n1403 2.24447
R26041 DVSS.n8390 DVSS.n8388 2.24447
R26042 DVSS.n8392 DVSS.n1402 2.24447
R26043 DVSS.n8388 DVSS.n1410 2.24447
R26044 DVSS.n8392 DVSS.n1400 2.24447
R26045 DVSS.n8388 DVSS.n1407 2.24447
R26046 DVSS.n8392 DVSS.n1399 2.24447
R26047 DVSS.n3703 DVSS.n3689 2.24447
R26048 DVSS.n4105 DVSS.n3973 2.24447
R26049 DVSS.n3184 DVSS.n3175 2.24447
R26050 DVSS.n8400 DVSS.n1391 2.24447
R26051 DVSS.n1377 DVSS.n1376 2.24447
R26052 DVSS.n8400 DVSS.n1390 2.24447
R26053 DVSS.n1377 DVSS.n1375 2.24447
R26054 DVSS.n8400 DVSS.n1389 2.24447
R26055 DVSS.n1377 DVSS.n1374 2.24447
R26056 DVSS.n8401 DVSS.n8400 2.24447
R26057 DVSS.n1377 DVSS.n1373 2.24447
R26058 DVSS.n2334 DVSS.n2310 2.24447
R26059 DVSS.n2304 DVSS.n2280 2.24447
R26060 DVSS.n3783 DVSS.n3781 2.24447
R26061 DVSS.n3783 DVSS.n3782 2.24447
R26062 DVSS.n4749 DVSS.n4619 2.24447
R26063 DVSS.n4749 DVSS.n4748 2.24447
R26064 DVSS.n9020 DVSS.n9018 2.24447
R26065 DVSS.n9379 DVSS.n384 2.24447
R26066 DVSS.n9023 DVSS.n9022 2.24447
R26067 DVSS.n9383 DVSS.n385 2.24447
R26068 DVSS.n9018 DVSS.n699 2.24447
R26069 DVSS.n387 DVSS.n384 2.24447
R26070 DVSS.n8866 DVSS.n8865 2.24447
R26071 DVSS.n377 DVSS.n376 2.24447
R26072 DVSS.n8869 DVSS.n8868 2.24447
R26073 DVSS.n9392 DVSS.n9391 2.24447
R26074 DVSS.n3235 DVSS.n3232 2.24447
R26075 DVSS.n5405 DVSS.n5402 2.24447
R26076 DVSS.n5692 DVSS.n5691 2.24447
R26077 DVSS.n5492 DVSS.n5491 2.24447
R26078 DVSS.n3237 DVSS.n3232 2.24447
R26079 DVSS.n5486 DVSS.n5402 2.24447
R26080 DVSS.n5695 DVSS.n5694 2.24447
R26081 DVSS.n5494 DVSS.n5403 2.24447
R26082 DVSS.n3278 DVSS.n3277 2.24447
R26083 DVSS.n5548 DVSS.n3288 2.24447
R26084 DVSS.n5645 DVSS.n3274 2.24447
R26085 DVSS.n5634 DVSS.n5633 2.24447
R26086 DVSS.n3277 DVSS.n3276 2.24447
R26087 DVSS.n5632 DVSS.n3288 2.24447
R26088 DVSS.n5643 DVSS.n3281 2.24447
R26089 DVSS.n5637 DVSS.n5636 2.24447
R26090 DVSS.n2696 DVSS.n2652 2.24447
R26091 DVSS.n2707 DVSS.n2706 2.24447
R26092 DVSS.n7268 DVSS.n2694 2.24447
R26093 DVSS.n2754 DVSS.n2703 2.24447
R26094 DVSS.n7267 DVSS.n2696 2.24447
R26095 DVSS.n2706 DVSS.n2705 2.24447
R26096 DVSS.n7270 DVSS.n2697 2.24447
R26097 DVSS.n2752 DVSS.n2751 2.24447
R26098 DVSS.n2618 DVSS.n2617 2.24447
R26099 DVSS.n2080 DVSS.n2078 2.24447
R26100 DVSS.n7333 DVSS.n2614 2.24447
R26101 DVSS.n7858 DVSS.n2079 2.24447
R26102 DVSS.n2617 DVSS.n2616 2.24447
R26103 DVSS.n7857 DVSS.n2080 2.24447
R26104 DVSS.n7331 DVSS.n2621 2.24447
R26105 DVSS.n7860 DVSS.n2081 2.24447
R26106 DVSS.n1878 DVSS.n1876 2.24447
R26107 DVSS.n1867 DVSS.n1864 2.24447
R26108 DVSS.n8091 DVSS.n8090 2.24447
R26109 DVSS.n8103 DVSS.n8102 2.24447
R26110 DVSS.n1880 DVSS.n1876 2.24447
R26111 DVSS.n1869 DVSS.n1864 2.24447
R26112 DVSS.n8094 DVSS.n8093 2.24447
R26113 DVSS.n8105 DVSS.n1865 2.24447
R26114 DVSS.n605 DVSS.n604 2.24447
R26115 DVSS.n9130 DVSS.n593 2.24447
R26116 DVSS.n615 DVSS.n605 2.24447
R26117 DVSS.n9130 DVSS.n592 2.24447
R26118 DVSS.n9112 DVSS.n605 2.24447
R26119 DVSS.n9130 DVSS.n591 2.24447
R26120 DVSS.n9114 DVSS.n605 2.24447
R26121 DVSS.n9130 DVSS.n590 2.24447
R26122 DVSS.n9116 DVSS.n605 2.24447
R26123 DVSS.n9118 DVSS.n605 2.24447
R26124 DVSS.n9130 DVSS.n599 2.24447
R26125 DVSS.n9120 DVSS.n605 2.24447
R26126 DVSS.n9130 DVSS.n600 2.24447
R26127 DVSS.n9122 DVSS.n605 2.24447
R26128 DVSS.n9130 DVSS.n601 2.24447
R26129 DVSS.n9124 DVSS.n605 2.24447
R26130 DVSS.n9130 DVSS.n602 2.24447
R26131 DVSS.n9126 DVSS.n605 2.24447
R26132 DVSS.n9153 DVSS.n9150 2.24447
R26133 DVSS.n9159 DVSS.n565 2.24447
R26134 DVSS.n9153 DVSS.n9149 2.24447
R26135 DVSS.n9159 DVSS.n564 2.24447
R26136 DVSS.n9153 DVSS.n9148 2.24447
R26137 DVSS.n9159 DVSS.n563 2.24447
R26138 DVSS.n9153 DVSS.n9147 2.24447
R26139 DVSS.n9159 DVSS.n562 2.24447
R26140 DVSS.n9153 DVSS.n9146 2.24447
R26141 DVSS.n9153 DVSS.n9145 2.24447
R26142 DVSS.n9159 DVSS.n571 2.24447
R26143 DVSS.n9153 DVSS.n9151 2.24447
R26144 DVSS.n9159 DVSS.n572 2.24447
R26145 DVSS.n9153 DVSS.n9152 2.24447
R26146 DVSS.n9159 DVSS.n573 2.24447
R26147 DVSS.n9154 DVSS.n9153 2.24447
R26148 DVSS.n9159 DVSS.n9158 2.24447
R26149 DVSS.n9153 DVSS.n574 2.24447
R26150 DVSS.n9065 DVSS.n649 2.24447
R26151 DVSS.n9060 DVSS.n9050 2.24447
R26152 DVSS.n9065 DVSS.n650 2.24447
R26153 DVSS.n9060 DVSS.n9051 2.24447
R26154 DVSS.n9065 DVSS.n651 2.24447
R26155 DVSS.n9060 DVSS.n9052 2.24447
R26156 DVSS.n9065 DVSS.n652 2.24447
R26157 DVSS.n9060 DVSS.n9053 2.24447
R26158 DVSS.n9065 DVSS.n653 2.24447
R26159 DVSS.n9060 DVSS.n9054 2.24447
R26160 DVSS.n9065 DVSS.n654 2.24447
R26161 DVSS.n9060 DVSS.n9055 2.24447
R26162 DVSS.n9065 DVSS.n655 2.24447
R26163 DVSS.n9060 DVSS.n9056 2.24447
R26164 DVSS.n9065 DVSS.n656 2.24447
R26165 DVSS.n9060 DVSS.n9057 2.24447
R26166 DVSS.n9065 DVSS.n657 2.24447
R26167 DVSS.n9060 DVSS.n9058 2.24447
R26168 DVSS.n9065 DVSS.n658 2.24447
R26169 DVSS.n9060 DVSS.n9059 2.24447
R26170 DVSS.n9065 DVSS.n659 2.24447
R26171 DVSS.n9061 DVSS.n9060 2.24447
R26172 DVSS.n9060 DVSS.n660 2.24447
R26173 DVSS.n517 DVSS.n502 2.24447
R26174 DVSS.n9208 DVSS.n9198 2.24447
R26175 DVSS.n519 DVSS.n502 2.24447
R26176 DVSS.n9208 DVSS.n9199 2.24447
R26177 DVSS.n521 DVSS.n502 2.24447
R26178 DVSS.n9208 DVSS.n9200 2.24447
R26179 DVSS.n523 DVSS.n502 2.24447
R26180 DVSS.n9208 DVSS.n9201 2.24447
R26181 DVSS.n525 DVSS.n502 2.24447
R26182 DVSS.n9208 DVSS.n9202 2.24447
R26183 DVSS.n527 DVSS.n502 2.24447
R26184 DVSS.n9208 DVSS.n9203 2.24447
R26185 DVSS.n529 DVSS.n502 2.24447
R26186 DVSS.n9208 DVSS.n9204 2.24447
R26187 DVSS.n531 DVSS.n502 2.24447
R26188 DVSS.n9208 DVSS.n9205 2.24447
R26189 DVSS.n533 DVSS.n502 2.24447
R26190 DVSS.n9208 DVSS.n9206 2.24447
R26191 DVSS.n535 DVSS.n502 2.24447
R26192 DVSS.n9208 DVSS.n9207 2.24447
R26193 DVSS.n9210 DVSS.n502 2.24447
R26194 DVSS.n9209 DVSS.n9208 2.24447
R26195 DVSS.n9208 DVSS.n501 2.24447
R26196 DVSS.n676 DVSS.n662 2.24447
R26197 DVSS.n8788 DVSS.n661 2.24447
R26198 DVSS.n678 DVSS.n662 2.24447
R26199 DVSS.n8788 DVSS.n8778 2.24447
R26200 DVSS.n680 DVSS.n662 2.24447
R26201 DVSS.n8788 DVSS.n8779 2.24447
R26202 DVSS.n682 DVSS.n662 2.24447
R26203 DVSS.n8788 DVSS.n8780 2.24447
R26204 DVSS.n684 DVSS.n662 2.24447
R26205 DVSS.n8788 DVSS.n8781 2.24447
R26206 DVSS.n686 DVSS.n662 2.24447
R26207 DVSS.n8788 DVSS.n8782 2.24447
R26208 DVSS.n688 DVSS.n662 2.24447
R26209 DVSS.n8788 DVSS.n8783 2.24447
R26210 DVSS.n690 DVSS.n662 2.24447
R26211 DVSS.n8788 DVSS.n8784 2.24447
R26212 DVSS.n692 DVSS.n662 2.24447
R26213 DVSS.n8788 DVSS.n8785 2.24447
R26214 DVSS.n694 DVSS.n662 2.24447
R26215 DVSS.n8788 DVSS.n8786 2.24447
R26216 DVSS.n696 DVSS.n662 2.24447
R26217 DVSS.n8788 DVSS.n8787 2.24447
R26218 DVSS.n8788 DVSS.n698 2.24447
R26219 DVSS.n9217 DVSS.n495 2.24447
R26220 DVSS.n9260 DVSS.n9215 2.24447
R26221 DVSS.n9221 DVSS.n495 2.24447
R26222 DVSS.n9260 DVSS.n9219 2.24447
R26223 DVSS.n9225 DVSS.n495 2.24447
R26224 DVSS.n9260 DVSS.n9223 2.24447
R26225 DVSS.n9229 DVSS.n495 2.24447
R26226 DVSS.n9260 DVSS.n9227 2.24447
R26227 DVSS.n9233 DVSS.n495 2.24447
R26228 DVSS.n9260 DVSS.n9231 2.24447
R26229 DVSS.n9237 DVSS.n495 2.24447
R26230 DVSS.n9260 DVSS.n9235 2.24447
R26231 DVSS.n9241 DVSS.n495 2.24447
R26232 DVSS.n9260 DVSS.n9239 2.24447
R26233 DVSS.n9245 DVSS.n495 2.24447
R26234 DVSS.n9260 DVSS.n9243 2.24447
R26235 DVSS.n9249 DVSS.n495 2.24447
R26236 DVSS.n9260 DVSS.n9247 2.24447
R26237 DVSS.n9253 DVSS.n495 2.24447
R26238 DVSS.n9260 DVSS.n9251 2.24447
R26239 DVSS.n9257 DVSS.n495 2.24447
R26240 DVSS.n9260 DVSS.n9255 2.24447
R26241 DVSS.n9260 DVSS.n9259 2.24447
R26242 DVSS.n7252 DVSS.n7251 2.24423
R26243 DVSS.n7136 DVSS.n6650 2.24423
R26244 DVSS.n7151 DVSS.n6649 2.24423
R26245 DVSS.n1538 DVSS.n1535 2.24423
R26246 DVSS.n8211 DVSS.n1532 2.24423
R26247 DVSS.n7241 DVSS.n6645 2.24423
R26248 DVSS.n8201 DVSS.n1540 2.24423
R26249 DVSS.n8194 DVSS.n1554 2.24423
R26250 DVSS.n8198 DVSS.n1558 2.24423
R26251 DVSS.n8205 DVSS.n1551 2.24423
R26252 DVSS.n1751 DVSS.n1561 2.24423
R26253 DVSS.n8189 DVSS.n8188 2.24423
R26254 DVSS.n4472 DVSS.n4471 2.24423
R26255 DVSS.n4471 DVSS.n4467 2.24423
R26256 DVSS.n3797 DVSS.n3792 2.24423
R26257 DVSS.n4592 DVSS.n3792 2.24423
R26258 DVSS.n4598 DVSS.n4597 2.24423
R26259 DVSS.n4598 DVSS.n3787 2.24423
R26260 DVSS.n4603 DVSS.n4602 2.24423
R26261 DVSS.n2765 DVSS.n2761 2.24423
R26262 DVSS.n6005 DVSS.n2769 2.24423
R26263 DVSS.n6005 DVSS.n2779 2.24423
R26264 DVSS.n2905 DVSS.n2904 2.24423
R26265 DVSS.n2905 DVSS.n2900 2.24423
R26266 DVSS.n2909 DVSS.n2908 2.24423
R26267 DVSS.n2909 DVSS.n2894 2.24423
R26268 DVSS.n4465 DVSS.n3826 2.24423
R26269 DVSS.n4469 DVSS.n3826 2.24423
R26270 DVSS.n4591 DVSS.n4590 2.24423
R26271 DVSS.n4590 DVSS.n3791 2.24423
R26272 DVSS.n3789 DVSS.n3744 2.24423
R26273 DVSS.n3785 DVSS.n3744 2.24423
R26274 DVSS.n4606 DVSS.n4605 2.24423
R26275 DVSS.n4606 DVSS.n3784 2.24423
R26276 DVSS.n4620 DVSS.n2760 2.24423
R26277 DVSS.n4620 DVSS.n2767 2.24423
R26278 DVSS.n2774 DVSS.n2768 2.24423
R26279 DVSS.n2776 DVSS.n2768 2.24423
R26280 DVSS.n2902 DVSS.n2831 2.24423
R26281 DVSS.n2898 DVSS.n2831 2.24423
R26282 DVSS.n2896 DVSS.n2864 2.24423
R26283 DVSS.n2892 DVSS.n2864 2.24423
R26284 DVSS.n5928 DVSS.n2891 2.24423
R26285 DVSS.n5926 DVSS.n2887 2.24423
R26286 DVSS.n6663 DVSS.n6659 2.24423
R26287 DVSS.n7069 DVSS.n6655 2.24423
R26288 DVSS.n7130 DVSS.n6654 2.24423
R26289 DVSS.n7064 DVSS.n6658 2.24423
R26290 DVSS.n6751 DVSS.n6745 2.24423
R26291 DVSS.n4476 DVSS.n4475 2.24423
R26292 DVSS.n4478 DVSS.n4462 2.24423
R26293 DVSS.n6753 DVSS.n6748 2.24423
R26294 DVSS.n8333 DVSS.n1442 2.24011
R26295 DVSS.n7097 DVSS.n7090 2.24011
R26296 DVSS.n8216 DVSS.n8215 2.24011
R26297 DVSS.n8223 DVSS.n1520 2.24011
R26298 DVSS.n8507 DVSS.n1087 2.24011
R26299 DVSS.n8507 DVSS.n8506 2.24011
R26300 DVSS.n8513 DVSS.n1085 2.24011
R26301 DVSS.n8513 DVSS.n8512 2.24011
R26302 DVSS.n8516 DVSS.n1083 2.24011
R26303 DVSS.n8518 DVSS.n1083 2.24011
R26304 DVSS.n8525 DVSS.n8524 2.24011
R26305 DVSS.n8532 DVSS.n8528 2.24011
R26306 DVSS.n8532 DVSS.n1079 2.24011
R26307 DVSS.n7148 DVSS.n7144 2.24011
R26308 DVSS.n7118 DVSS.n7115 2.24011
R26309 DVSS.n1547 DVSS.n1546 2.24011
R26310 DVSS.n8339 DVSS.n1439 2.24011
R26311 DVSS.n7123 DVSS.n7122 2.24011
R26312 DVSS.n7127 DVSS.n7125 2.24011
R26313 DVSS.n1296 DVSS.n1217 2.24011
R26314 DVSS.n1296 DVSS.n1219 2.24011
R26315 DVSS.n8331 DVSS.n8330 2.24011
R26316 DVSS.n8331 DVSS.n8329 2.24011
R26317 DVSS.n1528 DVSS.n1524 2.24011
R26318 DVSS.n8212 DVSS.n1529 2.24011
R26319 DVSS.n7083 DVSS.n7079 2.24011
R26320 DVSS.n8522 DVSS.n1080 2.24011
R26321 DVSS.n8523 DVSS.n8522 2.24011
R26322 DVSS.n8517 DVSS.n1082 2.24011
R26323 DVSS.n8510 DVSS.n1084 2.24011
R26324 DVSS.n8511 DVSS.n8510 2.24011
R26325 DVSS.n8504 DVSS.n1086 2.24011
R26326 DVSS.n8505 DVSS.n8504 2.24011
R26327 DVSS.n8530 DVSS.n1076 2.24011
R26328 DVSS.n7150 DVSS.n7140 2.24011
R26329 DVSS.n7116 DVSS.n1484 2.24011
R26330 DVSS.n7119 DVSS.n7075 2.24011
R26331 DVSS.n7109 DVSS.n7086 2.24011
R26332 DVSS.n7098 DVSS.n7088 2.24011
R26333 DVSS.n8337 DVSS.n8336 2.24011
R26334 DVSS.n1550 DVSS.n1544 2.24011
R26335 DVSS.n7129 DVSS.n7073 2.24011
R26336 DVSS.n1294 DVSS.n1214 2.24011
R26337 DVSS.n1218 DVSS.n1214 2.24011
R26338 DVSS.n5835 DVSS.n5834 2.23714
R26339 DVSS.n5837 DVSS.n3045 2.23714
R26340 DVSS.n5834 DVSS.n3053 2.23714
R26341 DVSS.n5837 DVSS.n3044 2.23714
R26342 DVSS.n5834 DVSS.n3052 2.23714
R26343 DVSS.n5837 DVSS.n3043 2.23714
R26344 DVSS.n5829 DVSS.n3055 2.23714
R26345 DVSS.n5831 DVSS.n3061 2.23714
R26346 DVSS.n5829 DVSS.n3068 2.23714
R26347 DVSS.n5831 DVSS.n3060 2.23714
R26348 DVSS.n5829 DVSS.n3067 2.23714
R26349 DVSS.n5674 DVSS.n5673 2.23714
R26350 DVSS.n5677 DVSS.n3256 2.23714
R26351 DVSS.n5675 DVSS.n5674 2.23714
R26352 DVSS.n5666 DVSS.n5665 2.23714
R26353 DVSS.n5668 DVSS.n3259 2.23714
R26354 DVSS.n5665 DVSS.n3258 2.23714
R26355 DVSS.n5899 DVSS.n2968 2.18432
R26356 DVSS.n5900 DVSS.n5899 2.18432
R26357 DVSS.n5897 DVSS.n2978 2.18432
R26358 DVSS.n5897 DVSS.n5896 2.18432
R26359 DVSS.n5671 DVSS.n5670 1.5539
R26360 DVSS.n5830 DVSS.n3066 1.53005
R26361 DVSS.n3871 DVSS.n3860 1.52689
R26362 DVSS.n9532 DVSS.n48 1.5005
R26363 DVSS.n9531 DVSS.n9530 1.5005
R26364 DVSS.n9529 DVSS.n9528 1.5005
R26365 DVSS.n9527 DVSS.n9526 1.5005
R26366 DVSS.n9525 DVSS.n9524 1.5005
R26367 DVSS.n9523 DVSS.n9522 1.5005
R26368 DVSS.n9521 DVSS.n9520 1.5005
R26369 DVSS.n9519 DVSS.n9518 1.5005
R26370 DVSS.n9517 DVSS.n9516 1.5005
R26371 DVSS.n9515 DVSS.n9514 1.5005
R26372 DVSS.n9513 DVSS.n9512 1.5005
R26373 DVSS.n9511 DVSS.n9510 1.5005
R26374 DVSS.n9509 DVSS.n9508 1.5005
R26375 DVSS.n9507 DVSS.n9506 1.5005
R26376 DVSS.n9505 DVSS.n9504 1.5005
R26377 DVSS.n9503 DVSS.n9502 1.5005
R26378 DVSS.n9501 DVSS.n9500 1.5005
R26379 DVSS.n9499 DVSS.n9498 1.5005
R26380 DVSS.n9497 DVSS.n9496 1.5005
R26381 DVSS.n9495 DVSS.n9494 1.5005
R26382 DVSS.n9493 DVSS.n9492 1.5005
R26383 DVSS.n9491 DVSS.n9490 1.5005
R26384 DVSS.n9489 DVSS.n9488 1.5005
R26385 DVSS.n9487 DVSS.n9486 1.5005
R26386 DVSS.n9485 DVSS.n9484 1.5005
R26387 DVSS.n9483 DVSS.n9482 1.5005
R26388 DVSS.n9481 DVSS.n9480 1.5005
R26389 DVSS.n9479 DVSS.n9478 1.5005
R26390 DVSS.n9477 DVSS.n9476 1.5005
R26391 DVSS.n9475 DVSS.n337 1.5005
R26392 DVSS.n9474 DVSS.n9473 1.5005
R26393 DVSS.n9469 DVSS.n338 1.5005
R26394 DVSS.n9468 DVSS.n9467 1.5005
R26395 DVSS.n9466 DVSS.n9465 1.5005
R26396 DVSS.n9464 DVSS.n9463 1.5005
R26397 DVSS.n9462 DVSS.n9461 1.5005
R26398 DVSS.n9460 DVSS.n9459 1.5005
R26399 DVSS.n9458 DVSS.n9457 1.5005
R26400 DVSS.n9456 DVSS.n9455 1.5005
R26401 DVSS.n9454 DVSS.n9453 1.5005
R26402 DVSS.n9452 DVSS.n9451 1.5005
R26403 DVSS.n9450 DVSS.n9449 1.5005
R26404 DVSS.n9448 DVSS.n9447 1.5005
R26405 DVSS.n9446 DVSS.n9445 1.5005
R26406 DVSS.n9444 DVSS.n9443 1.5005
R26407 DVSS.n9442 DVSS.n9441 1.5005
R26408 DVSS.n9440 DVSS.n9439 1.5005
R26409 DVSS.n9438 DVSS.n9437 1.5005
R26410 DVSS.n9436 DVSS.n9435 1.5005
R26411 DVSS.n9434 DVSS.n9433 1.5005
R26412 DVSS.n9432 DVSS.n9431 1.5005
R26413 DVSS.n9430 DVSS.n9429 1.5005
R26414 DVSS.n9428 DVSS.n9427 1.5005
R26415 DVSS.n9426 DVSS.n9425 1.5005
R26416 DVSS.n9424 DVSS.n9423 1.5005
R26417 DVSS.n9422 DVSS.n9421 1.5005
R26418 DVSS.n8999 DVSS.n8998 1.5005
R26419 DVSS.n722 DVSS.n721 1.5005
R26420 DVSS.n8994 DVSS.n8993 1.5005
R26421 DVSS.n8992 DVSS.n749 1.5005
R26422 DVSS.n8991 DVSS.n8990 1.5005
R26423 DVSS.n8989 DVSS.n8988 1.5005
R26424 DVSS.n8987 DVSS.n8986 1.5005
R26425 DVSS.n8985 DVSS.n8984 1.5005
R26426 DVSS.n8983 DVSS.n8982 1.5005
R26427 DVSS.n8981 DVSS.n8980 1.5005
R26428 DVSS.n8979 DVSS.n8978 1.5005
R26429 DVSS.n8977 DVSS.n8976 1.5005
R26430 DVSS.n8975 DVSS.n8974 1.5005
R26431 DVSS.n8973 DVSS.n8972 1.5005
R26432 DVSS.n8971 DVSS.n8970 1.5005
R26433 DVSS.n8969 DVSS.n8968 1.5005
R26434 DVSS.n8967 DVSS.n8966 1.5005
R26435 DVSS.n8965 DVSS.n8964 1.5005
R26436 DVSS.n8963 DVSS.n8962 1.5005
R26437 DVSS.n8961 DVSS.n8960 1.5005
R26438 DVSS.n8959 DVSS.n8958 1.5005
R26439 DVSS.n8957 DVSS.n8956 1.5005
R26440 DVSS.n8955 DVSS.n8954 1.5005
R26441 DVSS.n8953 DVSS.n8952 1.5005
R26442 DVSS.n8951 DVSS.n8950 1.5005
R26443 DVSS.n8949 DVSS.n8948 1.5005
R26444 DVSS.n8947 DVSS.n8946 1.5005
R26445 DVSS.n8945 DVSS.n8944 1.5005
R26446 DVSS.n8943 DVSS.n8942 1.5005
R26447 DVSS.n8941 DVSS.n752 1.5005
R26448 DVSS.n8940 DVSS.n8939 1.5005
R26449 DVSS.n8935 DVSS.n753 1.5005
R26450 DVSS.n8934 DVSS.n8933 1.5005
R26451 DVSS.n8932 DVSS.n8931 1.5005
R26452 DVSS.n8930 DVSS.n8929 1.5005
R26453 DVSS.n8928 DVSS.n8927 1.5005
R26454 DVSS.n8926 DVSS.n8925 1.5005
R26455 DVSS.n8924 DVSS.n8923 1.5005
R26456 DVSS.n8922 DVSS.n8921 1.5005
R26457 DVSS.n8920 DVSS.n8919 1.5005
R26458 DVSS.n8918 DVSS.n8917 1.5005
R26459 DVSS.n8916 DVSS.n8915 1.5005
R26460 DVSS.n8914 DVSS.n8913 1.5005
R26461 DVSS.n8912 DVSS.n8911 1.5005
R26462 DVSS.n8910 DVSS.n8909 1.5005
R26463 DVSS.n8908 DVSS.n8907 1.5005
R26464 DVSS.n8906 DVSS.n8905 1.5005
R26465 DVSS.n8904 DVSS.n8903 1.5005
R26466 DVSS.n8902 DVSS.n8901 1.5005
R26467 DVSS.n8900 DVSS.n8899 1.5005
R26468 DVSS.n8898 DVSS.n8897 1.5005
R26469 DVSS.n8896 DVSS.n8895 1.5005
R26470 DVSS.n8894 DVSS.n8893 1.5005
R26471 DVSS.n8892 DVSS.n8891 1.5005
R26472 DVSS.n8890 DVSS.n8889 1.5005
R26473 DVSS.n8888 DVSS.n8887 1.5005
R26474 DVSS.n6647 DVSS.n6646 1.49571
R26475 DVSS.n7244 DVSS.n7243 1.4956
R26476 DVSS.n1476 DVSS.n1474 1.35477
R26477 DVSS.n8256 DVSS.n1454 1.35477
R26478 DVSS.n8464 DVSS.n1147 1.35477
R26479 DVSS.n8465 DVSS.n1091 1.35477
R26480 DVSS.n7064 DVSS.n7063 1.3133
R26481 DVSS.n8198 DVSS.n1557 1.3133
R26482 DVSS.n1750 DVSS.n1749 1.3133
R26483 DVSS.n6755 DVSS.n6753 1.3133
R26484 DVSS.n8205 DVSS.n1550 1.17883
R26485 DVSS.n7130 DVSS.n7129 1.17883
R26486 DVSS.n5833 DVSS.n5832 0.8825
R26487 DVSS.n7117 DVSS.n1480 0.754554
R26488 DVSS.n8320 DVSS.n1443 0.754554
R26489 DVSS.n8316 DVSS.n1458 0.754554
R26490 DVSS.n7147 DVSS.n7146 0.754554
R26491 DVSS.n7112 DVSS.n7111 0.751716
R26492 DVSS.n7096 DVSS.n1444 0.751716
R26493 DVSS.n7149 DVSS.n7143 0.751716
R26494 DVSS.n8218 DVSS.n8217 0.751716
R26495 DVSS.n8527 DVSS.n8526 0.751716
R26496 DVSS.n8515 DVSS.n8514 0.751716
R26497 DVSS.n7106 DVSS.n7077 0.751716
R26498 DVSS.n8338 DVSS.n1440 0.751716
R26499 DVSS.n1216 DVSS.n1215 0.746446
R26500 DVSS.n8509 DVSS.n8508 0.746446
R26501 DVSS.n7128 DVSS.n7124 0.746446
R26502 DVSS.n1545 DVSS.n1438 0.746446
R26503 DVSS.n8320 DVSS.n8319 0.743357
R26504 DVSS.n8319 DVSS.n8318 0.743357
R26505 DVSS.n8296 DVSS.n8295 0.743357
R26506 DVSS.n8297 DVSS.n8296 0.743357
R26507 DVSS.n1480 DVSS.n1477 0.743357
R26508 DVSS.n8297 DVSS.n1477 0.743357
R26509 DVSS.n1455 DVSS.n1450 0.743357
R26510 DVSS.n8318 DVSS.n1455 0.743357
R26511 DVSS.n8298 DVSS.n1475 0.743357
R26512 DVSS.n8298 DVSS.n8297 0.743357
R26513 DVSS.n8317 DVSS.n8316 0.743357
R26514 DVSS.n8318 DVSS.n8317 0.743357
R26515 DVSS.n1459 DVSS.n1453 0.743357
R26516 DVSS.n8318 DVSS.n1453 0.743357
R26517 DVSS.n7146 DVSS.n1473 0.743357
R26518 DVSS.n8297 DVSS.n1473 0.743357
R26519 DVSS.n6436 DVSS.n6016 0.682336
R26520 DVSS.n6159 DVSS.n6158 0.682336
R26521 DVSS.n6045 DVSS.n6017 0.682078
R26522 DVSS.n6642 DVSS.n6641 0.682078
R26523 DVSS.n8070 DVSS 0.66425
R26524 DVSS.n1758 DVSS 0.66425
R26525 DVSS.n2582 DVSS 0.66425
R26526 DVSS.n2116 DVSS 0.66425
R26527 DVSS.n5672 DVSS 0.66425
R26528 DVSS.n2962 DVSS 0.66425
R26529 DVSS.n3025 DVSS 0.66425
R26530 DVSS.n2920 DVSS 0.66425
R26531 DVSS.n8192 DVSS 0.66425
R26532 DVSS.n4441 DVSS 0.66425
R26533 DVSS.n3593 DVSS 0.66425
R26534 DVSS.n3537 DVSS 0.66425
R26535 DVSS.n5379 DVSS 0.66425
R26536 DVSS.n2987 DVSS 0.66425
R26537 DVSS.n2971 DVSS 0.66425
R26538 DVSS.n7362 DVSS 0.66425
R26539 DVSS.n7709 DVSS 0.66425
R26540 DVSS.n6749 DVSS 0.66425
R26541 DVSS.n4934 DVSS.n2915 0.623413
R26542 DVSS.n5906 DVSS.n5905 0.623413
R26543 DVSS.n7707 DVSS.n7699 0.623413
R26544 DVSS.n4449 DVSS.n3020 0.623413
R26545 DVSS.n5891 DVSS.n5890 0.623413
R26546 DVSS.n7372 DVSS.n7371 0.623413
R26547 DVSS.n8183 DVSS.n1751 0.616858
R26548 DVSS.n8068 DVSS.n1914 0.616858
R26549 DVSS.n3626 DVSS.n3579 0.612075
R26550 DVSS.n5535 DVSS.n3301 0.612075
R26551 DVSS.n7723 DVSS.n2094 0.612075
R26552 DVSS.n4842 DVSS.n3569 0.612075
R26553 DVSS.n5545 DVSS.n3293 0.612075
R26554 DVSS.n7853 DVSS.n2086 0.612075
R26555 DVSS.n3999 DVSS.n3712 0.612075
R26556 DVSS.n5652 DVSS.n3241 0.612075
R26557 DVSS.n7340 DVSS.n2609 0.612075
R26558 DVSS.n4191 DVSS.n4190 0.612075
R26559 DVSS.n5662 DVSS.n3250 0.612075
R26560 DVSS.n7350 DVSS.n2601 0.612075
R26561 DVSS.n7359 DVSS.n2594 0.612075
R26562 DVSS.n4980 DVSS.n4979 0.612075
R26563 DVSS.n5526 DVSS.n5516 0.612075
R26564 DVSS.n7716 DVSS.n2102 0.612075
R26565 DVSS.n8201 DVSS.n1553 0.611189
R26566 DVSS.n1859 DVSS.n1538 0.611189
R26567 DVSS.n6650 DVSS.n1885 0.611189
R26568 DVSS.n6655 DVSS.n1895 0.611189
R26569 DVSS.n6659 DVSS.n1904 0.611189
R26570 DVSS.n8194 DVSS.n1560 0.611189
R26571 DVSS.n5911 DVSS.n5910 0.608354
R26572 DVSS.n5881 DVSS.n5880 0.608354
R26573 DVSS.n5129 DVSS.n3315 0.602685
R26574 DVSS.n5395 DVSS.n5394 0.602685
R26575 DVSS.n5776 DVSS.n3157 0.602685
R26576 DVSS.n5812 DVSS.n3113 0.602685
R26577 DVSS.n5365 DVSS.n3311 0.602685
R26578 DVSS.n4479 DVSS.n4461 0.513801
R26579 DVSS.n5936 DVSS.n2890 0.513519
R26580 DVSS.n5939 DVSS.n5935 0.5005
R26581 DVSS.n3833 DVSS.n3832 0.5005
R26582 DVSS.n4495 DVSS.n4494 0.5005
R26583 DVSS.n4496 DVSS.n3831 0.5005
R26584 DVSS.n4498 DVSS.n4497 0.5005
R26585 DVSS.n3829 DVSS.n3828 0.5005
R26586 DVSS.n4504 DVSS.n4503 0.5005
R26587 DVSS.n4505 DVSS.n3827 0.5005
R26588 DVSS.n4507 DVSS.n4506 0.5005
R26589 DVSS.n3814 DVSS.n3813 0.5005
R26590 DVSS.n4522 DVSS.n4521 0.5005
R26591 DVSS.n4523 DVSS.n3812 0.5005
R26592 DVSS.n4525 DVSS.n4524 0.5005
R26593 DVSS.n3810 DVSS.n3809 0.5005
R26594 DVSS.n4530 DVSS.n4529 0.5005
R26595 DVSS.n4531 DVSS.n3808 0.5005
R26596 DVSS.n4578 DVSS.n4532 0.5005
R26597 DVSS.n4577 DVSS.n4533 0.5005
R26598 DVSS.n4575 DVSS.n4534 0.5005
R26599 DVSS.n4573 DVSS.n4535 0.5005
R26600 DVSS.n4538 DVSS.n4536 0.5005
R26601 DVSS.n4569 DVSS.n4539 0.5005
R26602 DVSS.n4568 DVSS.n4540 0.5005
R26603 DVSS.n4567 DVSS.n4541 0.5005
R26604 DVSS.n4544 DVSS.n4542 0.5005
R26605 DVSS.n4563 DVSS.n4545 0.5005
R26606 DVSS.n4562 DVSS.n4546 0.5005
R26607 DVSS.n4561 DVSS.n4547 0.5005
R26608 DVSS.n4550 DVSS.n4548 0.5005
R26609 DVSS.n4557 DVSS.n4551 0.5005
R26610 DVSS.n4556 DVSS.n4552 0.5005
R26611 DVSS.n4555 DVSS.n4554 0.5005
R26612 DVSS.n4553 DVSS.n3747 0.5005
R26613 DVSS.n4780 DVSS.n3748 0.5005
R26614 DVSS.n4779 DVSS.n3749 0.5005
R26615 DVSS.n4777 DVSS.n3750 0.5005
R26616 DVSS.n3753 DVSS.n3751 0.5005
R26617 DVSS.n4773 DVSS.n3754 0.5005
R26618 DVSS.n4772 DVSS.n3755 0.5005
R26619 DVSS.n4771 DVSS.n3756 0.5005
R26620 DVSS.n3759 DVSS.n3757 0.5005
R26621 DVSS.n4767 DVSS.n3760 0.5005
R26622 DVSS.n4766 DVSS.n3761 0.5005
R26623 DVSS.n4765 DVSS.n3762 0.5005
R26624 DVSS.n3765 DVSS.n3763 0.5005
R26625 DVSS.n4761 DVSS.n3766 0.5005
R26626 DVSS.n4760 DVSS.n3767 0.5005
R26627 DVSS.n4759 DVSS.n3768 0.5005
R26628 DVSS.n4610 DVSS.n3769 0.5005
R26629 DVSS.n4611 DVSS.n4609 0.5005
R26630 DVSS.n4753 DVSS.n4612 0.5005
R26631 DVSS.n4752 DVSS.n4613 0.5005
R26632 DVSS.n4751 DVSS.n4614 0.5005
R26633 DVSS.n4706 DVSS.n4615 0.5005
R26634 DVSS.n4743 DVSS.n4707 0.5005
R26635 DVSS.n4742 DVSS.n4708 0.5005
R26636 DVSS.n4741 DVSS.n4709 0.5005
R26637 DVSS.n4712 DVSS.n4710 0.5005
R26638 DVSS.n4737 DVSS.n4713 0.5005
R26639 DVSS.n4736 DVSS.n4714 0.5005
R26640 DVSS.n4735 DVSS.n4715 0.5005
R26641 DVSS.n4718 DVSS.n4716 0.5005
R26642 DVSS.n4731 DVSS.n4719 0.5005
R26643 DVSS.n4730 DVSS.n4720 0.5005
R26644 DVSS.n4729 DVSS.n4721 0.5005
R26645 DVSS.n4726 DVSS.n4722 0.5005
R26646 DVSS.n4725 DVSS.n4724 0.5005
R26647 DVSS.n4723 DVSS.n2794 0.5005
R26648 DVSS.n5998 DVSS.n2795 0.5005
R26649 DVSS.n5997 DVSS.n2796 0.5005
R26650 DVSS.n5995 DVSS.n2797 0.5005
R26651 DVSS.n2800 DVSS.n2798 0.5005
R26652 DVSS.n5991 DVSS.n2801 0.5005
R26653 DVSS.n5990 DVSS.n2802 0.5005
R26654 DVSS.n5989 DVSS.n2803 0.5005
R26655 DVSS.n2806 DVSS.n2804 0.5005
R26656 DVSS.n5985 DVSS.n2807 0.5005
R26657 DVSS.n5984 DVSS.n2808 0.5005
R26658 DVSS.n5983 DVSS.n2809 0.5005
R26659 DVSS.n2812 DVSS.n2810 0.5005
R26660 DVSS.n5979 DVSS.n2813 0.5005
R26661 DVSS.n5978 DVSS.n2814 0.5005
R26662 DVSS.n5977 DVSS.n2815 0.5005
R26663 DVSS.n2837 DVSS.n2816 0.5005
R26664 DVSS.n5971 DVSS.n2838 0.5005
R26665 DVSS.n5970 DVSS.n2839 0.5005
R26666 DVSS.n5968 DVSS.n2840 0.5005
R26667 DVSS.n2843 DVSS.n2841 0.5005
R26668 DVSS.n5964 DVSS.n2844 0.5005
R26669 DVSS.n5963 DVSS.n2845 0.5005
R26670 DVSS.n5962 DVSS.n2846 0.5005
R26671 DVSS.n2866 DVSS.n2847 0.5005
R26672 DVSS.n5954 DVSS.n2867 0.5005
R26673 DVSS.n5953 DVSS.n2868 0.5005
R26674 DVSS.n5951 DVSS.n2869 0.5005
R26675 DVSS.n2872 DVSS.n2870 0.5005
R26676 DVSS.n5947 DVSS.n2873 0.5005
R26677 DVSS.n5946 DVSS.n2874 0.5005
R26678 DVSS.n5945 DVSS.n2875 0.5005
R26679 DVSS.n5934 DVSS.n2876 0.5005
R26680 DVSS.n5938 DVSS.n5937 0.5005
R26681 DVSS.n5940 DVSS.n5939 0.5005
R26682 DVSS.n4481 DVSS.n4480 0.5005
R26683 DVSS.n4489 DVSS.n3833 0.5005
R26684 DVSS.n4494 DVSS.n4493 0.5005
R26685 DVSS.n3831 DVSS.n3830 0.5005
R26686 DVSS.n4499 DVSS.n4498 0.5005
R26687 DVSS.n4500 DVSS.n3829 0.5005
R26688 DVSS.n4503 DVSS.n4502 0.5005
R26689 DVSS.n4501 DVSS.n3827 0.5005
R26690 DVSS.n4508 DVSS.n4507 0.5005
R26691 DVSS.n4516 DVSS.n3814 0.5005
R26692 DVSS.n4521 DVSS.n4520 0.5005
R26693 DVSS.n3812 DVSS.n3811 0.5005
R26694 DVSS.n4526 DVSS.n4525 0.5005
R26695 DVSS.n4527 DVSS.n3810 0.5005
R26696 DVSS.n4529 DVSS.n4528 0.5005
R26697 DVSS.n3808 DVSS.n3802 0.5005
R26698 DVSS.n4579 DVSS.n4578 0.5005
R26699 DVSS.n4577 DVSS.n4576 0.5005
R26700 DVSS.n4575 DVSS.n4574 0.5005
R26701 DVSS.n4573 DVSS.n4572 0.5005
R26702 DVSS.n4571 DVSS.n4536 0.5005
R26703 DVSS.n4570 DVSS.n4569 0.5005
R26704 DVSS.n4568 DVSS.n4537 0.5005
R26705 DVSS.n4567 DVSS.n4566 0.5005
R26706 DVSS.n4565 DVSS.n4542 0.5005
R26707 DVSS.n4564 DVSS.n4563 0.5005
R26708 DVSS.n4562 DVSS.n4543 0.5005
R26709 DVSS.n4561 DVSS.n4560 0.5005
R26710 DVSS.n4559 DVSS.n4548 0.5005
R26711 DVSS.n4558 DVSS.n4557 0.5005
R26712 DVSS.n4556 DVSS.n4549 0.5005
R26713 DVSS.n4555 DVSS.n3730 0.5005
R26714 DVSS.n3747 DVSS.n3735 0.5005
R26715 DVSS.n4781 DVSS.n4780 0.5005
R26716 DVSS.n4779 DVSS.n4778 0.5005
R26717 DVSS.n4777 DVSS.n4776 0.5005
R26718 DVSS.n4775 DVSS.n3751 0.5005
R26719 DVSS.n4774 DVSS.n4773 0.5005
R26720 DVSS.n4772 DVSS.n3752 0.5005
R26721 DVSS.n4771 DVSS.n4770 0.5005
R26722 DVSS.n4769 DVSS.n3757 0.5005
R26723 DVSS.n4768 DVSS.n4767 0.5005
R26724 DVSS.n4766 DVSS.n3758 0.5005
R26725 DVSS.n4765 DVSS.n4764 0.5005
R26726 DVSS.n4763 DVSS.n3763 0.5005
R26727 DVSS.n4762 DVSS.n4761 0.5005
R26728 DVSS.n4760 DVSS.n3764 0.5005
R26729 DVSS.n4759 DVSS.n4758 0.5005
R26730 DVSS.n3775 DVSS.n3769 0.5005
R26731 DVSS.n4609 DVSS.n4607 0.5005
R26732 DVSS.n4754 DVSS.n4753 0.5005
R26733 DVSS.n4752 DVSS.n4608 0.5005
R26734 DVSS.n4751 DVSS.n4750 0.5005
R26735 DVSS.n4622 DVSS.n4615 0.5005
R26736 DVSS.n4744 DVSS.n4743 0.5005
R26737 DVSS.n4742 DVSS.n4705 0.5005
R26738 DVSS.n4741 DVSS.n4740 0.5005
R26739 DVSS.n4739 DVSS.n4710 0.5005
R26740 DVSS.n4738 DVSS.n4737 0.5005
R26741 DVSS.n4736 DVSS.n4711 0.5005
R26742 DVSS.n4735 DVSS.n4734 0.5005
R26743 DVSS.n4733 DVSS.n4716 0.5005
R26744 DVSS.n4732 DVSS.n4731 0.5005
R26745 DVSS.n4730 DVSS.n4717 0.5005
R26746 DVSS.n4729 DVSS.n4728 0.5005
R26747 DVSS.n4727 DVSS.n4726 0.5005
R26748 DVSS.n4725 DVSS.n2783 0.5005
R26749 DVSS.n2794 DVSS.n2789 0.5005
R26750 DVSS.n5999 DVSS.n5998 0.5005
R26751 DVSS.n5997 DVSS.n5996 0.5005
R26752 DVSS.n5995 DVSS.n5994 0.5005
R26753 DVSS.n5993 DVSS.n2798 0.5005
R26754 DVSS.n5992 DVSS.n5991 0.5005
R26755 DVSS.n5990 DVSS.n2799 0.5005
R26756 DVSS.n5989 DVSS.n5988 0.5005
R26757 DVSS.n5987 DVSS.n2804 0.5005
R26758 DVSS.n5986 DVSS.n5985 0.5005
R26759 DVSS.n5984 DVSS.n2805 0.5005
R26760 DVSS.n5983 DVSS.n5982 0.5005
R26761 DVSS.n5981 DVSS.n2810 0.5005
R26762 DVSS.n5980 DVSS.n5979 0.5005
R26763 DVSS.n5978 DVSS.n2811 0.5005
R26764 DVSS.n5977 DVSS.n5976 0.5005
R26765 DVSS.n2822 DVSS.n2816 0.5005
R26766 DVSS.n5972 DVSS.n5971 0.5005
R26767 DVSS.n5970 DVSS.n5969 0.5005
R26768 DVSS.n5968 DVSS.n5967 0.5005
R26769 DVSS.n5966 DVSS.n2841 0.5005
R26770 DVSS.n5965 DVSS.n5964 0.5005
R26771 DVSS.n5963 DVSS.n2842 0.5005
R26772 DVSS.n5962 DVSS.n5961 0.5005
R26773 DVSS.n2853 DVSS.n2847 0.5005
R26774 DVSS.n5955 DVSS.n5954 0.5005
R26775 DVSS.n5953 DVSS.n5952 0.5005
R26776 DVSS.n5951 DVSS.n5950 0.5005
R26777 DVSS.n5949 DVSS.n2870 0.5005
R26778 DVSS.n5948 DVSS.n5947 0.5005
R26779 DVSS.n5946 DVSS.n2871 0.5005
R26780 DVSS.n5945 DVSS.n5944 0.5005
R26781 DVSS.n2882 DVSS.n2876 0.5005
R26782 DVSS.n4600 DVSS.n4599 0.466338
R26783 DVSS.n6009 DVSS.n6008 0.466338
R26784 DVSS.n4596 DVSS.n4595 0.46307
R26785 DVSS.n6006 DVSS.n2777 0.46307
R26786 DVSS.n6858 DVSS.n6738 0.462685
R26787 DVSS.n8060 DVSS.n1919 0.462685
R26788 DVSS.n5879 DVSS.n2997 0.462685
R26789 DVSS.n5864 DVSS.n3030 0.462685
R26790 DVSS.n4451 DVSS.n3839 0.462685
R26791 DVSS.n1742 DVSS.n1563 0.462428
R26792 DVSS.n8174 DVSS.n8170 0.462428
R26793 DVSS.n5094 DVSS.n2941 0.462428
R26794 DVSS.n5330 DVSS.n2923 0.462428
R26795 DVSS.n4939 DVSS.n4926 0.462428
R26796 DVSS.n6641 DVSS.n6018 0.455549
R26797 DVSS.n6437 DVSS.n6436 0.455549
R26798 DVSS.n6048 DVSS.n6045 0.455549
R26799 DVSS.n6159 DVSS.n6155 0.455549
R26800 DVSS.n4938 DVSS.n4936 0.4505
R26801 DVSS.n4237 DVSS.n4234 0.4505
R26802 DVSS.n4240 DVSS.n4239 0.4505
R26803 DVSS.n4241 DVSS.n4233 0.4505
R26804 DVSS.n4243 DVSS.n4242 0.4505
R26805 DVSS.n4231 DVSS.n4230 0.4505
R26806 DVSS.n4248 DVSS.n4247 0.4505
R26807 DVSS.n4249 DVSS.n4229 0.4505
R26808 DVSS.n4251 DVSS.n4250 0.4505
R26809 DVSS.n4214 DVSS.n4213 0.4505
R26810 DVSS.n4263 DVSS.n4262 0.4505
R26811 DVSS.n4264 DVSS.n4212 0.4505
R26812 DVSS.n4266 DVSS.n4265 0.4505
R26813 DVSS.n4210 DVSS.n4209 0.4505
R26814 DVSS.n4271 DVSS.n4270 0.4505
R26815 DVSS.n4272 DVSS.n4206 0.4505
R26816 DVSS.n4417 DVSS.n4416 0.4505
R26817 DVSS.n4415 DVSS.n4208 0.4505
R26818 DVSS.n4414 DVSS.n4413 0.4505
R26819 DVSS.n4411 DVSS.n4273 0.4505
R26820 DVSS.n4277 DVSS.n4274 0.4505
R26821 DVSS.n4407 DVSS.n4406 0.4505
R26822 DVSS.n4405 DVSS.n4276 0.4505
R26823 DVSS.n4404 DVSS.n4403 0.4505
R26824 DVSS.n4279 DVSS.n4278 0.4505
R26825 DVSS.n4399 DVSS.n4398 0.4505
R26826 DVSS.n4397 DVSS.n4281 0.4505
R26827 DVSS.n4396 DVSS.n4395 0.4505
R26828 DVSS.n4283 DVSS.n4282 0.4505
R26829 DVSS.n4391 DVSS.n4390 0.4505
R26830 DVSS.n4389 DVSS.n4285 0.4505
R26831 DVSS.n4388 DVSS.n4387 0.4505
R26832 DVSS.n4386 DVSS.n4286 0.4505
R26833 DVSS.n4385 DVSS.n4383 0.4505
R26834 DVSS.n4382 DVSS.n4288 0.4505
R26835 DVSS.n4381 DVSS.n4380 0.4505
R26836 DVSS.n4290 DVSS.n4289 0.4505
R26837 DVSS.n4376 DVSS.n4375 0.4505
R26838 DVSS.n4374 DVSS.n4292 0.4505
R26839 DVSS.n4373 DVSS.n4372 0.4505
R26840 DVSS.n4294 DVSS.n4293 0.4505
R26841 DVSS.n4368 DVSS.n4367 0.4505
R26842 DVSS.n4366 DVSS.n4296 0.4505
R26843 DVSS.n4365 DVSS.n4364 0.4505
R26844 DVSS.n4298 DVSS.n4297 0.4505
R26845 DVSS.n4360 DVSS.n4359 0.4505
R26846 DVSS.n4358 DVSS.n4300 0.4505
R26847 DVSS.n4357 DVSS.n4356 0.4505
R26848 DVSS.n4355 DVSS.n4301 0.4505
R26849 DVSS.n4354 DVSS.n4352 0.4505
R26850 DVSS.n4351 DVSS.n4303 0.4505
R26851 DVSS.n4350 DVSS.n4349 0.4505
R26852 DVSS.n4348 DVSS.n4304 0.4505
R26853 DVSS.n4347 DVSS.n4345 0.4505
R26854 DVSS.n4344 DVSS.n4305 0.4505
R26855 DVSS.n4343 DVSS.n4342 0.4505
R26856 DVSS.n4307 DVSS.n4306 0.4505
R26857 DVSS.n4338 DVSS.n4337 0.4505
R26858 DVSS.n4336 DVSS.n4310 0.4505
R26859 DVSS.n4335 DVSS.n4334 0.4505
R26860 DVSS.n4312 DVSS.n4311 0.4505
R26861 DVSS.n4330 DVSS.n4329 0.4505
R26862 DVSS.n4328 DVSS.n4314 0.4505
R26863 DVSS.n4327 DVSS.n4326 0.4505
R26864 DVSS.n4316 DVSS.n4315 0.4505
R26865 DVSS.n4322 DVSS.n4321 0.4505
R26866 DVSS.n4320 DVSS.n4317 0.4505
R26867 DVSS.n4319 DVSS.n4318 0.4505
R26868 DVSS.n3646 DVSS.n3645 0.4505
R26869 DVSS.n4853 DVSS.n4852 0.4505
R26870 DVSS.n4854 DVSS.n3644 0.4505
R26871 DVSS.n4856 DVSS.n4855 0.4505
R26872 DVSS.n3642 DVSS.n3641 0.4505
R26873 DVSS.n4861 DVSS.n4860 0.4505
R26874 DVSS.n4862 DVSS.n3640 0.4505
R26875 DVSS.n4864 DVSS.n4863 0.4505
R26876 DVSS.n3638 DVSS.n3637 0.4505
R26877 DVSS.n4869 DVSS.n4868 0.4505
R26878 DVSS.n4870 DVSS.n3636 0.4505
R26879 DVSS.n4872 DVSS.n4871 0.4505
R26880 DVSS.n3634 DVSS.n3633 0.4505
R26881 DVSS.n4877 DVSS.n4876 0.4505
R26882 DVSS.n4878 DVSS.n3632 0.4505
R26883 DVSS.n4880 DVSS.n4879 0.4505
R26884 DVSS.n3613 DVSS.n3612 0.4505
R26885 DVSS.n4891 DVSS.n4890 0.4505
R26886 DVSS.n4892 DVSS.n3611 0.4505
R26887 DVSS.n4894 DVSS.n4893 0.4505
R26888 DVSS.n3609 DVSS.n3608 0.4505
R26889 DVSS.n4899 DVSS.n4898 0.4505
R26890 DVSS.n4900 DVSS.n3605 0.4505
R26891 DVSS.n4960 DVSS.n4959 0.4505
R26892 DVSS.n4958 DVSS.n3607 0.4505
R26893 DVSS.n4957 DVSS.n4956 0.4505
R26894 DVSS.n4954 DVSS.n4901 0.4505
R26895 DVSS.n4905 DVSS.n4902 0.4505
R26896 DVSS.n4950 DVSS.n4949 0.4505
R26897 DVSS.n4948 DVSS.n4904 0.4505
R26898 DVSS.n4947 DVSS.n4946 0.4505
R26899 DVSS.n4937 DVSS.n4906 0.4505
R26900 DVSS.n1744 DVSS.n1743 0.4505
R26901 DVSS.n6769 DVSS.n6768 0.4505
R26902 DVSS.n6770 DVSS.n6764 0.4505
R26903 DVSS.n6849 DVSS.n6848 0.4505
R26904 DVSS.n6847 DVSS.n6765 0.4505
R26905 DVSS.n6846 DVSS.n6845 0.4505
R26906 DVSS.n6842 DVSS.n6771 0.4505
R26907 DVSS.n6841 DVSS.n6840 0.4505
R26908 DVSS.n6839 DVSS.n6772 0.4505
R26909 DVSS.n6838 DVSS.n6837 0.4505
R26910 DVSS.n6835 DVSS.n6773 0.4505
R26911 DVSS.n6833 DVSS.n6775 0.4505
R26912 DVSS.n6778 DVSS.n6774 0.4505
R26913 DVSS.n6829 DVSS.n6828 0.4505
R26914 DVSS.n6827 DVSS.n6777 0.4505
R26915 DVSS.n6826 DVSS.n6825 0.4505
R26916 DVSS.n6824 DVSS.n6779 0.4505
R26917 DVSS.n6823 DVSS.n6821 0.4505
R26918 DVSS.n6820 DVSS.n6781 0.4505
R26919 DVSS.n6819 DVSS.n6818 0.4505
R26920 DVSS.n6783 DVSS.n6782 0.4505
R26921 DVSS.n6814 DVSS.n6813 0.4505
R26922 DVSS.n6812 DVSS.n6785 0.4505
R26923 DVSS.n6811 DVSS.n6810 0.4505
R26924 DVSS.n6787 DVSS.n6786 0.4505
R26925 DVSS.n6806 DVSS.n6805 0.4505
R26926 DVSS.n6804 DVSS.n6789 0.4505
R26927 DVSS.n6803 DVSS.n6802 0.4505
R26928 DVSS.n6791 DVSS.n6790 0.4505
R26929 DVSS.n6798 DVSS.n6797 0.4505
R26930 DVSS.n6796 DVSS.n6793 0.4505
R26931 DVSS.n6795 DVSS.n6794 0.4505
R26932 DVSS.n1347 DVSS.n1344 0.4505
R26933 DVSS.n8433 DVSS.n8432 0.4505
R26934 DVSS.n8431 DVSS.n1346 0.4505
R26935 DVSS.n8430 DVSS.n8429 0.4505
R26936 DVSS.n1349 DVSS.n1348 0.4505
R26937 DVSS.n8425 DVSS.n8424 0.4505
R26938 DVSS.n8423 DVSS.n1351 0.4505
R26939 DVSS.n8422 DVSS.n8421 0.4505
R26940 DVSS.n1353 DVSS.n1352 0.4505
R26941 DVSS.n8417 DVSS.n8416 0.4505
R26942 DVSS.n8415 DVSS.n1355 0.4505
R26943 DVSS.n8414 DVSS.n8413 0.4505
R26944 DVSS.n1357 DVSS.n1356 0.4505
R26945 DVSS.n8409 DVSS.n8408 0.4505
R26946 DVSS.n8407 DVSS.n1359 0.4505
R26947 DVSS.n8406 DVSS.n8405 0.4505
R26948 DVSS.n1361 DVSS.n1360 0.4505
R26949 DVSS.n1395 DVSS.n1393 0.4505
R26950 DVSS.n8398 DVSS.n8397 0.4505
R26951 DVSS.n8396 DVSS.n1394 0.4505
R26952 DVSS.n8395 DVSS.n8394 0.4505
R26953 DVSS.n1397 DVSS.n1396 0.4505
R26954 DVSS.n1638 DVSS.n1637 0.4505
R26955 DVSS.n1640 DVSS.n1639 0.4505
R26956 DVSS.n1636 DVSS.n1635 0.4505
R26957 DVSS.n1645 DVSS.n1644 0.4505
R26958 DVSS.n1646 DVSS.n1634 0.4505
R26959 DVSS.n1648 DVSS.n1647 0.4505
R26960 DVSS.n1632 DVSS.n1631 0.4505
R26961 DVSS.n1653 DVSS.n1652 0.4505
R26962 DVSS.n1654 DVSS.n1630 0.4505
R26963 DVSS.n1656 DVSS.n1655 0.4505
R26964 DVSS.n1628 DVSS.n1627 0.4505
R26965 DVSS.n1661 DVSS.n1660 0.4505
R26966 DVSS.n1662 DVSS.n1626 0.4505
R26967 DVSS.n1664 DVSS.n1663 0.4505
R26968 DVSS.n1666 DVSS.n1625 0.4505
R26969 DVSS.n1669 DVSS.n1668 0.4505
R26970 DVSS.n1670 DVSS.n1624 0.4505
R26971 DVSS.n1672 DVSS.n1671 0.4505
R26972 DVSS.n1622 DVSS.n1621 0.4505
R26973 DVSS.n1677 DVSS.n1676 0.4505
R26974 DVSS.n1678 DVSS.n1620 0.4505
R26975 DVSS.n1680 DVSS.n1679 0.4505
R26976 DVSS.n1618 DVSS.n1617 0.4505
R26977 DVSS.n1685 DVSS.n1684 0.4505
R26978 DVSS.n1686 DVSS.n1616 0.4505
R26979 DVSS.n1688 DVSS.n1687 0.4505
R26980 DVSS.n1614 DVSS.n1613 0.4505
R26981 DVSS.n1693 DVSS.n1692 0.4505
R26982 DVSS.n1694 DVSS.n1612 0.4505
R26983 DVSS.n1696 DVSS.n1695 0.4505
R26984 DVSS.n1698 DVSS.n1611 0.4505
R26985 DVSS.n1701 DVSS.n1700 0.4505
R26986 DVSS.n1702 DVSS.n1610 0.4505
R26987 DVSS.n1704 DVSS.n1703 0.4505
R26988 DVSS.n1608 DVSS.n1607 0.4505
R26989 DVSS.n1709 DVSS.n1708 0.4505
R26990 DVSS.n1710 DVSS.n1606 0.4505
R26991 DVSS.n1712 DVSS.n1711 0.4505
R26992 DVSS.n1593 DVSS.n1592 0.4505
R26993 DVSS.n1730 DVSS.n1729 0.4505
R26994 DVSS.n1731 DVSS.n1591 0.4505
R26995 DVSS.n1734 DVSS.n1733 0.4505
R26996 DVSS.n1732 DVSS.n1589 0.4505
R26997 DVSS.n1738 DVSS.n1588 0.4505
R26998 DVSS.n1740 DVSS.n1739 0.4505
R26999 DVSS.n1741 DVSS.n1585 0.4505
R27000 DVSS.n1587 DVSS.n1586 0.4505
R27001 DVSS.n1745 DVSS.n1744 0.4505
R27002 DVSS.n6766 DVSS.n6744 0.4505
R27003 DVSS.n6768 DVSS.n6767 0.4505
R27004 DVSS.n6764 DVSS.n6762 0.4505
R27005 DVSS.n6850 DVSS.n6849 0.4505
R27006 DVSS.n6765 DVSS.n6763 0.4505
R27007 DVSS.n6845 DVSS.n6844 0.4505
R27008 DVSS.n6843 DVSS.n6842 0.4505
R27009 DVSS.n6841 DVSS.n6669 0.4505
R27010 DVSS.n6772 DVSS.n6675 0.4505
R27011 DVSS.n6837 DVSS.n6836 0.4505
R27012 DVSS.n6835 DVSS.n6834 0.4505
R27013 DVSS.n6833 DVSS.n6832 0.4505
R27014 DVSS.n6831 DVSS.n6774 0.4505
R27015 DVSS.n6830 DVSS.n6829 0.4505
R27016 DVSS.n6777 DVSS.n6776 0.4505
R27017 DVSS.n6825 DVSS.n1164 0.4505
R27018 DVSS.n6824 DVSS.n1171 0.4505
R27019 DVSS.n6823 DVSS.n6822 0.4505
R27020 DVSS.n6781 DVSS.n6780 0.4505
R27021 DVSS.n6818 DVSS.n6817 0.4505
R27022 DVSS.n6816 DVSS.n6783 0.4505
R27023 DVSS.n6815 DVSS.n6814 0.4505
R27024 DVSS.n6785 DVSS.n6784 0.4505
R27025 DVSS.n6810 DVSS.n6809 0.4505
R27026 DVSS.n6808 DVSS.n6787 0.4505
R27027 DVSS.n6807 DVSS.n6806 0.4505
R27028 DVSS.n6789 DVSS.n6788 0.4505
R27029 DVSS.n6802 DVSS.n6801 0.4505
R27030 DVSS.n6800 DVSS.n6791 0.4505
R27031 DVSS.n6799 DVSS.n6798 0.4505
R27032 DVSS.n6793 DVSS.n6792 0.4505
R27033 DVSS.n6794 DVSS.n1328 0.4505
R27034 DVSS.n1344 DVSS.n1334 0.4505
R27035 DVSS.n8434 DVSS.n8433 0.4505
R27036 DVSS.n1346 DVSS.n1345 0.4505
R27037 DVSS.n8429 DVSS.n8428 0.4505
R27038 DVSS.n8427 DVSS.n1349 0.4505
R27039 DVSS.n8426 DVSS.n8425 0.4505
R27040 DVSS.n1351 DVSS.n1350 0.4505
R27041 DVSS.n8421 DVSS.n8420 0.4505
R27042 DVSS.n8419 DVSS.n1353 0.4505
R27043 DVSS.n8418 DVSS.n8417 0.4505
R27044 DVSS.n1355 DVSS.n1354 0.4505
R27045 DVSS.n8413 DVSS.n8412 0.4505
R27046 DVSS.n8411 DVSS.n1357 0.4505
R27047 DVSS.n8410 DVSS.n8409 0.4505
R27048 DVSS.n1359 DVSS.n1358 0.4505
R27049 DVSS.n8405 DVSS.n8404 0.4505
R27050 DVSS.n1367 DVSS.n1361 0.4505
R27051 DVSS.n1393 DVSS.n1388 0.4505
R27052 DVSS.n8399 DVSS.n8398 0.4505
R27053 DVSS.n1394 DVSS.n1392 0.4505
R27054 DVSS.n8394 DVSS.n8393 0.4505
R27055 DVSS.n1404 DVSS.n1397 0.4505
R27056 DVSS.n1637 DVSS.n1414 0.4505
R27057 DVSS.n1641 DVSS.n1640 0.4505
R27058 DVSS.n1642 DVSS.n1636 0.4505
R27059 DVSS.n1644 DVSS.n1643 0.4505
R27060 DVSS.n1634 DVSS.n1633 0.4505
R27061 DVSS.n1649 DVSS.n1648 0.4505
R27062 DVSS.n1650 DVSS.n1632 0.4505
R27063 DVSS.n1652 DVSS.n1651 0.4505
R27064 DVSS.n1630 DVSS.n1629 0.4505
R27065 DVSS.n1657 DVSS.n1656 0.4505
R27066 DVSS.n1658 DVSS.n1628 0.4505
R27067 DVSS.n1660 DVSS.n1659 0.4505
R27068 DVSS.n1626 DVSS.n1428 0.4505
R27069 DVSS.n1664 DVSS.n1436 0.4505
R27070 DVSS.n1666 DVSS.n1665 0.4505
R27071 DVSS.n1668 DVSS.n1667 0.4505
R27072 DVSS.n1624 DVSS.n1623 0.4505
R27073 DVSS.n1673 DVSS.n1672 0.4505
R27074 DVSS.n1674 DVSS.n1622 0.4505
R27075 DVSS.n1676 DVSS.n1675 0.4505
R27076 DVSS.n1620 DVSS.n1619 0.4505
R27077 DVSS.n1681 DVSS.n1680 0.4505
R27078 DVSS.n1682 DVSS.n1618 0.4505
R27079 DVSS.n1684 DVSS.n1683 0.4505
R27080 DVSS.n1616 DVSS.n1615 0.4505
R27081 DVSS.n1689 DVSS.n1688 0.4505
R27082 DVSS.n1690 DVSS.n1614 0.4505
R27083 DVSS.n1692 DVSS.n1691 0.4505
R27084 DVSS.n1612 DVSS.n1108 0.4505
R27085 DVSS.n1696 DVSS.n1114 0.4505
R27086 DVSS.n1698 DVSS.n1697 0.4505
R27087 DVSS.n1700 DVSS.n1699 0.4505
R27088 DVSS.n1610 DVSS.n1609 0.4505
R27089 DVSS.n1705 DVSS.n1704 0.4505
R27090 DVSS.n1706 DVSS.n1608 0.4505
R27091 DVSS.n1708 DVSS.n1707 0.4505
R27092 DVSS.n1606 DVSS.n1601 0.4505
R27093 DVSS.n1713 DVSS.n1712 0.4505
R27094 DVSS.n1719 DVSS.n1593 0.4505
R27095 DVSS.n1729 DVSS.n1728 0.4505
R27096 DVSS.n1591 DVSS.n1590 0.4505
R27097 DVSS.n1735 DVSS.n1734 0.4505
R27098 DVSS.n1736 DVSS.n1589 0.4505
R27099 DVSS.n1738 DVSS.n1737 0.4505
R27100 DVSS.n1739 DVSS.n1565 0.4505
R27101 DVSS.n1585 DVSS.n1571 0.4505
R27102 DVSS.n8169 DVSS.n8168 0.4505
R27103 DVSS.n1941 DVSS.n1940 0.4505
R27104 DVSS.n1942 DVSS.n1936 0.4505
R27105 DVSS.n8051 DVSS.n8050 0.4505
R27106 DVSS.n8049 DVSS.n1937 0.4505
R27107 DVSS.n8048 DVSS.n8047 0.4505
R27108 DVSS.n1944 DVSS.n1943 0.4505
R27109 DVSS.n8043 DVSS.n8042 0.4505
R27110 DVSS.n8041 DVSS.n1946 0.4505
R27111 DVSS.n8040 DVSS.n8039 0.4505
R27112 DVSS.n1948 DVSS.n1947 0.4505
R27113 DVSS.n8028 DVSS.n8027 0.4505
R27114 DVSS.n8026 DVSS.n1968 0.4505
R27115 DVSS.n8025 DVSS.n8024 0.4505
R27116 DVSS.n1970 DVSS.n1969 0.4505
R27117 DVSS.n8020 DVSS.n8019 0.4505
R27118 DVSS.n8018 DVSS.n1972 0.4505
R27119 DVSS.n8017 DVSS.n8016 0.4505
R27120 DVSS.n1974 DVSS.n1973 0.4505
R27121 DVSS.n8005 DVSS.n8004 0.4505
R27122 DVSS.n8003 DVSS.n1994 0.4505
R27123 DVSS.n8002 DVSS.n8001 0.4505
R27124 DVSS.n1996 DVSS.n1995 0.4505
R27125 DVSS.n7997 DVSS.n7996 0.4505
R27126 DVSS.n7995 DVSS.n1998 0.4505
R27127 DVSS.n7994 DVSS.n7993 0.4505
R27128 DVSS.n2000 DVSS.n1999 0.4505
R27129 DVSS.n7989 DVSS.n7988 0.4505
R27130 DVSS.n7987 DVSS.n2002 0.4505
R27131 DVSS.n7986 DVSS.n7985 0.4505
R27132 DVSS.n2004 DVSS.n2003 0.4505
R27133 DVSS.n7981 DVSS.n7980 0.4505
R27134 DVSS.n7979 DVSS.n2006 0.4505
R27135 DVSS.n7978 DVSS.n7977 0.4505
R27136 DVSS.n2008 DVSS.n2007 0.4505
R27137 DVSS.n7966 DVSS.n7965 0.4505
R27138 DVSS.n7964 DVSS.n2028 0.4505
R27139 DVSS.n7963 DVSS.n7962 0.4505
R27140 DVSS.n2030 DVSS.n2029 0.4505
R27141 DVSS.n7958 DVSS.n7957 0.4505
R27142 DVSS.n7956 DVSS.n2032 0.4505
R27143 DVSS.n7955 DVSS.n7954 0.4505
R27144 DVSS.n2034 DVSS.n2033 0.4505
R27145 DVSS.n7950 DVSS.n7949 0.4505
R27146 DVSS.n7948 DVSS.n2036 0.4505
R27147 DVSS.n7947 DVSS.n7946 0.4505
R27148 DVSS.n2038 DVSS.n2037 0.4505
R27149 DVSS.n7942 DVSS.n7941 0.4505
R27150 DVSS.n7940 DVSS.n2040 0.4505
R27151 DVSS.n7939 DVSS.n7938 0.4505
R27152 DVSS.n2042 DVSS.n2041 0.4505
R27153 DVSS.n7768 DVSS.n7767 0.4505
R27154 DVSS.n7769 DVSS.n7766 0.4505
R27155 DVSS.n7772 DVSS.n7771 0.4505
R27156 DVSS.n7773 DVSS.n7765 0.4505
R27157 DVSS.n7775 DVSS.n7774 0.4505
R27158 DVSS.n7763 DVSS.n7762 0.4505
R27159 DVSS.n7780 DVSS.n7779 0.4505
R27160 DVSS.n7781 DVSS.n7761 0.4505
R27161 DVSS.n7783 DVSS.n7782 0.4505
R27162 DVSS.n7759 DVSS.n7758 0.4505
R27163 DVSS.n7788 DVSS.n7787 0.4505
R27164 DVSS.n7789 DVSS.n7757 0.4505
R27165 DVSS.n7792 DVSS.n7791 0.4505
R27166 DVSS.n7790 DVSS.n7755 0.4505
R27167 DVSS.n7796 DVSS.n7754 0.4505
R27168 DVSS.n7798 DVSS.n7797 0.4505
R27169 DVSS.n7799 DVSS.n7751 0.4505
R27170 DVSS.n7842 DVSS.n7841 0.4505
R27171 DVSS.n7840 DVSS.n7753 0.4505
R27172 DVSS.n7839 DVSS.n7838 0.4505
R27173 DVSS.n7801 DVSS.n7800 0.4505
R27174 DVSS.n7834 DVSS.n7833 0.4505
R27175 DVSS.n7832 DVSS.n7803 0.4505
R27176 DVSS.n7831 DVSS.n7830 0.4505
R27177 DVSS.n7805 DVSS.n7804 0.4505
R27178 DVSS.n7826 DVSS.n7825 0.4505
R27179 DVSS.n7824 DVSS.n7807 0.4505
R27180 DVSS.n7823 DVSS.n7822 0.4505
R27181 DVSS.n7809 DVSS.n7808 0.4505
R27182 DVSS.n7818 DVSS.n7817 0.4505
R27183 DVSS.n7816 DVSS.n7811 0.4505
R27184 DVSS.n7815 DVSS.n7814 0.4505
R27185 DVSS.n7813 DVSS.n7812 0.4505
R27186 DVSS.n1807 DVSS.n1806 0.4505
R27187 DVSS.n8126 DVSS.n8125 0.4505
R27188 DVSS.n8127 DVSS.n1805 0.4505
R27189 DVSS.n8129 DVSS.n8128 0.4505
R27190 DVSS.n1803 DVSS.n1802 0.4505
R27191 DVSS.n8134 DVSS.n8133 0.4505
R27192 DVSS.n8135 DVSS.n1801 0.4505
R27193 DVSS.n8137 DVSS.n8136 0.4505
R27194 DVSS.n1787 DVSS.n1786 0.4505
R27195 DVSS.n8155 DVSS.n8154 0.4505
R27196 DVSS.n8156 DVSS.n1785 0.4505
R27197 DVSS.n8158 DVSS.n8157 0.4505
R27198 DVSS.n1783 DVSS.n1782 0.4505
R27199 DVSS.n8163 DVSS.n8162 0.4505
R27200 DVSS.n8165 DVSS.n8164 0.4505
R27201 DVSS.n8166 DVSS.n1781 0.4505
R27202 DVSS.n1780 DVSS.n1779 0.4505
R27203 DVSS.n8168 DVSS.n8167 0.4505
R27204 DVSS.n1938 DVSS.n1925 0.4505
R27205 DVSS.n1940 DVSS.n1939 0.4505
R27206 DVSS.n1936 DVSS.n1934 0.4505
R27207 DVSS.n8052 DVSS.n8051 0.4505
R27208 DVSS.n1937 DVSS.n1935 0.4505
R27209 DVSS.n8047 DVSS.n8046 0.4505
R27210 DVSS.n8045 DVSS.n1944 0.4505
R27211 DVSS.n8044 DVSS.n8043 0.4505
R27212 DVSS.n1949 DVSS.n1946 0.4505
R27213 DVSS.n8039 DVSS.n8038 0.4505
R27214 DVSS.n1956 DVSS.n1948 0.4505
R27215 DVSS.n8029 DVSS.n8028 0.4505
R27216 DVSS.n1968 DVSS.n1967 0.4505
R27217 DVSS.n8024 DVSS.n8023 0.4505
R27218 DVSS.n8022 DVSS.n1970 0.4505
R27219 DVSS.n8021 DVSS.n8020 0.4505
R27220 DVSS.n1975 DVSS.n1972 0.4505
R27221 DVSS.n8016 DVSS.n8015 0.4505
R27222 DVSS.n1982 DVSS.n1974 0.4505
R27223 DVSS.n8006 DVSS.n8005 0.4505
R27224 DVSS.n1994 DVSS.n1993 0.4505
R27225 DVSS.n8001 DVSS.n8000 0.4505
R27226 DVSS.n7999 DVSS.n1996 0.4505
R27227 DVSS.n7998 DVSS.n7997 0.4505
R27228 DVSS.n1998 DVSS.n1997 0.4505
R27229 DVSS.n7993 DVSS.n7992 0.4505
R27230 DVSS.n7991 DVSS.n2000 0.4505
R27231 DVSS.n7990 DVSS.n7989 0.4505
R27232 DVSS.n2002 DVSS.n2001 0.4505
R27233 DVSS.n7985 DVSS.n7984 0.4505
R27234 DVSS.n7983 DVSS.n2004 0.4505
R27235 DVSS.n7982 DVSS.n7981 0.4505
R27236 DVSS.n2009 DVSS.n2006 0.4505
R27237 DVSS.n7977 DVSS.n7976 0.4505
R27238 DVSS.n2016 DVSS.n2008 0.4505
R27239 DVSS.n7967 DVSS.n7966 0.4505
R27240 DVSS.n2028 DVSS.n2027 0.4505
R27241 DVSS.n7962 DVSS.n7961 0.4505
R27242 DVSS.n7960 DVSS.n2030 0.4505
R27243 DVSS.n7959 DVSS.n7958 0.4505
R27244 DVSS.n2032 DVSS.n2031 0.4505
R27245 DVSS.n7954 DVSS.n7953 0.4505
R27246 DVSS.n7952 DVSS.n2034 0.4505
R27247 DVSS.n7951 DVSS.n7950 0.4505
R27248 DVSS.n2036 DVSS.n2035 0.4505
R27249 DVSS.n7946 DVSS.n7945 0.4505
R27250 DVSS.n7944 DVSS.n2038 0.4505
R27251 DVSS.n7943 DVSS.n7942 0.4505
R27252 DVSS.n2043 DVSS.n2040 0.4505
R27253 DVSS.n7938 DVSS.n7937 0.4505
R27254 DVSS.n2050 DVSS.n2042 0.4505
R27255 DVSS.n7768 DVSS.n2062 0.4505
R27256 DVSS.n7769 DVSS.n2068 0.4505
R27257 DVSS.n7771 DVSS.n7770 0.4505
R27258 DVSS.n7765 DVSS.n7764 0.4505
R27259 DVSS.n7776 DVSS.n7775 0.4505
R27260 DVSS.n7777 DVSS.n7763 0.4505
R27261 DVSS.n7779 DVSS.n7778 0.4505
R27262 DVSS.n7761 DVSS.n7760 0.4505
R27263 DVSS.n7784 DVSS.n7783 0.4505
R27264 DVSS.n7785 DVSS.n7759 0.4505
R27265 DVSS.n7787 DVSS.n7786 0.4505
R27266 DVSS.n7757 DVSS.n7756 0.4505
R27267 DVSS.n7793 DVSS.n7792 0.4505
R27268 DVSS.n7794 DVSS.n7755 0.4505
R27269 DVSS.n7796 DVSS.n7795 0.4505
R27270 DVSS.n7797 DVSS.n7731 0.4505
R27271 DVSS.n7751 DVSS.n7737 0.4505
R27272 DVSS.n7843 DVSS.n7842 0.4505
R27273 DVSS.n7753 DVSS.n7752 0.4505
R27274 DVSS.n7838 DVSS.n7837 0.4505
R27275 DVSS.n7836 DVSS.n7801 0.4505
R27276 DVSS.n7835 DVSS.n7834 0.4505
R27277 DVSS.n7803 DVSS.n7802 0.4505
R27278 DVSS.n7830 DVSS.n7829 0.4505
R27279 DVSS.n7828 DVSS.n7805 0.4505
R27280 DVSS.n7827 DVSS.n7826 0.4505
R27281 DVSS.n7807 DVSS.n7806 0.4505
R27282 DVSS.n7822 DVSS.n7821 0.4505
R27283 DVSS.n7820 DVSS.n7809 0.4505
R27284 DVSS.n7819 DVSS.n7818 0.4505
R27285 DVSS.n7811 DVSS.n7810 0.4505
R27286 DVSS.n7814 DVSS.n1816 0.4505
R27287 DVSS.n7813 DVSS.n1822 0.4505
R27288 DVSS.n1831 DVSS.n1807 0.4505
R27289 DVSS.n8125 DVSS.n8124 0.4505
R27290 DVSS.n1805 DVSS.n1804 0.4505
R27291 DVSS.n8130 DVSS.n8129 0.4505
R27292 DVSS.n8131 DVSS.n1803 0.4505
R27293 DVSS.n8133 DVSS.n8132 0.4505
R27294 DVSS.n1801 DVSS.n1796 0.4505
R27295 DVSS.n8138 DVSS.n8137 0.4505
R27296 DVSS.n8144 DVSS.n1787 0.4505
R27297 DVSS.n8154 DVSS.n8153 0.4505
R27298 DVSS.n1785 DVSS.n1784 0.4505
R27299 DVSS.n8159 DVSS.n8158 0.4505
R27300 DVSS.n8160 DVSS.n1783 0.4505
R27301 DVSS.n8162 DVSS.n8161 0.4505
R27302 DVSS.n8165 DVSS.n1764 0.4505
R27303 DVSS.n8166 DVSS.n1770 0.4505
R27304 DVSS.n5099 DVSS.n5098 0.4505
R27305 DVSS.n3079 DVSS.n3076 0.4505
R27306 DVSS.n3082 DVSS.n3081 0.4505
R27307 DVSS.n3083 DVSS.n3075 0.4505
R27308 DVSS.n3086 DVSS.n3085 0.4505
R27309 DVSS.n3084 DVSS.n3073 0.4505
R27310 DVSS.n3090 DVSS.n3072 0.4505
R27311 DVSS.n3092 DVSS.n3091 0.4505
R27312 DVSS.n3093 DVSS.n3070 0.4505
R27313 DVSS.n5827 DVSS.n5826 0.4505
R27314 DVSS.n5825 DVSS.n3071 0.4505
R27315 DVSS.n5824 DVSS.n5823 0.4505
R27316 DVSS.n3095 DVSS.n3094 0.4505
R27317 DVSS.n5819 DVSS.n5818 0.4505
R27318 DVSS.n5817 DVSS.n3097 0.4505
R27319 DVSS.n5816 DVSS.n5815 0.4505
R27320 DVSS.n3099 DVSS.n3098 0.4505
R27321 DVSS.n3124 DVSS.n3123 0.4505
R27322 DVSS.n3125 DVSS.n3120 0.4505
R27323 DVSS.n5807 DVSS.n5806 0.4505
R27324 DVSS.n5805 DVSS.n3121 0.4505
R27325 DVSS.n5804 DVSS.n5803 0.4505
R27326 DVSS.n3127 DVSS.n3126 0.4505
R27327 DVSS.n5799 DVSS.n5798 0.4505
R27328 DVSS.n5797 DVSS.n3129 0.4505
R27329 DVSS.n5796 DVSS.n5795 0.4505
R27330 DVSS.n3131 DVSS.n3130 0.4505
R27331 DVSS.n5791 DVSS.n5790 0.4505
R27332 DVSS.n5789 DVSS.n3133 0.4505
R27333 DVSS.n5788 DVSS.n5787 0.4505
R27334 DVSS.n3135 DVSS.n3134 0.4505
R27335 DVSS.n5783 DVSS.n5782 0.4505
R27336 DVSS.n5781 DVSS.n3137 0.4505
R27337 DVSS.n5780 DVSS.n5779 0.4505
R27338 DVSS.n3139 DVSS.n3138 0.4505
R27339 DVSS.n5771 DVSS.n5770 0.4505
R27340 DVSS.n5769 DVSS.n3159 0.4505
R27341 DVSS.n5768 DVSS.n5767 0.4505
R27342 DVSS.n3161 DVSS.n3160 0.4505
R27343 DVSS.n5763 DVSS.n5762 0.4505
R27344 DVSS.n5761 DVSS.n3163 0.4505
R27345 DVSS.n5760 DVSS.n5759 0.4505
R27346 DVSS.n3165 DVSS.n3164 0.4505
R27347 DVSS.n5755 DVSS.n5754 0.4505
R27348 DVSS.n5753 DVSS.n3167 0.4505
R27349 DVSS.n5752 DVSS.n5751 0.4505
R27350 DVSS.n3169 DVSS.n3168 0.4505
R27351 DVSS.n5747 DVSS.n5746 0.4505
R27352 DVSS.n5745 DVSS.n3171 0.4505
R27353 DVSS.n5744 DVSS.n5743 0.4505
R27354 DVSS.n3173 DVSS.n3172 0.4505
R27355 DVSS.n5034 DVSS.n5033 0.4505
R27356 DVSS.n5035 DVSS.n5031 0.4505
R27357 DVSS.n5192 DVSS.n5191 0.4505
R27358 DVSS.n5190 DVSS.n5032 0.4505
R27359 DVSS.n5189 DVSS.n5188 0.4505
R27360 DVSS.n5037 DVSS.n5036 0.4505
R27361 DVSS.n5184 DVSS.n5183 0.4505
R27362 DVSS.n5182 DVSS.n5040 0.4505
R27363 DVSS.n5181 DVSS.n5180 0.4505
R27364 DVSS.n5042 DVSS.n5041 0.4505
R27365 DVSS.n5176 DVSS.n5175 0.4505
R27366 DVSS.n5174 DVSS.n5044 0.4505
R27367 DVSS.n5173 DVSS.n5172 0.4505
R27368 DVSS.n5046 DVSS.n5045 0.4505
R27369 DVSS.n5168 DVSS.n5167 0.4505
R27370 DVSS.n5166 DVSS.n5048 0.4505
R27371 DVSS.n5165 DVSS.n5164 0.4505
R27372 DVSS.n5162 DVSS.n5049 0.4505
R27373 DVSS.n5160 DVSS.n5159 0.4505
R27374 DVSS.n5158 DVSS.n5050 0.4505
R27375 DVSS.n5157 DVSS.n5156 0.4505
R27376 DVSS.n5052 DVSS.n5051 0.4505
R27377 DVSS.n5152 DVSS.n5151 0.4505
R27378 DVSS.n5150 DVSS.n5054 0.4505
R27379 DVSS.n5149 DVSS.n5148 0.4505
R27380 DVSS.n5056 DVSS.n5055 0.4505
R27381 DVSS.n5144 DVSS.n5143 0.4505
R27382 DVSS.n5142 DVSS.n5058 0.4505
R27383 DVSS.n5141 DVSS.n5140 0.4505
R27384 DVSS.n5060 DVSS.n5059 0.4505
R27385 DVSS.n5136 DVSS.n5135 0.4505
R27386 DVSS.n5134 DVSS.n5062 0.4505
R27387 DVSS.n5133 DVSS.n5132 0.4505
R27388 DVSS.n5064 DVSS.n5063 0.4505
R27389 DVSS.n5085 DVSS.n5083 0.4505
R27390 DVSS.n5126 DVSS.n5125 0.4505
R27391 DVSS.n5124 DVSS.n5084 0.4505
R27392 DVSS.n5123 DVSS.n5122 0.4505
R27393 DVSS.n5087 DVSS.n5086 0.4505
R27394 DVSS.n5118 DVSS.n5117 0.4505
R27395 DVSS.n5116 DVSS.n5089 0.4505
R27396 DVSS.n5115 DVSS.n5114 0.4505
R27397 DVSS.n5112 DVSS.n5090 0.4505
R27398 DVSS.n5111 DVSS.n5110 0.4505
R27399 DVSS.n5109 DVSS.n5091 0.4505
R27400 DVSS.n5108 DVSS.n5107 0.4505
R27401 DVSS.n5103 DVSS.n5092 0.4505
R27402 DVSS.n5102 DVSS.n5101 0.4505
R27403 DVSS.n5100 DVSS.n5093 0.4505
R27404 DVSS.n5096 DVSS.n5095 0.4505
R27405 DVSS.n5098 DVSS.n5097 0.4505
R27406 DVSS.n3077 DVSS.n3003 0.4505
R27407 DVSS.n3079 DVSS.n3078 0.4505
R27408 DVSS.n3081 DVSS.n3080 0.4505
R27409 DVSS.n3075 DVSS.n3074 0.4505
R27410 DVSS.n3087 DVSS.n3086 0.4505
R27411 DVSS.n3088 DVSS.n3073 0.4505
R27412 DVSS.n3090 DVSS.n3089 0.4505
R27413 DVSS.n3091 DVSS.n3056 0.4505
R27414 DVSS.n3070 DVSS.n3062 0.4505
R27415 DVSS.n5828 DVSS.n5827 0.4505
R27416 DVSS.n3071 DVSS.n3069 0.4505
R27417 DVSS.n5823 DVSS.n5822 0.4505
R27418 DVSS.n5821 DVSS.n3095 0.4505
R27419 DVSS.n5820 DVSS.n5819 0.4505
R27420 DVSS.n3097 DVSS.n3096 0.4505
R27421 DVSS.n5815 DVSS.n5814 0.4505
R27422 DVSS.n3105 DVSS.n3099 0.4505
R27423 DVSS.n3123 DVSS.n3122 0.4505
R27424 DVSS.n3120 DVSS.n3118 0.4505
R27425 DVSS.n5808 DVSS.n5807 0.4505
R27426 DVSS.n3121 DVSS.n3119 0.4505
R27427 DVSS.n5803 DVSS.n5802 0.4505
R27428 DVSS.n5801 DVSS.n3127 0.4505
R27429 DVSS.n5800 DVSS.n5799 0.4505
R27430 DVSS.n3129 DVSS.n3128 0.4505
R27431 DVSS.n5795 DVSS.n5794 0.4505
R27432 DVSS.n5793 DVSS.n3131 0.4505
R27433 DVSS.n5792 DVSS.n5791 0.4505
R27434 DVSS.n3133 DVSS.n3132 0.4505
R27435 DVSS.n5787 DVSS.n5786 0.4505
R27436 DVSS.n5785 DVSS.n3135 0.4505
R27437 DVSS.n5784 DVSS.n5783 0.4505
R27438 DVSS.n3140 DVSS.n3137 0.4505
R27439 DVSS.n5779 DVSS.n5778 0.4505
R27440 DVSS.n3147 DVSS.n3139 0.4505
R27441 DVSS.n5772 DVSS.n5771 0.4505
R27442 DVSS.n3159 DVSS.n3158 0.4505
R27443 DVSS.n5767 DVSS.n5766 0.4505
R27444 DVSS.n5765 DVSS.n3161 0.4505
R27445 DVSS.n5764 DVSS.n5763 0.4505
R27446 DVSS.n3163 DVSS.n3162 0.4505
R27447 DVSS.n5759 DVSS.n5758 0.4505
R27448 DVSS.n5757 DVSS.n3165 0.4505
R27449 DVSS.n5756 DVSS.n5755 0.4505
R27450 DVSS.n3167 DVSS.n3166 0.4505
R27451 DVSS.n5751 DVSS.n5750 0.4505
R27452 DVSS.n5749 DVSS.n3169 0.4505
R27453 DVSS.n5748 DVSS.n5747 0.4505
R27454 DVSS.n3174 DVSS.n3171 0.4505
R27455 DVSS.n5743 DVSS.n5742 0.4505
R27456 DVSS.n3181 DVSS.n3173 0.4505
R27457 DVSS.n5033 DVSS.n5011 0.4505
R27458 DVSS.n5031 DVSS.n5016 0.4505
R27459 DVSS.n5193 DVSS.n5192 0.4505
R27460 DVSS.n5038 DVSS.n5032 0.4505
R27461 DVSS.n5188 DVSS.n5187 0.4505
R27462 DVSS.n5186 DVSS.n5037 0.4505
R27463 DVSS.n5185 DVSS.n5184 0.4505
R27464 DVSS.n5040 DVSS.n5039 0.4505
R27465 DVSS.n5180 DVSS.n5179 0.4505
R27466 DVSS.n5178 DVSS.n5042 0.4505
R27467 DVSS.n5177 DVSS.n5176 0.4505
R27468 DVSS.n5044 DVSS.n5043 0.4505
R27469 DVSS.n5172 DVSS.n5171 0.4505
R27470 DVSS.n5170 DVSS.n5046 0.4505
R27471 DVSS.n5169 DVSS.n5168 0.4505
R27472 DVSS.n5048 DVSS.n5047 0.4505
R27473 DVSS.n5164 DVSS.n5163 0.4505
R27474 DVSS.n5162 DVSS.n5161 0.4505
R27475 DVSS.n5160 DVSS.n3328 0.4505
R27476 DVSS.n5050 DVSS.n3332 0.4505
R27477 DVSS.n5156 DVSS.n5155 0.4505
R27478 DVSS.n5154 DVSS.n5052 0.4505
R27479 DVSS.n5153 DVSS.n5152 0.4505
R27480 DVSS.n5054 DVSS.n5053 0.4505
R27481 DVSS.n5148 DVSS.n5147 0.4505
R27482 DVSS.n5146 DVSS.n5056 0.4505
R27483 DVSS.n5145 DVSS.n5144 0.4505
R27484 DVSS.n5058 DVSS.n5057 0.4505
R27485 DVSS.n5140 DVSS.n5139 0.4505
R27486 DVSS.n5138 DVSS.n5060 0.4505
R27487 DVSS.n5137 DVSS.n5136 0.4505
R27488 DVSS.n5062 DVSS.n5061 0.4505
R27489 DVSS.n5132 DVSS.n5131 0.4505
R27490 DVSS.n5068 DVSS.n5064 0.4505
R27491 DVSS.n5083 DVSS.n5074 0.4505
R27492 DVSS.n5127 DVSS.n5126 0.4505
R27493 DVSS.n5084 DVSS.n5082 0.4505
R27494 DVSS.n5122 DVSS.n5121 0.4505
R27495 DVSS.n5120 DVSS.n5087 0.4505
R27496 DVSS.n5119 DVSS.n5118 0.4505
R27497 DVSS.n5089 DVSS.n5088 0.4505
R27498 DVSS.n5114 DVSS.n5113 0.4505
R27499 DVSS.n5112 DVSS.n3374 0.4505
R27500 DVSS.n5111 DVSS.n3376 0.4505
R27501 DVSS.n5104 DVSS.n5091 0.4505
R27502 DVSS.n5107 DVSS.n5106 0.4505
R27503 DVSS.n5105 DVSS.n5103 0.4505
R27504 DVSS.n5102 DVSS.n2943 0.4505
R27505 DVSS.n5093 DVSS.n2949 0.4505
R27506 DVSS.n5335 DVSS.n5334 0.4505
R27507 DVSS.n5852 DVSS.n5850 0.4505
R27508 DVSS.n5849 DVSS.n3036 0.4505
R27509 DVSS.n5848 DVSS.n5847 0.4505
R27510 DVSS.n3038 DVSS.n3037 0.4505
R27511 DVSS.n5843 DVSS.n5842 0.4505
R27512 DVSS.n5841 DVSS.n3040 0.4505
R27513 DVSS.n5840 DVSS.n5839 0.4505
R27514 DVSS.n3042 DVSS.n3041 0.4505
R27515 DVSS.n3903 DVSS.n3902 0.4505
R27516 DVSS.n3906 DVSS.n3905 0.4505
R27517 DVSS.n3907 DVSS.n3901 0.4505
R27518 DVSS.n3909 DVSS.n3908 0.4505
R27519 DVSS.n3899 DVSS.n3898 0.4505
R27520 DVSS.n3914 DVSS.n3913 0.4505
R27521 DVSS.n3915 DVSS.n3895 0.4505
R27522 DVSS.n4171 DVSS.n4170 0.4505
R27523 DVSS.n4169 DVSS.n3897 0.4505
R27524 DVSS.n4168 DVSS.n4167 0.4505
R27525 DVSS.n4165 DVSS.n3916 0.4505
R27526 DVSS.n3920 DVSS.n3917 0.4505
R27527 DVSS.n4161 DVSS.n4160 0.4505
R27528 DVSS.n4159 DVSS.n3919 0.4505
R27529 DVSS.n4158 DVSS.n4157 0.4505
R27530 DVSS.n3922 DVSS.n3921 0.4505
R27531 DVSS.n4153 DVSS.n4152 0.4505
R27532 DVSS.n4151 DVSS.n3924 0.4505
R27533 DVSS.n4150 DVSS.n4149 0.4505
R27534 DVSS.n3926 DVSS.n3925 0.4505
R27535 DVSS.n4145 DVSS.n4144 0.4505
R27536 DVSS.n4143 DVSS.n3928 0.4505
R27537 DVSS.n4142 DVSS.n4141 0.4505
R27538 DVSS.n3930 DVSS.n3929 0.4505
R27539 DVSS.n3953 DVSS.n3951 0.4505
R27540 DVSS.n4135 DVSS.n4134 0.4505
R27541 DVSS.n4133 DVSS.n3952 0.4505
R27542 DVSS.n4132 DVSS.n4131 0.4505
R27543 DVSS.n3955 DVSS.n3954 0.4505
R27544 DVSS.n4127 DVSS.n4126 0.4505
R27545 DVSS.n4125 DVSS.n3958 0.4505
R27546 DVSS.n4124 DVSS.n4123 0.4505
R27547 DVSS.n3960 DVSS.n3959 0.4505
R27548 DVSS.n4119 DVSS.n4118 0.4505
R27549 DVSS.n4117 DVSS.n3962 0.4505
R27550 DVSS.n4116 DVSS.n4115 0.4505
R27551 DVSS.n3964 DVSS.n3963 0.4505
R27552 DVSS.n4111 DVSS.n4110 0.4505
R27553 DVSS.n4109 DVSS.n3966 0.4505
R27554 DVSS.n4108 DVSS.n4107 0.4505
R27555 DVSS.n3968 DVSS.n3967 0.4505
R27556 DVSS.n3996 DVSS.n3995 0.4505
R27557 DVSS.n3473 DVSS.n3472 0.4505
R27558 DVSS.n5240 DVSS.n5239 0.4505
R27559 DVSS.n5241 DVSS.n3471 0.4505
R27560 DVSS.n5243 DVSS.n5242 0.4505
R27561 DVSS.n3469 DVSS.n3468 0.4505
R27562 DVSS.n5248 DVSS.n5247 0.4505
R27563 DVSS.n5249 DVSS.n3467 0.4505
R27564 DVSS.n5251 DVSS.n5250 0.4505
R27565 DVSS.n3465 DVSS.n3464 0.4505
R27566 DVSS.n5256 DVSS.n5255 0.4505
R27567 DVSS.n5257 DVSS.n3463 0.4505
R27568 DVSS.n5259 DVSS.n5258 0.4505
R27569 DVSS.n3461 DVSS.n3460 0.4505
R27570 DVSS.n5264 DVSS.n5263 0.4505
R27571 DVSS.n5265 DVSS.n3459 0.4505
R27572 DVSS.n5267 DVSS.n5266 0.4505
R27573 DVSS.n3439 DVSS.n3438 0.4505
R27574 DVSS.n5275 DVSS.n5274 0.4505
R27575 DVSS.n5276 DVSS.n3437 0.4505
R27576 DVSS.n5278 DVSS.n5277 0.4505
R27577 DVSS.n3435 DVSS.n3434 0.4505
R27578 DVSS.n5283 DVSS.n5282 0.4505
R27579 DVSS.n5284 DVSS.n3433 0.4505
R27580 DVSS.n5286 DVSS.n5285 0.4505
R27581 DVSS.n3431 DVSS.n3430 0.4505
R27582 DVSS.n5291 DVSS.n5290 0.4505
R27583 DVSS.n5292 DVSS.n3429 0.4505
R27584 DVSS.n5294 DVSS.n5293 0.4505
R27585 DVSS.n3427 DVSS.n3426 0.4505
R27586 DVSS.n5299 DVSS.n5298 0.4505
R27587 DVSS.n5300 DVSS.n3425 0.4505
R27588 DVSS.n5302 DVSS.n5301 0.4505
R27589 DVSS.n3404 DVSS.n3403 0.4505
R27590 DVSS.n5310 DVSS.n5309 0.4505
R27591 DVSS.n5311 DVSS.n3402 0.4505
R27592 DVSS.n5313 DVSS.n5312 0.4505
R27593 DVSS.n3400 DVSS.n3399 0.4505
R27594 DVSS.n5319 DVSS.n5318 0.4505
R27595 DVSS.n5320 DVSS.n3398 0.4505
R27596 DVSS.n5322 DVSS.n5321 0.4505
R27597 DVSS.n5323 DVSS.n3397 0.4505
R27598 DVSS.n5326 DVSS.n5325 0.4505
R27599 DVSS.n5327 DVSS.n3395 0.4505
R27600 DVSS.n5346 DVSS.n5345 0.4505
R27601 DVSS.n5344 DVSS.n3396 0.4505
R27602 DVSS.n5343 DVSS.n5342 0.4505
R27603 DVSS.n5339 DVSS.n5328 0.4505
R27604 DVSS.n5338 DVSS.n5337 0.4505
R27605 DVSS.n5336 DVSS.n5329 0.4505
R27606 DVSS.n5332 DVSS.n5331 0.4505
R27607 DVSS.n5334 DVSS.n5333 0.4505
R27608 DVSS.n5854 DVSS.n5853 0.4505
R27609 DVSS.n5852 DVSS.n5851 0.4505
R27610 DVSS.n3036 DVSS.n3035 0.4505
R27611 DVSS.n5847 DVSS.n5846 0.4505
R27612 DVSS.n5845 DVSS.n3038 0.4505
R27613 DVSS.n5844 DVSS.n5843 0.4505
R27614 DVSS.n3040 DVSS.n3039 0.4505
R27615 DVSS.n5839 DVSS.n5838 0.4505
R27616 DVSS.n3048 DVSS.n3042 0.4505
R27617 DVSS.n3903 DVSS.n3054 0.4505
R27618 DVSS.n3905 DVSS.n3904 0.4505
R27619 DVSS.n3901 DVSS.n3900 0.4505
R27620 DVSS.n3910 DVSS.n3909 0.4505
R27621 DVSS.n3911 DVSS.n3899 0.4505
R27622 DVSS.n3913 DVSS.n3912 0.4505
R27623 DVSS.n3895 DVSS.n3890 0.4505
R27624 DVSS.n4172 DVSS.n4171 0.4505
R27625 DVSS.n3897 DVSS.n3896 0.4505
R27626 DVSS.n4167 DVSS.n4166 0.4505
R27627 DVSS.n4165 DVSS.n4164 0.4505
R27628 DVSS.n4163 DVSS.n3917 0.4505
R27629 DVSS.n4162 DVSS.n4161 0.4505
R27630 DVSS.n3919 DVSS.n3918 0.4505
R27631 DVSS.n4157 DVSS.n4156 0.4505
R27632 DVSS.n4155 DVSS.n3922 0.4505
R27633 DVSS.n4154 DVSS.n4153 0.4505
R27634 DVSS.n3924 DVSS.n3923 0.4505
R27635 DVSS.n4149 DVSS.n4148 0.4505
R27636 DVSS.n4147 DVSS.n3926 0.4505
R27637 DVSS.n4146 DVSS.n4145 0.4505
R27638 DVSS.n3928 DVSS.n3927 0.4505
R27639 DVSS.n4141 DVSS.n4140 0.4505
R27640 DVSS.n3936 DVSS.n3930 0.4505
R27641 DVSS.n3951 DVSS.n3947 0.4505
R27642 DVSS.n4136 DVSS.n4135 0.4505
R27643 DVSS.n3956 DVSS.n3952 0.4505
R27644 DVSS.n4131 DVSS.n4130 0.4505
R27645 DVSS.n4129 DVSS.n3955 0.4505
R27646 DVSS.n4128 DVSS.n4127 0.4505
R27647 DVSS.n3958 DVSS.n3957 0.4505
R27648 DVSS.n4123 DVSS.n4122 0.4505
R27649 DVSS.n4121 DVSS.n3960 0.4505
R27650 DVSS.n4120 DVSS.n4119 0.4505
R27651 DVSS.n3962 DVSS.n3961 0.4505
R27652 DVSS.n4115 DVSS.n4114 0.4505
R27653 DVSS.n4113 DVSS.n3964 0.4505
R27654 DVSS.n4112 DVSS.n4111 0.4505
R27655 DVSS.n3966 DVSS.n3965 0.4505
R27656 DVSS.n4107 DVSS.n4106 0.4505
R27657 DVSS.n3976 DVSS.n3968 0.4505
R27658 DVSS.n3997 DVSS.n3996 0.4505
R27659 DVSS.n3994 DVSS.n3473 0.4505
R27660 DVSS.n5239 DVSS.n5238 0.4505
R27661 DVSS.n3480 DVSS.n3471 0.4505
R27662 DVSS.n5244 DVSS.n5243 0.4505
R27663 DVSS.n5245 DVSS.n3469 0.4505
R27664 DVSS.n5247 DVSS.n5246 0.4505
R27665 DVSS.n3467 DVSS.n3466 0.4505
R27666 DVSS.n5252 DVSS.n5251 0.4505
R27667 DVSS.n5253 DVSS.n3465 0.4505
R27668 DVSS.n5255 DVSS.n5254 0.4505
R27669 DVSS.n3463 DVSS.n3462 0.4505
R27670 DVSS.n5260 DVSS.n5259 0.4505
R27671 DVSS.n5261 DVSS.n3461 0.4505
R27672 DVSS.n5263 DVSS.n5262 0.4505
R27673 DVSS.n3459 DVSS.n3458 0.4505
R27674 DVSS.n5268 DVSS.n5267 0.4505
R27675 DVSS.n5269 DVSS.n3439 0.4505
R27676 DVSS.n5274 DVSS.n5273 0.4505
R27677 DVSS.n3446 DVSS.n3437 0.4505
R27678 DVSS.n5279 DVSS.n5278 0.4505
R27679 DVSS.n5280 DVSS.n3435 0.4505
R27680 DVSS.n5282 DVSS.n5281 0.4505
R27681 DVSS.n3433 DVSS.n3432 0.4505
R27682 DVSS.n5287 DVSS.n5286 0.4505
R27683 DVSS.n5288 DVSS.n3431 0.4505
R27684 DVSS.n5290 DVSS.n5289 0.4505
R27685 DVSS.n3429 DVSS.n3428 0.4505
R27686 DVSS.n5295 DVSS.n5294 0.4505
R27687 DVSS.n5296 DVSS.n3427 0.4505
R27688 DVSS.n5298 DVSS.n5297 0.4505
R27689 DVSS.n3425 DVSS.n3424 0.4505
R27690 DVSS.n5303 DVSS.n5302 0.4505
R27691 DVSS.n5304 DVSS.n3404 0.4505
R27692 DVSS.n5309 DVSS.n5308 0.4505
R27693 DVSS.n3411 DVSS.n3402 0.4505
R27694 DVSS.n5314 DVSS.n5313 0.4505
R27695 DVSS.n5315 DVSS.n3400 0.4505
R27696 DVSS.n5318 DVSS.n5317 0.4505
R27697 DVSS.n5316 DVSS.n3398 0.4505
R27698 DVSS.n5322 DVSS.n3380 0.4505
R27699 DVSS.n5323 DVSS.n3386 0.4505
R27700 DVSS.n5325 DVSS.n5324 0.4505
R27701 DVSS.n3395 DVSS.n3393 0.4505
R27702 DVSS.n5347 DVSS.n5346 0.4505
R27703 DVSS.n3396 DVSS.n3394 0.4505
R27704 DVSS.n5342 DVSS.n5341 0.4505
R27705 DVSS.n5340 DVSS.n5339 0.4505
R27706 DVSS.n5338 DVSS.n2925 0.4505
R27707 DVSS.n5329 DVSS.n2931 0.4505
R27708 DVSS.n4941 DVSS.n4940 0.4505
R27709 DVSS.n4936 DVSS.n4935 0.4505
R27710 DVSS.n4235 DVSS.n3845 0.4505
R27711 DVSS.n4237 DVSS.n4236 0.4505
R27712 DVSS.n4239 DVSS.n4238 0.4505
R27713 DVSS.n4233 DVSS.n4232 0.4505
R27714 DVSS.n4244 DVSS.n4243 0.4505
R27715 DVSS.n4245 DVSS.n4231 0.4505
R27716 DVSS.n4247 DVSS.n4246 0.4505
R27717 DVSS.n4229 DVSS.n4224 0.4505
R27718 DVSS.n4252 DVSS.n4251 0.4505
R27719 DVSS.n4222 DVSS.n4214 0.4505
R27720 DVSS.n4262 DVSS.n4261 0.4505
R27721 DVSS.n4212 DVSS.n4211 0.4505
R27722 DVSS.n4267 DVSS.n4266 0.4505
R27723 DVSS.n4268 DVSS.n4210 0.4505
R27724 DVSS.n4270 DVSS.n4269 0.4505
R27725 DVSS.n4206 DVSS.n4202 0.4505
R27726 DVSS.n4418 DVSS.n4417 0.4505
R27727 DVSS.n4208 DVSS.n4207 0.4505
R27728 DVSS.n4413 DVSS.n4412 0.4505
R27729 DVSS.n4411 DVSS.n4410 0.4505
R27730 DVSS.n4409 DVSS.n4274 0.4505
R27731 DVSS.n4408 DVSS.n4407 0.4505
R27732 DVSS.n4276 DVSS.n4275 0.4505
R27733 DVSS.n4403 DVSS.n4402 0.4505
R27734 DVSS.n4401 DVSS.n4279 0.4505
R27735 DVSS.n4400 DVSS.n4399 0.4505
R27736 DVSS.n4281 DVSS.n4280 0.4505
R27737 DVSS.n4395 DVSS.n4394 0.4505
R27738 DVSS.n4393 DVSS.n4283 0.4505
R27739 DVSS.n4392 DVSS.n4391 0.4505
R27740 DVSS.n4285 DVSS.n4284 0.4505
R27741 DVSS.n4387 DVSS.n3722 0.4505
R27742 DVSS.n4386 DVSS.n3726 0.4505
R27743 DVSS.n4385 DVSS.n4384 0.4505
R27744 DVSS.n4288 DVSS.n4287 0.4505
R27745 DVSS.n4380 DVSS.n4379 0.4505
R27746 DVSS.n4378 DVSS.n4290 0.4505
R27747 DVSS.n4377 DVSS.n4376 0.4505
R27748 DVSS.n4292 DVSS.n4291 0.4505
R27749 DVSS.n4372 DVSS.n4371 0.4505
R27750 DVSS.n4370 DVSS.n4294 0.4505
R27751 DVSS.n4369 DVSS.n4368 0.4505
R27752 DVSS.n4296 DVSS.n4295 0.4505
R27753 DVSS.n4364 DVSS.n4363 0.4505
R27754 DVSS.n4362 DVSS.n4298 0.4505
R27755 DVSS.n4361 DVSS.n4360 0.4505
R27756 DVSS.n4300 DVSS.n4299 0.4505
R27757 DVSS.n4356 DVSS.n3691 0.4505
R27758 DVSS.n4355 DVSS.n3697 0.4505
R27759 DVSS.n4354 DVSS.n4353 0.4505
R27760 DVSS.n4303 DVSS.n4302 0.4505
R27761 DVSS.n4349 DVSS.n3679 0.4505
R27762 DVSS.n4348 DVSS.n3683 0.4505
R27763 DVSS.n4347 DVSS.n4346 0.4505
R27764 DVSS.n4308 DVSS.n4305 0.4505
R27765 DVSS.n4342 DVSS.n4341 0.4505
R27766 DVSS.n4340 DVSS.n4307 0.4505
R27767 DVSS.n4339 DVSS.n4338 0.4505
R27768 DVSS.n4310 DVSS.n4309 0.4505
R27769 DVSS.n4334 DVSS.n4333 0.4505
R27770 DVSS.n4332 DVSS.n4312 0.4505
R27771 DVSS.n4331 DVSS.n4330 0.4505
R27772 DVSS.n4314 DVSS.n4313 0.4505
R27773 DVSS.n4326 DVSS.n4325 0.4505
R27774 DVSS.n4324 DVSS.n4316 0.4505
R27775 DVSS.n4323 DVSS.n4322 0.4505
R27776 DVSS.n4317 DVSS.n3656 0.4505
R27777 DVSS.n4318 DVSS.n3660 0.4505
R27778 DVSS.n3665 DVSS.n3646 0.4505
R27779 DVSS.n4852 DVSS.n4851 0.4505
R27780 DVSS.n3644 DVSS.n3643 0.4505
R27781 DVSS.n4857 DVSS.n4856 0.4505
R27782 DVSS.n4858 DVSS.n3642 0.4505
R27783 DVSS.n4860 DVSS.n4859 0.4505
R27784 DVSS.n3640 DVSS.n3639 0.4505
R27785 DVSS.n4865 DVSS.n4864 0.4505
R27786 DVSS.n4866 DVSS.n3638 0.4505
R27787 DVSS.n4868 DVSS.n4867 0.4505
R27788 DVSS.n3636 DVSS.n3635 0.4505
R27789 DVSS.n4873 DVSS.n4872 0.4505
R27790 DVSS.n4874 DVSS.n3634 0.4505
R27791 DVSS.n4876 DVSS.n4875 0.4505
R27792 DVSS.n3632 DVSS.n3627 0.4505
R27793 DVSS.n4881 DVSS.n4880 0.4505
R27794 DVSS.n3624 DVSS.n3613 0.4505
R27795 DVSS.n4890 DVSS.n4889 0.4505
R27796 DVSS.n3611 DVSS.n3610 0.4505
R27797 DVSS.n4895 DVSS.n4894 0.4505
R27798 DVSS.n4896 DVSS.n3609 0.4505
R27799 DVSS.n4898 DVSS.n4897 0.4505
R27800 DVSS.n3605 DVSS.n3601 0.4505
R27801 DVSS.n4961 DVSS.n4960 0.4505
R27802 DVSS.n3607 DVSS.n3606 0.4505
R27803 DVSS.n4956 DVSS.n4955 0.4505
R27804 DVSS.n4954 DVSS.n4953 0.4505
R27805 DVSS.n4952 DVSS.n4902 0.4505
R27806 DVSS.n4951 DVSS.n4950 0.4505
R27807 DVSS.n4904 DVSS.n4903 0.4505
R27808 DVSS.n4946 DVSS.n4945 0.4505
R27809 DVSS.n4912 DVSS.n4906 0.4505
R27810 DVSS.n6619 DVSS.n6618 0.4505
R27811 DVSS.n6031 DVSS.n6030 0.4505
R27812 DVSS.n6614 DVSS.n6613 0.4505
R27813 DVSS.n6612 DVSS.n6349 0.4505
R27814 DVSS.n6611 DVSS.n6610 0.4505
R27815 DVSS.n6351 DVSS.n6350 0.4505
R27816 DVSS.n6606 DVSS.n6605 0.4505
R27817 DVSS.n6604 DVSS.n6353 0.4505
R27818 DVSS.n6603 DVSS.n6602 0.4505
R27819 DVSS.n6355 DVSS.n6354 0.4505
R27820 DVSS.n6598 DVSS.n6597 0.4505
R27821 DVSS.n6596 DVSS.n6357 0.4505
R27822 DVSS.n6595 DVSS.n6594 0.4505
R27823 DVSS.n6359 DVSS.n6358 0.4505
R27824 DVSS.n6590 DVSS.n6589 0.4505
R27825 DVSS.n6588 DVSS.n6361 0.4505
R27826 DVSS.n6587 DVSS.n6586 0.4505
R27827 DVSS.n6363 DVSS.n6362 0.4505
R27828 DVSS.n6582 DVSS.n6581 0.4505
R27829 DVSS.n6580 DVSS.n6365 0.4505
R27830 DVSS.n6579 DVSS.n6578 0.4505
R27831 DVSS.n6367 DVSS.n6366 0.4505
R27832 DVSS.n6574 DVSS.n6573 0.4505
R27833 DVSS.n6572 DVSS.n6369 0.4505
R27834 DVSS.n6571 DVSS.n6570 0.4505
R27835 DVSS.n6371 DVSS.n6370 0.4505
R27836 DVSS.n6566 DVSS.n6565 0.4505
R27837 DVSS.n6564 DVSS.n6373 0.4505
R27838 DVSS.n6563 DVSS.n6562 0.4505
R27839 DVSS.n6375 DVSS.n6374 0.4505
R27840 DVSS.n6558 DVSS.n6557 0.4505
R27841 DVSS.n6556 DVSS.n6377 0.4505
R27842 DVSS.n6555 DVSS.n6554 0.4505
R27843 DVSS.n6379 DVSS.n6378 0.4505
R27844 DVSS.n6550 DVSS.n6549 0.4505
R27845 DVSS.n6548 DVSS.n6381 0.4505
R27846 DVSS.n6547 DVSS.n6546 0.4505
R27847 DVSS.n6383 DVSS.n6382 0.4505
R27848 DVSS.n6542 DVSS.n6541 0.4505
R27849 DVSS.n6540 DVSS.n6385 0.4505
R27850 DVSS.n6539 DVSS.n6538 0.4505
R27851 DVSS.n6387 DVSS.n6386 0.4505
R27852 DVSS.n6534 DVSS.n6533 0.4505
R27853 DVSS.n6532 DVSS.n6389 0.4505
R27854 DVSS.n6531 DVSS.n6530 0.4505
R27855 DVSS.n6391 DVSS.n6390 0.4505
R27856 DVSS.n6526 DVSS.n6525 0.4505
R27857 DVSS.n6524 DVSS.n6393 0.4505
R27858 DVSS.n6523 DVSS.n6522 0.4505
R27859 DVSS.n6395 DVSS.n6394 0.4505
R27860 DVSS.n6518 DVSS.n6517 0.4505
R27861 DVSS.n6516 DVSS.n6397 0.4505
R27862 DVSS.n6515 DVSS.n6514 0.4505
R27863 DVSS.n6399 DVSS.n6398 0.4505
R27864 DVSS.n6510 DVSS.n6509 0.4505
R27865 DVSS.n6508 DVSS.n6401 0.4505
R27866 DVSS.n6507 DVSS.n6506 0.4505
R27867 DVSS.n6403 DVSS.n6402 0.4505
R27868 DVSS.n6502 DVSS.n6501 0.4505
R27869 DVSS.n6500 DVSS.n6405 0.4505
R27870 DVSS.n6499 DVSS.n6498 0.4505
R27871 DVSS.n6407 DVSS.n6406 0.4505
R27872 DVSS.n6494 DVSS.n6493 0.4505
R27873 DVSS.n6492 DVSS.n6409 0.4505
R27874 DVSS.n6491 DVSS.n6490 0.4505
R27875 DVSS.n6411 DVSS.n6410 0.4505
R27876 DVSS.n6486 DVSS.n6485 0.4505
R27877 DVSS.n6484 DVSS.n6413 0.4505
R27878 DVSS.n6483 DVSS.n6482 0.4505
R27879 DVSS.n6415 DVSS.n6414 0.4505
R27880 DVSS.n6478 DVSS.n6477 0.4505
R27881 DVSS.n6476 DVSS.n6417 0.4505
R27882 DVSS.n6475 DVSS.n6474 0.4505
R27883 DVSS.n6419 DVSS.n6418 0.4505
R27884 DVSS.n6470 DVSS.n6469 0.4505
R27885 DVSS.n6468 DVSS.n6421 0.4505
R27886 DVSS.n6467 DVSS.n6466 0.4505
R27887 DVSS.n6423 DVSS.n6422 0.4505
R27888 DVSS.n6462 DVSS.n6461 0.4505
R27889 DVSS.n6460 DVSS.n6425 0.4505
R27890 DVSS.n6459 DVSS.n6458 0.4505
R27891 DVSS.n6427 DVSS.n6426 0.4505
R27892 DVSS.n6454 DVSS.n6453 0.4505
R27893 DVSS.n6452 DVSS.n6429 0.4505
R27894 DVSS.n6451 DVSS.n6450 0.4505
R27895 DVSS.n6431 DVSS.n6430 0.4505
R27896 DVSS.n6446 DVSS.n6445 0.4505
R27897 DVSS.n6444 DVSS.n6443 0.4505
R27898 DVSS.n6435 DVSS.n6432 0.4505
R27899 DVSS.n6439 DVSS.n6438 0.4505
R27900 DVSS.n6638 DVSS.n6637 0.4505
R27901 DVSS.n6636 DVSS.n6020 0.4505
R27902 DVSS.n6635 DVSS.n6634 0.4505
R27903 DVSS.n6022 DVSS.n6021 0.4505
R27904 DVSS.n6630 DVSS.n6629 0.4505
R27905 DVSS.n6628 DVSS.n6025 0.4505
R27906 DVSS.n6627 DVSS.n6626 0.4505
R27907 DVSS.n6027 DVSS.n6026 0.4505
R27908 DVSS.n6622 DVSS.n6621 0.4505
R27909 DVSS.n6620 DVSS.n6029 0.4505
R27910 DVSS.n6340 DVSS.n6036 0.4505
R27911 DVSS.n6339 DVSS.n6338 0.4505
R27912 DVSS.n6067 DVSS.n6066 0.4505
R27913 DVSS.n6334 DVSS.n6333 0.4505
R27914 DVSS.n6332 DVSS.n6070 0.4505
R27915 DVSS.n6331 DVSS.n6330 0.4505
R27916 DVSS.n6072 DVSS.n6071 0.4505
R27917 DVSS.n6326 DVSS.n6325 0.4505
R27918 DVSS.n6324 DVSS.n6074 0.4505
R27919 DVSS.n6323 DVSS.n6322 0.4505
R27920 DVSS.n6076 DVSS.n6075 0.4505
R27921 DVSS.n6318 DVSS.n6317 0.4505
R27922 DVSS.n6316 DVSS.n6078 0.4505
R27923 DVSS.n6315 DVSS.n6314 0.4505
R27924 DVSS.n6080 DVSS.n6079 0.4505
R27925 DVSS.n6310 DVSS.n6309 0.4505
R27926 DVSS.n6308 DVSS.n6082 0.4505
R27927 DVSS.n6307 DVSS.n6306 0.4505
R27928 DVSS.n6084 DVSS.n6083 0.4505
R27929 DVSS.n6302 DVSS.n6301 0.4505
R27930 DVSS.n6300 DVSS.n6086 0.4505
R27931 DVSS.n6299 DVSS.n6298 0.4505
R27932 DVSS.n6088 DVSS.n6087 0.4505
R27933 DVSS.n6294 DVSS.n6293 0.4505
R27934 DVSS.n6292 DVSS.n6090 0.4505
R27935 DVSS.n6291 DVSS.n6290 0.4505
R27936 DVSS.n6092 DVSS.n6091 0.4505
R27937 DVSS.n6286 DVSS.n6285 0.4505
R27938 DVSS.n6284 DVSS.n6094 0.4505
R27939 DVSS.n6283 DVSS.n6282 0.4505
R27940 DVSS.n6096 DVSS.n6095 0.4505
R27941 DVSS.n6278 DVSS.n6277 0.4505
R27942 DVSS.n6276 DVSS.n6098 0.4505
R27943 DVSS.n6275 DVSS.n6274 0.4505
R27944 DVSS.n6100 DVSS.n6099 0.4505
R27945 DVSS.n6270 DVSS.n6269 0.4505
R27946 DVSS.n6268 DVSS.n6102 0.4505
R27947 DVSS.n6267 DVSS.n6266 0.4505
R27948 DVSS.n6104 DVSS.n6103 0.4505
R27949 DVSS.n6262 DVSS.n6261 0.4505
R27950 DVSS.n6260 DVSS.n6106 0.4505
R27951 DVSS.n6259 DVSS.n6258 0.4505
R27952 DVSS.n6108 DVSS.n6107 0.4505
R27953 DVSS.n6254 DVSS.n6253 0.4505
R27954 DVSS.n6252 DVSS.n6110 0.4505
R27955 DVSS.n6251 DVSS.n6250 0.4505
R27956 DVSS.n6112 DVSS.n6111 0.4505
R27957 DVSS.n6246 DVSS.n6245 0.4505
R27958 DVSS.n6244 DVSS.n6114 0.4505
R27959 DVSS.n6243 DVSS.n6242 0.4505
R27960 DVSS.n6116 DVSS.n6115 0.4505
R27961 DVSS.n6238 DVSS.n6237 0.4505
R27962 DVSS.n6236 DVSS.n6118 0.4505
R27963 DVSS.n6235 DVSS.n6234 0.4505
R27964 DVSS.n6120 DVSS.n6119 0.4505
R27965 DVSS.n6230 DVSS.n6229 0.4505
R27966 DVSS.n6228 DVSS.n6122 0.4505
R27967 DVSS.n6227 DVSS.n6226 0.4505
R27968 DVSS.n6124 DVSS.n6123 0.4505
R27969 DVSS.n6222 DVSS.n6221 0.4505
R27970 DVSS.n6220 DVSS.n6126 0.4505
R27971 DVSS.n6219 DVSS.n6218 0.4505
R27972 DVSS.n6128 DVSS.n6127 0.4505
R27973 DVSS.n6214 DVSS.n6213 0.4505
R27974 DVSS.n6212 DVSS.n6130 0.4505
R27975 DVSS.n6211 DVSS.n6210 0.4505
R27976 DVSS.n6132 DVSS.n6131 0.4505
R27977 DVSS.n6206 DVSS.n6205 0.4505
R27978 DVSS.n6204 DVSS.n6134 0.4505
R27979 DVSS.n6203 DVSS.n6202 0.4505
R27980 DVSS.n6136 DVSS.n6135 0.4505
R27981 DVSS.n6198 DVSS.n6197 0.4505
R27982 DVSS.n6196 DVSS.n6138 0.4505
R27983 DVSS.n6195 DVSS.n6194 0.4505
R27984 DVSS.n6140 DVSS.n6139 0.4505
R27985 DVSS.n6190 DVSS.n6189 0.4505
R27986 DVSS.n6188 DVSS.n6142 0.4505
R27987 DVSS.n6187 DVSS.n6186 0.4505
R27988 DVSS.n6144 DVSS.n6143 0.4505
R27989 DVSS.n6182 DVSS.n6181 0.4505
R27990 DVSS.n6180 DVSS.n6146 0.4505
R27991 DVSS.n6179 DVSS.n6178 0.4505
R27992 DVSS.n6148 DVSS.n6147 0.4505
R27993 DVSS.n6174 DVSS.n6173 0.4505
R27994 DVSS.n6172 DVSS.n6150 0.4505
R27995 DVSS.n6171 DVSS.n6170 0.4505
R27996 DVSS.n6152 DVSS.n6151 0.4505
R27997 DVSS.n6166 DVSS.n6165 0.4505
R27998 DVSS.n6164 DVSS.n6154 0.4505
R27999 DVSS.n6163 DVSS.n6162 0.4505
R28000 DVSS.n6049 DVSS.n6044 0.4505
R28001 DVSS.n6051 DVSS.n6050 0.4505
R28002 DVSS.n6042 DVSS.n6041 0.4505
R28003 DVSS.n6056 DVSS.n6055 0.4505
R28004 DVSS.n6057 DVSS.n6040 0.4505
R28005 DVSS.n6059 DVSS.n6058 0.4505
R28006 DVSS.n6038 DVSS.n6037 0.4505
R28007 DVSS.n6064 DVSS.n6063 0.4505
R28008 DVSS.n6065 DVSS.n6035 0.4505
R28009 DVSS.n6342 DVSS.n6341 0.4505
R28010 DVSS.n6160 DVSS.n6156 0.4505
R28011 DVSS.n6162 DVSS.n6161 0.4505
R28012 DVSS.n6154 DVSS.n6153 0.4505
R28013 DVSS.n6167 DVSS.n6166 0.4505
R28014 DVSS.n6168 DVSS.n6152 0.4505
R28015 DVSS.n6170 DVSS.n6169 0.4505
R28016 DVSS.n6150 DVSS.n6149 0.4505
R28017 DVSS.n6175 DVSS.n6174 0.4505
R28018 DVSS.n6176 DVSS.n6148 0.4505
R28019 DVSS.n6178 DVSS.n6177 0.4505
R28020 DVSS.n6146 DVSS.n6145 0.4505
R28021 DVSS.n6183 DVSS.n6182 0.4505
R28022 DVSS.n6184 DVSS.n6144 0.4505
R28023 DVSS.n6186 DVSS.n6185 0.4505
R28024 DVSS.n6142 DVSS.n6141 0.4505
R28025 DVSS.n6191 DVSS.n6190 0.4505
R28026 DVSS.n6192 DVSS.n6140 0.4505
R28027 DVSS.n6194 DVSS.n6193 0.4505
R28028 DVSS.n6138 DVSS.n6137 0.4505
R28029 DVSS.n6199 DVSS.n6198 0.4505
R28030 DVSS.n6200 DVSS.n6136 0.4505
R28031 DVSS.n6202 DVSS.n6201 0.4505
R28032 DVSS.n6134 DVSS.n6133 0.4505
R28033 DVSS.n6207 DVSS.n6206 0.4505
R28034 DVSS.n6208 DVSS.n6132 0.4505
R28035 DVSS.n6210 DVSS.n6209 0.4505
R28036 DVSS.n6130 DVSS.n6129 0.4505
R28037 DVSS.n6215 DVSS.n6214 0.4505
R28038 DVSS.n6216 DVSS.n6128 0.4505
R28039 DVSS.n6218 DVSS.n6217 0.4505
R28040 DVSS.n6126 DVSS.n6125 0.4505
R28041 DVSS.n6223 DVSS.n6222 0.4505
R28042 DVSS.n6224 DVSS.n6124 0.4505
R28043 DVSS.n6226 DVSS.n6225 0.4505
R28044 DVSS.n6122 DVSS.n6121 0.4505
R28045 DVSS.n6231 DVSS.n6230 0.4505
R28046 DVSS.n6232 DVSS.n6120 0.4505
R28047 DVSS.n6234 DVSS.n6233 0.4505
R28048 DVSS.n6118 DVSS.n6117 0.4505
R28049 DVSS.n6239 DVSS.n6238 0.4505
R28050 DVSS.n6240 DVSS.n6116 0.4505
R28051 DVSS.n6242 DVSS.n6241 0.4505
R28052 DVSS.n6114 DVSS.n6113 0.4505
R28053 DVSS.n6247 DVSS.n6246 0.4505
R28054 DVSS.n6248 DVSS.n6112 0.4505
R28055 DVSS.n6250 DVSS.n6249 0.4505
R28056 DVSS.n6110 DVSS.n6109 0.4505
R28057 DVSS.n6255 DVSS.n6254 0.4505
R28058 DVSS.n6256 DVSS.n6108 0.4505
R28059 DVSS.n6258 DVSS.n6257 0.4505
R28060 DVSS.n6106 DVSS.n6105 0.4505
R28061 DVSS.n6263 DVSS.n6262 0.4505
R28062 DVSS.n6264 DVSS.n6104 0.4505
R28063 DVSS.n6266 DVSS.n6265 0.4505
R28064 DVSS.n6102 DVSS.n6101 0.4505
R28065 DVSS.n6271 DVSS.n6270 0.4505
R28066 DVSS.n6272 DVSS.n6100 0.4505
R28067 DVSS.n6274 DVSS.n6273 0.4505
R28068 DVSS.n6098 DVSS.n6097 0.4505
R28069 DVSS.n6279 DVSS.n6278 0.4505
R28070 DVSS.n6280 DVSS.n6096 0.4505
R28071 DVSS.n6282 DVSS.n6281 0.4505
R28072 DVSS.n6094 DVSS.n6093 0.4505
R28073 DVSS.n6287 DVSS.n6286 0.4505
R28074 DVSS.n6288 DVSS.n6092 0.4505
R28075 DVSS.n6290 DVSS.n6289 0.4505
R28076 DVSS.n6090 DVSS.n6089 0.4505
R28077 DVSS.n6295 DVSS.n6294 0.4505
R28078 DVSS.n6296 DVSS.n6088 0.4505
R28079 DVSS.n6298 DVSS.n6297 0.4505
R28080 DVSS.n6086 DVSS.n6085 0.4505
R28081 DVSS.n6303 DVSS.n6302 0.4505
R28082 DVSS.n6304 DVSS.n6084 0.4505
R28083 DVSS.n6306 DVSS.n6305 0.4505
R28084 DVSS.n6082 DVSS.n6081 0.4505
R28085 DVSS.n6311 DVSS.n6310 0.4505
R28086 DVSS.n6312 DVSS.n6080 0.4505
R28087 DVSS.n6314 DVSS.n6313 0.4505
R28088 DVSS.n6078 DVSS.n6077 0.4505
R28089 DVSS.n6319 DVSS.n6318 0.4505
R28090 DVSS.n6320 DVSS.n6076 0.4505
R28091 DVSS.n6322 DVSS.n6321 0.4505
R28092 DVSS.n6074 DVSS.n6073 0.4505
R28093 DVSS.n6327 DVSS.n6326 0.4505
R28094 DVSS.n6328 DVSS.n6072 0.4505
R28095 DVSS.n6330 DVSS.n6329 0.4505
R28096 DVSS.n6070 DVSS.n6069 0.4505
R28097 DVSS.n6335 DVSS.n6334 0.4505
R28098 DVSS.n6336 DVSS.n6067 0.4505
R28099 DVSS.n6338 DVSS.n6337 0.4505
R28100 DVSS.n6068 DVSS.n6036 0.4505
R28101 DVSS.n6047 DVSS.n6046 0.4505
R28102 DVSS.n6044 DVSS.n6043 0.4505
R28103 DVSS.n6052 DVSS.n6051 0.4505
R28104 DVSS.n6053 DVSS.n6042 0.4505
R28105 DVSS.n6055 DVSS.n6054 0.4505
R28106 DVSS.n6040 DVSS.n6039 0.4505
R28107 DVSS.n6060 DVSS.n6059 0.4505
R28108 DVSS.n6061 DVSS.n6038 0.4505
R28109 DVSS.n6063 DVSS.n6062 0.4505
R28110 DVSS.n6035 DVSS.n6034 0.4505
R28111 DVSS.n6343 DVSS.n6342 0.4505
R28112 DVSS.n6434 DVSS.n6433 0.4505
R28113 DVSS.n6440 DVSS.n6439 0.4505
R28114 DVSS.n6441 DVSS.n6432 0.4505
R28115 DVSS.n6443 DVSS.n6442 0.4505
R28116 DVSS.n6447 DVSS.n6446 0.4505
R28117 DVSS.n6448 DVSS.n6431 0.4505
R28118 DVSS.n6450 DVSS.n6449 0.4505
R28119 DVSS.n6429 DVSS.n6428 0.4505
R28120 DVSS.n6455 DVSS.n6454 0.4505
R28121 DVSS.n6456 DVSS.n6427 0.4505
R28122 DVSS.n6458 DVSS.n6457 0.4505
R28123 DVSS.n6425 DVSS.n6424 0.4505
R28124 DVSS.n6463 DVSS.n6462 0.4505
R28125 DVSS.n6464 DVSS.n6423 0.4505
R28126 DVSS.n6466 DVSS.n6465 0.4505
R28127 DVSS.n6421 DVSS.n6420 0.4505
R28128 DVSS.n6471 DVSS.n6470 0.4505
R28129 DVSS.n6472 DVSS.n6419 0.4505
R28130 DVSS.n6474 DVSS.n6473 0.4505
R28131 DVSS.n6417 DVSS.n6416 0.4505
R28132 DVSS.n6479 DVSS.n6478 0.4505
R28133 DVSS.n6480 DVSS.n6415 0.4505
R28134 DVSS.n6482 DVSS.n6481 0.4505
R28135 DVSS.n6413 DVSS.n6412 0.4505
R28136 DVSS.n6487 DVSS.n6486 0.4505
R28137 DVSS.n6488 DVSS.n6411 0.4505
R28138 DVSS.n6490 DVSS.n6489 0.4505
R28139 DVSS.n6409 DVSS.n6408 0.4505
R28140 DVSS.n6495 DVSS.n6494 0.4505
R28141 DVSS.n6496 DVSS.n6407 0.4505
R28142 DVSS.n6498 DVSS.n6497 0.4505
R28143 DVSS.n6405 DVSS.n6404 0.4505
R28144 DVSS.n6503 DVSS.n6502 0.4505
R28145 DVSS.n6504 DVSS.n6403 0.4505
R28146 DVSS.n6506 DVSS.n6505 0.4505
R28147 DVSS.n6401 DVSS.n6400 0.4505
R28148 DVSS.n6511 DVSS.n6510 0.4505
R28149 DVSS.n6512 DVSS.n6399 0.4505
R28150 DVSS.n6514 DVSS.n6513 0.4505
R28151 DVSS.n6397 DVSS.n6396 0.4505
R28152 DVSS.n6519 DVSS.n6518 0.4505
R28153 DVSS.n6520 DVSS.n6395 0.4505
R28154 DVSS.n6522 DVSS.n6521 0.4505
R28155 DVSS.n6393 DVSS.n6392 0.4505
R28156 DVSS.n6527 DVSS.n6526 0.4505
R28157 DVSS.n6528 DVSS.n6391 0.4505
R28158 DVSS.n6530 DVSS.n6529 0.4505
R28159 DVSS.n6389 DVSS.n6388 0.4505
R28160 DVSS.n6535 DVSS.n6534 0.4505
R28161 DVSS.n6536 DVSS.n6387 0.4505
R28162 DVSS.n6538 DVSS.n6537 0.4505
R28163 DVSS.n6385 DVSS.n6384 0.4505
R28164 DVSS.n6543 DVSS.n6542 0.4505
R28165 DVSS.n6544 DVSS.n6383 0.4505
R28166 DVSS.n6546 DVSS.n6545 0.4505
R28167 DVSS.n6381 DVSS.n6380 0.4505
R28168 DVSS.n6551 DVSS.n6550 0.4505
R28169 DVSS.n6552 DVSS.n6379 0.4505
R28170 DVSS.n6554 DVSS.n6553 0.4505
R28171 DVSS.n6377 DVSS.n6376 0.4505
R28172 DVSS.n6559 DVSS.n6558 0.4505
R28173 DVSS.n6560 DVSS.n6375 0.4505
R28174 DVSS.n6562 DVSS.n6561 0.4505
R28175 DVSS.n6373 DVSS.n6372 0.4505
R28176 DVSS.n6567 DVSS.n6566 0.4505
R28177 DVSS.n6568 DVSS.n6371 0.4505
R28178 DVSS.n6570 DVSS.n6569 0.4505
R28179 DVSS.n6369 DVSS.n6368 0.4505
R28180 DVSS.n6575 DVSS.n6574 0.4505
R28181 DVSS.n6576 DVSS.n6367 0.4505
R28182 DVSS.n6578 DVSS.n6577 0.4505
R28183 DVSS.n6365 DVSS.n6364 0.4505
R28184 DVSS.n6583 DVSS.n6582 0.4505
R28185 DVSS.n6584 DVSS.n6363 0.4505
R28186 DVSS.n6586 DVSS.n6585 0.4505
R28187 DVSS.n6361 DVSS.n6360 0.4505
R28188 DVSS.n6591 DVSS.n6590 0.4505
R28189 DVSS.n6592 DVSS.n6359 0.4505
R28190 DVSS.n6594 DVSS.n6593 0.4505
R28191 DVSS.n6357 DVSS.n6356 0.4505
R28192 DVSS.n6599 DVSS.n6598 0.4505
R28193 DVSS.n6600 DVSS.n6355 0.4505
R28194 DVSS.n6602 DVSS.n6601 0.4505
R28195 DVSS.n6353 DVSS.n6352 0.4505
R28196 DVSS.n6607 DVSS.n6606 0.4505
R28197 DVSS.n6608 DVSS.n6351 0.4505
R28198 DVSS.n6610 DVSS.n6609 0.4505
R28199 DVSS.n6349 DVSS.n6348 0.4505
R28200 DVSS.n6615 DVSS.n6614 0.4505
R28201 DVSS.n6616 DVSS.n6031 0.4505
R28202 DVSS.n6618 DVSS.n6617 0.4505
R28203 DVSS.n6640 DVSS.n6639 0.4505
R28204 DVSS.n6638 DVSS.n6019 0.4505
R28205 DVSS.n6023 DVSS.n6020 0.4505
R28206 DVSS.n6634 DVSS.n6633 0.4505
R28207 DVSS.n6632 DVSS.n6022 0.4505
R28208 DVSS.n6631 DVSS.n6630 0.4505
R28209 DVSS.n6025 DVSS.n6024 0.4505
R28210 DVSS.n6626 DVSS.n6625 0.4505
R28211 DVSS.n6624 DVSS.n6027 0.4505
R28212 DVSS.n6623 DVSS.n6622 0.4505
R28213 DVSS.n6032 DVSS.n6029 0.4505
R28214 DVSS.n8250 DVSS.n8249 0.444037
R28215 DVSS.n8274 DVSS.n8273 0.444037
R28216 DVSS.n8291 DVSS.n8290 0.444037
R28217 DVSS.n8281 DVSS.n1446 0.444037
R28218 DVSS.n8237 DVSS.n8231 0.444037
R28219 DVSS.n8308 DVSS.n8307 0.444037
R28220 DVSS.n1379 DVSS.n1324 0.444037
R28221 DVSS.n8476 DVSS.n8475 0.444037
R28222 DVSS.n1281 DVSS.n1280 0.444037
R28223 DVSS.n1268 DVSS.n1265 0.444037
R28224 DVSS.n8376 DVSS.n8372 0.444037
R28225 DVSS.n8355 DVSS.n8354 0.444037
R28226 DVSS.n8449 DVSS.n8448 0.440926
R28227 DVSS.n8482 DVSS.n8480 0.440926
R28228 DVSS.n1286 DVSS.n1285 0.440926
R28229 DVSS.n1261 DVSS.n1260 0.440926
R28230 DVSS.n8370 DVSS.n1158 0.440926
R28231 DVSS.n8494 DVSS.n1104 0.440926
R28232 DVSS.n8502 DVSS.n8501 0.433833
R28233 DVSS.n8501 DVSS.n8500 0.433833
R28234 DVSS.n1291 DVSS.n1146 0.433833
R28235 DVSS.n8462 DVSS.n1146 0.433833
R28236 DVSS.n1293 DVSS.n1150 0.433833
R28237 DVSS.n8462 DVSS.n1150 0.433833
R28238 DVSS.n8484 DVSS.n1092 0.433833
R28239 DVSS.n8500 DVSS.n1092 0.433833
R28240 DVSS.n8463 DVSS.n1149 0.433833
R28241 DVSS.n8463 DVSS.n8462 0.433833
R28242 DVSS.n8499 DVSS.n8498 0.433833
R28243 DVSS.n8500 DVSS.n8499 0.433833
R28244 DVSS.n1096 DVSS.n1090 0.433833
R28245 DVSS.n8500 DVSS.n1090 0.433833
R28246 DVSS.n8461 DVSS.n8460 0.433833
R28247 DVSS.n8462 DVSS.n8461 0.433833
R28248 DVSS.n6345 DVSS.n6033 0.412804
R28249 DVSS.n6345 DVSS.n6344 0.412569
R28250 DVSS.n6346 DVSS.n6028 0.412128
R28251 DVSS.n6347 DVSS.n6346 0.411993
R28252 DVSS.n7098 DVSS.n7097 0.400007
R28253 DVSS.n7110 DVSS.n7109 0.400007
R28254 DVSS DVSS.t11 0.391676
R28255 DVSS DVSS.t5 0.391676
R28256 DVSS DVSS.t0 0.391676
R28257 DVSS DVSS.t27 0.391676
R28258 DVSS DVSS.t7 0.391676
R28259 DVSS DVSS.t33 0.391676
R28260 DVSS DVSS.t31 0.391676
R28261 DVSS DVSS.t24 0.391676
R28262 DVSS DVSS.t22 0.391676
R28263 DVSS DVSS.t36 0.391676
R28264 DVSS DVSS.t29 0.391676
R28265 DVSS DVSS.t8 0.391676
R28266 DVSS DVSS.t2 0.391676
R28267 DVSS DVSS.t26 0.391676
R28268 DVSS DVSS.t19 0.391676
R28269 DVSS DVSS.t20 0.391676
R28270 DVSS DVSS.t18 0.391676
R28271 DVSS DVSS.t32 0.391676
R28272 DVSS.n8243 DVSS.n1479 0.384436
R28273 DVSS.n8271 DVSS.n8270 0.384436
R28274 DVSS.n8294 DVSS.n8293 0.384436
R28275 DVSS.n8327 DVSS.n8321 0.384436
R28276 DVSS.n7145 DVSS.n1513 0.384436
R28277 DVSS.n8315 DVSS.n8314 0.384436
R28278 DVSS.n7134 DVSS 0.37265
R28279 DVSS.n8207 DVSS 0.37265
R28280 DVSS.n9023 DVSS.n9016 0.369923
R28281 DVSS.n9381 DVSS.n9378 0.369923
R28282 DVSS.n8870 DVSS.n8869 0.369923
R28283 DVSS.n9397 DVSS.n9395 0.369923
R28284 DVSS.n9012 DVSS.n9010 0.365885
R28285 DVSS.n9376 DVSS.n325 0.365885
R28286 DVSS.n8875 DVSS.n8874 0.365885
R28287 DVSS.n9406 DVSS.n9404 0.365885
R28288 DVSS.n1295 DVSS.n1293 0.356041
R28289 DVSS.n8503 DVSS.n8502 0.356041
R28290 DVSS.n8498 DVSS.n1095 0.356041
R28291 DVSS.n8460 DVSS.n1151 0.356041
R28292 DVSS.n3620 DVSS.n2818 0.347921
R28293 DVSS.n4849 DVSS.n2786 0.347921
R28294 DVSS.n4787 DVSS.n4785 0.347921
R28295 DVSS.n4420 DVSS.n3805 0.347921
R28296 DVSS.n4217 DVSS.n3817 0.347921
R28297 DVSS.n4963 DVSS.n2849 0.347921
R28298 DVSS.n4913 DVSS.n2878 0.347921
R28299 DVSS.n4453 DVSS.n4452 0.347921
R28300 DVSS.n5306 DVSS.n3423 0.347744
R28301 DVSS.n5271 DVSS.n3333 0.347744
R28302 DVSS.n4138 DVSS.n3149 0.347744
R28303 DVSS.n4185 DVSS.n3106 0.347744
R28304 DVSS.n5355 DVSS.n5354 0.347744
R28305 DVSS.n5914 DVSS.n5913 0.347744
R28306 DVSS.n5863 DVSS.n3005 0.347744
R28307 DVSS.n7061 DVSS.n7060 0.346681
R28308 DVSS.n1599 DVSS.n155 0.346681
R28309 DVSS.n1747 DVSS.n112 0.346681
R28310 DVSS.n6860 DVSS.n6859 0.346681
R28311 DVSS.n8336 DVSS.n8333 0.33552
R28312 DVSS.n7119 DVSS.n7118 0.33552
R28313 DVSS.n8083 DVSS 0.332375
R28314 DVSS.n8112 DVSS 0.332375
R28315 DVSS.n2687 DVSS 0.332375
R28316 DVSS.n2744 DVSS 0.332375
R28317 DVSS.n5684 DVSS 0.332375
R28318 DVSS.n5501 DVSS 0.332375
R28319 DVSS.n3883 DVSS 0.332375
R28320 DVSS.n4995 DVSS 0.332375
R28321 DVSS.n4434 DVSS 0.332375
R28322 DVSS.n4840 DVSS 0.332375
R28323 DVSS.n3548 DVSS 0.332375
R28324 DVSS.n5386 DVSS 0.332375
R28325 DVSS.n5655 DVSS 0.332375
R28326 DVSS.n5538 DVSS 0.332375
R28327 DVSS.n7343 DVSS 0.332375
R28328 DVSS.n7726 DVSS 0.332375
R28329 DVSS.n7250 DVSS 0.330584
R28330 DVSS.n7242 DVSS 0.330584
R28331 DVSS.n1890 DVSS.t4 0.312926
R28332 DVSS.n1890 DVSS.t11 0.312926
R28333 DVSS.n1854 DVSS.t5 0.312926
R28334 DVSS.n1854 DVSS.t16 0.312926
R28335 DVSS.n2660 DVSS.t30 0.312926
R28336 DVSS.n2660 DVSS.t0 0.312926
R28337 DVSS.n2717 DVSS.t27 0.312926
R28338 DVSS.n2717 DVSS.t12 0.312926
R28339 DVSS.n3246 DVSS.t35 0.312926
R28340 DVSS.n3246 DVSS.t7 0.312926
R28341 DVSS.n3322 DVSS.t33 0.312926
R28342 DVSS.n3322 DVSS.t14 0.312926
R28343 DVSS.n3882 DVSS.t23 0.312926
R28344 DVSS.n3882 DVSS.t31 0.312926
R28345 DVSS.n3578 DVSS.t24 0.312926
R28346 DVSS.n3578 DVSS.t10 0.312926
R28347 DVSS.n7169 DVSS.t9 0.312926
R28348 DVSS.n7169 DVSS.t25 0.312926
R28349 DVSS.n6653 DVSS.t25 0.312926
R28350 DVSS.n6653 DVSS.t32 0.312926
R28351 DVSS.n4643 DVSS.t13 0.312926
R28352 DVSS.n4643 DVSS.t28 0.312926
R28353 DVSS.n4023 DVSS.t10 0.312926
R28354 DVSS.n4023 DVSS.t23 0.312926
R28355 DVSS.n3500 DVSS.t15 0.312926
R28356 DVSS.n3500 DVSS.t1 0.312926
R28357 DVSS.n5718 DVSS.t14 0.312926
R28358 DVSS.n5718 DVSS.t35 0.312926
R28359 DVSS.n5426 DVSS.t6 0.312926
R28360 DVSS.n5426 DVSS.t21 0.312926
R28361 DVSS.n5602 DVSS.t12 0.312926
R28362 DVSS.n5602 DVSS.t30 0.312926
R28363 DVSS.n2639 DVSS.t34 0.312926
R28364 DVSS.n2639 DVSS.t17 0.312926
R28365 DVSS.n7896 DVSS.t16 0.312926
R28366 DVSS.n7896 DVSS.t4 0.312926
R28367 DVSS.n1539 DVSS.t22 0.312926
R28368 DVSS.n1539 DVSS.t9 0.312926
R28369 DVSS.n4433 DVSS.t28 0.312926
R28370 DVSS.n4433 DVSS.t36 0.312926
R28371 DVSS.n4829 DVSS.t29 0.312926
R28372 DVSS.n4829 DVSS.t13 0.312926
R28373 DVSS.n3528 DVSS.t1 0.312926
R28374 DVSS.n3528 DVSS.t8 0.312926
R28375 DVSS.n3350 DVSS.t2 0.312926
R28376 DVSS.n3350 DVSS.t15 0.312926
R28377 DVSS.n3266 DVSS.t21 0.312926
R28378 DVSS.n3266 DVSS.t26 0.312926
R28379 DVSS.n3297 DVSS.t19 0.312926
R28380 DVSS.n3297 DVSS.t6 0.312926
R28381 DVSS.n2605 DVSS.t17 0.312926
R28382 DVSS.n2605 DVSS.t20 0.312926
R28383 DVSS.n2090 DVSS.t18 0.312926
R28384 DVSS.n2090 DVSS.t34 0.312926
R28385 DVSS.n8180 DVSS.n8179 0.288039
R28386 DVSS.n8062 DVSS.n8061 0.288039
R28387 DVSS.n8120 DVSS.n8119 0.28237
R28388 DVSS.n7845 DVSS.n1856 0.28237
R28389 DVSS.n7974 DVSS.n1882 0.28237
R28390 DVSS.n8013 DVSS.n1892 0.28237
R28391 DVSS.n8036 DVSS.n1901 0.28237
R28392 DVSS.n1849 DVSS.n1794 0.28237
R28393 DVSS.n6645 DVSS.n1528 0.27557
R28394 DVSS.n7252 DVSS.n1523 0.27557
R28395 DVSS.n4479 DVSS.n3832 0.256847
R28396 DVSS.n5936 DVSS.n5935 0.256847
R28397 DVSS.n4234 DVSS.n3839 0.231338
R28398 DVSS.n4939 DVSS.n4938 0.231338
R28399 DVSS.n6769 DVSS.n6738 0.231338
R28400 DVSS.n1743 DVSS.n1742 0.231338
R28401 DVSS.n1941 DVSS.n1919 0.231338
R28402 DVSS.n8170 DVSS.n8169 0.231338
R28403 DVSS.n3076 DVSS.n2997 0.231338
R28404 DVSS.n5099 DVSS.n5094 0.231338
R28405 DVSS.n5850 DVSS.n3030 0.231338
R28406 DVSS.n5335 DVSS.n5330 0.231338
R28407 DVSS.n6637 DVSS.n6018 0.231338
R28408 DVSS.n6438 DVSS.n6437 0.231338
R28409 DVSS.n6049 DVSS.n6048 0.231338
R28410 DVSS.n6163 DVSS.n6155 0.231338
R28411 DVSS.n8212 DVSS.n8211 0.231169
R28412 DVSS.n7151 DVSS.n7150 0.231169
R28413 DVSS.n8207 DVSS.n8206 0.225249
R28414 DVSS.n7134 DVSS.n7133 0.225249
R28415 DVSS.n8470 DVSS.n567 0.224444
R28416 DVSS.n1382 DVSS.n595 0.224444
R28417 DVSS.n8638 DVSS.n979 0.221476
R28418 DVSS.n8680 DVSS.n8642 0.221476
R28419 DVSS.n7378 DVSS.n2528 0.220739
R28420 DVSS.n6910 DVSS.n6874 0.220739
R28421 DVSS.n7674 DVSS.n2119 0.220619
R28422 DVSS.n9935 DVSS.n9934 0.220619
R28423 DVSS.n9846 DVSS.n84 0.220619
R28424 DVSS.n9785 DVSS.n98 0.220619
R28425 DVSS.n7677 DVSS.n7673 0.214786
R28426 DVSS.n7383 DVSS.n7382 0.214786
R28427 DVSS.n7384 DVSS.n2527 0.214786
R28428 DVSS.n7386 DVSS.n7385 0.214786
R28429 DVSS.n2525 DVSS.n2524 0.214786
R28430 DVSS.n7391 DVSS.n7390 0.214786
R28431 DVSS.n7392 DVSS.n2523 0.214786
R28432 DVSS.n7394 DVSS.n7393 0.214786
R28433 DVSS.n2472 DVSS.n2471 0.214786
R28434 DVSS.n7402 DVSS.n7401 0.214786
R28435 DVSS.n7403 DVSS.n2470 0.214786
R28436 DVSS.n7405 DVSS.n7404 0.214786
R28437 DVSS.n2468 DVSS.n2467 0.214786
R28438 DVSS.n7410 DVSS.n7409 0.214786
R28439 DVSS.n7411 DVSS.n2466 0.214786
R28440 DVSS.n7413 DVSS.n7412 0.214786
R28441 DVSS.n2416 DVSS.n2415 0.214786
R28442 DVSS.n7422 DVSS.n7421 0.214786
R28443 DVSS.n7423 DVSS.n2414 0.214786
R28444 DVSS.n7425 DVSS.n7424 0.214786
R28445 DVSS.n2412 DVSS.n2411 0.214786
R28446 DVSS.n7430 DVSS.n7429 0.214786
R28447 DVSS.n7431 DVSS.n2410 0.214786
R28448 DVSS.n7433 DVSS.n7432 0.214786
R28449 DVSS.n2408 DVSS.n2407 0.214786
R28450 DVSS.n7438 DVSS.n7437 0.214786
R28451 DVSS.n7439 DVSS.n2406 0.214786
R28452 DVSS.n7441 DVSS.n7440 0.214786
R28453 DVSS.n2404 DVSS.n2403 0.214786
R28454 DVSS.n7446 DVSS.n7445 0.214786
R28455 DVSS.n7447 DVSS.n2402 0.214786
R28456 DVSS.n7449 DVSS.n7448 0.214786
R28457 DVSS.n2351 DVSS.n2350 0.214786
R28458 DVSS.n7457 DVSS.n7456 0.214786
R28459 DVSS.n7458 DVSS.n2349 0.214786
R28460 DVSS.n7460 DVSS.n7459 0.214786
R28461 DVSS.n2347 DVSS.n2346 0.214786
R28462 DVSS.n7465 DVSS.n7464 0.214786
R28463 DVSS.n7466 DVSS.n2345 0.214786
R28464 DVSS.n7468 DVSS.n7467 0.214786
R28465 DVSS.n2343 DVSS.n2342 0.214786
R28466 DVSS.n7473 DVSS.n7472 0.214786
R28467 DVSS.n7474 DVSS.n2341 0.214786
R28468 DVSS.n7476 DVSS.n7475 0.214786
R28469 DVSS.n2339 DVSS.n2338 0.214786
R28470 DVSS.n7481 DVSS.n7480 0.214786
R28471 DVSS.n7482 DVSS.n2337 0.214786
R28472 DVSS.n7484 DVSS.n7483 0.214786
R28473 DVSS.n2309 DVSS.n2308 0.214786
R28474 DVSS.n7492 DVSS.n7491 0.214786
R28475 DVSS.n7493 DVSS.n2307 0.214786
R28476 DVSS.n7495 DVSS.n7494 0.214786
R28477 DVSS.n2279 DVSS.n2278 0.214786
R28478 DVSS.n7503 DVSS.n7502 0.214786
R28479 DVSS.n7504 DVSS.n2277 0.214786
R28480 DVSS.n7506 DVSS.n7505 0.214786
R28481 DVSS.n2275 DVSS.n2274 0.214786
R28482 DVSS.n7511 DVSS.n7510 0.214786
R28483 DVSS.n7512 DVSS.n2273 0.214786
R28484 DVSS.n7514 DVSS.n7513 0.214786
R28485 DVSS.n2271 DVSS.n2270 0.214786
R28486 DVSS.n7519 DVSS.n7518 0.214786
R28487 DVSS.n7520 DVSS.n2269 0.214786
R28488 DVSS.n7522 DVSS.n7521 0.214786
R28489 DVSS.n2267 DVSS.n2266 0.214786
R28490 DVSS.n7527 DVSS.n7526 0.214786
R28491 DVSS.n7528 DVSS.n2265 0.214786
R28492 DVSS.n7530 DVSS.n7529 0.214786
R28493 DVSS.n2237 DVSS.n2236 0.214786
R28494 DVSS.n7561 DVSS.n7560 0.214786
R28495 DVSS.n7562 DVSS.n2235 0.214786
R28496 DVSS.n7564 DVSS.n7563 0.214786
R28497 DVSS.n2233 DVSS.n2232 0.214786
R28498 DVSS.n7569 DVSS.n7568 0.214786
R28499 DVSS.n7570 DVSS.n2231 0.214786
R28500 DVSS.n7572 DVSS.n7571 0.214786
R28501 DVSS.n2229 DVSS.n2228 0.214786
R28502 DVSS.n7577 DVSS.n7576 0.214786
R28503 DVSS.n7578 DVSS.n2227 0.214786
R28504 DVSS.n7580 DVSS.n7579 0.214786
R28505 DVSS.n2225 DVSS.n2224 0.214786
R28506 DVSS.n7585 DVSS.n7584 0.214786
R28507 DVSS.n7586 DVSS.n2223 0.214786
R28508 DVSS.n7588 DVSS.n7587 0.214786
R28509 DVSS.n2195 DVSS.n2194 0.214786
R28510 DVSS.n7619 DVSS.n7618 0.214786
R28511 DVSS.n7620 DVSS.n2193 0.214786
R28512 DVSS.n7622 DVSS.n7621 0.214786
R28513 DVSS.n2191 DVSS.n2190 0.214786
R28514 DVSS.n7627 DVSS.n7626 0.214786
R28515 DVSS.n7628 DVSS.n2189 0.214786
R28516 DVSS.n7630 DVSS.n7629 0.214786
R28517 DVSS.n2161 DVSS.n2160 0.214786
R28518 DVSS.n7661 DVSS.n7660 0.214786
R28519 DVSS.n7662 DVSS.n2159 0.214786
R28520 DVSS.n7665 DVSS.n7664 0.214786
R28521 DVSS.n7663 DVSS.n2156 0.214786
R28522 DVSS.n7669 DVSS.n2157 0.214786
R28523 DVSS.n7671 DVSS.n7670 0.214786
R28524 DVSS.n7672 DVSS.n2155 0.214786
R28525 DVSS.n7676 DVSS.n7675 0.214786
R28526 DVSS.n7678 DVSS.n7677 0.214786
R28527 DVSS.n7377 DVSS.n2529 0.214786
R28528 DVSS.n7382 DVSS.n7381 0.214786
R28529 DVSS.n2543 DVSS.n2527 0.214786
R28530 DVSS.n7387 DVSS.n7386 0.214786
R28531 DVSS.n7388 DVSS.n2525 0.214786
R28532 DVSS.n7390 DVSS.n7389 0.214786
R28533 DVSS.n2523 DVSS.n2522 0.214786
R28534 DVSS.n7395 DVSS.n7394 0.214786
R28535 DVSS.n7396 DVSS.n2472 0.214786
R28536 DVSS.n7401 DVSS.n7400 0.214786
R28537 DVSS.n2486 DVSS.n2470 0.214786
R28538 DVSS.n7406 DVSS.n7405 0.214786
R28539 DVSS.n7407 DVSS.n2468 0.214786
R28540 DVSS.n7409 DVSS.n7408 0.214786
R28541 DVSS.n2466 DVSS.n2465 0.214786
R28542 DVSS.n7414 DVSS.n7413 0.214786
R28543 DVSS.n7415 DVSS.n2416 0.214786
R28544 DVSS.n7421 DVSS.n7420 0.214786
R28545 DVSS.n2430 DVSS.n2414 0.214786
R28546 DVSS.n7426 DVSS.n7425 0.214786
R28547 DVSS.n7427 DVSS.n2412 0.214786
R28548 DVSS.n7429 DVSS.n7428 0.214786
R28549 DVSS.n2410 DVSS.n2409 0.214786
R28550 DVSS.n7434 DVSS.n7433 0.214786
R28551 DVSS.n7435 DVSS.n2408 0.214786
R28552 DVSS.n7437 DVSS.n7436 0.214786
R28553 DVSS.n2406 DVSS.n2405 0.214786
R28554 DVSS.n7442 DVSS.n7441 0.214786
R28555 DVSS.n7443 DVSS.n2404 0.214786
R28556 DVSS.n7445 DVSS.n7444 0.214786
R28557 DVSS.n2402 DVSS.n2401 0.214786
R28558 DVSS.n7450 DVSS.n7449 0.214786
R28559 DVSS.n7451 DVSS.n2351 0.214786
R28560 DVSS.n7456 DVSS.n7455 0.214786
R28561 DVSS.n2365 DVSS.n2349 0.214786
R28562 DVSS.n7461 DVSS.n7460 0.214786
R28563 DVSS.n7462 DVSS.n2347 0.214786
R28564 DVSS.n7464 DVSS.n7463 0.214786
R28565 DVSS.n2345 DVSS.n2344 0.214786
R28566 DVSS.n7469 DVSS.n7468 0.214786
R28567 DVSS.n7470 DVSS.n2343 0.214786
R28568 DVSS.n7472 DVSS.n7471 0.214786
R28569 DVSS.n2341 DVSS.n2340 0.214786
R28570 DVSS.n7477 DVSS.n7476 0.214786
R28571 DVSS.n7478 DVSS.n2339 0.214786
R28572 DVSS.n7480 DVSS.n7479 0.214786
R28573 DVSS.n2337 DVSS.n2336 0.214786
R28574 DVSS.n7485 DVSS.n7484 0.214786
R28575 DVSS.n7486 DVSS.n2309 0.214786
R28576 DVSS.n7491 DVSS.n7490 0.214786
R28577 DVSS.n2307 DVSS.n2306 0.214786
R28578 DVSS.n7496 DVSS.n7495 0.214786
R28579 DVSS.n7497 DVSS.n2279 0.214786
R28580 DVSS.n7502 DVSS.n7501 0.214786
R28581 DVSS.n2277 DVSS.n2276 0.214786
R28582 DVSS.n7507 DVSS.n7506 0.214786
R28583 DVSS.n7508 DVSS.n2275 0.214786
R28584 DVSS.n7510 DVSS.n7509 0.214786
R28585 DVSS.n2273 DVSS.n2272 0.214786
R28586 DVSS.n7515 DVSS.n7514 0.214786
R28587 DVSS.n7516 DVSS.n2271 0.214786
R28588 DVSS.n7518 DVSS.n7517 0.214786
R28589 DVSS.n2269 DVSS.n2268 0.214786
R28590 DVSS.n7523 DVSS.n7522 0.214786
R28591 DVSS.n7524 DVSS.n2267 0.214786
R28592 DVSS.n7526 DVSS.n7525 0.214786
R28593 DVSS.n2265 DVSS.n2253 0.214786
R28594 DVSS.n7531 DVSS.n7530 0.214786
R28595 DVSS.n7542 DVSS.n2237 0.214786
R28596 DVSS.n7560 DVSS.n7559 0.214786
R28597 DVSS.n2235 DVSS.n2234 0.214786
R28598 DVSS.n7565 DVSS.n7564 0.214786
R28599 DVSS.n7566 DVSS.n2233 0.214786
R28600 DVSS.n7568 DVSS.n7567 0.214786
R28601 DVSS.n2231 DVSS.n2230 0.214786
R28602 DVSS.n7573 DVSS.n7572 0.214786
R28603 DVSS.n7574 DVSS.n2229 0.214786
R28604 DVSS.n7576 DVSS.n7575 0.214786
R28605 DVSS.n2227 DVSS.n2226 0.214786
R28606 DVSS.n7581 DVSS.n7580 0.214786
R28607 DVSS.n7582 DVSS.n2225 0.214786
R28608 DVSS.n7584 DVSS.n7583 0.214786
R28609 DVSS.n2223 DVSS.n2211 0.214786
R28610 DVSS.n7589 DVSS.n7588 0.214786
R28611 DVSS.n7600 DVSS.n2195 0.214786
R28612 DVSS.n7618 DVSS.n7617 0.214786
R28613 DVSS.n2193 DVSS.n2192 0.214786
R28614 DVSS.n7623 DVSS.n7622 0.214786
R28615 DVSS.n7624 DVSS.n2191 0.214786
R28616 DVSS.n7626 DVSS.n7625 0.214786
R28617 DVSS.n2189 DVSS.n2177 0.214786
R28618 DVSS.n7631 DVSS.n7630 0.214786
R28619 DVSS.n7642 DVSS.n2161 0.214786
R28620 DVSS.n7660 DVSS.n7659 0.214786
R28621 DVSS.n2159 DVSS.n2158 0.214786
R28622 DVSS.n7666 DVSS.n7665 0.214786
R28623 DVSS.n7667 DVSS.n2156 0.214786
R28624 DVSS.n7669 DVSS.n7668 0.214786
R28625 DVSS.n7670 DVSS.n2121 0.214786
R28626 DVSS.n2155 DVSS.n2134 0.214786
R28627 DVSS.n9936 DVSS.n5 0.214786
R28628 DVSS.n9937 DVSS.n4 0.214786
R28629 DVSS.n8655 DVSS.n8654 0.214786
R28630 DVSS.n8666 DVSS.n963 0.214786
R28631 DVSS.n8684 DVSS.n8683 0.214786
R28632 DVSS.n961 DVSS.n960 0.214786
R28633 DVSS.n8689 DVSS.n8688 0.214786
R28634 DVSS.n8690 DVSS.n959 0.214786
R28635 DVSS.n8693 DVSS.n8692 0.214786
R28636 DVSS.n8691 DVSS.n956 0.214786
R28637 DVSS.n8697 DVSS.n957 0.214786
R28638 DVSS.n8699 DVSS.n8698 0.214786
R28639 DVSS.n8700 DVSS.n726 0.214786
R28640 DVSS.n954 DVSS.n738 0.214786
R28641 DVSS.n8705 DVSS.n8704 0.214786
R28642 DVSS.n8706 DVSS.n953 0.214786
R28643 DVSS.n8708 DVSS.n8707 0.214786
R28644 DVSS.n8713 DVSS.n8712 0.214786
R28645 DVSS.n8714 DVSS.n901 0.214786
R28646 DVSS.n8719 DVSS.n8718 0.214786
R28647 DVSS.n916 DVSS.n899 0.214786
R28648 DVSS.n8724 DVSS.n8723 0.214786
R28649 DVSS.n8725 DVSS.n897 0.214786
R28650 DVSS.n8727 DVSS.n8726 0.214786
R28651 DVSS.n895 DVSS.n894 0.214786
R28652 DVSS.n8732 DVSS.n8731 0.214786
R28653 DVSS.n8733 DVSS.n893 0.214786
R28654 DVSS.n8735 DVSS.n8734 0.214786
R28655 DVSS.n891 DVSS.n890 0.214786
R28656 DVSS.n8740 DVSS.n8739 0.214786
R28657 DVSS.n8741 DVSS.n889 0.214786
R28658 DVSS.n8743 DVSS.n8742 0.214786
R28659 DVSS.n887 DVSS.n886 0.214786
R28660 DVSS.n8748 DVSS.n8747 0.214786
R28661 DVSS.n8749 DVSS.n838 0.214786
R28662 DVSS.n8754 DVSS.n8753 0.214786
R28663 DVSS.n853 DVSS.n836 0.214786
R28664 DVSS.n8760 DVSS.n8759 0.214786
R28665 DVSS.n8761 DVSS.n834 0.214786
R28666 DVSS.n8763 DVSS.n8762 0.214786
R28667 DVSS.n8764 DVSS.n830 0.214786
R28668 DVSS.n8810 DVSS.n8809 0.214786
R28669 DVSS.n832 DVSS.n831 0.214786
R28670 DVSS.n8805 DVSS.n8768 0.214786
R28671 DVSS.n8804 DVSS.n8769 0.214786
R28672 DVSS.n8803 DVSS.n8770 0.214786
R28673 DVSS.n8773 DVSS.n8771 0.214786
R28674 DVSS.n8799 DVSS.n8774 0.214786
R28675 DVSS.n8798 DVSS.n8775 0.214786
R28676 DVSS.n8797 DVSS.n663 0.214786
R28677 DVSS.n8776 DVSS.n675 0.214786
R28678 DVSS.n8793 DVSS.n8789 0.214786
R28679 DVSS.n8792 DVSS.n8791 0.214786
R28680 DVSS.n8790 DVSS.n498 0.214786
R28681 DVSS.n9262 DVSS.n9261 0.214786
R28682 DVSS.n500 DVSS.n496 0.214786
R28683 DVSS.n9267 DVSS.n9266 0.214786
R28684 DVSS.n9268 DVSS.n494 0.214786
R28685 DVSS.n9270 DVSS.n9269 0.214786
R28686 DVSS.n492 DVSS.n491 0.214786
R28687 DVSS.n9275 DVSS.n9274 0.214786
R28688 DVSS.n9276 DVSS.n490 0.214786
R28689 DVSS.n9279 DVSS.n9278 0.214786
R28690 DVSS.n9277 DVSS.n487 0.214786
R28691 DVSS.n9283 DVSS.n488 0.214786
R28692 DVSS.n9288 DVSS.n9287 0.214786
R28693 DVSS.n9289 DVSS.n485 0.214786
R28694 DVSS.n9291 DVSS.n9290 0.214786
R28695 DVSS.n9292 DVSS.n394 0.214786
R28696 DVSS.n481 DVSS.n460 0.214786
R28697 DVSS.n9352 DVSS.n9351 0.214786
R28698 DVSS.n483 DVSS.n482 0.214786
R28699 DVSS.n9347 DVSS.n9296 0.214786
R28700 DVSS.n9346 DVSS.n9297 0.214786
R28701 DVSS.n9345 DVSS.n9298 0.214786
R28702 DVSS.n9301 DVSS.n9299 0.214786
R28703 DVSS.n9341 DVSS.n9302 0.214786
R28704 DVSS.n9340 DVSS.n9303 0.214786
R28705 DVSS.n9339 DVSS.n9304 0.214786
R28706 DVSS.n9307 DVSS.n9305 0.214786
R28707 DVSS.n9335 DVSS.n9308 0.214786
R28708 DVSS.n9334 DVSS.n9309 0.214786
R28709 DVSS.n9333 DVSS.n9310 0.214786
R28710 DVSS.n9312 DVSS.n9311 0.214786
R28711 DVSS.n9329 DVSS.n288 0.214786
R28712 DVSS.n9328 DVSS.n300 0.214786
R28713 DVSS.n9327 DVSS.n9325 0.214786
R28714 DVSS.n286 DVSS.n61 0.214786
R28715 DVSS.n9870 DVSS.n62 0.214786
R28716 DVSS.n58 DVSS.n57 0.214786
R28717 DVSS.n9876 DVSS.n9875 0.214786
R28718 DVSS.n9877 DVSS.n56 0.214786
R28719 DVSS.n9879 DVSS.n9878 0.214786
R28720 DVSS.n53 DVSS.n52 0.214786
R28721 DVSS.n9885 DVSS.n9884 0.214786
R28722 DVSS.n54 DVSS.n24 0.214786
R28723 DVSS.n9889 DVSS.n23 0.214786
R28724 DVSS.n9891 DVSS.n9890 0.214786
R28725 DVSS.n21 DVSS.n20 0.214786
R28726 DVSS.n9896 DVSS.n9895 0.214786
R28727 DVSS.n9897 DVSS.n2 0.214786
R28728 DVSS.n9938 DVSS.n3 0.214786
R28729 DVSS.n9845 DVSS.n9844 0.214786
R28730 DVSS.n85 DVSS.n83 0.214786
R28731 DVSS.n9849 DVSS.n82 0.214786
R28732 DVSS.n9850 DVSS.n81 0.214786
R28733 DVSS.n9851 DVSS.n80 0.214786
R28734 DVSS.n79 DVSS.n77 0.214786
R28735 DVSS.n9855 DVSS.n76 0.214786
R28736 DVSS.n9856 DVSS.n75 0.214786
R28737 DVSS.n9857 DVSS.n74 0.214786
R28738 DVSS.n342 DVSS.n72 0.214786
R28739 DVSS.n9861 DVSS.n71 0.214786
R28740 DVSS.n9862 DVSS.n70 0.214786
R28741 DVSS.n9863 DVSS.n69 0.214786
R28742 DVSS.n68 DVSS.n66 0.214786
R28743 DVSS.n9867 DVSS.n65 0.214786
R28744 DVSS.n271 DVSS.n64 0.214786
R28745 DVSS.n9587 DVSS.n9584 0.214786
R28746 DVSS.n9588 DVSS.n266 0.214786
R28747 DVSS.n9589 DVSS.n265 0.214786
R28748 DVSS.n9548 DVSS.n263 0.214786
R28749 DVSS.n9593 DVSS.n262 0.214786
R28750 DVSS.n9594 DVSS.n261 0.214786
R28751 DVSS.n9595 DVSS.n260 0.214786
R28752 DVSS.n259 DVSS.n257 0.214786
R28753 DVSS.n9599 DVSS.n256 0.214786
R28754 DVSS.n9600 DVSS.n255 0.214786
R28755 DVSS.n9601 DVSS.n254 0.214786
R28756 DVSS.n253 DVSS.n251 0.214786
R28757 DVSS.n9605 DVSS.n250 0.214786
R28758 DVSS.n9606 DVSS.n249 0.214786
R28759 DVSS.n9607 DVSS.n248 0.214786
R28760 DVSS.n443 DVSS.n246 0.214786
R28761 DVSS.n9611 DVSS.n245 0.214786
R28762 DVSS.n9612 DVSS.n244 0.214786
R28763 DVSS.n9613 DVSS.n243 0.214786
R28764 DVSS.n409 DVSS.n241 0.214786
R28765 DVSS.n9617 DVSS.n240 0.214786
R28766 DVSS.n9618 DVSS.n239 0.214786
R28767 DVSS.n9619 DVSS.n238 0.214786
R28768 DVSS.n9182 DVSS.n9181 0.214786
R28769 DVSS.n9184 DVSS.n550 0.214786
R28770 DVSS.n9185 DVSS.n549 0.214786
R28771 DVSS.n9186 DVSS.n548 0.214786
R28772 DVSS.n547 DVSS.n545 0.214786
R28773 DVSS.n9190 DVSS.n544 0.214786
R28774 DVSS.n9191 DVSS.n543 0.214786
R28775 DVSS.n9192 DVSS.n542 0.214786
R28776 DVSS.n541 DVSS.n538 0.214786
R28777 DVSS.n9197 DVSS.n9196 0.214786
R28778 DVSS.n537 DVSS.n516 0.214786
R28779 DVSS.n9068 DVSS.n503 0.214786
R28780 DVSS.n9069 DVSS.n9066 0.214786
R28781 DVSS.n9070 DVSS.n647 0.214786
R28782 DVSS.n9039 DVSS.n645 0.214786
R28783 DVSS.n9074 DVSS.n644 0.214786
R28784 DVSS.n9075 DVSS.n643 0.214786
R28785 DVSS.n9076 DVSS.n642 0.214786
R28786 DVSS.n641 DVSS.n639 0.214786
R28787 DVSS.n9080 DVSS.n638 0.214786
R28788 DVSS.n9081 DVSS.n637 0.214786
R28789 DVSS.n9082 DVSS.n636 0.214786
R28790 DVSS.n635 DVSS.n633 0.214786
R28791 DVSS.n9086 DVSS.n632 0.214786
R28792 DVSS.n8814 DVSS.n631 0.214786
R28793 DVSS.n8818 DVSS.n8815 0.214786
R28794 DVSS.n8819 DVSS.n829 0.214786
R28795 DVSS.n8820 DVSS.n810 0.214786
R28796 DVSS.n826 DVSS.n809 0.214786
R28797 DVSS.n8825 DVSS.n8824 0.214786
R28798 DVSS.n825 DVSS.n824 0.214786
R28799 DVSS.n7004 DVSS.n7003 0.214786
R28800 DVSS.n7007 DVSS.n7002 0.214786
R28801 DVSS.n7008 DVSS.n7001 0.214786
R28802 DVSS.n7009 DVSS.n7000 0.214786
R28803 DVSS.n6999 DVSS.n6997 0.214786
R28804 DVSS.n7013 DVSS.n6996 0.214786
R28805 DVSS.n7014 DVSS.n6995 0.214786
R28806 DVSS.n7015 DVSS.n6994 0.214786
R28807 DVSS.n6993 DVSS.n6991 0.214786
R28808 DVSS.n7019 DVSS.n6990 0.214786
R28809 DVSS.n7020 DVSS.n6989 0.214786
R28810 DVSS.n7021 DVSS.n6988 0.214786
R28811 DVSS.n6987 DVSS.n6981 0.214786
R28812 DVSS.n7026 DVSS.n7025 0.214786
R28813 DVSS.n6980 DVSS.n6968 0.214786
R28814 DVSS.n6983 DVSS.n6943 0.214786
R28815 DVSS.n7031 DVSS.n1031 0.214786
R28816 DVSS.n8601 DVSS.n1030 0.214786
R28817 DVSS.n8604 DVSS.n1029 0.214786
R28818 DVSS.n8605 DVSS.n1028 0.214786
R28819 DVSS.n8606 DVSS.n1027 0.214786
R28820 DVSS.n1025 DVSS.n1024 0.214786
R28821 DVSS.n8610 DVSS.n1023 0.214786
R28822 DVSS.n8611 DVSS.n770 0.214786
R28823 DVSS.n8612 DVSS.n758 0.214786
R28824 DVSS.n1021 DVSS.n1020 0.214786
R28825 DVSS.n8616 DVSS.n1019 0.214786
R28826 DVSS.n8617 DVSS.n1018 0.214786
R28827 DVSS.n8618 DVSS.n1017 0.214786
R28828 DVSS.n1015 DVSS.n1014 0.214786
R28829 DVSS.n8623 DVSS.n8622 0.214786
R28830 DVSS.n1013 DVSS.n992 0.214786
R28831 DVSS.n136 DVSS.n135 0.214786
R28832 DVSS.n9788 DVSS.n9787 0.214786
R28833 DVSS.n134 DVSS.n113 0.214786
R28834 DVSS.n9782 DVSS.n100 0.214786
R28835 DVSS.n9781 DVSS.n9780 0.214786
R28836 DVSS.n9779 DVSS.n138 0.214786
R28837 DVSS.n9778 DVSS.n9777 0.214786
R28838 DVSS.n140 DVSS.n139 0.214786
R28839 DVSS.n9772 DVSS.n9771 0.214786
R28840 DVSS.n9735 DVSS.n142 0.214786
R28841 DVSS.n9733 DVSS.n9732 0.214786
R28842 DVSS.n9726 DVSS.n159 0.214786
R28843 DVSS.n9728 DVSS.n9727 0.214786
R28844 DVSS.n9725 DVSS.n161 0.214786
R28845 DVSS.n9724 DVSS.n9723 0.214786
R28846 DVSS.n9719 DVSS.n9718 0.214786
R28847 DVSS.n165 DVSS.n164 0.214786
R28848 DVSS.n9691 DVSS.n9690 0.214786
R28849 DVSS.n189 DVSS.n186 0.214786
R28850 DVSS.n9686 DVSS.n9685 0.214786
R28851 DVSS.n9684 DVSS.n191 0.214786
R28852 DVSS.n9683 DVSS.n9682 0.214786
R28853 DVSS.n193 DVSS.n192 0.214786
R28854 DVSS.n9678 DVSS.n9677 0.214786
R28855 DVSS.n9676 DVSS.n195 0.214786
R28856 DVSS.n9675 DVSS.n9674 0.214786
R28857 DVSS.n197 DVSS.n196 0.214786
R28858 DVSS.n9670 DVSS.n9669 0.214786
R28859 DVSS.n9668 DVSS.n199 0.214786
R28860 DVSS.n9667 DVSS.n9666 0.214786
R28861 DVSS.n201 DVSS.n200 0.214786
R28862 DVSS.n9662 DVSS.n9661 0.214786
R28863 DVSS.n204 DVSS.n203 0.214786
R28864 DVSS.n9634 DVSS.n9633 0.214786
R28865 DVSS.n228 DVSS.n225 0.214786
R28866 DVSS.n9629 DVSS.n9628 0.214786
R28867 DVSS.n9627 DVSS.n230 0.214786
R28868 DVSS.n9626 DVSS.n9625 0.214786
R28869 DVSS.n232 DVSS.n231 0.214786
R28870 DVSS.n9178 DVSS.n9177 0.214786
R28871 DVSS.n9175 DVSS.n551 0.214786
R28872 DVSS.n9169 DVSS.n552 0.214786
R28873 DVSS.n9171 DVSS.n9170 0.214786
R28874 DVSS.n9168 DVSS.n554 0.214786
R28875 DVSS.n9167 DVSS.n9166 0.214786
R28876 DVSS.n556 DVSS.n555 0.214786
R28877 DVSS.n9162 DVSS.n9161 0.214786
R28878 DVSS.n9160 DVSS.n558 0.214786
R28879 DVSS.n584 DVSS.n559 0.214786
R28880 DVSS.n9138 DVSS.n9137 0.214786
R28881 DVSS.n583 DVSS.n575 0.214786
R28882 DVSS.n9132 DVSS.n9131 0.214786
R28883 DVSS.n587 DVSS.n586 0.214786
R28884 DVSS.n9111 DVSS.n9110 0.214786
R28885 DVSS.n617 DVSS.n607 0.214786
R28886 DVSS.n9106 DVSS.n9105 0.214786
R28887 DVSS.n9104 DVSS.n619 0.214786
R28888 DVSS.n9103 DVSS.n9102 0.214786
R28889 DVSS.n621 DVSS.n620 0.214786
R28890 DVSS.n9098 DVSS.n9097 0.214786
R28891 DVSS.n9096 DVSS.n623 0.214786
R28892 DVSS.n9095 DVSS.n9094 0.214786
R28893 DVSS.n625 DVSS.n624 0.214786
R28894 DVSS.n9089 DVSS.n629 0.214786
R28895 DVSS.n8563 DVSS.n628 0.214786
R28896 DVSS.n8565 DVSS.n8564 0.214786
R28897 DVSS.n8568 DVSS.n8562 0.214786
R28898 DVSS.n8569 DVSS.n1061 0.214786
R28899 DVSS.n8570 DVSS.n1060 0.214786
R28900 DVSS.n8542 DVSS.n1058 0.214786
R28901 DVSS.n8574 DVSS.n1057 0.214786
R28902 DVSS.n8575 DVSS.n1056 0.214786
R28903 DVSS.n8576 DVSS.n1055 0.214786
R28904 DVSS.n1054 DVSS.n1052 0.214786
R28905 DVSS.n8580 DVSS.n1051 0.214786
R28906 DVSS.n8581 DVSS.n1050 0.214786
R28907 DVSS.n8582 DVSS.n1049 0.214786
R28908 DVSS.n1048 DVSS.n1046 0.214786
R28909 DVSS.n8586 DVSS.n1045 0.214786
R28910 DVSS.n8587 DVSS.n1044 0.214786
R28911 DVSS.n8588 DVSS.n1043 0.214786
R28912 DVSS.n1042 DVSS.n1040 0.214786
R28913 DVSS.n8592 DVSS.n1039 0.214786
R28914 DVSS.n8593 DVSS.n1038 0.214786
R28915 DVSS.n8594 DVSS.n1037 0.214786
R28916 DVSS.n1202 DVSS.n1034 0.214786
R28917 DVSS.n8598 DVSS.n1033 0.214786
R28918 DVSS.n7034 DVSS.n1032 0.214786
R28919 DVSS.n7038 DVSS.n7035 0.214786
R28920 DVSS.n7039 DVSS.n6930 0.214786
R28921 DVSS.n7040 DVSS.n6929 0.214786
R28922 DVSS.n6727 DVSS.n6726 0.214786
R28923 DVSS.n7045 DVSS.n7044 0.214786
R28924 DVSS.n6725 DVSS.n6704 0.214786
R28925 DVSS.n6925 DVSS.n6693 0.214786
R28926 DVSS.n6924 DVSS.n6923 0.214786
R28927 DVSS.n6922 DVSS.n6729 0.214786
R28928 DVSS.n6921 DVSS.n6920 0.214786
R28929 DVSS.n6731 DVSS.n6730 0.214786
R28930 DVSS.n6915 DVSS.n6914 0.214786
R28931 DVSS.n6905 DVSS.n6733 0.214786
R28932 DVSS.n6886 DVSS.n6885 0.214786
R28933 DVSS.n6733 DVSS.n6732 0.214786
R28934 DVSS.n6916 DVSS.n6915 0.214786
R28935 DVSS.n6917 DVSS.n6731 0.214786
R28936 DVSS.n6920 DVSS.n6919 0.214786
R28937 DVSS.n6918 DVSS.n6729 0.214786
R28938 DVSS.n6924 DVSS.n6728 0.214786
R28939 DVSS.n6926 DVSS.n6925 0.214786
R28940 DVSS.n6927 DVSS.n6725 0.214786
R28941 DVSS.n7044 DVSS.n7043 0.214786
R28942 DVSS.n7042 DVSS.n6727 0.214786
R28943 DVSS.n7041 DVSS.n7040 0.214786
R28944 DVSS.n7039 DVSS.n6928 0.214786
R28945 DVSS.n7038 DVSS.n7037 0.214786
R28946 DVSS.n7036 DVSS.n1032 0.214786
R28947 DVSS.n8598 DVSS.n8597 0.214786
R28948 DVSS.n8596 DVSS.n1034 0.214786
R28949 DVSS.n8595 DVSS.n8594 0.214786
R28950 DVSS.n8593 DVSS.n1036 0.214786
R28951 DVSS.n8592 DVSS.n8591 0.214786
R28952 DVSS.n8590 DVSS.n1040 0.214786
R28953 DVSS.n8589 DVSS.n8588 0.214786
R28954 DVSS.n8587 DVSS.n1041 0.214786
R28955 DVSS.n8586 DVSS.n8585 0.214786
R28956 DVSS.n8584 DVSS.n1046 0.214786
R28957 DVSS.n8583 DVSS.n8582 0.214786
R28958 DVSS.n8581 DVSS.n1047 0.214786
R28959 DVSS.n8580 DVSS.n8579 0.214786
R28960 DVSS.n8578 DVSS.n1052 0.214786
R28961 DVSS.n8577 DVSS.n8576 0.214786
R28962 DVSS.n8575 DVSS.n1053 0.214786
R28963 DVSS.n8574 DVSS.n8573 0.214786
R28964 DVSS.n8572 DVSS.n1058 0.214786
R28965 DVSS.n8571 DVSS.n8570 0.214786
R28966 DVSS.n8569 DVSS.n1059 0.214786
R28967 DVSS.n8568 DVSS.n8567 0.214786
R28968 DVSS.n8566 DVSS.n8565 0.214786
R28969 DVSS.n628 DVSS.n627 0.214786
R28970 DVSS.n9090 DVSS.n9089 0.214786
R28971 DVSS.n9092 DVSS.n625 0.214786
R28972 DVSS.n9094 DVSS.n9093 0.214786
R28973 DVSS.n623 DVSS.n622 0.214786
R28974 DVSS.n9099 DVSS.n9098 0.214786
R28975 DVSS.n9100 DVSS.n621 0.214786
R28976 DVSS.n9102 DVSS.n9101 0.214786
R28977 DVSS.n619 DVSS.n618 0.214786
R28978 DVSS.n9107 DVSS.n9106 0.214786
R28979 DVSS.n9108 DVSS.n617 0.214786
R28980 DVSS.n9110 DVSS.n9109 0.214786
R28981 DVSS.n586 DVSS.n585 0.214786
R28982 DVSS.n9133 DVSS.n9132 0.214786
R28983 DVSS.n9134 DVSS.n583 0.214786
R28984 DVSS.n9137 DVSS.n9136 0.214786
R28985 DVSS.n9135 DVSS.n584 0.214786
R28986 DVSS.n558 DVSS.n557 0.214786
R28987 DVSS.n9163 DVSS.n9162 0.214786
R28988 DVSS.n9164 DVSS.n556 0.214786
R28989 DVSS.n9166 DVSS.n9165 0.214786
R28990 DVSS.n554 DVSS.n553 0.214786
R28991 DVSS.n9172 DVSS.n9171 0.214786
R28992 DVSS.n9173 DVSS.n552 0.214786
R28993 DVSS.n9175 DVSS.n9174 0.214786
R28994 DVSS.n9177 DVSS.n233 0.214786
R28995 DVSS.n9623 DVSS.n232 0.214786
R28996 DVSS.n9625 DVSS.n9624 0.214786
R28997 DVSS.n230 DVSS.n229 0.214786
R28998 DVSS.n9630 DVSS.n9629 0.214786
R28999 DVSS.n9631 DVSS.n228 0.214786
R29000 DVSS.n9633 DVSS.n9632 0.214786
R29001 DVSS.n203 DVSS.n202 0.214786
R29002 DVSS.n9663 DVSS.n9662 0.214786
R29003 DVSS.n9664 DVSS.n201 0.214786
R29004 DVSS.n9666 DVSS.n9665 0.214786
R29005 DVSS.n199 DVSS.n198 0.214786
R29006 DVSS.n9671 DVSS.n9670 0.214786
R29007 DVSS.n9672 DVSS.n197 0.214786
R29008 DVSS.n9674 DVSS.n9673 0.214786
R29009 DVSS.n195 DVSS.n194 0.214786
R29010 DVSS.n9679 DVSS.n9678 0.214786
R29011 DVSS.n9680 DVSS.n193 0.214786
R29012 DVSS.n9682 DVSS.n9681 0.214786
R29013 DVSS.n191 DVSS.n190 0.214786
R29014 DVSS.n9687 DVSS.n9686 0.214786
R29015 DVSS.n9688 DVSS.n189 0.214786
R29016 DVSS.n9690 DVSS.n9689 0.214786
R29017 DVSS.n164 DVSS.n163 0.214786
R29018 DVSS.n9720 DVSS.n9719 0.214786
R29019 DVSS.n9723 DVSS.n9722 0.214786
R29020 DVSS.n161 DVSS.n160 0.214786
R29021 DVSS.n9729 DVSS.n9728 0.214786
R29022 DVSS.n9730 DVSS.n159 0.214786
R29023 DVSS.n9732 DVSS.n9731 0.214786
R29024 DVSS.n142 DVSS.n141 0.214786
R29025 DVSS.n9773 DVSS.n9772 0.214786
R29026 DVSS.n9774 DVSS.n140 0.214786
R29027 DVSS.n9777 DVSS.n9776 0.214786
R29028 DVSS.n9775 DVSS.n138 0.214786
R29029 DVSS.n9781 DVSS.n137 0.214786
R29030 DVSS.n9783 DVSS.n9782 0.214786
R29031 DVSS.n9784 DVSS.n134 0.214786
R29032 DVSS.n9787 DVSS.n9786 0.214786
R29033 DVSS.n8622 DVSS.n8621 0.214786
R29034 DVSS.n8620 DVSS.n1015 0.214786
R29035 DVSS.n8619 DVSS.n8618 0.214786
R29036 DVSS.n8617 DVSS.n1016 0.214786
R29037 DVSS.n8616 DVSS.n8615 0.214786
R29038 DVSS.n8614 DVSS.n1021 0.214786
R29039 DVSS.n8613 DVSS.n8612 0.214786
R29040 DVSS.n8611 DVSS.n1022 0.214786
R29041 DVSS.n8610 DVSS.n8609 0.214786
R29042 DVSS.n8608 DVSS.n1025 0.214786
R29043 DVSS.n8607 DVSS.n8606 0.214786
R29044 DVSS.n8605 DVSS.n1026 0.214786
R29045 DVSS.n8604 DVSS.n8603 0.214786
R29046 DVSS.n8602 DVSS.n8601 0.214786
R29047 DVSS.n6982 DVSS.n1031 0.214786
R29048 DVSS.n6984 DVSS.n6983 0.214786
R29049 DVSS.n6985 DVSS.n6980 0.214786
R29050 DVSS.n7025 DVSS.n7024 0.214786
R29051 DVSS.n7023 DVSS.n6981 0.214786
R29052 DVSS.n7022 DVSS.n7021 0.214786
R29053 DVSS.n7020 DVSS.n6986 0.214786
R29054 DVSS.n7019 DVSS.n7018 0.214786
R29055 DVSS.n7017 DVSS.n6991 0.214786
R29056 DVSS.n7016 DVSS.n7015 0.214786
R29057 DVSS.n7014 DVSS.n6992 0.214786
R29058 DVSS.n7013 DVSS.n7012 0.214786
R29059 DVSS.n7011 DVSS.n6997 0.214786
R29060 DVSS.n7010 DVSS.n7009 0.214786
R29061 DVSS.n7008 DVSS.n6998 0.214786
R29062 DVSS.n7007 DVSS.n7006 0.214786
R29063 DVSS.n7005 DVSS.n7004 0.214786
R29064 DVSS.n827 DVSS.n825 0.214786
R29065 DVSS.n8824 DVSS.n8823 0.214786
R29066 DVSS.n8822 DVSS.n826 0.214786
R29067 DVSS.n8821 DVSS.n8820 0.214786
R29068 DVSS.n8819 DVSS.n828 0.214786
R29069 DVSS.n8818 DVSS.n8817 0.214786
R29070 DVSS.n8816 DVSS.n631 0.214786
R29071 DVSS.n9086 DVSS.n9085 0.214786
R29072 DVSS.n9084 DVSS.n633 0.214786
R29073 DVSS.n9083 DVSS.n9082 0.214786
R29074 DVSS.n9081 DVSS.n634 0.214786
R29075 DVSS.n9080 DVSS.n9079 0.214786
R29076 DVSS.n9078 DVSS.n639 0.214786
R29077 DVSS.n9077 DVSS.n9076 0.214786
R29078 DVSS.n9075 DVSS.n640 0.214786
R29079 DVSS.n9074 DVSS.n9073 0.214786
R29080 DVSS.n9072 DVSS.n645 0.214786
R29081 DVSS.n9071 DVSS.n9070 0.214786
R29082 DVSS.n9069 DVSS.n646 0.214786
R29083 DVSS.n9068 DVSS.n9067 0.214786
R29084 DVSS.n539 DVSS.n537 0.214786
R29085 DVSS.n9196 DVSS.n9195 0.214786
R29086 DVSS.n9194 DVSS.n538 0.214786
R29087 DVSS.n9193 DVSS.n9192 0.214786
R29088 DVSS.n9191 DVSS.n540 0.214786
R29089 DVSS.n9190 DVSS.n9189 0.214786
R29090 DVSS.n9188 DVSS.n545 0.214786
R29091 DVSS.n9187 DVSS.n9186 0.214786
R29092 DVSS.n9185 DVSS.n546 0.214786
R29093 DVSS.n9184 DVSS.n9183 0.214786
R29094 DVSS.n9182 DVSS.n235 0.214786
R29095 DVSS.n9620 DVSS.n9619 0.214786
R29096 DVSS.n9618 DVSS.n236 0.214786
R29097 DVSS.n9617 DVSS.n9616 0.214786
R29098 DVSS.n9615 DVSS.n241 0.214786
R29099 DVSS.n9614 DVSS.n9613 0.214786
R29100 DVSS.n9612 DVSS.n242 0.214786
R29101 DVSS.n9611 DVSS.n9610 0.214786
R29102 DVSS.n9609 DVSS.n246 0.214786
R29103 DVSS.n9608 DVSS.n9607 0.214786
R29104 DVSS.n9606 DVSS.n247 0.214786
R29105 DVSS.n9605 DVSS.n9604 0.214786
R29106 DVSS.n9603 DVSS.n251 0.214786
R29107 DVSS.n9602 DVSS.n9601 0.214786
R29108 DVSS.n9600 DVSS.n252 0.214786
R29109 DVSS.n9599 DVSS.n9598 0.214786
R29110 DVSS.n9597 DVSS.n257 0.214786
R29111 DVSS.n9596 DVSS.n9595 0.214786
R29112 DVSS.n9594 DVSS.n258 0.214786
R29113 DVSS.n9593 DVSS.n9592 0.214786
R29114 DVSS.n9591 DVSS.n263 0.214786
R29115 DVSS.n9590 DVSS.n9589 0.214786
R29116 DVSS.n9588 DVSS.n264 0.214786
R29117 DVSS.n9587 DVSS.n9586 0.214786
R29118 DVSS.n9585 DVSS.n64 0.214786
R29119 DVSS.n9867 DVSS.n9866 0.214786
R29120 DVSS.n9865 DVSS.n66 0.214786
R29121 DVSS.n9864 DVSS.n9863 0.214786
R29122 DVSS.n9862 DVSS.n67 0.214786
R29123 DVSS.n9861 DVSS.n9860 0.214786
R29124 DVSS.n9859 DVSS.n72 0.214786
R29125 DVSS.n9858 DVSS.n9857 0.214786
R29126 DVSS.n9856 DVSS.n73 0.214786
R29127 DVSS.n9855 DVSS.n9854 0.214786
R29128 DVSS.n9853 DVSS.n77 0.214786
R29129 DVSS.n9852 DVSS.n9851 0.214786
R29130 DVSS.n9850 DVSS.n78 0.214786
R29131 DVSS.n9849 DVSS.n9848 0.214786
R29132 DVSS.n9847 DVSS.n83 0.214786
R29133 DVSS.n9937 DVSS.n1 0.214786
R29134 DVSS.n963 DVSS.n962 0.214786
R29135 DVSS.n8685 DVSS.n8684 0.214786
R29136 DVSS.n8686 DVSS.n961 0.214786
R29137 DVSS.n8688 DVSS.n8687 0.214786
R29138 DVSS.n959 DVSS.n958 0.214786
R29139 DVSS.n8694 DVSS.n8693 0.214786
R29140 DVSS.n8695 DVSS.n956 0.214786
R29141 DVSS.n8697 DVSS.n8696 0.214786
R29142 DVSS.n8699 DVSS.n955 0.214786
R29143 DVSS.n8701 DVSS.n8700 0.214786
R29144 DVSS.n8702 DVSS.n954 0.214786
R29145 DVSS.n8704 DVSS.n8703 0.214786
R29146 DVSS.n953 DVSS.n952 0.214786
R29147 DVSS.n8709 DVSS.n8708 0.214786
R29148 DVSS.n8712 DVSS.n8711 0.214786
R29149 DVSS.n901 DVSS.n900 0.214786
R29150 DVSS.n8720 DVSS.n8719 0.214786
R29151 DVSS.n8721 DVSS.n899 0.214786
R29152 DVSS.n8723 DVSS.n8722 0.214786
R29153 DVSS.n897 DVSS.n896 0.214786
R29154 DVSS.n8728 DVSS.n8727 0.214786
R29155 DVSS.n8729 DVSS.n895 0.214786
R29156 DVSS.n8731 DVSS.n8730 0.214786
R29157 DVSS.n893 DVSS.n892 0.214786
R29158 DVSS.n8736 DVSS.n8735 0.214786
R29159 DVSS.n8737 DVSS.n891 0.214786
R29160 DVSS.n8739 DVSS.n8738 0.214786
R29161 DVSS.n889 DVSS.n888 0.214786
R29162 DVSS.n8744 DVSS.n8743 0.214786
R29163 DVSS.n8745 DVSS.n887 0.214786
R29164 DVSS.n8747 DVSS.n8746 0.214786
R29165 DVSS.n838 DVSS.n837 0.214786
R29166 DVSS.n8755 DVSS.n8754 0.214786
R29167 DVSS.n8756 DVSS.n836 0.214786
R29168 DVSS.n8759 DVSS.n8758 0.214786
R29169 DVSS.n8757 DVSS.n834 0.214786
R29170 DVSS.n8763 DVSS.n833 0.214786
R29171 DVSS.n8765 DVSS.n8764 0.214786
R29172 DVSS.n8809 DVSS.n8808 0.214786
R29173 DVSS.n8807 DVSS.n832 0.214786
R29174 DVSS.n8806 DVSS.n8805 0.214786
R29175 DVSS.n8804 DVSS.n8767 0.214786
R29176 DVSS.n8803 DVSS.n8802 0.214786
R29177 DVSS.n8801 DVSS.n8771 0.214786
R29178 DVSS.n8800 DVSS.n8799 0.214786
R29179 DVSS.n8798 DVSS.n8772 0.214786
R29180 DVSS.n8797 DVSS.n8796 0.214786
R29181 DVSS.n8795 DVSS.n8776 0.214786
R29182 DVSS.n8794 DVSS.n8793 0.214786
R29183 DVSS.n8792 DVSS.n8777 0.214786
R29184 DVSS.n498 DVSS.n497 0.214786
R29185 DVSS.n9263 DVSS.n9262 0.214786
R29186 DVSS.n9264 DVSS.n496 0.214786
R29187 DVSS.n9266 DVSS.n9265 0.214786
R29188 DVSS.n494 DVSS.n493 0.214786
R29189 DVSS.n9271 DVSS.n9270 0.214786
R29190 DVSS.n9272 DVSS.n492 0.214786
R29191 DVSS.n9274 DVSS.n9273 0.214786
R29192 DVSS.n490 DVSS.n489 0.214786
R29193 DVSS.n9280 DVSS.n9279 0.214786
R29194 DVSS.n9281 DVSS.n487 0.214786
R29195 DVSS.n9283 DVSS.n9282 0.214786
R29196 DVSS.n9287 DVSS.n9286 0.214786
R29197 DVSS.n9285 DVSS.n485 0.214786
R29198 DVSS.n9291 DVSS.n484 0.214786
R29199 DVSS.n9293 DVSS.n9292 0.214786
R29200 DVSS.n9294 DVSS.n481 0.214786
R29201 DVSS.n9351 DVSS.n9350 0.214786
R29202 DVSS.n9349 DVSS.n483 0.214786
R29203 DVSS.n9348 DVSS.n9347 0.214786
R29204 DVSS.n9346 DVSS.n9295 0.214786
R29205 DVSS.n9345 DVSS.n9344 0.214786
R29206 DVSS.n9343 DVSS.n9299 0.214786
R29207 DVSS.n9342 DVSS.n9341 0.214786
R29208 DVSS.n9340 DVSS.n9300 0.214786
R29209 DVSS.n9339 DVSS.n9338 0.214786
R29210 DVSS.n9337 DVSS.n9305 0.214786
R29211 DVSS.n9336 DVSS.n9335 0.214786
R29212 DVSS.n9334 DVSS.n9306 0.214786
R29213 DVSS.n9333 DVSS.n9332 0.214786
R29214 DVSS.n9331 DVSS.n9312 0.214786
R29215 DVSS.n9330 DVSS.n9329 0.214786
R29216 DVSS.n9328 DVSS.n9313 0.214786
R29217 DVSS.n9327 DVSS.n9326 0.214786
R29218 DVSS.n61 DVSS.n60 0.214786
R29219 DVSS.n9871 DVSS.n9870 0.214786
R29220 DVSS.n9873 DVSS.n58 0.214786
R29221 DVSS.n9875 DVSS.n9874 0.214786
R29222 DVSS.n56 DVSS.n55 0.214786
R29223 DVSS.n9880 DVSS.n9879 0.214786
R29224 DVSS.n9881 DVSS.n53 0.214786
R29225 DVSS.n9884 DVSS.n9883 0.214786
R29226 DVSS.n9882 DVSS.n54 0.214786
R29227 DVSS.n23 DVSS.n22 0.214786
R29228 DVSS.n9892 DVSS.n9891 0.214786
R29229 DVSS.n9893 DVSS.n21 0.214786
R29230 DVSS.n9895 DVSS.n9894 0.214786
R29231 DVSS.n2 DVSS.n0 0.214786
R29232 DVSS.n9939 DVSS.n9938 0.214786
R29233 DVSS.n8459 DVSS.n1149 0.208878
R29234 DVSS.n1188 DVSS.n1149 0.208878
R29235 DVSS.n1293 DVSS.n1292 0.208878
R29236 DVSS.n8485 DVSS.n8484 0.208878
R29237 DVSS.n8484 DVSS.n1088 0.208878
R29238 DVSS.n8502 DVSS.n1088 0.208878
R29239 DVSS.n1291 DVSS.n1188 0.208878
R29240 DVSS.n1292 DVSS.n1291 0.208878
R29241 DVSS.n8498 DVSS.n8497 0.208878
R29242 DVSS.n8497 DVSS.n1096 0.208878
R29243 DVSS.n8485 DVSS.n1096 0.208878
R29244 DVSS.n8460 DVSS.n8459 0.208878
R29245 DVSS.n4474 DVSS.n4473 0.188545
R29246 DVSS.n5927 DVSS.n2910 0.188545
R29247 DVSS.n8481 DVSS.n177 0.188295
R29248 DVSS.n8477 DVSS.n216 0.188295
R29249 DVSS.n8447 DVSS.n1073 0.188295
R29250 DVSS.n1317 DVSS.n1316 0.188295
R29251 DVSS.n4804 DVSS 0.188139
R29252 DVSS DVSS.n4823 0.188139
R29253 DVSS.n4099 DVSS 0.188139
R29254 DVSS.n5001 DVSS 0.188139
R29255 DVSS.n3558 DVSS 0.188139
R29256 DVSS.n5029 DVSS 0.188139
R29257 DVSS.n5691 DVSS 0.188139
R29258 DVSS DVSS.n5494 0.188139
R29259 DVSS DVSS.n5645 0.188139
R29260 DVSS.n5636 DVSS 0.188139
R29261 DVSS.n2694 DVSS 0.188139
R29262 DVSS.n2751 DVSS 0.188139
R29263 DVSS DVSS.n7333 0.188139
R29264 DVSS.n7860 DVSS 0.188139
R29265 DVSS.n8090 DVSS 0.188139
R29266 DVSS DVSS.n8105 0.188139
R29267 DVSS.n4470 DVSS.n3798 0.177483
R29268 DVSS.n2907 DVSS.n2906 0.177483
R29269 DVSS.n8193 DVSS.n8192 0.169941
R29270 DVSS.n6749 DVSS.n6662 0.169941
R29271 DVSS.n1479 DVSS.n1476 0.167502
R29272 DVSS.n8270 DVSS.n1454 0.167502
R29273 DVSS.n4435 DVSS.n4434 0.156611
R29274 DVSS.n4840 DVSS.n4839 0.156611
R29275 DVSS.n4189 DVSS.n3883 0.156611
R29276 DVSS.n4995 DVSS.n4994 0.156611
R29277 DVSS.n3548 DVSS.n3547 0.156611
R29278 DVSS.n5386 DVSS.n5385 0.156611
R29279 DVSS.n5684 DVSS.n5683 0.156611
R29280 DVSS.n5503 DVSS.n5501 0.156611
R29281 DVSS.n5661 DVSS.n5655 0.156611
R29282 DVSS.n5538 DVSS.n5537 0.156611
R29283 DVSS.n2687 DVSS.n2686 0.156611
R29284 DVSS.n2744 DVSS.n2743 0.156611
R29285 DVSS.n7349 DVSS.n7343 0.156611
R29286 DVSS.n7726 DVSS.n7725 0.156611
R29287 DVSS.n8083 DVSS.n8082 0.156611
R29288 DVSS.n8114 DVSS.n8112 0.156611
R29289 DVSS.n9006 DVSS.n9004 0.148192
R29290 DVSS.n9541 DVSS.n9537 0.148192
R29291 DVSS.n8883 DVSS.n8879 0.148192
R29292 DVSS.n9415 DVSS.n9413 0.148192
R29293 DVSS.n8474 DVSS.n1143 0.143739
R29294 DVSS.n8402 DVSS.n1387 0.143739
R29295 DVSS.n8306 DVSS.n1471 0.139092
R29296 DVSS.n8280 DVSS.n8279 0.139092
R29297 DVSS.n1518 DVSS.n1507 0.139092
R29298 DVSS.n8254 DVSS.n1497 0.139092
R29299 DVSS.n7102 DVSS.n1415 0.138035
R29300 DVSS.n7107 DVSS.n1368 0.138035
R29301 DVSS.n7135 DVSS.n7134 0.137763
R29302 DVSS.n8208 DVSS.n8207 0.137763
R29303 DVSS DVSS.n7154 0.136254
R29304 DVSS.n8210 DVSS 0.136254
R29305 DVSS.n8219 DVSS.n1467 0.135923
R29306 DVSS.n7095 DVSS.n1499 0.135923
R29307 DVSS.n8224 DVSS.n8223 0.135923
R29308 DVSS.n7083 DVSS.n1492 0.135923
R29309 DVSS DVSS.n8199 0.129215
R29310 DVSS DVSS.n7067 0.129215
R29311 DVSS.n8488 DVSS.n8487 0.120618
R29312 DVSS.n8479 DVSS.n1135 0.120618
R29313 DVSS.n8442 DVSS.n8440 0.120618
R29314 DVSS.n8451 DVSS.n8450 0.120618
R29315 DVSS.n8313 DVSS.n1465 0.11672
R29316 DVSS.n8272 DVSS.n1449 0.11672
R29317 DVSS.n8239 DVSS.n8238 0.11672
R29318 DVSS.n8248 DVSS.n1490 0.11672
R29319 DVSS.n7704 DVSS.n1772 0.116189
R29320 DVSS.n7367 DVSS.n1927 0.116189
R29321 DVSS.n1546 DVSS.n1116 0.115835
R29322 DVSS.n8341 DVSS.n8339 0.115835
R29323 DVSS.n7123 DVSS.n1335 0.115835
R29324 DVSS.n7127 DVSS.n1173 0.115835
R29325 DVSS DVSS.n3877 0.114389
R29326 DVSS DVSS.n3540 0.114389
R29327 DVSS DVSS.n5677 0.114389
R29328 DVSS.n5668 DVSS 0.114389
R29329 DVSS.n8216 DVSS.n1461 0.114063
R29330 DVSS.n8331 DVSS.n8328 0.114063
R29331 DVSS.n7148 DVSS.n1516 0.114063
R29332 DVSS.n8292 DVSS.n1484 0.114063
R29333 DVSS.n8621 DVSS.n979 0.110647
R29334 DVSS.n8642 DVSS.n962 0.110647
R29335 DVSS.n7383 DVSS.n2528 0.110634
R29336 DVSS.n7674 DVSS.n7673 0.110634
R29337 DVSS.n6874 DVSS.n6732 0.110634
R29338 DVSS.n9786 DVSS.n9785 0.110634
R29339 DVSS.n9847 DVSS.n9846 0.110634
R29340 DVSS.n9935 DVSS.n1 0.110634
R29341 DVSS.n8122 DVSS.n1814 0.11052
R29342 DVSS.n7848 DVSS.n7847 0.11052
R29343 DVSS.n7335 DVSS.n2018 0.11052
R29344 DVSS.n7345 DVSS.n1984 0.11052
R29345 DVSS.n7354 DVSS.n1958 0.11052
R29346 DVSS.n7711 DVSS.n1789 0.11052
R29347 DVSS.n1188 DVSS.n1147 0.110159
R29348 DVSS.n8485 DVSS.n1091 0.110159
R29349 DVSS.n4434 DVSS.n3716 0.108278
R29350 DVSS.n4845 DVSS.n4840 0.108278
R29351 DVSS.n4004 DVSS.n3883 0.108278
R29352 DVSS.n4996 DVSS.n4995 0.108278
R29353 DVSS.n3549 DVSS.n3548 0.108278
R29354 DVSS.n5387 DVSS.n5386 0.108278
R29355 DVSS.n5686 DVSS.n5684 0.108278
R29356 DVSS.n5501 DVSS.n5500 0.108278
R29357 DVSS.n5655 DVSS.n5654 0.108278
R29358 DVSS.n5544 DVSS.n5538 0.108278
R29359 DVSS.n2689 DVSS.n2687 0.108278
R29360 DVSS.n2746 DVSS.n2744 0.108278
R29361 DVSS.n7343 DVSS.n7342 0.108278
R29362 DVSS.n7852 DVSS.n7726 0.108278
R29363 DVSS.n8085 DVSS.n8083 0.108278
R29364 DVSS.n8112 DVSS.n8111 0.108278
R29365 DVSS.n7145 DVSS.n1475 0.101041
R29366 DVSS.n1479 DVSS.n1475 0.101041
R29367 DVSS.n8294 DVSS.n1480 0.101041
R29368 DVSS.n8270 DVSS.n1450 0.101041
R29369 DVSS.n8321 DVSS.n1450 0.101041
R29370 DVSS.n8321 DVSS.n8320 0.101041
R29371 DVSS.n8295 DVSS.n1479 0.101041
R29372 DVSS.n8295 DVSS.n8294 0.101041
R29373 DVSS.n8316 DVSS.n8315 0.101041
R29374 DVSS.n8315 DVSS.n1459 0.101041
R29375 DVSS.n8270 DVSS.n1459 0.101041
R29376 DVSS.n7146 DVSS.n7145 0.101041
R29377 DVSS.n4441 DVSS.n4440 0.0982778
R29378 DVSS.n4978 DVSS.n3593 0.0982778
R29379 DVSS.n4989 DVSS.n2920 0.0982778
R29380 DVSS.n5380 DVSS.n5379 0.0982778
R29381 DVSS.n5515 DVSS.n2962 0.0982778
R29382 DVSS.n5525 DVSS.n2971 0.0982778
R29383 DVSS.n2676 DVSS.n2582 0.0982778
R29384 DVSS.n2735 DVSS.n2116 0.0982778
R29385 DVSS.n7362 DVSS.n7361 0.0982778
R29386 DVSS.n7715 DVSS.n7709 0.0982778
R29387 DVSS.n8072 DVSS.n8070 0.0982778
R29388 DVSS.n1848 DVSS.n1758 0.0982778
R29389 DVSS.n5901 DVSS.n2133 0.0967008
R29390 DVSS.n5894 DVSS.n2542 0.0967008
R29391 DVSS.n3875 DVSS.n3025 0.0941111
R29392 DVSS.n3538 DVSS.n3537 0.0941111
R29393 DVSS.n5674 DVSS.n5672 0.0941111
R29394 DVSS.n5665 DVSS.n2987 0.0941111
R29395 DVSS.n5530 DVSS.n2208 0.0910315
R29396 DVSS.n5540 DVSS.n2250 0.0910315
R29397 DVSS.n5647 DVSS.n2364 0.0910315
R29398 DVSS.n5657 DVSS.n2429 0.0910315
R29399 DVSS.n5521 DVSS.n2174 0.0910315
R29400 DVSS.n1318 DVSS.n1188 0.0873883
R29401 DVSS.n8486 DVSS.n8485 0.0873883
R29402 DVSS.n1292 DVSS.n1290 0.0873883
R29403 DVSS.n1256 DVSS.n1088 0.0873883
R29404 DVSS.n8459 DVSS.n8458 0.0873883
R29405 DVSS.n8497 DVSS.n8496 0.0873883
R29406 DVSS DVSS.n4803 0.0796667
R29407 DVSS.n4824 DVSS 0.0796667
R29408 DVSS DVSS.n4010 0.0796667
R29409 DVSS DVSS.n4998 0.0796667
R29410 DVSS DVSS.n3555 0.0796667
R29411 DVSS DVSS.n3346 0.0796667
R29412 DVSS DVSS.n5690 0.0796667
R29413 DVSS.n5496 DVSS 0.0796667
R29414 DVSS.n5651 DVSS 0.0796667
R29415 DVSS DVSS.n5547 0.0796667
R29416 DVSS DVSS.n2693 0.0796667
R29417 DVSS DVSS.n2749 0.0796667
R29418 DVSS.n7339 DVSS 0.0796667
R29419 DVSS DVSS.n7855 0.0796667
R29420 DVSS DVSS.n8089 0.0796667
R29421 DVSS.n8107 DVSS 0.0796667
R29422 DVSS.n7254 DVSS.n7253 0.0786237
R29423 DVSS.n4438 DVSS 0.0757778
R29424 DVSS DVSS.n3590 0.0757778
R29425 DVSS DVSS.n4991 0.0757778
R29426 DVSS DVSS.n5382 0.0757778
R29427 DVSS.n5509 DVSS 0.0757778
R29428 DVSS DVSS.n5528 0.0757778
R29429 DVSS DVSS.n2680 0.0757778
R29430 DVSS DVSS.n2738 0.0757778
R29431 DVSS.n7358 DVSS 0.0757778
R29432 DVSS DVSS.n7718 0.0757778
R29433 DVSS DVSS.n8076 0.0757778
R29434 DVSS DVSS.n1851 0.0757778
R29435 DVSS.n9214 DVSS.n9213 0.0740211
R29436 DVSS.n9064 DVSS.n9027 0.0740211
R29437 DVSS.n6013 DVSS.n6012 0.0702987
R29438 DVSS.n3675 DVSS.n2758 0.0702987
R29439 DVSS.n5005 DVSS.n5004 0.0702987
R29440 DVSS.n5007 DVSS.n5006 0.0702987
R29441 DVSS.n3234 DVSS.n2977 0.0702987
R29442 DVSS.n3284 DVSS.n2755 0.0702987
R29443 DVSS.n7265 DVSS.n7264 0.0702987
R29444 DVSS.n7263 DVSS.n2624 0.0702987
R29445 DVSS.n2757 DVSS.n1870 0.0702987
R29446 DVSS.n9546 DVSS.n9545 0.0621535
R29447 DVSS.n459 DVSS.n458 0.0621535
R29448 DVSS.n852 DVSS.n822 0.0621535
R29449 DVSS.n7029 DVSS.n915 0.0621535
R29450 DVSS.n9805 DVSS.n9804 0.0621535
R29451 DVSS.n9842 DVSS.n17 0.0621535
R29452 DVSS.n6872 DVSS.n991 0.0621535
R29453 DVSS.n8640 DVSS.n8639 0.0621535
R29454 DVSS.n7247 DVSS.n7156 0.059675
R29455 DVSS.n4036 DVSS.n3670 0.0571197
R29456 DVSS.n4089 DVSS.n3563 0.0571197
R29457 DVSS.n5488 DVSS.n5487 0.0571197
R29458 DVSS.n5485 DVSS.n5484 0.0571197
R29459 DVSS.n5639 DVSS.n5638 0.0571197
R29460 DVSS.n5631 DVSS.n5630 0.0571197
R29461 DVSS.n2704 DVSS.n2650 0.0571197
R29462 DVSS.n7327 DVSS.n7326 0.0571197
R29463 DVSS.n7862 DVSS.n7861 0.0571197
R29464 DVSS.n8099 DVSS.n8098 0.0571197
R29465 DVSS.n7184 DVSS.n1868 0.0571197
R29466 DVSS.n4807 DVSS.n3705 0.0571197
R29467 DVSS.n4094 DVSS.n4093 0.0571197
R29468 DVSS.n5697 DVSS.n5696 0.0571197
R29469 DVSS.n5482 DVSS.n3236 0.0571197
R29470 DVSS.n5642 DVSS.n5641 0.0571197
R29471 DVSS.n5628 DVSS.n3275 0.0571197
R29472 DVSS.n7272 DVSS.n7271 0.0571197
R29473 DVSS.n7330 DVSS.n7329 0.0571197
R29474 DVSS.n2615 DVSS.n2076 0.0571197
R29475 DVSS.n8096 DVSS.n8095 0.0571197
R29476 DVSS.n7182 DVSS.n1879 0.0571197
R29477 DVSS.n5835 DVSS.n3045 0.0569562
R29478 DVSS.n3053 DVSS.n3044 0.0569562
R29479 DVSS.n3052 DVSS.n3043 0.0569562
R29480 DVSS.n3061 DVSS.n3055 0.0569562
R29481 DVSS.n3068 DVSS.n3060 0.0569562
R29482 DVSS.n5675 DVSS.n3256 0.0569562
R29483 DVSS.n5673 DVSS.n3256 0.0569562
R29484 DVSS.n3259 DVSS.n3258 0.0569562
R29485 DVSS.n5666 DVSS.n3259 0.0569562
R29486 DVSS.n3053 DVSS.n3045 0.0569562
R29487 DVSS.n3052 DVSS.n3044 0.0569562
R29488 DVSS.n3068 DVSS.n3061 0.0569562
R29489 DVSS.n3067 DVSS.n3060 0.0569562
R29490 DVSS.n5676 DVSS.n3066 0.0563
R29491 DVSS.n5670 DVSS.n5669 0.0563
R29492 DVSS.n7246 DVSS.n7239 0.0560634
R29493 DVSS.n7248 DVSS.n7155 0.0560634
R29494 DVSS.n8200 DVSS 0.0487682
R29495 DVSS.n7068 DVSS 0.0487682
R29496 DVSS.n5195 DVSS.n3190 0.0459225
R29497 DVSS.n5740 DVSS.n5739 0.0459225
R29498 DVSS.n7116 DVSS.n7115 0.0450718
R29499 DVSS.n8330 DVSS.n1442 0.0450718
R29500 DVSS.n8329 DVSS.n1442 0.0450718
R29501 DVSS.n7144 DVSS.n7140 0.0450718
R29502 DVSS.n8215 DVSS.n1529 0.0450718
R29503 DVSS.n1294 DVSS.n1219 0.0450718
R29504 DVSS.n1219 DVSS.n1218 0.0450718
R29505 DVSS.n1218 DVSS.n1217 0.0450718
R29506 DVSS.n8530 DVSS.n8528 0.0450718
R29507 DVSS.n8524 DVSS.n1080 0.0450718
R29508 DVSS.n8524 DVSS.n8523 0.0450718
R29509 DVSS.n8518 DVSS.n8517 0.0450718
R29510 DVSS.n8517 DVSS.n8516 0.0450718
R29511 DVSS.n8512 DVSS.n1084 0.0450718
R29512 DVSS.n8512 DVSS.n8511 0.0450718
R29513 DVSS.n8511 DVSS.n1085 0.0450718
R29514 DVSS.n8506 DVSS.n1086 0.0450718
R29515 DVSS.n8506 DVSS.n8505 0.0450718
R29516 DVSS.n8505 DVSS.n1087 0.0450718
R29517 DVSS.n7125 DVSS.n7073 0.0450718
R29518 DVSS.n7122 DVSS.n7075 0.0450718
R29519 DVSS.n8337 DVSS.n1439 0.0450718
R29520 DVSS.n1547 DVSS.n1544 0.0450718
R29521 DVSS.n7114 DVSS.n7113 0.0442838
R29522 DVSS.n7113 DVSS.n7112 0.0442838
R29523 DVSS.n7082 DVSS.n7081 0.0442838
R29524 DVSS.n7084 DVSS.n7082 0.0442838
R29525 DVSS.n7094 DVSS.n7091 0.0442838
R29526 DVSS.n7096 DVSS.n7091 0.0442838
R29527 DVSS.n1444 DVSS.n1441 0.0442838
R29528 DVSS.n7142 DVSS.n7141 0.0442838
R29529 DVSS.n7149 DVSS.n7142 0.0442838
R29530 DVSS.n1522 DVSS.n1521 0.0442838
R29531 DVSS.n8222 DVSS.n1521 0.0442838
R29532 DVSS.n1527 DVSS.n1526 0.0442838
R29533 DVSS.n8218 DVSS.n1527 0.0442838
R29534 DVSS.n8214 DVSS.n8213 0.0442838
R29535 DVSS.n8213 DVSS.n1458 0.0442838
R29536 DVSS.n8531 DVSS.n8529 0.0442838
R29537 DVSS.n7126 DVSS.n7074 0.0442838
R29538 DVSS.n7128 DVSS.n7074 0.0442838
R29539 DVSS.n7121 DVSS.n7120 0.0442838
R29540 DVSS.n7120 DVSS.n7077 0.0442838
R29541 DVSS.n7105 DVSS.n7087 0.0442838
R29542 DVSS.n7108 DVSS.n7087 0.0442838
R29543 DVSS.n7101 DVSS.n7100 0.0442838
R29544 DVSS.n7100 DVSS.n1440 0.0442838
R29545 DVSS.n8335 DVSS.n8334 0.0442838
R29546 DVSS.n8334 DVSS.n1438 0.0442838
R29547 DVSS.n1549 DVSS.n1548 0.0442838
R29548 DVSS.n1548 DVSS.n1095 0.0442838
R29549 DVSS.n4812 DVSS.n3675 0.0437
R29550 DVSS.n5004 DVSS.n3561 0.0437
R29551 DVSS.n5199 DVSS.n5007 0.0437
R29552 DVSS.n3234 DVSS.n3229 0.0437
R29553 DVSS.n5640 DVSS.n3284 0.0437
R29554 DVSS.n7265 DVSS.n2701 0.0437
R29555 DVSS.n7328 DVSS.n2624 0.0437
R29556 DVSS.n8097 DVSS.n1870 0.0437
R29557 DVSS DVSS.n1890 0.039875
R29558 DVSS DVSS.n1854 0.039875
R29559 DVSS DVSS.n2660 0.039875
R29560 DVSS DVSS.n2717 0.039875
R29561 DVSS DVSS.n3246 0.039875
R29562 DVSS DVSS.n3322 0.039875
R29563 DVSS DVSS.n3882 0.039875
R29564 DVSS DVSS.n3578 0.039875
R29565 DVSS DVSS.n6653 0.039875
R29566 DVSS DVSS.n1539 0.039875
R29567 DVSS DVSS.n4433 0.039875
R29568 DVSS DVSS.n4829 0.039875
R29569 DVSS DVSS.n3528 0.039875
R29570 DVSS DVSS.n3350 0.039875
R29571 DVSS DVSS.n3266 0.039875
R29572 DVSS DVSS.n3297 0.039875
R29573 DVSS DVSS.n2605 0.039875
R29574 DVSS DVSS.n2090 0.039875
R29575 DVSS.n7092 DVSS.n7084 0.0333378
R29576 DVSS.n7093 DVSS.n7092 0.0333378
R29577 DVSS.n8222 DVSS.n8221 0.0333378
R29578 DVSS.n8221 DVSS.n8220 0.0333378
R29579 DVSS.n8521 DVSS.n8520 0.0333378
R29580 DVSS.n8520 DVSS.n8519 0.0333378
R29581 DVSS.n7108 DVSS.n7104 0.0333378
R29582 DVSS.n7104 DVSS.n7103 0.0333378
R29583 DVSS.n3533 DVSS.n3059 0.03245
R29584 DVSS.n3539 DVSS.n3063 0.03245
R29585 DVSS.n3536 DVSS.n3058 0.03245
R29586 DVSS.n3534 DVSS.n3064 0.03245
R29587 DVSS.n3065 DVSS.n3057 0.03245
R29588 DVSS DVSS.n4437 0.0313333
R29589 DVSS.n4837 DVSS 0.0313333
R29590 DVSS.n3878 DVSS 0.0313333
R29591 DVSS.n4992 DVSS 0.0313333
R29592 DVSS.n3541 DVSS 0.0313333
R29593 DVSS.n5383 DVSS 0.0313333
R29594 DVSS.n5679 DVSS 0.0313333
R29595 DVSS DVSS.n5507 0.0313333
R29596 DVSS DVSS.n5664 0.0313333
R29597 DVSS.n5534 DVSS 0.0313333
R29598 DVSS.n2682 DVSS 0.0313333
R29599 DVSS.n2740 DVSS 0.0313333
R29600 DVSS DVSS.n7352 0.0313333
R29601 DVSS.n7722 DVSS 0.0313333
R29602 DVSS.n8078 DVSS 0.0313333
R29603 DVSS.n8118 DVSS 0.0313333
R29604 DVSS.n3876 DVSS.n3049 0.03065
R29605 DVSS.n3874 DVSS.n3047 0.03065
R29606 DVSS.n3872 DVSS.n3050 0.03065
R29607 DVSS.n3051 DVSS.n3046 0.03065
R29608 DVSS.n7092 DVSS.n1452 0.0292293
R29609 DVSS.t3 DVSS.n1452 0.0292293
R29610 DVSS.n8221 DVSS.n1456 0.0292293
R29611 DVSS.n1456 DVSS.t3 0.0292293
R29612 DVSS.n3067 DVSS.n3059 0.0287281
R29613 DVSS.n5673 DVSS.n5671 0.0287281
R29614 DVSS.n5667 DVSS.n5666 0.0287281
R29615 DVSS.n5836 DVSS.n5835 0.0287281
R29616 DVSS.n5833 DVSS.n3043 0.0287281
R29617 DVSS.n5832 DVSS.n3055 0.0287281
R29618 DVSS.n5676 DVSS.n5675 0.0287281
R29619 DVSS.n5669 DVSS.n3258 0.0287281
R29620 DVSS.n751 DVSS.n750 0.0286081
R29621 DVSS.n9386 DVSS.n336 0.0286081
R29622 DVSS.n5899 DVSS.n5898 0.0279406
R29623 DVSS.n5898 DVSS.n5897 0.0279406
R29624 DVSS.n7152 DVSS.n7137 0.0276508
R29625 DVSS.n7152 DVSS.n7138 0.0276508
R29626 DVSS.n1534 DVSS.n1533 0.0276508
R29627 DVSS.n1536 DVSS.n1533 0.0276508
R29628 DVSS.n8204 DVSS.n1552 0.0276508
R29629 DVSS.n8204 DVSS.n8203 0.0276508
R29630 DVSS.n8197 DVSS.n1559 0.0276508
R29631 DVSS.n8197 DVSS.n8196 0.0276508
R29632 DVSS.n7065 DVSS.n6664 0.0276508
R29633 DVSS.n7065 DVSS.n6665 0.0276508
R29634 DVSS.n7131 DVSS.n7070 0.0276508
R29635 DVSS.n7131 DVSS.n7071 0.0276508
R29636 DVSS.n8246 DVSS.n8245 0.0263511
R29637 DVSS.n8249 DVSS.n1511 0.0263511
R29638 DVSS.n8255 DVSS.n1506 0.0263511
R29639 DVSS.n8266 DVSS.n8265 0.0263511
R29640 DVSS.n8271 DVSS.n8269 0.0263511
R29641 DVSS.n1489 DVSS.n1488 0.0263511
R29642 DVSS.n8291 DVSS.n1486 0.0263511
R29643 DVSS.n8287 DVSS.n1496 0.0263511
R29644 DVSS.n8281 DVSS.n1503 0.0263511
R29645 DVSS.n8325 DVSS.n8324 0.0263511
R29646 DVSS.n8327 DVSS.n1448 0.0263511
R29647 DVSS.n8235 DVSS.n8234 0.0263511
R29648 DVSS.n8237 DVSS.n1515 0.0263511
R29649 DVSS.n8226 DVSS.n1472 0.0263511
R29650 DVSS.n8307 DVSS.n1466 0.0263511
R29651 DVSS.n8311 DVSS.n8310 0.0263511
R29652 DVSS.n8314 DVSS.n1460 0.0263511
R29653 DVSS.n1186 DVSS.n1183 0.0263511
R29654 DVSS.n1184 DVSS.n1183 0.0263511
R29655 DVSS.n8448 DVSS.n1320 0.0263511
R29656 DVSS.n1385 DVSS.n1380 0.0263511
R29657 DVSS.n8472 DVSS.n8469 0.0263511
R29658 DVSS.n8478 DVSS.n1138 0.0263511
R29659 DVSS.n8478 DVSS.n1139 0.0263511
R29660 DVSS.n1131 DVSS.n1128 0.0263511
R29661 DVSS.n1129 DVSS.n1128 0.0263511
R29662 DVSS.n1288 DVSS.n1225 0.0263511
R29663 DVSS.n1283 DVSS.n1232 0.0263511
R29664 DVSS.n1237 DVSS.n1236 0.0263511
R29665 DVSS.n1241 DVSS.n1240 0.0263511
R29666 DVSS.n1263 DVSS.n1247 0.0263511
R29667 DVSS.n1258 DVSS.n1254 0.0263511
R29668 DVSS.n8456 DVSS.n1159 0.0263511
R29669 DVSS.n8368 DVSS.n8366 0.0263511
R29670 DVSS.n8376 DVSS.n8375 0.0263511
R29671 DVSS.n8385 DVSS.n8384 0.0263511
R29672 DVSS.n8352 DVSS.n1423 0.0263511
R29673 DVSS.n8492 DVSS.n1103 0.0263511
R29674 DVSS.n3871 DVSS.n3049 0.02615
R29675 DVSS.n3876 DVSS.n3047 0.02615
R29676 DVSS.n3874 DVSS.n3050 0.02615
R29677 DVSS.n3872 DVSS.n3046 0.02615
R29678 DVSS.n5836 DVSS.n3051 0.02615
R29679 DVSS.n1083 DVSS.n560 0.0256408
R29680 DVSS.n8525 DVSS.n588 0.0256408
R29681 DVSS.n4702 DVSS.n4700 0.0248
R29682 DVSS.n4700 DVSS.n4698 0.0248
R29683 DVSS.n4698 DVSS.n4696 0.0248
R29684 DVSS.n4696 DVSS.n4694 0.0248
R29685 DVSS.n4694 DVSS.n4629 0.0248
R29686 DVSS.n4690 DVSS.n4629 0.0248
R29687 DVSS.n4690 DVSS.n4689 0.0248
R29688 DVSS.n4689 DVSS.n4688 0.0248
R29689 DVSS.n4688 DVSS.n4635 0.0248
R29690 DVSS.n4684 DVSS.n4635 0.0248
R29691 DVSS.n4684 DVSS.n4683 0.0248
R29692 DVSS.n4683 DVSS.n4682 0.0248
R29693 DVSS.n4682 DVSS.n4641 0.0248
R29694 DVSS.n4678 DVSS.n4677 0.0248
R29695 DVSS.n4676 DVSS.n4648 0.0248
R29696 DVSS.n4672 DVSS.n4648 0.0248
R29697 DVSS.n4672 DVSS.n4671 0.0248
R29698 DVSS.n4671 DVSS.n4670 0.0248
R29699 DVSS.n4670 DVSS.n4654 0.0248
R29700 DVSS.n4666 DVSS.n4654 0.0248
R29701 DVSS.n4666 DVSS.n4665 0.0248
R29702 DVSS.n4665 DVSS.n4663 0.0248
R29703 DVSS.n4663 DVSS.n4661 0.0248
R29704 DVSS.n4661 DVSS.n3687 0.0248
R29705 DVSS.n4812 DVSS.n3687 0.0248
R29706 DVSS.n4039 DVSS.n4037 0.0248
R29707 DVSS.n4039 DVSS.n4035 0.0248
R29708 DVSS.n4043 DVSS.n4035 0.0248
R29709 DVSS.n4043 DVSS.n4033 0.0248
R29710 DVSS.n4047 DVSS.n4033 0.0248
R29711 DVSS.n4047 DVSS.n4031 0.0248
R29712 DVSS.n4051 DVSS.n4031 0.0248
R29713 DVSS.n4051 DVSS.n4029 0.0248
R29714 DVSS.n4055 DVSS.n4029 0.0248
R29715 DVSS.n4055 DVSS.n4027 0.0248
R29716 DVSS.n4059 DVSS.n4027 0.0248
R29717 DVSS.n4059 DVSS.n4025 0.0248
R29718 DVSS.n4063 DVSS.n4025 0.0248
R29719 DVSS.n4067 DVSS.n4066 0.0248
R29720 DVSS.n4070 DVSS.n4020 0.0248
R29721 DVSS.n4074 DVSS.n4020 0.0248
R29722 DVSS.n4074 DVSS.n4018 0.0248
R29723 DVSS.n4078 DVSS.n4018 0.0248
R29724 DVSS.n4078 DVSS.n4016 0.0248
R29725 DVSS.n4082 DVSS.n4016 0.0248
R29726 DVSS.n4082 DVSS.n4014 0.0248
R29727 DVSS.n4086 DVSS.n4014 0.0248
R29728 DVSS.n4086 DVSS.n4012 0.0248
R29729 DVSS.n4091 DVSS.n4012 0.0248
R29730 DVSS.n4091 DVSS.n3561 0.0248
R29731 DVSS.n3991 DVSS.n3990 0.0248
R29732 DVSS.n3990 DVSS.n3988 0.0248
R29733 DVSS.n3988 DVSS.n3987 0.0248
R29734 DVSS.n3987 DVSS.n3487 0.0248
R29735 DVSS.n5234 DVSS.n3487 0.0248
R29736 DVSS.n5234 DVSS.n3488 0.0248
R29737 DVSS.n5230 DVSS.n3488 0.0248
R29738 DVSS.n5230 DVSS.n5229 0.0248
R29739 DVSS.n5229 DVSS.n5228 0.0248
R29740 DVSS.n5228 DVSS.n3494 0.0248
R29741 DVSS.n5224 DVSS.n3494 0.0248
R29742 DVSS.n5224 DVSS.n5223 0.0248
R29743 DVSS.n5223 DVSS.n5222 0.0248
R29744 DVSS.n5219 DVSS.n5218 0.0248
R29745 DVSS.n5217 DVSS.n3505 0.0248
R29746 DVSS.n5213 DVSS.n3505 0.0248
R29747 DVSS.n5213 DVSS.n5212 0.0248
R29748 DVSS.n5212 DVSS.n5211 0.0248
R29749 DVSS.n5211 DVSS.n3511 0.0248
R29750 DVSS.n5207 DVSS.n3511 0.0248
R29751 DVSS.n5207 DVSS.n5206 0.0248
R29752 DVSS.n5206 DVSS.n5205 0.0248
R29753 DVSS.n5205 DVSS.n5203 0.0248
R29754 DVSS.n5203 DVSS.n5201 0.0248
R29755 DVSS.n5201 DVSS.n5199 0.0248
R29756 DVSS.n5738 DVSS.n5737 0.0248
R29757 DVSS.n5737 DVSS.n5736 0.0248
R29758 DVSS.n5736 DVSS.n3193 0.0248
R29759 DVSS.n5732 DVSS.n3193 0.0248
R29760 DVSS.n5732 DVSS.n5731 0.0248
R29761 DVSS.n5731 DVSS.n5730 0.0248
R29762 DVSS.n5730 DVSS.n3199 0.0248
R29763 DVSS.n5726 DVSS.n3199 0.0248
R29764 DVSS.n5726 DVSS.n5725 0.0248
R29765 DVSS.n5725 DVSS.n5724 0.0248
R29766 DVSS.n5724 DVSS.n3205 0.0248
R29767 DVSS.n5720 DVSS.n3205 0.0248
R29768 DVSS.n5720 DVSS.n5719 0.0248
R29769 DVSS.n5717 DVSS.n3211 0.0248
R29770 DVSS.n5713 DVSS.n5712 0.0248
R29771 DVSS.n5712 DVSS.n5711 0.0248
R29772 DVSS.n5711 DVSS.n3217 0.0248
R29773 DVSS.n5707 DVSS.n3217 0.0248
R29774 DVSS.n5707 DVSS.n5706 0.0248
R29775 DVSS.n5706 DVSS.n5705 0.0248
R29776 DVSS.n5705 DVSS.n3223 0.0248
R29777 DVSS.n5701 DVSS.n3223 0.0248
R29778 DVSS.n5701 DVSS.n5700 0.0248
R29779 DVSS.n5700 DVSS.n5699 0.0248
R29780 DVSS.n5699 DVSS.n3229 0.0248
R29781 DVSS.n5483 DVSS.n5407 0.0248
R29782 DVSS.n5479 DVSS.n5407 0.0248
R29783 DVSS.n5479 DVSS.n5478 0.0248
R29784 DVSS.n5478 DVSS.n5477 0.0248
R29785 DVSS.n5477 DVSS.n5412 0.0248
R29786 DVSS.n5473 DVSS.n5412 0.0248
R29787 DVSS.n5473 DVSS.n5472 0.0248
R29788 DVSS.n5472 DVSS.n5471 0.0248
R29789 DVSS.n5471 DVSS.n5418 0.0248
R29790 DVSS.n5467 DVSS.n5418 0.0248
R29791 DVSS.n5467 DVSS.n5466 0.0248
R29792 DVSS.n5466 DVSS.n5465 0.0248
R29793 DVSS.n5465 DVSS.n5424 0.0248
R29794 DVSS.n5461 DVSS.n5460 0.0248
R29795 DVSS.n5459 DVSS.n5431 0.0248
R29796 DVSS.n5455 DVSS.n5431 0.0248
R29797 DVSS.n5455 DVSS.n5454 0.0248
R29798 DVSS.n5454 DVSS.n5453 0.0248
R29799 DVSS.n5453 DVSS.n5437 0.0248
R29800 DVSS.n5449 DVSS.n5437 0.0248
R29801 DVSS.n5449 DVSS.n5448 0.0248
R29802 DVSS.n5448 DVSS.n5447 0.0248
R29803 DVSS.n5447 DVSS.n5444 0.0248
R29804 DVSS.n5444 DVSS.n3283 0.0248
R29805 DVSS.n5640 DVSS.n3283 0.0248
R29806 DVSS.n5629 DVSS.n5550 0.0248
R29807 DVSS.n5625 DVSS.n5550 0.0248
R29808 DVSS.n5625 DVSS.n5624 0.0248
R29809 DVSS.n5624 DVSS.n5622 0.0248
R29810 DVSS.n5622 DVSS.n5620 0.0248
R29811 DVSS.n5620 DVSS.n5618 0.0248
R29812 DVSS.n5618 DVSS.n5616 0.0248
R29813 DVSS.n5616 DVSS.n5614 0.0248
R29814 DVSS.n5614 DVSS.n5611 0.0248
R29815 DVSS.n5611 DVSS.n5610 0.0248
R29816 DVSS.n5610 DVSS.n5608 0.0248
R29817 DVSS.n5608 DVSS.n5606 0.0248
R29818 DVSS.n5606 DVSS.n5604 0.0248
R29819 DVSS.n5601 DVSS.n5599 0.0248
R29820 DVSS.n5596 DVSS.n5595 0.0248
R29821 DVSS.n5595 DVSS.n5593 0.0248
R29822 DVSS.n5593 DVSS.n5591 0.0248
R29823 DVSS.n5591 DVSS.n5589 0.0248
R29824 DVSS.n5589 DVSS.n5587 0.0248
R29825 DVSS.n5587 DVSS.n5585 0.0248
R29826 DVSS.n5585 DVSS.n5583 0.0248
R29827 DVSS.n5583 DVSS.n5580 0.0248
R29828 DVSS.n5580 DVSS.n5579 0.0248
R29829 DVSS.n5579 DVSS.n5577 0.0248
R29830 DVSS.n5577 DVSS.n2701 0.0248
R29831 DVSS.n7274 DVSS.n2651 0.0248
R29832 DVSS.n7274 DVSS.n2649 0.0248
R29833 DVSS.n7278 DVSS.n2649 0.0248
R29834 DVSS.n7278 DVSS.n2647 0.0248
R29835 DVSS.n7282 DVSS.n2647 0.0248
R29836 DVSS.n7282 DVSS.n2645 0.0248
R29837 DVSS.n7286 DVSS.n2645 0.0248
R29838 DVSS.n7286 DVSS.n2643 0.0248
R29839 DVSS.n7290 DVSS.n2643 0.0248
R29840 DVSS.n7290 DVSS.n2641 0.0248
R29841 DVSS.n7294 DVSS.n2641 0.0248
R29842 DVSS.n7294 DVSS.n2638 0.0248
R29843 DVSS.n7298 DVSS.n2638 0.0248
R29844 DVSS.n7302 DVSS.n2636 0.0248
R29845 DVSS.n7306 DVSS.n2634 0.0248
R29846 DVSS.n7306 DVSS.n2632 0.0248
R29847 DVSS.n7310 DVSS.n2632 0.0248
R29848 DVSS.n7310 DVSS.n2630 0.0248
R29849 DVSS.n7314 DVSS.n2630 0.0248
R29850 DVSS.n7314 DVSS.n2628 0.0248
R29851 DVSS.n7318 DVSS.n2628 0.0248
R29852 DVSS.n7318 DVSS.n2626 0.0248
R29853 DVSS.n7322 DVSS.n2626 0.0248
R29854 DVSS.n7322 DVSS.n2623 0.0248
R29855 DVSS.n7328 DVSS.n2623 0.0248
R29856 DVSS.n7865 DVSS.n2077 0.0248
R29857 DVSS.n7865 DVSS.n2074 0.0248
R29858 DVSS.n7869 DVSS.n2074 0.0248
R29859 DVSS.n7872 DVSS.n7869 0.0248
R29860 DVSS.n7875 DVSS.n7872 0.0248
R29861 DVSS.n7878 DVSS.n7875 0.0248
R29862 DVSS.n7881 DVSS.n7878 0.0248
R29863 DVSS.n7882 DVSS.n7881 0.0248
R29864 DVSS.n7887 DVSS.n7882 0.0248
R29865 DVSS.n7890 DVSS.n7887 0.0248
R29866 DVSS.n7893 DVSS.n7890 0.0248
R29867 DVSS.n7895 DVSS.n7893 0.0248
R29868 DVSS.n7898 DVSS.n7895 0.0248
R29869 DVSS.n7933 DVSS.n2058 0.0248
R29870 DVSS.n7932 DVSS.n7931 0.0248
R29871 DVSS.n7931 DVSS.n7906 0.0248
R29872 DVSS.n7927 DVSS.n7906 0.0248
R29873 DVSS.n7927 DVSS.n7926 0.0248
R29874 DVSS.n7926 DVSS.n7925 0.0248
R29875 DVSS.n7925 DVSS.n7912 0.0248
R29876 DVSS.n7921 DVSS.n7912 0.0248
R29877 DVSS.n7921 DVSS.n7920 0.0248
R29878 DVSS.n7920 DVSS.n7919 0.0248
R29879 DVSS.n7919 DVSS.n1872 0.0248
R29880 DVSS.n8097 DVSS.n1872 0.0248
R29881 DVSS.n7186 DVSS.n7183 0.0248
R29882 DVSS.n7186 DVSS.n7181 0.0248
R29883 DVSS.n7190 DVSS.n7181 0.0248
R29884 DVSS.n7190 DVSS.n7179 0.0248
R29885 DVSS.n7194 DVSS.n7179 0.0248
R29886 DVSS.n7194 DVSS.n7177 0.0248
R29887 DVSS.n7198 DVSS.n7177 0.0248
R29888 DVSS.n7198 DVSS.n7175 0.0248
R29889 DVSS.n7202 DVSS.n7175 0.0248
R29890 DVSS.n7202 DVSS.n7173 0.0248
R29891 DVSS.n7206 DVSS.n7173 0.0248
R29892 DVSS.n7206 DVSS.n7171 0.0248
R29893 DVSS.n7210 DVSS.n7171 0.0248
R29894 DVSS.n7214 DVSS.n7213 0.0248
R29895 DVSS.n7217 DVSS.n7166 0.0248
R29896 DVSS.n7221 DVSS.n7166 0.0248
R29897 DVSS.n7221 DVSS.n7164 0.0248
R29898 DVSS.n7225 DVSS.n7164 0.0248
R29899 DVSS.n7225 DVSS.n7162 0.0248
R29900 DVSS.n7229 DVSS.n7162 0.0248
R29901 DVSS.n7229 DVSS.n7160 0.0248
R29902 DVSS.n7233 DVSS.n7160 0.0248
R29903 DVSS.n7233 DVSS.n7158 0.0248
R29904 DVSS.n7237 DVSS.n7158 0.0248
R29905 DVSS.n7237 DVSS.n7156 0.0248
R29906 DVSS.n7247 DVSS.n6644 0.0248
R29907 DVSS.n7253 DVSS.n6644 0.0248
R29908 DVSS.n3533 DVSS.n3063 0.02435
R29909 DVSS.n3539 DVSS.n3058 0.02435
R29910 DVSS.n3536 DVSS.n3064 0.02435
R29911 DVSS.n3534 DVSS.n3057 0.02435
R29912 DVSS.n5830 DVSS.n3065 0.02435
R29913 DVSS.n9008 DVSS.n707 0.0243462
R29914 DVSS.n9010 DVSS.n707 0.0243462
R29915 DVSS.n9014 DVSS.n700 0.0243462
R29916 DVSS.n9016 DVSS.n700 0.0243462
R29917 DVSS.n9023 DVSS.n9018 0.0243462
R29918 DVSS.n9018 DVSS.n382 0.0243462
R29919 DVSS.n9383 DVSS.n384 0.0243462
R29920 DVSS.n9381 DVSS.n384 0.0243462
R29921 DVSS.n9371 DVSS.n9370 0.0243462
R29922 DVSS.n9376 DVSS.n9371 0.0243462
R29923 DVSS.n327 DVSS.n326 0.0243462
R29924 DVSS.n9541 DVSS.n327 0.0243462
R29925 DVSS.n8520 DVSS.n1081 0.0237143
R29926 DVSS.t37 DVSS.n1081 0.0237143
R29927 DVSS.n7104 DVSS.n1093 0.0237143
R29928 DVSS.n1093 DVSS.t37 0.0237143
R29929 DVSS.n9384 DVSS.n382 0.0233846
R29930 DVSS.n9384 DVSS.n9383 0.0233846
R29931 DVSS.n9389 DVSS.n378 0.0233846
R29932 DVSS.n9392 DVSS.n9389 0.0233846
R29933 DVSS.n4631 DVSS.n4628 0.0233169
R29934 DVSS.n4632 DVSS.n4631 0.0233169
R29935 DVSS.n4633 DVSS.n4632 0.0233169
R29936 DVSS.n4634 DVSS.n4633 0.0233169
R29937 DVSS.n4637 DVSS.n4634 0.0233169
R29938 DVSS.n4638 DVSS.n4637 0.0233169
R29939 DVSS.n4639 DVSS.n4638 0.0233169
R29940 DVSS.n4640 DVSS.n4639 0.0233169
R29941 DVSS.n4644 DVSS.n4640 0.0233169
R29942 DVSS.n4645 DVSS.n4644 0.0233169
R29943 DVSS.n4646 DVSS.n4645 0.0233169
R29944 DVSS.n4647 DVSS.n4646 0.0233169
R29945 DVSS.n4650 DVSS.n4647 0.0233169
R29946 DVSS.n4651 DVSS.n4650 0.0233169
R29947 DVSS.n4652 DVSS.n4651 0.0233169
R29948 DVSS.n4653 DVSS.n4652 0.0233169
R29949 DVSS.n4655 DVSS.n4653 0.0233169
R29950 DVSS.n4656 DVSS.n4655 0.0233169
R29951 DVSS.n4040 DVSS.n4036 0.0233169
R29952 DVSS.n4041 DVSS.n4040 0.0233169
R29953 DVSS.n4042 DVSS.n4041 0.0233169
R29954 DVSS.n4042 DVSS.n4032 0.0233169
R29955 DVSS.n4048 DVSS.n4032 0.0233169
R29956 DVSS.n4049 DVSS.n4048 0.0233169
R29957 DVSS.n4050 DVSS.n4049 0.0233169
R29958 DVSS.n4050 DVSS.n4028 0.0233169
R29959 DVSS.n4056 DVSS.n4028 0.0233169
R29960 DVSS.n4057 DVSS.n4056 0.0233169
R29961 DVSS.n4058 DVSS.n4057 0.0233169
R29962 DVSS.n4058 DVSS.n4024 0.0233169
R29963 DVSS.n4064 DVSS.n4024 0.0233169
R29964 DVSS.n4065 DVSS.n4064 0.0233169
R29965 DVSS.n4065 DVSS.n4021 0.0233169
R29966 DVSS.n4071 DVSS.n4021 0.0233169
R29967 DVSS.n4072 DVSS.n4071 0.0233169
R29968 DVSS.n4073 DVSS.n4072 0.0233169
R29969 DVSS.n4073 DVSS.n4017 0.0233169
R29970 DVSS.n4079 DVSS.n4017 0.0233169
R29971 DVSS.n4080 DVSS.n4079 0.0233169
R29972 DVSS.n4081 DVSS.n4080 0.0233169
R29973 DVSS.n4081 DVSS.n4013 0.0233169
R29974 DVSS.n4087 DVSS.n4013 0.0233169
R29975 DVSS.n4088 DVSS.n4087 0.0233169
R29976 DVSS.n4090 DVSS.n4088 0.0233169
R29977 DVSS.n4090 DVSS.n4089 0.0233169
R29978 DVSS.n5235 DVSS.n3486 0.0233169
R29979 DVSS.n3491 DVSS.n3486 0.0233169
R29980 DVSS.n3492 DVSS.n3491 0.0233169
R29981 DVSS.n3493 DVSS.n3492 0.0233169
R29982 DVSS.n3496 DVSS.n3493 0.0233169
R29983 DVSS.n3497 DVSS.n3496 0.0233169
R29984 DVSS.n3498 DVSS.n3497 0.0233169
R29985 DVSS.n3499 DVSS.n3498 0.0233169
R29986 DVSS.n3502 DVSS.n3499 0.0233169
R29987 DVSS.n3503 DVSS.n3502 0.0233169
R29988 DVSS.n3504 DVSS.n3503 0.0233169
R29989 DVSS.n3507 DVSS.n3504 0.0233169
R29990 DVSS.n3508 DVSS.n3507 0.0233169
R29991 DVSS.n3509 DVSS.n3508 0.0233169
R29992 DVSS.n3510 DVSS.n3509 0.0233169
R29993 DVSS.n3513 DVSS.n3510 0.0233169
R29994 DVSS.n3514 DVSS.n3513 0.0233169
R29995 DVSS.n3515 DVSS.n3514 0.0233169
R29996 DVSS.n3191 DVSS.n3190 0.0233169
R29997 DVSS.n3192 DVSS.n3191 0.0233169
R29998 DVSS.n3195 DVSS.n3192 0.0233169
R29999 DVSS.n3196 DVSS.n3195 0.0233169
R30000 DVSS.n3197 DVSS.n3196 0.0233169
R30001 DVSS.n3198 DVSS.n3197 0.0233169
R30002 DVSS.n3201 DVSS.n3198 0.0233169
R30003 DVSS.n3202 DVSS.n3201 0.0233169
R30004 DVSS.n3203 DVSS.n3202 0.0233169
R30005 DVSS.n3204 DVSS.n3203 0.0233169
R30006 DVSS.n3207 DVSS.n3204 0.0233169
R30007 DVSS.n3208 DVSS.n3207 0.0233169
R30008 DVSS.n3209 DVSS.n3208 0.0233169
R30009 DVSS.n3210 DVSS.n3209 0.0233169
R30010 DVSS.n3213 DVSS.n3210 0.0233169
R30011 DVSS.n3214 DVSS.n3213 0.0233169
R30012 DVSS.n3215 DVSS.n3214 0.0233169
R30013 DVSS.n3216 DVSS.n3215 0.0233169
R30014 DVSS.n3219 DVSS.n3216 0.0233169
R30015 DVSS.n3220 DVSS.n3219 0.0233169
R30016 DVSS.n3221 DVSS.n3220 0.0233169
R30017 DVSS.n3222 DVSS.n3221 0.0233169
R30018 DVSS.n3225 DVSS.n3222 0.0233169
R30019 DVSS.n3226 DVSS.n3225 0.0233169
R30020 DVSS.n3227 DVSS.n3226 0.0233169
R30021 DVSS.n3228 DVSS.n3227 0.0233169
R30022 DVSS.n5487 DVSS.n3228 0.0233169
R30023 DVSS.n5484 DVSS.n5406 0.0233169
R30024 DVSS.n5409 DVSS.n5406 0.0233169
R30025 DVSS.n5410 DVSS.n5409 0.0233169
R30026 DVSS.n5411 DVSS.n5410 0.0233169
R30027 DVSS.n5414 DVSS.n5411 0.0233169
R30028 DVSS.n5415 DVSS.n5414 0.0233169
R30029 DVSS.n5416 DVSS.n5415 0.0233169
R30030 DVSS.n5417 DVSS.n5416 0.0233169
R30031 DVSS.n5420 DVSS.n5417 0.0233169
R30032 DVSS.n5421 DVSS.n5420 0.0233169
R30033 DVSS.n5422 DVSS.n5421 0.0233169
R30034 DVSS.n5423 DVSS.n5422 0.0233169
R30035 DVSS.n5427 DVSS.n5423 0.0233169
R30036 DVSS.n5428 DVSS.n5427 0.0233169
R30037 DVSS.n5429 DVSS.n5428 0.0233169
R30038 DVSS.n5430 DVSS.n5429 0.0233169
R30039 DVSS.n5433 DVSS.n5430 0.0233169
R30040 DVSS.n5434 DVSS.n5433 0.0233169
R30041 DVSS.n5435 DVSS.n5434 0.0233169
R30042 DVSS.n5436 DVSS.n5435 0.0233169
R30043 DVSS.n5439 DVSS.n5436 0.0233169
R30044 DVSS.n5440 DVSS.n5439 0.0233169
R30045 DVSS.n5441 DVSS.n5440 0.0233169
R30046 DVSS.n5442 DVSS.n5441 0.0233169
R30047 DVSS.n5443 DVSS.n5442 0.0233169
R30048 DVSS.n5443 DVSS.n3285 0.0233169
R30049 DVSS.n5639 DVSS.n3285 0.0233169
R30050 DVSS.n5630 DVSS.n5549 0.0233169
R30051 DVSS.n5551 DVSS.n5549 0.0233169
R30052 DVSS.n5558 DVSS.n5557 0.0233169
R30053 DVSS.n5565 DVSS.n5564 0.0233169
R30054 DVSS.n5573 DVSS.n5572 0.0233169
R30055 DVSS.n7275 DVSS.n2650 0.0233169
R30056 DVSS.n7276 DVSS.n7275 0.0233169
R30057 DVSS.n7277 DVSS.n7276 0.0233169
R30058 DVSS.n7277 DVSS.n2646 0.0233169
R30059 DVSS.n7283 DVSS.n2646 0.0233169
R30060 DVSS.n7284 DVSS.n7283 0.0233169
R30061 DVSS.n7285 DVSS.n7284 0.0233169
R30062 DVSS.n7285 DVSS.n2642 0.0233169
R30063 DVSS.n7291 DVSS.n2642 0.0233169
R30064 DVSS.n7292 DVSS.n7291 0.0233169
R30065 DVSS.n7293 DVSS.n7292 0.0233169
R30066 DVSS.n7293 DVSS.n2637 0.0233169
R30067 DVSS.n7299 DVSS.n2637 0.0233169
R30068 DVSS.n7300 DVSS.n7299 0.0233169
R30069 DVSS.n7301 DVSS.n7300 0.0233169
R30070 DVSS.n7301 DVSS.n2633 0.0233169
R30071 DVSS.n7307 DVSS.n2633 0.0233169
R30072 DVSS.n7308 DVSS.n7307 0.0233169
R30073 DVSS.n7309 DVSS.n7308 0.0233169
R30074 DVSS.n7309 DVSS.n2629 0.0233169
R30075 DVSS.n7315 DVSS.n2629 0.0233169
R30076 DVSS.n7316 DVSS.n7315 0.0233169
R30077 DVSS.n7317 DVSS.n7316 0.0233169
R30078 DVSS.n7317 DVSS.n2625 0.0233169
R30079 DVSS.n7323 DVSS.n2625 0.0233169
R30080 DVSS.n7324 DVSS.n7323 0.0233169
R30081 DVSS.n7327 DVSS.n7324 0.0233169
R30082 DVSS.n7864 DVSS.n7862 0.0233169
R30083 DVSS.n7864 DVSS.n7863 0.0233169
R30084 DVSS.n7863 DVSS.n2075 0.0233169
R30085 DVSS.n7884 DVSS.n7883 0.0233169
R30086 DVSS.n7904 DVSS.n7903 0.0233169
R30087 DVSS.n7905 DVSS.n7904 0.0233169
R30088 DVSS.n7908 DVSS.n7905 0.0233169
R30089 DVSS.n7909 DVSS.n7908 0.0233169
R30090 DVSS.n7910 DVSS.n7909 0.0233169
R30091 DVSS.n7911 DVSS.n7910 0.0233169
R30092 DVSS.n7914 DVSS.n7911 0.0233169
R30093 DVSS.n7915 DVSS.n7914 0.0233169
R30094 DVSS.n7916 DVSS.n7915 0.0233169
R30095 DVSS.n7917 DVSS.n7916 0.0233169
R30096 DVSS.n7917 DVSS.n1871 0.0233169
R30097 DVSS.n8098 DVSS.n1871 0.0233169
R30098 DVSS.n7185 DVSS.n7184 0.0233169
R30099 DVSS.n7185 DVSS.n7180 0.0233169
R30100 DVSS.n7191 DVSS.n7180 0.0233169
R30101 DVSS.n7192 DVSS.n7191 0.0233169
R30102 DVSS.n7193 DVSS.n7192 0.0233169
R30103 DVSS.n7193 DVSS.n7176 0.0233169
R30104 DVSS.n7199 DVSS.n7176 0.0233169
R30105 DVSS.n7200 DVSS.n7199 0.0233169
R30106 DVSS.n7201 DVSS.n7200 0.0233169
R30107 DVSS.n7201 DVSS.n7172 0.0233169
R30108 DVSS.n7207 DVSS.n7172 0.0233169
R30109 DVSS.n7208 DVSS.n7207 0.0233169
R30110 DVSS.n7209 DVSS.n7208 0.0233169
R30111 DVSS.n7209 DVSS.n7168 0.0233169
R30112 DVSS.n7215 DVSS.n7168 0.0233169
R30113 DVSS.n7216 DVSS.n7215 0.0233169
R30114 DVSS.n7216 DVSS.n7165 0.0233169
R30115 DVSS.n7222 DVSS.n7165 0.0233169
R30116 DVSS.n7223 DVSS.n7222 0.0233169
R30117 DVSS.n7224 DVSS.n7223 0.0233169
R30118 DVSS.n7224 DVSS.n7161 0.0233169
R30119 DVSS.n7230 DVSS.n7161 0.0233169
R30120 DVSS.n7231 DVSS.n7230 0.0233169
R30121 DVSS.n7232 DVSS.n7231 0.0233169
R30122 DVSS.n7232 DVSS.n7157 0.0233169
R30123 DVSS.n7238 DVSS.n7157 0.0233169
R30124 DVSS.n7239 DVSS.n7238 0.0233169
R30125 DVSS.n7244 DVSS.n6645 0.0233169
R30126 DVSS.n4693 DVSS.n4692 0.0233169
R30127 DVSS.n4692 DVSS.n4691 0.0233169
R30128 DVSS.n4691 DVSS.n4630 0.0233169
R30129 DVSS.n4687 DVSS.n4630 0.0233169
R30130 DVSS.n4687 DVSS.n4686 0.0233169
R30131 DVSS.n4686 DVSS.n4685 0.0233169
R30132 DVSS.n4685 DVSS.n4636 0.0233169
R30133 DVSS.n4681 DVSS.n4636 0.0233169
R30134 DVSS.n4681 DVSS.n4680 0.0233169
R30135 DVSS.n4680 DVSS.n4679 0.0233169
R30136 DVSS.n4679 DVSS.n4642 0.0233169
R30137 DVSS.n4675 DVSS.n4642 0.0233169
R30138 DVSS.n4675 DVSS.n4674 0.0233169
R30139 DVSS.n4674 DVSS.n4673 0.0233169
R30140 DVSS.n4673 DVSS.n4649 0.0233169
R30141 DVSS.n4669 DVSS.n4649 0.0233169
R30142 DVSS.n4669 DVSS.n4668 0.0233169
R30143 DVSS.n4668 DVSS.n4667 0.0233169
R30144 DVSS.n4038 DVSS.n3705 0.0233169
R30145 DVSS.n4038 DVSS.n4034 0.0233169
R30146 DVSS.n4044 DVSS.n4034 0.0233169
R30147 DVSS.n4045 DVSS.n4044 0.0233169
R30148 DVSS.n4046 DVSS.n4045 0.0233169
R30149 DVSS.n4046 DVSS.n4030 0.0233169
R30150 DVSS.n4052 DVSS.n4030 0.0233169
R30151 DVSS.n4053 DVSS.n4052 0.0233169
R30152 DVSS.n4054 DVSS.n4053 0.0233169
R30153 DVSS.n4054 DVSS.n4026 0.0233169
R30154 DVSS.n4060 DVSS.n4026 0.0233169
R30155 DVSS.n4061 DVSS.n4060 0.0233169
R30156 DVSS.n4062 DVSS.n4061 0.0233169
R30157 DVSS.n4062 DVSS.n4022 0.0233169
R30158 DVSS.n4068 DVSS.n4022 0.0233169
R30159 DVSS.n4069 DVSS.n4068 0.0233169
R30160 DVSS.n4069 DVSS.n4019 0.0233169
R30161 DVSS.n4075 DVSS.n4019 0.0233169
R30162 DVSS.n4076 DVSS.n4075 0.0233169
R30163 DVSS.n4077 DVSS.n4076 0.0233169
R30164 DVSS.n4077 DVSS.n4015 0.0233169
R30165 DVSS.n4083 DVSS.n4015 0.0233169
R30166 DVSS.n4084 DVSS.n4083 0.0233169
R30167 DVSS.n4085 DVSS.n4084 0.0233169
R30168 DVSS.n4085 DVSS.n4011 0.0233169
R30169 DVSS.n4092 DVSS.n4011 0.0233169
R30170 DVSS.n4093 DVSS.n4092 0.0233169
R30171 DVSS.n5233 DVSS.n5232 0.0233169
R30172 DVSS.n5232 DVSS.n5231 0.0233169
R30173 DVSS.n5231 DVSS.n3490 0.0233169
R30174 DVSS.n5227 DVSS.n3490 0.0233169
R30175 DVSS.n5227 DVSS.n5226 0.0233169
R30176 DVSS.n5226 DVSS.n5225 0.0233169
R30177 DVSS.n5225 DVSS.n3495 0.0233169
R30178 DVSS.n5221 DVSS.n3495 0.0233169
R30179 DVSS.n5221 DVSS.n5220 0.0233169
R30180 DVSS.n5220 DVSS.n3501 0.0233169
R30181 DVSS.n5216 DVSS.n3501 0.0233169
R30182 DVSS.n5216 DVSS.n5215 0.0233169
R30183 DVSS.n5215 DVSS.n5214 0.0233169
R30184 DVSS.n5214 DVSS.n3506 0.0233169
R30185 DVSS.n5210 DVSS.n3506 0.0233169
R30186 DVSS.n5210 DVSS.n5209 0.0233169
R30187 DVSS.n5209 DVSS.n5208 0.0233169
R30188 DVSS.n5208 DVSS.n3512 0.0233169
R30189 DVSS.n5739 DVSS.n3189 0.0233169
R30190 DVSS.n5735 DVSS.n3189 0.0233169
R30191 DVSS.n5735 DVSS.n5734 0.0233169
R30192 DVSS.n5734 DVSS.n5733 0.0233169
R30193 DVSS.n5733 DVSS.n3194 0.0233169
R30194 DVSS.n5729 DVSS.n3194 0.0233169
R30195 DVSS.n5729 DVSS.n5728 0.0233169
R30196 DVSS.n5728 DVSS.n5727 0.0233169
R30197 DVSS.n5727 DVSS.n3200 0.0233169
R30198 DVSS.n5723 DVSS.n3200 0.0233169
R30199 DVSS.n5723 DVSS.n5722 0.0233169
R30200 DVSS.n5722 DVSS.n5721 0.0233169
R30201 DVSS.n5721 DVSS.n3206 0.0233169
R30202 DVSS.n5716 DVSS.n3206 0.0233169
R30203 DVSS.n5716 DVSS.n5715 0.0233169
R30204 DVSS.n5715 DVSS.n5714 0.0233169
R30205 DVSS.n5714 DVSS.n3212 0.0233169
R30206 DVSS.n5710 DVSS.n3212 0.0233169
R30207 DVSS.n5710 DVSS.n5709 0.0233169
R30208 DVSS.n5709 DVSS.n5708 0.0233169
R30209 DVSS.n5708 DVSS.n3218 0.0233169
R30210 DVSS.n5704 DVSS.n3218 0.0233169
R30211 DVSS.n5704 DVSS.n5703 0.0233169
R30212 DVSS.n5703 DVSS.n5702 0.0233169
R30213 DVSS.n5702 DVSS.n3224 0.0233169
R30214 DVSS.n5698 DVSS.n3224 0.0233169
R30215 DVSS.n5698 DVSS.n5697 0.0233169
R30216 DVSS.n5482 DVSS.n5481 0.0233169
R30217 DVSS.n5481 DVSS.n5480 0.0233169
R30218 DVSS.n5480 DVSS.n5408 0.0233169
R30219 DVSS.n5476 DVSS.n5408 0.0233169
R30220 DVSS.n5476 DVSS.n5475 0.0233169
R30221 DVSS.n5475 DVSS.n5474 0.0233169
R30222 DVSS.n5474 DVSS.n5413 0.0233169
R30223 DVSS.n5470 DVSS.n5413 0.0233169
R30224 DVSS.n5470 DVSS.n5469 0.0233169
R30225 DVSS.n5469 DVSS.n5468 0.0233169
R30226 DVSS.n5468 DVSS.n5419 0.0233169
R30227 DVSS.n5464 DVSS.n5419 0.0233169
R30228 DVSS.n5464 DVSS.n5463 0.0233169
R30229 DVSS.n5463 DVSS.n5462 0.0233169
R30230 DVSS.n5462 DVSS.n5425 0.0233169
R30231 DVSS.n5458 DVSS.n5425 0.0233169
R30232 DVSS.n5458 DVSS.n5457 0.0233169
R30233 DVSS.n5457 DVSS.n5456 0.0233169
R30234 DVSS.n5456 DVSS.n5432 0.0233169
R30235 DVSS.n5452 DVSS.n5432 0.0233169
R30236 DVSS.n5452 DVSS.n5451 0.0233169
R30237 DVSS.n5451 DVSS.n5450 0.0233169
R30238 DVSS.n5450 DVSS.n5438 0.0233169
R30239 DVSS.n5446 DVSS.n5438 0.0233169
R30240 DVSS.n5446 DVSS.n5445 0.0233169
R30241 DVSS.n5445 DVSS.n3282 0.0233169
R30242 DVSS.n5641 DVSS.n3282 0.0233169
R30243 DVSS.n5628 DVSS.n5627 0.0233169
R30244 DVSS.n5627 DVSS.n5626 0.0233169
R30245 DVSS.n5613 DVSS.n5612 0.0233169
R30246 DVSS.n5598 DVSS.n5597 0.0233169
R30247 DVSS.n5582 DVSS.n5581 0.0233169
R30248 DVSS.n7273 DVSS.n7272 0.0233169
R30249 DVSS.n7273 DVSS.n2648 0.0233169
R30250 DVSS.n7279 DVSS.n2648 0.0233169
R30251 DVSS.n7280 DVSS.n7279 0.0233169
R30252 DVSS.n7281 DVSS.n7280 0.0233169
R30253 DVSS.n7281 DVSS.n2644 0.0233169
R30254 DVSS.n7287 DVSS.n2644 0.0233169
R30255 DVSS.n7288 DVSS.n7287 0.0233169
R30256 DVSS.n7289 DVSS.n7288 0.0233169
R30257 DVSS.n7289 DVSS.n2640 0.0233169
R30258 DVSS.n7295 DVSS.n2640 0.0233169
R30259 DVSS.n7296 DVSS.n7295 0.0233169
R30260 DVSS.n7297 DVSS.n7296 0.0233169
R30261 DVSS.n7297 DVSS.n2635 0.0233169
R30262 DVSS.n7303 DVSS.n2635 0.0233169
R30263 DVSS.n7304 DVSS.n7303 0.0233169
R30264 DVSS.n7305 DVSS.n7304 0.0233169
R30265 DVSS.n7305 DVSS.n2631 0.0233169
R30266 DVSS.n7311 DVSS.n2631 0.0233169
R30267 DVSS.n7312 DVSS.n7311 0.0233169
R30268 DVSS.n7313 DVSS.n7312 0.0233169
R30269 DVSS.n7313 DVSS.n2627 0.0233169
R30270 DVSS.n7319 DVSS.n2627 0.0233169
R30271 DVSS.n7320 DVSS.n7319 0.0233169
R30272 DVSS.n7321 DVSS.n7320 0.0233169
R30273 DVSS.n7321 DVSS.n2622 0.0233169
R30274 DVSS.n7329 DVSS.n2622 0.0233169
R30275 DVSS.n7866 DVSS.n2076 0.0233169
R30276 DVSS.n7867 DVSS.n7866 0.0233169
R30277 DVSS.n7868 DVSS.n7867 0.0233169
R30278 DVSS.n7886 DVSS.n7885 0.0233169
R30279 DVSS.n7934 DVSS.n2057 0.0233169
R30280 DVSS.n7930 DVSS.n2057 0.0233169
R30281 DVSS.n7930 DVSS.n7929 0.0233169
R30282 DVSS.n7929 DVSS.n7928 0.0233169
R30283 DVSS.n7928 DVSS.n7907 0.0233169
R30284 DVSS.n7924 DVSS.n7907 0.0233169
R30285 DVSS.n7924 DVSS.n7923 0.0233169
R30286 DVSS.n7923 DVSS.n7922 0.0233169
R30287 DVSS.n7922 DVSS.n7913 0.0233169
R30288 DVSS.n7918 DVSS.n7913 0.0233169
R30289 DVSS.n7918 DVSS.n1873 0.0233169
R30290 DVSS.n8096 DVSS.n1873 0.0233169
R30291 DVSS.n7187 DVSS.n7182 0.0233169
R30292 DVSS.n7188 DVSS.n7187 0.0233169
R30293 DVSS.n7189 DVSS.n7188 0.0233169
R30294 DVSS.n7189 DVSS.n7178 0.0233169
R30295 DVSS.n7195 DVSS.n7178 0.0233169
R30296 DVSS.n7196 DVSS.n7195 0.0233169
R30297 DVSS.n7197 DVSS.n7196 0.0233169
R30298 DVSS.n7197 DVSS.n7174 0.0233169
R30299 DVSS.n7203 DVSS.n7174 0.0233169
R30300 DVSS.n7204 DVSS.n7203 0.0233169
R30301 DVSS.n7205 DVSS.n7204 0.0233169
R30302 DVSS.n7205 DVSS.n7170 0.0233169
R30303 DVSS.n7211 DVSS.n7170 0.0233169
R30304 DVSS.n7212 DVSS.n7211 0.0233169
R30305 DVSS.n7212 DVSS.n7167 0.0233169
R30306 DVSS.n7218 DVSS.n7167 0.0233169
R30307 DVSS.n7219 DVSS.n7218 0.0233169
R30308 DVSS.n7220 DVSS.n7219 0.0233169
R30309 DVSS.n7220 DVSS.n7163 0.0233169
R30310 DVSS.n7226 DVSS.n7163 0.0233169
R30311 DVSS.n7227 DVSS.n7226 0.0233169
R30312 DVSS.n7228 DVSS.n7227 0.0233169
R30313 DVSS.n7228 DVSS.n7159 0.0233169
R30314 DVSS.n7234 DVSS.n7159 0.0233169
R30315 DVSS.n7235 DVSS.n7234 0.0233169
R30316 DVSS.n7236 DVSS.n7235 0.0233169
R30317 DVSS.n7236 DVSS.n7155 0.0233169
R30318 DVSS.n7252 DVSS.n6646 0.0233169
R30319 DVSS.n5556 DVSS.n2295 0.0231056
R30320 DVSS.n7888 DVSS.n2065 0.0231056
R30321 DVSS.n5615 DVSS.n2325 0.0231056
R30322 DVSS.n7889 DVSS.n2047 0.0231056
R30323 DVSS.n1405 DVSS.n1401 0.0228944
R30324 DVSS.n8358 DVSS.n1364 0.0228944
R30325 DVSS.n7115 DVSS.n7114 0.0227859
R30326 DVSS.n7111 DVSS.n7079 0.0227859
R30327 DVSS.n7094 DVSS.n7090 0.0227859
R30328 DVSS.n8329 DVSS.n1443 0.0227859
R30329 DVSS.n8330 DVSS.n1441 0.0227859
R30330 DVSS.n7093 DVSS.n7090 0.0227859
R30331 DVSS.n7144 DVSS.n7141 0.0227859
R30332 DVSS.n1522 DVSS.n1520 0.0227859
R30333 DVSS.n8220 DVSS.n1524 0.0227859
R30334 DVSS.n8215 DVSS.n8214 0.0227859
R30335 DVSS.n1526 DVSS.n1524 0.0227859
R30336 DVSS.n8217 DVSS.n1529 0.0227859
R30337 DVSS.n7143 DVSS.n1520 0.0227859
R30338 DVSS.n7081 DVSS.n7079 0.0227859
R30339 DVSS.n1217 DVSS.n1216 0.0227859
R30340 DVSS.n8529 DVSS.n1079 0.0227859
R30341 DVSS.n8528 DVSS.n8527 0.0227859
R30342 DVSS.n8523 DVSS.n8521 0.0227859
R30343 DVSS.n8516 DVSS.n8515 0.0227859
R30344 DVSS.n8509 DVSS.n1085 0.0227859
R30345 DVSS.n8503 DVSS.n1087 0.0227859
R30346 DVSS.n8526 DVSS.n1080 0.0227859
R30347 DVSS.n8514 DVSS.n1084 0.0227859
R30348 DVSS.n8508 DVSS.n1086 0.0227859
R30349 DVSS.n8519 DVSS.n8518 0.0227859
R30350 DVSS.n8531 DVSS.n8530 0.0227859
R30351 DVSS.n1215 DVSS.n1079 0.0227859
R30352 DVSS.n7147 DVSS.n7140 0.0227859
R30353 DVSS.n7117 DVSS.n7116 0.0227859
R30354 DVSS.n7122 DVSS.n7121 0.0227859
R30355 DVSS.n7106 DVSS.n7086 0.0227859
R30356 DVSS.n7103 DVSS.n7088 0.0227859
R30357 DVSS.n8335 DVSS.n1439 0.0227859
R30358 DVSS.n1549 DVSS.n1547 0.0227859
R30359 DVSS.n7124 DVSS.n7075 0.0227859
R30360 DVSS.n7105 DVSS.n7086 0.0227859
R30361 DVSS.n7101 DVSS.n7088 0.0227859
R30362 DVSS.n8338 DVSS.n8337 0.0227859
R30363 DVSS.n1545 DVSS.n1544 0.0227859
R30364 DVSS.n7126 DVSS.n7073 0.0227859
R30365 DVSS.n7125 DVSS.n1151 0.0227859
R30366 DVSS.n1295 DVSS.n1294 0.0227859
R30367 DVSS.n5566 DVSS.n2286 0.0226831
R30368 DVSS.n5594 DVSS.n2316 0.0226831
R30369 DVSS.n4627 DVSS.n4617 0.0224718
R30370 DVSS.n4695 DVSS.n3771 0.0224718
R30371 DVSS.n1082 DVSS.n570 0.0222606
R30372 DVSS.n8522 DVSS.n598 0.0222606
R30373 DVSS.n7695 DVSS.n7694 0.021937
R30374 DVSS.n7379 DVSS.n7376 0.021937
R30375 DVSS DVSS.n4676 0.021875
R30376 DVSS.n4070 DVSS 0.021875
R30377 DVSS DVSS.n5217 0.021875
R30378 DVSS.n5713 DVSS 0.021875
R30379 DVSS DVSS.n5459 0.021875
R30380 DVSS.n5596 DVSS 0.021875
R30381 DVSS DVSS.n2634 0.021875
R30382 DVSS DVSS.n7932 0.021875
R30383 DVSS.n7217 DVSS 0.021875
R30384 DVSS.n5236 DVSS.n3485 0.021838
R30385 DVSS.n5574 DVSS.n2302 0.021838
R30386 DVSS.n3970 DVSS.n3489 0.021838
R30387 DVSS.n5578 DVSS.n2332 0.021838
R30388 DVSS.n8507 DVSS.n170 0.0215827
R30389 DVSS.n8513 DVSS.n209 0.0215827
R30390 DVSS.n8532 DVSS.n1066 0.0215827
R30391 DVSS.n1296 DVSS.n1195 0.0215827
R30392 DVSS.n5017 DVSS.n3516 0.0214155
R30393 DVSS.n5571 DVSS.n2283 0.0214155
R30394 DVSS.n5204 DVSS.n3182 0.0214155
R30395 DVSS.n5584 DVSS.n2313 0.0214155
R30396 DVSS.n9424 DVSS.n9422 0.0212692
R30397 DVSS.n9426 DVSS.n9424 0.0212692
R30398 DVSS.n9428 DVSS.n9426 0.0212692
R30399 DVSS.n9429 DVSS.n9428 0.0212692
R30400 DVSS.n9432 DVSS.n9429 0.0212692
R30401 DVSS.n9434 DVSS.n9432 0.0212692
R30402 DVSS.n9436 DVSS.n9434 0.0212692
R30403 DVSS.n9438 DVSS.n9436 0.0212692
R30404 DVSS.n9440 DVSS.n9438 0.0212692
R30405 DVSS.n9442 DVSS.n9440 0.0212692
R30406 DVSS.n9444 DVSS.n9442 0.0212692
R30407 DVSS.n9445 DVSS.n9444 0.0212692
R30408 DVSS.n9448 DVSS.n9445 0.0212692
R30409 DVSS.n9450 DVSS.n9448 0.0212692
R30410 DVSS.n9452 DVSS.n9450 0.0212692
R30411 DVSS.n9454 DVSS.n9452 0.0212692
R30412 DVSS.n9456 DVSS.n9454 0.0212692
R30413 DVSS.n9458 DVSS.n9456 0.0212692
R30414 DVSS.n9459 DVSS.n9458 0.0212692
R30415 DVSS.n9462 DVSS.n9459 0.0212692
R30416 DVSS.n9464 DVSS.n9462 0.0212692
R30417 DVSS.n9466 DVSS.n9464 0.0212692
R30418 DVSS.n9467 DVSS.n9466 0.0212692
R30419 DVSS.n9467 DVSS.n338 0.0212692
R30420 DVSS.n9474 DVSS.n338 0.0212692
R30421 DVSS.n9475 DVSS.n9474 0.0212692
R30422 DVSS.n9476 DVSS.n9475 0.0212692
R30423 DVSS.n9480 DVSS.n9479 0.0212692
R30424 DVSS.n9483 DVSS.n9480 0.0212692
R30425 DVSS.n9485 DVSS.n9483 0.0212692
R30426 DVSS.n9487 DVSS.n9485 0.0212692
R30427 DVSS.n9489 DVSS.n9487 0.0212692
R30428 DVSS.n9491 DVSS.n9489 0.0212692
R30429 DVSS.n9493 DVSS.n9491 0.0212692
R30430 DVSS.n9494 DVSS.n9493 0.0212692
R30431 DVSS.n9497 DVSS.n9494 0.0212692
R30432 DVSS.n9499 DVSS.n9497 0.0212692
R30433 DVSS.n9501 DVSS.n9499 0.0212692
R30434 DVSS.n9503 DVSS.n9501 0.0212692
R30435 DVSS.n9505 DVSS.n9503 0.0212692
R30436 DVSS.n9507 DVSS.n9505 0.0212692
R30437 DVSS.n9509 DVSS.n9507 0.0212692
R30438 DVSS.n9510 DVSS.n9509 0.0212692
R30439 DVSS.n9513 DVSS.n9510 0.0212692
R30440 DVSS.n9515 DVSS.n9513 0.0212692
R30441 DVSS.n9517 DVSS.n9515 0.0212692
R30442 DVSS.n9519 DVSS.n9517 0.0212692
R30443 DVSS.n9521 DVSS.n9519 0.0212692
R30444 DVSS.n9523 DVSS.n9521 0.0212692
R30445 DVSS.n9525 DVSS.n9523 0.0212692
R30446 DVSS.n9526 DVSS.n9525 0.0212692
R30447 DVSS.n9529 DVSS.n9526 0.0212692
R30448 DVSS.n9531 DVSS.n9529 0.0212692
R30449 DVSS.n9532 DVSS.n9531 0.0212692
R30450 DVSS.n9004 DVSS.n714 0.0212692
R30451 DVSS.n9537 DVSS.n332 0.0212692
R30452 DVSS.n8890 DVSS.n8888 0.0212692
R30453 DVSS.n8892 DVSS.n8890 0.0212692
R30454 DVSS.n8894 DVSS.n8892 0.0212692
R30455 DVSS.n8895 DVSS.n8894 0.0212692
R30456 DVSS.n8898 DVSS.n8895 0.0212692
R30457 DVSS.n8900 DVSS.n8898 0.0212692
R30458 DVSS.n8902 DVSS.n8900 0.0212692
R30459 DVSS.n8904 DVSS.n8902 0.0212692
R30460 DVSS.n8906 DVSS.n8904 0.0212692
R30461 DVSS.n8908 DVSS.n8906 0.0212692
R30462 DVSS.n8910 DVSS.n8908 0.0212692
R30463 DVSS.n8911 DVSS.n8910 0.0212692
R30464 DVSS.n8914 DVSS.n8911 0.0212692
R30465 DVSS.n8916 DVSS.n8914 0.0212692
R30466 DVSS.n8918 DVSS.n8916 0.0212692
R30467 DVSS.n8920 DVSS.n8918 0.0212692
R30468 DVSS.n8922 DVSS.n8920 0.0212692
R30469 DVSS.n8924 DVSS.n8922 0.0212692
R30470 DVSS.n8925 DVSS.n8924 0.0212692
R30471 DVSS.n8928 DVSS.n8925 0.0212692
R30472 DVSS.n8930 DVSS.n8928 0.0212692
R30473 DVSS.n8932 DVSS.n8930 0.0212692
R30474 DVSS.n8933 DVSS.n8932 0.0212692
R30475 DVSS.n8933 DVSS.n753 0.0212692
R30476 DVSS.n8940 DVSS.n753 0.0212692
R30477 DVSS.n8941 DVSS.n8940 0.0212692
R30478 DVSS.n8942 DVSS.n8941 0.0212692
R30479 DVSS.n8946 DVSS.n8945 0.0212692
R30480 DVSS.n8949 DVSS.n8946 0.0212692
R30481 DVSS.n8951 DVSS.n8949 0.0212692
R30482 DVSS.n8953 DVSS.n8951 0.0212692
R30483 DVSS.n8955 DVSS.n8953 0.0212692
R30484 DVSS.n8957 DVSS.n8955 0.0212692
R30485 DVSS.n8959 DVSS.n8957 0.0212692
R30486 DVSS.n8960 DVSS.n8959 0.0212692
R30487 DVSS.n8963 DVSS.n8960 0.0212692
R30488 DVSS.n8965 DVSS.n8963 0.0212692
R30489 DVSS.n8967 DVSS.n8965 0.0212692
R30490 DVSS.n8969 DVSS.n8967 0.0212692
R30491 DVSS.n8971 DVSS.n8969 0.0212692
R30492 DVSS.n8973 DVSS.n8971 0.0212692
R30493 DVSS.n8975 DVSS.n8973 0.0212692
R30494 DVSS.n8976 DVSS.n8975 0.0212692
R30495 DVSS.n8979 DVSS.n8976 0.0212692
R30496 DVSS.n8981 DVSS.n8979 0.0212692
R30497 DVSS.n8983 DVSS.n8981 0.0212692
R30498 DVSS.n8985 DVSS.n8983 0.0212692
R30499 DVSS.n8987 DVSS.n8985 0.0212692
R30500 DVSS.n8989 DVSS.n8987 0.0212692
R30501 DVSS.n8991 DVSS.n8989 0.0212692
R30502 DVSS.n8992 DVSS.n8991 0.0212692
R30503 DVSS.n8993 DVSS.n8992 0.0212692
R30504 DVSS.n8993 DVSS.n721 0.0212692
R30505 DVSS.n8999 DVSS.n721 0.0212692
R30506 DVSS.n6012 DVSS.n2759 0.0208631
R30507 DVSS.n6012 DVSS.n6011 0.0208631
R30508 DVSS.n1270 DVSS.n566 0.0207817
R30509 DVSS.n1279 DVSS.n594 0.0207817
R30510 DVSS.n4657 DVSS.n3684 0.0205704
R30511 DVSS.n5563 DVSS.n2298 0.0205704
R30512 DVSS.n4664 DVSS.n3698 0.0205704
R30513 DVSS.n5600 DVSS.n2328 0.0205704
R30514 DVSS.n8286 DVSS.n8285 0.020197
R30515 DVSS.n8285 DVSS.t3 0.020197
R30516 DVSS.n8258 DVSS.n8257 0.020197
R30517 DVSS.n8257 DVSS.t3 0.020197
R30518 DVSS.n8301 DVSS.n8300 0.020197
R30519 DVSS.n8300 DVSS.t3 0.020197
R30520 DVSS.n4813 DVSS.n3680 0.0201479
R30521 DVSS.n5559 DVSS.n2289 0.0201479
R30522 DVSS.n7879 DVSS.n2071 0.0201479
R30523 DVSS.n4811 DVSS.n4810 0.0201479
R30524 DVSS.n5609 DVSS.n2319 0.0201479
R30525 DVSS.n7880 DVSS.n2053 0.0201479
R30526 DVSS.n8258 DVSS.n8255 0.0198883
R30527 DVSS.n8259 DVSS.n8258 0.0198883
R30528 DVSS.n8287 DVSS.n8286 0.0198883
R30529 DVSS.n8286 DVSS.n8284 0.0198883
R30530 DVSS.n8301 DVSS.n1472 0.0198883
R30531 DVSS.n8302 DVSS.n8301 0.0198883
R30532 DVSS.n8467 DVSS.n1145 0.0198883
R30533 DVSS.n8468 DVSS.n8467 0.0198883
R30534 DVSS.n1277 DVSS.n1274 0.0198883
R30535 DVSS.n1274 DVSS.n1271 0.0198883
R30536 DVSS.n8380 DVSS.n8378 0.0198883
R30537 DVSS.n8385 DVSS.n8380 0.0198883
R30538 DVSS.n8884 DVSS.n784 0.019811
R30539 DVSS.n9734 DVSS.n156 0.019811
R30540 DVSS.n5555 DVSS.n2290 0.0197254
R30541 DVSS.n7891 DVSS.n2072 0.0197254
R30542 DVSS.n5617 DVSS.n2320 0.0197254
R30543 DVSS.n7892 DVSS.n2054 0.0197254
R30544 DVSS.n8897 DVSS.n8896 0.0196339
R30545 DVSS.n8913 DVSS.n8912 0.0196339
R30546 DVSS.n8927 DVSS.n8926 0.0196339
R30547 DVSS.n8943 DVSS.n752 0.0196339
R30548 DVSS.n8944 DVSS.n8943 0.0196339
R30549 DVSS.n8948 DVSS.n8947 0.0196339
R30550 DVSS.n8962 DVSS.n8961 0.0196339
R30551 DVSS.n8978 DVSS.n8977 0.0196339
R30552 DVSS.n8994 DVSS.n749 0.0196339
R30553 DVSS.n9431 DVSS.n9430 0.0196339
R30554 DVSS.n9447 DVSS.n9446 0.0196339
R30555 DVSS.n9461 DVSS.n9460 0.0196339
R30556 DVSS.n9477 DVSS.n337 0.0196339
R30557 DVSS.n9478 DVSS.n9477 0.0196339
R30558 DVSS.n9482 DVSS.n9481 0.0196339
R30559 DVSS.n9496 DVSS.n9495 0.0196339
R30560 DVSS.n9512 DVSS.n9511 0.0196339
R30561 DVSS.n9528 DVSS.n9527 0.0196339
R30562 DVSS.n5908 DVSS.n2965 0.0196339
R30563 DVSS.n5908 DVSS.n2966 0.0196339
R30564 DVSS.n5903 DVSS.n2974 0.0196339
R30565 DVSS.n5903 DVSS.n2975 0.0196339
R30566 DVSS.n7697 DVSS.n2114 0.0196339
R30567 DVSS.n7697 DVSS.n2115 0.0196339
R30568 DVSS.n7701 DVSS.n2108 0.0196339
R30569 DVSS.n7702 DVSS.n2108 0.0196339
R30570 DVSS.n1759 DVSS.n1755 0.0196339
R30571 DVSS.n1757 DVSS.n1755 0.0196339
R30572 DVSS.n8189 DVSS.n1751 0.0196339
R30573 DVSS.n6753 DVSS.n6745 0.0196339
R30574 DVSS.n8909 DVSS.n776 0.0194567
R30575 DVSS.n8944 DVSS.n737 0.0194567
R30576 DVSS.n9443 DVSS.n360 0.0194567
R30577 DVSS.n9478 DVSS.n36 0.0194567
R30578 DVSS.n5567 DVSS.n2299 0.0193028
R30579 DVSS.n7499 DVSS.n2305 0.0193028
R30580 DVSS.n5592 DVSS.n2329 0.0193028
R30581 DVSS.n7488 DVSS.n2335 0.0193028
R30582 DVSS.n8490 DVSS.n1098 0.0192795
R30583 DVSS.n8350 DVSS.n8349 0.0192795
R30584 DVSS.n8362 DVSS.n1331 0.0192795
R30585 DVSS.n8454 DVSS.n8453 0.0192795
R30586 DVSS.n8192 DVSS.n8191 0.0191034
R30587 DVSS.n6752 DVSS.n6749 0.0191034
R30588 DVSS.n8929 DVSS.n760 0.0191024
R30589 DVSS.n8964 DVSS.n742 0.0191024
R30590 DVSS.n9463 DVSS.n345 0.0191024
R30591 DVSS.n9498 DVSS.n40 0.0191024
R30592 DVSS.n4626 DVSS.n4624 0.0190915
R30593 DVSS.n4697 DVSS.n3778 0.0190915
R30594 DVSS.n3983 DVSS.n3982 0.0188803
R30595 DVSS.n3993 DVSS.n3992 0.0188803
R30596 DVSS.n8504 DVSS.n180 0.018748
R30597 DVSS.n8510 DVSS.n219 0.018748
R30598 DVSS.n8560 DVSS.n1076 0.018748
R30599 DVSS.n1297 DVSS.n1214 0.018748
R30600 DVSS.n8893 DVSS.n767 0.018748
R30601 DVSS.n8990 DVSS.n727 0.018748
R30602 DVSS.n9427 DVSS.n352 0.018748
R30603 DVSS.n9524 DVSS.n26 0.018748
R30604 DVSS.n5377 DVSS.n2946 0.018748
R30605 DVSS.n5875 DVSS.n3000 0.018748
R30606 DVSS.n6010 DVSS.n2762 0.0184577
R30607 DVSS.n3986 DVSS.n3475 0.0184577
R30608 DVSS.n5575 DVSS.n2282 0.0184577
R30609 DVSS.n3780 DVSS.n3779 0.0184577
R30610 DVSS.n3981 DVSS.n3971 0.0184577
R30611 DVSS.n5576 DVSS.n2312 0.0184577
R30612 DVSS.n8980 DVSS.n730 0.0183937
R30613 DVSS.n9514 DVSS.n29 0.0183937
R30614 DVSS.n9389 DVSS.n9388 0.0181271
R30615 DVSS.n9385 DVSS.n9384 0.0181271
R30616 DVSS.n8974 DVSS.n745 0.0180394
R30617 DVSS.n9508 DVSS.n43 0.0180394
R30618 DVSS.n5015 DVSS.n3517 0.0180352
R30619 DVSS.n5570 DVSS.n2301 0.0180352
R30620 DVSS.n5202 DVSS.n3180 0.0180352
R30621 DVSS.n5586 DVSS.n2331 0.0180352
R30622 DVSS.n6648 DVSS.n6647 0.0178648
R30623 DVSS.n5683 DVSS.n3247 0.0177222
R30624 DVSS.n5690 DVSS.n3238 0.0177222
R30625 DVSS.n5694 DVSS.n3232 0.0177222
R30626 DVSS.n5494 DVSS.n5402 0.0177222
R30627 DVSS.n5500 DVSS.n3323 0.0177222
R30628 DVSS.n5507 DVSS.n3314 0.0177222
R30629 DVSS.n5515 DVSS.n3310 0.0177222
R30630 DVSS.n5661 DVSS.n3264 0.0177222
R30631 DVSS.n5651 DVSS.n3271 0.0177222
R30632 DVSS.n3281 DVSS.n3277 0.0177222
R30633 DVSS.n5636 DVSS.n3288 0.0177222
R30634 DVSS.n5544 DVSS.n3295 0.0177222
R30635 DVSS.n5534 DVSS.n3303 0.0177222
R30636 DVSS.n5525 DVSS.n5518 0.0177222
R30637 DVSS.n2680 DVSS.n2668 0.0177222
R30638 DVSS.n2686 DVSS.n2661 0.0177222
R30639 DVSS.n2693 DVSS.n2653 0.0177222
R30640 DVSS.n7270 DVSS.n2696 0.0177222
R30641 DVSS.n2751 DVSS.n2706 0.0177222
R30642 DVSS.n2746 DVSS.n2714 0.0177222
R30643 DVSS.n2740 DVSS.n2723 0.0177222
R30644 DVSS.n2735 DVSS.n2731 0.0177222
R30645 DVSS.n7358 DVSS.n2596 0.0177222
R30646 DVSS.n7349 DVSS.n2603 0.0177222
R30647 DVSS.n7339 DVSS.n2611 0.0177222
R30648 DVSS.n2621 DVSS.n2617 0.0177222
R30649 DVSS.n7860 DVSS.n2080 0.0177222
R30650 DVSS.n7852 DVSS.n2088 0.0177222
R30651 DVSS.n7722 DVSS.n2096 0.0177222
R30652 DVSS.n7715 DVSS.n2104 0.0177222
R30653 DVSS.n8076 DVSS.n1900 0.0177222
R30654 DVSS.n8082 DVSS.n1891 0.0177222
R30655 DVSS.n8089 DVSS.n1881 0.0177222
R30656 DVSS.n8093 DVSS.n1876 0.0177222
R30657 DVSS.n8105 DVSS.n1864 0.0177222
R30658 DVSS.n8111 DVSS.n1855 0.0177222
R30659 DVSS.n8118 DVSS.n1835 0.0177222
R30660 DVSS.n1848 DVSS.n1842 0.0177222
R30661 DVSS.n8899 DVSS.n773 0.017685
R30662 DVSS.n8995 DVSS.n722 0.017685
R30663 DVSS.n9433 DVSS.n357 0.017685
R30664 DVSS.n9530 DVSS.n47 0.017685
R30665 DVSS.n5552 DVSS.n2292 0.0176127
R30666 DVSS.n7902 DVSS.n2059 0.0176127
R30667 DVSS.n5623 DVSS.n2322 0.0176127
R30668 DVSS.n7935 DVSS.n2056 0.0176127
R30669 DVSS.n1259 DVSS.n176 0.0175079
R30670 DVSS.n1264 DVSS.n215 0.0175079
R30671 DVSS.n1284 DVSS.n1072 0.0175079
R30672 DVSS.n1289 DVSS.n1201 0.0175079
R30673 DVSS.n8923 DVSS.n779 0.0173307
R30674 DVSS.n8958 DVSS.n734 0.0173307
R30675 DVSS.n9457 DVSS.n363 0.0173307
R30676 DVSS.n9492 DVSS.n33 0.0173307
R30677 DVSS.n7243 DVSS.n7240 0.0171985
R30678 DVSS.n4658 DVSS.n3682 0.0171901
R30679 DVSS.n5562 DVSS.n2287 0.0171901
R30680 DVSS.n7870 DVSS.n2069 0.0171901
R30681 DVSS.n4662 DVSS.n3696 0.0171901
R30682 DVSS.n5603 DVSS.n2317 0.0171901
R30683 DVSS.n7871 DVSS.n2051 0.0171901
R30684 DVSS.n7258 DVSS.n6015 0.0171667
R30685 DVSS.n6015 DVSS.n381 0.0171667
R30686 DVSS.n6157 DVSS.n6014 0.0171667
R30687 DVSS.n4806 DVSS.n3675 0.0170278
R30688 DVSS.n4821 DVSS.n3675 0.0170278
R30689 DVSS.n5004 DVSS.n3562 0.0170278
R30690 DVSS.n5004 DVSS.n5003 0.0170278
R30691 DVSS.n5007 DVSS.n3560 0.0170278
R30692 DVSS.n5027 DVSS.n5007 0.0170278
R30693 DVSS.n5694 DVSS.n3234 0.0170278
R30694 DVSS.n5491 DVSS.n3234 0.0170278
R30695 DVSS.n3284 DVSS.n3281 0.0170278
R30696 DVSS.n5633 DVSS.n3284 0.0170278
R30697 DVSS.n7270 DVSS.n7265 0.0170278
R30698 DVSS.n7265 DVSS.n2754 0.0170278
R30699 DVSS.n2624 DVSS.n2621 0.0170278
R30700 DVSS.n2624 DVSS.n2079 0.0170278
R30701 DVSS.n8093 DVSS.n1870 0.0170278
R30702 DVSS.n8102 DVSS.n1870 0.0170278
R30703 DVSS.n8880 DVSS.n785 0.0169764
R30704 DVSS.n8915 DVSS.n763 0.0169764
R30705 DVSS.n8950 DVSS.n739 0.0169764
R30706 DVSS.n9769 DVSS.n158 0.0169764
R30707 DVSS.n9449 DVSS.n348 0.0169764
R30708 DVSS.n9484 DVSS.n37 0.0169764
R30709 DVSS.n4814 DVSS.n3686 0.0167676
R30710 DVSS.n5560 DVSS.n2296 0.0167676
R30711 DVSS.n7876 DVSS.n2066 0.0167676
R30712 DVSS.n3694 DVSS.n3688 0.0167676
R30713 DVSS.n5607 DVSS.n2326 0.0167676
R30714 DVSS.n7877 DVSS.n2048 0.0167676
R30715 DVSS.n8907 DVSS.n764 0.016622
R30716 DVSS.n9441 DVSS.n349 0.016622
R30717 DVSS.n5554 DVSS.n2294 0.0163451
R30718 DVSS.n2073 DVSS.n2064 0.0163451
R30719 DVSS.n9394 DVSS.n374 0.0163451
R30720 DVSS.n9390 DVSS.n375 0.0163451
R30721 DVSS.n5619 DVSS.n2324 0.0163451
R30722 DVSS.n7894 DVSS.n2046 0.0163451
R30723 DVSS.n608 DVSS.n603 0.0163451
R30724 DVSS.n9129 DVSS.n606 0.0163451
R30725 DVSS.n7615 DVSS.n2210 0.0162677
R30726 DVSS.n7557 DVSS.n2252 0.0162677
R30727 DVSS.n7453 DVSS.n2400 0.0162677
R30728 DVSS.n7418 DVSS.n2464 0.0162677
R30729 DVSS.n7398 DVSS.n2521 0.0162677
R30730 DVSS.n8931 DVSS.n780 0.0162677
R30731 DVSS.n8966 DVSS.n733 0.0162677
R30732 DVSS.n7657 DVSS.n2176 0.0162677
R30733 DVSS.n9465 DVSS.n364 0.0162677
R30734 DVSS.n9500 DVSS.n32 0.0162677
R30735 DVSS.n4943 DVSS.n4918 0.0162677
R30736 DVSS.n5919 DVSS.n2919 0.0162677
R30737 DVSS.n4450 DVSS.n3853 0.0162677
R30738 DVSS.n5868 DVSS.n3023 0.0162677
R30739 DVSS.n1274 DVSS.n1273 0.0162576
R30740 DVSS.n1273 DVSS.t37 0.0162576
R30741 DVSS.n8467 DVSS.n8466 0.0162576
R30742 DVSS.n8466 DVSS.t37 0.0162576
R30743 DVSS.n8380 DVSS.n8379 0.0162576
R30744 DVSS.n8379 DVSS.t37 0.0162576
R30745 DVSS.n3672 DVSS.n3668 0.0159225
R30746 DVSS.n4822 DVSS.n3674 0.0159225
R30747 DVSS.n3676 DVSS.n3671 0.0159225
R30748 DVSS.n4819 DVSS.n4818 0.0159225
R30749 DVSS.n5198 DVSS.n5197 0.0159225
R30750 DVSS.n5568 DVSS.n2285 0.0159225
R30751 DVSS.n3706 DVSS.n3693 0.0159225
R30752 DVSS.n4805 DVSS.n3701 0.0159225
R30753 DVSS.n3708 DVSS.n3692 0.0159225
R30754 DVSS.n4808 DVSS.n3702 0.0159225
R30755 DVSS.n3519 DVSS.n3185 0.0159225
R30756 DVSS.n5590 DVSS.n2315 0.0159225
R30757 DVSS.n8891 DVSS.n772 0.0159134
R30758 DVSS.n8988 DVSS.n748 0.0159134
R30759 DVSS.n9425 DVSS.n356 0.0159134
R30760 DVSS.n9522 DVSS.n46 0.0159134
R30761 DVSS.n5375 DVSS.n2954 0.0159134
R30762 DVSS.n5873 DVSS.n3012 0.0159134
R30763 DVSS.n4625 DVSS.n4618 0.0157113
R30764 DVSS.n4699 DVSS.n3772 0.0157113
R30765 DVSS.n2827 DVSS.n2826 0.0155591
R30766 DVSS.n6007 DVSS.n2770 0.0155591
R30767 DVSS.n3743 DVSS.n3742 0.0155591
R30768 DVSS.n4594 DVSS.n3793 0.0155591
R30769 DVSS.n8982 DVSS.n746 0.0155591
R30770 DVSS.n3824 DVSS.n3823 0.0155591
R30771 DVSS.n2858 DVSS.n2857 0.0155591
R30772 DVSS.n9516 DVSS.n44 0.0155591
R30773 DVSS.n2887 DVSS.n2886 0.0155591
R30774 DVSS.n5911 DVSS.n2956 0.0155591
R30775 DVSS.n4460 DVSS.n4459 0.0155591
R30776 DVSS.n5880 DVSS.n2993 0.0155591
R30777 DVSS.n4745 DVSS.n2761 0.0155
R30778 DVSS.n3984 DVSS.n3483 0.0155
R30779 DVSS.n5022 DVSS.n5014 0.0155
R30780 DVSS.n5028 DVSS.n5019 0.0155
R30781 DVSS.n5024 DVSS.n5013 0.0155
R30782 DVSS.n5026 DVSS.n5020 0.0155
R30783 DVSS.n5030 DVSS.n5012 0.0155
R30784 DVSS.n4602 DVSS.n3776 0.0155
R30785 DVSS.n3989 DVSS.n3979 0.0155
R30786 DVSS.n3520 DVSS.n3178 0.0155
R30787 DVSS.n3559 DVSS.n3186 0.0155
R30788 DVSS.n3522 DVSS.n3177 0.0155
R30789 DVSS.n3556 DVSS.n3187 0.0155
R30790 DVSS.n3188 DVSS.n3176 0.0155
R30791 DVSS.n5889 DVSS.n5883 0.0155
R30792 DVSS.n5895 DVSS.n2982 0.0155
R30793 DVSS.n2585 DVSS.n2579 0.0155
R30794 DVSS.n7365 DVSS.n2588 0.0155
R30795 DVSS.n8067 DVSS.n8065 0.0155
R30796 DVSS.n8939 DVSS.n8938 0.0152047
R30797 DVSS.n8972 DVSS.n731 0.0152047
R30798 DVSS.n9473 DVSS.n9472 0.0152047
R30799 DVSS.n9506 DVSS.n30 0.0152047
R30800 DVSS.n4932 DVSS.n4916 0.0152047
R30801 DVSS.n2932 DVSS.n2914 0.0152047
R30802 DVSS.n4447 DVSS.n3851 0.0152047
R30803 DVSS.n5855 DVSS.n3018 0.0152047
R30804 DVSS.n4620 DVSS.n2764 0.0150775
R30805 DVSS.n3985 DVSS.n3484 0.0150775
R30806 DVSS.n2700 DVSS.n2303 0.0150775
R30807 DVSS.n4756 DVSS.n4606 0.0150775
R30808 DVSS.n4104 DVSS.n3980 0.0150775
R30809 DVSS.n2699 DVSS.n2333 0.0150775
R30810 DVSS.n4704 DVSS.n4703 0.0148662
R30811 DVSS.n4701 DVSS.n3773 0.0148662
R30812 DVSS.n8901 DVSS.n766 0.0148504
R30813 DVSS.n8998 DVSS.n8997 0.0148504
R30814 DVSS.n9435 DVSS.n351 0.0148504
R30815 DVSS.n48 DVSS.n25 0.0148504
R30816 DVSS.n5002 DVSS.n3481 0.0146549
R30817 DVSS.n3566 DVSS.n3479 0.0146549
R30818 DVSS.n3564 DVSS.n3482 0.0146549
R30819 DVSS.n5000 DVSS.n3478 0.0146549
R30820 DVSS.n5018 DVSS.n3518 0.0146549
R30821 DVSS.n5569 DVSS.n2284 0.0146549
R30822 DVSS.n4098 DVSS.n3977 0.0146549
R30823 DVSS.n4097 DVSS.n3975 0.0146549
R30824 DVSS.n4096 DVSS.n3978 0.0146549
R30825 DVSS.n4101 DVSS.n3974 0.0146549
R30826 DVSS.n5200 DVSS.n3183 0.0146549
R30827 DVSS.n5588 DVSS.n2314 0.0146549
R30828 DVSS.n7137 DVSS.n7136 0.0145346
R30829 DVSS.n7154 DVSS.n6649 0.0145346
R30830 DVSS.n7251 DVSS.n6648 0.0145346
R30831 DVSS.n7251 DVSS.n7250 0.0145346
R30832 DVSS.n7136 DVSS.n7135 0.0145346
R30833 DVSS.n7138 DVSS.n6649 0.0145346
R30834 DVSS.n7242 DVSS.n7241 0.0145346
R30835 DVSS.n1535 DVSS.n1534 0.0145346
R30836 DVSS.n8208 DVSS.n1532 0.0145346
R30837 DVSS.n8210 DVSS.n1535 0.0145346
R30838 DVSS.n1536 DVSS.n1532 0.0145346
R30839 DVSS.n7241 DVSS.n7240 0.0145346
R30840 DVSS.n1552 DVSS.n1540 0.0145346
R30841 DVSS.n8200 DVSS.n1551 0.0145346
R30842 DVSS.n1559 DVSS.n1554 0.0145346
R30843 DVSS.n8193 DVSS.n1558 0.0145346
R30844 DVSS.n8187 DVSS.n1561 0.0145346
R30845 DVSS.n8188 DVSS.n8186 0.0145346
R30846 DVSS.n8206 DVSS.n1540 0.0145346
R30847 DVSS.n8199 DVSS.n1554 0.0145346
R30848 DVSS.n8196 DVSS.n1558 0.0145346
R30849 DVSS.n8203 DVSS.n1551 0.0145346
R30850 DVSS.n8188 DVSS.n8187 0.0145346
R30851 DVSS.n8191 DVSS.n1561 0.0145346
R30852 DVSS.n4476 DVSS.n4463 0.0145346
R30853 DVSS.n4463 DVSS.n4462 0.0145346
R30854 DVSS.n4472 DVSS.n4464 0.0145346
R30855 DVSS.n4465 DVSS.n4464 0.0145346
R30856 DVSS.n4468 DVSS.n4467 0.0145346
R30857 DVSS.n4469 DVSS.n4468 0.0145346
R30858 DVSS.n3797 DVSS.n3795 0.0145346
R30859 DVSS.n4591 DVSS.n3795 0.0145346
R30860 DVSS.n4592 DVSS.n3794 0.0145346
R30861 DVSS.n3794 DVSS.n3791 0.0145346
R30862 DVSS.n4597 DVSS.n3790 0.0145346
R30863 DVSS.n3790 DVSS.n3789 0.0145346
R30864 DVSS.n3787 DVSS.n3786 0.0145346
R30865 DVSS.n3786 DVSS.n3785 0.0145346
R30866 DVSS.n4605 DVSS.n4600 0.0145346
R30867 DVSS.n4603 DVSS.n4601 0.0145346
R30868 DVSS.n4601 DVSS.n3784 0.0145346
R30869 DVSS.n6011 DVSS.n2760 0.0145346
R30870 DVSS.n2765 DVSS.n2763 0.0145346
R30871 DVSS.n2767 DVSS.n2763 0.0145346
R30872 DVSS.n2772 DVSS.n2769 0.0145346
R30873 DVSS.n2774 DVSS.n2772 0.0145346
R30874 DVSS.n2779 DVSS.n2771 0.0145346
R30875 DVSS.n2776 DVSS.n2771 0.0145346
R30876 DVSS.n2904 DVSS.n2903 0.0145346
R30877 DVSS.n2903 DVSS.n2902 0.0145346
R30878 DVSS.n2900 DVSS.n2899 0.0145346
R30879 DVSS.n2899 DVSS.n2898 0.0145346
R30880 DVSS.n2908 DVSS.n2897 0.0145346
R30881 DVSS.n2897 DVSS.n2896 0.0145346
R30882 DVSS.n2894 DVSS.n2893 0.0145346
R30883 DVSS.n2893 DVSS.n2892 0.0145346
R30884 DVSS.n5926 DVSS.n5925 0.0145346
R30885 DVSS.n5925 DVSS.n2891 0.0145346
R30886 DVSS.n4473 DVSS.n4472 0.0145346
R30887 DVSS.n4467 DVSS.n4466 0.0145346
R30888 DVSS.n3798 DVSS.n3797 0.0145346
R30889 DVSS.n4593 DVSS.n4592 0.0145346
R30890 DVSS.n4597 DVSS.n4596 0.0145346
R30891 DVSS.n3788 DVSS.n3787 0.0145346
R30892 DVSS.n4604 DVSS.n4603 0.0145346
R30893 DVSS.n2766 DVSS.n2765 0.0145346
R30894 DVSS.n6008 DVSS.n2769 0.0145346
R30895 DVSS.n2779 DVSS.n2775 0.0145346
R30896 DVSS.n2904 DVSS.n2777 0.0145346
R30897 DVSS.n2901 DVSS.n2900 0.0145346
R30898 DVSS.n2908 DVSS.n2907 0.0145346
R30899 DVSS.n2895 DVSS.n2894 0.0145346
R30900 DVSS.n4466 DVSS.n4465 0.0145346
R30901 DVSS.n4470 DVSS.n4469 0.0145346
R30902 DVSS.n4593 DVSS.n4591 0.0145346
R30903 DVSS.n4595 DVSS.n3791 0.0145346
R30904 DVSS.n3789 DVSS.n3788 0.0145346
R30905 DVSS.n4599 DVSS.n3785 0.0145346
R30906 DVSS.n4605 DVSS.n4604 0.0145346
R30907 DVSS.n3784 DVSS.n2759 0.0145346
R30908 DVSS.n2766 DVSS.n2760 0.0145346
R30909 DVSS.n6009 DVSS.n2767 0.0145346
R30910 DVSS.n2775 DVSS.n2774 0.0145346
R30911 DVSS.n6006 DVSS.n2776 0.0145346
R30912 DVSS.n2902 DVSS.n2901 0.0145346
R30913 DVSS.n2906 DVSS.n2898 0.0145346
R30914 DVSS.n2896 DVSS.n2895 0.0145346
R30915 DVSS.n2910 DVSS.n2892 0.0145346
R30916 DVSS.n5923 DVSS.n2891 0.0145346
R30917 DVSS.n5927 DVSS.n5926 0.0145346
R30918 DVSS.n6750 DVSS.n6748 0.0145346
R30919 DVSS.n6751 DVSS.n6750 0.0145346
R30920 DVSS.n6664 DVSS.n6663 0.0145346
R30921 DVSS.n7067 DVSS.n6658 0.0145346
R30922 DVSS.n7070 DVSS.n7069 0.0145346
R30923 DVSS.n7133 DVSS.n6654 0.0145346
R30924 DVSS.n6663 DVSS.n6662 0.0145346
R30925 DVSS.n7069 DVSS.n7068 0.0145346
R30926 DVSS.n7071 DVSS.n6654 0.0145346
R30927 DVSS.n6665 DVSS.n6658 0.0145346
R30928 DVSS.n6752 DVSS.n6751 0.0145346
R30929 DVSS.n4477 DVSS.n4476 0.0145346
R30930 DVSS.n4474 DVSS.n4462 0.0145346
R30931 DVSS.n6748 DVSS.n6747 0.0145346
R30932 DVSS.n8921 DVSS.n761 0.0144961
R30933 DVSS.n8956 DVSS.n741 0.0144961
R30934 DVSS.n9455 DVSS.n346 0.0144961
R30935 DVSS.n9490 DVSS.n39 0.0144961
R30936 DVSS.n5553 DVSS.n2293 0.0142324
R30937 DVSS.n7899 DVSS.n2063 0.0142324
R30938 DVSS.n5621 DVSS.n2323 0.0142324
R30939 DVSS.n7897 DVSS.n2045 0.0142324
R30940 DVSS.n8917 DVSS.n777 0.0141417
R30941 DVSS.n8952 DVSS.n736 0.0141417
R30942 DVSS.n9451 DVSS.n361 0.0141417
R30943 DVSS.n9486 DVSS.n35 0.0141417
R30944 DVSS.n4748 DVSS.n2762 0.0140606
R30945 DVSS.n4704 DVSS.n4619 0.0140606
R30946 DVSS.n4816 DVSS.n4815 0.0140606
R30947 DVSS.n3982 DVSS.n3477 0.0140606
R30948 DVSS.n5014 DVSS.n5009 0.0140606
R30949 DVSS.n5488 DVSS.n5403 0.0140606
R30950 DVSS.n5493 DVSS.n5486 0.0140606
R30951 DVSS.n5492 DVSS.n5404 0.0140606
R30952 DVSS.n5485 DVSS.n5405 0.0140606
R30953 DVSS.n5638 DVSS.n5637 0.0140606
R30954 DVSS.n5635 DVSS.n5632 0.0140606
R30955 DVSS.n5634 DVSS.n3289 0.0140606
R30956 DVSS.n5631 DVSS.n5548 0.0140606
R30957 DVSS.n7499 DVSS.n2304 0.0140606
R30958 DVSS.n2752 DVSS.n2305 0.0140606
R30959 DVSS.n2750 DVSS.n2705 0.0140606
R30960 DVSS.n2708 DVSS.n2703 0.0140606
R30961 DVSS.n2707 DVSS.n2704 0.0140606
R30962 DVSS.n7326 DVSS.n2081 0.0140606
R30963 DVSS.n7859 DVSS.n7857 0.0140606
R30964 DVSS.n7858 DVSS.n2082 0.0140606
R30965 DVSS.n7861 DVSS.n2078 0.0140606
R30966 DVSS.n8099 DVSS.n1865 0.0140606
R30967 DVSS.n8104 DVSS.n1869 0.0140606
R30968 DVSS.n8103 DVSS.n1866 0.0140606
R30969 DVSS.n1868 DVSS.n1867 0.0140606
R30970 DVSS.n1412 DVSS.n1403 0.0140606
R30971 DVSS.n1413 DVSS.n1412 0.0140606
R30972 DVSS.n8389 DVSS.n1402 0.0140606
R30973 DVSS.n8390 DVSS.n8389 0.0140606
R30974 DVSS.n1409 DVSS.n1400 0.0140606
R30975 DVSS.n1410 DVSS.n1409 0.0140606
R30976 DVSS.n1406 DVSS.n1399 0.0140606
R30977 DVSS.n1407 DVSS.n1406 0.0140606
R30978 DVSS.n9150 DVSS.n568 0.0140606
R30979 DVSS.n9149 DVSS.n582 0.0140606
R30980 DVSS.n582 DVSS.n565 0.0140606
R30981 DVSS.n9148 DVSS.n581 0.0140606
R30982 DVSS.n581 DVSS.n564 0.0140606
R30983 DVSS.n9147 DVSS.n580 0.0140606
R30984 DVSS.n580 DVSS.n563 0.0140606
R30985 DVSS.n9146 DVSS.n579 0.0140606
R30986 DVSS.n579 DVSS.n562 0.0140606
R30987 DVSS.n9145 DVSS.n561 0.0140606
R30988 DVSS.n9151 DVSS.n9143 0.0140606
R30989 DVSS.n9143 DVSS.n571 0.0140606
R30990 DVSS.n9152 DVSS.n9144 0.0140606
R30991 DVSS.n9144 DVSS.n572 0.0140606
R30992 DVSS.n9155 DVSS.n9154 0.0140606
R30993 DVSS.n9155 DVSS.n573 0.0140606
R30994 DVSS.n9157 DVSS.n574 0.0140606
R30995 DVSS.n9158 DVSS.n9157 0.0140606
R30996 DVSS.n9391 DVSS.n373 0.0140606
R30997 DVSS.n376 DVSS.n372 0.0140606
R30998 DVSS.n9198 DVSS.n518 0.0140606
R30999 DVSS.n518 DVSS.n517 0.0140606
R31000 DVSS.n9199 DVSS.n520 0.0140606
R31001 DVSS.n520 DVSS.n519 0.0140606
R31002 DVSS.n9200 DVSS.n522 0.0140606
R31003 DVSS.n522 DVSS.n521 0.0140606
R31004 DVSS.n9201 DVSS.n524 0.0140606
R31005 DVSS.n524 DVSS.n523 0.0140606
R31006 DVSS.n9202 DVSS.n526 0.0140606
R31007 DVSS.n526 DVSS.n525 0.0140606
R31008 DVSS.n9203 DVSS.n528 0.0140606
R31009 DVSS.n528 DVSS.n527 0.0140606
R31010 DVSS.n9204 DVSS.n530 0.0140606
R31011 DVSS.n530 DVSS.n529 0.0140606
R31012 DVSS.n9205 DVSS.n532 0.0140606
R31013 DVSS.n532 DVSS.n531 0.0140606
R31014 DVSS.n9206 DVSS.n534 0.0140606
R31015 DVSS.n534 DVSS.n533 0.0140606
R31016 DVSS.n9207 DVSS.n536 0.0140606
R31017 DVSS.n536 DVSS.n535 0.0140606
R31018 DVSS.n9211 DVSS.n9209 0.0140606
R31019 DVSS.n9211 DVSS.n9210 0.0140606
R31020 DVSS.n9213 DVSS.n501 0.0140606
R31021 DVSS.n9216 DVSS.n9215 0.0140606
R31022 DVSS.n9217 DVSS.n9216 0.0140606
R31023 DVSS.n9220 DVSS.n9219 0.0140606
R31024 DVSS.n9221 DVSS.n9220 0.0140606
R31025 DVSS.n9224 DVSS.n9223 0.0140606
R31026 DVSS.n9225 DVSS.n9224 0.0140606
R31027 DVSS.n9228 DVSS.n9227 0.0140606
R31028 DVSS.n9229 DVSS.n9228 0.0140606
R31029 DVSS.n9232 DVSS.n9231 0.0140606
R31030 DVSS.n9233 DVSS.n9232 0.0140606
R31031 DVSS.n9236 DVSS.n9235 0.0140606
R31032 DVSS.n9237 DVSS.n9236 0.0140606
R31033 DVSS.n9240 DVSS.n9239 0.0140606
R31034 DVSS.n9241 DVSS.n9240 0.0140606
R31035 DVSS.n9244 DVSS.n9243 0.0140606
R31036 DVSS.n9245 DVSS.n9244 0.0140606
R31037 DVSS.n9248 DVSS.n9247 0.0140606
R31038 DVSS.n9249 DVSS.n9248 0.0140606
R31039 DVSS.n9252 DVSS.n9251 0.0140606
R31040 DVSS.n9253 DVSS.n9252 0.0140606
R31041 DVSS.n9256 DVSS.n9255 0.0140606
R31042 DVSS.n9257 DVSS.n9256 0.0140606
R31043 DVSS.n9259 DVSS.n386 0.0140606
R31044 DVSS.n388 DVSS.n387 0.0140606
R31045 DVSS.n9380 DVSS.n385 0.0140606
R31046 DVSS.n9379 DVSS.n383 0.0140606
R31047 DVSS.n4815 DVSS.n3680 0.0140606
R31048 DVSS.n4999 DVSS.n3477 0.0140606
R31049 DVSS.n5197 DVSS.n5009 0.0140606
R31050 DVSS.n1415 DVSS.n1403 0.0140606
R31051 DVSS.n1413 DVSS.n1411 0.0140606
R31052 DVSS.n1411 DVSS.n1402 0.0140606
R31053 DVSS.n8391 DVSS.n8390 0.0140606
R31054 DVSS.n8387 DVSS.n1400 0.0140606
R31055 DVSS.n1410 DVSS.n1408 0.0140606
R31056 DVSS.n1408 DVSS.n1399 0.0140606
R31057 DVSS.n1407 DVSS.n1143 0.0140606
R31058 DVSS.n3782 DVSS.n3779 0.0140606
R31059 DVSS.n3781 DVSS.n3773 0.0140606
R31060 DVSS.n3700 DVSS.n3689 0.0140606
R31061 DVSS.n3993 DVSS.n3973 0.0140606
R31062 DVSS.n3184 DVSS.n3178 0.0140606
R31063 DVSS.n5696 DVSS.n5695 0.0140606
R31064 DVSS.n5693 DVSS.n3237 0.0140606
R31065 DVSS.n5692 DVSS.n3233 0.0140606
R31066 DVSS.n3236 DVSS.n3235 0.0140606
R31067 DVSS.n5643 DVSS.n5642 0.0140606
R31068 DVSS.n3280 DVSS.n3276 0.0140606
R31069 DVSS.n3279 DVSS.n3274 0.0140606
R31070 DVSS.n3278 DVSS.n3275 0.0140606
R31071 DVSS.n7488 DVSS.n2334 0.0140606
R31072 DVSS.n2697 DVSS.n2335 0.0140606
R31073 DVSS.n7269 DVSS.n7267 0.0140606
R31074 DVSS.n7268 DVSS.n2698 0.0140606
R31075 DVSS.n7271 DVSS.n2652 0.0140606
R31076 DVSS.n7331 DVSS.n7330 0.0140606
R31077 DVSS.n2620 DVSS.n2616 0.0140606
R31078 DVSS.n2619 DVSS.n2614 0.0140606
R31079 DVSS.n2618 DVSS.n2615 0.0140606
R31080 DVSS.n8095 DVSS.n8094 0.0140606
R31081 DVSS.n8092 DVSS.n1880 0.0140606
R31082 DVSS.n8091 DVSS.n1877 0.0140606
R31083 DVSS.n1879 DVSS.n1878 0.0140606
R31084 DVSS.n1376 DVSS.n1366 0.0140606
R31085 DVSS.n1391 DVSS.n1366 0.0140606
R31086 DVSS.n1375 DVSS.n1365 0.0140606
R31087 DVSS.n1390 DVSS.n1365 0.0140606
R31088 DVSS.n1374 DVSS.n1363 0.0140606
R31089 DVSS.n1389 DVSS.n1363 0.0140606
R31090 DVSS.n1373 DVSS.n1362 0.0140606
R31091 DVSS.n8401 DVSS.n1362 0.0140606
R31092 DVSS.n604 DVSS.n596 0.0140606
R31093 DVSS.n616 DVSS.n615 0.0140606
R31094 DVSS.n616 DVSS.n593 0.0140606
R31095 DVSS.n9112 DVSS.n614 0.0140606
R31096 DVSS.n614 DVSS.n592 0.0140606
R31097 DVSS.n9114 DVSS.n613 0.0140606
R31098 DVSS.n613 DVSS.n591 0.0140606
R31099 DVSS.n9116 DVSS.n612 0.0140606
R31100 DVSS.n612 DVSS.n590 0.0140606
R31101 DVSS.n9118 DVSS.n589 0.0140606
R31102 DVSS.n9121 DVSS.n9120 0.0140606
R31103 DVSS.n9121 DVSS.n599 0.0140606
R31104 DVSS.n9123 DVSS.n9122 0.0140606
R31105 DVSS.n9123 DVSS.n600 0.0140606
R31106 DVSS.n9125 DVSS.n9124 0.0140606
R31107 DVSS.n9125 DVSS.n601 0.0140606
R31108 DVSS.n9127 DVSS.n9126 0.0140606
R31109 DVSS.n9127 DVSS.n602 0.0140606
R31110 DVSS.n8868 DVSS.n8867 0.0140606
R31111 DVSS.n8866 DVSS.n8862 0.0140606
R31112 DVSS.n9050 DVSS.n9040 0.0140606
R31113 DVSS.n9040 DVSS.n649 0.0140606
R31114 DVSS.n9051 DVSS.n9041 0.0140606
R31115 DVSS.n9041 DVSS.n650 0.0140606
R31116 DVSS.n9052 DVSS.n9042 0.0140606
R31117 DVSS.n9042 DVSS.n651 0.0140606
R31118 DVSS.n9053 DVSS.n9043 0.0140606
R31119 DVSS.n9043 DVSS.n652 0.0140606
R31120 DVSS.n9054 DVSS.n9044 0.0140606
R31121 DVSS.n9044 DVSS.n653 0.0140606
R31122 DVSS.n9055 DVSS.n9045 0.0140606
R31123 DVSS.n9045 DVSS.n654 0.0140606
R31124 DVSS.n9056 DVSS.n9046 0.0140606
R31125 DVSS.n9046 DVSS.n655 0.0140606
R31126 DVSS.n9057 DVSS.n9047 0.0140606
R31127 DVSS.n9047 DVSS.n656 0.0140606
R31128 DVSS.n9058 DVSS.n9048 0.0140606
R31129 DVSS.n9048 DVSS.n657 0.0140606
R31130 DVSS.n9059 DVSS.n9049 0.0140606
R31131 DVSS.n9049 DVSS.n658 0.0140606
R31132 DVSS.n9062 DVSS.n9061 0.0140606
R31133 DVSS.n9062 DVSS.n659 0.0140606
R31134 DVSS.n9064 DVSS.n660 0.0140606
R31135 DVSS.n677 DVSS.n661 0.0140606
R31136 DVSS.n677 DVSS.n676 0.0140606
R31137 DVSS.n8778 DVSS.n679 0.0140606
R31138 DVSS.n679 DVSS.n678 0.0140606
R31139 DVSS.n8779 DVSS.n681 0.0140606
R31140 DVSS.n681 DVSS.n680 0.0140606
R31141 DVSS.n8780 DVSS.n683 0.0140606
R31142 DVSS.n683 DVSS.n682 0.0140606
R31143 DVSS.n8781 DVSS.n685 0.0140606
R31144 DVSS.n685 DVSS.n684 0.0140606
R31145 DVSS.n8782 DVSS.n687 0.0140606
R31146 DVSS.n687 DVSS.n686 0.0140606
R31147 DVSS.n8783 DVSS.n689 0.0140606
R31148 DVSS.n689 DVSS.n688 0.0140606
R31149 DVSS.n8784 DVSS.n691 0.0140606
R31150 DVSS.n691 DVSS.n690 0.0140606
R31151 DVSS.n8785 DVSS.n693 0.0140606
R31152 DVSS.n693 DVSS.n692 0.0140606
R31153 DVSS.n8786 DVSS.n695 0.0140606
R31154 DVSS.n695 DVSS.n694 0.0140606
R31155 DVSS.n8787 DVSS.n697 0.0140606
R31156 DVSS.n697 DVSS.n696 0.0140606
R31157 DVSS.n9025 DVSS.n698 0.0140606
R31158 DVSS.n9019 DVSS.n699 0.0140606
R31159 DVSS.n9022 DVSS.n9021 0.0140606
R31160 DVSS.n9020 DVSS.n9017 0.0140606
R31161 DVSS.n4810 DVSS.n3689 0.0140606
R31162 DVSS.n4102 DVSS.n3973 0.0140606
R31163 DVSS.n3185 DVSS.n3184 0.0140606
R31164 DVSS.n1376 DVSS.n1368 0.0140606
R31165 DVSS.n1391 DVSS.n1369 0.0140606
R31166 DVSS.n1375 DVSS.n1369 0.0140606
R31167 DVSS.n1390 DVSS.n1370 0.0140606
R31168 DVSS.n1374 DVSS.n1371 0.0140606
R31169 DVSS.n1389 DVSS.n1372 0.0140606
R31170 DVSS.n1373 DVSS.n1372 0.0140606
R31171 DVSS.n8402 DVSS.n8401 0.0140606
R31172 DVSS.n2334 DVSS.n2311 0.0140606
R31173 DVSS.n2304 DVSS.n2281 0.0140606
R31174 DVSS.n3781 DVSS.n3776 0.0140606
R31175 DVSS.n3782 DVSS.n3770 0.0140606
R31176 DVSS.n4745 DVSS.n4619 0.0140606
R31177 DVSS.n4748 DVSS.n4747 0.0140606
R31178 DVSS.n9021 DVSS.n9020 0.0140606
R31179 DVSS.n9380 DVSS.n9379 0.0140606
R31180 DVSS.n9022 DVSS.n9019 0.0140606
R31181 DVSS.n388 DVSS.n385 0.0140606
R31182 DVSS.n9024 DVSS.n699 0.0140606
R31183 DVSS.n9382 DVSS.n387 0.0140606
R31184 DVSS.n8867 DVSS.n8866 0.0140606
R31185 DVSS.n376 DVSS.n373 0.0140606
R31186 DVSS.n8868 DVSS.n606 0.0140606
R31187 DVSS.n9391 DVSS.n9390 0.0140606
R31188 DVSS.n3235 DVSS.n3233 0.0140606
R31189 DVSS.n5405 DVSS.n5404 0.0140606
R31190 DVSS.n5693 DVSS.n5692 0.0140606
R31191 DVSS.n5493 DVSS.n5492 0.0140606
R31192 DVSS.n3237 DVSS.n3231 0.0140606
R31193 DVSS.n5695 DVSS.n3231 0.0140606
R31194 DVSS.n5490 DVSS.n5486 0.0140606
R31195 DVSS.n5490 DVSS.n5403 0.0140606
R31196 DVSS.n3279 DVSS.n3278 0.0140606
R31197 DVSS.n5548 DVSS.n3289 0.0140606
R31198 DVSS.n3280 DVSS.n3274 0.0140606
R31199 DVSS.n5635 DVSS.n5634 0.0140606
R31200 DVSS.n5644 DVSS.n3276 0.0140606
R31201 DVSS.n5644 DVSS.n5643 0.0140606
R31202 DVSS.n5632 DVSS.n3287 0.0140606
R31203 DVSS.n5637 DVSS.n3287 0.0140606
R31204 DVSS.n2698 DVSS.n2652 0.0140606
R31205 DVSS.n2708 DVSS.n2707 0.0140606
R31206 DVSS.n7269 DVSS.n7268 0.0140606
R31207 DVSS.n2750 DVSS.n2703 0.0140606
R31208 DVSS.n7267 DVSS.n7266 0.0140606
R31209 DVSS.n7266 DVSS.n2697 0.0140606
R31210 DVSS.n2753 DVSS.n2705 0.0140606
R31211 DVSS.n2753 DVSS.n2752 0.0140606
R31212 DVSS.n2619 DVSS.n2618 0.0140606
R31213 DVSS.n2082 DVSS.n2078 0.0140606
R31214 DVSS.n2620 DVSS.n2614 0.0140606
R31215 DVSS.n7859 DVSS.n7858 0.0140606
R31216 DVSS.n7332 DVSS.n2616 0.0140606
R31217 DVSS.n7332 DVSS.n7331 0.0140606
R31218 DVSS.n7857 DVSS.n7856 0.0140606
R31219 DVSS.n7856 DVSS.n2081 0.0140606
R31220 DVSS.n1878 DVSS.n1877 0.0140606
R31221 DVSS.n1867 DVSS.n1866 0.0140606
R31222 DVSS.n8092 DVSS.n8091 0.0140606
R31223 DVSS.n8104 DVSS.n8103 0.0140606
R31224 DVSS.n1880 DVSS.n1875 0.0140606
R31225 DVSS.n8094 DVSS.n1875 0.0140606
R31226 DVSS.n8101 DVSS.n1869 0.0140606
R31227 DVSS.n8101 DVSS.n1865 0.0140606
R31228 DVSS.n604 DVSS.n595 0.0140606
R31229 DVSS.n615 DVSS.n597 0.0140606
R31230 DVSS.n9113 DVSS.n593 0.0140606
R31231 DVSS.n9113 DVSS.n9112 0.0140606
R31232 DVSS.n9115 DVSS.n592 0.0140606
R31233 DVSS.n9115 DVSS.n9114 0.0140606
R31234 DVSS.n9117 DVSS.n591 0.0140606
R31235 DVSS.n9117 DVSS.n9116 0.0140606
R31236 DVSS.n9119 DVSS.n590 0.0140606
R31237 DVSS.n9119 DVSS.n9118 0.0140606
R31238 DVSS.n9120 DVSS.n588 0.0140606
R31239 DVSS.n611 DVSS.n599 0.0140606
R31240 DVSS.n9122 DVSS.n611 0.0140606
R31241 DVSS.n610 DVSS.n600 0.0140606
R31242 DVSS.n9124 DVSS.n610 0.0140606
R31243 DVSS.n609 DVSS.n601 0.0140606
R31244 DVSS.n9126 DVSS.n609 0.0140606
R31245 DVSS.n608 DVSS.n602 0.0140606
R31246 DVSS.n9150 DVSS.n567 0.0140606
R31247 DVSS.n9149 DVSS.n569 0.0140606
R31248 DVSS.n9139 DVSS.n565 0.0140606
R31249 DVSS.n9148 DVSS.n9139 0.0140606
R31250 DVSS.n9140 DVSS.n564 0.0140606
R31251 DVSS.n9147 DVSS.n9140 0.0140606
R31252 DVSS.n9141 DVSS.n563 0.0140606
R31253 DVSS.n9146 DVSS.n9141 0.0140606
R31254 DVSS.n9142 DVSS.n562 0.0140606
R31255 DVSS.n9145 DVSS.n9142 0.0140606
R31256 DVSS.n9151 DVSS.n560 0.0140606
R31257 DVSS.n578 DVSS.n571 0.0140606
R31258 DVSS.n9152 DVSS.n578 0.0140606
R31259 DVSS.n577 DVSS.n572 0.0140606
R31260 DVSS.n9154 DVSS.n577 0.0140606
R31261 DVSS.n576 DVSS.n573 0.0140606
R31262 DVSS.n576 DVSS.n574 0.0140606
R31263 DVSS.n9158 DVSS.n374 0.0140606
R31264 DVSS.n9050 DVSS.n648 0.0140606
R31265 DVSS.n9038 DVSS.n649 0.0140606
R31266 DVSS.n9051 DVSS.n9038 0.0140606
R31267 DVSS.n9037 DVSS.n650 0.0140606
R31268 DVSS.n9052 DVSS.n9037 0.0140606
R31269 DVSS.n9036 DVSS.n651 0.0140606
R31270 DVSS.n9053 DVSS.n9036 0.0140606
R31271 DVSS.n9035 DVSS.n652 0.0140606
R31272 DVSS.n9054 DVSS.n9035 0.0140606
R31273 DVSS.n9034 DVSS.n653 0.0140606
R31274 DVSS.n9055 DVSS.n9034 0.0140606
R31275 DVSS.n9033 DVSS.n654 0.0140606
R31276 DVSS.n9056 DVSS.n9033 0.0140606
R31277 DVSS.n9032 DVSS.n655 0.0140606
R31278 DVSS.n9057 DVSS.n9032 0.0140606
R31279 DVSS.n9031 DVSS.n656 0.0140606
R31280 DVSS.n9058 DVSS.n9031 0.0140606
R31281 DVSS.n9030 DVSS.n657 0.0140606
R31282 DVSS.n9059 DVSS.n9030 0.0140606
R31283 DVSS.n9029 DVSS.n658 0.0140606
R31284 DVSS.n9061 DVSS.n9029 0.0140606
R31285 DVSS.n9028 DVSS.n659 0.0140606
R31286 DVSS.n9028 DVSS.n660 0.0140606
R31287 DVSS.n9198 DVSS.n515 0.0140606
R31288 DVSS.n517 DVSS.n514 0.0140606
R31289 DVSS.n9199 DVSS.n514 0.0140606
R31290 DVSS.n519 DVSS.n513 0.0140606
R31291 DVSS.n9200 DVSS.n513 0.0140606
R31292 DVSS.n521 DVSS.n512 0.0140606
R31293 DVSS.n9201 DVSS.n512 0.0140606
R31294 DVSS.n523 DVSS.n511 0.0140606
R31295 DVSS.n9202 DVSS.n511 0.0140606
R31296 DVSS.n525 DVSS.n510 0.0140606
R31297 DVSS.n9203 DVSS.n510 0.0140606
R31298 DVSS.n527 DVSS.n509 0.0140606
R31299 DVSS.n9204 DVSS.n509 0.0140606
R31300 DVSS.n529 DVSS.n508 0.0140606
R31301 DVSS.n9205 DVSS.n508 0.0140606
R31302 DVSS.n531 DVSS.n507 0.0140606
R31303 DVSS.n9206 DVSS.n507 0.0140606
R31304 DVSS.n533 DVSS.n506 0.0140606
R31305 DVSS.n9207 DVSS.n506 0.0140606
R31306 DVSS.n535 DVSS.n505 0.0140606
R31307 DVSS.n9209 DVSS.n505 0.0140606
R31308 DVSS.n9210 DVSS.n504 0.0140606
R31309 DVSS.n504 DVSS.n501 0.0140606
R31310 DVSS.n9027 DVSS.n661 0.0140606
R31311 DVSS.n676 DVSS.n674 0.0140606
R31312 DVSS.n8778 DVSS.n674 0.0140606
R31313 DVSS.n678 DVSS.n673 0.0140606
R31314 DVSS.n8779 DVSS.n673 0.0140606
R31315 DVSS.n680 DVSS.n672 0.0140606
R31316 DVSS.n8780 DVSS.n672 0.0140606
R31317 DVSS.n682 DVSS.n671 0.0140606
R31318 DVSS.n8781 DVSS.n671 0.0140606
R31319 DVSS.n684 DVSS.n670 0.0140606
R31320 DVSS.n8782 DVSS.n670 0.0140606
R31321 DVSS.n686 DVSS.n669 0.0140606
R31322 DVSS.n8783 DVSS.n669 0.0140606
R31323 DVSS.n688 DVSS.n668 0.0140606
R31324 DVSS.n8784 DVSS.n668 0.0140606
R31325 DVSS.n690 DVSS.n667 0.0140606
R31326 DVSS.n8785 DVSS.n667 0.0140606
R31327 DVSS.n692 DVSS.n666 0.0140606
R31328 DVSS.n8786 DVSS.n666 0.0140606
R31329 DVSS.n694 DVSS.n665 0.0140606
R31330 DVSS.n8787 DVSS.n665 0.0140606
R31331 DVSS.n696 DVSS.n664 0.0140606
R31332 DVSS.n698 DVSS.n664 0.0140606
R31333 DVSS.n9215 DVSS.n9214 0.0140606
R31334 DVSS.n9218 DVSS.n9217 0.0140606
R31335 DVSS.n9219 DVSS.n9218 0.0140606
R31336 DVSS.n9222 DVSS.n9221 0.0140606
R31337 DVSS.n9223 DVSS.n9222 0.0140606
R31338 DVSS.n9226 DVSS.n9225 0.0140606
R31339 DVSS.n9227 DVSS.n9226 0.0140606
R31340 DVSS.n9230 DVSS.n9229 0.0140606
R31341 DVSS.n9231 DVSS.n9230 0.0140606
R31342 DVSS.n9234 DVSS.n9233 0.0140606
R31343 DVSS.n9235 DVSS.n9234 0.0140606
R31344 DVSS.n9238 DVSS.n9237 0.0140606
R31345 DVSS.n9239 DVSS.n9238 0.0140606
R31346 DVSS.n9242 DVSS.n9241 0.0140606
R31347 DVSS.n9243 DVSS.n9242 0.0140606
R31348 DVSS.n9246 DVSS.n9245 0.0140606
R31349 DVSS.n9247 DVSS.n9246 0.0140606
R31350 DVSS.n9250 DVSS.n9249 0.0140606
R31351 DVSS.n9251 DVSS.n9250 0.0140606
R31352 DVSS.n9254 DVSS.n9253 0.0140606
R31353 DVSS.n9255 DVSS.n9254 0.0140606
R31354 DVSS.n9258 DVSS.n9257 0.0140606
R31355 DVSS.n9259 DVSS.n9258 0.0140606
R31356 DVSS.n8245 DVSS.n8244 0.0138885
R31357 DVSS.n8251 DVSS.n8250 0.0138885
R31358 DVSS.n8260 DVSS.n8259 0.0138885
R31359 DVSS.n8277 DVSS.n8261 0.0138885
R31360 DVSS.n8265 DVSS.n8262 0.0138885
R31361 DVSS.n8278 DVSS.n8277 0.0138885
R31362 DVSS.n8278 DVSS.n8260 0.0138885
R31363 DVSS.n8273 DVSS.n8262 0.0138885
R31364 DVSS.n1488 DVSS.n1481 0.0138885
R31365 DVSS.n8290 DVSS.n1491 0.0138885
R31366 DVSS.n8284 DVSS.n1498 0.0138885
R31367 DVSS.n8324 DVSS.n8323 0.0138885
R31368 DVSS.n1501 DVSS.n1498 0.0138885
R31369 DVSS.n8323 DVSS.n1446 0.0138885
R31370 DVSS.n8234 DVSS.n8233 0.0138885
R31371 DVSS.n8231 DVSS.n1517 0.0138885
R31372 DVSS.n8303 DVSS.n8302 0.0138885
R31373 DVSS.n8310 DVSS.n8309 0.0138885
R31374 DVSS.n8304 DVSS.n8303 0.0138885
R31375 DVSS.n8309 DVSS.n8308 0.0138885
R31376 DVSS.n1494 DVSS.n1491 0.0138885
R31377 DVSS.n8252 DVSS.n8251 0.0138885
R31378 DVSS.n8228 DVSS.n1517 0.0138885
R31379 DVSS.n8293 DVSS.n1481 0.0138885
R31380 DVSS.n8244 DVSS.n8243 0.0138885
R31381 DVSS.n8233 DVSS.n1513 0.0138885
R31382 DVSS.n1186 DVSS.n1182 0.0138885
R31383 DVSS.n8446 DVSS.n8443 0.0138885
R31384 DVSS.n8445 DVSS.n1323 0.0138885
R31385 DVSS.n8441 DVSS.n1324 0.0138885
R31386 DVSS.n1386 DVSS.n1379 0.0138885
R31387 DVSS.n8473 DVSS.n8468 0.0138885
R31388 DVSS.n1138 DVSS.n1137 0.0138885
R31389 DVSS.n1131 DVSS.n1127 0.0138885
R31390 DVSS.n8443 DVSS.n1320 0.0138885
R31391 DVSS.n8441 DVSS.n1323 0.0138885
R31392 DVSS.n1386 DVSS.n1385 0.0138885
R31393 DVSS.n8473 DVSS.n8472 0.0138885
R31394 DVSS.n8476 DVSS.n1137 0.0138885
R31395 DVSS.n8482 DVSS.n1127 0.0138885
R31396 DVSS.n8446 DVSS.n8445 0.0138885
R31397 DVSS.n1222 DVSS.n1221 0.0138885
R31398 DVSS.n1224 DVSS.n1222 0.0138885
R31399 DVSS.n1229 DVSS.n1228 0.0138885
R31400 DVSS.n1231 DVSS.n1229 0.0138885
R31401 DVSS.n1280 DVSS.n1235 0.0138885
R31402 DVSS.n1271 DVSS.n1239 0.0138885
R31403 DVSS.n1244 DVSS.n1243 0.0138885
R31404 DVSS.n1246 DVSS.n1244 0.0138885
R31405 DVSS.n1251 DVSS.n1250 0.0138885
R31406 DVSS.n1253 DVSS.n1251 0.0138885
R31407 DVSS.n1285 DVSS.n1228 0.0138885
R31408 DVSS.n1236 DVSS.n1235 0.0138885
R31409 DVSS.n1240 DVSS.n1239 0.0138885
R31410 DVSS.n1265 DVSS.n1243 0.0138885
R31411 DVSS.n1260 DVSS.n1250 0.0138885
R31412 DVSS.n1258 DVSS.n1253 0.0138885
R31413 DVSS.n1263 DVSS.n1246 0.0138885
R31414 DVSS.n1283 DVSS.n1231 0.0138885
R31415 DVSS.n1159 DVSS.n1153 0.0138885
R31416 DVSS.n8455 DVSS.n1155 0.0138885
R31417 DVSS.n1157 DVSS.n1155 0.0138885
R31418 DVSS.n8369 DVSS.n8368 0.0138885
R31419 DVSS.n8365 DVSS.n8364 0.0138885
R31420 DVSS.n8364 DVSS.n8361 0.0138885
R31421 DVSS.n8374 DVSS.n8360 0.0138885
R31422 DVSS.n8378 DVSS.n8357 0.0138885
R31423 DVSS.n8383 DVSS.n8356 0.0138885
R31424 DVSS.n8381 DVSS.n8355 0.0138885
R31425 DVSS.n1423 DVSS.n1418 0.0138885
R31426 DVSS.n8351 DVSS.n1421 0.0138885
R31427 DVSS.n1421 DVSS.n1420 0.0138885
R31428 DVSS.n8493 DVSS.n8492 0.0138885
R31429 DVSS.n1102 DVSS.n1100 0.0138885
R31430 DVSS.n1100 DVSS.n1097 0.0138885
R31431 DVSS.n8370 DVSS.n8369 0.0138885
R31432 DVSS.n8366 DVSS.n8365 0.0138885
R31433 DVSS.n8375 DVSS.n8374 0.0138885
R31434 DVSS.n8384 DVSS.n8383 0.0138885
R31435 DVSS.n8354 DVSS.n1418 0.0138885
R31436 DVSS.n8352 DVSS.n8351 0.0138885
R31437 DVSS.n8494 DVSS.n8493 0.0138885
R31438 DVSS.n1103 DVSS.n1102 0.0138885
R31439 DVSS.n8496 DVSS.n1097 0.0138885
R31440 DVSS.n1420 DVSS.n1104 0.0138885
R31441 DVSS.n8381 DVSS.n8356 0.0138885
R31442 DVSS.n8360 DVSS.n8357 0.0138885
R31443 DVSS.n8372 DVSS.n8361 0.0138885
R31444 DVSS.n8458 DVSS.n1153 0.0138885
R31445 DVSS.n8456 DVSS.n8455 0.0138885
R31446 DVSS.n1158 DVSS.n1157 0.0138885
R31447 DVSS.n1318 DVSS.n1182 0.0138885
R31448 DVSS.n1290 DVSS.n1221 0.0138885
R31449 DVSS.n1288 DVSS.n1224 0.0138885
R31450 DVSS.n8247 DVSS.n8246 0.0138885
R31451 DVSS.n8253 DVSS.n8252 0.0138885
R31452 DVSS.n8261 DVSS.n1504 0.0138885
R31453 DVSS.n8267 DVSS.n8266 0.0138885
R31454 DVSS.n8274 DVSS.n1504 0.0138885
R31455 DVSS.n8269 DVSS.n8267 0.0138885
R31456 DVSS.n1489 DVSS.n1485 0.0138885
R31457 DVSS.n1495 DVSS.n1494 0.0138885
R31458 DVSS.n1502 DVSS.n1501 0.0138885
R31459 DVSS.n8325 DVSS.n1447 0.0138885
R31460 DVSS.n1503 DVSS.n1502 0.0138885
R31461 DVSS.n1448 DVSS.n1447 0.0138885
R31462 DVSS.n8235 DVSS.n1514 0.0138885
R31463 DVSS.n8228 DVSS.n8227 0.0138885
R31464 DVSS.n8305 DVSS.n8304 0.0138885
R31465 DVSS.n8312 DVSS.n8311 0.0138885
R31466 DVSS.n8305 DVSS.n1466 0.0138885
R31467 DVSS.n8312 DVSS.n1460 0.0138885
R31468 DVSS.n8227 DVSS.n8226 0.0138885
R31469 DVSS.n8253 DVSS.n1506 0.0138885
R31470 DVSS.n1496 DVSS.n1495 0.0138885
R31471 DVSS.n1515 DVSS.n1514 0.0138885
R31472 DVSS.n8247 DVSS.n1511 0.0138885
R31473 DVSS.n1486 DVSS.n1485 0.0138885
R31474 DVSS.n8449 DVSS.n1185 0.0138885
R31475 DVSS.n1381 DVSS.n1145 0.0138885
R31476 DVSS.n8475 DVSS.n1141 0.0138885
R31477 DVSS.n8480 DVSS.n1133 0.0138885
R31478 DVSS.n8486 DVSS.n1130 0.0138885
R31479 DVSS.n1130 DVSS.n1129 0.0138885
R31480 DVSS.n1139 DVSS.n1133 0.0138885
R31481 DVSS.n8469 DVSS.n1141 0.0138885
R31482 DVSS.n1381 DVSS.n1380 0.0138885
R31483 DVSS.n1286 DVSS.n1223 0.0138885
R31484 DVSS.n1281 DVSS.n1230 0.0138885
R31485 DVSS.n1278 DVSS.n1277 0.0138885
R31486 DVSS.n1269 DVSS.n1268 0.0138885
R31487 DVSS.n1261 DVSS.n1245 0.0138885
R31488 DVSS.n1256 DVSS.n1252 0.0138885
R31489 DVSS.n1254 DVSS.n1252 0.0138885
R31490 DVSS.n1247 DVSS.n1245 0.0138885
R31491 DVSS.n1269 DVSS.n1241 0.0138885
R31492 DVSS.n1278 DVSS.n1237 0.0138885
R31493 DVSS.n1232 DVSS.n1230 0.0138885
R31494 DVSS.n1185 DVSS.n1184 0.0138885
R31495 DVSS.n1225 DVSS.n1223 0.0138885
R31496 DVSS.n4659 DVSS.n3685 0.0138099
R31497 DVSS.n5561 DVSS.n2297 0.0138099
R31498 DVSS.n7873 DVSS.n2067 0.0138099
R31499 DVSS.n4660 DVSS.n3699 0.0138099
R31500 DVSS.n5605 DVSS.n2327 0.0138099
R31501 DVSS.n7874 DVSS.n2049 0.0138099
R31502 DVSS.n187 DVSS.n181 0.0137874
R31503 DVSS.n9716 DVSS.n185 0.0137874
R31504 DVSS.n226 DVSS.n220 0.0137874
R31505 DVSS.n9659 DVSS.n224 0.0137874
R31506 DVSS.n8873 DVSS.n799 0.0137874
R31507 DVSS.n805 DVSS.n801 0.0137874
R31508 DVSS.n8878 DVSS.n789 0.0137874
R31509 DVSS.n795 DVSS.n791 0.0137874
R31510 DVSS.n8905 DVSS.n775 0.0137874
R31511 DVSS.n9439 DVSS.n359 0.0137874
R31512 DVSS.n4830 DVSS.n3616 0.0134331
R31513 DVSS.n4838 DVSS.n3622 0.0134331
R31514 DVSS.n4832 DVSS.n3615 0.0134331
R31515 DVSS.n4887 DVSS.n3623 0.0134331
R31516 DVSS.n4846 DVSS.n3651 0.0134331
R31517 DVSS.n4844 DVSS.n3650 0.0134331
R31518 DVSS.n4843 DVSS.n3649 0.0134331
R31519 DVSS.n4827 DVSS.n3648 0.0134331
R31520 DVSS.n3714 DVSS.n3710 0.0134331
R31521 DVSS.n4802 DVSS.n3717 0.0134331
R31522 DVSS.n3718 DVSS.n3713 0.0134331
R31523 DVSS.n4798 DVSS.n4797 0.0134331
R31524 DVSS.n4193 DVSS.n3868 0.0134331
R31525 DVSS.n4436 DVSS.n4195 0.0134331
R31526 DVSS.n4198 DVSS.n4192 0.0134331
R31527 DVSS.n4431 DVSS.n4430 0.0134331
R31528 DVSS.n8934 DVSS.n759 0.0134331
R31529 DVSS.n8968 DVSS.n743 0.0134331
R31530 DVSS.n3862 DVSS.n3858 0.0134331
R31531 DVSS.n4439 DVSS.n3864 0.0134331
R31532 DVSS.n4216 DVSS.n3861 0.0134331
R31533 DVSS.n4259 DVSS.n4221 0.0134331
R31534 DVSS.n3595 DVSS.n3591 0.0134331
R31535 DVSS.n4977 DVSS.n3597 0.0134331
R31536 DVSS.n4973 DVSS.n3594 0.0134331
R31537 DVSS.n4974 DVSS.n3588 0.0134331
R31538 DVSS.n9468 DVSS.n344 0.0134331
R31539 DVSS.n9502 DVSS.n41 0.0134331
R31540 DVSS.n4931 DVSS.n4907 0.0134331
R31541 DVSS.n5917 DVSS.n2917 0.0134331
R31542 DVSS.n4445 DVSS.n3840 0.0134331
R31543 DVSS.n3021 DVSS.n3017 0.0134331
R31544 DVSS.n4659 DVSS.n3681 0.0133873
R31545 DVSS.n5561 DVSS.n2288 0.0133873
R31546 DVSS.n7873 DVSS.n2070 0.0133873
R31547 DVSS.n4660 DVSS.n3695 0.0133873
R31548 DVSS.n5605 DVSS.n2318 0.0133873
R31549 DVSS.n7874 DVSS.n2052 0.0133873
R31550 DVSS.n2905 DVSS.n2823 0.0130787
R31551 DVSS.n5067 DVSS.n3351 0.0130787
R31552 DVSS.n5384 DVSS.n3355 0.0130787
R31553 DVSS.n3357 DVSS.n3354 0.0130787
R31554 DVSS.n5072 DVSS.n5071 0.0130787
R31555 DVSS.n5066 DVSS.n3353 0.0130787
R31556 DVSS.n6005 DVSS.n6004 0.0130787
R31557 DVSS.n3347 DVSS.n3331 0.0130787
R31558 DVSS.n5388 DVSS.n3343 0.0130787
R31559 DVSS.n3344 DVSS.n3330 0.0130787
R31560 DVSS.n5392 DVSS.n5391 0.0130787
R31561 DVSS.n3329 DVSS.n3324 0.0130787
R31562 DVSS.n4598 DVSS.n3736 0.0130787
R31563 DVSS.n3524 DVSS.n3144 0.0130787
R31564 DVSS.n3554 DVSS.n3154 0.0130787
R31565 DVSS.n3526 DVSS.n3143 0.0130787
R31566 DVSS.n3550 DVSS.n3155 0.0130787
R31567 DVSS.n3156 DVSS.n3142 0.0130787
R31568 DVSS.n4581 DVSS.n3792 0.0130787
R31569 DVSS.n3529 DVSS.n3102 0.0130787
R31570 DVSS.n3546 DVSS.n3109 0.0130787
R31571 DVSS.n3531 DVSS.n3101 0.0130787
R31572 DVSS.n3542 DVSS.n3110 0.0130787
R31573 DVSS.n3111 DVSS.n3100 0.0130787
R31574 DVSS.n8889 DVSS.n768 0.0130787
R31575 DVSS.n8986 DVSS.n728 0.0130787
R31576 DVSS.n4471 DVSS.n3819 0.0130787
R31577 DVSS.n2909 DVSS.n2854 0.0130787
R31578 DVSS.n3375 DVSS.n3361 0.0130787
R31579 DVSS.n5381 DVSS.n3365 0.0130787
R31580 DVSS.n3367 DVSS.n3364 0.0130787
R31581 DVSS.n5368 DVSS.n3370 0.0130787
R31582 DVSS.n5367 DVSS.n3363 0.0130787
R31583 DVSS.n9423 DVSS.n353 0.0130787
R31584 DVSS.n9520 DVSS.n27 0.0130787
R31585 DVSS.n5924 DVSS.n2883 0.0130787
R31586 DVSS.n5372 DVSS.n2945 0.0130787
R31587 DVSS.n4475 DVSS.n4455 0.0130787
R31588 DVSS.n3013 DVSS.n2999 0.0130787
R31589 DVSS.n5553 DVSS.n2291 0.0129648
R31590 DVSS.n7900 DVSS.n7899 0.0129648
R31591 DVSS.n5621 DVSS.n2321 0.0129648
R31592 DVSS.n7897 DVSS.n2055 0.0129648
R31593 DVSS.n9007 DVSS.n9006 0.0128916
R31594 DVSS.n9013 DVSS.n9012 0.0128916
R31595 DVSS.n9378 DVSS.n389 0.0128916
R31596 DVSS.n329 DVSS.n325 0.0128916
R31597 DVSS.n9008 DVSS.n9007 0.0128916
R31598 DVSS.n9014 DVSS.n9013 0.0128916
R31599 DVSS.n9370 DVSS.n389 0.0128916
R31600 DVSS.n329 DVSS.n326 0.0128916
R31601 DVSS.n8879 DVSS.n787 0.0128916
R31602 DVSS.n793 DVSS.n792 0.0128916
R31603 DVSS.n793 DVSS.n790 0.0128916
R31604 DVSS.n8874 DVSS.n797 0.0128916
R31605 DVSS.n803 DVSS.n802 0.0128916
R31606 DVSS.n803 DVSS.n800 0.0128916
R31607 DVSS.n8869 DVSS.n8863 0.0128916
R31608 DVSS.n8865 DVSS.n8864 0.0128916
R31609 DVSS.n9393 DVSS.n9392 0.0128916
R31610 DVSS.n377 DVSS.n371 0.0128916
R31611 DVSS.n9398 DVSS.n9397 0.0128916
R31612 DVSS.n9402 DVSS.n9400 0.0128916
R31613 DVSS.n9403 DVSS.n9402 0.0128916
R31614 DVSS.n9407 DVSS.n9406 0.0128916
R31615 DVSS.n9411 DVSS.n9409 0.0128916
R31616 DVSS.n9412 DVSS.n9411 0.0128916
R31617 DVSS.n8877 DVSS.n787 0.0128916
R31618 DVSS.n8872 DVSS.n797 0.0128916
R31619 DVSS.n9399 DVSS.n9398 0.0128916
R31620 DVSS.n9408 DVSS.n9407 0.0128916
R31621 DVSS.n8877 DVSS.n792 0.0128916
R31622 DVSS.n8872 DVSS.n802 0.0128916
R31623 DVSS.n8864 DVSS.n378 0.0128916
R31624 DVSS.n9395 DVSS.n371 0.0128916
R31625 DVSS.n9400 DVSS.n9399 0.0128916
R31626 DVSS.n9409 DVSS.n9408 0.0128916
R31627 DVSS.n8875 DVSS.n790 0.0128916
R31628 DVSS.n8870 DVSS.n800 0.0128916
R31629 DVSS.n8865 DVSS.n8863 0.0128916
R31630 DVSS.n9393 DVSS.n377 0.0128916
R31631 DVSS.n9404 DVSS.n9403 0.0128916
R31632 DVSS.n9413 DVSS.n9412 0.0128916
R31633 DVSS.n5974 DVSS.n2831 0.0127244
R31634 DVSS.n2773 DVSS.n2768 0.0127244
R31635 DVSS.n4783 DVSS.n3744 0.0127244
R31636 DVSS.n4590 DVSS.n3796 0.0127244
R31637 DVSS.n8887 DVSS.n769 0.0127244
R31638 DVSS.n8984 DVSS.n729 0.0127244
R31639 DVSS.n4518 DVSS.n3826 0.0127244
R31640 DVSS.n5959 DVSS.n2864 0.0127244
R31641 DVSS.n9421 DVSS.n354 0.0127244
R31642 DVSS.n9518 DVSS.n28 0.0127244
R31643 DVSS.n5942 DVSS.n5928 0.0127244
R31644 DVSS.n5371 DVSS.n2944 0.0127244
R31645 DVSS.n4491 DVSS.n4478 0.0127244
R31646 DVSS.n5877 DVSS.n2998 0.0127244
R31647 DVSS.n4643 DVSS.n4641 0.01265
R31648 DVSS.n4678 DVSS.n4643 0.01265
R31649 DVSS.n4063 DVSS.n4023 0.01265
R31650 DVSS.n4066 DVSS.n4023 0.01265
R31651 DVSS.n5222 DVSS.n3500 0.01265
R31652 DVSS.n5219 DVSS.n3500 0.01265
R31653 DVSS.n5719 DVSS.n5718 0.01265
R31654 DVSS.n5718 DVSS.n5717 0.01265
R31655 DVSS.n5426 DVSS.n5424 0.01265
R31656 DVSS.n5461 DVSS.n5426 0.01265
R31657 DVSS.n5604 DVSS.n5602 0.01265
R31658 DVSS.n5602 DVSS.n5601 0.01265
R31659 DVSS.n7298 DVSS.n2639 0.01265
R31660 DVSS.n2639 DVSS.n2636 0.01265
R31661 DVSS.n7898 DVSS.n7896 0.01265
R31662 DVSS.n7896 DVSS.n2058 0.01265
R31663 DVSS.n7210 DVSS.n7169 0.01265
R31664 DVSS.n7213 DVSS.n7169 0.01265
R31665 DVSS.n3563 DVSS.n3481 0.0125423
R31666 DVSS.n5002 DVSS.n3479 0.0125423
R31667 DVSS.n3566 DVSS.n3482 0.0125423
R31668 DVSS.n3564 DVSS.n3478 0.0125423
R31669 DVSS.n5000 DVSS.n4999 0.0125423
R31670 DVSS.n5008 DVSS.n3518 0.0125423
R31671 DVSS.n5569 DVSS.n2300 0.0125423
R31672 DVSS.n4094 DVSS.n3977 0.0125423
R31673 DVSS.n4098 DVSS.n3975 0.0125423
R31674 DVSS.n4097 DVSS.n3978 0.0125423
R31675 DVSS.n4096 DVSS.n3974 0.0125423
R31676 DVSS.n4102 DVSS.n4101 0.0125423
R31677 DVSS.n5200 DVSS.n3179 0.0125423
R31678 DVSS.n5588 DVSS.n2330 0.0125423
R31679 DVSS.n9002 DVSS.n9000 0.0124231
R31680 DVSS.n9534 DVSS.n9533 0.0124231
R31681 DVSS.n8886 DVSS.n781 0.0124231
R31682 DVSS.n9420 DVSS.n9419 0.0124231
R31683 DVSS.n7245 DVSS.n7244 0.0123796
R31684 DVSS.n8219 DVSS.n1525 0.0123796
R31685 DVSS.n1469 DVSS.n1468 0.0123796
R31686 DVSS.n8306 DVSS.n1470 0.0123796
R31687 DVSS.n8276 DVSS.n8275 0.0123796
R31688 DVSS.n8276 DVSS.n1505 0.0123796
R31689 DVSS.n8282 DVSS.n1500 0.0123796
R31690 DVSS.n8283 DVSS.n1499 0.0123796
R31691 DVSS.n7097 DVSS.n7089 0.0123796
R31692 DVSS.n7102 DVSS.n7099 0.0123796
R31693 DVSS.n8386 DVSS.n1416 0.0123796
R31694 DVSS.n1144 DVSS.n1142 0.0123796
R31695 DVSS.n8471 DVSS.n8470 0.0123796
R31696 DVSS.n1266 DVSS.n1238 0.0123796
R31697 DVSS.n7095 DVSS.n7089 0.0123796
R31698 DVSS.n8275 DVSS.n1471 0.0123796
R31699 DVSS.n8279 DVSS.n1505 0.0123796
R31700 DVSS.n8283 DVSS.n8282 0.0123796
R31701 DVSS.n8280 DVSS.n1500 0.0123796
R31702 DVSS.n1470 DVSS.n1469 0.0123796
R31703 DVSS.n1468 DVSS.n1467 0.0123796
R31704 DVSS.n1528 DVSS.n1525 0.0123796
R31705 DVSS.n8223 DVSS.n1519 0.0123796
R31706 DVSS.n8229 DVSS.n8225 0.0123796
R31707 DVSS.n8230 DVSS.n1518 0.0123796
R31708 DVSS.n1509 DVSS.n1508 0.0123796
R31709 DVSS.n8254 DVSS.n1510 0.0123796
R31710 DVSS.n8288 DVSS.n1493 0.0123796
R31711 DVSS.n8289 DVSS.n1492 0.0123796
R31712 DVSS.n7110 DVSS.n7080 0.0123796
R31713 DVSS.n7107 DVSS.n7085 0.0123796
R31714 DVSS.n8377 DVSS.n8359 0.0123796
R31715 DVSS.n1383 DVSS.n1378 0.0123796
R31716 DVSS.n1384 DVSS.n1382 0.0123796
R31717 DVSS.n1275 DVSS.n1234 0.0123796
R31718 DVSS.n1523 DVSS.n1519 0.0123796
R31719 DVSS.n7083 DVSS.n7080 0.0123796
R31720 DVSS.n8289 DVSS.n8288 0.0123796
R31721 DVSS.n1497 DVSS.n1493 0.0123796
R31722 DVSS.n1510 DVSS.n1509 0.0123796
R31723 DVSS.n1508 DVSS.n1507 0.0123796
R31724 DVSS.n8230 DVSS.n8229 0.0123796
R31725 DVSS.n8225 DVSS.n8224 0.0123796
R31726 DVSS.n1387 DVSS.n1378 0.0123796
R31727 DVSS.n8474 DVSS.n1144 0.0123796
R31728 DVSS.n8471 DVSS.n1142 0.0123796
R31729 DVSS.n1384 DVSS.n1383 0.0123796
R31730 DVSS.n1276 DVSS.n1275 0.0123796
R31731 DVSS.n1267 DVSS.n1266 0.0123796
R31732 DVSS.n8382 DVSS.n1416 0.0123796
R31733 DVSS.n8373 DVSS.n8359 0.0123796
R31734 DVSS.n7109 DVSS.n7085 0.0123796
R31735 DVSS.n7099 DVSS.n7098 0.0123796
R31736 DVSS.n7246 DVSS.n7245 0.0123796
R31737 DVSS.n7249 DVSS.n7248 0.0123796
R31738 DVSS.n7249 DVSS.n6646 0.0123796
R31739 DVSS.n4993 DVSS.n3412 0.0123701
R31740 DVSS.n3582 DVSS.n3410 0.0123701
R31741 DVSS.n3586 DVSS.n3413 0.0123701
R31742 DVSS.n3581 DVSS.n3409 0.0123701
R31743 DVSS.n4997 DVSS.n3447 0.0123701
R31744 DVSS.n3572 DVSS.n3445 0.0123701
R31745 DVSS.n3576 DVSS.n3448 0.0123701
R31746 DVSS.n3571 DVSS.n3444 0.0123701
R31747 DVSS.n4009 DVSS.n3937 0.0123701
R31748 DVSS.n4002 DVSS.n3935 0.0123701
R31749 DVSS.n4005 DVSS.n3938 0.0123701
R31750 DVSS.n4001 DVSS.n3934 0.0123701
R31751 DVSS.n4188 DVSS.n3879 0.0123701
R31752 DVSS.n4187 DVSS.n3886 0.0123701
R31753 DVSS.n4175 DVSS.n4174 0.0123701
R31754 DVSS.n3894 DVSS.n3885 0.0123701
R31755 DVSS.n8935 DVSS.n754 0.0123701
R31756 DVSS.n8970 DVSS.n744 0.0123701
R31757 DVSS.n4990 DVSS.n3387 0.0123701
R31758 DVSS.n4983 DVSS.n3385 0.0123701
R31759 DVSS.n4987 DVSS.n3388 0.0123701
R31760 DVSS.n4982 DVSS.n3384 0.0123701
R31761 DVSS.n9469 DVSS.n339 0.0123701
R31762 DVSS.n9504 DVSS.n42 0.0123701
R31763 DVSS.n4929 DVSS.n4908 0.0123701
R31764 DVSS.n2930 DVSS.n2916 0.0123701
R31765 DVSS.n4444 DVSS.n3841 0.0123701
R31766 DVSS.n5866 DVSS.n3026 0.0123701
R31767 DVSS.n4703 DVSS.n4623 0.012331
R31768 DVSS.n4701 DVSS.n3777 0.012331
R31769 DVSS.n4621 DVSS.n4620 0.0121197
R31770 DVSS.n3985 DVSS.n3476 0.0121197
R31771 DVSS.n2700 DVSS.n2281 0.0121197
R31772 DVSS.n4606 DVSS.n3774 0.0121197
R31773 DVSS.n3980 DVSS.n3972 0.0121197
R31774 DVSS.n2699 DVSS.n2311 0.0121197
R31775 DVSS.n8903 DVSS.n774 0.0120157
R31776 DVSS.n9003 DVSS.n719 0.0120157
R31777 DVSS.n9437 DVSS.n358 0.0120157
R31778 DVSS.n9887 DVSS.n51 0.0120157
R31779 DVSS.n2832 DVSS.n2826 0.0119575
R31780 DVSS.n2836 DVSS.n2820 0.0119575
R31781 DVSS.n2828 DVSS.n2824 0.0119575
R31782 DVSS.n2835 DVSS.n2819 0.0119575
R31783 DVSS.n2829 DVSS.n2825 0.0119575
R31784 DVSS.n2834 DVSS.n2818 0.0119575
R31785 DVSS.n3631 DVSS.n3619 0.0119575
R31786 DVSS.n4883 DVSS.n4882 0.0119575
R31787 DVSS.n3630 DVSS.n3618 0.0119575
R31788 DVSS.n4885 DVSS.n4884 0.0119575
R31789 DVSS.n3629 DVSS.n3617 0.0119575
R31790 DVSS.n3628 DVSS.n3621 0.0119575
R31791 DVSS.n3414 DVSS.n3408 0.0119575
R31792 DVSS.n3418 DVSS.n3416 0.0119575
R31793 DVSS.n3417 DVSS.n3407 0.0119575
R31794 DVSS.n3421 DVSS.n3419 0.0119575
R31795 DVSS.n3420 DVSS.n3406 0.0119575
R31796 DVSS.n5306 DVSS.n3422 0.0119575
R31797 DVSS.n5081 DVSS.n5080 0.0119575
R31798 DVSS.n5078 DVSS.n5069 0.0119575
R31799 DVSS.n5079 DVSS.n5077 0.0119575
R31800 DVSS.n5075 DVSS.n5070 0.0119575
R31801 DVSS.n5076 DVSS.n5067 0.0119575
R31802 DVSS.n5506 DVSS.n3319 0.0119575
R31803 DVSS.n3320 DVSS.n3318 0.0119575
R31804 DVSS.n5502 DVSS.n3317 0.0119575
R31805 DVSS.n3316 DVSS.n3301 0.0119575
R31806 DVSS.n5536 DVSS.n3300 0.0119575
R31807 DVSS.n5533 DVSS.n5531 0.0119575
R31808 DVSS.n3304 DVSS.n3298 0.0119575
R31809 DVSS.n5530 DVSS.n5529 0.0119575
R31810 DVSS.n7601 DVSS.n7590 0.0119575
R31811 DVSS.n2222 DVSS.n2207 0.0119575
R31812 DVSS.n7602 DVSS.n7591 0.0119575
R31813 DVSS.n2221 DVSS.n2206 0.0119575
R31814 DVSS.n7603 DVSS.n7592 0.0119575
R31815 DVSS.n2220 DVSS.n2205 0.0119575
R31816 DVSS.n7604 DVSS.n7593 0.0119575
R31817 DVSS.n2219 DVSS.n2204 0.0119575
R31818 DVSS.n7605 DVSS.n7594 0.0119575
R31819 DVSS.n2218 DVSS.n2203 0.0119575
R31820 DVSS.n7606 DVSS.n7595 0.0119575
R31821 DVSS.n2217 DVSS.n2202 0.0119575
R31822 DVSS.n7607 DVSS.n7596 0.0119575
R31823 DVSS.n2216 DVSS.n2201 0.0119575
R31824 DVSS.n7608 DVSS.n7597 0.0119575
R31825 DVSS.n2215 DVSS.n2200 0.0119575
R31826 DVSS.n7609 DVSS.n7598 0.0119575
R31827 DVSS.n2214 DVSS.n2199 0.0119575
R31828 DVSS.n7610 DVSS.n7599 0.0119575
R31829 DVSS.n2213 DVSS.n2198 0.0119575
R31830 DVSS.n7613 DVSS.n7612 0.0119575
R31831 DVSS.n2212 DVSS.n2197 0.0119575
R31832 DVSS.n7615 DVSS.n2209 0.0119575
R31833 DVSS.n2742 DVSS.n2741 0.0119575
R31834 DVSS.n2739 DVSS.n2720 0.0119575
R31835 DVSS.n2725 DVSS.n2718 0.0119575
R31836 DVSS.n2724 DVSS.n2094 0.0119575
R31837 DVSS.n7724 DVSS.n2093 0.0119575
R31838 DVSS.n7721 DVSS.n7719 0.0119575
R31839 DVSS.n2098 DVSS.n2091 0.0119575
R31840 DVSS.n2097 DVSS.n1814 0.0119575
R31841 DVSS.n1821 DVSS.n1815 0.0119575
R31842 DVSS.n1823 DVSS.n1813 0.0119575
R31843 DVSS.n1830 DVSS.n1820 0.0119575
R31844 DVSS.n1824 DVSS.n1812 0.0119575
R31845 DVSS.n1829 DVSS.n1819 0.0119575
R31846 DVSS.n1825 DVSS.n1811 0.0119575
R31847 DVSS.n1828 DVSS.n1818 0.0119575
R31848 DVSS.n1826 DVSS.n1810 0.0119575
R31849 DVSS.n1827 DVSS.n1817 0.0119575
R31850 DVSS.n8120 DVSS.n1809 0.0119575
R31851 DVSS.n8117 DVSS.n1834 0.0119575
R31852 DVSS.n1853 DVSS.n1852 0.0119575
R31853 DVSS.n8113 DVSS.n1837 0.0119575
R31854 DVSS.n1836 DVSS.n1553 0.0119575
R31855 DVSS.n1115 DVSS.n1113 0.0119575
R31856 DVSS.n1119 DVSS.n1117 0.0119575
R31857 DVSS.n1118 DVSS.n1112 0.0119575
R31858 DVSS.n1121 DVSS.n1120 0.0119575
R31859 DVSS.n1111 DVSS.n1110 0.0119575
R31860 DVSS.n1124 DVSS.n1122 0.0119575
R31861 DVSS.n1123 DVSS.n1109 0.0119575
R31862 DVSS.n8488 DVSS.n1125 0.0119575
R31863 DVSS.n9692 DVSS.n178 0.0119575
R31864 DVSS.n182 DVSS.n175 0.0119575
R31865 DVSS.n9694 DVSS.n9693 0.0119575
R31866 DVSS.n9696 DVSS.n174 0.0119575
R31867 DVSS.n9697 DVSS.n9695 0.0119575
R31868 DVSS.n9699 DVSS.n173 0.0119575
R31869 DVSS.n9700 DVSS.n9698 0.0119575
R31870 DVSS.n9702 DVSS.n172 0.0119575
R31871 DVSS.n9703 DVSS.n9701 0.0119575
R31872 DVSS.n188 DVSS.n171 0.0119575
R31873 DVSS.n9705 DVSS.n9704 0.0119575
R31874 DVSS.n9707 DVSS.n169 0.0119575
R31875 DVSS.n9708 DVSS.n9706 0.0119575
R31876 DVSS.n9710 DVSS.n168 0.0119575
R31877 DVSS.n9711 DVSS.n9709 0.0119575
R31878 DVSS.n9713 DVSS.n167 0.0119575
R31879 DVSS.n9714 DVSS.n9712 0.0119575
R31880 DVSS.n187 DVSS.n166 0.0119575
R31881 DVSS.n9405 DVSS.n368 0.0119575
R31882 DVSS.n9410 DVSS.n367 0.0119575
R31883 DVSS.n273 DVSS.n272 0.0119575
R31884 DVSS.n9575 DVSS.n9558 0.0119575
R31885 DVSS.n9559 DVSS.n274 0.0119575
R31886 DVSS.n9574 DVSS.n9557 0.0119575
R31887 DVSS.n9560 DVSS.n275 0.0119575
R31888 DVSS.n9573 DVSS.n9556 0.0119575
R31889 DVSS.n9561 DVSS.n276 0.0119575
R31890 DVSS.n9572 DVSS.n9555 0.0119575
R31891 DVSS.n9562 DVSS.n277 0.0119575
R31892 DVSS.n9571 DVSS.n9554 0.0119575
R31893 DVSS.n9563 DVSS.n278 0.0119575
R31894 DVSS.n9570 DVSS.n9553 0.0119575
R31895 DVSS.n9564 DVSS.n279 0.0119575
R31896 DVSS.n9569 DVSS.n9552 0.0119575
R31897 DVSS.n9565 DVSS.n280 0.0119575
R31898 DVSS.n9568 DVSS.n9551 0.0119575
R31899 DVSS.n9566 DVSS.n281 0.0119575
R31900 DVSS.n9567 DVSS.n9550 0.0119575
R31901 DVSS.n9578 DVSS.n282 0.0119575
R31902 DVSS.n9577 DVSS.n9549 0.0119575
R31903 DVSS.n9579 DVSS.n283 0.0119575
R31904 DVSS.n9581 DVSS.n9547 0.0119575
R31905 DVSS.n9582 DVSS.n9546 0.0119575
R31906 DVSS.n302 DVSS.n284 0.0119575
R31907 DVSS.n301 DVSS.n299 0.0119575
R31908 DVSS.n9314 DVSS.n304 0.0119575
R31909 DVSS.n303 DVSS.n298 0.0119575
R31910 DVSS.n9315 DVSS.n306 0.0119575
R31911 DVSS.n305 DVSS.n297 0.0119575
R31912 DVSS.n9316 DVSS.n308 0.0119575
R31913 DVSS.n307 DVSS.n296 0.0119575
R31914 DVSS.n9317 DVSS.n310 0.0119575
R31915 DVSS.n309 DVSS.n295 0.0119575
R31916 DVSS.n9318 DVSS.n312 0.0119575
R31917 DVSS.n311 DVSS.n294 0.0119575
R31918 DVSS.n9319 DVSS.n314 0.0119575
R31919 DVSS.n313 DVSS.n293 0.0119575
R31920 DVSS.n9320 DVSS.n316 0.0119575
R31921 DVSS.n315 DVSS.n292 0.0119575
R31922 DVSS.n9321 DVSS.n318 0.0119575
R31923 DVSS.n317 DVSS.n291 0.0119575
R31924 DVSS.n9322 DVSS.n320 0.0119575
R31925 DVSS.n319 DVSS.n290 0.0119575
R31926 DVSS.n9323 DVSS.n322 0.0119575
R31927 DVSS.n321 DVSS.n289 0.0119575
R31928 DVSS.n9543 DVSS.n323 0.0119575
R31929 DVSS.n328 DVSS.n324 0.0119575
R31930 DVSS.n9540 DVSS.n9538 0.0119575
R31931 DVSS.n9539 DVSS.n330 0.0119575
R31932 DVSS.n3415 DVSS.n3414 0.0119575
R31933 DVSS.n3416 DVSS.n3408 0.0119575
R31934 DVSS.n3418 DVSS.n3417 0.0119575
R31935 DVSS.n3419 DVSS.n3407 0.0119575
R31936 DVSS.n3421 DVSS.n3420 0.0119575
R31937 DVSS.n3422 DVSS.n3406 0.0119575
R31938 DVSS.n5081 DVSS.n3423 0.0119575
R31939 DVSS.n5080 DVSS.n5069 0.0119575
R31940 DVSS.n5079 DVSS.n5078 0.0119575
R31941 DVSS.n5077 DVSS.n5070 0.0119575
R31942 DVSS.n5076 DVSS.n5075 0.0119575
R31943 DVSS.n8122 DVSS.n1815 0.0119575
R31944 DVSS.n1821 DVSS.n1813 0.0119575
R31945 DVSS.n1830 DVSS.n1823 0.0119575
R31946 DVSS.n1820 DVSS.n1812 0.0119575
R31947 DVSS.n1829 DVSS.n1824 0.0119575
R31948 DVSS.n1819 DVSS.n1811 0.0119575
R31949 DVSS.n1828 DVSS.n1825 0.0119575
R31950 DVSS.n1818 DVSS.n1810 0.0119575
R31951 DVSS.n1827 DVSS.n1826 0.0119575
R31952 DVSS.n1817 DVSS.n1809 0.0119575
R31953 DVSS.n1116 DVSS.n1115 0.0119575
R31954 DVSS.n1117 DVSS.n1113 0.0119575
R31955 DVSS.n1119 DVSS.n1118 0.0119575
R31956 DVSS.n1120 DVSS.n1112 0.0119575
R31957 DVSS.n1110 DVSS.n1101 0.0119575
R31958 DVSS.n1122 DVSS.n1111 0.0119575
R31959 DVSS.n1124 DVSS.n1123 0.0119575
R31960 DVSS.n1125 DVSS.n1109 0.0119575
R31961 DVSS.n3631 DVSS.n3620 0.0119575
R31962 DVSS.n4882 DVSS.n3619 0.0119575
R31963 DVSS.n4883 DVSS.n3618 0.0119575
R31964 DVSS.n4884 DVSS.n3630 0.0119575
R31965 DVSS.n4885 DVSS.n3617 0.0119575
R31966 DVSS.n3629 DVSS.n3628 0.0119575
R31967 DVSS.n2784 DVSS.n2770 0.0119575
R31968 DVSS.n2788 DVSS.n2780 0.0119575
R31969 DVSS.n2791 DVSS.n2790 0.0119575
R31970 DVSS.n2793 DVSS.n2787 0.0119575
R31971 DVSS.n6002 DVSS.n2792 0.0119575
R31972 DVSS.n6001 DVSS.n2786 0.0119575
R31973 DVSS.n3659 DVSS.n3655 0.0119575
R31974 DVSS.n3661 DVSS.n3654 0.0119575
R31975 DVSS.n3664 DVSS.n3658 0.0119575
R31976 DVSS.n3662 DVSS.n3653 0.0119575
R31977 DVSS.n3663 DVSS.n3657 0.0119575
R31978 DVSS.n4847 DVSS.n3652 0.0119575
R31979 DVSS.n3449 DVSS.n3443 0.0119575
R31980 DVSS.n3453 DVSS.n3451 0.0119575
R31981 DVSS.n3452 DVSS.n3442 0.0119575
R31982 DVSS.n3456 DVSS.n3454 0.0119575
R31983 DVSS.n3455 DVSS.n3441 0.0119575
R31984 DVSS.n5271 DVSS.n3457 0.0119575
R31985 DVSS.n3335 DVSS.n3334 0.0119575
R31986 DVSS.n3339 DVSS.n3336 0.0119575
R31987 DVSS.n3341 DVSS.n3340 0.0119575
R31988 DVSS.n3342 DVSS.n3338 0.0119575
R31989 DVSS.n3337 DVSS.n3331 0.0119575
R31990 DVSS.n5499 DVSS.n5399 0.0119575
R31991 DVSS.n5400 DVSS.n5398 0.0119575
R31992 DVSS.n5495 DVSS.n5397 0.0119575
R31993 DVSS.n5396 DVSS.n3293 0.0119575
R31994 DVSS.n5546 DVSS.n3292 0.0119575
R31995 DVSS.n5543 DVSS.n5541 0.0119575
R31996 DVSS.n3296 DVSS.n3290 0.0119575
R31997 DVSS.n5540 DVSS.n5539 0.0119575
R31998 DVSS.n7543 DVSS.n7532 0.0119575
R31999 DVSS.n2264 DVSS.n2249 0.0119575
R32000 DVSS.n7544 DVSS.n7533 0.0119575
R32001 DVSS.n2263 DVSS.n2248 0.0119575
R32002 DVSS.n7545 DVSS.n7534 0.0119575
R32003 DVSS.n2262 DVSS.n2247 0.0119575
R32004 DVSS.n7546 DVSS.n7535 0.0119575
R32005 DVSS.n2261 DVSS.n2246 0.0119575
R32006 DVSS.n7547 DVSS.n7536 0.0119575
R32007 DVSS.n2260 DVSS.n2245 0.0119575
R32008 DVSS.n7548 DVSS.n7537 0.0119575
R32009 DVSS.n2259 DVSS.n2244 0.0119575
R32010 DVSS.n7549 DVSS.n7538 0.0119575
R32011 DVSS.n2258 DVSS.n2243 0.0119575
R32012 DVSS.n7550 DVSS.n7539 0.0119575
R32013 DVSS.n2257 DVSS.n2242 0.0119575
R32014 DVSS.n7551 DVSS.n7540 0.0119575
R32015 DVSS.n2256 DVSS.n2241 0.0119575
R32016 DVSS.n7552 DVSS.n7541 0.0119575
R32017 DVSS.n2255 DVSS.n2240 0.0119575
R32018 DVSS.n7555 DVSS.n7554 0.0119575
R32019 DVSS.n2254 DVSS.n2239 0.0119575
R32020 DVSS.n7557 DVSS.n2251 0.0119575
R32021 DVSS.n2748 DVSS.n2747 0.0119575
R32022 DVSS.n2745 DVSS.n2711 0.0119575
R32023 DVSS.n2716 DVSS.n2709 0.0119575
R32024 DVSS.n2715 DVSS.n2086 0.0119575
R32025 DVSS.n7854 DVSS.n2085 0.0119575
R32026 DVSS.n7851 DVSS.n7849 0.0119575
R32027 DVSS.n2089 DVSS.n2083 0.0119575
R32028 DVSS.n7848 DVSS.n7727 0.0119575
R32029 DVSS.n7736 DVSS.n7728 0.0119575
R32030 DVSS.n7739 DVSS.n7738 0.0119575
R32031 DVSS.n7750 DVSS.n7735 0.0119575
R32032 DVSS.n7741 DVSS.n7740 0.0119575
R32033 DVSS.n7749 DVSS.n7734 0.0119575
R32034 DVSS.n7743 DVSS.n7742 0.0119575
R32035 DVSS.n7748 DVSS.n7733 0.0119575
R32036 DVSS.n7745 DVSS.n7744 0.0119575
R32037 DVSS.n7747 DVSS.n7732 0.0119575
R32038 DVSS.n7845 DVSS.n7746 0.0119575
R32039 DVSS.n8110 DVSS.n1861 0.0119575
R32040 DVSS.n1862 DVSS.n1860 0.0119575
R32041 DVSS.n8106 DVSS.n1857 0.0119575
R32042 DVSS.n1859 DVSS.n1858 0.0119575
R32043 DVSS.n8340 DVSS.n1435 0.0119575
R32044 DVSS.n8344 DVSS.n8342 0.0119575
R32045 DVSS.n8343 DVSS.n1434 0.0119575
R32046 DVSS.n1433 DVSS.n1424 0.0119575
R32047 DVSS.n1432 DVSS.n1431 0.0119575
R32048 DVSS.n8347 DVSS.n8345 0.0119575
R32049 DVSS.n8346 DVSS.n1430 0.0119575
R32050 DVSS.n1429 DVSS.n1135 0.0119575
R32051 DVSS.n9635 DVSS.n217 0.0119575
R32052 DVSS.n221 DVSS.n214 0.0119575
R32053 DVSS.n9637 DVSS.n9636 0.0119575
R32054 DVSS.n9639 DVSS.n213 0.0119575
R32055 DVSS.n9640 DVSS.n9638 0.0119575
R32056 DVSS.n9642 DVSS.n212 0.0119575
R32057 DVSS.n9643 DVSS.n9641 0.0119575
R32058 DVSS.n9645 DVSS.n211 0.0119575
R32059 DVSS.n9646 DVSS.n9644 0.0119575
R32060 DVSS.n227 DVSS.n210 0.0119575
R32061 DVSS.n9648 DVSS.n9647 0.0119575
R32062 DVSS.n9650 DVSS.n208 0.0119575
R32063 DVSS.n9651 DVSS.n9649 0.0119575
R32064 DVSS.n9653 DVSS.n207 0.0119575
R32065 DVSS.n9654 DVSS.n9652 0.0119575
R32066 DVSS.n9656 DVSS.n206 0.0119575
R32067 DVSS.n9657 DVSS.n9655 0.0119575
R32068 DVSS.n226 DVSS.n205 0.0119575
R32069 DVSS.n9396 DVSS.n370 0.0119575
R32070 DVSS.n9401 DVSS.n369 0.0119575
R32071 DVSS.n424 DVSS.n422 0.0119575
R32072 DVSS.n423 DVSS.n420 0.0119575
R32073 DVSS.n444 DVSS.n426 0.0119575
R32074 DVSS.n425 DVSS.n419 0.0119575
R32075 DVSS.n445 DVSS.n428 0.0119575
R32076 DVSS.n427 DVSS.n418 0.0119575
R32077 DVSS.n446 DVSS.n430 0.0119575
R32078 DVSS.n429 DVSS.n417 0.0119575
R32079 DVSS.n447 DVSS.n432 0.0119575
R32080 DVSS.n431 DVSS.n416 0.0119575
R32081 DVSS.n448 DVSS.n434 0.0119575
R32082 DVSS.n433 DVSS.n415 0.0119575
R32083 DVSS.n449 DVSS.n436 0.0119575
R32084 DVSS.n435 DVSS.n414 0.0119575
R32085 DVSS.n450 DVSS.n438 0.0119575
R32086 DVSS.n437 DVSS.n413 0.0119575
R32087 DVSS.n451 DVSS.n440 0.0119575
R32088 DVSS.n439 DVSS.n412 0.0119575
R32089 DVSS.n452 DVSS.n442 0.0119575
R32090 DVSS.n441 DVSS.n411 0.0119575
R32091 DVSS.n456 DVSS.n454 0.0119575
R32092 DVSS.n455 DVSS.n410 0.0119575
R32093 DVSS.n458 DVSS.n406 0.0119575
R32094 DVSS.n9353 DVSS.n462 0.0119575
R32095 DVSS.n461 DVSS.n405 0.0119575
R32096 DVSS.n9354 DVSS.n464 0.0119575
R32097 DVSS.n463 DVSS.n404 0.0119575
R32098 DVSS.n9355 DVSS.n466 0.0119575
R32099 DVSS.n465 DVSS.n403 0.0119575
R32100 DVSS.n9356 DVSS.n468 0.0119575
R32101 DVSS.n467 DVSS.n402 0.0119575
R32102 DVSS.n9357 DVSS.n470 0.0119575
R32103 DVSS.n469 DVSS.n401 0.0119575
R32104 DVSS.n9358 DVSS.n472 0.0119575
R32105 DVSS.n471 DVSS.n400 0.0119575
R32106 DVSS.n9359 DVSS.n474 0.0119575
R32107 DVSS.n473 DVSS.n399 0.0119575
R32108 DVSS.n9360 DVSS.n476 0.0119575
R32109 DVSS.n475 DVSS.n398 0.0119575
R32110 DVSS.n9361 DVSS.n478 0.0119575
R32111 DVSS.n477 DVSS.n397 0.0119575
R32112 DVSS.n9362 DVSS.n480 0.0119575
R32113 DVSS.n479 DVSS.n396 0.0119575
R32114 DVSS.n9366 DVSS.n9364 0.0119575
R32115 DVSS.n9365 DVSS.n395 0.0119575
R32116 DVSS.n9368 DVSS.n391 0.0119575
R32117 DVSS.n9372 DVSS.n9369 0.0119575
R32118 DVSS.n9375 DVSS.n390 0.0119575
R32119 DVSS.n9374 DVSS.n9373 0.0119575
R32120 DVSS.n4849 DVSS.n3655 0.0119575
R32121 DVSS.n3659 DVSS.n3654 0.0119575
R32122 DVSS.n3664 DVSS.n3661 0.0119575
R32123 DVSS.n3658 DVSS.n3653 0.0119575
R32124 DVSS.n3663 DVSS.n3662 0.0119575
R32125 DVSS.n3657 DVSS.n3652 0.0119575
R32126 DVSS.n3450 DVSS.n3449 0.0119575
R32127 DVSS.n3451 DVSS.n3443 0.0119575
R32128 DVSS.n3453 DVSS.n3452 0.0119575
R32129 DVSS.n3454 DVSS.n3442 0.0119575
R32130 DVSS.n3456 DVSS.n3455 0.0119575
R32131 DVSS.n3457 DVSS.n3441 0.0119575
R32132 DVSS.n3334 DVSS.n3333 0.0119575
R32133 DVSS.n3336 DVSS.n3335 0.0119575
R32134 DVSS.n3340 DVSS.n3339 0.0119575
R32135 DVSS.n3342 DVSS.n3341 0.0119575
R32136 DVSS.n3338 DVSS.n3337 0.0119575
R32137 DVSS.n7847 DVSS.n7728 0.0119575
R32138 DVSS.n7738 DVSS.n7736 0.0119575
R32139 DVSS.n7750 DVSS.n7739 0.0119575
R32140 DVSS.n7740 DVSS.n7735 0.0119575
R32141 DVSS.n7749 DVSS.n7741 0.0119575
R32142 DVSS.n7742 DVSS.n7734 0.0119575
R32143 DVSS.n7748 DVSS.n7743 0.0119575
R32144 DVSS.n7744 DVSS.n7733 0.0119575
R32145 DVSS.n7747 DVSS.n7745 0.0119575
R32146 DVSS.n7746 DVSS.n7732 0.0119575
R32147 DVSS.n8341 DVSS.n8340 0.0119575
R32148 DVSS.n8342 DVSS.n1435 0.0119575
R32149 DVSS.n8344 DVSS.n8343 0.0119575
R32150 DVSS.n1434 DVSS.n1433 0.0119575
R32151 DVSS.n1431 DVSS.n1422 0.0119575
R32152 DVSS.n8345 DVSS.n1432 0.0119575
R32153 DVSS.n8347 DVSS.n8346 0.0119575
R32154 DVSS.n1430 DVSS.n1429 0.0119575
R32155 DVSS.n3742 DVSS.n3741 0.0119575
R32156 DVSS.n3746 DVSS.n3733 0.0119575
R32157 DVSS.n3738 DVSS.n3737 0.0119575
R32158 DVSS.n3745 DVSS.n3732 0.0119575
R32159 DVSS.n3740 DVSS.n3739 0.0119575
R32160 DVSS.n4785 DVSS.n3727 0.0119575
R32161 DVSS.n4786 DVSS.n3725 0.0119575
R32162 DVSS.n4790 DVSS.n4788 0.0119575
R32163 DVSS.n4789 DVSS.n3724 0.0119575
R32164 DVSS.n4793 DVSS.n4791 0.0119575
R32165 DVSS.n4792 DVSS.n3723 0.0119575
R32166 DVSS.n4795 DVSS.n4794 0.0119575
R32167 DVSS.n3945 DVSS.n3933 0.0119575
R32168 DVSS.n3948 DVSS.n3940 0.0119575
R32169 DVSS.n3944 DVSS.n3932 0.0119575
R32170 DVSS.n3949 DVSS.n3941 0.0119575
R32171 DVSS.n3943 DVSS.n3931 0.0119575
R32172 DVSS.n4138 DVSS.n3942 0.0119575
R32173 DVSS.n3148 DVSS.n3146 0.0119575
R32174 DVSS.n5773 DVSS.n3151 0.0119575
R32175 DVSS.n3150 DVSS.n3145 0.0119575
R32176 DVSS.n5774 DVSS.n3153 0.0119575
R32177 DVSS.n3152 DVSS.n3144 0.0119575
R32178 DVSS.n5689 DVSS.n3243 0.0119575
R32179 DVSS.n3244 DVSS.n3242 0.0119575
R32180 DVSS.n5685 DVSS.n3239 0.0119575
R32181 DVSS.n3241 DVSS.n3240 0.0119575
R32182 DVSS.n5653 DVSS.n3269 0.0119575
R32183 DVSS.n5650 DVSS.n5648 0.0119575
R32184 DVSS.n3272 DVSS.n3267 0.0119575
R32185 DVSS.n5647 DVSS.n5646 0.0119575
R32186 DVSS.n2368 DVSS.n2366 0.0119575
R32187 DVSS.n2367 DVSS.n2363 0.0119575
R32188 DVSS.n2371 DVSS.n2369 0.0119575
R32189 DVSS.n2370 DVSS.n2362 0.0119575
R32190 DVSS.n2374 DVSS.n2372 0.0119575
R32191 DVSS.n2373 DVSS.n2361 0.0119575
R32192 DVSS.n2377 DVSS.n2375 0.0119575
R32193 DVSS.n2376 DVSS.n2360 0.0119575
R32194 DVSS.n2380 DVSS.n2378 0.0119575
R32195 DVSS.n2379 DVSS.n2359 0.0119575
R32196 DVSS.n2383 DVSS.n2381 0.0119575
R32197 DVSS.n2382 DVSS.n2358 0.0119575
R32198 DVSS.n2386 DVSS.n2384 0.0119575
R32199 DVSS.n2385 DVSS.n2357 0.0119575
R32200 DVSS.n2389 DVSS.n2387 0.0119575
R32201 DVSS.n2388 DVSS.n2356 0.0119575
R32202 DVSS.n2392 DVSS.n2390 0.0119575
R32203 DVSS.n2391 DVSS.n2355 0.0119575
R32204 DVSS.n2395 DVSS.n2393 0.0119575
R32205 DVSS.n2394 DVSS.n2354 0.0119575
R32206 DVSS.n2398 DVSS.n2396 0.0119575
R32207 DVSS.n2397 DVSS.n2353 0.0119575
R32208 DVSS.n7453 DVSS.n2399 0.0119575
R32209 DVSS.n2692 DVSS.n2657 0.0119575
R32210 DVSS.n2658 DVSS.n2656 0.0119575
R32211 DVSS.n2688 DVSS.n2655 0.0119575
R32212 DVSS.n2654 DVSS.n2609 0.0119575
R32213 DVSS.n7341 DVSS.n2608 0.0119575
R32214 DVSS.n7338 DVSS.n7336 0.0119575
R32215 DVSS.n2612 DVSS.n2606 0.0119575
R32216 DVSS.n7335 DVSS.n7334 0.0119575
R32217 DVSS.n2017 DVSS.n2015 0.0119575
R32218 DVSS.n7968 DVSS.n2020 0.0119575
R32219 DVSS.n2019 DVSS.n2014 0.0119575
R32220 DVSS.n7969 DVSS.n2022 0.0119575
R32221 DVSS.n2021 DVSS.n2013 0.0119575
R32222 DVSS.n7970 DVSS.n2024 0.0119575
R32223 DVSS.n2023 DVSS.n2012 0.0119575
R32224 DVSS.n7971 DVSS.n2026 0.0119575
R32225 DVSS.n2025 DVSS.n2011 0.0119575
R32226 DVSS.n7974 DVSS.n7973 0.0119575
R32227 DVSS.n8088 DVSS.n1887 0.0119575
R32228 DVSS.n1888 DVSS.n1886 0.0119575
R32229 DVSS.n8084 DVSS.n1883 0.0119575
R32230 DVSS.n1885 DVSS.n1884 0.0119575
R32231 DVSS.n1343 DVSS.n1333 0.0119575
R32232 DVSS.n1337 DVSS.n1336 0.0119575
R32233 DVSS.n1342 DVSS.n1332 0.0119575
R32234 DVSS.n1339 DVSS.n1338 0.0119575
R32235 DVSS.n1340 DVSS.n1330 0.0119575
R32236 DVSS.n8438 DVSS.n8436 0.0119575
R32237 DVSS.n8437 DVSS.n1329 0.0119575
R32238 DVSS.n8440 DVSS.n1325 0.0119575
R32239 DVSS.n1077 DVSS.n1074 0.0119575
R32240 DVSS.n8533 DVSS.n1071 0.0119575
R32241 DVSS.n8544 DVSS.n8543 0.0119575
R32242 DVSS.n8541 DVSS.n1070 0.0119575
R32243 DVSS.n8546 DVSS.n8545 0.0119575
R32244 DVSS.n8540 DVSS.n1069 0.0119575
R32245 DVSS.n8548 DVSS.n8547 0.0119575
R32246 DVSS.n8539 DVSS.n1068 0.0119575
R32247 DVSS.n8550 DVSS.n8549 0.0119575
R32248 DVSS.n8538 DVSS.n1067 0.0119575
R32249 DVSS.n8552 DVSS.n8551 0.0119575
R32250 DVSS.n8537 DVSS.n1065 0.0119575
R32251 DVSS.n8554 DVSS.n8553 0.0119575
R32252 DVSS.n8536 DVSS.n1064 0.0119575
R32253 DVSS.n8556 DVSS.n8555 0.0119575
R32254 DVSS.n8535 DVSS.n1063 0.0119575
R32255 DVSS.n8558 DVSS.n8557 0.0119575
R32256 DVSS.n1062 DVSS.n799 0.0119575
R32257 DVSS.n8871 DVSS.n798 0.0119575
R32258 DVSS.n8861 DVSS.n804 0.0119575
R32259 DVSS.n811 DVSS.n806 0.0119575
R32260 DVSS.n8836 DVSS.n8835 0.0119575
R32261 DVSS.n8838 DVSS.n812 0.0119575
R32262 DVSS.n8837 DVSS.n8834 0.0119575
R32263 DVSS.n8840 DVSS.n813 0.0119575
R32264 DVSS.n8839 DVSS.n8833 0.0119575
R32265 DVSS.n8842 DVSS.n814 0.0119575
R32266 DVSS.n8841 DVSS.n8832 0.0119575
R32267 DVSS.n8844 DVSS.n815 0.0119575
R32268 DVSS.n8843 DVSS.n8831 0.0119575
R32269 DVSS.n8846 DVSS.n816 0.0119575
R32270 DVSS.n8845 DVSS.n8830 0.0119575
R32271 DVSS.n8848 DVSS.n817 0.0119575
R32272 DVSS.n8847 DVSS.n8829 0.0119575
R32273 DVSS.n8850 DVSS.n818 0.0119575
R32274 DVSS.n8849 DVSS.n8828 0.0119575
R32275 DVSS.n8852 DVSS.n819 0.0119575
R32276 DVSS.n8851 DVSS.n8827 0.0119575
R32277 DVSS.n8854 DVSS.n820 0.0119575
R32278 DVSS.n8853 DVSS.n8826 0.0119575
R32279 DVSS.n8855 DVSS.n821 0.0119575
R32280 DVSS.n8857 DVSS.n823 0.0119575
R32281 DVSS.n8858 DVSS.n822 0.0119575
R32282 DVSS.n856 DVSS.n854 0.0119575
R32283 DVSS.n855 DVSS.n851 0.0119575
R32284 DVSS.n859 DVSS.n857 0.0119575
R32285 DVSS.n858 DVSS.n850 0.0119575
R32286 DVSS.n862 DVSS.n860 0.0119575
R32287 DVSS.n861 DVSS.n849 0.0119575
R32288 DVSS.n865 DVSS.n863 0.0119575
R32289 DVSS.n864 DVSS.n848 0.0119575
R32290 DVSS.n868 DVSS.n866 0.0119575
R32291 DVSS.n867 DVSS.n847 0.0119575
R32292 DVSS.n871 DVSS.n869 0.0119575
R32293 DVSS.n870 DVSS.n846 0.0119575
R32294 DVSS.n874 DVSS.n872 0.0119575
R32295 DVSS.n873 DVSS.n845 0.0119575
R32296 DVSS.n877 DVSS.n875 0.0119575
R32297 DVSS.n876 DVSS.n844 0.0119575
R32298 DVSS.n880 DVSS.n878 0.0119575
R32299 DVSS.n879 DVSS.n843 0.0119575
R32300 DVSS.n883 DVSS.n881 0.0119575
R32301 DVSS.n882 DVSS.n842 0.0119575
R32302 DVSS.n8751 DVSS.n884 0.0119575
R32303 DVSS.n885 DVSS.n841 0.0119575
R32304 DVSS.n840 DVSS.n705 0.0119575
R32305 DVSS.n706 DVSS.n701 0.0119575
R32306 DVSS.n9011 DVSS.n704 0.0119575
R32307 DVSS.n703 DVSS.n702 0.0119575
R32308 DVSS.n4787 DVSS.n4786 0.0119575
R32309 DVSS.n4788 DVSS.n3725 0.0119575
R32310 DVSS.n4790 DVSS.n4789 0.0119575
R32311 DVSS.n4791 DVSS.n3724 0.0119575
R32312 DVSS.n4793 DVSS.n4792 0.0119575
R32313 DVSS.n4794 DVSS.n3723 0.0119575
R32314 DVSS.n3945 DVSS.n3939 0.0119575
R32315 DVSS.n3948 DVSS.n3933 0.0119575
R32316 DVSS.n3944 DVSS.n3940 0.0119575
R32317 DVSS.n3949 DVSS.n3932 0.0119575
R32318 DVSS.n3943 DVSS.n3941 0.0119575
R32319 DVSS.n3942 DVSS.n3931 0.0119575
R32320 DVSS.n3149 DVSS.n3148 0.0119575
R32321 DVSS.n5773 DVSS.n3146 0.0119575
R32322 DVSS.n3151 DVSS.n3150 0.0119575
R32323 DVSS.n5774 DVSS.n3145 0.0119575
R32324 DVSS.n3153 DVSS.n3152 0.0119575
R32325 DVSS.n2018 DVSS.n2017 0.0119575
R32326 DVSS.n7968 DVSS.n2015 0.0119575
R32327 DVSS.n2020 DVSS.n2019 0.0119575
R32328 DVSS.n7969 DVSS.n2014 0.0119575
R32329 DVSS.n2022 DVSS.n2021 0.0119575
R32330 DVSS.n7970 DVSS.n2013 0.0119575
R32331 DVSS.n2024 DVSS.n2023 0.0119575
R32332 DVSS.n7971 DVSS.n2012 0.0119575
R32333 DVSS.n2026 DVSS.n2025 0.0119575
R32334 DVSS.n7973 DVSS.n2011 0.0119575
R32335 DVSS.n1343 DVSS.n1335 0.0119575
R32336 DVSS.n1336 DVSS.n1333 0.0119575
R32337 DVSS.n1342 DVSS.n1337 0.0119575
R32338 DVSS.n1338 DVSS.n1332 0.0119575
R32339 DVSS.n1341 DVSS.n1340 0.0119575
R32340 DVSS.n8436 DVSS.n1330 0.0119575
R32341 DVSS.n8438 DVSS.n8437 0.0119575
R32342 DVSS.n1329 DVSS.n1325 0.0119575
R32343 DVSS.n3803 DVSS.n3793 0.0119575
R32344 DVSS.n4580 DVSS.n3807 0.0119575
R32345 DVSS.n4584 DVSS.n4582 0.0119575
R32346 DVSS.n4583 DVSS.n3806 0.0119575
R32347 DVSS.n4587 DVSS.n4585 0.0119575
R32348 DVSS.n4586 DVSS.n3805 0.0119575
R32349 DVSS.n4419 DVSS.n4205 0.0119575
R32350 DVSS.n4423 DVSS.n4421 0.0119575
R32351 DVSS.n4422 DVSS.n4204 0.0119575
R32352 DVSS.n4426 DVSS.n4424 0.0119575
R32353 DVSS.n4425 DVSS.n4203 0.0119575
R32354 DVSS.n4428 DVSS.n4427 0.0119575
R32355 DVSS.n4176 DVSS.n3893 0.0119575
R32356 DVSS.n4180 DVSS.n4178 0.0119575
R32357 DVSS.n4179 DVSS.n3892 0.0119575
R32358 DVSS.n4183 DVSS.n4181 0.0119575
R32359 DVSS.n4182 DVSS.n3891 0.0119575
R32360 DVSS.n4185 DVSS.n4184 0.0119575
R32361 DVSS.n3116 DVSS.n3104 0.0119575
R32362 DVSS.n5809 DVSS.n3107 0.0119575
R32363 DVSS.n3115 DVSS.n3103 0.0119575
R32364 DVSS.n5810 DVSS.n3108 0.0119575
R32365 DVSS.n3114 DVSS.n3102 0.0119575
R32366 DVSS.n5682 DVSS.n3252 0.0119575
R32367 DVSS.n3253 DVSS.n3251 0.0119575
R32368 DVSS.n5678 DVSS.n3248 0.0119575
R32369 DVSS.n3250 DVSS.n3249 0.0119575
R32370 DVSS.n5663 DVSS.n3262 0.0119575
R32371 DVSS.n5660 DVSS.n5658 0.0119575
R32372 DVSS.n3265 DVSS.n3260 0.0119575
R32373 DVSS.n5657 DVSS.n5656 0.0119575
R32374 DVSS.n7416 DVSS.n2432 0.0119575
R32375 DVSS.n2431 DVSS.n2428 0.0119575
R32376 DVSS.n2435 DVSS.n2433 0.0119575
R32377 DVSS.n2434 DVSS.n2427 0.0119575
R32378 DVSS.n2438 DVSS.n2436 0.0119575
R32379 DVSS.n2437 DVSS.n2426 0.0119575
R32380 DVSS.n2441 DVSS.n2439 0.0119575
R32381 DVSS.n2440 DVSS.n2425 0.0119575
R32382 DVSS.n2444 DVSS.n2442 0.0119575
R32383 DVSS.n2443 DVSS.n2424 0.0119575
R32384 DVSS.n2447 DVSS.n2445 0.0119575
R32385 DVSS.n2446 DVSS.n2423 0.0119575
R32386 DVSS.n2450 DVSS.n2448 0.0119575
R32387 DVSS.n2449 DVSS.n2422 0.0119575
R32388 DVSS.n2453 DVSS.n2451 0.0119575
R32389 DVSS.n2452 DVSS.n2421 0.0119575
R32390 DVSS.n2456 DVSS.n2454 0.0119575
R32391 DVSS.n2455 DVSS.n2420 0.0119575
R32392 DVSS.n2459 DVSS.n2457 0.0119575
R32393 DVSS.n2458 DVSS.n2419 0.0119575
R32394 DVSS.n2462 DVSS.n2460 0.0119575
R32395 DVSS.n2461 DVSS.n2418 0.0119575
R32396 DVSS.n7418 DVSS.n2463 0.0119575
R32397 DVSS.n2685 DVSS.n2665 0.0119575
R32398 DVSS.n2666 DVSS.n2664 0.0119575
R32399 DVSS.n2681 DVSS.n2663 0.0119575
R32400 DVSS.n2662 DVSS.n2601 0.0119575
R32401 DVSS.n7351 DVSS.n2600 0.0119575
R32402 DVSS.n7348 DVSS.n7346 0.0119575
R32403 DVSS.n2604 DVSS.n2598 0.0119575
R32404 DVSS.n7345 DVSS.n7344 0.0119575
R32405 DVSS.n1983 DVSS.n1981 0.0119575
R32406 DVSS.n8007 DVSS.n1986 0.0119575
R32407 DVSS.n1985 DVSS.n1980 0.0119575
R32408 DVSS.n8008 DVSS.n1988 0.0119575
R32409 DVSS.n1987 DVSS.n1979 0.0119575
R32410 DVSS.n8009 DVSS.n1990 0.0119575
R32411 DVSS.n1989 DVSS.n1978 0.0119575
R32412 DVSS.n8010 DVSS.n1992 0.0119575
R32413 DVSS.n1991 DVSS.n1977 0.0119575
R32414 DVSS.n8013 DVSS.n8012 0.0119575
R32415 DVSS.n8081 DVSS.n1897 0.0119575
R32416 DVSS.n1898 DVSS.n1896 0.0119575
R32417 DVSS.n8077 DVSS.n1893 0.0119575
R32418 DVSS.n1895 DVSS.n1894 0.0119575
R32419 DVSS.n1172 DVSS.n1170 0.0119575
R32420 DVSS.n1176 DVSS.n1174 0.0119575
R32421 DVSS.n1175 DVSS.n1169 0.0119575
R32422 DVSS.n1168 DVSS.n1160 0.0119575
R32423 DVSS.n1167 DVSS.n1166 0.0119575
R32424 DVSS.n1179 DVSS.n1177 0.0119575
R32425 DVSS.n1178 DVSS.n1165 0.0119575
R32426 DVSS.n8451 DVSS.n1180 0.0119575
R32427 DVSS.n1203 DVSS.n1189 0.0119575
R32428 DVSS.n1204 DVSS.n1200 0.0119575
R32429 DVSS.n1304 DVSS.n1207 0.0119575
R32430 DVSS.n1206 DVSS.n1199 0.0119575
R32431 DVSS.n1305 DVSS.n1209 0.0119575
R32432 DVSS.n1208 DVSS.n1198 0.0119575
R32433 DVSS.n1306 DVSS.n1211 0.0119575
R32434 DVSS.n1210 DVSS.n1197 0.0119575
R32435 DVSS.n1307 DVSS.n1213 0.0119575
R32436 DVSS.n1212 DVSS.n1196 0.0119575
R32437 DVSS.n1308 DVSS.n1299 0.0119575
R32438 DVSS.n1298 DVSS.n1194 0.0119575
R32439 DVSS.n1309 DVSS.n1301 0.0119575
R32440 DVSS.n1300 DVSS.n1193 0.0119575
R32441 DVSS.n1310 DVSS.n1303 0.0119575
R32442 DVSS.n1302 DVSS.n1192 0.0119575
R32443 DVSS.n1314 DVSS.n1312 0.0119575
R32444 DVSS.n1313 DVSS.n789 0.0119575
R32445 DVSS.n8876 DVSS.n788 0.0119575
R32446 DVSS.n796 DVSS.n794 0.0119575
R32447 DVSS.n7027 DVSS.n6944 0.0119575
R32448 DVSS.n6966 DVSS.n6941 0.0119575
R32449 DVSS.n6969 DVSS.n6945 0.0119575
R32450 DVSS.n6965 DVSS.n6940 0.0119575
R32451 DVSS.n6970 DVSS.n6946 0.0119575
R32452 DVSS.n6964 DVSS.n6939 0.0119575
R32453 DVSS.n6971 DVSS.n6947 0.0119575
R32454 DVSS.n6963 DVSS.n6938 0.0119575
R32455 DVSS.n6972 DVSS.n6948 0.0119575
R32456 DVSS.n6962 DVSS.n6937 0.0119575
R32457 DVSS.n6973 DVSS.n6949 0.0119575
R32458 DVSS.n6961 DVSS.n6936 0.0119575
R32459 DVSS.n6974 DVSS.n6950 0.0119575
R32460 DVSS.n6960 DVSS.n6935 0.0119575
R32461 DVSS.n6975 DVSS.n6951 0.0119575
R32462 DVSS.n6959 DVSS.n6934 0.0119575
R32463 DVSS.n6976 DVSS.n6952 0.0119575
R32464 DVSS.n6958 DVSS.n6933 0.0119575
R32465 DVSS.n6977 DVSS.n6953 0.0119575
R32466 DVSS.n6957 DVSS.n6932 0.0119575
R32467 DVSS.n6978 DVSS.n6954 0.0119575
R32468 DVSS.n6956 DVSS.n6931 0.0119575
R32469 DVSS.n7029 DVSS.n6955 0.0119575
R32470 DVSS.n919 DVSS.n917 0.0119575
R32471 DVSS.n918 DVSS.n914 0.0119575
R32472 DVSS.n922 DVSS.n920 0.0119575
R32473 DVSS.n921 DVSS.n913 0.0119575
R32474 DVSS.n925 DVSS.n923 0.0119575
R32475 DVSS.n924 DVSS.n912 0.0119575
R32476 DVSS.n928 DVSS.n926 0.0119575
R32477 DVSS.n927 DVSS.n911 0.0119575
R32478 DVSS.n931 DVSS.n929 0.0119575
R32479 DVSS.n930 DVSS.n910 0.0119575
R32480 DVSS.n934 DVSS.n932 0.0119575
R32481 DVSS.n933 DVSS.n909 0.0119575
R32482 DVSS.n937 DVSS.n935 0.0119575
R32483 DVSS.n936 DVSS.n908 0.0119575
R32484 DVSS.n940 DVSS.n938 0.0119575
R32485 DVSS.n939 DVSS.n907 0.0119575
R32486 DVSS.n943 DVSS.n941 0.0119575
R32487 DVSS.n942 DVSS.n906 0.0119575
R32488 DVSS.n946 DVSS.n944 0.0119575
R32489 DVSS.n945 DVSS.n905 0.0119575
R32490 DVSS.n8716 DVSS.n947 0.0119575
R32491 DVSS.n948 DVSS.n904 0.0119575
R32492 DVSS.n903 DVSS.n712 0.0119575
R32493 DVSS.n713 DVSS.n708 0.0119575
R32494 DVSS.n9005 DVSS.n711 0.0119575
R32495 DVSS.n710 DVSS.n709 0.0119575
R32496 DVSS.n4420 DVSS.n4419 0.0119575
R32497 DVSS.n4421 DVSS.n4205 0.0119575
R32498 DVSS.n4423 DVSS.n4422 0.0119575
R32499 DVSS.n4424 DVSS.n4204 0.0119575
R32500 DVSS.n4426 DVSS.n4425 0.0119575
R32501 DVSS.n4427 DVSS.n4203 0.0119575
R32502 DVSS.n4177 DVSS.n4176 0.0119575
R32503 DVSS.n4178 DVSS.n3893 0.0119575
R32504 DVSS.n4180 DVSS.n4179 0.0119575
R32505 DVSS.n4181 DVSS.n3892 0.0119575
R32506 DVSS.n4183 DVSS.n4182 0.0119575
R32507 DVSS.n4184 DVSS.n3891 0.0119575
R32508 DVSS.n3116 DVSS.n3106 0.0119575
R32509 DVSS.n5809 DVSS.n3104 0.0119575
R32510 DVSS.n3115 DVSS.n3107 0.0119575
R32511 DVSS.n5810 DVSS.n3103 0.0119575
R32512 DVSS.n3114 DVSS.n3108 0.0119575
R32513 DVSS.n1984 DVSS.n1983 0.0119575
R32514 DVSS.n8007 DVSS.n1981 0.0119575
R32515 DVSS.n1986 DVSS.n1985 0.0119575
R32516 DVSS.n8008 DVSS.n1980 0.0119575
R32517 DVSS.n1988 DVSS.n1987 0.0119575
R32518 DVSS.n8009 DVSS.n1979 0.0119575
R32519 DVSS.n1990 DVSS.n1989 0.0119575
R32520 DVSS.n8010 DVSS.n1978 0.0119575
R32521 DVSS.n1992 DVSS.n1991 0.0119575
R32522 DVSS.n8012 DVSS.n1977 0.0119575
R32523 DVSS.n1173 DVSS.n1172 0.0119575
R32524 DVSS.n1174 DVSS.n1170 0.0119575
R32525 DVSS.n1176 DVSS.n1175 0.0119575
R32526 DVSS.n1169 DVSS.n1168 0.0119575
R32527 DVSS.n1166 DVSS.n1156 0.0119575
R32528 DVSS.n1177 DVSS.n1167 0.0119575
R32529 DVSS.n1179 DVSS.n1178 0.0119575
R32530 DVSS.n1180 DVSS.n1165 0.0119575
R32531 DVSS.n7416 DVSS.n2429 0.0119575
R32532 DVSS.n2432 DVSS.n2431 0.0119575
R32533 DVSS.n2433 DVSS.n2428 0.0119575
R32534 DVSS.n2435 DVSS.n2434 0.0119575
R32535 DVSS.n2436 DVSS.n2427 0.0119575
R32536 DVSS.n2438 DVSS.n2437 0.0119575
R32537 DVSS.n2439 DVSS.n2426 0.0119575
R32538 DVSS.n2441 DVSS.n2440 0.0119575
R32539 DVSS.n2442 DVSS.n2425 0.0119575
R32540 DVSS.n2444 DVSS.n2443 0.0119575
R32541 DVSS.n2445 DVSS.n2424 0.0119575
R32542 DVSS.n2447 DVSS.n2446 0.0119575
R32543 DVSS.n2448 DVSS.n2423 0.0119575
R32544 DVSS.n2450 DVSS.n2449 0.0119575
R32545 DVSS.n2451 DVSS.n2422 0.0119575
R32546 DVSS.n2453 DVSS.n2452 0.0119575
R32547 DVSS.n2454 DVSS.n2421 0.0119575
R32548 DVSS.n2456 DVSS.n2455 0.0119575
R32549 DVSS.n2457 DVSS.n2420 0.0119575
R32550 DVSS.n2459 DVSS.n2458 0.0119575
R32551 DVSS.n2460 DVSS.n2419 0.0119575
R32552 DVSS.n2462 DVSS.n2461 0.0119575
R32553 DVSS.n2463 DVSS.n2418 0.0119575
R32554 DVSS.n2366 DVSS.n2364 0.0119575
R32555 DVSS.n2368 DVSS.n2367 0.0119575
R32556 DVSS.n2369 DVSS.n2363 0.0119575
R32557 DVSS.n2371 DVSS.n2370 0.0119575
R32558 DVSS.n2372 DVSS.n2362 0.0119575
R32559 DVSS.n2374 DVSS.n2373 0.0119575
R32560 DVSS.n2375 DVSS.n2361 0.0119575
R32561 DVSS.n2377 DVSS.n2376 0.0119575
R32562 DVSS.n2378 DVSS.n2360 0.0119575
R32563 DVSS.n2380 DVSS.n2379 0.0119575
R32564 DVSS.n2381 DVSS.n2359 0.0119575
R32565 DVSS.n2383 DVSS.n2382 0.0119575
R32566 DVSS.n2384 DVSS.n2358 0.0119575
R32567 DVSS.n2386 DVSS.n2385 0.0119575
R32568 DVSS.n2387 DVSS.n2357 0.0119575
R32569 DVSS.n2389 DVSS.n2388 0.0119575
R32570 DVSS.n2390 DVSS.n2356 0.0119575
R32571 DVSS.n2392 DVSS.n2391 0.0119575
R32572 DVSS.n2393 DVSS.n2355 0.0119575
R32573 DVSS.n2395 DVSS.n2394 0.0119575
R32574 DVSS.n2396 DVSS.n2354 0.0119575
R32575 DVSS.n2398 DVSS.n2397 0.0119575
R32576 DVSS.n2399 DVSS.n2353 0.0119575
R32577 DVSS.n7543 DVSS.n2250 0.0119575
R32578 DVSS.n7532 DVSS.n2249 0.0119575
R32579 DVSS.n7544 DVSS.n2264 0.0119575
R32580 DVSS.n7533 DVSS.n2248 0.0119575
R32581 DVSS.n7545 DVSS.n2263 0.0119575
R32582 DVSS.n7534 DVSS.n2247 0.0119575
R32583 DVSS.n7546 DVSS.n2262 0.0119575
R32584 DVSS.n7535 DVSS.n2246 0.0119575
R32585 DVSS.n7547 DVSS.n2261 0.0119575
R32586 DVSS.n7536 DVSS.n2245 0.0119575
R32587 DVSS.n7548 DVSS.n2260 0.0119575
R32588 DVSS.n7537 DVSS.n2244 0.0119575
R32589 DVSS.n7549 DVSS.n2259 0.0119575
R32590 DVSS.n7538 DVSS.n2243 0.0119575
R32591 DVSS.n7550 DVSS.n2258 0.0119575
R32592 DVSS.n7539 DVSS.n2242 0.0119575
R32593 DVSS.n7551 DVSS.n2257 0.0119575
R32594 DVSS.n7540 DVSS.n2241 0.0119575
R32595 DVSS.n7552 DVSS.n2256 0.0119575
R32596 DVSS.n7541 DVSS.n2240 0.0119575
R32597 DVSS.n7554 DVSS.n2255 0.0119575
R32598 DVSS.n7555 DVSS.n2239 0.0119575
R32599 DVSS.n2254 DVSS.n2251 0.0119575
R32600 DVSS.n7601 DVSS.n2208 0.0119575
R32601 DVSS.n7590 DVSS.n2207 0.0119575
R32602 DVSS.n7602 DVSS.n2222 0.0119575
R32603 DVSS.n7591 DVSS.n2206 0.0119575
R32604 DVSS.n7603 DVSS.n2221 0.0119575
R32605 DVSS.n7592 DVSS.n2205 0.0119575
R32606 DVSS.n7604 DVSS.n2220 0.0119575
R32607 DVSS.n7593 DVSS.n2204 0.0119575
R32608 DVSS.n7605 DVSS.n2219 0.0119575
R32609 DVSS.n7594 DVSS.n2203 0.0119575
R32610 DVSS.n7606 DVSS.n2218 0.0119575
R32611 DVSS.n7595 DVSS.n2202 0.0119575
R32612 DVSS.n7607 DVSS.n2217 0.0119575
R32613 DVSS.n7596 DVSS.n2201 0.0119575
R32614 DVSS.n7608 DVSS.n2216 0.0119575
R32615 DVSS.n7597 DVSS.n2200 0.0119575
R32616 DVSS.n7609 DVSS.n2215 0.0119575
R32617 DVSS.n7598 DVSS.n2199 0.0119575
R32618 DVSS.n7610 DVSS.n2214 0.0119575
R32619 DVSS.n7599 DVSS.n2198 0.0119575
R32620 DVSS.n7612 DVSS.n2213 0.0119575
R32621 DVSS.n7613 DVSS.n2197 0.0119575
R32622 DVSS.n2212 DVSS.n2209 0.0119575
R32623 DVSS.n2489 DVSS.n2487 0.0119575
R32624 DVSS.n2488 DVSS.n2484 0.0119575
R32625 DVSS.n2492 DVSS.n2490 0.0119575
R32626 DVSS.n2491 DVSS.n2483 0.0119575
R32627 DVSS.n2495 DVSS.n2493 0.0119575
R32628 DVSS.n2494 DVSS.n2482 0.0119575
R32629 DVSS.n2498 DVSS.n2496 0.0119575
R32630 DVSS.n2497 DVSS.n2481 0.0119575
R32631 DVSS.n2501 DVSS.n2499 0.0119575
R32632 DVSS.n2500 DVSS.n2480 0.0119575
R32633 DVSS.n2504 DVSS.n2502 0.0119575
R32634 DVSS.n2503 DVSS.n2479 0.0119575
R32635 DVSS.n2507 DVSS.n2505 0.0119575
R32636 DVSS.n2506 DVSS.n2478 0.0119575
R32637 DVSS.n2510 DVSS.n2508 0.0119575
R32638 DVSS.n2509 DVSS.n2477 0.0119575
R32639 DVSS.n2513 DVSS.n2511 0.0119575
R32640 DVSS.n2512 DVSS.n2476 0.0119575
R32641 DVSS.n2516 DVSS.n2514 0.0119575
R32642 DVSS.n2515 DVSS.n2475 0.0119575
R32643 DVSS.n2519 DVSS.n2517 0.0119575
R32644 DVSS.n2518 DVSS.n2474 0.0119575
R32645 DVSS.n7398 DVSS.n2520 0.0119575
R32646 DVSS.n2679 DVSS.n2672 0.0119575
R32647 DVSS.n2673 DVSS.n2671 0.0119575
R32648 DVSS.n2675 DVSS.n2670 0.0119575
R32649 DVSS.n2669 DVSS.n2594 0.0119575
R32650 DVSS.n7360 DVSS.n2593 0.0119575
R32651 DVSS.n7357 DVSS.n7355 0.0119575
R32652 DVSS.n2597 DVSS.n2591 0.0119575
R32653 DVSS.n7354 DVSS.n7353 0.0119575
R32654 DVSS.n1957 DVSS.n1955 0.0119575
R32655 DVSS.n8030 DVSS.n1960 0.0119575
R32656 DVSS.n1959 DVSS.n1954 0.0119575
R32657 DVSS.n8031 DVSS.n1962 0.0119575
R32658 DVSS.n1961 DVSS.n1953 0.0119575
R32659 DVSS.n8032 DVSS.n1964 0.0119575
R32660 DVSS.n1963 DVSS.n1952 0.0119575
R32661 DVSS.n8033 DVSS.n1966 0.0119575
R32662 DVSS.n1965 DVSS.n1951 0.0119575
R32663 DVSS.n8036 DVSS.n8035 0.0119575
R32664 DVSS.n8075 DVSS.n1906 0.0119575
R32665 DVSS.n1907 DVSS.n1905 0.0119575
R32666 DVSS.n8071 DVSS.n1902 0.0119575
R32667 DVSS.n1904 DVSS.n1903 0.0119575
R32668 DVSS.n6674 DVSS.n6666 0.0119575
R32669 DVSS.n6677 DVSS.n6676 0.0119575
R32670 DVSS.n6688 DVSS.n6673 0.0119575
R32671 DVSS.n6679 DVSS.n6678 0.0119575
R32672 DVSS.n6687 DVSS.n6672 0.0119575
R32673 DVSS.n6681 DVSS.n6680 0.0119575
R32674 DVSS.n6686 DVSS.n6671 0.0119575
R32675 DVSS.n6683 DVSS.n6682 0.0119575
R32676 DVSS.n6685 DVSS.n6670 0.0119575
R32677 DVSS.n7061 DVSS.n6684 0.0119575
R32678 DVSS.n6706 DVSS.n6690 0.0119575
R32679 DVSS.n6705 DVSS.n6703 0.0119575
R32680 DVSS.n7046 DVSS.n6708 0.0119575
R32681 DVSS.n6707 DVSS.n6702 0.0119575
R32682 DVSS.n7047 DVSS.n6710 0.0119575
R32683 DVSS.n6709 DVSS.n6701 0.0119575
R32684 DVSS.n7048 DVSS.n6712 0.0119575
R32685 DVSS.n6711 DVSS.n6700 0.0119575
R32686 DVSS.n7049 DVSS.n6714 0.0119575
R32687 DVSS.n6713 DVSS.n6699 0.0119575
R32688 DVSS.n7050 DVSS.n6716 0.0119575
R32689 DVSS.n6715 DVSS.n6698 0.0119575
R32690 DVSS.n7051 DVSS.n6718 0.0119575
R32691 DVSS.n6717 DVSS.n6697 0.0119575
R32692 DVSS.n7052 DVSS.n6720 0.0119575
R32693 DVSS.n6719 DVSS.n6696 0.0119575
R32694 DVSS.n7053 DVSS.n6722 0.0119575
R32695 DVSS.n6721 DVSS.n6695 0.0119575
R32696 DVSS.n7054 DVSS.n6724 0.0119575
R32697 DVSS.n6723 DVSS.n6694 0.0119575
R32698 DVSS.n7058 DVSS.n7056 0.0119575
R32699 DVSS.n7057 DVSS.n784 0.0119575
R32700 DVSS.n2487 DVSS.n2485 0.0119575
R32701 DVSS.n2489 DVSS.n2488 0.0119575
R32702 DVSS.n2490 DVSS.n2484 0.0119575
R32703 DVSS.n2492 DVSS.n2491 0.0119575
R32704 DVSS.n2493 DVSS.n2483 0.0119575
R32705 DVSS.n2495 DVSS.n2494 0.0119575
R32706 DVSS.n2496 DVSS.n2482 0.0119575
R32707 DVSS.n2498 DVSS.n2497 0.0119575
R32708 DVSS.n2499 DVSS.n2481 0.0119575
R32709 DVSS.n2501 DVSS.n2500 0.0119575
R32710 DVSS.n2502 DVSS.n2480 0.0119575
R32711 DVSS.n2504 DVSS.n2503 0.0119575
R32712 DVSS.n2505 DVSS.n2479 0.0119575
R32713 DVSS.n2507 DVSS.n2506 0.0119575
R32714 DVSS.n2508 DVSS.n2478 0.0119575
R32715 DVSS.n2510 DVSS.n2509 0.0119575
R32716 DVSS.n2511 DVSS.n2477 0.0119575
R32717 DVSS.n2513 DVSS.n2512 0.0119575
R32718 DVSS.n2514 DVSS.n2476 0.0119575
R32719 DVSS.n2516 DVSS.n2515 0.0119575
R32720 DVSS.n2517 DVSS.n2475 0.0119575
R32721 DVSS.n2519 DVSS.n2518 0.0119575
R32722 DVSS.n2520 DVSS.n2474 0.0119575
R32723 DVSS.n1958 DVSS.n1957 0.0119575
R32724 DVSS.n8030 DVSS.n1955 0.0119575
R32725 DVSS.n1960 DVSS.n1959 0.0119575
R32726 DVSS.n8031 DVSS.n1954 0.0119575
R32727 DVSS.n1962 DVSS.n1961 0.0119575
R32728 DVSS.n8032 DVSS.n1953 0.0119575
R32729 DVSS.n1964 DVSS.n1963 0.0119575
R32730 DVSS.n8033 DVSS.n1952 0.0119575
R32731 DVSS.n1966 DVSS.n1965 0.0119575
R32732 DVSS.n8035 DVSS.n1951 0.0119575
R32733 DVSS.n7063 DVSS.n6666 0.0119575
R32734 DVSS.n6676 DVSS.n6674 0.0119575
R32735 DVSS.n6688 DVSS.n6677 0.0119575
R32736 DVSS.n6678 DVSS.n6673 0.0119575
R32737 DVSS.n6687 DVSS.n6679 0.0119575
R32738 DVSS.n6680 DVSS.n6672 0.0119575
R32739 DVSS.n6686 DVSS.n6681 0.0119575
R32740 DVSS.n6682 DVSS.n6671 0.0119575
R32741 DVSS.n6685 DVSS.n6683 0.0119575
R32742 DVSS.n6684 DVSS.n6670 0.0119575
R32743 DVSS.n3823 DVSS.n3822 0.0119575
R32744 DVSS.n4515 DVSS.n4514 0.0119575
R32745 DVSS.n4512 DVSS.n3820 0.0119575
R32746 DVSS.n4513 DVSS.n4511 0.0119575
R32747 DVSS.n4509 DVSS.n3821 0.0119575
R32748 DVSS.n4510 DVSS.n3817 0.0119575
R32749 DVSS.n4228 DVSS.n4227 0.0119575
R32750 DVSS.n4254 DVSS.n4218 0.0119575
R32751 DVSS.n4253 DVSS.n4226 0.0119575
R32752 DVSS.n4256 DVSS.n4219 0.0119575
R32753 DVSS.n4255 DVSS.n4225 0.0119575
R32754 DVSS.n4257 DVSS.n4220 0.0119575
R32755 DVSS.n4227 DVSS.n4217 0.0119575
R32756 DVSS.n4228 DVSS.n4218 0.0119575
R32757 DVSS.n4254 DVSS.n4253 0.0119575
R32758 DVSS.n4226 DVSS.n4219 0.0119575
R32759 DVSS.n4256 DVSS.n4255 0.0119575
R32760 DVSS.n4225 DVSS.n4220 0.0119575
R32761 DVSS.n4515 DVSS.n3819 0.0119575
R32762 DVSS.n4514 DVSS.n3820 0.0119575
R32763 DVSS.n4513 DVSS.n4512 0.0119575
R32764 DVSS.n4511 DVSS.n3821 0.0119575
R32765 DVSS.n4510 DVSS.n4509 0.0119575
R32766 DVSS.n3822 DVSS.n3816 0.0119575
R32767 DVSS.n4581 DVSS.n4580 0.0119575
R32768 DVSS.n4582 DVSS.n3807 0.0119575
R32769 DVSS.n4584 DVSS.n4583 0.0119575
R32770 DVSS.n4585 DVSS.n3806 0.0119575
R32771 DVSS.n4587 DVSS.n4586 0.0119575
R32772 DVSS.n3804 DVSS.n3803 0.0119575
R32773 DVSS.n3746 DVSS.n3736 0.0119575
R32774 DVSS.n3737 DVSS.n3733 0.0119575
R32775 DVSS.n3745 DVSS.n3738 0.0119575
R32776 DVSS.n3739 DVSS.n3732 0.0119575
R32777 DVSS.n3740 DVSS.n3727 0.0119575
R32778 DVSS.n3741 DVSS.n3731 0.0119575
R32779 DVSS.n6004 DVSS.n2780 0.0119575
R32780 DVSS.n2790 DVSS.n2788 0.0119575
R32781 DVSS.n2793 DVSS.n2791 0.0119575
R32782 DVSS.n2792 DVSS.n2787 0.0119575
R32783 DVSS.n6002 DVSS.n6001 0.0119575
R32784 DVSS.n2785 DVSS.n2784 0.0119575
R32785 DVSS.n2836 DVSS.n2823 0.0119575
R32786 DVSS.n2828 DVSS.n2820 0.0119575
R32787 DVSS.n2835 DVSS.n2824 0.0119575
R32788 DVSS.n2829 DVSS.n2819 0.0119575
R32789 DVSS.n2834 DVSS.n2825 0.0119575
R32790 DVSS.n2832 DVSS.n2817 0.0119575
R32791 DVSS.n2859 DVSS.n2848 0.0119575
R32792 DVSS.n2862 DVSS.n2851 0.0119575
R32793 DVSS.n5956 DVSS.n2855 0.0119575
R32794 DVSS.n2861 DVSS.n2850 0.0119575
R32795 DVSS.n5957 DVSS.n2856 0.0119575
R32796 DVSS.n2860 DVSS.n2849 0.0119575
R32797 DVSS.n4962 DVSS.n3604 0.0119575
R32798 DVSS.n4966 DVSS.n4964 0.0119575
R32799 DVSS.n4965 DVSS.n3603 0.0119575
R32800 DVSS.n4969 DVSS.n4967 0.0119575
R32801 DVSS.n4968 DVSS.n3602 0.0119575
R32802 DVSS.n4971 DVSS.n4970 0.0119575
R32803 DVSS.n3389 DVSS.n3383 0.0119575
R32804 DVSS.n5348 DVSS.n3392 0.0119575
R32805 DVSS.n3391 DVSS.n3382 0.0119575
R32806 DVSS.n5352 DVSS.n5350 0.0119575
R32807 DVSS.n5351 DVSS.n3381 0.0119575
R32808 DVSS.n5354 DVSS.n3377 0.0119575
R32809 DVSS.n5357 DVSS.n5356 0.0119575
R32810 DVSS.n5361 DVSS.n5358 0.0119575
R32811 DVSS.n5363 DVSS.n5362 0.0119575
R32812 DVSS.n5364 DVSS.n5360 0.0119575
R32813 DVSS.n5359 DVSS.n3375 0.0119575
R32814 DVSS.n5514 DVSS.n5510 0.0119575
R32815 DVSS.n5511 DVSS.n3313 0.0119575
R32816 DVSS.n5508 DVSS.n3312 0.0119575
R32817 DVSS.n5516 DVSS.n3308 0.0119575
R32818 DVSS.n5527 DVSS.n3307 0.0119575
R32819 DVSS.n5524 DVSS.n5522 0.0119575
R32820 DVSS.n5519 DVSS.n3305 0.0119575
R32821 DVSS.n5521 DVSS.n5520 0.0119575
R32822 DVSS.n7643 DVSS.n7632 0.0119575
R32823 DVSS.n2188 DVSS.n2173 0.0119575
R32824 DVSS.n7644 DVSS.n7633 0.0119575
R32825 DVSS.n2187 DVSS.n2172 0.0119575
R32826 DVSS.n7645 DVSS.n7634 0.0119575
R32827 DVSS.n2186 DVSS.n2171 0.0119575
R32828 DVSS.n7646 DVSS.n7635 0.0119575
R32829 DVSS.n2185 DVSS.n2170 0.0119575
R32830 DVSS.n7647 DVSS.n7636 0.0119575
R32831 DVSS.n2184 DVSS.n2169 0.0119575
R32832 DVSS.n7648 DVSS.n7637 0.0119575
R32833 DVSS.n2183 DVSS.n2168 0.0119575
R32834 DVSS.n7649 DVSS.n7638 0.0119575
R32835 DVSS.n2182 DVSS.n2167 0.0119575
R32836 DVSS.n7650 DVSS.n7639 0.0119575
R32837 DVSS.n2181 DVSS.n2166 0.0119575
R32838 DVSS.n7651 DVSS.n7640 0.0119575
R32839 DVSS.n2180 DVSS.n2165 0.0119575
R32840 DVSS.n7652 DVSS.n7641 0.0119575
R32841 DVSS.n2179 DVSS.n2164 0.0119575
R32842 DVSS.n7655 DVSS.n7654 0.0119575
R32843 DVSS.n2178 DVSS.n2163 0.0119575
R32844 DVSS.n7657 DVSS.n2175 0.0119575
R32845 DVSS.n2737 DVSS.n2736 0.0119575
R32846 DVSS.n2734 DVSS.n2728 0.0119575
R32847 DVSS.n2733 DVSS.n2726 0.0119575
R32848 DVSS.n2732 DVSS.n2102 0.0119575
R32849 DVSS.n7717 DVSS.n2101 0.0119575
R32850 DVSS.n7714 DVSS.n7712 0.0119575
R32851 DVSS.n2105 DVSS.n2099 0.0119575
R32852 DVSS.n7711 DVSS.n7710 0.0119575
R32853 DVSS.n8143 DVSS.n1800 0.0119575
R32854 DVSS.n8139 DVSS.n1790 0.0119575
R32855 DVSS.n8142 DVSS.n1799 0.0119575
R32856 DVSS.n8140 DVSS.n1791 0.0119575
R32857 DVSS.n8141 DVSS.n1798 0.0119575
R32858 DVSS.n8147 DVSS.n1792 0.0119575
R32859 DVSS.n8146 DVSS.n1797 0.0119575
R32860 DVSS.n8148 DVSS.n1793 0.0119575
R32861 DVSS.n8150 DVSS.n1795 0.0119575
R32862 DVSS.n8151 DVSS.n1794 0.0119575
R32863 DVSS.n1850 DVSS.n1840 0.0119575
R32864 DVSS.n1847 DVSS.n1845 0.0119575
R32865 DVSS.n1844 DVSS.n1838 0.0119575
R32866 DVSS.n1843 DVSS.n1560 0.0119575
R32867 DVSS.n1718 DVSS.n1605 0.0119575
R32868 DVSS.n1714 DVSS.n1595 0.0119575
R32869 DVSS.n1717 DVSS.n1604 0.0119575
R32870 DVSS.n1715 DVSS.n1596 0.0119575
R32871 DVSS.n1716 DVSS.n1603 0.0119575
R32872 DVSS.n1722 DVSS.n1597 0.0119575
R32873 DVSS.n1721 DVSS.n1602 0.0119575
R32874 DVSS.n1723 DVSS.n1598 0.0119575
R32875 DVSS.n1725 DVSS.n1600 0.0119575
R32876 DVSS.n1726 DVSS.n1599 0.0119575
R32877 DVSS.n9737 DVSS.n9736 0.0119575
R32878 DVSS.n9739 DVSS.n154 0.0119575
R32879 DVSS.n9740 DVSS.n9738 0.0119575
R32880 DVSS.n9742 DVSS.n153 0.0119575
R32881 DVSS.n9743 DVSS.n9741 0.0119575
R32882 DVSS.n9745 DVSS.n152 0.0119575
R32883 DVSS.n9746 DVSS.n9744 0.0119575
R32884 DVSS.n9748 DVSS.n151 0.0119575
R32885 DVSS.n9749 DVSS.n9747 0.0119575
R32886 DVSS.n9751 DVSS.n150 0.0119575
R32887 DVSS.n9752 DVSS.n9750 0.0119575
R32888 DVSS.n9754 DVSS.n149 0.0119575
R32889 DVSS.n9755 DVSS.n9753 0.0119575
R32890 DVSS.n9757 DVSS.n148 0.0119575
R32891 DVSS.n9758 DVSS.n9756 0.0119575
R32892 DVSS.n9760 DVSS.n147 0.0119575
R32893 DVSS.n9761 DVSS.n9759 0.0119575
R32894 DVSS.n9763 DVSS.n146 0.0119575
R32895 DVSS.n9764 DVSS.n9762 0.0119575
R32896 DVSS.n9766 DVSS.n145 0.0119575
R32897 DVSS.n9767 DVSS.n9765 0.0119575
R32898 DVSS.n9734 DVSS.n144 0.0119575
R32899 DVSS.n2862 DVSS.n2854 0.0119575
R32900 DVSS.n5956 DVSS.n2851 0.0119575
R32901 DVSS.n2861 DVSS.n2855 0.0119575
R32902 DVSS.n5957 DVSS.n2850 0.0119575
R32903 DVSS.n2860 DVSS.n2856 0.0119575
R32904 DVSS.n4963 DVSS.n4962 0.0119575
R32905 DVSS.n4964 DVSS.n3604 0.0119575
R32906 DVSS.n4966 DVSS.n4965 0.0119575
R32907 DVSS.n4967 DVSS.n3603 0.0119575
R32908 DVSS.n4969 DVSS.n4968 0.0119575
R32909 DVSS.n4970 DVSS.n3602 0.0119575
R32910 DVSS.n3390 DVSS.n3389 0.0119575
R32911 DVSS.n5348 DVSS.n3383 0.0119575
R32912 DVSS.n3392 DVSS.n3391 0.0119575
R32913 DVSS.n5350 DVSS.n3382 0.0119575
R32914 DVSS.n5352 DVSS.n5351 0.0119575
R32915 DVSS.n3381 DVSS.n3377 0.0119575
R32916 DVSS.n5356 DVSS.n5355 0.0119575
R32917 DVSS.n5358 DVSS.n5357 0.0119575
R32918 DVSS.n5362 DVSS.n5361 0.0119575
R32919 DVSS.n5364 DVSS.n5363 0.0119575
R32920 DVSS.n5360 DVSS.n5359 0.0119575
R32921 DVSS.n7643 DVSS.n2174 0.0119575
R32922 DVSS.n7632 DVSS.n2173 0.0119575
R32923 DVSS.n7644 DVSS.n2188 0.0119575
R32924 DVSS.n7633 DVSS.n2172 0.0119575
R32925 DVSS.n7645 DVSS.n2187 0.0119575
R32926 DVSS.n7634 DVSS.n2171 0.0119575
R32927 DVSS.n7646 DVSS.n2186 0.0119575
R32928 DVSS.n7635 DVSS.n2170 0.0119575
R32929 DVSS.n7647 DVSS.n2185 0.0119575
R32930 DVSS.n7636 DVSS.n2169 0.0119575
R32931 DVSS.n7648 DVSS.n2184 0.0119575
R32932 DVSS.n7637 DVSS.n2168 0.0119575
R32933 DVSS.n7649 DVSS.n2183 0.0119575
R32934 DVSS.n7638 DVSS.n2167 0.0119575
R32935 DVSS.n7650 DVSS.n2182 0.0119575
R32936 DVSS.n7639 DVSS.n2166 0.0119575
R32937 DVSS.n7651 DVSS.n2181 0.0119575
R32938 DVSS.n7640 DVSS.n2165 0.0119575
R32939 DVSS.n7652 DVSS.n2180 0.0119575
R32940 DVSS.n7641 DVSS.n2164 0.0119575
R32941 DVSS.n7654 DVSS.n2179 0.0119575
R32942 DVSS.n7655 DVSS.n2163 0.0119575
R32943 DVSS.n2178 DVSS.n2175 0.0119575
R32944 DVSS.n8143 DVSS.n1789 0.0119575
R32945 DVSS.n1800 DVSS.n1790 0.0119575
R32946 DVSS.n8142 DVSS.n8139 0.0119575
R32947 DVSS.n1799 DVSS.n1791 0.0119575
R32948 DVSS.n8141 DVSS.n8140 0.0119575
R32949 DVSS.n1798 DVSS.n1792 0.0119575
R32950 DVSS.n8147 DVSS.n8146 0.0119575
R32951 DVSS.n1797 DVSS.n1793 0.0119575
R32952 DVSS.n8148 DVSS.n1795 0.0119575
R32953 DVSS.n8151 DVSS.n8150 0.0119575
R32954 DVSS.n1718 DVSS.n1557 0.0119575
R32955 DVSS.n1605 DVSS.n1595 0.0119575
R32956 DVSS.n1717 DVSS.n1714 0.0119575
R32957 DVSS.n1604 DVSS.n1596 0.0119575
R32958 DVSS.n1716 DVSS.n1715 0.0119575
R32959 DVSS.n1603 DVSS.n1597 0.0119575
R32960 DVSS.n1722 DVSS.n1721 0.0119575
R32961 DVSS.n1602 DVSS.n1598 0.0119575
R32962 DVSS.n1723 DVSS.n1600 0.0119575
R32963 DVSS.n1726 DVSS.n1725 0.0119575
R32964 DVSS.n2859 DVSS.n2857 0.0119575
R32965 DVSS.n711 DVSS.n710 0.0119575
R32966 DVSS.n704 DVSS.n703 0.0119575
R32967 DVSS.n9375 DVSS.n9374 0.0119575
R32968 DVSS.n9540 DVSS.n9539 0.0119575
R32969 DVSS.n9005 DVSS.n708 0.0119575
R32970 DVSS.n9011 DVSS.n701 0.0119575
R32971 DVSS.n9372 DVSS.n390 0.0119575
R32972 DVSS.n9538 DVSS.n328 0.0119575
R32973 DVSS.n9009 DVSS.n713 0.0119575
R32974 DVSS.n9015 DVSS.n706 0.0119575
R32975 DVSS.n9377 DVSS.n9369 0.0119575
R32976 DVSS.n9542 DVSS.n324 0.0119575
R32977 DVSS.n8876 DVSS.n794 0.0119575
R32978 DVSS.n8871 DVSS.n804 0.0119575
R32979 DVSS.n9401 DVSS.n370 0.0119575
R32980 DVSS.n9410 DVSS.n368 0.0119575
R32981 DVSS.n795 DVSS.n788 0.0119575
R32982 DVSS.n805 DVSS.n798 0.0119575
R32983 DVSS.n9396 DVSS.n224 0.0119575
R32984 DVSS.n9405 DVSS.n185 0.0119575
R32985 DVSS.n5929 DVSS.n2886 0.0119575
R32986 DVSS.n5933 DVSS.n2880 0.0119575
R32987 DVSS.n2888 DVSS.n2884 0.0119575
R32988 DVSS.n5932 DVSS.n2879 0.0119575
R32989 DVSS.n2889 DVSS.n2885 0.0119575
R32990 DVSS.n5931 DVSS.n2878 0.0119575
R32991 DVSS.n4921 DVSS.n4911 0.0119575
R32992 DVSS.n4923 DVSS.n4914 0.0119575
R32993 DVSS.n4920 DVSS.n4910 0.0119575
R32994 DVSS.n4924 DVSS.n4915 0.0119575
R32995 DVSS.n4919 DVSS.n4909 0.0119575
R32996 DVSS.n4925 DVSS.n4916 0.0119575
R32997 DVSS.n2929 DVSS.n2928 0.0119575
R32998 DVSS.n2935 DVSS.n2933 0.0119575
R32999 DVSS.n2934 DVSS.n2927 0.0119575
R33000 DVSS.n2938 DVSS.n2936 0.0119575
R33001 DVSS.n2937 DVSS.n2926 0.0119575
R33002 DVSS.n5914 DVSS.n2939 0.0119575
R33003 DVSS.n2948 DVSS.n2940 0.0119575
R33004 DVSS.n2951 DVSS.n2950 0.0119575
R33005 DVSS.n2958 DVSS.n2947 0.0119575
R33006 DVSS.n2953 DVSS.n2952 0.0119575
R33007 DVSS.n2957 DVSS.n2946 0.0119575
R33008 DVSS.n7679 DVSS.n2136 0.0119575
R33009 DVSS.n2135 DVSS.n2132 0.0119575
R33010 DVSS.n7680 DVSS.n2138 0.0119575
R33011 DVSS.n2137 DVSS.n2131 0.0119575
R33012 DVSS.n7681 DVSS.n2140 0.0119575
R33013 DVSS.n2139 DVSS.n2130 0.0119575
R33014 DVSS.n7682 DVSS.n2142 0.0119575
R33015 DVSS.n2141 DVSS.n2129 0.0119575
R33016 DVSS.n7683 DVSS.n2144 0.0119575
R33017 DVSS.n2143 DVSS.n2128 0.0119575
R33018 DVSS.n7684 DVSS.n2146 0.0119575
R33019 DVSS.n2145 DVSS.n2127 0.0119575
R33020 DVSS.n7685 DVSS.n2148 0.0119575
R33021 DVSS.n2147 DVSS.n2126 0.0119575
R33022 DVSS.n7686 DVSS.n2150 0.0119575
R33023 DVSS.n2149 DVSS.n2125 0.0119575
R33024 DVSS.n7687 DVSS.n2152 0.0119575
R33025 DVSS.n2151 DVSS.n2124 0.0119575
R33026 DVSS.n7688 DVSS.n2154 0.0119575
R33027 DVSS.n2153 DVSS.n2123 0.0119575
R33028 DVSS.n7692 DVSS.n7690 0.0119575
R33029 DVSS.n7691 DVSS.n2122 0.0119575
R33030 DVSS.n7694 DVSS.n2118 0.0119575
R33031 DVSS.n1771 DVSS.n1769 0.0119575
R33032 DVSS.n8171 DVSS.n1774 0.0119575
R33033 DVSS.n1773 DVSS.n1768 0.0119575
R33034 DVSS.n8172 DVSS.n1776 0.0119575
R33035 DVSS.n1775 DVSS.n1767 0.0119575
R33036 DVSS.n8173 DVSS.n1778 0.0119575
R33037 DVSS.n1777 DVSS.n1766 0.0119575
R33038 DVSS.n8177 DVSS.n8175 0.0119575
R33039 DVSS.n8176 DVSS.n1765 0.0119575
R33040 DVSS.n8179 DVSS.n1761 0.0119575
R33041 DVSS.n1570 DVSS.n1562 0.0119575
R33042 DVSS.n1573 DVSS.n1572 0.0119575
R33043 DVSS.n1584 DVSS.n1569 0.0119575
R33044 DVSS.n1575 DVSS.n1574 0.0119575
R33045 DVSS.n1583 DVSS.n1568 0.0119575
R33046 DVSS.n1577 DVSS.n1576 0.0119575
R33047 DVSS.n1582 DVSS.n1567 0.0119575
R33048 DVSS.n1579 DVSS.n1578 0.0119575
R33049 DVSS.n1581 DVSS.n1566 0.0119575
R33050 DVSS.n1747 DVSS.n1580 0.0119575
R33051 DVSS.n9789 DVSS.n115 0.0119575
R33052 DVSS.n114 DVSS.n111 0.0119575
R33053 DVSS.n9790 DVSS.n117 0.0119575
R33054 DVSS.n116 DVSS.n110 0.0119575
R33055 DVSS.n9791 DVSS.n119 0.0119575
R33056 DVSS.n118 DVSS.n109 0.0119575
R33057 DVSS.n9792 DVSS.n121 0.0119575
R33058 DVSS.n120 DVSS.n108 0.0119575
R33059 DVSS.n9793 DVSS.n123 0.0119575
R33060 DVSS.n122 DVSS.n107 0.0119575
R33061 DVSS.n9794 DVSS.n125 0.0119575
R33062 DVSS.n124 DVSS.n106 0.0119575
R33063 DVSS.n9795 DVSS.n127 0.0119575
R33064 DVSS.n126 DVSS.n105 0.0119575
R33065 DVSS.n9796 DVSS.n129 0.0119575
R33066 DVSS.n128 DVSS.n104 0.0119575
R33067 DVSS.n9797 DVSS.n131 0.0119575
R33068 DVSS.n130 DVSS.n103 0.0119575
R33069 DVSS.n9798 DVSS.n133 0.0119575
R33070 DVSS.n132 DVSS.n102 0.0119575
R33071 DVSS.n9802 DVSS.n9800 0.0119575
R33072 DVSS.n9801 DVSS.n101 0.0119575
R33073 DVSS.n9804 DVSS.n97 0.0119575
R33074 DVSS.n9828 DVSS.n9807 0.0119575
R33075 DVSS.n9806 DVSS.n96 0.0119575
R33076 DVSS.n9829 DVSS.n9809 0.0119575
R33077 DVSS.n9808 DVSS.n95 0.0119575
R33078 DVSS.n9830 DVSS.n9811 0.0119575
R33079 DVSS.n9810 DVSS.n94 0.0119575
R33080 DVSS.n9831 DVSS.n9813 0.0119575
R33081 DVSS.n9812 DVSS.n93 0.0119575
R33082 DVSS.n9832 DVSS.n9815 0.0119575
R33083 DVSS.n9814 DVSS.n92 0.0119575
R33084 DVSS.n9833 DVSS.n9817 0.0119575
R33085 DVSS.n9816 DVSS.n91 0.0119575
R33086 DVSS.n9834 DVSS.n9819 0.0119575
R33087 DVSS.n9818 DVSS.n90 0.0119575
R33088 DVSS.n9835 DVSS.n9821 0.0119575
R33089 DVSS.n9820 DVSS.n89 0.0119575
R33090 DVSS.n9836 DVSS.n9823 0.0119575
R33091 DVSS.n9822 DVSS.n88 0.0119575
R33092 DVSS.n9837 DVSS.n9825 0.0119575
R33093 DVSS.n9824 DVSS.n87 0.0119575
R33094 DVSS.n9838 DVSS.n9827 0.0119575
R33095 DVSS.n9826 DVSS.n86 0.0119575
R33096 DVSS.n9842 DVSS.n9840 0.0119575
R33097 DVSS.n9919 DVSS.n9909 0.0119575
R33098 DVSS.n9908 DVSS.n16 0.0119575
R33099 DVSS.n9920 DVSS.n9910 0.0119575
R33100 DVSS.n9907 DVSS.n15 0.0119575
R33101 DVSS.n9921 DVSS.n9911 0.0119575
R33102 DVSS.n9906 DVSS.n14 0.0119575
R33103 DVSS.n9922 DVSS.n9912 0.0119575
R33104 DVSS.n9905 DVSS.n13 0.0119575
R33105 DVSS.n9923 DVSS.n9913 0.0119575
R33106 DVSS.n9904 DVSS.n12 0.0119575
R33107 DVSS.n9924 DVSS.n9914 0.0119575
R33108 DVSS.n9903 DVSS.n11 0.0119575
R33109 DVSS.n9925 DVSS.n9915 0.0119575
R33110 DVSS.n9902 DVSS.n10 0.0119575
R33111 DVSS.n9926 DVSS.n9916 0.0119575
R33112 DVSS.n9901 DVSS.n9 0.0119575
R33113 DVSS.n9927 DVSS.n9917 0.0119575
R33114 DVSS.n9900 DVSS.n8 0.0119575
R33115 DVSS.n9928 DVSS.n9918 0.0119575
R33116 DVSS.n9899 DVSS.n7 0.0119575
R33117 DVSS.n9931 DVSS.n9930 0.0119575
R33118 DVSS.n9898 DVSS.n6 0.0119575
R33119 DVSS.n9933 DVSS.n18 0.0119575
R33120 DVSS.n5933 DVSS.n2883 0.0119575
R33121 DVSS.n2888 DVSS.n2880 0.0119575
R33122 DVSS.n5932 DVSS.n2884 0.0119575
R33123 DVSS.n2889 DVSS.n2879 0.0119575
R33124 DVSS.n5931 DVSS.n2885 0.0119575
R33125 DVSS.n4921 DVSS.n4913 0.0119575
R33126 DVSS.n4923 DVSS.n4911 0.0119575
R33127 DVSS.n4920 DVSS.n4914 0.0119575
R33128 DVSS.n4924 DVSS.n4910 0.0119575
R33129 DVSS.n4919 DVSS.n4915 0.0119575
R33130 DVSS.n4925 DVSS.n4909 0.0119575
R33131 DVSS.n2928 DVSS.n2919 0.0119575
R33132 DVSS.n2933 DVSS.n2929 0.0119575
R33133 DVSS.n2935 DVSS.n2934 0.0119575
R33134 DVSS.n2936 DVSS.n2927 0.0119575
R33135 DVSS.n2938 DVSS.n2937 0.0119575
R33136 DVSS.n2939 DVSS.n2926 0.0119575
R33137 DVSS.n5913 DVSS.n2940 0.0119575
R33138 DVSS.n2950 DVSS.n2948 0.0119575
R33139 DVSS.n2958 DVSS.n2951 0.0119575
R33140 DVSS.n2952 DVSS.n2947 0.0119575
R33141 DVSS.n2957 DVSS.n2953 0.0119575
R33142 DVSS.n7679 DVSS.n2133 0.0119575
R33143 DVSS.n2136 DVSS.n2135 0.0119575
R33144 DVSS.n7680 DVSS.n2132 0.0119575
R33145 DVSS.n2138 DVSS.n2137 0.0119575
R33146 DVSS.n7681 DVSS.n2131 0.0119575
R33147 DVSS.n2140 DVSS.n2139 0.0119575
R33148 DVSS.n7682 DVSS.n2130 0.0119575
R33149 DVSS.n2142 DVSS.n2141 0.0119575
R33150 DVSS.n7683 DVSS.n2129 0.0119575
R33151 DVSS.n2144 DVSS.n2143 0.0119575
R33152 DVSS.n7684 DVSS.n2128 0.0119575
R33153 DVSS.n2146 DVSS.n2145 0.0119575
R33154 DVSS.n7685 DVSS.n2127 0.0119575
R33155 DVSS.n2148 DVSS.n2147 0.0119575
R33156 DVSS.n7686 DVSS.n2126 0.0119575
R33157 DVSS.n2150 DVSS.n2149 0.0119575
R33158 DVSS.n7687 DVSS.n2125 0.0119575
R33159 DVSS.n2152 DVSS.n2151 0.0119575
R33160 DVSS.n7688 DVSS.n2124 0.0119575
R33161 DVSS.n2154 DVSS.n2153 0.0119575
R33162 DVSS.n7690 DVSS.n2123 0.0119575
R33163 DVSS.n7692 DVSS.n7691 0.0119575
R33164 DVSS.n2122 DVSS.n2118 0.0119575
R33165 DVSS.n1772 DVSS.n1771 0.0119575
R33166 DVSS.n8171 DVSS.n1769 0.0119575
R33167 DVSS.n1774 DVSS.n1773 0.0119575
R33168 DVSS.n8172 DVSS.n1768 0.0119575
R33169 DVSS.n1776 DVSS.n1775 0.0119575
R33170 DVSS.n8173 DVSS.n1767 0.0119575
R33171 DVSS.n1778 DVSS.n1777 0.0119575
R33172 DVSS.n8175 DVSS.n1766 0.0119575
R33173 DVSS.n8177 DVSS.n8176 0.0119575
R33174 DVSS.n1765 DVSS.n1761 0.0119575
R33175 DVSS.n1749 DVSS.n1562 0.0119575
R33176 DVSS.n1572 DVSS.n1570 0.0119575
R33177 DVSS.n1584 DVSS.n1573 0.0119575
R33178 DVSS.n1574 DVSS.n1569 0.0119575
R33179 DVSS.n1583 DVSS.n1575 0.0119575
R33180 DVSS.n1576 DVSS.n1568 0.0119575
R33181 DVSS.n1582 DVSS.n1577 0.0119575
R33182 DVSS.n1578 DVSS.n1567 0.0119575
R33183 DVSS.n1581 DVSS.n1579 0.0119575
R33184 DVSS.n1580 DVSS.n1566 0.0119575
R33185 DVSS.n5929 DVSS.n2877 0.0119575
R33186 DVSS.n3249 DVSS.n3248 0.0119575
R33187 DVSS.n3240 DVSS.n3239 0.0119575
R33188 DVSS.n5397 DVSS.n5396 0.0119575
R33189 DVSS.n3317 DVSS.n3316 0.0119575
R33190 DVSS.n3312 DVSS.n3308 0.0119575
R33191 DVSS.n5678 DVSS.n3251 0.0119575
R33192 DVSS.n5685 DVSS.n3242 0.0119575
R33193 DVSS.n5495 DVSS.n5398 0.0119575
R33194 DVSS.n5502 DVSS.n3318 0.0119575
R33195 DVSS.n5508 DVSS.n3313 0.0119575
R33196 DVSS.n3252 DVSS.n3113 0.0119575
R33197 DVSS.n3243 DVSS.n3157 0.0119575
R33198 DVSS.n5399 DVSS.n5395 0.0119575
R33199 DVSS.n3319 DVSS.n3315 0.0119575
R33200 DVSS.n5510 DVSS.n3311 0.0119575
R33201 DVSS.n5682 DVSS.n3253 0.0119575
R33202 DVSS.n5689 DVSS.n3244 0.0119575
R33203 DVSS.n5499 DVSS.n5400 0.0119575
R33204 DVSS.n5506 DVSS.n3320 0.0119575
R33205 DVSS.n5514 DVSS.n5511 0.0119575
R33206 DVSS.n5656 DVSS.n3265 0.0119575
R33207 DVSS.n5646 DVSS.n3272 0.0119575
R33208 DVSS.n5539 DVSS.n3296 0.0119575
R33209 DVSS.n5529 DVSS.n3304 0.0119575
R33210 DVSS.n5520 DVSS.n5519 0.0119575
R33211 DVSS.n5660 DVSS.n3260 0.0119575
R33212 DVSS.n5650 DVSS.n3267 0.0119575
R33213 DVSS.n5543 DVSS.n3290 0.0119575
R33214 DVSS.n5533 DVSS.n3298 0.0119575
R33215 DVSS.n5524 DVSS.n3305 0.0119575
R33216 DVSS.n5663 DVSS.n5662 0.0119575
R33217 DVSS.n5653 DVSS.n5652 0.0119575
R33218 DVSS.n5546 DVSS.n5545 0.0119575
R33219 DVSS.n5536 DVSS.n5535 0.0119575
R33220 DVSS.n5527 DVSS.n5526 0.0119575
R33221 DVSS.n5658 DVSS.n3262 0.0119575
R33222 DVSS.n5648 DVSS.n3269 0.0119575
R33223 DVSS.n5541 DVSS.n3292 0.0119575
R33224 DVSS.n5531 DVSS.n3300 0.0119575
R33225 DVSS.n5522 DVSS.n3307 0.0119575
R33226 DVSS.n2670 DVSS.n2669 0.0119575
R33227 DVSS.n2663 DVSS.n2662 0.0119575
R33228 DVSS.n2655 DVSS.n2654 0.0119575
R33229 DVSS.n2716 DVSS.n2715 0.0119575
R33230 DVSS.n2725 DVSS.n2724 0.0119575
R33231 DVSS.n2733 DVSS.n2732 0.0119575
R33232 DVSS.n2675 DVSS.n2671 0.0119575
R33233 DVSS.n2681 DVSS.n2664 0.0119575
R33234 DVSS.n2688 DVSS.n2656 0.0119575
R33235 DVSS.n2745 DVSS.n2709 0.0119575
R33236 DVSS.n2739 DVSS.n2718 0.0119575
R33237 DVSS.n2734 DVSS.n2726 0.0119575
R33238 DVSS.n2672 DVSS.n2521 0.0119575
R33239 DVSS.n2665 DVSS.n2464 0.0119575
R33240 DVSS.n2657 DVSS.n2400 0.0119575
R33241 DVSS.n2748 DVSS.n2252 0.0119575
R33242 DVSS.n2742 DVSS.n2210 0.0119575
R33243 DVSS.n2737 DVSS.n2176 0.0119575
R33244 DVSS.n2679 DVSS.n2673 0.0119575
R33245 DVSS.n2685 DVSS.n2666 0.0119575
R33246 DVSS.n2692 DVSS.n2658 0.0119575
R33247 DVSS.n2747 DVSS.n2711 0.0119575
R33248 DVSS.n2741 DVSS.n2720 0.0119575
R33249 DVSS.n2736 DVSS.n2728 0.0119575
R33250 DVSS.n7353 DVSS.n2597 0.0119575
R33251 DVSS.n7344 DVSS.n2604 0.0119575
R33252 DVSS.n7334 DVSS.n2612 0.0119575
R33253 DVSS.n7727 DVSS.n2089 0.0119575
R33254 DVSS.n2098 DVSS.n2097 0.0119575
R33255 DVSS.n7710 DVSS.n2105 0.0119575
R33256 DVSS.n7357 DVSS.n2591 0.0119575
R33257 DVSS.n7348 DVSS.n2598 0.0119575
R33258 DVSS.n7338 DVSS.n2606 0.0119575
R33259 DVSS.n7851 DVSS.n2083 0.0119575
R33260 DVSS.n7721 DVSS.n2091 0.0119575
R33261 DVSS.n7714 DVSS.n2099 0.0119575
R33262 DVSS.n7360 DVSS.n7359 0.0119575
R33263 DVSS.n7351 DVSS.n7350 0.0119575
R33264 DVSS.n7341 DVSS.n7340 0.0119575
R33265 DVSS.n7854 DVSS.n7853 0.0119575
R33266 DVSS.n7724 DVSS.n7723 0.0119575
R33267 DVSS.n7717 DVSS.n7716 0.0119575
R33268 DVSS.n7355 DVSS.n2593 0.0119575
R33269 DVSS.n7346 DVSS.n2600 0.0119575
R33270 DVSS.n7336 DVSS.n2608 0.0119575
R33271 DVSS.n7849 DVSS.n2085 0.0119575
R33272 DVSS.n7719 DVSS.n2093 0.0119575
R33273 DVSS.n7712 DVSS.n2101 0.0119575
R33274 DVSS.n1903 DVSS.n1902 0.0119575
R33275 DVSS.n1894 DVSS.n1893 0.0119575
R33276 DVSS.n1884 DVSS.n1883 0.0119575
R33277 DVSS.n1858 DVSS.n1857 0.0119575
R33278 DVSS.n1837 DVSS.n1836 0.0119575
R33279 DVSS.n1844 DVSS.n1843 0.0119575
R33280 DVSS.n8071 DVSS.n1905 0.0119575
R33281 DVSS.n8077 DVSS.n1896 0.0119575
R33282 DVSS.n8084 DVSS.n1886 0.0119575
R33283 DVSS.n8106 DVSS.n1860 0.0119575
R33284 DVSS.n8113 DVSS.n1852 0.0119575
R33285 DVSS.n1847 DVSS.n1838 0.0119575
R33286 DVSS.n1906 DVSS.n1901 0.0119575
R33287 DVSS.n1897 DVSS.n1892 0.0119575
R33288 DVSS.n1887 DVSS.n1882 0.0119575
R33289 DVSS.n1861 DVSS.n1856 0.0119575
R33290 DVSS.n8119 DVSS.n1834 0.0119575
R33291 DVSS.n1850 DVSS.n1849 0.0119575
R33292 DVSS.n8075 DVSS.n1907 0.0119575
R33293 DVSS.n8081 DVSS.n1898 0.0119575
R33294 DVSS.n8088 DVSS.n1888 0.0119575
R33295 DVSS.n8110 DVSS.n1862 0.0119575
R33296 DVSS.n8117 DVSS.n1853 0.0119575
R33297 DVSS.n1845 DVSS.n1840 0.0119575
R33298 DVSS.n4459 DVSS.n4458 0.0119575
R33299 DVSS.n4488 DVSS.n4487 0.0119575
R33300 DVSS.n4485 DVSS.n4456 0.0119575
R33301 DVSS.n4486 DVSS.n4484 0.0119575
R33302 DVSS.n4482 DVSS.n4457 0.0119575
R33303 DVSS.n4483 DVSS.n4453 0.0119575
R33304 DVSS.n3844 DVSS.n3836 0.0119575
R33305 DVSS.n3847 DVSS.n3846 0.0119575
R33306 DVSS.n3855 DVSS.n3843 0.0119575
R33307 DVSS.n3849 DVSS.n3848 0.0119575
R33308 DVSS.n3854 DVSS.n3842 0.0119575
R33309 DVSS.n3851 DVSS.n3850 0.0119575
R33310 DVSS.n3034 DVSS.n3033 0.0119575
R33311 DVSS.n5858 DVSS.n5856 0.0119575
R33312 DVSS.n5857 DVSS.n3032 0.0119575
R33313 DVSS.n5861 DVSS.n5859 0.0119575
R33314 DVSS.n5860 DVSS.n3031 0.0119575
R33315 DVSS.n5863 DVSS.n5862 0.0119575
R33316 DVSS.n3004 DVSS.n3002 0.0119575
R33317 DVSS.n3008 DVSS.n3006 0.0119575
R33318 DVSS.n3007 DVSS.n3001 0.0119575
R33319 DVSS.n3011 DVSS.n3009 0.0119575
R33320 DVSS.n3010 DVSS.n3000 0.0119575
R33321 DVSS.n2546 DVSS.n2544 0.0119575
R33322 DVSS.n2545 DVSS.n2541 0.0119575
R33323 DVSS.n2549 DVSS.n2547 0.0119575
R33324 DVSS.n2548 DVSS.n2540 0.0119575
R33325 DVSS.n2552 DVSS.n2550 0.0119575
R33326 DVSS.n2551 DVSS.n2539 0.0119575
R33327 DVSS.n2555 DVSS.n2553 0.0119575
R33328 DVSS.n2554 DVSS.n2538 0.0119575
R33329 DVSS.n2558 DVSS.n2556 0.0119575
R33330 DVSS.n2557 DVSS.n2537 0.0119575
R33331 DVSS.n2561 DVSS.n2559 0.0119575
R33332 DVSS.n2560 DVSS.n2536 0.0119575
R33333 DVSS.n2564 DVSS.n2562 0.0119575
R33334 DVSS.n2563 DVSS.n2535 0.0119575
R33335 DVSS.n2567 DVSS.n2565 0.0119575
R33336 DVSS.n2566 DVSS.n2534 0.0119575
R33337 DVSS.n2570 DVSS.n2568 0.0119575
R33338 DVSS.n2569 DVSS.n2533 0.0119575
R33339 DVSS.n2573 DVSS.n2571 0.0119575
R33340 DVSS.n2572 DVSS.n2532 0.0119575
R33341 DVSS.n2576 DVSS.n2574 0.0119575
R33342 DVSS.n2575 DVSS.n2531 0.0119575
R33343 DVSS.n7379 DVSS.n2577 0.0119575
R33344 DVSS.n1926 DVSS.n1924 0.0119575
R33345 DVSS.n8053 DVSS.n1929 0.0119575
R33346 DVSS.n1928 DVSS.n1923 0.0119575
R33347 DVSS.n8054 DVSS.n1931 0.0119575
R33348 DVSS.n1930 DVSS.n1922 0.0119575
R33349 DVSS.n8055 DVSS.n1933 0.0119575
R33350 DVSS.n1932 DVSS.n1921 0.0119575
R33351 DVSS.n8059 DVSS.n8057 0.0119575
R33352 DVSS.n8058 DVSS.n1920 0.0119575
R33353 DVSS.n8061 DVSS.n1916 0.0119575
R33354 DVSS.n6754 DVSS.n6743 0.0119575
R33355 DVSS.n6851 DVSS.n6757 0.0119575
R33356 DVSS.n6756 DVSS.n6742 0.0119575
R33357 DVSS.n6852 DVSS.n6759 0.0119575
R33358 DVSS.n6758 DVSS.n6741 0.0119575
R33359 DVSS.n6853 DVSS.n6761 0.0119575
R33360 DVSS.n6760 DVSS.n6740 0.0119575
R33361 DVSS.n6857 DVSS.n6855 0.0119575
R33362 DVSS.n6856 DVSS.n6739 0.0119575
R33363 DVSS.n6859 DVSS.n6735 0.0119575
R33364 DVSS.n6887 DVSS.n6861 0.0119575
R33365 DVSS.n6904 DVSS.n6884 0.0119575
R33366 DVSS.n6888 DVSS.n6862 0.0119575
R33367 DVSS.n6903 DVSS.n6883 0.0119575
R33368 DVSS.n6889 DVSS.n6863 0.0119575
R33369 DVSS.n6902 DVSS.n6882 0.0119575
R33370 DVSS.n6890 DVSS.n6864 0.0119575
R33371 DVSS.n6901 DVSS.n6881 0.0119575
R33372 DVSS.n6891 DVSS.n6865 0.0119575
R33373 DVSS.n6900 DVSS.n6880 0.0119575
R33374 DVSS.n6892 DVSS.n6866 0.0119575
R33375 DVSS.n6899 DVSS.n6879 0.0119575
R33376 DVSS.n6893 DVSS.n6867 0.0119575
R33377 DVSS.n6898 DVSS.n6878 0.0119575
R33378 DVSS.n6894 DVSS.n6868 0.0119575
R33379 DVSS.n6897 DVSS.n6877 0.0119575
R33380 DVSS.n6895 DVSS.n6869 0.0119575
R33381 DVSS.n6896 DVSS.n6876 0.0119575
R33382 DVSS.n6908 DVSS.n6870 0.0119575
R33383 DVSS.n6907 DVSS.n6875 0.0119575
R33384 DVSS.n6909 DVSS.n6871 0.0119575
R33385 DVSS.n6911 DVSS.n6873 0.0119575
R33386 DVSS.n6912 DVSS.n6872 0.0119575
R33387 DVSS.n8624 DVSS.n994 0.0119575
R33388 DVSS.n993 DVSS.n990 0.0119575
R33389 DVSS.n8625 DVSS.n996 0.0119575
R33390 DVSS.n995 DVSS.n989 0.0119575
R33391 DVSS.n8626 DVSS.n998 0.0119575
R33392 DVSS.n997 DVSS.n988 0.0119575
R33393 DVSS.n8627 DVSS.n1000 0.0119575
R33394 DVSS.n999 DVSS.n987 0.0119575
R33395 DVSS.n8628 DVSS.n1002 0.0119575
R33396 DVSS.n1001 DVSS.n986 0.0119575
R33397 DVSS.n8629 DVSS.n1004 0.0119575
R33398 DVSS.n1003 DVSS.n985 0.0119575
R33399 DVSS.n8630 DVSS.n1006 0.0119575
R33400 DVSS.n1005 DVSS.n984 0.0119575
R33401 DVSS.n8631 DVSS.n1008 0.0119575
R33402 DVSS.n1007 DVSS.n983 0.0119575
R33403 DVSS.n8632 DVSS.n1010 0.0119575
R33404 DVSS.n1009 DVSS.n982 0.0119575
R33405 DVSS.n8633 DVSS.n1012 0.0119575
R33406 DVSS.n1011 DVSS.n981 0.0119575
R33407 DVSS.n8637 DVSS.n8635 0.0119575
R33408 DVSS.n8636 DVSS.n980 0.0119575
R33409 DVSS.n8639 DVSS.n976 0.0119575
R33410 DVSS.n8667 DVSS.n8656 0.0119575
R33411 DVSS.n8653 DVSS.n975 0.0119575
R33412 DVSS.n8668 DVSS.n8657 0.0119575
R33413 DVSS.n8652 DVSS.n974 0.0119575
R33414 DVSS.n8669 DVSS.n8658 0.0119575
R33415 DVSS.n8651 DVSS.n973 0.0119575
R33416 DVSS.n8670 DVSS.n8659 0.0119575
R33417 DVSS.n8650 DVSS.n972 0.0119575
R33418 DVSS.n8671 DVSS.n8660 0.0119575
R33419 DVSS.n8649 DVSS.n971 0.0119575
R33420 DVSS.n8672 DVSS.n8661 0.0119575
R33421 DVSS.n8648 DVSS.n970 0.0119575
R33422 DVSS.n8673 DVSS.n8662 0.0119575
R33423 DVSS.n8647 DVSS.n969 0.0119575
R33424 DVSS.n8674 DVSS.n8663 0.0119575
R33425 DVSS.n8646 DVSS.n968 0.0119575
R33426 DVSS.n8675 DVSS.n8664 0.0119575
R33427 DVSS.n8645 DVSS.n967 0.0119575
R33428 DVSS.n8676 DVSS.n8665 0.0119575
R33429 DVSS.n8644 DVSS.n966 0.0119575
R33430 DVSS.n8679 DVSS.n8678 0.0119575
R33431 DVSS.n8643 DVSS.n965 0.0119575
R33432 DVSS.n8681 DVSS.n8641 0.0119575
R33433 DVSS.n4488 DVSS.n4455 0.0119575
R33434 DVSS.n4487 DVSS.n4456 0.0119575
R33435 DVSS.n4486 DVSS.n4485 0.0119575
R33436 DVSS.n4484 DVSS.n4457 0.0119575
R33437 DVSS.n4483 DVSS.n4482 0.0119575
R33438 DVSS.n4452 DVSS.n3836 0.0119575
R33439 DVSS.n3846 DVSS.n3844 0.0119575
R33440 DVSS.n3855 DVSS.n3847 0.0119575
R33441 DVSS.n3848 DVSS.n3843 0.0119575
R33442 DVSS.n3854 DVSS.n3849 0.0119575
R33443 DVSS.n3850 DVSS.n3842 0.0119575
R33444 DVSS.n3033 DVSS.n3023 0.0119575
R33445 DVSS.n5856 DVSS.n3034 0.0119575
R33446 DVSS.n5858 DVSS.n5857 0.0119575
R33447 DVSS.n5859 DVSS.n3032 0.0119575
R33448 DVSS.n5861 DVSS.n5860 0.0119575
R33449 DVSS.n5862 DVSS.n3031 0.0119575
R33450 DVSS.n3005 DVSS.n3004 0.0119575
R33451 DVSS.n3006 DVSS.n3002 0.0119575
R33452 DVSS.n3008 DVSS.n3007 0.0119575
R33453 DVSS.n3009 DVSS.n3001 0.0119575
R33454 DVSS.n3011 DVSS.n3010 0.0119575
R33455 DVSS.n2544 DVSS.n2542 0.0119575
R33456 DVSS.n2546 DVSS.n2545 0.0119575
R33457 DVSS.n2547 DVSS.n2541 0.0119575
R33458 DVSS.n2549 DVSS.n2548 0.0119575
R33459 DVSS.n2550 DVSS.n2540 0.0119575
R33460 DVSS.n2552 DVSS.n2551 0.0119575
R33461 DVSS.n2553 DVSS.n2539 0.0119575
R33462 DVSS.n2555 DVSS.n2554 0.0119575
R33463 DVSS.n2556 DVSS.n2538 0.0119575
R33464 DVSS.n2558 DVSS.n2557 0.0119575
R33465 DVSS.n2559 DVSS.n2537 0.0119575
R33466 DVSS.n2561 DVSS.n2560 0.0119575
R33467 DVSS.n2562 DVSS.n2536 0.0119575
R33468 DVSS.n2564 DVSS.n2563 0.0119575
R33469 DVSS.n2565 DVSS.n2535 0.0119575
R33470 DVSS.n2567 DVSS.n2566 0.0119575
R33471 DVSS.n2568 DVSS.n2534 0.0119575
R33472 DVSS.n2570 DVSS.n2569 0.0119575
R33473 DVSS.n2571 DVSS.n2533 0.0119575
R33474 DVSS.n2573 DVSS.n2572 0.0119575
R33475 DVSS.n2574 DVSS.n2532 0.0119575
R33476 DVSS.n2576 DVSS.n2575 0.0119575
R33477 DVSS.n2577 DVSS.n2531 0.0119575
R33478 DVSS.n1927 DVSS.n1926 0.0119575
R33479 DVSS.n8053 DVSS.n1924 0.0119575
R33480 DVSS.n1929 DVSS.n1928 0.0119575
R33481 DVSS.n8054 DVSS.n1923 0.0119575
R33482 DVSS.n1931 DVSS.n1930 0.0119575
R33483 DVSS.n8055 DVSS.n1922 0.0119575
R33484 DVSS.n1933 DVSS.n1932 0.0119575
R33485 DVSS.n8057 DVSS.n1921 0.0119575
R33486 DVSS.n8059 DVSS.n8058 0.0119575
R33487 DVSS.n1920 DVSS.n1916 0.0119575
R33488 DVSS.n6755 DVSS.n6754 0.0119575
R33489 DVSS.n6851 DVSS.n6743 0.0119575
R33490 DVSS.n6757 DVSS.n6756 0.0119575
R33491 DVSS.n6852 DVSS.n6742 0.0119575
R33492 DVSS.n6759 DVSS.n6758 0.0119575
R33493 DVSS.n6853 DVSS.n6741 0.0119575
R33494 DVSS.n6761 DVSS.n6760 0.0119575
R33495 DVSS.n6855 DVSS.n6740 0.0119575
R33496 DVSS.n6857 DVSS.n6856 0.0119575
R33497 DVSS.n6739 DVSS.n6735 0.0119575
R33498 DVSS.n4458 DVSS.n3835 0.0119575
R33499 DVSS.n6887 DVSS.n6860 0.0119575
R33500 DVSS.n6904 DVSS.n6861 0.0119575
R33501 DVSS.n6884 DVSS.n6862 0.0119575
R33502 DVSS.n6903 DVSS.n6888 0.0119575
R33503 DVSS.n6883 DVSS.n6863 0.0119575
R33504 DVSS.n6902 DVSS.n6889 0.0119575
R33505 DVSS.n6882 DVSS.n6864 0.0119575
R33506 DVSS.n6901 DVSS.n6890 0.0119575
R33507 DVSS.n6881 DVSS.n6865 0.0119575
R33508 DVSS.n6900 DVSS.n6891 0.0119575
R33509 DVSS.n6880 DVSS.n6866 0.0119575
R33510 DVSS.n6899 DVSS.n6892 0.0119575
R33511 DVSS.n6879 DVSS.n6867 0.0119575
R33512 DVSS.n6898 DVSS.n6893 0.0119575
R33513 DVSS.n6878 DVSS.n6868 0.0119575
R33514 DVSS.n6897 DVSS.n6894 0.0119575
R33515 DVSS.n6877 DVSS.n6869 0.0119575
R33516 DVSS.n6896 DVSS.n6895 0.0119575
R33517 DVSS.n6876 DVSS.n6870 0.0119575
R33518 DVSS.n6908 DVSS.n6907 0.0119575
R33519 DVSS.n6875 DVSS.n6871 0.0119575
R33520 DVSS.n6909 DVSS.n6873 0.0119575
R33521 DVSS.n6912 DVSS.n6911 0.0119575
R33522 DVSS.n7060 DVSS.n6690 0.0119575
R33523 DVSS.n6706 DVSS.n6705 0.0119575
R33524 DVSS.n7046 DVSS.n6703 0.0119575
R33525 DVSS.n6708 DVSS.n6707 0.0119575
R33526 DVSS.n7047 DVSS.n6702 0.0119575
R33527 DVSS.n6710 DVSS.n6709 0.0119575
R33528 DVSS.n7048 DVSS.n6701 0.0119575
R33529 DVSS.n6712 DVSS.n6711 0.0119575
R33530 DVSS.n7049 DVSS.n6700 0.0119575
R33531 DVSS.n6714 DVSS.n6713 0.0119575
R33532 DVSS.n7050 DVSS.n6699 0.0119575
R33533 DVSS.n6716 DVSS.n6715 0.0119575
R33534 DVSS.n7051 DVSS.n6698 0.0119575
R33535 DVSS.n6718 DVSS.n6717 0.0119575
R33536 DVSS.n7052 DVSS.n6697 0.0119575
R33537 DVSS.n6720 DVSS.n6719 0.0119575
R33538 DVSS.n7053 DVSS.n6696 0.0119575
R33539 DVSS.n6722 DVSS.n6721 0.0119575
R33540 DVSS.n7054 DVSS.n6695 0.0119575
R33541 DVSS.n6724 DVSS.n6723 0.0119575
R33542 DVSS.n7056 DVSS.n6694 0.0119575
R33543 DVSS.n7058 DVSS.n7057 0.0119575
R33544 DVSS.n1316 DVSS.n1189 0.0119575
R33545 DVSS.n1205 DVSS.n1204 0.0119575
R33546 DVSS.n1304 DVSS.n1200 0.0119575
R33547 DVSS.n1207 DVSS.n1206 0.0119575
R33548 DVSS.n1305 DVSS.n1199 0.0119575
R33549 DVSS.n1209 DVSS.n1208 0.0119575
R33550 DVSS.n1306 DVSS.n1198 0.0119575
R33551 DVSS.n1211 DVSS.n1210 0.0119575
R33552 DVSS.n1307 DVSS.n1197 0.0119575
R33553 DVSS.n1213 DVSS.n1212 0.0119575
R33554 DVSS.n1308 DVSS.n1195 0.0119575
R33555 DVSS.n1299 DVSS.n1298 0.0119575
R33556 DVSS.n1309 DVSS.n1194 0.0119575
R33557 DVSS.n1301 DVSS.n1300 0.0119575
R33558 DVSS.n1310 DVSS.n1193 0.0119575
R33559 DVSS.n1303 DVSS.n1302 0.0119575
R33560 DVSS.n1312 DVSS.n1192 0.0119575
R33561 DVSS.n1314 DVSS.n1313 0.0119575
R33562 DVSS.n1077 DVSS.n1073 0.0119575
R33563 DVSS.n8533 DVSS.n1075 0.0119575
R33564 DVSS.n8543 DVSS.n1071 0.0119575
R33565 DVSS.n8544 DVSS.n1070 0.0119575
R33566 DVSS.n8545 DVSS.n8541 0.0119575
R33567 DVSS.n8546 DVSS.n1069 0.0119575
R33568 DVSS.n8547 DVSS.n8540 0.0119575
R33569 DVSS.n8548 DVSS.n1068 0.0119575
R33570 DVSS.n8549 DVSS.n8539 0.0119575
R33571 DVSS.n8550 DVSS.n1067 0.0119575
R33572 DVSS.n8551 DVSS.n1066 0.0119575
R33573 DVSS.n8552 DVSS.n1065 0.0119575
R33574 DVSS.n8553 DVSS.n8537 0.0119575
R33575 DVSS.n8554 DVSS.n1064 0.0119575
R33576 DVSS.n8555 DVSS.n8536 0.0119575
R33577 DVSS.n8556 DVSS.n1063 0.0119575
R33578 DVSS.n8557 DVSS.n8535 0.0119575
R33579 DVSS.n8558 DVSS.n1062 0.0119575
R33580 DVSS.n9635 DVSS.n216 0.0119575
R33581 DVSS.n221 DVSS.n218 0.0119575
R33582 DVSS.n9637 DVSS.n214 0.0119575
R33583 DVSS.n9636 DVSS.n213 0.0119575
R33584 DVSS.n9640 DVSS.n9639 0.0119575
R33585 DVSS.n9638 DVSS.n212 0.0119575
R33586 DVSS.n9643 DVSS.n9642 0.0119575
R33587 DVSS.n9641 DVSS.n211 0.0119575
R33588 DVSS.n9646 DVSS.n9645 0.0119575
R33589 DVSS.n9644 DVSS.n210 0.0119575
R33590 DVSS.n9648 DVSS.n209 0.0119575
R33591 DVSS.n9647 DVSS.n208 0.0119575
R33592 DVSS.n9651 DVSS.n9650 0.0119575
R33593 DVSS.n9649 DVSS.n207 0.0119575
R33594 DVSS.n9654 DVSS.n9653 0.0119575
R33595 DVSS.n9652 DVSS.n206 0.0119575
R33596 DVSS.n9657 DVSS.n9656 0.0119575
R33597 DVSS.n9655 DVSS.n205 0.0119575
R33598 DVSS.n9692 DVSS.n177 0.0119575
R33599 DVSS.n182 DVSS.n179 0.0119575
R33600 DVSS.n9694 DVSS.n175 0.0119575
R33601 DVSS.n9693 DVSS.n174 0.0119575
R33602 DVSS.n9697 DVSS.n9696 0.0119575
R33603 DVSS.n9695 DVSS.n173 0.0119575
R33604 DVSS.n9700 DVSS.n9699 0.0119575
R33605 DVSS.n9698 DVSS.n172 0.0119575
R33606 DVSS.n9703 DVSS.n9702 0.0119575
R33607 DVSS.n9701 DVSS.n171 0.0119575
R33608 DVSS.n9705 DVSS.n170 0.0119575
R33609 DVSS.n9704 DVSS.n169 0.0119575
R33610 DVSS.n9708 DVSS.n9707 0.0119575
R33611 DVSS.n9706 DVSS.n168 0.0119575
R33612 DVSS.n9711 DVSS.n9710 0.0119575
R33613 DVSS.n9709 DVSS.n167 0.0119575
R33614 DVSS.n9714 DVSS.n9713 0.0119575
R33615 DVSS.n9712 DVSS.n166 0.0119575
R33616 DVSS.n9737 DVSS.n155 0.0119575
R33617 DVSS.n9736 DVSS.n154 0.0119575
R33618 DVSS.n9740 DVSS.n9739 0.0119575
R33619 DVSS.n9738 DVSS.n153 0.0119575
R33620 DVSS.n9743 DVSS.n9742 0.0119575
R33621 DVSS.n9741 DVSS.n152 0.0119575
R33622 DVSS.n9746 DVSS.n9745 0.0119575
R33623 DVSS.n9744 DVSS.n151 0.0119575
R33624 DVSS.n9749 DVSS.n9748 0.0119575
R33625 DVSS.n9747 DVSS.n150 0.0119575
R33626 DVSS.n9752 DVSS.n9751 0.0119575
R33627 DVSS.n9750 DVSS.n149 0.0119575
R33628 DVSS.n9755 DVSS.n9754 0.0119575
R33629 DVSS.n9753 DVSS.n148 0.0119575
R33630 DVSS.n9758 DVSS.n9757 0.0119575
R33631 DVSS.n9756 DVSS.n147 0.0119575
R33632 DVSS.n9761 DVSS.n9760 0.0119575
R33633 DVSS.n9759 DVSS.n146 0.0119575
R33634 DVSS.n9764 DVSS.n9763 0.0119575
R33635 DVSS.n9762 DVSS.n145 0.0119575
R33636 DVSS.n9767 DVSS.n9766 0.0119575
R33637 DVSS.n9765 DVSS.n144 0.0119575
R33638 DVSS.n9789 DVSS.n112 0.0119575
R33639 DVSS.n115 DVSS.n114 0.0119575
R33640 DVSS.n9790 DVSS.n111 0.0119575
R33641 DVSS.n117 DVSS.n116 0.0119575
R33642 DVSS.n9791 DVSS.n110 0.0119575
R33643 DVSS.n119 DVSS.n118 0.0119575
R33644 DVSS.n9792 DVSS.n109 0.0119575
R33645 DVSS.n121 DVSS.n120 0.0119575
R33646 DVSS.n9793 DVSS.n108 0.0119575
R33647 DVSS.n123 DVSS.n122 0.0119575
R33648 DVSS.n9794 DVSS.n107 0.0119575
R33649 DVSS.n125 DVSS.n124 0.0119575
R33650 DVSS.n9795 DVSS.n106 0.0119575
R33651 DVSS.n127 DVSS.n126 0.0119575
R33652 DVSS.n9796 DVSS.n105 0.0119575
R33653 DVSS.n129 DVSS.n128 0.0119575
R33654 DVSS.n9797 DVSS.n104 0.0119575
R33655 DVSS.n131 DVSS.n130 0.0119575
R33656 DVSS.n9798 DVSS.n103 0.0119575
R33657 DVSS.n133 DVSS.n132 0.0119575
R33658 DVSS.n9800 DVSS.n102 0.0119575
R33659 DVSS.n9802 DVSS.n9801 0.0119575
R33660 DVSS.n101 DVSS.n97 0.0119575
R33661 DVSS.n8624 DVSS.n991 0.0119575
R33662 DVSS.n994 DVSS.n993 0.0119575
R33663 DVSS.n8625 DVSS.n990 0.0119575
R33664 DVSS.n996 DVSS.n995 0.0119575
R33665 DVSS.n8626 DVSS.n989 0.0119575
R33666 DVSS.n998 DVSS.n997 0.0119575
R33667 DVSS.n8627 DVSS.n988 0.0119575
R33668 DVSS.n1000 DVSS.n999 0.0119575
R33669 DVSS.n8628 DVSS.n987 0.0119575
R33670 DVSS.n1002 DVSS.n1001 0.0119575
R33671 DVSS.n8629 DVSS.n986 0.0119575
R33672 DVSS.n1004 DVSS.n1003 0.0119575
R33673 DVSS.n8630 DVSS.n985 0.0119575
R33674 DVSS.n1006 DVSS.n1005 0.0119575
R33675 DVSS.n8631 DVSS.n984 0.0119575
R33676 DVSS.n1008 DVSS.n1007 0.0119575
R33677 DVSS.n8632 DVSS.n983 0.0119575
R33678 DVSS.n1010 DVSS.n1009 0.0119575
R33679 DVSS.n8633 DVSS.n982 0.0119575
R33680 DVSS.n1012 DVSS.n1011 0.0119575
R33681 DVSS.n8635 DVSS.n981 0.0119575
R33682 DVSS.n8637 DVSS.n8636 0.0119575
R33683 DVSS.n980 DVSS.n976 0.0119575
R33684 DVSS.n7027 DVSS.n6942 0.0119575
R33685 DVSS.n6966 DVSS.n6944 0.0119575
R33686 DVSS.n6969 DVSS.n6941 0.0119575
R33687 DVSS.n6965 DVSS.n6945 0.0119575
R33688 DVSS.n6970 DVSS.n6940 0.0119575
R33689 DVSS.n6964 DVSS.n6946 0.0119575
R33690 DVSS.n6971 DVSS.n6939 0.0119575
R33691 DVSS.n6963 DVSS.n6947 0.0119575
R33692 DVSS.n6972 DVSS.n6938 0.0119575
R33693 DVSS.n6962 DVSS.n6948 0.0119575
R33694 DVSS.n6973 DVSS.n6937 0.0119575
R33695 DVSS.n6961 DVSS.n6949 0.0119575
R33696 DVSS.n6974 DVSS.n6936 0.0119575
R33697 DVSS.n6960 DVSS.n6950 0.0119575
R33698 DVSS.n6975 DVSS.n6935 0.0119575
R33699 DVSS.n6959 DVSS.n6951 0.0119575
R33700 DVSS.n6976 DVSS.n6934 0.0119575
R33701 DVSS.n6958 DVSS.n6952 0.0119575
R33702 DVSS.n6977 DVSS.n6933 0.0119575
R33703 DVSS.n6957 DVSS.n6953 0.0119575
R33704 DVSS.n6978 DVSS.n6932 0.0119575
R33705 DVSS.n6956 DVSS.n6954 0.0119575
R33706 DVSS.n6955 DVSS.n6931 0.0119575
R33707 DVSS.n8860 DVSS.n806 0.0119575
R33708 DVSS.n8835 DVSS.n811 0.0119575
R33709 DVSS.n8836 DVSS.n812 0.0119575
R33710 DVSS.n8838 DVSS.n8837 0.0119575
R33711 DVSS.n8834 DVSS.n813 0.0119575
R33712 DVSS.n8840 DVSS.n8839 0.0119575
R33713 DVSS.n8833 DVSS.n814 0.0119575
R33714 DVSS.n8842 DVSS.n8841 0.0119575
R33715 DVSS.n8832 DVSS.n815 0.0119575
R33716 DVSS.n8844 DVSS.n8843 0.0119575
R33717 DVSS.n8831 DVSS.n816 0.0119575
R33718 DVSS.n8846 DVSS.n8845 0.0119575
R33719 DVSS.n8830 DVSS.n817 0.0119575
R33720 DVSS.n8848 DVSS.n8847 0.0119575
R33721 DVSS.n8829 DVSS.n818 0.0119575
R33722 DVSS.n8850 DVSS.n8849 0.0119575
R33723 DVSS.n8828 DVSS.n819 0.0119575
R33724 DVSS.n8852 DVSS.n8851 0.0119575
R33725 DVSS.n8827 DVSS.n820 0.0119575
R33726 DVSS.n8854 DVSS.n8853 0.0119575
R33727 DVSS.n8826 DVSS.n821 0.0119575
R33728 DVSS.n8855 DVSS.n823 0.0119575
R33729 DVSS.n8858 DVSS.n8857 0.0119575
R33730 DVSS.n422 DVSS.n421 0.0119575
R33731 DVSS.n424 DVSS.n423 0.0119575
R33732 DVSS.n444 DVSS.n420 0.0119575
R33733 DVSS.n426 DVSS.n425 0.0119575
R33734 DVSS.n445 DVSS.n419 0.0119575
R33735 DVSS.n428 DVSS.n427 0.0119575
R33736 DVSS.n446 DVSS.n418 0.0119575
R33737 DVSS.n430 DVSS.n429 0.0119575
R33738 DVSS.n447 DVSS.n417 0.0119575
R33739 DVSS.n432 DVSS.n431 0.0119575
R33740 DVSS.n448 DVSS.n416 0.0119575
R33741 DVSS.n434 DVSS.n433 0.0119575
R33742 DVSS.n449 DVSS.n415 0.0119575
R33743 DVSS.n436 DVSS.n435 0.0119575
R33744 DVSS.n450 DVSS.n414 0.0119575
R33745 DVSS.n438 DVSS.n437 0.0119575
R33746 DVSS.n451 DVSS.n413 0.0119575
R33747 DVSS.n440 DVSS.n439 0.0119575
R33748 DVSS.n452 DVSS.n412 0.0119575
R33749 DVSS.n442 DVSS.n441 0.0119575
R33750 DVSS.n454 DVSS.n411 0.0119575
R33751 DVSS.n456 DVSS.n455 0.0119575
R33752 DVSS.n410 DVSS.n406 0.0119575
R33753 DVSS.n272 DVSS.n268 0.0119575
R33754 DVSS.n9575 DVSS.n273 0.0119575
R33755 DVSS.n9558 DVSS.n274 0.0119575
R33756 DVSS.n9574 DVSS.n9559 0.0119575
R33757 DVSS.n9557 DVSS.n275 0.0119575
R33758 DVSS.n9573 DVSS.n9560 0.0119575
R33759 DVSS.n9556 DVSS.n276 0.0119575
R33760 DVSS.n9572 DVSS.n9561 0.0119575
R33761 DVSS.n9555 DVSS.n277 0.0119575
R33762 DVSS.n9571 DVSS.n9562 0.0119575
R33763 DVSS.n9554 DVSS.n278 0.0119575
R33764 DVSS.n9570 DVSS.n9563 0.0119575
R33765 DVSS.n9553 DVSS.n279 0.0119575
R33766 DVSS.n9569 DVSS.n9564 0.0119575
R33767 DVSS.n9552 DVSS.n280 0.0119575
R33768 DVSS.n9568 DVSS.n9565 0.0119575
R33769 DVSS.n9551 DVSS.n281 0.0119575
R33770 DVSS.n9567 DVSS.n9566 0.0119575
R33771 DVSS.n9550 DVSS.n282 0.0119575
R33772 DVSS.n9578 DVSS.n9577 0.0119575
R33773 DVSS.n9549 DVSS.n283 0.0119575
R33774 DVSS.n9579 DVSS.n9547 0.0119575
R33775 DVSS.n9582 DVSS.n9581 0.0119575
R33776 DVSS.n9828 DVSS.n9805 0.0119575
R33777 DVSS.n9807 DVSS.n9806 0.0119575
R33778 DVSS.n9829 DVSS.n96 0.0119575
R33779 DVSS.n9809 DVSS.n9808 0.0119575
R33780 DVSS.n9830 DVSS.n95 0.0119575
R33781 DVSS.n9811 DVSS.n9810 0.0119575
R33782 DVSS.n9831 DVSS.n94 0.0119575
R33783 DVSS.n9813 DVSS.n9812 0.0119575
R33784 DVSS.n9832 DVSS.n93 0.0119575
R33785 DVSS.n9815 DVSS.n9814 0.0119575
R33786 DVSS.n9833 DVSS.n92 0.0119575
R33787 DVSS.n9817 DVSS.n9816 0.0119575
R33788 DVSS.n9834 DVSS.n91 0.0119575
R33789 DVSS.n9819 DVSS.n9818 0.0119575
R33790 DVSS.n9835 DVSS.n90 0.0119575
R33791 DVSS.n9821 DVSS.n9820 0.0119575
R33792 DVSS.n9836 DVSS.n89 0.0119575
R33793 DVSS.n9823 DVSS.n9822 0.0119575
R33794 DVSS.n9837 DVSS.n88 0.0119575
R33795 DVSS.n9825 DVSS.n9824 0.0119575
R33796 DVSS.n9838 DVSS.n87 0.0119575
R33797 DVSS.n9827 DVSS.n9826 0.0119575
R33798 DVSS.n9840 DVSS.n86 0.0119575
R33799 DVSS.n8667 DVSS.n8640 0.0119575
R33800 DVSS.n8656 DVSS.n975 0.0119575
R33801 DVSS.n8668 DVSS.n8653 0.0119575
R33802 DVSS.n8657 DVSS.n974 0.0119575
R33803 DVSS.n8669 DVSS.n8652 0.0119575
R33804 DVSS.n8658 DVSS.n973 0.0119575
R33805 DVSS.n8670 DVSS.n8651 0.0119575
R33806 DVSS.n8659 DVSS.n972 0.0119575
R33807 DVSS.n8671 DVSS.n8650 0.0119575
R33808 DVSS.n8660 DVSS.n971 0.0119575
R33809 DVSS.n8672 DVSS.n8649 0.0119575
R33810 DVSS.n8661 DVSS.n970 0.0119575
R33811 DVSS.n8673 DVSS.n8648 0.0119575
R33812 DVSS.n8662 DVSS.n969 0.0119575
R33813 DVSS.n8674 DVSS.n8647 0.0119575
R33814 DVSS.n8663 DVSS.n968 0.0119575
R33815 DVSS.n8675 DVSS.n8646 0.0119575
R33816 DVSS.n8664 DVSS.n967 0.0119575
R33817 DVSS.n8676 DVSS.n8645 0.0119575
R33818 DVSS.n8665 DVSS.n966 0.0119575
R33819 DVSS.n8678 DVSS.n8644 0.0119575
R33820 DVSS.n8679 DVSS.n965 0.0119575
R33821 DVSS.n8643 DVSS.n8641 0.0119575
R33822 DVSS.n917 DVSS.n915 0.0119575
R33823 DVSS.n919 DVSS.n918 0.0119575
R33824 DVSS.n920 DVSS.n914 0.0119575
R33825 DVSS.n922 DVSS.n921 0.0119575
R33826 DVSS.n923 DVSS.n913 0.0119575
R33827 DVSS.n925 DVSS.n924 0.0119575
R33828 DVSS.n926 DVSS.n912 0.0119575
R33829 DVSS.n928 DVSS.n927 0.0119575
R33830 DVSS.n929 DVSS.n911 0.0119575
R33831 DVSS.n931 DVSS.n930 0.0119575
R33832 DVSS.n932 DVSS.n910 0.0119575
R33833 DVSS.n934 DVSS.n933 0.0119575
R33834 DVSS.n935 DVSS.n909 0.0119575
R33835 DVSS.n937 DVSS.n936 0.0119575
R33836 DVSS.n938 DVSS.n908 0.0119575
R33837 DVSS.n940 DVSS.n939 0.0119575
R33838 DVSS.n941 DVSS.n907 0.0119575
R33839 DVSS.n943 DVSS.n942 0.0119575
R33840 DVSS.n944 DVSS.n906 0.0119575
R33841 DVSS.n946 DVSS.n945 0.0119575
R33842 DVSS.n947 DVSS.n905 0.0119575
R33843 DVSS.n8716 DVSS.n948 0.0119575
R33844 DVSS.n904 DVSS.n903 0.0119575
R33845 DVSS.n854 DVSS.n852 0.0119575
R33846 DVSS.n856 DVSS.n855 0.0119575
R33847 DVSS.n857 DVSS.n851 0.0119575
R33848 DVSS.n859 DVSS.n858 0.0119575
R33849 DVSS.n860 DVSS.n850 0.0119575
R33850 DVSS.n862 DVSS.n861 0.0119575
R33851 DVSS.n863 DVSS.n849 0.0119575
R33852 DVSS.n865 DVSS.n864 0.0119575
R33853 DVSS.n866 DVSS.n848 0.0119575
R33854 DVSS.n868 DVSS.n867 0.0119575
R33855 DVSS.n869 DVSS.n847 0.0119575
R33856 DVSS.n871 DVSS.n870 0.0119575
R33857 DVSS.n872 DVSS.n846 0.0119575
R33858 DVSS.n874 DVSS.n873 0.0119575
R33859 DVSS.n875 DVSS.n845 0.0119575
R33860 DVSS.n877 DVSS.n876 0.0119575
R33861 DVSS.n878 DVSS.n844 0.0119575
R33862 DVSS.n880 DVSS.n879 0.0119575
R33863 DVSS.n881 DVSS.n843 0.0119575
R33864 DVSS.n883 DVSS.n882 0.0119575
R33865 DVSS.n884 DVSS.n842 0.0119575
R33866 DVSS.n8751 DVSS.n885 0.0119575
R33867 DVSS.n841 DVSS.n840 0.0119575
R33868 DVSS.n9353 DVSS.n459 0.0119575
R33869 DVSS.n462 DVSS.n461 0.0119575
R33870 DVSS.n9354 DVSS.n405 0.0119575
R33871 DVSS.n464 DVSS.n463 0.0119575
R33872 DVSS.n9355 DVSS.n404 0.0119575
R33873 DVSS.n466 DVSS.n465 0.0119575
R33874 DVSS.n9356 DVSS.n403 0.0119575
R33875 DVSS.n468 DVSS.n467 0.0119575
R33876 DVSS.n9357 DVSS.n402 0.0119575
R33877 DVSS.n470 DVSS.n469 0.0119575
R33878 DVSS.n9358 DVSS.n401 0.0119575
R33879 DVSS.n472 DVSS.n471 0.0119575
R33880 DVSS.n9359 DVSS.n400 0.0119575
R33881 DVSS.n474 DVSS.n473 0.0119575
R33882 DVSS.n9360 DVSS.n399 0.0119575
R33883 DVSS.n476 DVSS.n475 0.0119575
R33884 DVSS.n9361 DVSS.n398 0.0119575
R33885 DVSS.n478 DVSS.n477 0.0119575
R33886 DVSS.n9362 DVSS.n397 0.0119575
R33887 DVSS.n480 DVSS.n479 0.0119575
R33888 DVSS.n9364 DVSS.n396 0.0119575
R33889 DVSS.n9366 DVSS.n9365 0.0119575
R33890 DVSS.n395 DVSS.n391 0.0119575
R33891 DVSS.n9545 DVSS.n284 0.0119575
R33892 DVSS.n302 DVSS.n301 0.0119575
R33893 DVSS.n9314 DVSS.n299 0.0119575
R33894 DVSS.n304 DVSS.n303 0.0119575
R33895 DVSS.n9315 DVSS.n298 0.0119575
R33896 DVSS.n306 DVSS.n305 0.0119575
R33897 DVSS.n9316 DVSS.n297 0.0119575
R33898 DVSS.n308 DVSS.n307 0.0119575
R33899 DVSS.n9317 DVSS.n296 0.0119575
R33900 DVSS.n310 DVSS.n309 0.0119575
R33901 DVSS.n9318 DVSS.n295 0.0119575
R33902 DVSS.n312 DVSS.n311 0.0119575
R33903 DVSS.n9319 DVSS.n294 0.0119575
R33904 DVSS.n314 DVSS.n313 0.0119575
R33905 DVSS.n9320 DVSS.n293 0.0119575
R33906 DVSS.n316 DVSS.n315 0.0119575
R33907 DVSS.n9321 DVSS.n292 0.0119575
R33908 DVSS.n318 DVSS.n317 0.0119575
R33909 DVSS.n9322 DVSS.n291 0.0119575
R33910 DVSS.n320 DVSS.n319 0.0119575
R33911 DVSS.n9323 DVSS.n290 0.0119575
R33912 DVSS.n322 DVSS.n321 0.0119575
R33913 DVSS.n323 DVSS.n289 0.0119575
R33914 DVSS.n9919 DVSS.n17 0.0119575
R33915 DVSS.n9909 DVSS.n16 0.0119575
R33916 DVSS.n9920 DVSS.n9908 0.0119575
R33917 DVSS.n9910 DVSS.n15 0.0119575
R33918 DVSS.n9921 DVSS.n9907 0.0119575
R33919 DVSS.n9911 DVSS.n14 0.0119575
R33920 DVSS.n9922 DVSS.n9906 0.0119575
R33921 DVSS.n9912 DVSS.n13 0.0119575
R33922 DVSS.n9923 DVSS.n9905 0.0119575
R33923 DVSS.n9913 DVSS.n12 0.0119575
R33924 DVSS.n9924 DVSS.n9904 0.0119575
R33925 DVSS.n9914 DVSS.n11 0.0119575
R33926 DVSS.n9925 DVSS.n9903 0.0119575
R33927 DVSS.n9915 DVSS.n10 0.0119575
R33928 DVSS.n9926 DVSS.n9902 0.0119575
R33929 DVSS.n9916 DVSS.n9 0.0119575
R33930 DVSS.n9927 DVSS.n9901 0.0119575
R33931 DVSS.n9917 DVSS.n8 0.0119575
R33932 DVSS.n9928 DVSS.n9900 0.0119575
R33933 DVSS.n9918 DVSS.n7 0.0119575
R33934 DVSS.n9930 DVSS.n9899 0.0119575
R33935 DVSS.n9931 DVSS.n6 0.0119575
R33936 DVSS.n9898 DVSS.n18 0.0119575
R33937 DVSS.n4621 DVSS.n2761 0.0116972
R33938 DVSS.n3984 DVSS.n3476 0.0116972
R33939 DVSS.n5022 DVSS.n5019 0.0116972
R33940 DVSS.n5028 DVSS.n5013 0.0116972
R33941 DVSS.n5024 DVSS.n5020 0.0116972
R33942 DVSS.n5026 DVSS.n5012 0.0116972
R33943 DVSS.n5195 DVSS.n5030 0.0116972
R33944 DVSS.n4602 DVSS.n3774 0.0116972
R33945 DVSS.n3989 DVSS.n3972 0.0116972
R33946 DVSS.n3520 DVSS.n3186 0.0116972
R33947 DVSS.n3559 DVSS.n3177 0.0116972
R33948 DVSS.n3522 DVSS.n3187 0.0116972
R33949 DVSS.n3556 DVSS.n3176 0.0116972
R33950 DVSS.n5740 DVSS.n3188 0.0116972
R33951 DVSS.n8919 DVSS.n778 0.0116614
R33952 DVSS.n8954 DVSS.n735 0.0116614
R33953 DVSS.n9453 DVSS.n362 0.0116614
R33954 DVSS.n9488 DVSS.n34 0.0116614
R33955 DVSS.n4625 DVSS.n4623 0.0114859
R33956 DVSS.n4699 DVSS.n3777 0.0114859
R33957 DVSS.n8885 DVSS.n783 0.0113607
R33958 DVSS.n9415 DVSS.n9414 0.0113607
R33959 DVSS.n8883 DVSS.n783 0.0113607
R33960 DVSS.n9414 DVSS.n365 0.0113607
R33961 DVSS.n8919 DVSS.n762 0.0113071
R33962 DVSS.n8954 DVSS.n740 0.0113071
R33963 DVSS.n9453 DVSS.n347 0.0113071
R33964 DVSS.n9488 DVSS.n38 0.0113071
R33965 DVSS.n4816 DVSS.n3668 0.0112746
R33966 DVSS.n4822 DVSS.n3672 0.0112746
R33967 DVSS.n3674 DVSS.n3671 0.0112746
R33968 DVSS.n4819 DVSS.n3676 0.0112746
R33969 DVSS.n4818 DVSS.n3670 0.0112746
R33970 DVSS.n5198 DVSS.n5008 0.0112746
R33971 DVSS.n5568 DVSS.n2300 0.0112746
R33972 DVSS.n9382 DVSS.n386 0.0112746
R33973 DVSS.n3706 DVSS.n3700 0.0112746
R33974 DVSS.n4805 DVSS.n3693 0.0112746
R33975 DVSS.n3708 DVSS.n3701 0.0112746
R33976 DVSS.n3702 DVSS.n3692 0.0112746
R33977 DVSS.n4808 DVSS.n4807 0.0112746
R33978 DVSS.n3519 DVSS.n3179 0.0112746
R33979 DVSS.n5590 DVSS.n2330 0.0112746
R33980 DVSS.n9025 DVSS.n9024 0.0112746
R33981 DVSS.n8903 DVSS.n765 0.0109528
R33982 DVSS.n9437 DVSS.n350 0.0109528
R33983 DVSS.n9476 DVSS.n336 0.0108846
R33984 DVSS.n9479 DVSS.n336 0.0108846
R33985 DVSS.n8942 DVSS.n751 0.0108846
R33986 DVSS.n8945 DVSS.n751 0.0108846
R33987 DVSS.n5554 DVSS.n2291 0.0108521
R33988 DVSS.n7900 DVSS.n2073 0.0108521
R33989 DVSS.n9394 DVSS.n375 0.0108521
R33990 DVSS.n5619 DVSS.n2321 0.0108521
R33991 DVSS.n7894 DVSS.n2055 0.0108521
R33992 DVSS.n9129 DVSS.n603 0.0108521
R33993 DVSS.n4442 DVSS.n4441 0.0107778
R33994 DVSS.n4933 DVSS.n3593 0.0107778
R33995 DVSS.n5867 DVSS.n3025 0.0107778
R33996 DVSS.n5918 DVSS.n2920 0.0107778
R33997 DVSS.n3537 DVSS.n3015 0.0107778
R33998 DVSS.n5379 DVSS.n5378 0.0107778
R33999 DVSS.n5672 DVSS.n2991 0.0107778
R34000 DVSS.n5909 DVSS.n2962 0.0107778
R34001 DVSS.n5893 DVSS.n2987 0.0107778
R34002 DVSS.n5904 DVSS.n2971 0.0107778
R34003 DVSS.n7373 DVSS.n2582 0.0107778
R34004 DVSS.n7696 DVSS.n2116 0.0107778
R34005 DVSS.n7368 DVSS.n7362 0.0107778
R34006 DVSS.n7709 DVSS.n7708 0.0107778
R34007 DVSS.n8070 DVSS.n8069 0.0107778
R34008 DVSS.n8181 DVSS.n1758 0.0107778
R34009 DVSS.n3579 DVSS.n3412 0.0105984
R34010 DVSS.n4993 DVSS.n3410 0.0105984
R34011 DVSS.n3582 DVSS.n3413 0.0105984
R34012 DVSS.n3586 DVSS.n3409 0.0105984
R34013 DVSS.n3581 DVSS.n3415 0.0105984
R34014 DVSS.n3569 DVSS.n3447 0.0105984
R34015 DVSS.n4997 DVSS.n3445 0.0105984
R34016 DVSS.n3572 DVSS.n3448 0.0105984
R34017 DVSS.n3576 DVSS.n3444 0.0105984
R34018 DVSS.n3571 DVSS.n3450 0.0105984
R34019 DVSS.n3999 DVSS.n3937 0.0105984
R34020 DVSS.n4009 DVSS.n3935 0.0105984
R34021 DVSS.n4002 DVSS.n3938 0.0105984
R34022 DVSS.n4005 DVSS.n3934 0.0105984
R34023 DVSS.n4001 DVSS.n3939 0.0105984
R34024 DVSS.n4190 DVSS.n3879 0.0105984
R34025 DVSS.n4188 DVSS.n4187 0.0105984
R34026 DVSS.n4175 DVSS.n3886 0.0105984
R34027 DVSS.n4174 DVSS.n3894 0.0105984
R34028 DVSS.n4177 DVSS.n3885 0.0105984
R34029 DVSS.n8936 DVSS.n8935 0.0105984
R34030 DVSS.n8970 DVSS.n732 0.0105984
R34031 DVSS.n4980 DVSS.n3387 0.0105984
R34032 DVSS.n4990 DVSS.n3385 0.0105984
R34033 DVSS.n4983 DVSS.n3388 0.0105984
R34034 DVSS.n4987 DVSS.n3384 0.0105984
R34035 DVSS.n4982 DVSS.n3390 0.0105984
R34036 DVSS.n9470 DVSS.n9469 0.0105984
R34037 DVSS.n9504 DVSS.n31 0.0105984
R34038 DVSS.n4929 DVSS.n4917 0.0105984
R34039 DVSS.n5916 DVSS.n2916 0.0105984
R34040 DVSS.n4444 DVSS.n3852 0.0105984
R34041 DVSS.n5866 DVSS.n5865 0.0105984
R34042 DVSS.n8202 DVSS.n1541 0.0105466
R34043 DVSS.n8205 DVSS.n1542 0.0105466
R34044 DVSS.n1546 DVSS.n1543 0.0105466
R34045 DVSS.n8495 DVSS.n1099 0.0105466
R34046 DVSS.n8483 DVSS.n1126 0.0105466
R34047 DVSS.n8481 DVSS.n1132 0.0105466
R34048 DVSS.n1255 DVSS.n1249 0.0105466
R34049 DVSS.n8209 DVSS.n1537 0.0105466
R34050 DVSS.n8211 DVSS.n1531 0.0105466
R34051 DVSS.n8216 DVSS.n1530 0.0105466
R34052 DVSS.n1463 DVSS.n1462 0.0105466
R34053 DVSS.n8313 DVSS.n1464 0.0105466
R34054 DVSS.n8268 DVSS.n8263 0.0105466
R34055 DVSS.n8272 DVSS.n8264 0.0105466
R34056 DVSS.n8326 DVSS.n8322 0.0105466
R34057 DVSS.n8328 DVSS.n1445 0.0105466
R34058 DVSS.n8332 DVSS.n8331 0.0105466
R34059 DVSS.n8339 DVSS.n1437 0.0105466
R34060 DVSS.n8353 DVSS.n1419 0.0105466
R34061 DVSS.n1136 DVSS.n1134 0.0105466
R34062 DVSS.n8477 DVSS.n1140 0.0105466
R34063 DVSS.n1248 DVSS.n1242 0.0105466
R34064 DVSS.n8333 DVSS.n8332 0.0105466
R34065 DVSS.n8264 DVSS.n8263 0.0105466
R34066 DVSS.n8268 DVSS.n1465 0.0105466
R34067 DVSS.n8326 DVSS.n1445 0.0105466
R34068 DVSS.n8322 DVSS.n1449 0.0105466
R34069 DVSS.n1464 DVSS.n1463 0.0105466
R34070 DVSS.n1462 DVSS.n1461 0.0105466
R34071 DVSS.n8212 DVSS.n1530 0.0105466
R34072 DVSS.n7153 DVSS.n6651 0.0105466
R34073 DVSS.n7151 DVSS.n6652 0.0105466
R34074 DVSS.n7148 DVSS.n7139 0.0105466
R34075 DVSS.n8236 DVSS.n8232 0.0105466
R34076 DVSS.n8238 DVSS.n1512 0.0105466
R34077 DVSS.n8241 DVSS.n8240 0.0105466
R34078 DVSS.n8248 DVSS.n8242 0.0105466
R34079 DVSS.n1487 DVSS.n1482 0.0105466
R34080 DVSS.n8292 DVSS.n1483 0.0105466
R34081 DVSS.n7118 DVSS.n7078 0.0105466
R34082 DVSS.n7123 DVSS.n7076 0.0105466
R34083 DVSS.n8371 DVSS.n8363 0.0105466
R34084 DVSS.n8442 DVSS.n1321 0.0105466
R34085 DVSS.n8447 DVSS.n1322 0.0105466
R34086 DVSS.n1233 DVSS.n1227 0.0105466
R34087 DVSS.n7150 DVSS.n7139 0.0105466
R34088 DVSS.n7078 DVSS.n1484 0.0105466
R34089 DVSS.n1483 DVSS.n1482 0.0105466
R34090 DVSS.n1490 DVSS.n1487 0.0105466
R34091 DVSS.n8242 DVSS.n8241 0.0105466
R34092 DVSS.n8240 DVSS.n8239 0.0105466
R34093 DVSS.n8236 DVSS.n1512 0.0105466
R34094 DVSS.n8232 DVSS.n1516 0.0105466
R34095 DVSS.n7153 DVSS.n6652 0.0105466
R34096 DVSS.n6651 DVSS.n6650 0.0105466
R34097 DVSS.n8479 DVSS.n1136 0.0105466
R34098 DVSS.n8487 DVSS.n1126 0.0105466
R34099 DVSS.n8483 DVSS.n1132 0.0105466
R34100 DVSS.n1140 DVSS.n1134 0.0105466
R34101 DVSS.n8444 DVSS.n1322 0.0105466
R34102 DVSS.n8444 DVSS.n1321 0.0105466
R34103 DVSS.n1282 DVSS.n1233 0.0105466
R34104 DVSS.n1262 DVSS.n1248 0.0105466
R34105 DVSS.n1257 DVSS.n1255 0.0105466
R34106 DVSS.n8491 DVSS.n1099 0.0105466
R34107 DVSS.n1419 DVSS.n1417 0.0105466
R34108 DVSS.n8367 DVSS.n8363 0.0105466
R34109 DVSS.n7119 DVSS.n7076 0.0105466
R34110 DVSS.n8336 DVSS.n1437 0.0105466
R34111 DVSS.n1550 DVSS.n1543 0.0105466
R34112 DVSS.n7132 DVSS.n6656 0.0105466
R34113 DVSS.n7130 DVSS.n6657 0.0105466
R34114 DVSS.n7127 DVSS.n7072 0.0105466
R34115 DVSS.n8457 DVSS.n1154 0.0105466
R34116 DVSS.n1319 DVSS.n1181 0.0105466
R34117 DVSS.n1317 DVSS.n1187 0.0105466
R34118 DVSS.n1226 DVSS.n1220 0.0105466
R34119 DVSS.n7129 DVSS.n7072 0.0105466
R34120 DVSS.n1154 DVSS.n1152 0.0105466
R34121 DVSS.n8450 DVSS.n1181 0.0105466
R34122 DVSS.n1319 DVSS.n1187 0.0105466
R34123 DVSS.n1287 DVSS.n1226 0.0105466
R34124 DVSS.n7066 DVSS.n6660 0.0105466
R34125 DVSS.n7064 DVSS.n6661 0.0105466
R34126 DVSS.n8882 DVSS.n8881 0.0105466
R34127 DVSS.n786 DVSS.n782 0.0105466
R34128 DVSS.n720 DVSS.n715 0.0105466
R34129 DVSS.n9001 DVSS.n718 0.0105466
R34130 DVSS.n717 DVSS.n716 0.0105466
R34131 DVSS.n8195 DVSS.n1555 0.0105466
R34132 DVSS.n8198 DVSS.n1556 0.0105466
R34133 DVSS.n9418 DVSS.n9416 0.0105466
R34134 DVSS.n9417 DVSS.n366 0.0105466
R34135 DVSS.n334 DVSS.n333 0.0105466
R34136 DVSS.n9536 DVSS.n9535 0.0105466
R34137 DVSS.n335 DVSS.n331 0.0105466
R34138 DVSS.n718 DVSS.n717 0.0105466
R34139 DVSS.n9001 DVSS.n715 0.0105466
R34140 DVSS.n9003 DVSS.n720 0.0105466
R34141 DVSS.n9535 DVSS.n335 0.0105466
R34142 DVSS.n9536 DVSS.n334 0.0105466
R34143 DVSS.n333 DVSS.n51 0.0105466
R34144 DVSS.n8882 DVSS.n782 0.0105466
R34145 DVSS.n8881 DVSS.n8880 0.0105466
R34146 DVSS.n9418 DVSS.n9417 0.0105466
R34147 DVSS.n9416 DVSS.n158 0.0105466
R34148 DVSS.n8209 DVSS.n1531 0.0105466
R34149 DVSS.n1538 DVSS.n1537 0.0105466
R34150 DVSS.n1542 DVSS.n1541 0.0105466
R34151 DVSS.n1556 DVSS.n1555 0.0105466
R34152 DVSS.n8202 DVSS.n8201 0.0105466
R34153 DVSS.n8195 DVSS.n8194 0.0105466
R34154 DVSS.n5910 DVSS.n2961 0.0105466
R34155 DVSS.n2966 DVSS.n2964 0.0105466
R34156 DVSS.n5905 DVSS.n2970 0.0105466
R34157 DVSS.n2975 DVSS.n2973 0.0105466
R34158 DVSS.n7695 DVSS.n2113 0.0105466
R34159 DVSS.n2115 DVSS.n2110 0.0105466
R34160 DVSS.n7707 DVSS.n7706 0.0105466
R34161 DVSS.n7702 DVSS.n2107 0.0105466
R34162 DVSS.n8180 DVSS.n1754 0.0105466
R34163 DVSS.n8182 DVSS.n1757 0.0105466
R34164 DVSS.n8190 DVSS.n8189 0.0105466
R34165 DVSS.n8190 DVSS.n1750 0.0105466
R34166 DVSS.n5906 DVSS.n2964 0.0105466
R34167 DVSS.n2965 DVSS.n2961 0.0105466
R34168 DVSS.n5901 DVSS.n2973 0.0105466
R34169 DVSS.n2974 DVSS.n2970 0.0105466
R34170 DVSS.n7699 DVSS.n2110 0.0105466
R34171 DVSS.n2114 DVSS.n2113 0.0105466
R34172 DVSS.n7704 DVSS.n2107 0.0105466
R34173 DVSS.n7706 DVSS.n7701 0.0105466
R34174 DVSS.n8183 DVSS.n8182 0.0105466
R34175 DVSS.n1759 DVSS.n1754 0.0105466
R34176 DVSS.n7066 DVSS.n6661 0.0105466
R34177 DVSS.n7132 DVSS.n6657 0.0105466
R34178 DVSS.n6660 DVSS.n6659 0.0105466
R34179 DVSS.n6656 DVSS.n6655 0.0105466
R34180 DVSS.n5885 DVSS.n2992 0.0105466
R34181 DVSS.n5887 DVSS.n5886 0.0105466
R34182 DVSS.n5888 DVSS.n5887 0.0105466
R34183 DVSS.n5890 DVSS.n2990 0.0105466
R34184 DVSS.n2986 DVSS.n2981 0.0105466
R34185 DVSS.n2989 DVSS.n2988 0.0105466
R34186 DVSS.n2989 DVSS.n2983 0.0105466
R34187 DVSS.n5894 DVSS.n2984 0.0105466
R34188 DVSS.n7375 DVSS.n7374 0.0105466
R34189 DVSS.n2584 DVSS.n2580 0.0105466
R34190 DVSS.n2584 DVSS.n2583 0.0105466
R34191 DVSS.n7372 DVSS.n2586 0.0105466
R34192 DVSS.n7370 DVSS.n7369 0.0105466
R34193 DVSS.n7364 DVSS.n2589 0.0105466
R34194 DVSS.n7364 DVSS.n7363 0.0105466
R34195 DVSS.n7367 DVSS.n7366 0.0105466
R34196 DVSS.n8063 DVSS.n1910 0.0105466
R34197 DVSS.n8064 DVSS.n1911 0.0105466
R34198 DVSS.n8066 DVSS.n1911 0.0105466
R34199 DVSS.n8068 DVSS.n1913 0.0105466
R34200 DVSS.n6746 DVSS.n1914 0.0105466
R34201 DVSS.n6746 DVSS.n6745 0.0105466
R34202 DVSS.n8064 DVSS.n1910 0.0105466
R34203 DVSS.n8063 DVSS.n8062 0.0105466
R34204 DVSS.n7369 DVSS.n2589 0.0105466
R34205 DVSS.n7371 DVSS.n7370 0.0105466
R34206 DVSS.n7374 DVSS.n2580 0.0105466
R34207 DVSS.n7376 DVSS.n7375 0.0105466
R34208 DVSS.n2988 DVSS.n2986 0.0105466
R34209 DVSS.n5891 DVSS.n2981 0.0105466
R34210 DVSS.n5886 DVSS.n5885 0.0105466
R34211 DVSS.n5881 DVSS.n2992 0.0105466
R34212 DVSS.n5884 DVSS.n2990 0.0105466
R34213 DVSS.n5888 DVSS.n5884 0.0105466
R34214 DVSS.n2985 DVSS.n2984 0.0105466
R34215 DVSS.n2985 DVSS.n2983 0.0105466
R34216 DVSS.n2586 DVSS.n2581 0.0105466
R34217 DVSS.n2583 DVSS.n2581 0.0105466
R34218 DVSS.n7366 DVSS.n2590 0.0105466
R34219 DVSS.n7363 DVSS.n2590 0.0105466
R34220 DVSS.n1913 DVSS.n1909 0.0105466
R34221 DVSS.n8066 DVSS.n1909 0.0105466
R34222 DVSS.n4480 DVSS.n3833 0.0105
R34223 DVSS.n4494 DVSS.n3833 0.0105
R34224 DVSS.n4494 DVSS.n3831 0.0105
R34225 DVSS.n4498 DVSS.n3831 0.0105
R34226 DVSS.n4498 DVSS.n3829 0.0105
R34227 DVSS.n4503 DVSS.n3829 0.0105
R34228 DVSS.n4503 DVSS.n3827 0.0105
R34229 DVSS.n4507 DVSS.n3827 0.0105
R34230 DVSS.n4507 DVSS.n3814 0.0105
R34231 DVSS.n4521 DVSS.n3814 0.0105
R34232 DVSS.n4521 DVSS.n3812 0.0105
R34233 DVSS.n4525 DVSS.n3812 0.0105
R34234 DVSS.n4525 DVSS.n3810 0.0105
R34235 DVSS.n4529 DVSS.n3810 0.0105
R34236 DVSS.n4529 DVSS.n3808 0.0105
R34237 DVSS.n4578 DVSS.n3808 0.0105
R34238 DVSS.n4578 DVSS.n4577 0.0105
R34239 DVSS.n4577 DVSS.n4575 0.0105
R34240 DVSS.n4575 DVSS.n4573 0.0105
R34241 DVSS.n4573 DVSS.n4536 0.0105
R34242 DVSS.n4569 DVSS.n4536 0.0105
R34243 DVSS.n4569 DVSS.n4568 0.0105
R34244 DVSS.n4568 DVSS.n4567 0.0105
R34245 DVSS.n4567 DVSS.n4542 0.0105
R34246 DVSS.n4563 DVSS.n4542 0.0105
R34247 DVSS.n4563 DVSS.n4562 0.0105
R34248 DVSS.n4562 DVSS.n4561 0.0105
R34249 DVSS.n4561 DVSS.n4548 0.0105
R34250 DVSS.n4557 DVSS.n4548 0.0105
R34251 DVSS.n4557 DVSS.n4556 0.0105
R34252 DVSS.n4556 DVSS.n4555 0.0105
R34253 DVSS.n4555 DVSS.n3747 0.0105
R34254 DVSS.n4780 DVSS.n3747 0.0105
R34255 DVSS.n4780 DVSS.n4779 0.0105
R34256 DVSS.n4779 DVSS.n4777 0.0105
R34257 DVSS.n4777 DVSS.n3751 0.0105
R34258 DVSS.n4773 DVSS.n3751 0.0105
R34259 DVSS.n4773 DVSS.n4772 0.0105
R34260 DVSS.n4772 DVSS.n4771 0.0105
R34261 DVSS.n4771 DVSS.n3757 0.0105
R34262 DVSS.n4767 DVSS.n3757 0.0105
R34263 DVSS.n4767 DVSS.n4766 0.0105
R34264 DVSS.n4766 DVSS.n4765 0.0105
R34265 DVSS.n4765 DVSS.n3763 0.0105
R34266 DVSS.n4761 DVSS.n3763 0.0105
R34267 DVSS.n4761 DVSS.n4760 0.0105
R34268 DVSS.n4760 DVSS.n4759 0.0105
R34269 DVSS.n4759 DVSS.n3769 0.0105
R34270 DVSS.n4609 DVSS.n3769 0.0105
R34271 DVSS.n4753 DVSS.n4609 0.0105
R34272 DVSS.n4753 DVSS.n4752 0.0105
R34273 DVSS.n4752 DVSS.n4751 0.0105
R34274 DVSS.n4751 DVSS.n4615 0.0105
R34275 DVSS.n4743 DVSS.n4615 0.0105
R34276 DVSS.n4743 DVSS.n4742 0.0105
R34277 DVSS.n4742 DVSS.n4741 0.0105
R34278 DVSS.n4741 DVSS.n4710 0.0105
R34279 DVSS.n4737 DVSS.n4710 0.0105
R34280 DVSS.n4737 DVSS.n4736 0.0105
R34281 DVSS.n4736 DVSS.n4735 0.0105
R34282 DVSS.n4735 DVSS.n4716 0.0105
R34283 DVSS.n4731 DVSS.n4716 0.0105
R34284 DVSS.n4731 DVSS.n4730 0.0105
R34285 DVSS.n4730 DVSS.n4729 0.0105
R34286 DVSS.n4729 DVSS.n4726 0.0105
R34287 DVSS.n4726 DVSS.n4725 0.0105
R34288 DVSS.n4725 DVSS.n2794 0.0105
R34289 DVSS.n5998 DVSS.n2794 0.0105
R34290 DVSS.n5998 DVSS.n5997 0.0105
R34291 DVSS.n5997 DVSS.n5995 0.0105
R34292 DVSS.n5995 DVSS.n2798 0.0105
R34293 DVSS.n5991 DVSS.n2798 0.0105
R34294 DVSS.n5991 DVSS.n5990 0.0105
R34295 DVSS.n5990 DVSS.n5989 0.0105
R34296 DVSS.n5989 DVSS.n2804 0.0105
R34297 DVSS.n5985 DVSS.n2804 0.0105
R34298 DVSS.n5985 DVSS.n5984 0.0105
R34299 DVSS.n5984 DVSS.n5983 0.0105
R34300 DVSS.n5983 DVSS.n2810 0.0105
R34301 DVSS.n5979 DVSS.n2810 0.0105
R34302 DVSS.n5979 DVSS.n5978 0.0105
R34303 DVSS.n5978 DVSS.n5977 0.0105
R34304 DVSS.n5977 DVSS.n2816 0.0105
R34305 DVSS.n5971 DVSS.n2816 0.0105
R34306 DVSS.n5971 DVSS.n5970 0.0105
R34307 DVSS.n5970 DVSS.n5968 0.0105
R34308 DVSS.n5968 DVSS.n2841 0.0105
R34309 DVSS.n5964 DVSS.n2841 0.0105
R34310 DVSS.n5964 DVSS.n5963 0.0105
R34311 DVSS.n5963 DVSS.n5962 0.0105
R34312 DVSS.n5962 DVSS.n2847 0.0105
R34313 DVSS.n5954 DVSS.n2847 0.0105
R34314 DVSS.n5954 DVSS.n5953 0.0105
R34315 DVSS.n5953 DVSS.n5951 0.0105
R34316 DVSS.n5951 DVSS.n2870 0.0105
R34317 DVSS.n5947 DVSS.n2870 0.0105
R34318 DVSS.n5947 DVSS.n5946 0.0105
R34319 DVSS.n5945 DVSS.n2876 0.0105
R34320 DVSS.n5939 DVSS.n2876 0.0105
R34321 DVSS.n5939 DVSS.n5938 0.0105
R34322 DVSS.n4499 DVSS.n3830 0.0105
R34323 DVSS.n4500 DVSS.n4499 0.0105
R34324 DVSS.n4502 DVSS.n4500 0.0105
R34325 DVSS.n4502 DVSS.n4501 0.0105
R34326 DVSS.n4526 DVSS.n3811 0.0105
R34327 DVSS.n4527 DVSS.n4526 0.0105
R34328 DVSS.n4528 DVSS.n4527 0.0105
R34329 DVSS.n4528 DVSS.n3802 0.0105
R34330 DVSS.n4572 DVSS.n4571 0.0105
R34331 DVSS.n4571 DVSS.n4570 0.0105
R34332 DVSS.n4570 DVSS.n4537 0.0105
R34333 DVSS.n4566 DVSS.n4537 0.0105
R34334 DVSS.n4566 DVSS.n4565 0.0105
R34335 DVSS.n4565 DVSS.n4564 0.0105
R34336 DVSS.n4564 DVSS.n4543 0.0105
R34337 DVSS.n4560 DVSS.n4543 0.0105
R34338 DVSS.n4560 DVSS.n4559 0.0105
R34339 DVSS.n4559 DVSS.n4558 0.0105
R34340 DVSS.n4558 DVSS.n4549 0.0105
R34341 DVSS.n4549 DVSS.n3730 0.0105
R34342 DVSS.n4776 DVSS.n4775 0.0105
R34343 DVSS.n4775 DVSS.n4774 0.0105
R34344 DVSS.n4774 DVSS.n3752 0.0105
R34345 DVSS.n4770 DVSS.n3752 0.0105
R34346 DVSS.n4770 DVSS.n4769 0.0105
R34347 DVSS.n4769 DVSS.n4768 0.0105
R34348 DVSS.n4768 DVSS.n3758 0.0105
R34349 DVSS.n4764 DVSS.n3758 0.0105
R34350 DVSS.n4764 DVSS.n4763 0.0105
R34351 DVSS.n4763 DVSS.n4762 0.0105
R34352 DVSS.n4762 DVSS.n3764 0.0105
R34353 DVSS.n4758 DVSS.n3764 0.0105
R34354 DVSS.n4754 DVSS.n4608 0.0105
R34355 DVSS.n4744 DVSS.n4705 0.0105
R34356 DVSS.n4740 DVSS.n4705 0.0105
R34357 DVSS.n4740 DVSS.n4739 0.0105
R34358 DVSS.n4739 DVSS.n4738 0.0105
R34359 DVSS.n4738 DVSS.n4711 0.0105
R34360 DVSS.n4734 DVSS.n4711 0.0105
R34361 DVSS.n4734 DVSS.n4733 0.0105
R34362 DVSS.n4733 DVSS.n4732 0.0105
R34363 DVSS.n4732 DVSS.n4717 0.0105
R34364 DVSS.n4728 DVSS.n4717 0.0105
R34365 DVSS.n4728 DVSS.n4727 0.0105
R34366 DVSS.n4727 DVSS.n2783 0.0105
R34367 DVSS.n5994 DVSS.n5993 0.0105
R34368 DVSS.n5993 DVSS.n5992 0.0105
R34369 DVSS.n5992 DVSS.n2799 0.0105
R34370 DVSS.n5988 DVSS.n2799 0.0105
R34371 DVSS.n5988 DVSS.n5987 0.0105
R34372 DVSS.n5987 DVSS.n5986 0.0105
R34373 DVSS.n5986 DVSS.n2805 0.0105
R34374 DVSS.n5982 DVSS.n2805 0.0105
R34375 DVSS.n5982 DVSS.n5981 0.0105
R34376 DVSS.n5981 DVSS.n5980 0.0105
R34377 DVSS.n5980 DVSS.n2811 0.0105
R34378 DVSS.n5976 DVSS.n2811 0.0105
R34379 DVSS.n5967 DVSS.n5966 0.0105
R34380 DVSS.n5966 DVSS.n5965 0.0105
R34381 DVSS.n5965 DVSS.n2842 0.0105
R34382 DVSS.n5961 DVSS.n2842 0.0105
R34383 DVSS.n5950 DVSS.n5949 0.0105
R34384 DVSS.n5949 DVSS.n5948 0.0105
R34385 DVSS.n5948 DVSS.n2871 0.0105
R34386 DVSS.n3686 DVSS.n3681 0.0104296
R34387 DVSS.n5560 DVSS.n2288 0.0104296
R34388 DVSS.n7876 DVSS.n2070 0.0104296
R34389 DVSS.n3695 DVSS.n3694 0.0104296
R34390 DVSS.n5607 DVSS.n2318 0.0104296
R34391 DVSS.n7877 DVSS.n2052 0.0104296
R34392 DVSS.n2831 DVSS.n2821 0.0102441
R34393 DVSS.n2778 DVSS.n2768 0.0102441
R34394 DVSS.n3744 DVSS.n3734 0.0102441
R34395 DVSS.n4590 DVSS.n4589 0.0102441
R34396 DVSS.n8887 DVSS.n771 0.0102441
R34397 DVSS.n8984 DVSS.n747 0.0102441
R34398 DVSS.n3826 DVSS.n3818 0.0102441
R34399 DVSS.n2864 DVSS.n2852 0.0102441
R34400 DVSS.n9421 DVSS.n355 0.0102441
R34401 DVSS.n9518 DVSS.n45 0.0102441
R34402 DVSS.n5928 DVSS.n2881 0.0102441
R34403 DVSS.n5371 DVSS.n2955 0.0102441
R34404 DVSS.n4478 DVSS.n4454 0.0102441
R34405 DVSS.n5878 DVSS.n5877 0.0102441
R34406 DVSS.n4658 DVSS.n3685 0.010007
R34407 DVSS.n5562 DVSS.n2297 0.010007
R34408 DVSS.n7870 DVSS.n2067 0.010007
R34409 DVSS.n4662 DVSS.n3699 0.010007
R34410 DVSS.n5603 DVSS.n2327 0.010007
R34411 DVSS.n7871 DVSS.n2049 0.010007
R34412 DVSS.n2905 DVSS.n2821 0.00988976
R34413 DVSS.n3355 DVSS.n3351 0.00988976
R34414 DVSS.n5384 DVSS.n3357 0.00988976
R34415 DVSS.n5072 DVSS.n3354 0.00988976
R34416 DVSS.n5071 DVSS.n5066 0.00988976
R34417 DVSS.n5129 DVSS.n3353 0.00988976
R34418 DVSS.n6005 DVSS.n2778 0.00988976
R34419 DVSS.n3347 DVSS.n3343 0.00988976
R34420 DVSS.n5388 DVSS.n3330 0.00988976
R34421 DVSS.n5392 DVSS.n3344 0.00988976
R34422 DVSS.n5391 DVSS.n3329 0.00988976
R34423 DVSS.n5394 DVSS.n3324 0.00988976
R34424 DVSS.n4598 DVSS.n3734 0.00988976
R34425 DVSS.n3524 DVSS.n3154 0.00988976
R34426 DVSS.n3554 DVSS.n3143 0.00988976
R34427 DVSS.n3526 DVSS.n3155 0.00988976
R34428 DVSS.n3550 DVSS.n3142 0.00988976
R34429 DVSS.n5776 DVSS.n3156 0.00988976
R34430 DVSS.n4589 DVSS.n3792 0.00988976
R34431 DVSS.n3529 DVSS.n3109 0.00988976
R34432 DVSS.n3546 DVSS.n3101 0.00988976
R34433 DVSS.n3531 DVSS.n3110 0.00988976
R34434 DVSS.n3542 DVSS.n3100 0.00988976
R34435 DVSS.n5812 DVSS.n3111 0.00988976
R34436 DVSS.n8889 DVSS.n771 0.00988976
R34437 DVSS.n8986 DVSS.n747 0.00988976
R34438 DVSS.n4471 DVSS.n3818 0.00988976
R34439 DVSS.n2909 DVSS.n2852 0.00988976
R34440 DVSS.n3365 DVSS.n3361 0.00988976
R34441 DVSS.n5381 DVSS.n3367 0.00988976
R34442 DVSS.n3370 DVSS.n3364 0.00988976
R34443 DVSS.n5368 DVSS.n5367 0.00988976
R34444 DVSS.n5365 DVSS.n3363 0.00988976
R34445 DVSS.n9423 DVSS.n355 0.00988976
R34446 DVSS.n9520 DVSS.n45 0.00988976
R34447 DVSS.n5924 DVSS.n2881 0.00988976
R34448 DVSS.n5372 DVSS.n2955 0.00988976
R34449 DVSS.n4475 DVSS.n4454 0.00988976
R34450 DVSS.n5878 DVSS.n3013 0.00988976
R34451 DVSS.n4758 DVSS.n4757 0.00979577
R34452 DVSS.n4237 DVSS.n4235 0.00962857
R34453 DVSS.n4239 DVSS.n4237 0.00962857
R34454 DVSS.n4239 DVSS.n4233 0.00962857
R34455 DVSS.n4243 DVSS.n4233 0.00962857
R34456 DVSS.n4243 DVSS.n4231 0.00962857
R34457 DVSS.n4247 DVSS.n4231 0.00962857
R34458 DVSS.n4247 DVSS.n4229 0.00962857
R34459 DVSS.n4251 DVSS.n4229 0.00962857
R34460 DVSS.n4251 DVSS.n4214 0.00962857
R34461 DVSS.n4262 DVSS.n4214 0.00962857
R34462 DVSS.n4262 DVSS.n4212 0.00962857
R34463 DVSS.n4266 DVSS.n4212 0.00962857
R34464 DVSS.n4266 DVSS.n4210 0.00962857
R34465 DVSS.n4270 DVSS.n4210 0.00962857
R34466 DVSS.n4270 DVSS.n4206 0.00962857
R34467 DVSS.n4417 DVSS.n4206 0.00962857
R34468 DVSS.n4417 DVSS.n4208 0.00962857
R34469 DVSS.n4413 DVSS.n4208 0.00962857
R34470 DVSS.n4413 DVSS.n4411 0.00962857
R34471 DVSS.n4411 DVSS.n4274 0.00962857
R34472 DVSS.n4407 DVSS.n4274 0.00962857
R34473 DVSS.n4407 DVSS.n4276 0.00962857
R34474 DVSS.n4403 DVSS.n4276 0.00962857
R34475 DVSS.n4403 DVSS.n4279 0.00962857
R34476 DVSS.n4399 DVSS.n4279 0.00962857
R34477 DVSS.n4399 DVSS.n4281 0.00962857
R34478 DVSS.n4395 DVSS.n4281 0.00962857
R34479 DVSS.n4395 DVSS.n4283 0.00962857
R34480 DVSS.n4391 DVSS.n4283 0.00962857
R34481 DVSS.n4391 DVSS.n4285 0.00962857
R34482 DVSS.n4387 DVSS.n4285 0.00962857
R34483 DVSS.n4387 DVSS.n4386 0.00962857
R34484 DVSS.n4386 DVSS.n4385 0.00962857
R34485 DVSS.n4385 DVSS.n4288 0.00962857
R34486 DVSS.n4380 DVSS.n4288 0.00962857
R34487 DVSS.n4380 DVSS.n4290 0.00962857
R34488 DVSS.n4376 DVSS.n4290 0.00962857
R34489 DVSS.n4376 DVSS.n4292 0.00962857
R34490 DVSS.n4372 DVSS.n4292 0.00962857
R34491 DVSS.n4372 DVSS.n4294 0.00962857
R34492 DVSS.n4368 DVSS.n4294 0.00962857
R34493 DVSS.n4368 DVSS.n4296 0.00962857
R34494 DVSS.n4364 DVSS.n4296 0.00962857
R34495 DVSS.n4364 DVSS.n4298 0.00962857
R34496 DVSS.n4360 DVSS.n4298 0.00962857
R34497 DVSS.n4360 DVSS.n4300 0.00962857
R34498 DVSS.n4356 DVSS.n4300 0.00962857
R34499 DVSS.n4356 DVSS.n4355 0.00962857
R34500 DVSS.n4355 DVSS.n4354 0.00962857
R34501 DVSS.n4354 DVSS.n4303 0.00962857
R34502 DVSS.n4349 DVSS.n4303 0.00962857
R34503 DVSS.n4349 DVSS.n4348 0.00962857
R34504 DVSS.n4348 DVSS.n4347 0.00962857
R34505 DVSS.n4347 DVSS.n4305 0.00962857
R34506 DVSS.n4342 DVSS.n4305 0.00962857
R34507 DVSS.n4342 DVSS.n4307 0.00962857
R34508 DVSS.n4338 DVSS.n4307 0.00962857
R34509 DVSS.n4338 DVSS.n4310 0.00962857
R34510 DVSS.n4334 DVSS.n4310 0.00962857
R34511 DVSS.n4334 DVSS.n4312 0.00962857
R34512 DVSS.n4330 DVSS.n4312 0.00962857
R34513 DVSS.n4330 DVSS.n4314 0.00962857
R34514 DVSS.n4326 DVSS.n4314 0.00962857
R34515 DVSS.n4326 DVSS.n4316 0.00962857
R34516 DVSS.n4322 DVSS.n4316 0.00962857
R34517 DVSS.n4322 DVSS.n4317 0.00962857
R34518 DVSS.n4318 DVSS.n4317 0.00962857
R34519 DVSS.n4318 DVSS.n3646 0.00962857
R34520 DVSS.n4852 DVSS.n3646 0.00962857
R34521 DVSS.n4852 DVSS.n3644 0.00962857
R34522 DVSS.n4856 DVSS.n3644 0.00962857
R34523 DVSS.n4856 DVSS.n3642 0.00962857
R34524 DVSS.n4860 DVSS.n3642 0.00962857
R34525 DVSS.n4860 DVSS.n3640 0.00962857
R34526 DVSS.n4864 DVSS.n3640 0.00962857
R34527 DVSS.n4864 DVSS.n3638 0.00962857
R34528 DVSS.n4868 DVSS.n3638 0.00962857
R34529 DVSS.n4868 DVSS.n3636 0.00962857
R34530 DVSS.n4872 DVSS.n3636 0.00962857
R34531 DVSS.n4872 DVSS.n3634 0.00962857
R34532 DVSS.n4876 DVSS.n3634 0.00962857
R34533 DVSS.n4876 DVSS.n3632 0.00962857
R34534 DVSS.n4880 DVSS.n3632 0.00962857
R34535 DVSS.n4880 DVSS.n3613 0.00962857
R34536 DVSS.n4890 DVSS.n3613 0.00962857
R34537 DVSS.n4890 DVSS.n3611 0.00962857
R34538 DVSS.n4894 DVSS.n3611 0.00962857
R34539 DVSS.n4894 DVSS.n3609 0.00962857
R34540 DVSS.n4898 DVSS.n3609 0.00962857
R34541 DVSS.n4898 DVSS.n3605 0.00962857
R34542 DVSS.n4960 DVSS.n3605 0.00962857
R34543 DVSS.n4960 DVSS.n3607 0.00962857
R34544 DVSS.n4956 DVSS.n3607 0.00962857
R34545 DVSS.n4956 DVSS.n4954 0.00962857
R34546 DVSS.n4954 DVSS.n4902 0.00962857
R34547 DVSS.n4950 DVSS.n4902 0.00962857
R34548 DVSS.n4950 DVSS.n4904 0.00962857
R34549 DVSS.n4946 DVSS.n4906 0.00962857
R34550 DVSS.n4936 DVSS.n4906 0.00962857
R34551 DVSS.n4940 DVSS.n4936 0.00962857
R34552 DVSS.n6768 DVSS.n6766 0.00962857
R34553 DVSS.n6768 DVSS.n6764 0.00962857
R34554 DVSS.n6849 DVSS.n6764 0.00962857
R34555 DVSS.n6849 DVSS.n6765 0.00962857
R34556 DVSS.n6845 DVSS.n6765 0.00962857
R34557 DVSS.n6845 DVSS.n6842 0.00962857
R34558 DVSS.n6842 DVSS.n6841 0.00962857
R34559 DVSS.n6841 DVSS.n6772 0.00962857
R34560 DVSS.n6837 DVSS.n6772 0.00962857
R34561 DVSS.n6837 DVSS.n6835 0.00962857
R34562 DVSS.n6835 DVSS.n6833 0.00962857
R34563 DVSS.n6833 DVSS.n6774 0.00962857
R34564 DVSS.n6829 DVSS.n6774 0.00962857
R34565 DVSS.n6829 DVSS.n6777 0.00962857
R34566 DVSS.n6825 DVSS.n6777 0.00962857
R34567 DVSS.n6825 DVSS.n6824 0.00962857
R34568 DVSS.n6824 DVSS.n6823 0.00962857
R34569 DVSS.n6823 DVSS.n6781 0.00962857
R34570 DVSS.n6818 DVSS.n6781 0.00962857
R34571 DVSS.n6818 DVSS.n6783 0.00962857
R34572 DVSS.n6814 DVSS.n6783 0.00962857
R34573 DVSS.n6814 DVSS.n6785 0.00962857
R34574 DVSS.n6810 DVSS.n6785 0.00962857
R34575 DVSS.n6810 DVSS.n6787 0.00962857
R34576 DVSS.n6806 DVSS.n6787 0.00962857
R34577 DVSS.n6806 DVSS.n6789 0.00962857
R34578 DVSS.n6802 DVSS.n6789 0.00962857
R34579 DVSS.n6802 DVSS.n6791 0.00962857
R34580 DVSS.n6798 DVSS.n6791 0.00962857
R34581 DVSS.n6798 DVSS.n6793 0.00962857
R34582 DVSS.n6794 DVSS.n6793 0.00962857
R34583 DVSS.n6794 DVSS.n1344 0.00962857
R34584 DVSS.n8433 DVSS.n1344 0.00962857
R34585 DVSS.n8433 DVSS.n1346 0.00962857
R34586 DVSS.n8429 DVSS.n1346 0.00962857
R34587 DVSS.n8429 DVSS.n1349 0.00962857
R34588 DVSS.n8425 DVSS.n1349 0.00962857
R34589 DVSS.n8425 DVSS.n1351 0.00962857
R34590 DVSS.n8421 DVSS.n1351 0.00962857
R34591 DVSS.n8421 DVSS.n1353 0.00962857
R34592 DVSS.n8417 DVSS.n1353 0.00962857
R34593 DVSS.n8417 DVSS.n1355 0.00962857
R34594 DVSS.n8413 DVSS.n1355 0.00962857
R34595 DVSS.n8413 DVSS.n1357 0.00962857
R34596 DVSS.n8409 DVSS.n1357 0.00962857
R34597 DVSS.n8409 DVSS.n1359 0.00962857
R34598 DVSS.n8405 DVSS.n1359 0.00962857
R34599 DVSS.n8405 DVSS.n1361 0.00962857
R34600 DVSS.n1393 DVSS.n1361 0.00962857
R34601 DVSS.n8398 DVSS.n1393 0.00962857
R34602 DVSS.n8398 DVSS.n1394 0.00962857
R34603 DVSS.n8394 DVSS.n1394 0.00962857
R34604 DVSS.n8394 DVSS.n1397 0.00962857
R34605 DVSS.n1637 DVSS.n1397 0.00962857
R34606 DVSS.n1640 DVSS.n1637 0.00962857
R34607 DVSS.n1640 DVSS.n1636 0.00962857
R34608 DVSS.n1644 DVSS.n1636 0.00962857
R34609 DVSS.n1644 DVSS.n1634 0.00962857
R34610 DVSS.n1648 DVSS.n1634 0.00962857
R34611 DVSS.n1648 DVSS.n1632 0.00962857
R34612 DVSS.n1652 DVSS.n1632 0.00962857
R34613 DVSS.n1652 DVSS.n1630 0.00962857
R34614 DVSS.n1656 DVSS.n1630 0.00962857
R34615 DVSS.n1656 DVSS.n1628 0.00962857
R34616 DVSS.n1660 DVSS.n1628 0.00962857
R34617 DVSS.n1660 DVSS.n1626 0.00962857
R34618 DVSS.n1664 DVSS.n1626 0.00962857
R34619 DVSS.n1666 DVSS.n1664 0.00962857
R34620 DVSS.n1668 DVSS.n1666 0.00962857
R34621 DVSS.n1668 DVSS.n1624 0.00962857
R34622 DVSS.n1672 DVSS.n1624 0.00962857
R34623 DVSS.n1672 DVSS.n1622 0.00962857
R34624 DVSS.n1676 DVSS.n1622 0.00962857
R34625 DVSS.n1676 DVSS.n1620 0.00962857
R34626 DVSS.n1680 DVSS.n1620 0.00962857
R34627 DVSS.n1680 DVSS.n1618 0.00962857
R34628 DVSS.n1684 DVSS.n1618 0.00962857
R34629 DVSS.n1684 DVSS.n1616 0.00962857
R34630 DVSS.n1688 DVSS.n1616 0.00962857
R34631 DVSS.n1688 DVSS.n1614 0.00962857
R34632 DVSS.n1692 DVSS.n1614 0.00962857
R34633 DVSS.n1692 DVSS.n1612 0.00962857
R34634 DVSS.n1696 DVSS.n1612 0.00962857
R34635 DVSS.n1698 DVSS.n1696 0.00962857
R34636 DVSS.n1700 DVSS.n1698 0.00962857
R34637 DVSS.n1700 DVSS.n1610 0.00962857
R34638 DVSS.n1704 DVSS.n1610 0.00962857
R34639 DVSS.n1704 DVSS.n1608 0.00962857
R34640 DVSS.n1708 DVSS.n1608 0.00962857
R34641 DVSS.n1708 DVSS.n1606 0.00962857
R34642 DVSS.n1712 DVSS.n1606 0.00962857
R34643 DVSS.n1712 DVSS.n1593 0.00962857
R34644 DVSS.n1729 DVSS.n1593 0.00962857
R34645 DVSS.n1729 DVSS.n1591 0.00962857
R34646 DVSS.n1734 DVSS.n1591 0.00962857
R34647 DVSS.n1734 DVSS.n1589 0.00962857
R34648 DVSS.n1738 DVSS.n1589 0.00962857
R34649 DVSS.n1739 DVSS.n1585 0.00962857
R34650 DVSS.n1744 DVSS.n1585 0.00962857
R34651 DVSS.n1744 DVSS.n1587 0.00962857
R34652 DVSS.n6850 DVSS.n6763 0.00962857
R34653 DVSS.n6844 DVSS.n6763 0.00962857
R34654 DVSS.n6844 DVSS.n6843 0.00962857
R34655 DVSS.n6843 DVSS.n6669 0.00962857
R34656 DVSS.n6832 DVSS.n6831 0.00962857
R34657 DVSS.n6831 DVSS.n6830 0.00962857
R34658 DVSS.n6830 DVSS.n6776 0.00962857
R34659 DVSS.n6776 DVSS.n1164 0.00962857
R34660 DVSS.n6817 DVSS.n6816 0.00962857
R34661 DVSS.n6816 DVSS.n6815 0.00962857
R34662 DVSS.n6815 DVSS.n6784 0.00962857
R34663 DVSS.n6809 DVSS.n6784 0.00962857
R34664 DVSS.n6809 DVSS.n6808 0.00962857
R34665 DVSS.n6808 DVSS.n6807 0.00962857
R34666 DVSS.n6807 DVSS.n6788 0.00962857
R34667 DVSS.n6801 DVSS.n6788 0.00962857
R34668 DVSS.n6801 DVSS.n6800 0.00962857
R34669 DVSS.n6800 DVSS.n6799 0.00962857
R34670 DVSS.n6799 DVSS.n6792 0.00962857
R34671 DVSS.n6792 DVSS.n1328 0.00962857
R34672 DVSS.n8428 DVSS.n8427 0.00962857
R34673 DVSS.n8427 DVSS.n8426 0.00962857
R34674 DVSS.n8426 DVSS.n1350 0.00962857
R34675 DVSS.n8420 DVSS.n1350 0.00962857
R34676 DVSS.n8420 DVSS.n8419 0.00962857
R34677 DVSS.n8419 DVSS.n8418 0.00962857
R34678 DVSS.n8418 DVSS.n1354 0.00962857
R34679 DVSS.n8412 DVSS.n1354 0.00962857
R34680 DVSS.n8412 DVSS.n8411 0.00962857
R34681 DVSS.n8411 DVSS.n8410 0.00962857
R34682 DVSS.n8410 DVSS.n1358 0.00962857
R34683 DVSS.n8404 DVSS.n1358 0.00962857
R34684 DVSS.n8399 DVSS.n1392 0.00962857
R34685 DVSS.n1641 DVSS.n1414 0.00962857
R34686 DVSS.n1642 DVSS.n1641 0.00962857
R34687 DVSS.n1643 DVSS.n1642 0.00962857
R34688 DVSS.n1643 DVSS.n1633 0.00962857
R34689 DVSS.n1649 DVSS.n1633 0.00962857
R34690 DVSS.n1650 DVSS.n1649 0.00962857
R34691 DVSS.n1651 DVSS.n1650 0.00962857
R34692 DVSS.n1651 DVSS.n1629 0.00962857
R34693 DVSS.n1657 DVSS.n1629 0.00962857
R34694 DVSS.n1658 DVSS.n1657 0.00962857
R34695 DVSS.n1659 DVSS.n1658 0.00962857
R34696 DVSS.n1659 DVSS.n1428 0.00962857
R34697 DVSS.n1673 DVSS.n1623 0.00962857
R34698 DVSS.n1674 DVSS.n1673 0.00962857
R34699 DVSS.n1675 DVSS.n1674 0.00962857
R34700 DVSS.n1675 DVSS.n1619 0.00962857
R34701 DVSS.n1681 DVSS.n1619 0.00962857
R34702 DVSS.n1682 DVSS.n1681 0.00962857
R34703 DVSS.n1683 DVSS.n1682 0.00962857
R34704 DVSS.n1683 DVSS.n1615 0.00962857
R34705 DVSS.n1689 DVSS.n1615 0.00962857
R34706 DVSS.n1690 DVSS.n1689 0.00962857
R34707 DVSS.n1691 DVSS.n1690 0.00962857
R34708 DVSS.n1691 DVSS.n1108 0.00962857
R34709 DVSS.n1705 DVSS.n1609 0.00962857
R34710 DVSS.n1706 DVSS.n1705 0.00962857
R34711 DVSS.n1707 DVSS.n1706 0.00962857
R34712 DVSS.n1707 DVSS.n1601 0.00962857
R34713 DVSS.n1735 DVSS.n1590 0.00962857
R34714 DVSS.n1736 DVSS.n1735 0.00962857
R34715 DVSS.n1737 DVSS.n1736 0.00962857
R34716 DVSS.n1940 DVSS.n1938 0.00962857
R34717 DVSS.n1940 DVSS.n1936 0.00962857
R34718 DVSS.n8051 DVSS.n1936 0.00962857
R34719 DVSS.n8051 DVSS.n1937 0.00962857
R34720 DVSS.n8047 DVSS.n1937 0.00962857
R34721 DVSS.n8047 DVSS.n1944 0.00962857
R34722 DVSS.n8043 DVSS.n1944 0.00962857
R34723 DVSS.n8043 DVSS.n1946 0.00962857
R34724 DVSS.n8039 DVSS.n1946 0.00962857
R34725 DVSS.n8039 DVSS.n1948 0.00962857
R34726 DVSS.n8028 DVSS.n1948 0.00962857
R34727 DVSS.n8028 DVSS.n1968 0.00962857
R34728 DVSS.n8024 DVSS.n1968 0.00962857
R34729 DVSS.n8024 DVSS.n1970 0.00962857
R34730 DVSS.n8020 DVSS.n1970 0.00962857
R34731 DVSS.n8020 DVSS.n1972 0.00962857
R34732 DVSS.n8016 DVSS.n1972 0.00962857
R34733 DVSS.n8016 DVSS.n1974 0.00962857
R34734 DVSS.n8005 DVSS.n1974 0.00962857
R34735 DVSS.n8005 DVSS.n1994 0.00962857
R34736 DVSS.n8001 DVSS.n1994 0.00962857
R34737 DVSS.n8001 DVSS.n1996 0.00962857
R34738 DVSS.n7997 DVSS.n1996 0.00962857
R34739 DVSS.n7997 DVSS.n1998 0.00962857
R34740 DVSS.n7993 DVSS.n1998 0.00962857
R34741 DVSS.n7993 DVSS.n2000 0.00962857
R34742 DVSS.n7989 DVSS.n2000 0.00962857
R34743 DVSS.n7989 DVSS.n2002 0.00962857
R34744 DVSS.n7985 DVSS.n2002 0.00962857
R34745 DVSS.n7985 DVSS.n2004 0.00962857
R34746 DVSS.n7981 DVSS.n2004 0.00962857
R34747 DVSS.n7981 DVSS.n2006 0.00962857
R34748 DVSS.n7977 DVSS.n2006 0.00962857
R34749 DVSS.n7977 DVSS.n2008 0.00962857
R34750 DVSS.n7966 DVSS.n2008 0.00962857
R34751 DVSS.n7966 DVSS.n2028 0.00962857
R34752 DVSS.n7962 DVSS.n2028 0.00962857
R34753 DVSS.n7962 DVSS.n2030 0.00962857
R34754 DVSS.n7958 DVSS.n2030 0.00962857
R34755 DVSS.n7958 DVSS.n2032 0.00962857
R34756 DVSS.n7954 DVSS.n2032 0.00962857
R34757 DVSS.n7954 DVSS.n2034 0.00962857
R34758 DVSS.n7950 DVSS.n2034 0.00962857
R34759 DVSS.n7950 DVSS.n2036 0.00962857
R34760 DVSS.n7946 DVSS.n2036 0.00962857
R34761 DVSS.n7946 DVSS.n2038 0.00962857
R34762 DVSS.n7942 DVSS.n2038 0.00962857
R34763 DVSS.n7942 DVSS.n2040 0.00962857
R34764 DVSS.n7938 DVSS.n2040 0.00962857
R34765 DVSS.n7938 DVSS.n2042 0.00962857
R34766 DVSS.n7768 DVSS.n2042 0.00962857
R34767 DVSS.n7769 DVSS.n7768 0.00962857
R34768 DVSS.n7771 DVSS.n7769 0.00962857
R34769 DVSS.n7771 DVSS.n7765 0.00962857
R34770 DVSS.n7775 DVSS.n7765 0.00962857
R34771 DVSS.n7775 DVSS.n7763 0.00962857
R34772 DVSS.n7779 DVSS.n7763 0.00962857
R34773 DVSS.n7779 DVSS.n7761 0.00962857
R34774 DVSS.n7783 DVSS.n7761 0.00962857
R34775 DVSS.n7783 DVSS.n7759 0.00962857
R34776 DVSS.n7787 DVSS.n7759 0.00962857
R34777 DVSS.n7787 DVSS.n7757 0.00962857
R34778 DVSS.n7792 DVSS.n7757 0.00962857
R34779 DVSS.n7792 DVSS.n7755 0.00962857
R34780 DVSS.n7796 DVSS.n7755 0.00962857
R34781 DVSS.n7797 DVSS.n7796 0.00962857
R34782 DVSS.n7797 DVSS.n7751 0.00962857
R34783 DVSS.n7842 DVSS.n7751 0.00962857
R34784 DVSS.n7842 DVSS.n7753 0.00962857
R34785 DVSS.n7838 DVSS.n7753 0.00962857
R34786 DVSS.n7838 DVSS.n7801 0.00962857
R34787 DVSS.n7834 DVSS.n7801 0.00962857
R34788 DVSS.n7834 DVSS.n7803 0.00962857
R34789 DVSS.n7830 DVSS.n7803 0.00962857
R34790 DVSS.n7830 DVSS.n7805 0.00962857
R34791 DVSS.n7826 DVSS.n7805 0.00962857
R34792 DVSS.n7826 DVSS.n7807 0.00962857
R34793 DVSS.n7822 DVSS.n7807 0.00962857
R34794 DVSS.n7822 DVSS.n7809 0.00962857
R34795 DVSS.n7818 DVSS.n7809 0.00962857
R34796 DVSS.n7818 DVSS.n7811 0.00962857
R34797 DVSS.n7814 DVSS.n7811 0.00962857
R34798 DVSS.n7814 DVSS.n7813 0.00962857
R34799 DVSS.n7813 DVSS.n1807 0.00962857
R34800 DVSS.n8125 DVSS.n1807 0.00962857
R34801 DVSS.n8125 DVSS.n1805 0.00962857
R34802 DVSS.n8129 DVSS.n1805 0.00962857
R34803 DVSS.n8129 DVSS.n1803 0.00962857
R34804 DVSS.n8133 DVSS.n1803 0.00962857
R34805 DVSS.n8133 DVSS.n1801 0.00962857
R34806 DVSS.n8137 DVSS.n1801 0.00962857
R34807 DVSS.n8137 DVSS.n1787 0.00962857
R34808 DVSS.n8154 DVSS.n1787 0.00962857
R34809 DVSS.n8154 DVSS.n1785 0.00962857
R34810 DVSS.n8158 DVSS.n1785 0.00962857
R34811 DVSS.n8158 DVSS.n1783 0.00962857
R34812 DVSS.n8162 DVSS.n1783 0.00962857
R34813 DVSS.n8166 DVSS.n8165 0.00962857
R34814 DVSS.n8168 DVSS.n8166 0.00962857
R34815 DVSS.n8168 DVSS.n1780 0.00962857
R34816 DVSS.n8052 DVSS.n1935 0.00962857
R34817 DVSS.n8046 DVSS.n1935 0.00962857
R34818 DVSS.n8046 DVSS.n8045 0.00962857
R34819 DVSS.n8045 DVSS.n8044 0.00962857
R34820 DVSS.n8029 DVSS.n1967 0.00962857
R34821 DVSS.n8023 DVSS.n1967 0.00962857
R34822 DVSS.n8023 DVSS.n8022 0.00962857
R34823 DVSS.n8022 DVSS.n8021 0.00962857
R34824 DVSS.n8006 DVSS.n1993 0.00962857
R34825 DVSS.n8000 DVSS.n1993 0.00962857
R34826 DVSS.n8000 DVSS.n7999 0.00962857
R34827 DVSS.n7999 DVSS.n7998 0.00962857
R34828 DVSS.n7998 DVSS.n1997 0.00962857
R34829 DVSS.n7992 DVSS.n1997 0.00962857
R34830 DVSS.n7992 DVSS.n7991 0.00962857
R34831 DVSS.n7991 DVSS.n7990 0.00962857
R34832 DVSS.n7990 DVSS.n2001 0.00962857
R34833 DVSS.n7984 DVSS.n2001 0.00962857
R34834 DVSS.n7984 DVSS.n7983 0.00962857
R34835 DVSS.n7983 DVSS.n7982 0.00962857
R34836 DVSS.n7967 DVSS.n2027 0.00962857
R34837 DVSS.n7961 DVSS.n2027 0.00962857
R34838 DVSS.n7961 DVSS.n7960 0.00962857
R34839 DVSS.n7960 DVSS.n7959 0.00962857
R34840 DVSS.n7959 DVSS.n2031 0.00962857
R34841 DVSS.n7953 DVSS.n2031 0.00962857
R34842 DVSS.n7953 DVSS.n7952 0.00962857
R34843 DVSS.n7952 DVSS.n7951 0.00962857
R34844 DVSS.n7951 DVSS.n2035 0.00962857
R34845 DVSS.n7945 DVSS.n2035 0.00962857
R34846 DVSS.n7945 DVSS.n7944 0.00962857
R34847 DVSS.n7944 DVSS.n7943 0.00962857
R34848 DVSS.n2062 DVSS.n2050 0.00962857
R34849 DVSS.n7776 DVSS.n7764 0.00962857
R34850 DVSS.n7777 DVSS.n7776 0.00962857
R34851 DVSS.n7778 DVSS.n7777 0.00962857
R34852 DVSS.n7778 DVSS.n7760 0.00962857
R34853 DVSS.n7784 DVSS.n7760 0.00962857
R34854 DVSS.n7785 DVSS.n7784 0.00962857
R34855 DVSS.n7786 DVSS.n7785 0.00962857
R34856 DVSS.n7786 DVSS.n7756 0.00962857
R34857 DVSS.n7793 DVSS.n7756 0.00962857
R34858 DVSS.n7794 DVSS.n7793 0.00962857
R34859 DVSS.n7795 DVSS.n7794 0.00962857
R34860 DVSS.n7795 DVSS.n7731 0.00962857
R34861 DVSS.n7837 DVSS.n7836 0.00962857
R34862 DVSS.n7836 DVSS.n7835 0.00962857
R34863 DVSS.n7835 DVSS.n7802 0.00962857
R34864 DVSS.n7829 DVSS.n7802 0.00962857
R34865 DVSS.n7829 DVSS.n7828 0.00962857
R34866 DVSS.n7828 DVSS.n7827 0.00962857
R34867 DVSS.n7827 DVSS.n7806 0.00962857
R34868 DVSS.n7821 DVSS.n7806 0.00962857
R34869 DVSS.n7821 DVSS.n7820 0.00962857
R34870 DVSS.n7820 DVSS.n7819 0.00962857
R34871 DVSS.n7819 DVSS.n7810 0.00962857
R34872 DVSS.n7810 DVSS.n1816 0.00962857
R34873 DVSS.n8130 DVSS.n1804 0.00962857
R34874 DVSS.n8131 DVSS.n8130 0.00962857
R34875 DVSS.n8132 DVSS.n8131 0.00962857
R34876 DVSS.n8132 DVSS.n1796 0.00962857
R34877 DVSS.n8159 DVSS.n1784 0.00962857
R34878 DVSS.n8160 DVSS.n8159 0.00962857
R34879 DVSS.n8161 DVSS.n8160 0.00962857
R34880 DVSS.n3079 DVSS.n3077 0.00962857
R34881 DVSS.n3081 DVSS.n3079 0.00962857
R34882 DVSS.n3081 DVSS.n3075 0.00962857
R34883 DVSS.n3086 DVSS.n3075 0.00962857
R34884 DVSS.n3086 DVSS.n3073 0.00962857
R34885 DVSS.n3090 DVSS.n3073 0.00962857
R34886 DVSS.n3091 DVSS.n3090 0.00962857
R34887 DVSS.n3091 DVSS.n3070 0.00962857
R34888 DVSS.n5827 DVSS.n3070 0.00962857
R34889 DVSS.n5827 DVSS.n3071 0.00962857
R34890 DVSS.n5823 DVSS.n3071 0.00962857
R34891 DVSS.n5823 DVSS.n3095 0.00962857
R34892 DVSS.n5819 DVSS.n3095 0.00962857
R34893 DVSS.n5819 DVSS.n3097 0.00962857
R34894 DVSS.n5815 DVSS.n3097 0.00962857
R34895 DVSS.n5815 DVSS.n3099 0.00962857
R34896 DVSS.n3123 DVSS.n3099 0.00962857
R34897 DVSS.n3123 DVSS.n3120 0.00962857
R34898 DVSS.n5807 DVSS.n3120 0.00962857
R34899 DVSS.n5807 DVSS.n3121 0.00962857
R34900 DVSS.n5803 DVSS.n3121 0.00962857
R34901 DVSS.n5803 DVSS.n3127 0.00962857
R34902 DVSS.n5799 DVSS.n3127 0.00962857
R34903 DVSS.n5799 DVSS.n3129 0.00962857
R34904 DVSS.n5795 DVSS.n3129 0.00962857
R34905 DVSS.n5795 DVSS.n3131 0.00962857
R34906 DVSS.n5791 DVSS.n3131 0.00962857
R34907 DVSS.n5791 DVSS.n3133 0.00962857
R34908 DVSS.n5787 DVSS.n3133 0.00962857
R34909 DVSS.n5787 DVSS.n3135 0.00962857
R34910 DVSS.n5783 DVSS.n3135 0.00962857
R34911 DVSS.n5783 DVSS.n3137 0.00962857
R34912 DVSS.n5779 DVSS.n3137 0.00962857
R34913 DVSS.n5779 DVSS.n3139 0.00962857
R34914 DVSS.n5771 DVSS.n3139 0.00962857
R34915 DVSS.n5771 DVSS.n3159 0.00962857
R34916 DVSS.n5767 DVSS.n3159 0.00962857
R34917 DVSS.n5767 DVSS.n3161 0.00962857
R34918 DVSS.n5763 DVSS.n3161 0.00962857
R34919 DVSS.n5763 DVSS.n3163 0.00962857
R34920 DVSS.n5759 DVSS.n3163 0.00962857
R34921 DVSS.n5759 DVSS.n3165 0.00962857
R34922 DVSS.n5755 DVSS.n3165 0.00962857
R34923 DVSS.n5755 DVSS.n3167 0.00962857
R34924 DVSS.n5751 DVSS.n3167 0.00962857
R34925 DVSS.n5751 DVSS.n3169 0.00962857
R34926 DVSS.n5747 DVSS.n3169 0.00962857
R34927 DVSS.n5747 DVSS.n3171 0.00962857
R34928 DVSS.n5743 DVSS.n3171 0.00962857
R34929 DVSS.n5743 DVSS.n3173 0.00962857
R34930 DVSS.n5033 DVSS.n3173 0.00962857
R34931 DVSS.n5033 DVSS.n5031 0.00962857
R34932 DVSS.n5192 DVSS.n5031 0.00962857
R34933 DVSS.n5192 DVSS.n5032 0.00962857
R34934 DVSS.n5188 DVSS.n5032 0.00962857
R34935 DVSS.n5188 DVSS.n5037 0.00962857
R34936 DVSS.n5184 DVSS.n5037 0.00962857
R34937 DVSS.n5184 DVSS.n5040 0.00962857
R34938 DVSS.n5180 DVSS.n5040 0.00962857
R34939 DVSS.n5180 DVSS.n5042 0.00962857
R34940 DVSS.n5176 DVSS.n5042 0.00962857
R34941 DVSS.n5176 DVSS.n5044 0.00962857
R34942 DVSS.n5172 DVSS.n5044 0.00962857
R34943 DVSS.n5172 DVSS.n5046 0.00962857
R34944 DVSS.n5168 DVSS.n5046 0.00962857
R34945 DVSS.n5168 DVSS.n5048 0.00962857
R34946 DVSS.n5164 DVSS.n5048 0.00962857
R34947 DVSS.n5164 DVSS.n5162 0.00962857
R34948 DVSS.n5162 DVSS.n5160 0.00962857
R34949 DVSS.n5160 DVSS.n5050 0.00962857
R34950 DVSS.n5156 DVSS.n5050 0.00962857
R34951 DVSS.n5156 DVSS.n5052 0.00962857
R34952 DVSS.n5152 DVSS.n5052 0.00962857
R34953 DVSS.n5152 DVSS.n5054 0.00962857
R34954 DVSS.n5148 DVSS.n5054 0.00962857
R34955 DVSS.n5148 DVSS.n5056 0.00962857
R34956 DVSS.n5144 DVSS.n5056 0.00962857
R34957 DVSS.n5144 DVSS.n5058 0.00962857
R34958 DVSS.n5140 DVSS.n5058 0.00962857
R34959 DVSS.n5140 DVSS.n5060 0.00962857
R34960 DVSS.n5136 DVSS.n5060 0.00962857
R34961 DVSS.n5136 DVSS.n5062 0.00962857
R34962 DVSS.n5132 DVSS.n5062 0.00962857
R34963 DVSS.n5132 DVSS.n5064 0.00962857
R34964 DVSS.n5083 DVSS.n5064 0.00962857
R34965 DVSS.n5126 DVSS.n5083 0.00962857
R34966 DVSS.n5126 DVSS.n5084 0.00962857
R34967 DVSS.n5122 DVSS.n5084 0.00962857
R34968 DVSS.n5122 DVSS.n5087 0.00962857
R34969 DVSS.n5118 DVSS.n5087 0.00962857
R34970 DVSS.n5118 DVSS.n5089 0.00962857
R34971 DVSS.n5114 DVSS.n5089 0.00962857
R34972 DVSS.n5114 DVSS.n5112 0.00962857
R34973 DVSS.n5112 DVSS.n5111 0.00962857
R34974 DVSS.n5111 DVSS.n5091 0.00962857
R34975 DVSS.n5107 DVSS.n5091 0.00962857
R34976 DVSS.n5107 DVSS.n5103 0.00962857
R34977 DVSS.n5102 DVSS.n5093 0.00962857
R34978 DVSS.n5098 DVSS.n5093 0.00962857
R34979 DVSS.n5098 DVSS.n5096 0.00962857
R34980 DVSS.n3087 DVSS.n3074 0.00962857
R34981 DVSS.n3088 DVSS.n3087 0.00962857
R34982 DVSS.n3089 DVSS.n3088 0.00962857
R34983 DVSS.n3089 DVSS.n3056 0.00962857
R34984 DVSS.n5828 DVSS.n3069 0.00962857
R34985 DVSS.n5822 DVSS.n3069 0.00962857
R34986 DVSS.n5822 DVSS.n5821 0.00962857
R34987 DVSS.n5821 DVSS.n5820 0.00962857
R34988 DVSS.n5820 DVSS.n3096 0.00962857
R34989 DVSS.n5814 DVSS.n3096 0.00962857
R34990 DVSS.n5808 DVSS.n3119 0.00962857
R34991 DVSS.n5802 DVSS.n3119 0.00962857
R34992 DVSS.n5802 DVSS.n5801 0.00962857
R34993 DVSS.n5801 DVSS.n5800 0.00962857
R34994 DVSS.n5800 DVSS.n3128 0.00962857
R34995 DVSS.n5794 DVSS.n3128 0.00962857
R34996 DVSS.n5794 DVSS.n5793 0.00962857
R34997 DVSS.n5793 DVSS.n5792 0.00962857
R34998 DVSS.n5792 DVSS.n3132 0.00962857
R34999 DVSS.n5786 DVSS.n3132 0.00962857
R35000 DVSS.n5786 DVSS.n5785 0.00962857
R35001 DVSS.n5785 DVSS.n5784 0.00962857
R35002 DVSS.n5772 DVSS.n3158 0.00962857
R35003 DVSS.n5766 DVSS.n3158 0.00962857
R35004 DVSS.n5766 DVSS.n5765 0.00962857
R35005 DVSS.n5765 DVSS.n5764 0.00962857
R35006 DVSS.n5764 DVSS.n3162 0.00962857
R35007 DVSS.n5758 DVSS.n3162 0.00962857
R35008 DVSS.n5758 DVSS.n5757 0.00962857
R35009 DVSS.n5757 DVSS.n5756 0.00962857
R35010 DVSS.n5756 DVSS.n3166 0.00962857
R35011 DVSS.n5750 DVSS.n3166 0.00962857
R35012 DVSS.n5750 DVSS.n5749 0.00962857
R35013 DVSS.n5749 DVSS.n5748 0.00962857
R35014 DVSS.n5011 DVSS.n3181 0.00962857
R35015 DVSS.n5187 DVSS.n5038 0.00962857
R35016 DVSS.n5187 DVSS.n5186 0.00962857
R35017 DVSS.n5186 DVSS.n5185 0.00962857
R35018 DVSS.n5185 DVSS.n5039 0.00962857
R35019 DVSS.n5179 DVSS.n5039 0.00962857
R35020 DVSS.n5179 DVSS.n5178 0.00962857
R35021 DVSS.n5178 DVSS.n5177 0.00962857
R35022 DVSS.n5177 DVSS.n5043 0.00962857
R35023 DVSS.n5171 DVSS.n5043 0.00962857
R35024 DVSS.n5171 DVSS.n5170 0.00962857
R35025 DVSS.n5170 DVSS.n5169 0.00962857
R35026 DVSS.n5169 DVSS.n5047 0.00962857
R35027 DVSS.n5155 DVSS.n3332 0.00962857
R35028 DVSS.n5155 DVSS.n5154 0.00962857
R35029 DVSS.n5154 DVSS.n5153 0.00962857
R35030 DVSS.n5153 DVSS.n5053 0.00962857
R35031 DVSS.n5147 DVSS.n5053 0.00962857
R35032 DVSS.n5147 DVSS.n5146 0.00962857
R35033 DVSS.n5146 DVSS.n5145 0.00962857
R35034 DVSS.n5145 DVSS.n5057 0.00962857
R35035 DVSS.n5139 DVSS.n5057 0.00962857
R35036 DVSS.n5139 DVSS.n5138 0.00962857
R35037 DVSS.n5138 DVSS.n5137 0.00962857
R35038 DVSS.n5137 DVSS.n5061 0.00962857
R35039 DVSS.n5127 DVSS.n5082 0.00962857
R35040 DVSS.n5121 DVSS.n5082 0.00962857
R35041 DVSS.n5121 DVSS.n5120 0.00962857
R35042 DVSS.n5120 DVSS.n5119 0.00962857
R35043 DVSS.n5104 DVSS.n3376 0.00962857
R35044 DVSS.n5106 DVSS.n5104 0.00962857
R35045 DVSS.n5106 DVSS.n5105 0.00962857
R35046 DVSS.n5853 DVSS.n5852 0.00962857
R35047 DVSS.n5852 DVSS.n3036 0.00962857
R35048 DVSS.n5847 DVSS.n3036 0.00962857
R35049 DVSS.n5847 DVSS.n3038 0.00962857
R35050 DVSS.n5843 DVSS.n3038 0.00962857
R35051 DVSS.n5843 DVSS.n3040 0.00962857
R35052 DVSS.n5839 DVSS.n3040 0.00962857
R35053 DVSS.n5839 DVSS.n3042 0.00962857
R35054 DVSS.n3903 DVSS.n3042 0.00962857
R35055 DVSS.n3905 DVSS.n3903 0.00962857
R35056 DVSS.n3905 DVSS.n3901 0.00962857
R35057 DVSS.n3909 DVSS.n3901 0.00962857
R35058 DVSS.n3909 DVSS.n3899 0.00962857
R35059 DVSS.n3913 DVSS.n3899 0.00962857
R35060 DVSS.n3913 DVSS.n3895 0.00962857
R35061 DVSS.n4171 DVSS.n3895 0.00962857
R35062 DVSS.n4171 DVSS.n3897 0.00962857
R35063 DVSS.n4167 DVSS.n3897 0.00962857
R35064 DVSS.n4167 DVSS.n4165 0.00962857
R35065 DVSS.n4165 DVSS.n3917 0.00962857
R35066 DVSS.n4161 DVSS.n3917 0.00962857
R35067 DVSS.n4161 DVSS.n3919 0.00962857
R35068 DVSS.n4157 DVSS.n3919 0.00962857
R35069 DVSS.n4157 DVSS.n3922 0.00962857
R35070 DVSS.n4153 DVSS.n3922 0.00962857
R35071 DVSS.n4153 DVSS.n3924 0.00962857
R35072 DVSS.n4149 DVSS.n3924 0.00962857
R35073 DVSS.n4149 DVSS.n3926 0.00962857
R35074 DVSS.n4145 DVSS.n3926 0.00962857
R35075 DVSS.n4145 DVSS.n3928 0.00962857
R35076 DVSS.n4141 DVSS.n3928 0.00962857
R35077 DVSS.n4141 DVSS.n3930 0.00962857
R35078 DVSS.n3951 DVSS.n3930 0.00962857
R35079 DVSS.n4135 DVSS.n3951 0.00962857
R35080 DVSS.n4135 DVSS.n3952 0.00962857
R35081 DVSS.n4131 DVSS.n3952 0.00962857
R35082 DVSS.n4131 DVSS.n3955 0.00962857
R35083 DVSS.n4127 DVSS.n3955 0.00962857
R35084 DVSS.n4127 DVSS.n3958 0.00962857
R35085 DVSS.n4123 DVSS.n3958 0.00962857
R35086 DVSS.n4123 DVSS.n3960 0.00962857
R35087 DVSS.n4119 DVSS.n3960 0.00962857
R35088 DVSS.n4119 DVSS.n3962 0.00962857
R35089 DVSS.n4115 DVSS.n3962 0.00962857
R35090 DVSS.n4115 DVSS.n3964 0.00962857
R35091 DVSS.n4111 DVSS.n3964 0.00962857
R35092 DVSS.n4111 DVSS.n3966 0.00962857
R35093 DVSS.n4107 DVSS.n3966 0.00962857
R35094 DVSS.n4107 DVSS.n3968 0.00962857
R35095 DVSS.n3996 DVSS.n3968 0.00962857
R35096 DVSS.n3996 DVSS.n3473 0.00962857
R35097 DVSS.n5239 DVSS.n3473 0.00962857
R35098 DVSS.n5239 DVSS.n3471 0.00962857
R35099 DVSS.n5243 DVSS.n3471 0.00962857
R35100 DVSS.n5243 DVSS.n3469 0.00962857
R35101 DVSS.n5247 DVSS.n3469 0.00962857
R35102 DVSS.n5247 DVSS.n3467 0.00962857
R35103 DVSS.n5251 DVSS.n3467 0.00962857
R35104 DVSS.n5251 DVSS.n3465 0.00962857
R35105 DVSS.n5255 DVSS.n3465 0.00962857
R35106 DVSS.n5255 DVSS.n3463 0.00962857
R35107 DVSS.n5259 DVSS.n3463 0.00962857
R35108 DVSS.n5259 DVSS.n3461 0.00962857
R35109 DVSS.n5263 DVSS.n3461 0.00962857
R35110 DVSS.n5263 DVSS.n3459 0.00962857
R35111 DVSS.n5267 DVSS.n3459 0.00962857
R35112 DVSS.n5267 DVSS.n3439 0.00962857
R35113 DVSS.n5274 DVSS.n3439 0.00962857
R35114 DVSS.n5274 DVSS.n3437 0.00962857
R35115 DVSS.n5278 DVSS.n3437 0.00962857
R35116 DVSS.n5278 DVSS.n3435 0.00962857
R35117 DVSS.n5282 DVSS.n3435 0.00962857
R35118 DVSS.n5282 DVSS.n3433 0.00962857
R35119 DVSS.n5286 DVSS.n3433 0.00962857
R35120 DVSS.n5286 DVSS.n3431 0.00962857
R35121 DVSS.n5290 DVSS.n3431 0.00962857
R35122 DVSS.n5290 DVSS.n3429 0.00962857
R35123 DVSS.n5294 DVSS.n3429 0.00962857
R35124 DVSS.n5294 DVSS.n3427 0.00962857
R35125 DVSS.n5298 DVSS.n3427 0.00962857
R35126 DVSS.n5298 DVSS.n3425 0.00962857
R35127 DVSS.n5302 DVSS.n3425 0.00962857
R35128 DVSS.n5302 DVSS.n3404 0.00962857
R35129 DVSS.n5309 DVSS.n3404 0.00962857
R35130 DVSS.n5309 DVSS.n3402 0.00962857
R35131 DVSS.n5313 DVSS.n3402 0.00962857
R35132 DVSS.n5313 DVSS.n3400 0.00962857
R35133 DVSS.n5318 DVSS.n3400 0.00962857
R35134 DVSS.n5318 DVSS.n3398 0.00962857
R35135 DVSS.n5322 DVSS.n3398 0.00962857
R35136 DVSS.n5323 DVSS.n5322 0.00962857
R35137 DVSS.n5325 DVSS.n5323 0.00962857
R35138 DVSS.n5325 DVSS.n3395 0.00962857
R35139 DVSS.n5346 DVSS.n3395 0.00962857
R35140 DVSS.n5346 DVSS.n3396 0.00962857
R35141 DVSS.n5342 DVSS.n3396 0.00962857
R35142 DVSS.n5342 DVSS.n5339 0.00962857
R35143 DVSS.n5338 DVSS.n5329 0.00962857
R35144 DVSS.n5334 DVSS.n5329 0.00962857
R35145 DVSS.n5334 DVSS.n5332 0.00962857
R35146 DVSS.n5846 DVSS.n5845 0.00962857
R35147 DVSS.n5845 DVSS.n5844 0.00962857
R35148 DVSS.n5844 DVSS.n3039 0.00962857
R35149 DVSS.n5838 DVSS.n3039 0.00962857
R35150 DVSS.n3904 DVSS.n3054 0.00962857
R35151 DVSS.n3904 DVSS.n3900 0.00962857
R35152 DVSS.n3910 DVSS.n3900 0.00962857
R35153 DVSS.n3911 DVSS.n3910 0.00962857
R35154 DVSS.n3912 DVSS.n3911 0.00962857
R35155 DVSS.n3912 DVSS.n3890 0.00962857
R35156 DVSS.n4164 DVSS.n4163 0.00962857
R35157 DVSS.n4163 DVSS.n4162 0.00962857
R35158 DVSS.n4162 DVSS.n3918 0.00962857
R35159 DVSS.n4156 DVSS.n3918 0.00962857
R35160 DVSS.n4156 DVSS.n4155 0.00962857
R35161 DVSS.n4155 DVSS.n4154 0.00962857
R35162 DVSS.n4154 DVSS.n3923 0.00962857
R35163 DVSS.n4148 DVSS.n3923 0.00962857
R35164 DVSS.n4148 DVSS.n4147 0.00962857
R35165 DVSS.n4147 DVSS.n4146 0.00962857
R35166 DVSS.n4146 DVSS.n3927 0.00962857
R35167 DVSS.n4140 DVSS.n3927 0.00962857
R35168 DVSS.n4130 DVSS.n3956 0.00962857
R35169 DVSS.n4130 DVSS.n4129 0.00962857
R35170 DVSS.n4129 DVSS.n4128 0.00962857
R35171 DVSS.n4128 DVSS.n3957 0.00962857
R35172 DVSS.n4122 DVSS.n3957 0.00962857
R35173 DVSS.n4122 DVSS.n4121 0.00962857
R35174 DVSS.n4121 DVSS.n4120 0.00962857
R35175 DVSS.n4120 DVSS.n3961 0.00962857
R35176 DVSS.n4114 DVSS.n3961 0.00962857
R35177 DVSS.n4114 DVSS.n4113 0.00962857
R35178 DVSS.n4113 DVSS.n4112 0.00962857
R35179 DVSS.n4112 DVSS.n3965 0.00962857
R35180 DVSS.n3997 DVSS.n3994 0.00962857
R35181 DVSS.n5245 DVSS.n5244 0.00962857
R35182 DVSS.n5246 DVSS.n5245 0.00962857
R35183 DVSS.n5246 DVSS.n3466 0.00962857
R35184 DVSS.n5252 DVSS.n3466 0.00962857
R35185 DVSS.n5253 DVSS.n5252 0.00962857
R35186 DVSS.n5254 DVSS.n5253 0.00962857
R35187 DVSS.n5254 DVSS.n3462 0.00962857
R35188 DVSS.n5260 DVSS.n3462 0.00962857
R35189 DVSS.n5261 DVSS.n5260 0.00962857
R35190 DVSS.n5262 DVSS.n5261 0.00962857
R35191 DVSS.n5262 DVSS.n3458 0.00962857
R35192 DVSS.n5268 DVSS.n3458 0.00962857
R35193 DVSS.n5280 DVSS.n5279 0.00962857
R35194 DVSS.n5281 DVSS.n5280 0.00962857
R35195 DVSS.n5281 DVSS.n3432 0.00962857
R35196 DVSS.n5287 DVSS.n3432 0.00962857
R35197 DVSS.n5288 DVSS.n5287 0.00962857
R35198 DVSS.n5289 DVSS.n5288 0.00962857
R35199 DVSS.n5289 DVSS.n3428 0.00962857
R35200 DVSS.n5295 DVSS.n3428 0.00962857
R35201 DVSS.n5296 DVSS.n5295 0.00962857
R35202 DVSS.n5297 DVSS.n5296 0.00962857
R35203 DVSS.n5297 DVSS.n3424 0.00962857
R35204 DVSS.n5303 DVSS.n3424 0.00962857
R35205 DVSS.n5315 DVSS.n5314 0.00962857
R35206 DVSS.n5317 DVSS.n5315 0.00962857
R35207 DVSS.n5317 DVSS.n5316 0.00962857
R35208 DVSS.n5316 DVSS.n3380 0.00962857
R35209 DVSS.n5347 DVSS.n3394 0.00962857
R35210 DVSS.n5341 DVSS.n3394 0.00962857
R35211 DVSS.n5341 DVSS.n5340 0.00962857
R35212 DVSS.n4244 DVSS.n4232 0.00962857
R35213 DVSS.n4245 DVSS.n4244 0.00962857
R35214 DVSS.n4246 DVSS.n4245 0.00962857
R35215 DVSS.n4246 DVSS.n4224 0.00962857
R35216 DVSS.n4267 DVSS.n4211 0.00962857
R35217 DVSS.n4268 DVSS.n4267 0.00962857
R35218 DVSS.n4269 DVSS.n4268 0.00962857
R35219 DVSS.n4269 DVSS.n4202 0.00962857
R35220 DVSS.n4410 DVSS.n4409 0.00962857
R35221 DVSS.n4409 DVSS.n4408 0.00962857
R35222 DVSS.n4408 DVSS.n4275 0.00962857
R35223 DVSS.n4402 DVSS.n4275 0.00962857
R35224 DVSS.n4402 DVSS.n4401 0.00962857
R35225 DVSS.n4401 DVSS.n4400 0.00962857
R35226 DVSS.n4400 DVSS.n4280 0.00962857
R35227 DVSS.n4394 DVSS.n4280 0.00962857
R35228 DVSS.n4394 DVSS.n4393 0.00962857
R35229 DVSS.n4393 DVSS.n4392 0.00962857
R35230 DVSS.n4392 DVSS.n4284 0.00962857
R35231 DVSS.n4284 DVSS.n3722 0.00962857
R35232 DVSS.n4379 DVSS.n4378 0.00962857
R35233 DVSS.n4378 DVSS.n4377 0.00962857
R35234 DVSS.n4377 DVSS.n4291 0.00962857
R35235 DVSS.n4371 DVSS.n4291 0.00962857
R35236 DVSS.n4371 DVSS.n4370 0.00962857
R35237 DVSS.n4370 DVSS.n4369 0.00962857
R35238 DVSS.n4369 DVSS.n4295 0.00962857
R35239 DVSS.n4363 DVSS.n4295 0.00962857
R35240 DVSS.n4363 DVSS.n4362 0.00962857
R35241 DVSS.n4362 DVSS.n4361 0.00962857
R35242 DVSS.n4361 DVSS.n4299 0.00962857
R35243 DVSS.n4299 DVSS.n3691 0.00962857
R35244 DVSS.n4302 DVSS.n3679 0.00962857
R35245 DVSS.n4341 DVSS.n4308 0.00962857
R35246 DVSS.n4341 DVSS.n4340 0.00962857
R35247 DVSS.n4340 DVSS.n4339 0.00962857
R35248 DVSS.n4339 DVSS.n4309 0.00962857
R35249 DVSS.n4333 DVSS.n4309 0.00962857
R35250 DVSS.n4333 DVSS.n4332 0.00962857
R35251 DVSS.n4332 DVSS.n4331 0.00962857
R35252 DVSS.n4331 DVSS.n4313 0.00962857
R35253 DVSS.n4325 DVSS.n4313 0.00962857
R35254 DVSS.n4325 DVSS.n4324 0.00962857
R35255 DVSS.n4324 DVSS.n4323 0.00962857
R35256 DVSS.n4323 DVSS.n3656 0.00962857
R35257 DVSS.n4857 DVSS.n3643 0.00962857
R35258 DVSS.n4858 DVSS.n4857 0.00962857
R35259 DVSS.n4859 DVSS.n4858 0.00962857
R35260 DVSS.n4859 DVSS.n3639 0.00962857
R35261 DVSS.n4865 DVSS.n3639 0.00962857
R35262 DVSS.n4866 DVSS.n4865 0.00962857
R35263 DVSS.n4867 DVSS.n4866 0.00962857
R35264 DVSS.n4867 DVSS.n3635 0.00962857
R35265 DVSS.n4873 DVSS.n3635 0.00962857
R35266 DVSS.n4874 DVSS.n4873 0.00962857
R35267 DVSS.n4875 DVSS.n4874 0.00962857
R35268 DVSS.n4875 DVSS.n3627 0.00962857
R35269 DVSS.n4895 DVSS.n3610 0.00962857
R35270 DVSS.n4896 DVSS.n4895 0.00962857
R35271 DVSS.n4897 DVSS.n4896 0.00962857
R35272 DVSS.n4897 DVSS.n3601 0.00962857
R35273 DVSS.n4953 DVSS.n4952 0.00962857
R35274 DVSS.n4952 DVSS.n4951 0.00962857
R35275 DVSS.n4951 DVSS.n4903 0.00962857
R35276 DVSS.n6639 DVSS.n6638 0.00962857
R35277 DVSS.n6638 DVSS.n6020 0.00962857
R35278 DVSS.n6634 DVSS.n6020 0.00962857
R35279 DVSS.n6634 DVSS.n6022 0.00962857
R35280 DVSS.n6630 DVSS.n6022 0.00962857
R35281 DVSS.n6630 DVSS.n6025 0.00962857
R35282 DVSS.n6626 DVSS.n6025 0.00962857
R35283 DVSS.n6626 DVSS.n6027 0.00962857
R35284 DVSS.n6622 DVSS.n6027 0.00962857
R35285 DVSS.n6622 DVSS.n6029 0.00962857
R35286 DVSS.n6618 DVSS.n6029 0.00962857
R35287 DVSS.n6618 DVSS.n6031 0.00962857
R35288 DVSS.n6614 DVSS.n6031 0.00962857
R35289 DVSS.n6614 DVSS.n6349 0.00962857
R35290 DVSS.n6610 DVSS.n6349 0.00962857
R35291 DVSS.n6610 DVSS.n6351 0.00962857
R35292 DVSS.n6606 DVSS.n6351 0.00962857
R35293 DVSS.n6606 DVSS.n6353 0.00962857
R35294 DVSS.n6602 DVSS.n6353 0.00962857
R35295 DVSS.n6602 DVSS.n6355 0.00962857
R35296 DVSS.n6598 DVSS.n6355 0.00962857
R35297 DVSS.n6598 DVSS.n6357 0.00962857
R35298 DVSS.n6594 DVSS.n6357 0.00962857
R35299 DVSS.n6594 DVSS.n6359 0.00962857
R35300 DVSS.n6590 DVSS.n6359 0.00962857
R35301 DVSS.n6590 DVSS.n6361 0.00962857
R35302 DVSS.n6586 DVSS.n6361 0.00962857
R35303 DVSS.n6586 DVSS.n6363 0.00962857
R35304 DVSS.n6582 DVSS.n6363 0.00962857
R35305 DVSS.n6582 DVSS.n6365 0.00962857
R35306 DVSS.n6578 DVSS.n6365 0.00962857
R35307 DVSS.n6578 DVSS.n6367 0.00962857
R35308 DVSS.n6574 DVSS.n6367 0.00962857
R35309 DVSS.n6574 DVSS.n6369 0.00962857
R35310 DVSS.n6570 DVSS.n6369 0.00962857
R35311 DVSS.n6570 DVSS.n6371 0.00962857
R35312 DVSS.n6566 DVSS.n6371 0.00962857
R35313 DVSS.n6566 DVSS.n6373 0.00962857
R35314 DVSS.n6562 DVSS.n6373 0.00962857
R35315 DVSS.n6562 DVSS.n6375 0.00962857
R35316 DVSS.n6558 DVSS.n6375 0.00962857
R35317 DVSS.n6558 DVSS.n6377 0.00962857
R35318 DVSS.n6554 DVSS.n6377 0.00962857
R35319 DVSS.n6554 DVSS.n6379 0.00962857
R35320 DVSS.n6550 DVSS.n6379 0.00962857
R35321 DVSS.n6550 DVSS.n6381 0.00962857
R35322 DVSS.n6546 DVSS.n6381 0.00962857
R35323 DVSS.n6546 DVSS.n6383 0.00962857
R35324 DVSS.n6542 DVSS.n6383 0.00962857
R35325 DVSS.n6542 DVSS.n6385 0.00962857
R35326 DVSS.n6538 DVSS.n6385 0.00962857
R35327 DVSS.n6538 DVSS.n6387 0.00962857
R35328 DVSS.n6534 DVSS.n6387 0.00962857
R35329 DVSS.n6534 DVSS.n6389 0.00962857
R35330 DVSS.n6530 DVSS.n6389 0.00962857
R35331 DVSS.n6530 DVSS.n6391 0.00962857
R35332 DVSS.n6526 DVSS.n6391 0.00962857
R35333 DVSS.n6526 DVSS.n6393 0.00962857
R35334 DVSS.n6522 DVSS.n6393 0.00962857
R35335 DVSS.n6522 DVSS.n6395 0.00962857
R35336 DVSS.n6518 DVSS.n6395 0.00962857
R35337 DVSS.n6518 DVSS.n6397 0.00962857
R35338 DVSS.n6514 DVSS.n6397 0.00962857
R35339 DVSS.n6514 DVSS.n6399 0.00962857
R35340 DVSS.n6510 DVSS.n6399 0.00962857
R35341 DVSS.n6510 DVSS.n6401 0.00962857
R35342 DVSS.n6506 DVSS.n6401 0.00962857
R35343 DVSS.n6506 DVSS.n6403 0.00962857
R35344 DVSS.n6502 DVSS.n6403 0.00962857
R35345 DVSS.n6502 DVSS.n6405 0.00962857
R35346 DVSS.n6498 DVSS.n6405 0.00962857
R35347 DVSS.n6498 DVSS.n6407 0.00962857
R35348 DVSS.n6494 DVSS.n6407 0.00962857
R35349 DVSS.n6494 DVSS.n6409 0.00962857
R35350 DVSS.n6490 DVSS.n6409 0.00962857
R35351 DVSS.n6490 DVSS.n6411 0.00962857
R35352 DVSS.n6486 DVSS.n6411 0.00962857
R35353 DVSS.n6486 DVSS.n6413 0.00962857
R35354 DVSS.n6482 DVSS.n6413 0.00962857
R35355 DVSS.n6482 DVSS.n6415 0.00962857
R35356 DVSS.n6478 DVSS.n6415 0.00962857
R35357 DVSS.n6478 DVSS.n6417 0.00962857
R35358 DVSS.n6474 DVSS.n6417 0.00962857
R35359 DVSS.n6474 DVSS.n6419 0.00962857
R35360 DVSS.n6470 DVSS.n6419 0.00962857
R35361 DVSS.n6470 DVSS.n6421 0.00962857
R35362 DVSS.n6466 DVSS.n6421 0.00962857
R35363 DVSS.n6466 DVSS.n6423 0.00962857
R35364 DVSS.n6462 DVSS.n6423 0.00962857
R35365 DVSS.n6462 DVSS.n6425 0.00962857
R35366 DVSS.n6458 DVSS.n6425 0.00962857
R35367 DVSS.n6458 DVSS.n6427 0.00962857
R35368 DVSS.n6454 DVSS.n6427 0.00962857
R35369 DVSS.n6454 DVSS.n6429 0.00962857
R35370 DVSS.n6450 DVSS.n6429 0.00962857
R35371 DVSS.n6450 DVSS.n6431 0.00962857
R35372 DVSS.n6446 DVSS.n6431 0.00962857
R35373 DVSS.n6443 DVSS.n6432 0.00962857
R35374 DVSS.n6439 DVSS.n6432 0.00962857
R35375 DVSS.n6439 DVSS.n6434 0.00962857
R35376 DVSS.n6047 DVSS.n6044 0.00962857
R35377 DVSS.n6051 DVSS.n6044 0.00962857
R35378 DVSS.n6051 DVSS.n6042 0.00962857
R35379 DVSS.n6055 DVSS.n6042 0.00962857
R35380 DVSS.n6055 DVSS.n6040 0.00962857
R35381 DVSS.n6059 DVSS.n6040 0.00962857
R35382 DVSS.n6059 DVSS.n6038 0.00962857
R35383 DVSS.n6063 DVSS.n6038 0.00962857
R35384 DVSS.n6063 DVSS.n6035 0.00962857
R35385 DVSS.n6342 DVSS.n6035 0.00962857
R35386 DVSS.n6342 DVSS.n6036 0.00962857
R35387 DVSS.n6338 DVSS.n6036 0.00962857
R35388 DVSS.n6338 DVSS.n6067 0.00962857
R35389 DVSS.n6334 DVSS.n6067 0.00962857
R35390 DVSS.n6334 DVSS.n6070 0.00962857
R35391 DVSS.n6330 DVSS.n6070 0.00962857
R35392 DVSS.n6330 DVSS.n6072 0.00962857
R35393 DVSS.n6326 DVSS.n6072 0.00962857
R35394 DVSS.n6326 DVSS.n6074 0.00962857
R35395 DVSS.n6322 DVSS.n6074 0.00962857
R35396 DVSS.n6322 DVSS.n6076 0.00962857
R35397 DVSS.n6318 DVSS.n6076 0.00962857
R35398 DVSS.n6318 DVSS.n6078 0.00962857
R35399 DVSS.n6314 DVSS.n6078 0.00962857
R35400 DVSS.n6314 DVSS.n6080 0.00962857
R35401 DVSS.n6310 DVSS.n6080 0.00962857
R35402 DVSS.n6310 DVSS.n6082 0.00962857
R35403 DVSS.n6306 DVSS.n6082 0.00962857
R35404 DVSS.n6306 DVSS.n6084 0.00962857
R35405 DVSS.n6302 DVSS.n6084 0.00962857
R35406 DVSS.n6302 DVSS.n6086 0.00962857
R35407 DVSS.n6298 DVSS.n6086 0.00962857
R35408 DVSS.n6298 DVSS.n6088 0.00962857
R35409 DVSS.n6294 DVSS.n6088 0.00962857
R35410 DVSS.n6294 DVSS.n6090 0.00962857
R35411 DVSS.n6290 DVSS.n6090 0.00962857
R35412 DVSS.n6290 DVSS.n6092 0.00962857
R35413 DVSS.n6286 DVSS.n6092 0.00962857
R35414 DVSS.n6286 DVSS.n6094 0.00962857
R35415 DVSS.n6282 DVSS.n6094 0.00962857
R35416 DVSS.n6282 DVSS.n6096 0.00962857
R35417 DVSS.n6278 DVSS.n6096 0.00962857
R35418 DVSS.n6278 DVSS.n6098 0.00962857
R35419 DVSS.n6274 DVSS.n6098 0.00962857
R35420 DVSS.n6274 DVSS.n6100 0.00962857
R35421 DVSS.n6270 DVSS.n6100 0.00962857
R35422 DVSS.n6270 DVSS.n6102 0.00962857
R35423 DVSS.n6266 DVSS.n6102 0.00962857
R35424 DVSS.n6266 DVSS.n6104 0.00962857
R35425 DVSS.n6262 DVSS.n6104 0.00962857
R35426 DVSS.n6262 DVSS.n6106 0.00962857
R35427 DVSS.n6258 DVSS.n6106 0.00962857
R35428 DVSS.n6258 DVSS.n6108 0.00962857
R35429 DVSS.n6254 DVSS.n6108 0.00962857
R35430 DVSS.n6254 DVSS.n6110 0.00962857
R35431 DVSS.n6250 DVSS.n6110 0.00962857
R35432 DVSS.n6250 DVSS.n6112 0.00962857
R35433 DVSS.n6246 DVSS.n6112 0.00962857
R35434 DVSS.n6246 DVSS.n6114 0.00962857
R35435 DVSS.n6242 DVSS.n6114 0.00962857
R35436 DVSS.n6242 DVSS.n6116 0.00962857
R35437 DVSS.n6238 DVSS.n6116 0.00962857
R35438 DVSS.n6238 DVSS.n6118 0.00962857
R35439 DVSS.n6234 DVSS.n6118 0.00962857
R35440 DVSS.n6234 DVSS.n6120 0.00962857
R35441 DVSS.n6230 DVSS.n6120 0.00962857
R35442 DVSS.n6230 DVSS.n6122 0.00962857
R35443 DVSS.n6226 DVSS.n6122 0.00962857
R35444 DVSS.n6226 DVSS.n6124 0.00962857
R35445 DVSS.n6222 DVSS.n6124 0.00962857
R35446 DVSS.n6222 DVSS.n6126 0.00962857
R35447 DVSS.n6218 DVSS.n6126 0.00962857
R35448 DVSS.n6218 DVSS.n6128 0.00962857
R35449 DVSS.n6214 DVSS.n6128 0.00962857
R35450 DVSS.n6214 DVSS.n6130 0.00962857
R35451 DVSS.n6210 DVSS.n6130 0.00962857
R35452 DVSS.n6210 DVSS.n6132 0.00962857
R35453 DVSS.n6206 DVSS.n6132 0.00962857
R35454 DVSS.n6206 DVSS.n6134 0.00962857
R35455 DVSS.n6202 DVSS.n6134 0.00962857
R35456 DVSS.n6202 DVSS.n6136 0.00962857
R35457 DVSS.n6198 DVSS.n6136 0.00962857
R35458 DVSS.n6198 DVSS.n6138 0.00962857
R35459 DVSS.n6194 DVSS.n6138 0.00962857
R35460 DVSS.n6194 DVSS.n6140 0.00962857
R35461 DVSS.n6190 DVSS.n6140 0.00962857
R35462 DVSS.n6190 DVSS.n6142 0.00962857
R35463 DVSS.n6186 DVSS.n6142 0.00962857
R35464 DVSS.n6186 DVSS.n6144 0.00962857
R35465 DVSS.n6182 DVSS.n6144 0.00962857
R35466 DVSS.n6182 DVSS.n6146 0.00962857
R35467 DVSS.n6178 DVSS.n6146 0.00962857
R35468 DVSS.n6178 DVSS.n6148 0.00962857
R35469 DVSS.n6174 DVSS.n6148 0.00962857
R35470 DVSS.n6174 DVSS.n6150 0.00962857
R35471 DVSS.n6170 DVSS.n6150 0.00962857
R35472 DVSS.n6170 DVSS.n6152 0.00962857
R35473 DVSS.n6166 DVSS.n6154 0.00962857
R35474 DVSS.n6162 DVSS.n6154 0.00962857
R35475 DVSS.n6162 DVSS.n6156 0.00962857
R35476 DVSS.n6046 DVSS.n6045 0.00962857
R35477 DVSS.n6046 DVSS.n6043 0.00962857
R35478 DVSS.n6052 DVSS.n6043 0.00962857
R35479 DVSS.n6053 DVSS.n6052 0.00962857
R35480 DVSS.n6054 DVSS.n6053 0.00962857
R35481 DVSS.n6054 DVSS.n6039 0.00962857
R35482 DVSS.n6060 DVSS.n6039 0.00962857
R35483 DVSS.n6061 DVSS.n6060 0.00962857
R35484 DVSS.n6062 DVSS.n6061 0.00962857
R35485 DVSS.n6062 DVSS.n6034 0.00962857
R35486 DVSS.n6337 DVSS.n6068 0.00962857
R35487 DVSS.n6337 DVSS.n6336 0.00962857
R35488 DVSS.n6336 DVSS.n6335 0.00962857
R35489 DVSS.n6335 DVSS.n6069 0.00962857
R35490 DVSS.n6329 DVSS.n6069 0.00962857
R35491 DVSS.n6329 DVSS.n6328 0.00962857
R35492 DVSS.n6328 DVSS.n6327 0.00962857
R35493 DVSS.n6327 DVSS.n6073 0.00962857
R35494 DVSS.n6321 DVSS.n6073 0.00962857
R35495 DVSS.n6321 DVSS.n6320 0.00962857
R35496 DVSS.n6320 DVSS.n6319 0.00962857
R35497 DVSS.n6319 DVSS.n6077 0.00962857
R35498 DVSS.n6313 DVSS.n6077 0.00962857
R35499 DVSS.n6313 DVSS.n6312 0.00962857
R35500 DVSS.n6312 DVSS.n6311 0.00962857
R35501 DVSS.n6311 DVSS.n6081 0.00962857
R35502 DVSS.n6305 DVSS.n6081 0.00962857
R35503 DVSS.n6305 DVSS.n6304 0.00962857
R35504 DVSS.n6304 DVSS.n6303 0.00962857
R35505 DVSS.n6303 DVSS.n6085 0.00962857
R35506 DVSS.n6297 DVSS.n6085 0.00962857
R35507 DVSS.n6297 DVSS.n6296 0.00962857
R35508 DVSS.n6296 DVSS.n6295 0.00962857
R35509 DVSS.n6295 DVSS.n6089 0.00962857
R35510 DVSS.n6289 DVSS.n6089 0.00962857
R35511 DVSS.n6289 DVSS.n6288 0.00962857
R35512 DVSS.n6288 DVSS.n6287 0.00962857
R35513 DVSS.n6287 DVSS.n6093 0.00962857
R35514 DVSS.n6281 DVSS.n6093 0.00962857
R35515 DVSS.n6281 DVSS.n6280 0.00962857
R35516 DVSS.n6280 DVSS.n6279 0.00962857
R35517 DVSS.n6279 DVSS.n6097 0.00962857
R35518 DVSS.n6273 DVSS.n6097 0.00962857
R35519 DVSS.n6273 DVSS.n6272 0.00962857
R35520 DVSS.n6272 DVSS.n6271 0.00962857
R35521 DVSS.n6271 DVSS.n6101 0.00962857
R35522 DVSS.n6265 DVSS.n6101 0.00962857
R35523 DVSS.n6265 DVSS.n6264 0.00962857
R35524 DVSS.n6264 DVSS.n6263 0.00962857
R35525 DVSS.n6263 DVSS.n6105 0.00962857
R35526 DVSS.n6257 DVSS.n6105 0.00962857
R35527 DVSS.n6257 DVSS.n6256 0.00962857
R35528 DVSS.n6256 DVSS.n6255 0.00962857
R35529 DVSS.n6255 DVSS.n6109 0.00962857
R35530 DVSS.n6249 DVSS.n6109 0.00962857
R35531 DVSS.n6249 DVSS.n6248 0.00962857
R35532 DVSS.n6248 DVSS.n6247 0.00962857
R35533 DVSS.n6247 DVSS.n6113 0.00962857
R35534 DVSS.n6241 DVSS.n6113 0.00962857
R35535 DVSS.n6241 DVSS.n6240 0.00962857
R35536 DVSS.n6240 DVSS.n6239 0.00962857
R35537 DVSS.n6239 DVSS.n6117 0.00962857
R35538 DVSS.n6233 DVSS.n6117 0.00962857
R35539 DVSS.n6233 DVSS.n6232 0.00962857
R35540 DVSS.n6232 DVSS.n6231 0.00962857
R35541 DVSS.n6231 DVSS.n6121 0.00962857
R35542 DVSS.n6225 DVSS.n6121 0.00962857
R35543 DVSS.n6225 DVSS.n6224 0.00962857
R35544 DVSS.n6224 DVSS.n6223 0.00962857
R35545 DVSS.n6223 DVSS.n6125 0.00962857
R35546 DVSS.n6217 DVSS.n6125 0.00962857
R35547 DVSS.n6217 DVSS.n6216 0.00962857
R35548 DVSS.n6216 DVSS.n6215 0.00962857
R35549 DVSS.n6215 DVSS.n6129 0.00962857
R35550 DVSS.n6209 DVSS.n6129 0.00962857
R35551 DVSS.n6209 DVSS.n6208 0.00962857
R35552 DVSS.n6208 DVSS.n6207 0.00962857
R35553 DVSS.n6207 DVSS.n6133 0.00962857
R35554 DVSS.n6201 DVSS.n6133 0.00962857
R35555 DVSS.n6201 DVSS.n6200 0.00962857
R35556 DVSS.n6200 DVSS.n6199 0.00962857
R35557 DVSS.n6199 DVSS.n6137 0.00962857
R35558 DVSS.n6193 DVSS.n6137 0.00962857
R35559 DVSS.n6193 DVSS.n6192 0.00962857
R35560 DVSS.n6192 DVSS.n6191 0.00962857
R35561 DVSS.n6191 DVSS.n6141 0.00962857
R35562 DVSS.n6185 DVSS.n6141 0.00962857
R35563 DVSS.n6185 DVSS.n6184 0.00962857
R35564 DVSS.n6184 DVSS.n6183 0.00962857
R35565 DVSS.n6183 DVSS.n6145 0.00962857
R35566 DVSS.n6177 DVSS.n6145 0.00962857
R35567 DVSS.n6177 DVSS.n6176 0.00962857
R35568 DVSS.n6176 DVSS.n6175 0.00962857
R35569 DVSS.n6175 DVSS.n6149 0.00962857
R35570 DVSS.n6169 DVSS.n6149 0.00962857
R35571 DVSS.n6169 DVSS.n6168 0.00962857
R35572 DVSS.n6167 DVSS.n6153 0.00962857
R35573 DVSS.n6161 DVSS.n6153 0.00962857
R35574 DVSS.n6161 DVSS.n6160 0.00962857
R35575 DVSS.n6160 DVSS.n6159 0.00962857
R35576 DVSS.n6641 DVSS.n6640 0.00962857
R35577 DVSS.n6640 DVSS.n6019 0.00962857
R35578 DVSS.n6023 DVSS.n6019 0.00962857
R35579 DVSS.n6633 DVSS.n6023 0.00962857
R35580 DVSS.n6633 DVSS.n6632 0.00962857
R35581 DVSS.n6632 DVSS.n6631 0.00962857
R35582 DVSS.n6631 DVSS.n6024 0.00962857
R35583 DVSS.n6625 DVSS.n6024 0.00962857
R35584 DVSS.n6625 DVSS.n6624 0.00962857
R35585 DVSS.n6624 DVSS.n6623 0.00962857
R35586 DVSS.n6617 DVSS.n6616 0.00962857
R35587 DVSS.n6616 DVSS.n6615 0.00962857
R35588 DVSS.n6615 DVSS.n6348 0.00962857
R35589 DVSS.n6609 DVSS.n6348 0.00962857
R35590 DVSS.n6609 DVSS.n6608 0.00962857
R35591 DVSS.n6608 DVSS.n6607 0.00962857
R35592 DVSS.n6607 DVSS.n6352 0.00962857
R35593 DVSS.n6601 DVSS.n6352 0.00962857
R35594 DVSS.n6601 DVSS.n6600 0.00962857
R35595 DVSS.n6600 DVSS.n6599 0.00962857
R35596 DVSS.n6599 DVSS.n6356 0.00962857
R35597 DVSS.n6593 DVSS.n6356 0.00962857
R35598 DVSS.n6593 DVSS.n6592 0.00962857
R35599 DVSS.n6592 DVSS.n6591 0.00962857
R35600 DVSS.n6591 DVSS.n6360 0.00962857
R35601 DVSS.n6585 DVSS.n6360 0.00962857
R35602 DVSS.n6585 DVSS.n6584 0.00962857
R35603 DVSS.n6584 DVSS.n6583 0.00962857
R35604 DVSS.n6583 DVSS.n6364 0.00962857
R35605 DVSS.n6577 DVSS.n6364 0.00962857
R35606 DVSS.n6577 DVSS.n6576 0.00962857
R35607 DVSS.n6576 DVSS.n6575 0.00962857
R35608 DVSS.n6575 DVSS.n6368 0.00962857
R35609 DVSS.n6569 DVSS.n6368 0.00962857
R35610 DVSS.n6569 DVSS.n6568 0.00962857
R35611 DVSS.n6568 DVSS.n6567 0.00962857
R35612 DVSS.n6567 DVSS.n6372 0.00962857
R35613 DVSS.n6561 DVSS.n6372 0.00962857
R35614 DVSS.n6561 DVSS.n6560 0.00962857
R35615 DVSS.n6560 DVSS.n6559 0.00962857
R35616 DVSS.n6559 DVSS.n6376 0.00962857
R35617 DVSS.n6553 DVSS.n6376 0.00962857
R35618 DVSS.n6553 DVSS.n6552 0.00962857
R35619 DVSS.n6552 DVSS.n6551 0.00962857
R35620 DVSS.n6551 DVSS.n6380 0.00962857
R35621 DVSS.n6545 DVSS.n6380 0.00962857
R35622 DVSS.n6545 DVSS.n6544 0.00962857
R35623 DVSS.n6544 DVSS.n6543 0.00962857
R35624 DVSS.n6543 DVSS.n6384 0.00962857
R35625 DVSS.n6537 DVSS.n6384 0.00962857
R35626 DVSS.n6537 DVSS.n6536 0.00962857
R35627 DVSS.n6536 DVSS.n6535 0.00962857
R35628 DVSS.n6535 DVSS.n6388 0.00962857
R35629 DVSS.n6529 DVSS.n6388 0.00962857
R35630 DVSS.n6529 DVSS.n6528 0.00962857
R35631 DVSS.n6528 DVSS.n6527 0.00962857
R35632 DVSS.n6527 DVSS.n6392 0.00962857
R35633 DVSS.n6521 DVSS.n6392 0.00962857
R35634 DVSS.n6521 DVSS.n6520 0.00962857
R35635 DVSS.n6520 DVSS.n6519 0.00962857
R35636 DVSS.n6519 DVSS.n6396 0.00962857
R35637 DVSS.n6513 DVSS.n6396 0.00962857
R35638 DVSS.n6513 DVSS.n6512 0.00962857
R35639 DVSS.n6512 DVSS.n6511 0.00962857
R35640 DVSS.n6511 DVSS.n6400 0.00962857
R35641 DVSS.n6505 DVSS.n6400 0.00962857
R35642 DVSS.n6505 DVSS.n6504 0.00962857
R35643 DVSS.n6504 DVSS.n6503 0.00962857
R35644 DVSS.n6503 DVSS.n6404 0.00962857
R35645 DVSS.n6497 DVSS.n6404 0.00962857
R35646 DVSS.n6497 DVSS.n6496 0.00962857
R35647 DVSS.n6496 DVSS.n6495 0.00962857
R35648 DVSS.n6495 DVSS.n6408 0.00962857
R35649 DVSS.n6489 DVSS.n6408 0.00962857
R35650 DVSS.n6489 DVSS.n6488 0.00962857
R35651 DVSS.n6488 DVSS.n6487 0.00962857
R35652 DVSS.n6487 DVSS.n6412 0.00962857
R35653 DVSS.n6481 DVSS.n6412 0.00962857
R35654 DVSS.n6481 DVSS.n6480 0.00962857
R35655 DVSS.n6480 DVSS.n6479 0.00962857
R35656 DVSS.n6479 DVSS.n6416 0.00962857
R35657 DVSS.n6473 DVSS.n6416 0.00962857
R35658 DVSS.n6473 DVSS.n6472 0.00962857
R35659 DVSS.n6472 DVSS.n6471 0.00962857
R35660 DVSS.n6471 DVSS.n6420 0.00962857
R35661 DVSS.n6465 DVSS.n6420 0.00962857
R35662 DVSS.n6465 DVSS.n6464 0.00962857
R35663 DVSS.n6464 DVSS.n6463 0.00962857
R35664 DVSS.n6463 DVSS.n6424 0.00962857
R35665 DVSS.n6457 DVSS.n6424 0.00962857
R35666 DVSS.n6457 DVSS.n6456 0.00962857
R35667 DVSS.n6456 DVSS.n6455 0.00962857
R35668 DVSS.n6455 DVSS.n6428 0.00962857
R35669 DVSS.n6449 DVSS.n6428 0.00962857
R35670 DVSS.n6449 DVSS.n6448 0.00962857
R35671 DVSS.n6448 DVSS.n6447 0.00962857
R35672 DVSS.n6442 DVSS.n6441 0.00962857
R35673 DVSS.n6441 DVSS.n6440 0.00962857
R35674 DVSS.n6440 DVSS.n6433 0.00962857
R35675 DVSS.n6436 DVSS.n6433 0.00962857
R35676 DVSS.n4440 DVSS.n3859 0.00959466
R35677 DVSS.n3865 DVSS.n3863 0.00959466
R35678 DVSS.n3867 DVSS.n3863 0.00959466
R35679 DVSS.n4437 DVSS.n3869 0.00959466
R35680 DVSS.n4196 DVSS.n4194 0.00959466
R35681 DVSS.n4432 DVSS.n4194 0.00959466
R35682 DVSS.n4799 DVSS.n3716 0.00959466
R35683 DVSS.n4800 DVSS.n3715 0.00959466
R35684 DVSS.n3715 DVSS.n3711 0.00959466
R35685 DVSS.n3709 DVSS.n3704 0.00959466
R35686 DVSS.n3709 DVSS.n3707 0.00959466
R35687 DVSS.n4820 DVSS.n3673 0.00959466
R35688 DVSS.n3673 DVSS.n3669 0.00959466
R35689 DVSS.n4826 DVSS.n4824 0.00959466
R35690 DVSS.n4841 DVSS.n3667 0.00959466
R35691 DVSS.n4828 DVSS.n3667 0.00959466
R35692 DVSS.n4839 DVSS.n4831 0.00959466
R35693 DVSS.n4834 DVSS.n4833 0.00959466
R35694 DVSS.n4836 DVSS.n4833 0.00959466
R35695 DVSS.n4975 DVSS.n3590 0.00959466
R35696 DVSS.n3596 DVSS.n3589 0.00959466
R35697 DVSS.n3596 DVSS.n3592 0.00959466
R35698 DVSS.n3866 DVSS.n3865 0.00959466
R35699 DVSS.n4197 DVSS.n4196 0.00959466
R35700 DVSS.n4801 DVSS.n4800 0.00959466
R35701 DVSS.n4804 DVSS.n3704 0.00959466
R35702 DVSS.n4821 DVSS.n4820 0.00959466
R35703 DVSS.n4841 DVSS.n4825 0.00959466
R35704 DVSS.n4835 DVSS.n4834 0.00959466
R35705 DVSS.n4976 DVSS.n3589 0.00959466
R35706 DVSS.n3866 DVSS.n3859 0.00959466
R35707 DVSS.n4438 DVSS.n3867 0.00959466
R35708 DVSS.n4197 DVSS.n3869 0.00959466
R35709 DVSS.n4435 DVSS.n4432 0.00959466
R35710 DVSS.n4801 DVSS.n4799 0.00959466
R35711 DVSS.n4803 DVSS.n3711 0.00959466
R35712 DVSS.n4806 DVSS.n3707 0.00959466
R35713 DVSS.n4823 DVSS.n3669 0.00959466
R35714 DVSS.n4826 DVSS.n4825 0.00959466
R35715 DVSS.n4845 DVSS.n4828 0.00959466
R35716 DVSS.n4835 DVSS.n4831 0.00959466
R35717 DVSS.n4837 DVSS.n4836 0.00959466
R35718 DVSS.n4976 DVSS.n4975 0.00959466
R35719 DVSS.n4978 DVSS.n3592 0.00959466
R35720 DVSS.n3875 DVSS.n3873 0.00959466
R35721 DVSS.n4173 DVSS.n3878 0.00959466
R35722 DVSS.n3884 DVSS.n3870 0.00959466
R35723 DVSS.n3881 DVSS.n3870 0.00959466
R35724 DVSS.n4006 DVSS.n4004 0.00959466
R35725 DVSS.n4007 DVSS.n4003 0.00959466
R35726 DVSS.n4003 DVSS.n4000 0.00959466
R35727 DVSS.n4100 DVSS.n3998 0.00959466
R35728 DVSS.n4095 DVSS.n3998 0.00959466
R35729 DVSS.n3567 DVSS.n3565 0.00959466
R35730 DVSS.n3568 DVSS.n3567 0.00959466
R35731 DVSS.n4998 DVSS.n3570 0.00959466
R35732 DVSS.n3574 DVSS.n3573 0.00959466
R35733 DVSS.n3577 DVSS.n3573 0.00959466
R35734 DVSS.n4994 DVSS.n3580 0.00959466
R35735 DVSS.n3584 DVSS.n3583 0.00959466
R35736 DVSS.n3587 DVSS.n3583 0.00959466
R35737 DVSS.n4991 DVSS.n4981 0.00959466
R35738 DVSS.n4985 DVSS.n4984 0.00959466
R35739 DVSS.n4988 DVSS.n4984 0.00959466
R35740 DVSS.n3877 DVSS.n3873 0.00959466
R35741 DVSS.n3884 DVSS.n3880 0.00959466
R35742 DVSS.n4008 DVSS.n4007 0.00959466
R35743 DVSS.n4100 DVSS.n4099 0.00959466
R35744 DVSS.n5003 DVSS.n3565 0.00959466
R35745 DVSS.n3575 DVSS.n3574 0.00959466
R35746 DVSS.n3585 DVSS.n3584 0.00959466
R35747 DVSS.n4986 DVSS.n4985 0.00959466
R35748 DVSS.n4173 DVSS.n3880 0.00959466
R35749 DVSS.n4189 DVSS.n3881 0.00959466
R35750 DVSS.n4008 DVSS.n4006 0.00959466
R35751 DVSS.n4010 DVSS.n4000 0.00959466
R35752 DVSS.n4095 DVSS.n3562 0.00959466
R35753 DVSS.n5001 DVSS.n3568 0.00959466
R35754 DVSS.n3575 DVSS.n3570 0.00959466
R35755 DVSS.n4996 DVSS.n3577 0.00959466
R35756 DVSS.n3585 DVSS.n3580 0.00959466
R35757 DVSS.n4992 DVSS.n3587 0.00959466
R35758 DVSS.n4986 DVSS.n4981 0.00959466
R35759 DVSS.n4989 DVSS.n4988 0.00959466
R35760 DVSS.n3538 DVSS.n3535 0.00959466
R35761 DVSS.n3543 DVSS.n3541 0.00959466
R35762 DVSS.n3544 DVSS.n3532 0.00959466
R35763 DVSS.n3532 DVSS.n3530 0.00959466
R35764 DVSS.n3551 DVSS.n3549 0.00959466
R35765 DVSS.n3552 DVSS.n3527 0.00959466
R35766 DVSS.n3527 DVSS.n3525 0.00959466
R35767 DVSS.n3557 DVSS.n3523 0.00959466
R35768 DVSS.n3523 DVSS.n3521 0.00959466
R35769 DVSS.n5025 DVSS.n5021 0.00959466
R35770 DVSS.n5025 DVSS.n5023 0.00959466
R35771 DVSS.n5390 DVSS.n3346 0.00959466
R35772 DVSS.n3349 DVSS.n3348 0.00959466
R35773 DVSS.n3349 DVSS.n3345 0.00959466
R35774 DVSS.n5385 DVSS.n3352 0.00959466
R35775 DVSS.n3358 DVSS.n3356 0.00959466
R35776 DVSS.n3360 DVSS.n3356 0.00959466
R35777 DVSS.n5382 DVSS.n3362 0.00959466
R35778 DVSS.n3368 DVSS.n3366 0.00959466
R35779 DVSS.n5369 DVSS.n3366 0.00959466
R35780 DVSS.n3540 DVSS.n3535 0.00959466
R35781 DVSS.n3545 DVSS.n3544 0.00959466
R35782 DVSS.n3553 DVSS.n3552 0.00959466
R35783 DVSS.n3558 DVSS.n3557 0.00959466
R35784 DVSS.n5027 DVSS.n5021 0.00959466
R35785 DVSS.n5389 DVSS.n3348 0.00959466
R35786 DVSS.n3359 DVSS.n3358 0.00959466
R35787 DVSS.n3369 DVSS.n3368 0.00959466
R35788 DVSS.n3545 DVSS.n3543 0.00959466
R35789 DVSS.n3547 DVSS.n3530 0.00959466
R35790 DVSS.n3553 DVSS.n3551 0.00959466
R35791 DVSS.n3555 DVSS.n3525 0.00959466
R35792 DVSS.n3560 DVSS.n3521 0.00959466
R35793 DVSS.n5029 DVSS.n5023 0.00959466
R35794 DVSS.n5390 DVSS.n5389 0.00959466
R35795 DVSS.n5387 DVSS.n3345 0.00959466
R35796 DVSS.n3359 DVSS.n3352 0.00959466
R35797 DVSS.n5383 DVSS.n3360 0.00959466
R35798 DVSS.n3369 DVSS.n3362 0.00959466
R35799 DVSS.n5380 DVSS.n5369 0.00959466
R35800 DVSS.n5674 DVSS.n3255 0.00959466
R35801 DVSS.n5680 DVSS.n5679 0.00959466
R35802 DVSS.n3254 DVSS.n3247 0.00959466
R35803 DVSS.n5687 DVSS.n5686 0.00959466
R35804 DVSS.n3245 DVSS.n3238 0.00959466
R35805 DVSS.n3232 DVSS.n3230 0.00959466
R35806 DVSS.n5489 DVSS.n5402 0.00959466
R35807 DVSS.n5497 DVSS.n5496 0.00959466
R35808 DVSS.n5401 DVSS.n3323 0.00959466
R35809 DVSS.n5504 DVSS.n5503 0.00959466
R35810 DVSS.n3321 DVSS.n3314 0.00959466
R35811 DVSS.n5509 DVSS.n3309 0.00959466
R35812 DVSS.n5512 DVSS.n3310 0.00959466
R35813 DVSS.n5681 DVSS.n5680 0.00959466
R35814 DVSS.n5688 DVSS.n5687 0.00959466
R35815 DVSS.n5498 DVSS.n5497 0.00959466
R35816 DVSS.n5505 DVSS.n5504 0.00959466
R35817 DVSS.n5513 DVSS.n3309 0.00959466
R35818 DVSS.n5677 DVSS.n3255 0.00959466
R35819 DVSS.n5681 DVSS.n3254 0.00959466
R35820 DVSS.n5688 DVSS.n3245 0.00959466
R35821 DVSS.n5691 DVSS.n3230 0.00959466
R35822 DVSS.n5491 DVSS.n5489 0.00959466
R35823 DVSS.n5498 DVSS.n5401 0.00959466
R35824 DVSS.n5505 DVSS.n3321 0.00959466
R35825 DVSS.n5513 DVSS.n5512 0.00959466
R35826 DVSS.n5665 DVSS.n3257 0.00959466
R35827 DVSS.n5664 DVSS.n3261 0.00959466
R35828 DVSS.n3264 DVSS.n3263 0.00959466
R35829 DVSS.n5654 DVSS.n3268 0.00959466
R35830 DVSS.n3271 DVSS.n3270 0.00959466
R35831 DVSS.n3277 DVSS.n3273 0.00959466
R35832 DVSS.n3288 DVSS.n3286 0.00959466
R35833 DVSS.n5547 DVSS.n3291 0.00959466
R35834 DVSS.n3295 DVSS.n3294 0.00959466
R35835 DVSS.n5537 DVSS.n3299 0.00959466
R35836 DVSS.n3303 DVSS.n3302 0.00959466
R35837 DVSS.n5528 DVSS.n3306 0.00959466
R35838 DVSS.n5518 DVSS.n5517 0.00959466
R35839 DVSS.n5659 DVSS.n3261 0.00959466
R35840 DVSS.n5649 DVSS.n3268 0.00959466
R35841 DVSS.n5542 DVSS.n3291 0.00959466
R35842 DVSS.n5532 DVSS.n3299 0.00959466
R35843 DVSS.n5523 DVSS.n3306 0.00959466
R35844 DVSS.n5668 DVSS.n3257 0.00959466
R35845 DVSS.n5659 DVSS.n3263 0.00959466
R35846 DVSS.n5649 DVSS.n3270 0.00959466
R35847 DVSS.n5645 DVSS.n3273 0.00959466
R35848 DVSS.n5633 DVSS.n3286 0.00959466
R35849 DVSS.n5542 DVSS.n3294 0.00959466
R35850 DVSS.n5532 DVSS.n3302 0.00959466
R35851 DVSS.n5523 DVSS.n5517 0.00959466
R35852 DVSS.n2677 DVSS.n2676 0.00959466
R35853 DVSS.n2674 DVSS.n2668 0.00959466
R35854 DVSS.n2683 DVSS.n2682 0.00959466
R35855 DVSS.n2667 DVSS.n2661 0.00959466
R35856 DVSS.n2690 DVSS.n2689 0.00959466
R35857 DVSS.n2659 DVSS.n2653 0.00959466
R35858 DVSS.n2696 DVSS.n2695 0.00959466
R35859 DVSS.n2706 DVSS.n2702 0.00959466
R35860 DVSS.n2749 DVSS.n2710 0.00959466
R35861 DVSS.n2714 DVSS.n2713 0.00959466
R35862 DVSS.n2743 DVSS.n2719 0.00959466
R35863 DVSS.n2723 DVSS.n2722 0.00959466
R35864 DVSS.n2738 DVSS.n2727 0.00959466
R35865 DVSS.n2731 DVSS.n2730 0.00959466
R35866 DVSS.n2678 DVSS.n2677 0.00959466
R35867 DVSS.n2684 DVSS.n2683 0.00959466
R35868 DVSS.n2691 DVSS.n2690 0.00959466
R35869 DVSS.n2712 DVSS.n2710 0.00959466
R35870 DVSS.n2721 DVSS.n2719 0.00959466
R35871 DVSS.n2729 DVSS.n2727 0.00959466
R35872 DVSS.n2678 DVSS.n2674 0.00959466
R35873 DVSS.n2684 DVSS.n2667 0.00959466
R35874 DVSS.n2691 DVSS.n2659 0.00959466
R35875 DVSS.n2695 DVSS.n2694 0.00959466
R35876 DVSS.n2754 DVSS.n2702 0.00959466
R35877 DVSS.n2713 DVSS.n2712 0.00959466
R35878 DVSS.n2722 DVSS.n2721 0.00959466
R35879 DVSS.n2730 DVSS.n2729 0.00959466
R35880 DVSS.n7361 DVSS.n2592 0.00959466
R35881 DVSS.n2596 DVSS.n2595 0.00959466
R35882 DVSS.n7352 DVSS.n2599 0.00959466
R35883 DVSS.n2603 DVSS.n2602 0.00959466
R35884 DVSS.n7342 DVSS.n2607 0.00959466
R35885 DVSS.n2611 DVSS.n2610 0.00959466
R35886 DVSS.n2617 DVSS.n2613 0.00959466
R35887 DVSS.n7325 DVSS.n2080 0.00959466
R35888 DVSS.n7855 DVSS.n2084 0.00959466
R35889 DVSS.n2088 DVSS.n2087 0.00959466
R35890 DVSS.n7725 DVSS.n2092 0.00959466
R35891 DVSS.n2096 DVSS.n2095 0.00959466
R35892 DVSS.n7718 DVSS.n2100 0.00959466
R35893 DVSS.n2104 DVSS.n2103 0.00959466
R35894 DVSS.n7356 DVSS.n2592 0.00959466
R35895 DVSS.n7347 DVSS.n2599 0.00959466
R35896 DVSS.n7337 DVSS.n2607 0.00959466
R35897 DVSS.n7850 DVSS.n2084 0.00959466
R35898 DVSS.n7720 DVSS.n2092 0.00959466
R35899 DVSS.n7713 DVSS.n2100 0.00959466
R35900 DVSS.n7356 DVSS.n2595 0.00959466
R35901 DVSS.n7347 DVSS.n2602 0.00959466
R35902 DVSS.n7337 DVSS.n2610 0.00959466
R35903 DVSS.n7333 DVSS.n2613 0.00959466
R35904 DVSS.n7325 DVSS.n2079 0.00959466
R35905 DVSS.n7850 DVSS.n2087 0.00959466
R35906 DVSS.n7720 DVSS.n2095 0.00959466
R35907 DVSS.n7713 DVSS.n2103 0.00959466
R35908 DVSS.n8073 DVSS.n8072 0.00959466
R35909 DVSS.n1908 DVSS.n1900 0.00959466
R35910 DVSS.n8079 DVSS.n8078 0.00959466
R35911 DVSS.n1899 DVSS.n1891 0.00959466
R35912 DVSS.n8086 DVSS.n8085 0.00959466
R35913 DVSS.n1889 DVSS.n1881 0.00959466
R35914 DVSS.n1876 DVSS.n1874 0.00959466
R35915 DVSS.n8100 DVSS.n1864 0.00959466
R35916 DVSS.n8108 DVSS.n8107 0.00959466
R35917 DVSS.n1863 DVSS.n1855 0.00959466
R35918 DVSS.n8115 DVSS.n8114 0.00959466
R35919 DVSS.n1835 DVSS.n1833 0.00959466
R35920 DVSS.n1851 DVSS.n1839 0.00959466
R35921 DVSS.n1842 DVSS.n1841 0.00959466
R35922 DVSS.n8074 DVSS.n8073 0.00959466
R35923 DVSS.n8080 DVSS.n8079 0.00959466
R35924 DVSS.n8087 DVSS.n8086 0.00959466
R35925 DVSS.n8109 DVSS.n8108 0.00959466
R35926 DVSS.n8116 DVSS.n8115 0.00959466
R35927 DVSS.n1846 DVSS.n1839 0.00959466
R35928 DVSS.n8074 DVSS.n1908 0.00959466
R35929 DVSS.n8080 DVSS.n1899 0.00959466
R35930 DVSS.n8087 DVSS.n1889 0.00959466
R35931 DVSS.n8090 DVSS.n1874 0.00959466
R35932 DVSS.n8102 DVSS.n8100 0.00959466
R35933 DVSS.n8109 DVSS.n1863 0.00959466
R35934 DVSS.n8116 DVSS.n1833 0.00959466
R35935 DVSS.n1846 DVSS.n1841 0.00959466
R35936 DVSS.n5552 DVSS.n2293 0.00958451
R35937 DVSS.n2063 DVSS.n2059 0.00958451
R35938 DVSS.n5623 DVSS.n2323 0.00958451
R35939 DVSS.n2056 DVSS.n2045 0.00958451
R35940 DVSS.n4830 DVSS.n3621 0.00953543
R35941 DVSS.n4838 DVSS.n3616 0.00953543
R35942 DVSS.n4832 DVSS.n3622 0.00953543
R35943 DVSS.n3623 DVSS.n3615 0.00953543
R35944 DVSS.n4887 DVSS.n3626 0.00953543
R35945 DVSS.n9543 DVSS.n9542 0.00953543
R35946 DVSS.n4847 DVSS.n4846 0.00953543
R35947 DVSS.n4844 DVSS.n3651 0.00953543
R35948 DVSS.n4843 DVSS.n3650 0.00953543
R35949 DVSS.n4827 DVSS.n3649 0.00953543
R35950 DVSS.n4842 DVSS.n3648 0.00953543
R35951 DVSS.n9377 DVSS.n9368 0.00953543
R35952 DVSS.n4795 DVSS.n3710 0.00953543
R35953 DVSS.n4802 DVSS.n3714 0.00953543
R35954 DVSS.n3717 DVSS.n3713 0.00953543
R35955 DVSS.n4798 DVSS.n3718 0.00953543
R35956 DVSS.n4797 DVSS.n3712 0.00953543
R35957 DVSS.n9015 DVSS.n705 0.00953543
R35958 DVSS.n4428 DVSS.n3868 0.00953543
R35959 DVSS.n4436 DVSS.n4193 0.00953543
R35960 DVSS.n4195 DVSS.n4192 0.00953543
R35961 DVSS.n4431 DVSS.n4198 0.00953543
R35962 DVSS.n4430 DVSS.n4191 0.00953543
R35963 DVSS.n9009 DVSS.n712 0.00953543
R35964 DVSS.n8936 DVSS.n8934 0.00953543
R35965 DVSS.n8968 DVSS.n732 0.00953543
R35966 DVSS.n4257 DVSS.n3858 0.00953543
R35967 DVSS.n4439 DVSS.n3862 0.00953543
R35968 DVSS.n3864 DVSS.n3861 0.00953543
R35969 DVSS.n4221 DVSS.n4216 0.00953543
R35970 DVSS.n4259 DVSS.n3860 0.00953543
R35971 DVSS.n4971 DVSS.n3591 0.00953543
R35972 DVSS.n4977 DVSS.n3595 0.00953543
R35973 DVSS.n3597 DVSS.n3594 0.00953543
R35974 DVSS.n4974 DVSS.n4973 0.00953543
R35975 DVSS.n4979 DVSS.n3588 0.00953543
R35976 DVSS.n9470 DVSS.n9468 0.00953543
R35977 DVSS.n9502 DVSS.n31 0.00953543
R35978 DVSS.n4931 DVSS.n4917 0.00953543
R35979 DVSS.n5917 DVSS.n5916 0.00953543
R35980 DVSS.n4445 DVSS.n3852 0.00953543
R35981 DVSS.n5865 DVSS.n3017 0.00953543
R35982 DVSS.n4746 DVSS.n4744 0.00951408
R35983 DVSS.n6647 DVSS.n6644 0.00943102
R35984 DVSS.n9422 DVSS.n9420 0.00934615
R35985 DVSS.n9533 DVSS.n9532 0.00934615
R35986 DVSS.n9000 DVSS.n714 0.00934615
R35987 DVSS.n9533 DVSS.n332 0.00934615
R35988 DVSS.n8888 DVSS.n8886 0.00934615
R35989 DVSS.n9000 DVSS.n8999 0.00934615
R35990 DVSS.n8886 DVSS.n8885 0.00934615
R35991 DVSS.n9420 DVSS.n365 0.00934615
R35992 DVSS.n9716 DVSS.n181 0.0091811
R35993 DVSS.n9659 DVSS.n220 0.0091811
R35994 DVSS.n8873 DVSS.n801 0.0091811
R35995 DVSS.n8878 DVSS.n791 0.0091811
R35996 DVSS.n8905 DVSS.n765 0.0091811
R35997 DVSS.n9439 DVSS.n350 0.0091811
R35998 DVSS.n5018 DVSS.n3517 0.00916197
R35999 DVSS.n5570 DVSS.n2284 0.00916197
R36000 DVSS.n5202 DVSS.n3183 0.00916197
R36001 DVSS.n5586 DVSS.n2314 0.00916197
R36002 DVSS.n6643 DVSS.n2756 0.00910927
R36003 DVSS.n7262 DVSS.n2756 0.00910927
R36004 DVSS.n7261 DVSS.n7260 0.00910927
R36005 DVSS.n7262 DVSS.n7261 0.00910927
R36006 DVSS.n7243 DVSS.n6644 0.00909923
R36007 DVSS.n8404 DVSS.n8403 0.00898571
R36008 DVSS.n7943 DVSS.n2039 0.00898571
R36009 DVSS.n5748 DVSS.n3170 0.00898571
R36010 DVSS.n3969 DVSS.n3965 0.00898571
R36011 DVSS.n4809 DVSS.n3691 0.00898571
R36012 DVSS.n8917 DVSS.n762 0.00882677
R36013 DVSS.n8952 DVSS.n740 0.00882677
R36014 DVSS.n9451 DVSS.n347 0.00882677
R36015 DVSS.n9486 DVSS.n38 0.00882677
R36016 DVSS.n6010 DVSS.n2764 0.00873944
R36017 DVSS.n3986 DVSS.n3484 0.00873944
R36018 DVSS.n5575 DVSS.n2303 0.00873944
R36019 DVSS.n4756 DVSS.n3780 0.00873944
R36020 DVSS.n4104 DVSS.n3981 0.00873944
R36021 DVSS.n5576 DVSS.n2333 0.00873944
R36022 DVSS.n8388 DVSS.n1414 0.00872857
R36023 DVSS.n7764 DVSS.n2061 0.00872857
R36024 DVSS.n5038 DVSS.n5010 0.00872857
R36025 DVSS.n5244 DVSS.n3470 0.00872857
R36026 DVSS.n4308 DVSS.n3678 0.00872857
R36027 DVSS.n5946 DVSS 0.00852817
R36028 DVSS.n3783 DVSS.n3775 0.00852817
R36029 DVSS DVSS.n2871 0.00852817
R36030 DVSS.n4446 DVSS.n3857 0.00848752
R36031 DVSS.n4443 DVSS.n3857 0.00848752
R36032 DVSS.n4930 DVSS.n4928 0.00848752
R36033 DVSS.n4927 DVSS.n2911 0.00848752
R36034 DVSS.n4928 DVSS.n4927 0.00848752
R36035 DVSS.n4933 DVSS.n4930 0.00848752
R36036 DVSS.n3022 DVSS.n3019 0.00848752
R36037 DVSS.n3024 DVSS.n3022 0.00848752
R36038 DVSS.n2921 DVSS.n2918 0.00848752
R36039 DVSS.n5920 DVSS.n2913 0.00848752
R36040 DVSS.n2918 DVSS.n2913 0.00848752
R36041 DVSS.n5918 DVSS.n2921 0.00848752
R36042 DVSS.n5874 DVSS.n3014 0.00848752
R36043 DVSS.n5872 DVSS.n3014 0.00848752
R36044 DVSS.n5373 DVSS.n5370 0.00848752
R36045 DVSS.n5376 DVSS.n5374 0.00848752
R36046 DVSS.n5374 DVSS.n5373 0.00848752
R36047 DVSS.n5378 DVSS.n5370 0.00848752
R36048 DVSS.n5883 DVSS.n5882 0.00848752
R36049 DVSS.n2963 DVSS.n2960 0.00848752
R36050 DVSS.n5907 DVSS.n2967 0.00848752
R36051 DVSS.n2967 DVSS.n2960 0.00848752
R36052 DVSS.n5909 DVSS.n2963 0.00848752
R36053 DVSS.n5892 DVSS.n2982 0.00848752
R36054 DVSS.n2972 DVSS.n2969 0.00848752
R36055 DVSS.n5902 DVSS.n2976 0.00848752
R36056 DVSS.n2976 DVSS.n2969 0.00848752
R36057 DVSS.n5904 DVSS.n2972 0.00848752
R36058 DVSS.n2585 DVSS.n2578 0.00848752
R36059 DVSS.n2117 DVSS.n2109 0.00848752
R36060 DVSS.n7698 DVSS.n2111 0.00848752
R36061 DVSS.n2111 DVSS.n2109 0.00848752
R36062 DVSS.n7696 DVSS.n2117 0.00848752
R36063 DVSS.n7365 DVSS.n2587 0.00848752
R36064 DVSS.n7700 DVSS.n2106 0.00848752
R36065 DVSS.n7705 DVSS.n7703 0.00848752
R36066 DVSS.n7703 DVSS.n7700 0.00848752
R36067 DVSS.n7708 DVSS.n2106 0.00848752
R36068 DVSS.n8065 DVSS.n1912 0.00848752
R36069 DVSS.n1760 DVSS.n1756 0.00848752
R36070 DVSS.n8184 DVSS.n1753 0.00848752
R36071 DVSS.n1756 DVSS.n1753 0.00848752
R36072 DVSS.n8181 DVSS.n1760 0.00848752
R36073 DVSS.n8069 DVSS.n1912 0.00848752
R36074 DVSS.n7368 DVSS.n2587 0.00848752
R36075 DVSS.n7373 DVSS.n2578 0.00848752
R36076 DVSS.n5893 DVSS.n5892 0.00848752
R36077 DVSS.n5882 DVSS.n2991 0.00848752
R36078 DVSS.n5876 DVSS.n5874 0.00848752
R36079 DVSS.n5872 DVSS.n3015 0.00848752
R36080 DVSS.n5869 DVSS.n3019 0.00848752
R36081 DVSS.n5867 DVSS.n3024 0.00848752
R36082 DVSS.n4448 DVSS.n4446 0.00848752
R36083 DVSS.n4443 DVSS.n4442 0.00848752
R36084 DVSS.n8921 DVSS.n778 0.00847244
R36085 DVSS.n8956 DVSS.n735 0.00847244
R36086 DVSS.n9455 DVSS.n362 0.00847244
R36087 DVSS.n9490 DVSS.n34 0.00847244
R36088 DVSS.n3983 DVSS.n3483 0.0083169
R36089 DVSS.n3992 DVSS.n3979 0.0083169
R36090 DVSS.n4501 DVSS.n3825 0.0083169
R36091 DVSS.n4588 DVSS.n3802 0.0083169
R36092 DVSS.n4784 DVSS.n3730 0.0083169
R36093 DVSS.n4749 DVSS.n4622 0.00824648
R36094 DVSS.n8901 DVSS.n774 0.00811811
R36095 DVSS.n8998 DVSS.n719 0.00811811
R36096 DVSS.n9435 DVSS.n358 0.00811811
R36097 DVSS.n9887 DVSS.n48 0.00811811
R36098 DVSS.n4626 DVSS.n4618 0.00810563
R36099 DVSS.n4697 DVSS.n3772 0.00810563
R36100 DVSS.n5994 DVSS.n2781 0.00803521
R36101 DVSS.n5967 DVSS.n2830 0.00803521
R36102 DVSS.n5950 DVSS.n2863 0.00803521
R36103 DVSS.n5567 DVSS.n2285 0.00789437
R36104 DVSS.n5592 DVSS.n2315 0.00789437
R36105 DVSS DVSS.n4904 0.00782857
R36106 DVSS DVSS.n1738 0.00782857
R36107 DVSS.n1377 DVSS.n1367 0.00782857
R36108 DVSS.n1737 DVSS 0.00782857
R36109 DVSS.n8162 DVSS 0.00782857
R36110 DVSS.n2044 DVSS.n2043 0.00782857
R36111 DVSS.n8161 DVSS 0.00782857
R36112 DVSS.n5103 DVSS 0.00782857
R36113 DVSS.n3175 DVSS.n3174 0.00782857
R36114 DVSS.n5105 DVSS 0.00782857
R36115 DVSS.n5339 DVSS 0.00782857
R36116 DVSS.n4106 DVSS.n4105 0.00782857
R36117 DVSS.n5340 DVSS 0.00782857
R36118 DVSS.n3703 DVSS.n3697 0.00782857
R36119 DVSS DVSS.n4903 0.00782857
R36120 DVSS.n6446 VSS 0.00782857
R36121 VSS DVSS.n6152 0.00782857
R36122 DVSS.n6168 VSS 0.00782857
R36123 DVSS.n6447 VSS 0.00782857
R36124 DVSS.n8939 DVSS.n754 0.00776378
R36125 DVSS.n8972 DVSS.n744 0.00776378
R36126 DVSS.n9473 DVSS.n339 0.00776378
R36127 DVSS.n9506 DVSS.n42 0.00776378
R36128 DVSS.n4932 DVSS.n4908 0.00776378
R36129 DVSS.n2930 DVSS.n2914 0.00776378
R36130 DVSS.n4447 DVSS.n3841 0.00776378
R36131 DVSS.n3026 DVSS.n3018 0.00776378
R36132 DVSS.n7062 DVSS.n6669 0.00763571
R36133 DVSS.n8452 DVSS.n1164 0.00763571
R36134 DVSS.n8439 DVSS.n1328 0.00763571
R36135 DVSS.n8044 DVSS.n1945 0.00763571
R36136 DVSS.n8021 DVSS.n1971 0.00763571
R36137 DVSS.n7982 DVSS.n2005 0.00763571
R36138 DVSS.n5814 DVSS.n5813 0.00763571
R36139 DVSS.n5784 DVSS.n3136 0.00763571
R36140 DVSS.n4186 DVSS.n3890 0.00763571
R36141 DVSS.n4140 DVSS.n4139 0.00763571
R36142 DVSS.n4258 DVSS.n4224 0.00763571
R36143 DVSS.n4429 DVSS.n4202 0.00763571
R36144 DVSS.n4796 DVSS.n3722 0.00763571
R36145 DVSS.n8392 DVSS.n1404 0.00757143
R36146 DVSS.n7770 DVSS.n2060 0.00757143
R36147 DVSS.n5194 DVSS.n5193 0.00757143
R36148 DVSS.n5237 DVSS.n3480 0.00757143
R36149 DVSS.n4346 DVSS.n3677 0.00757143
R36150 DVSS.n5555 DVSS.n2294 0.00747183
R36151 DVSS.n7891 DVSS.n2064 0.00747183
R36152 DVSS.n5617 DVSS.n2324 0.00747183
R36153 DVSS.n7892 DVSS.n2046 0.00747183
R36154 DVSS.n5974 DVSS.n2827 0.00740945
R36155 DVSS.n6007 DVSS.n2773 0.00740945
R36156 DVSS.n4783 DVSS.n3743 0.00740945
R36157 DVSS.n4594 DVSS.n3796 0.00740945
R36158 DVSS.n786 DVSS.n769 0.00740945
R36159 DVSS.n8982 DVSS.n729 0.00740945
R36160 DVSS.n4518 DVSS.n3824 0.00740945
R36161 DVSS.n5959 DVSS.n2858 0.00740945
R36162 DVSS.n366 DVSS.n354 0.00740945
R36163 DVSS.n9516 DVSS.n28 0.00740945
R36164 DVSS.n5942 DVSS.n2887 0.00740945
R36165 DVSS.n2956 DVSS.n2944 0.00740945
R36166 DVSS.n4491 DVSS.n4460 0.00740945
R36167 DVSS.n2998 DVSS.n2993 0.00740945
R36168 DVSS.n1623 DVSS.n1426 0.00737857
R36169 DVSS.n1609 DVSS.n1106 0.00737857
R36170 DVSS.n1727 DVSS.n1590 0.00737857
R36171 DVSS.n7837 DVSS.n7729 0.00737857
R36172 DVSS.n8123 DVSS.n1804 0.00737857
R36173 DVSS.n8152 DVSS.n1784 0.00737857
R36174 DVSS.n5393 DVSS.n3332 0.00737857
R36175 DVSS.n5128 DVSS.n5127 0.00737857
R36176 DVSS.n5366 DVSS.n3376 0.00737857
R36177 DVSS.n5279 DVSS.n3436 0.00737857
R36178 DVSS.n5314 DVSS.n3401 0.00737857
R36179 DVSS.n5349 DVSS.n5347 0.00737857
R36180 DVSS.n4850 DVSS.n3643 0.00737857
R36181 DVSS.n4888 DVSS.n3610 0.00737857
R36182 DVSS.n4953 DVSS.n3599 0.00737857
R36183 DVSS.n4755 DVSS.n4607 0.00726056
R36184 DVSS.n6344 DVSS.n6034 0.00725
R36185 DVSS.n6623 DVSS.n6028 0.00725
R36186 DVSS.n4495 DVSS.n3832 0.00716667
R36187 DVSS.n4496 DVSS.n4495 0.00716667
R36188 DVSS.n4497 DVSS.n4496 0.00716667
R36189 DVSS.n4497 DVSS.n3828 0.00716667
R36190 DVSS.n4504 DVSS.n3828 0.00716667
R36191 DVSS.n4505 DVSS.n4504 0.00716667
R36192 DVSS.n4506 DVSS.n4505 0.00716667
R36193 DVSS.n4506 DVSS.n3813 0.00716667
R36194 DVSS.n4522 DVSS.n3813 0.00716667
R36195 DVSS.n4523 DVSS.n4522 0.00716667
R36196 DVSS.n4524 DVSS.n4523 0.00716667
R36197 DVSS.n4524 DVSS.n3809 0.00716667
R36198 DVSS.n4530 DVSS.n3809 0.00716667
R36199 DVSS.n4531 DVSS.n4530 0.00716667
R36200 DVSS.n4532 DVSS.n4531 0.00716667
R36201 DVSS.n4533 DVSS.n4532 0.00716667
R36202 DVSS.n4534 DVSS.n4533 0.00716667
R36203 DVSS.n4535 DVSS.n4534 0.00716667
R36204 DVSS.n4538 DVSS.n4535 0.00716667
R36205 DVSS.n4539 DVSS.n4538 0.00716667
R36206 DVSS.n4540 DVSS.n4539 0.00716667
R36207 DVSS.n4541 DVSS.n4540 0.00716667
R36208 DVSS.n4544 DVSS.n4541 0.00716667
R36209 DVSS.n4545 DVSS.n4544 0.00716667
R36210 DVSS.n4546 DVSS.n4545 0.00716667
R36211 DVSS.n4547 DVSS.n4546 0.00716667
R36212 DVSS.n4550 DVSS.n4547 0.00716667
R36213 DVSS.n4551 DVSS.n4550 0.00716667
R36214 DVSS.n4552 DVSS.n4551 0.00716667
R36215 DVSS.n4554 DVSS.n4552 0.00716667
R36216 DVSS.n4554 DVSS.n4553 0.00716667
R36217 DVSS.n4553 DVSS.n3748 0.00716667
R36218 DVSS.n3749 DVSS.n3748 0.00716667
R36219 DVSS.n3750 DVSS.n3749 0.00716667
R36220 DVSS.n3753 DVSS.n3750 0.00716667
R36221 DVSS.n3754 DVSS.n3753 0.00716667
R36222 DVSS.n3755 DVSS.n3754 0.00716667
R36223 DVSS.n3756 DVSS.n3755 0.00716667
R36224 DVSS.n3759 DVSS.n3756 0.00716667
R36225 DVSS.n3760 DVSS.n3759 0.00716667
R36226 DVSS.n3761 DVSS.n3760 0.00716667
R36227 DVSS.n3762 DVSS.n3761 0.00716667
R36228 DVSS.n3765 DVSS.n3762 0.00716667
R36229 DVSS.n3766 DVSS.n3765 0.00716667
R36230 DVSS.n3767 DVSS.n3766 0.00716667
R36231 DVSS.n3768 DVSS.n3767 0.00716667
R36232 DVSS.n4610 DVSS.n3768 0.00716667
R36233 DVSS.n4611 DVSS.n4610 0.00716667
R36234 DVSS.n4612 DVSS.n4611 0.00716667
R36235 DVSS.n4613 DVSS.n4612 0.00716667
R36236 DVSS.n4614 DVSS.n4613 0.00716667
R36237 DVSS.n4706 DVSS.n4614 0.00716667
R36238 DVSS.n4707 DVSS.n4706 0.00716667
R36239 DVSS.n4708 DVSS.n4707 0.00716667
R36240 DVSS.n4709 DVSS.n4708 0.00716667
R36241 DVSS.n4712 DVSS.n4709 0.00716667
R36242 DVSS.n4713 DVSS.n4712 0.00716667
R36243 DVSS.n4714 DVSS.n4713 0.00716667
R36244 DVSS.n4715 DVSS.n4714 0.00716667
R36245 DVSS.n4718 DVSS.n4715 0.00716667
R36246 DVSS.n4719 DVSS.n4718 0.00716667
R36247 DVSS.n4720 DVSS.n4719 0.00716667
R36248 DVSS.n4721 DVSS.n4720 0.00716667
R36249 DVSS.n4722 DVSS.n4721 0.00716667
R36250 DVSS.n4724 DVSS.n4722 0.00716667
R36251 DVSS.n4724 DVSS.n4723 0.00716667
R36252 DVSS.n4723 DVSS.n2795 0.00716667
R36253 DVSS.n2796 DVSS.n2795 0.00716667
R36254 DVSS.n2797 DVSS.n2796 0.00716667
R36255 DVSS.n2800 DVSS.n2797 0.00716667
R36256 DVSS.n2801 DVSS.n2800 0.00716667
R36257 DVSS.n2802 DVSS.n2801 0.00716667
R36258 DVSS.n2803 DVSS.n2802 0.00716667
R36259 DVSS.n2806 DVSS.n2803 0.00716667
R36260 DVSS.n2807 DVSS.n2806 0.00716667
R36261 DVSS.n2808 DVSS.n2807 0.00716667
R36262 DVSS.n2809 DVSS.n2808 0.00716667
R36263 DVSS.n2812 DVSS.n2809 0.00716667
R36264 DVSS.n2813 DVSS.n2812 0.00716667
R36265 DVSS.n2814 DVSS.n2813 0.00716667
R36266 DVSS.n2815 DVSS.n2814 0.00716667
R36267 DVSS.n2837 DVSS.n2815 0.00716667
R36268 DVSS.n2838 DVSS.n2837 0.00716667
R36269 DVSS.n2839 DVSS.n2838 0.00716667
R36270 DVSS.n2840 DVSS.n2839 0.00716667
R36271 DVSS.n2843 DVSS.n2840 0.00716667
R36272 DVSS.n2844 DVSS.n2843 0.00716667
R36273 DVSS.n2845 DVSS.n2844 0.00716667
R36274 DVSS.n2846 DVSS.n2845 0.00716667
R36275 DVSS.n2866 DVSS.n2846 0.00716667
R36276 DVSS.n2867 DVSS.n2866 0.00716667
R36277 DVSS.n2868 DVSS.n2867 0.00716667
R36278 DVSS.n2869 DVSS.n2868 0.00716667
R36279 DVSS.n2872 DVSS.n2869 0.00716667
R36280 DVSS.n2873 DVSS.n2872 0.00716667
R36281 DVSS.n2874 DVSS.n2873 0.00716667
R36282 DVSS.n2875 DVSS.n2874 0.00716667
R36283 DVSS.n5935 DVSS.n5934 0.00716667
R36284 DVSS.n4448 DVSS.n3016 0.00716667
R36285 DVSS.n5922 DVSS.n2911 0.00716667
R36286 DVSS.n5870 DVSS.n5869 0.00716667
R36287 DVSS.n5921 DVSS.n5920 0.00716667
R36288 DVSS.n5876 DVSS.n5871 0.00716667
R36289 DVSS.n5376 DVSS.n2912 0.00716667
R36290 DVSS.n5889 DVSS.n2978 0.00716667
R36291 DVSS.n5907 DVSS.n2968 0.00716667
R36292 DVSS.n5896 DVSS.n5895 0.00716667
R36293 DVSS.n5902 DVSS.n5900 0.00716667
R36294 DVSS.n2980 DVSS.n2579 0.00716667
R36295 DVSS.n7698 DVSS.n2112 0.00716667
R36296 DVSS.n2979 DVSS.n2588 0.00716667
R36297 DVSS.n7705 DVSS.n1752 0.00716667
R36298 DVSS.n8067 DVSS.n1915 0.00716667
R36299 DVSS.n8185 DVSS.n8184 0.00716667
R36300 DVSS.n8891 DVSS.n768 0.00705512
R36301 DVSS.n8988 DVSS.n728 0.00705512
R36302 DVSS.n9425 DVSS.n353 0.00705512
R36303 DVSS.n9522 DVSS.n27 0.00705512
R36304 DVSS.n5375 DVSS.n2945 0.00705512
R36305 DVSS.n5873 DVSS.n2999 0.00705512
R36306 DVSS.n4814 DVSS.n4813 0.0070493
R36307 DVSS.n5559 DVSS.n2296 0.0070493
R36308 DVSS.n7879 DVSS.n2066 0.0070493
R36309 DVSS.n4811 DVSS.n3688 0.0070493
R36310 DVSS.n5609 DVSS.n2326 0.0070493
R36311 DVSS.n7880 DVSS.n2048 0.0070493
R36312 DVSS.n4490 DVSS.n4481 0.0070493
R36313 DVSS.n4517 DVSS.n4508 0.0070493
R36314 DVSS.n4579 DVSS.n3799 0.0070493
R36315 DVSS.n4782 DVSS.n3735 0.0070493
R36316 DVSS.n5934 DVSS 0.00697887
R36317 DVSS.n4750 DVSS.n4616 0.00697887
R36318 DVSS.n7257 DVSS.n7256 0.00678019
R36319 DVSS.n7259 DVSS.n380 0.00678019
R36320 DVSS.n6003 DVSS.n2783 0.00676761
R36321 DVSS.n5996 DVSS.n2782 0.00676761
R36322 DVSS.n5976 DVSS.n5975 0.00676761
R36323 DVSS.n5969 DVSS.n2833 0.00676761
R36324 DVSS.n5961 DVSS.n5960 0.00676761
R36325 DVSS.n5952 DVSS.n2865 0.00676761
R36326 DVSS.n5944 DVSS.n5943 0.00676761
R36327 DVSS.n5937 DVSS.n5930 0.00676761
R36328 DVSS.n8931 DVSS.n759 0.00670079
R36329 DVSS.n8966 DVSS.n743 0.00670079
R36330 DVSS.n9465 DVSS.n344 0.00670079
R36331 DVSS.n9500 DVSS.n41 0.00670079
R36332 DVSS.n4918 DVSS.n4907 0.00670079
R36333 DVSS.n5919 DVSS.n2917 0.00670079
R36334 DVSS.n3853 DVSS.n3840 0.00670079
R36335 DVSS.n5868 DVSS.n3021 0.00670079
R36336 DVSS.n8400 DVSS.n1388 0.00667143
R36337 DVSS.n7937 DVSS.n7936 0.00667143
R36338 DVSS.n5742 DVSS.n5741 0.00667143
R36339 DVSS.n4103 DVSS.n3976 0.00667143
R36340 DVSS.n4353 DVSS.n3690 0.00667143
R36341 DVSS.n4657 DVSS.n3682 0.00662676
R36342 DVSS.n5563 DVSS.n2287 0.00662676
R36343 DVSS.n2075 DVSS.n2069 0.00662676
R36344 DVSS.n4664 DVSS.n3696 0.00662676
R36345 DVSS.n5600 DVSS.n2317 0.00662676
R36346 DVSS.n7868 DVSS.n2051 0.00662676
R36347 DVSS.n4240 DVSS.n4234 0.00658571
R36348 DVSS.n4241 DVSS.n4240 0.00658571
R36349 DVSS.n4242 DVSS.n4241 0.00658571
R36350 DVSS.n4242 DVSS.n4230 0.00658571
R36351 DVSS.n4248 DVSS.n4230 0.00658571
R36352 DVSS.n4249 DVSS.n4248 0.00658571
R36353 DVSS.n4250 DVSS.n4249 0.00658571
R36354 DVSS.n4250 DVSS.n4213 0.00658571
R36355 DVSS.n4263 DVSS.n4213 0.00658571
R36356 DVSS.n4264 DVSS.n4263 0.00658571
R36357 DVSS.n4265 DVSS.n4264 0.00658571
R36358 DVSS.n4265 DVSS.n4209 0.00658571
R36359 DVSS.n4271 DVSS.n4209 0.00658571
R36360 DVSS.n4272 DVSS.n4271 0.00658571
R36361 DVSS.n4416 DVSS.n4272 0.00658571
R36362 DVSS.n4416 DVSS.n4415 0.00658571
R36363 DVSS.n4415 DVSS.n4414 0.00658571
R36364 DVSS.n4414 DVSS.n4273 0.00658571
R36365 DVSS.n4277 DVSS.n4273 0.00658571
R36366 DVSS.n4406 DVSS.n4277 0.00658571
R36367 DVSS.n4406 DVSS.n4405 0.00658571
R36368 DVSS.n4405 DVSS.n4404 0.00658571
R36369 DVSS.n4404 DVSS.n4278 0.00658571
R36370 DVSS.n4398 DVSS.n4278 0.00658571
R36371 DVSS.n4398 DVSS.n4397 0.00658571
R36372 DVSS.n4397 DVSS.n4396 0.00658571
R36373 DVSS.n4396 DVSS.n4282 0.00658571
R36374 DVSS.n4390 DVSS.n4282 0.00658571
R36375 DVSS.n4390 DVSS.n4389 0.00658571
R36376 DVSS.n4389 DVSS.n4388 0.00658571
R36377 DVSS.n4388 DVSS.n4286 0.00658571
R36378 DVSS.n4383 DVSS.n4286 0.00658571
R36379 DVSS.n4383 DVSS.n4382 0.00658571
R36380 DVSS.n4382 DVSS.n4381 0.00658571
R36381 DVSS.n4381 DVSS.n4289 0.00658571
R36382 DVSS.n4375 DVSS.n4289 0.00658571
R36383 DVSS.n4375 DVSS.n4374 0.00658571
R36384 DVSS.n4374 DVSS.n4373 0.00658571
R36385 DVSS.n4373 DVSS.n4293 0.00658571
R36386 DVSS.n4367 DVSS.n4293 0.00658571
R36387 DVSS.n4367 DVSS.n4366 0.00658571
R36388 DVSS.n4366 DVSS.n4365 0.00658571
R36389 DVSS.n4365 DVSS.n4297 0.00658571
R36390 DVSS.n4359 DVSS.n4297 0.00658571
R36391 DVSS.n4359 DVSS.n4358 0.00658571
R36392 DVSS.n4358 DVSS.n4357 0.00658571
R36393 DVSS.n4357 DVSS.n4301 0.00658571
R36394 DVSS.n4352 DVSS.n4301 0.00658571
R36395 DVSS.n4352 DVSS.n4351 0.00658571
R36396 DVSS.n4351 DVSS.n4350 0.00658571
R36397 DVSS.n4350 DVSS.n4304 0.00658571
R36398 DVSS.n4345 DVSS.n4304 0.00658571
R36399 DVSS.n4345 DVSS.n4344 0.00658571
R36400 DVSS.n4344 DVSS.n4343 0.00658571
R36401 DVSS.n4343 DVSS.n4306 0.00658571
R36402 DVSS.n4337 DVSS.n4306 0.00658571
R36403 DVSS.n4337 DVSS.n4336 0.00658571
R36404 DVSS.n4336 DVSS.n4335 0.00658571
R36405 DVSS.n4335 DVSS.n4311 0.00658571
R36406 DVSS.n4329 DVSS.n4311 0.00658571
R36407 DVSS.n4329 DVSS.n4328 0.00658571
R36408 DVSS.n4328 DVSS.n4327 0.00658571
R36409 DVSS.n4327 DVSS.n4315 0.00658571
R36410 DVSS.n4321 DVSS.n4315 0.00658571
R36411 DVSS.n4321 DVSS.n4320 0.00658571
R36412 DVSS.n4320 DVSS.n4319 0.00658571
R36413 DVSS.n4319 DVSS.n3645 0.00658571
R36414 DVSS.n4853 DVSS.n3645 0.00658571
R36415 DVSS.n4854 DVSS.n4853 0.00658571
R36416 DVSS.n4855 DVSS.n4854 0.00658571
R36417 DVSS.n4855 DVSS.n3641 0.00658571
R36418 DVSS.n4861 DVSS.n3641 0.00658571
R36419 DVSS.n4862 DVSS.n4861 0.00658571
R36420 DVSS.n4863 DVSS.n4862 0.00658571
R36421 DVSS.n4863 DVSS.n3637 0.00658571
R36422 DVSS.n4869 DVSS.n3637 0.00658571
R36423 DVSS.n4870 DVSS.n4869 0.00658571
R36424 DVSS.n4871 DVSS.n4870 0.00658571
R36425 DVSS.n4871 DVSS.n3633 0.00658571
R36426 DVSS.n4877 DVSS.n3633 0.00658571
R36427 DVSS.n4878 DVSS.n4877 0.00658571
R36428 DVSS.n4879 DVSS.n4878 0.00658571
R36429 DVSS.n4879 DVSS.n3612 0.00658571
R36430 DVSS.n4891 DVSS.n3612 0.00658571
R36431 DVSS.n4892 DVSS.n4891 0.00658571
R36432 DVSS.n4893 DVSS.n4892 0.00658571
R36433 DVSS.n4893 DVSS.n3608 0.00658571
R36434 DVSS.n4899 DVSS.n3608 0.00658571
R36435 DVSS.n4900 DVSS.n4899 0.00658571
R36436 DVSS.n4959 DVSS.n4900 0.00658571
R36437 DVSS.n4959 DVSS.n4958 0.00658571
R36438 DVSS.n4958 DVSS.n4957 0.00658571
R36439 DVSS.n4957 DVSS.n4901 0.00658571
R36440 DVSS.n4905 DVSS.n4901 0.00658571
R36441 DVSS.n4949 DVSS.n4905 0.00658571
R36442 DVSS.n4949 DVSS.n4948 0.00658571
R36443 DVSS.n4948 DVSS.n4947 0.00658571
R36444 DVSS.n4938 DVSS.n4937 0.00658571
R36445 DVSS.n6770 DVSS.n6769 0.00658571
R36446 DVSS.n6848 DVSS.n6770 0.00658571
R36447 DVSS.n6848 DVSS.n6847 0.00658571
R36448 DVSS.n6847 DVSS.n6846 0.00658571
R36449 DVSS.n6846 DVSS.n6771 0.00658571
R36450 DVSS.n6840 DVSS.n6771 0.00658571
R36451 DVSS.n6840 DVSS.n6839 0.00658571
R36452 DVSS.n6839 DVSS.n6838 0.00658571
R36453 DVSS.n6838 DVSS.n6773 0.00658571
R36454 DVSS.n6775 DVSS.n6773 0.00658571
R36455 DVSS.n6778 DVSS.n6775 0.00658571
R36456 DVSS.n6828 DVSS.n6778 0.00658571
R36457 DVSS.n6828 DVSS.n6827 0.00658571
R36458 DVSS.n6827 DVSS.n6826 0.00658571
R36459 DVSS.n6826 DVSS.n6779 0.00658571
R36460 DVSS.n6821 DVSS.n6779 0.00658571
R36461 DVSS.n6821 DVSS.n6820 0.00658571
R36462 DVSS.n6820 DVSS.n6819 0.00658571
R36463 DVSS.n6819 DVSS.n6782 0.00658571
R36464 DVSS.n6813 DVSS.n6782 0.00658571
R36465 DVSS.n6813 DVSS.n6812 0.00658571
R36466 DVSS.n6812 DVSS.n6811 0.00658571
R36467 DVSS.n6811 DVSS.n6786 0.00658571
R36468 DVSS.n6805 DVSS.n6786 0.00658571
R36469 DVSS.n6805 DVSS.n6804 0.00658571
R36470 DVSS.n6804 DVSS.n6803 0.00658571
R36471 DVSS.n6803 DVSS.n6790 0.00658571
R36472 DVSS.n6797 DVSS.n6790 0.00658571
R36473 DVSS.n6797 DVSS.n6796 0.00658571
R36474 DVSS.n6796 DVSS.n6795 0.00658571
R36475 DVSS.n6795 DVSS.n1347 0.00658571
R36476 DVSS.n8432 DVSS.n1347 0.00658571
R36477 DVSS.n8432 DVSS.n8431 0.00658571
R36478 DVSS.n8431 DVSS.n8430 0.00658571
R36479 DVSS.n8430 DVSS.n1348 0.00658571
R36480 DVSS.n8424 DVSS.n1348 0.00658571
R36481 DVSS.n8424 DVSS.n8423 0.00658571
R36482 DVSS.n8423 DVSS.n8422 0.00658571
R36483 DVSS.n8422 DVSS.n1352 0.00658571
R36484 DVSS.n8416 DVSS.n1352 0.00658571
R36485 DVSS.n8416 DVSS.n8415 0.00658571
R36486 DVSS.n8415 DVSS.n8414 0.00658571
R36487 DVSS.n8414 DVSS.n1356 0.00658571
R36488 DVSS.n8408 DVSS.n1356 0.00658571
R36489 DVSS.n8408 DVSS.n8407 0.00658571
R36490 DVSS.n8407 DVSS.n8406 0.00658571
R36491 DVSS.n8406 DVSS.n1360 0.00658571
R36492 DVSS.n1395 DVSS.n1360 0.00658571
R36493 DVSS.n8397 DVSS.n1395 0.00658571
R36494 DVSS.n8397 DVSS.n8396 0.00658571
R36495 DVSS.n8396 DVSS.n8395 0.00658571
R36496 DVSS.n8395 DVSS.n1396 0.00658571
R36497 DVSS.n1638 DVSS.n1396 0.00658571
R36498 DVSS.n1639 DVSS.n1638 0.00658571
R36499 DVSS.n1639 DVSS.n1635 0.00658571
R36500 DVSS.n1645 DVSS.n1635 0.00658571
R36501 DVSS.n1646 DVSS.n1645 0.00658571
R36502 DVSS.n1647 DVSS.n1646 0.00658571
R36503 DVSS.n1647 DVSS.n1631 0.00658571
R36504 DVSS.n1653 DVSS.n1631 0.00658571
R36505 DVSS.n1654 DVSS.n1653 0.00658571
R36506 DVSS.n1655 DVSS.n1654 0.00658571
R36507 DVSS.n1655 DVSS.n1627 0.00658571
R36508 DVSS.n1661 DVSS.n1627 0.00658571
R36509 DVSS.n1662 DVSS.n1661 0.00658571
R36510 DVSS.n1663 DVSS.n1662 0.00658571
R36511 DVSS.n1663 DVSS.n1625 0.00658571
R36512 DVSS.n1669 DVSS.n1625 0.00658571
R36513 DVSS.n1670 DVSS.n1669 0.00658571
R36514 DVSS.n1671 DVSS.n1670 0.00658571
R36515 DVSS.n1671 DVSS.n1621 0.00658571
R36516 DVSS.n1677 DVSS.n1621 0.00658571
R36517 DVSS.n1678 DVSS.n1677 0.00658571
R36518 DVSS.n1679 DVSS.n1678 0.00658571
R36519 DVSS.n1679 DVSS.n1617 0.00658571
R36520 DVSS.n1685 DVSS.n1617 0.00658571
R36521 DVSS.n1686 DVSS.n1685 0.00658571
R36522 DVSS.n1687 DVSS.n1686 0.00658571
R36523 DVSS.n1687 DVSS.n1613 0.00658571
R36524 DVSS.n1693 DVSS.n1613 0.00658571
R36525 DVSS.n1694 DVSS.n1693 0.00658571
R36526 DVSS.n1695 DVSS.n1694 0.00658571
R36527 DVSS.n1695 DVSS.n1611 0.00658571
R36528 DVSS.n1701 DVSS.n1611 0.00658571
R36529 DVSS.n1702 DVSS.n1701 0.00658571
R36530 DVSS.n1703 DVSS.n1702 0.00658571
R36531 DVSS.n1703 DVSS.n1607 0.00658571
R36532 DVSS.n1709 DVSS.n1607 0.00658571
R36533 DVSS.n1710 DVSS.n1709 0.00658571
R36534 DVSS.n1711 DVSS.n1710 0.00658571
R36535 DVSS.n1711 DVSS.n1592 0.00658571
R36536 DVSS.n1730 DVSS.n1592 0.00658571
R36537 DVSS.n1731 DVSS.n1730 0.00658571
R36538 DVSS.n1733 DVSS.n1731 0.00658571
R36539 DVSS.n1733 DVSS.n1732 0.00658571
R36540 DVSS.n1732 DVSS.n1588 0.00658571
R36541 DVSS.n1740 DVSS.n1588 0.00658571
R36542 DVSS.n1743 DVSS.n1741 0.00658571
R36543 DVSS.n1942 DVSS.n1941 0.00658571
R36544 DVSS.n8050 DVSS.n1942 0.00658571
R36545 DVSS.n8050 DVSS.n8049 0.00658571
R36546 DVSS.n8049 DVSS.n8048 0.00658571
R36547 DVSS.n8048 DVSS.n1943 0.00658571
R36548 DVSS.n8042 DVSS.n1943 0.00658571
R36549 DVSS.n8042 DVSS.n8041 0.00658571
R36550 DVSS.n8041 DVSS.n8040 0.00658571
R36551 DVSS.n8040 DVSS.n1947 0.00658571
R36552 DVSS.n8027 DVSS.n1947 0.00658571
R36553 DVSS.n8027 DVSS.n8026 0.00658571
R36554 DVSS.n8026 DVSS.n8025 0.00658571
R36555 DVSS.n8025 DVSS.n1969 0.00658571
R36556 DVSS.n8019 DVSS.n1969 0.00658571
R36557 DVSS.n8019 DVSS.n8018 0.00658571
R36558 DVSS.n8018 DVSS.n8017 0.00658571
R36559 DVSS.n8017 DVSS.n1973 0.00658571
R36560 DVSS.n8004 DVSS.n1973 0.00658571
R36561 DVSS.n8004 DVSS.n8003 0.00658571
R36562 DVSS.n8003 DVSS.n8002 0.00658571
R36563 DVSS.n8002 DVSS.n1995 0.00658571
R36564 DVSS.n7996 DVSS.n1995 0.00658571
R36565 DVSS.n7996 DVSS.n7995 0.00658571
R36566 DVSS.n7995 DVSS.n7994 0.00658571
R36567 DVSS.n7994 DVSS.n1999 0.00658571
R36568 DVSS.n7988 DVSS.n1999 0.00658571
R36569 DVSS.n7988 DVSS.n7987 0.00658571
R36570 DVSS.n7987 DVSS.n7986 0.00658571
R36571 DVSS.n7986 DVSS.n2003 0.00658571
R36572 DVSS.n7980 DVSS.n2003 0.00658571
R36573 DVSS.n7980 DVSS.n7979 0.00658571
R36574 DVSS.n7979 DVSS.n7978 0.00658571
R36575 DVSS.n7978 DVSS.n2007 0.00658571
R36576 DVSS.n7965 DVSS.n2007 0.00658571
R36577 DVSS.n7965 DVSS.n7964 0.00658571
R36578 DVSS.n7964 DVSS.n7963 0.00658571
R36579 DVSS.n7963 DVSS.n2029 0.00658571
R36580 DVSS.n7957 DVSS.n2029 0.00658571
R36581 DVSS.n7957 DVSS.n7956 0.00658571
R36582 DVSS.n7956 DVSS.n7955 0.00658571
R36583 DVSS.n7955 DVSS.n2033 0.00658571
R36584 DVSS.n7949 DVSS.n2033 0.00658571
R36585 DVSS.n7949 DVSS.n7948 0.00658571
R36586 DVSS.n7948 DVSS.n7947 0.00658571
R36587 DVSS.n7947 DVSS.n2037 0.00658571
R36588 DVSS.n7941 DVSS.n2037 0.00658571
R36589 DVSS.n7941 DVSS.n7940 0.00658571
R36590 DVSS.n7940 DVSS.n7939 0.00658571
R36591 DVSS.n7939 DVSS.n2041 0.00658571
R36592 DVSS.n7767 DVSS.n2041 0.00658571
R36593 DVSS.n7767 DVSS.n7766 0.00658571
R36594 DVSS.n7772 DVSS.n7766 0.00658571
R36595 DVSS.n7773 DVSS.n7772 0.00658571
R36596 DVSS.n7774 DVSS.n7773 0.00658571
R36597 DVSS.n7774 DVSS.n7762 0.00658571
R36598 DVSS.n7780 DVSS.n7762 0.00658571
R36599 DVSS.n7781 DVSS.n7780 0.00658571
R36600 DVSS.n7782 DVSS.n7781 0.00658571
R36601 DVSS.n7782 DVSS.n7758 0.00658571
R36602 DVSS.n7788 DVSS.n7758 0.00658571
R36603 DVSS.n7789 DVSS.n7788 0.00658571
R36604 DVSS.n7791 DVSS.n7789 0.00658571
R36605 DVSS.n7791 DVSS.n7790 0.00658571
R36606 DVSS.n7790 DVSS.n7754 0.00658571
R36607 DVSS.n7798 DVSS.n7754 0.00658571
R36608 DVSS.n7799 DVSS.n7798 0.00658571
R36609 DVSS.n7841 DVSS.n7799 0.00658571
R36610 DVSS.n7841 DVSS.n7840 0.00658571
R36611 DVSS.n7840 DVSS.n7839 0.00658571
R36612 DVSS.n7839 DVSS.n7800 0.00658571
R36613 DVSS.n7833 DVSS.n7800 0.00658571
R36614 DVSS.n7833 DVSS.n7832 0.00658571
R36615 DVSS.n7832 DVSS.n7831 0.00658571
R36616 DVSS.n7831 DVSS.n7804 0.00658571
R36617 DVSS.n7825 DVSS.n7804 0.00658571
R36618 DVSS.n7825 DVSS.n7824 0.00658571
R36619 DVSS.n7824 DVSS.n7823 0.00658571
R36620 DVSS.n7823 DVSS.n7808 0.00658571
R36621 DVSS.n7817 DVSS.n7808 0.00658571
R36622 DVSS.n7817 DVSS.n7816 0.00658571
R36623 DVSS.n7816 DVSS.n7815 0.00658571
R36624 DVSS.n7815 DVSS.n7812 0.00658571
R36625 DVSS.n7812 DVSS.n1806 0.00658571
R36626 DVSS.n8126 DVSS.n1806 0.00658571
R36627 DVSS.n8127 DVSS.n8126 0.00658571
R36628 DVSS.n8128 DVSS.n8127 0.00658571
R36629 DVSS.n8128 DVSS.n1802 0.00658571
R36630 DVSS.n8134 DVSS.n1802 0.00658571
R36631 DVSS.n8135 DVSS.n8134 0.00658571
R36632 DVSS.n8136 DVSS.n8135 0.00658571
R36633 DVSS.n8136 DVSS.n1786 0.00658571
R36634 DVSS.n8155 DVSS.n1786 0.00658571
R36635 DVSS.n8156 DVSS.n8155 0.00658571
R36636 DVSS.n8157 DVSS.n8156 0.00658571
R36637 DVSS.n8157 DVSS.n1782 0.00658571
R36638 DVSS.n8163 DVSS.n1782 0.00658571
R36639 DVSS.n8164 DVSS.n8163 0.00658571
R36640 DVSS.n8169 DVSS.n1781 0.00658571
R36641 DVSS.n3082 DVSS.n3076 0.00658571
R36642 DVSS.n3083 DVSS.n3082 0.00658571
R36643 DVSS.n3085 DVSS.n3083 0.00658571
R36644 DVSS.n3085 DVSS.n3084 0.00658571
R36645 DVSS.n3084 DVSS.n3072 0.00658571
R36646 DVSS.n3092 DVSS.n3072 0.00658571
R36647 DVSS.n3093 DVSS.n3092 0.00658571
R36648 DVSS.n5826 DVSS.n3093 0.00658571
R36649 DVSS.n5826 DVSS.n5825 0.00658571
R36650 DVSS.n5825 DVSS.n5824 0.00658571
R36651 DVSS.n5824 DVSS.n3094 0.00658571
R36652 DVSS.n5818 DVSS.n3094 0.00658571
R36653 DVSS.n5818 DVSS.n5817 0.00658571
R36654 DVSS.n5817 DVSS.n5816 0.00658571
R36655 DVSS.n5816 DVSS.n3098 0.00658571
R36656 DVSS.n3124 DVSS.n3098 0.00658571
R36657 DVSS.n3125 DVSS.n3124 0.00658571
R36658 DVSS.n5806 DVSS.n3125 0.00658571
R36659 DVSS.n5806 DVSS.n5805 0.00658571
R36660 DVSS.n5805 DVSS.n5804 0.00658571
R36661 DVSS.n5804 DVSS.n3126 0.00658571
R36662 DVSS.n5798 DVSS.n3126 0.00658571
R36663 DVSS.n5798 DVSS.n5797 0.00658571
R36664 DVSS.n5797 DVSS.n5796 0.00658571
R36665 DVSS.n5796 DVSS.n3130 0.00658571
R36666 DVSS.n5790 DVSS.n3130 0.00658571
R36667 DVSS.n5790 DVSS.n5789 0.00658571
R36668 DVSS.n5789 DVSS.n5788 0.00658571
R36669 DVSS.n5788 DVSS.n3134 0.00658571
R36670 DVSS.n5782 DVSS.n3134 0.00658571
R36671 DVSS.n5782 DVSS.n5781 0.00658571
R36672 DVSS.n5781 DVSS.n5780 0.00658571
R36673 DVSS.n5780 DVSS.n3138 0.00658571
R36674 DVSS.n5770 DVSS.n3138 0.00658571
R36675 DVSS.n5770 DVSS.n5769 0.00658571
R36676 DVSS.n5769 DVSS.n5768 0.00658571
R36677 DVSS.n5768 DVSS.n3160 0.00658571
R36678 DVSS.n5762 DVSS.n3160 0.00658571
R36679 DVSS.n5762 DVSS.n5761 0.00658571
R36680 DVSS.n5761 DVSS.n5760 0.00658571
R36681 DVSS.n5760 DVSS.n3164 0.00658571
R36682 DVSS.n5754 DVSS.n3164 0.00658571
R36683 DVSS.n5754 DVSS.n5753 0.00658571
R36684 DVSS.n5753 DVSS.n5752 0.00658571
R36685 DVSS.n5752 DVSS.n3168 0.00658571
R36686 DVSS.n5746 DVSS.n3168 0.00658571
R36687 DVSS.n5746 DVSS.n5745 0.00658571
R36688 DVSS.n5745 DVSS.n5744 0.00658571
R36689 DVSS.n5744 DVSS.n3172 0.00658571
R36690 DVSS.n5034 DVSS.n3172 0.00658571
R36691 DVSS.n5035 DVSS.n5034 0.00658571
R36692 DVSS.n5191 DVSS.n5035 0.00658571
R36693 DVSS.n5191 DVSS.n5190 0.00658571
R36694 DVSS.n5190 DVSS.n5189 0.00658571
R36695 DVSS.n5189 DVSS.n5036 0.00658571
R36696 DVSS.n5183 DVSS.n5036 0.00658571
R36697 DVSS.n5183 DVSS.n5182 0.00658571
R36698 DVSS.n5182 DVSS.n5181 0.00658571
R36699 DVSS.n5181 DVSS.n5041 0.00658571
R36700 DVSS.n5175 DVSS.n5041 0.00658571
R36701 DVSS.n5175 DVSS.n5174 0.00658571
R36702 DVSS.n5174 DVSS.n5173 0.00658571
R36703 DVSS.n5173 DVSS.n5045 0.00658571
R36704 DVSS.n5167 DVSS.n5045 0.00658571
R36705 DVSS.n5167 DVSS.n5166 0.00658571
R36706 DVSS.n5166 DVSS.n5165 0.00658571
R36707 DVSS.n5165 DVSS.n5049 0.00658571
R36708 DVSS.n5159 DVSS.n5049 0.00658571
R36709 DVSS.n5159 DVSS.n5158 0.00658571
R36710 DVSS.n5158 DVSS.n5157 0.00658571
R36711 DVSS.n5157 DVSS.n5051 0.00658571
R36712 DVSS.n5151 DVSS.n5051 0.00658571
R36713 DVSS.n5151 DVSS.n5150 0.00658571
R36714 DVSS.n5150 DVSS.n5149 0.00658571
R36715 DVSS.n5149 DVSS.n5055 0.00658571
R36716 DVSS.n5143 DVSS.n5055 0.00658571
R36717 DVSS.n5143 DVSS.n5142 0.00658571
R36718 DVSS.n5142 DVSS.n5141 0.00658571
R36719 DVSS.n5141 DVSS.n5059 0.00658571
R36720 DVSS.n5135 DVSS.n5059 0.00658571
R36721 DVSS.n5135 DVSS.n5134 0.00658571
R36722 DVSS.n5134 DVSS.n5133 0.00658571
R36723 DVSS.n5133 DVSS.n5063 0.00658571
R36724 DVSS.n5085 DVSS.n5063 0.00658571
R36725 DVSS.n5125 DVSS.n5085 0.00658571
R36726 DVSS.n5125 DVSS.n5124 0.00658571
R36727 DVSS.n5124 DVSS.n5123 0.00658571
R36728 DVSS.n5123 DVSS.n5086 0.00658571
R36729 DVSS.n5117 DVSS.n5086 0.00658571
R36730 DVSS.n5117 DVSS.n5116 0.00658571
R36731 DVSS.n5116 DVSS.n5115 0.00658571
R36732 DVSS.n5115 DVSS.n5090 0.00658571
R36733 DVSS.n5110 DVSS.n5090 0.00658571
R36734 DVSS.n5110 DVSS.n5109 0.00658571
R36735 DVSS.n5109 DVSS.n5108 0.00658571
R36736 DVSS.n5108 DVSS.n5092 0.00658571
R36737 DVSS.n5101 DVSS.n5092 0.00658571
R36738 DVSS.n5100 DVSS.n5099 0.00658571
R36739 DVSS.n5850 DVSS.n5849 0.00658571
R36740 DVSS.n5849 DVSS.n5848 0.00658571
R36741 DVSS.n5848 DVSS.n3037 0.00658571
R36742 DVSS.n5842 DVSS.n3037 0.00658571
R36743 DVSS.n5842 DVSS.n5841 0.00658571
R36744 DVSS.n5841 DVSS.n5840 0.00658571
R36745 DVSS.n5840 DVSS.n3041 0.00658571
R36746 DVSS.n3902 DVSS.n3041 0.00658571
R36747 DVSS.n3906 DVSS.n3902 0.00658571
R36748 DVSS.n3907 DVSS.n3906 0.00658571
R36749 DVSS.n3908 DVSS.n3907 0.00658571
R36750 DVSS.n3908 DVSS.n3898 0.00658571
R36751 DVSS.n3914 DVSS.n3898 0.00658571
R36752 DVSS.n3915 DVSS.n3914 0.00658571
R36753 DVSS.n4170 DVSS.n3915 0.00658571
R36754 DVSS.n4170 DVSS.n4169 0.00658571
R36755 DVSS.n4169 DVSS.n4168 0.00658571
R36756 DVSS.n4168 DVSS.n3916 0.00658571
R36757 DVSS.n3920 DVSS.n3916 0.00658571
R36758 DVSS.n4160 DVSS.n3920 0.00658571
R36759 DVSS.n4160 DVSS.n4159 0.00658571
R36760 DVSS.n4159 DVSS.n4158 0.00658571
R36761 DVSS.n4158 DVSS.n3921 0.00658571
R36762 DVSS.n4152 DVSS.n3921 0.00658571
R36763 DVSS.n4152 DVSS.n4151 0.00658571
R36764 DVSS.n4151 DVSS.n4150 0.00658571
R36765 DVSS.n4150 DVSS.n3925 0.00658571
R36766 DVSS.n4144 DVSS.n3925 0.00658571
R36767 DVSS.n4144 DVSS.n4143 0.00658571
R36768 DVSS.n4143 DVSS.n4142 0.00658571
R36769 DVSS.n4142 DVSS.n3929 0.00658571
R36770 DVSS.n3953 DVSS.n3929 0.00658571
R36771 DVSS.n4134 DVSS.n3953 0.00658571
R36772 DVSS.n4134 DVSS.n4133 0.00658571
R36773 DVSS.n4133 DVSS.n4132 0.00658571
R36774 DVSS.n4132 DVSS.n3954 0.00658571
R36775 DVSS.n4126 DVSS.n3954 0.00658571
R36776 DVSS.n4126 DVSS.n4125 0.00658571
R36777 DVSS.n4125 DVSS.n4124 0.00658571
R36778 DVSS.n4124 DVSS.n3959 0.00658571
R36779 DVSS.n4118 DVSS.n3959 0.00658571
R36780 DVSS.n4118 DVSS.n4117 0.00658571
R36781 DVSS.n4117 DVSS.n4116 0.00658571
R36782 DVSS.n4116 DVSS.n3963 0.00658571
R36783 DVSS.n4110 DVSS.n3963 0.00658571
R36784 DVSS.n4110 DVSS.n4109 0.00658571
R36785 DVSS.n4109 DVSS.n4108 0.00658571
R36786 DVSS.n4108 DVSS.n3967 0.00658571
R36787 DVSS.n3995 DVSS.n3967 0.00658571
R36788 DVSS.n3995 DVSS.n3472 0.00658571
R36789 DVSS.n5240 DVSS.n3472 0.00658571
R36790 DVSS.n5241 DVSS.n5240 0.00658571
R36791 DVSS.n5242 DVSS.n5241 0.00658571
R36792 DVSS.n5242 DVSS.n3468 0.00658571
R36793 DVSS.n5248 DVSS.n3468 0.00658571
R36794 DVSS.n5249 DVSS.n5248 0.00658571
R36795 DVSS.n5250 DVSS.n5249 0.00658571
R36796 DVSS.n5250 DVSS.n3464 0.00658571
R36797 DVSS.n5256 DVSS.n3464 0.00658571
R36798 DVSS.n5257 DVSS.n5256 0.00658571
R36799 DVSS.n5258 DVSS.n5257 0.00658571
R36800 DVSS.n5258 DVSS.n3460 0.00658571
R36801 DVSS.n5264 DVSS.n3460 0.00658571
R36802 DVSS.n5265 DVSS.n5264 0.00658571
R36803 DVSS.n5266 DVSS.n5265 0.00658571
R36804 DVSS.n5266 DVSS.n3438 0.00658571
R36805 DVSS.n5275 DVSS.n3438 0.00658571
R36806 DVSS.n5276 DVSS.n5275 0.00658571
R36807 DVSS.n5277 DVSS.n5276 0.00658571
R36808 DVSS.n5277 DVSS.n3434 0.00658571
R36809 DVSS.n5283 DVSS.n3434 0.00658571
R36810 DVSS.n5284 DVSS.n5283 0.00658571
R36811 DVSS.n5285 DVSS.n5284 0.00658571
R36812 DVSS.n5285 DVSS.n3430 0.00658571
R36813 DVSS.n5291 DVSS.n3430 0.00658571
R36814 DVSS.n5292 DVSS.n5291 0.00658571
R36815 DVSS.n5293 DVSS.n5292 0.00658571
R36816 DVSS.n5293 DVSS.n3426 0.00658571
R36817 DVSS.n5299 DVSS.n3426 0.00658571
R36818 DVSS.n5300 DVSS.n5299 0.00658571
R36819 DVSS.n5301 DVSS.n5300 0.00658571
R36820 DVSS.n5301 DVSS.n3403 0.00658571
R36821 DVSS.n5310 DVSS.n3403 0.00658571
R36822 DVSS.n5311 DVSS.n5310 0.00658571
R36823 DVSS.n5312 DVSS.n5311 0.00658571
R36824 DVSS.n5312 DVSS.n3399 0.00658571
R36825 DVSS.n5319 DVSS.n3399 0.00658571
R36826 DVSS.n5320 DVSS.n5319 0.00658571
R36827 DVSS.n5321 DVSS.n5320 0.00658571
R36828 DVSS.n5321 DVSS.n3397 0.00658571
R36829 DVSS.n5326 DVSS.n3397 0.00658571
R36830 DVSS.n5327 DVSS.n5326 0.00658571
R36831 DVSS.n5345 DVSS.n5327 0.00658571
R36832 DVSS.n5345 DVSS.n5344 0.00658571
R36833 DVSS.n5344 DVSS.n5343 0.00658571
R36834 DVSS.n5343 DVSS.n5328 0.00658571
R36835 DVSS.n5337 DVSS.n5328 0.00658571
R36836 DVSS.n5336 DVSS.n5335 0.00658571
R36837 DVSS.n6637 DVSS.n6636 0.00658571
R36838 DVSS.n6636 DVSS.n6635 0.00658571
R36839 DVSS.n6635 DVSS.n6021 0.00658571
R36840 DVSS.n6629 DVSS.n6021 0.00658571
R36841 DVSS.n6629 DVSS.n6628 0.00658571
R36842 DVSS.n6628 DVSS.n6627 0.00658571
R36843 DVSS.n6627 DVSS.n6026 0.00658571
R36844 DVSS.n6621 DVSS.n6026 0.00658571
R36845 DVSS.n6621 DVSS.n6620 0.00658571
R36846 DVSS.n6620 DVSS.n6619 0.00658571
R36847 DVSS.n6619 DVSS.n6030 0.00658571
R36848 DVSS.n6613 DVSS.n6030 0.00658571
R36849 DVSS.n6613 DVSS.n6612 0.00658571
R36850 DVSS.n6612 DVSS.n6611 0.00658571
R36851 DVSS.n6611 DVSS.n6350 0.00658571
R36852 DVSS.n6605 DVSS.n6350 0.00658571
R36853 DVSS.n6605 DVSS.n6604 0.00658571
R36854 DVSS.n6604 DVSS.n6603 0.00658571
R36855 DVSS.n6603 DVSS.n6354 0.00658571
R36856 DVSS.n6597 DVSS.n6354 0.00658571
R36857 DVSS.n6597 DVSS.n6596 0.00658571
R36858 DVSS.n6596 DVSS.n6595 0.00658571
R36859 DVSS.n6595 DVSS.n6358 0.00658571
R36860 DVSS.n6589 DVSS.n6358 0.00658571
R36861 DVSS.n6589 DVSS.n6588 0.00658571
R36862 DVSS.n6588 DVSS.n6587 0.00658571
R36863 DVSS.n6587 DVSS.n6362 0.00658571
R36864 DVSS.n6581 DVSS.n6362 0.00658571
R36865 DVSS.n6581 DVSS.n6580 0.00658571
R36866 DVSS.n6580 DVSS.n6579 0.00658571
R36867 DVSS.n6579 DVSS.n6366 0.00658571
R36868 DVSS.n6573 DVSS.n6366 0.00658571
R36869 DVSS.n6573 DVSS.n6572 0.00658571
R36870 DVSS.n6572 DVSS.n6571 0.00658571
R36871 DVSS.n6571 DVSS.n6370 0.00658571
R36872 DVSS.n6565 DVSS.n6370 0.00658571
R36873 DVSS.n6565 DVSS.n6564 0.00658571
R36874 DVSS.n6564 DVSS.n6563 0.00658571
R36875 DVSS.n6563 DVSS.n6374 0.00658571
R36876 DVSS.n6557 DVSS.n6374 0.00658571
R36877 DVSS.n6557 DVSS.n6556 0.00658571
R36878 DVSS.n6556 DVSS.n6555 0.00658571
R36879 DVSS.n6555 DVSS.n6378 0.00658571
R36880 DVSS.n6549 DVSS.n6378 0.00658571
R36881 DVSS.n6549 DVSS.n6548 0.00658571
R36882 DVSS.n6548 DVSS.n6547 0.00658571
R36883 DVSS.n6547 DVSS.n6382 0.00658571
R36884 DVSS.n6541 DVSS.n6382 0.00658571
R36885 DVSS.n6541 DVSS.n6540 0.00658571
R36886 DVSS.n6540 DVSS.n6539 0.00658571
R36887 DVSS.n6539 DVSS.n6386 0.00658571
R36888 DVSS.n6533 DVSS.n6386 0.00658571
R36889 DVSS.n6533 DVSS.n6532 0.00658571
R36890 DVSS.n6532 DVSS.n6531 0.00658571
R36891 DVSS.n6531 DVSS.n6390 0.00658571
R36892 DVSS.n6525 DVSS.n6390 0.00658571
R36893 DVSS.n6525 DVSS.n6524 0.00658571
R36894 DVSS.n6524 DVSS.n6523 0.00658571
R36895 DVSS.n6523 DVSS.n6394 0.00658571
R36896 DVSS.n6517 DVSS.n6394 0.00658571
R36897 DVSS.n6517 DVSS.n6516 0.00658571
R36898 DVSS.n6516 DVSS.n6515 0.00658571
R36899 DVSS.n6515 DVSS.n6398 0.00658571
R36900 DVSS.n6509 DVSS.n6398 0.00658571
R36901 DVSS.n6509 DVSS.n6508 0.00658571
R36902 DVSS.n6508 DVSS.n6507 0.00658571
R36903 DVSS.n6507 DVSS.n6402 0.00658571
R36904 DVSS.n6501 DVSS.n6402 0.00658571
R36905 DVSS.n6501 DVSS.n6500 0.00658571
R36906 DVSS.n6500 DVSS.n6499 0.00658571
R36907 DVSS.n6499 DVSS.n6406 0.00658571
R36908 DVSS.n6493 DVSS.n6406 0.00658571
R36909 DVSS.n6493 DVSS.n6492 0.00658571
R36910 DVSS.n6492 DVSS.n6491 0.00658571
R36911 DVSS.n6491 DVSS.n6410 0.00658571
R36912 DVSS.n6485 DVSS.n6410 0.00658571
R36913 DVSS.n6485 DVSS.n6484 0.00658571
R36914 DVSS.n6484 DVSS.n6483 0.00658571
R36915 DVSS.n6483 DVSS.n6414 0.00658571
R36916 DVSS.n6477 DVSS.n6414 0.00658571
R36917 DVSS.n6477 DVSS.n6476 0.00658571
R36918 DVSS.n6476 DVSS.n6475 0.00658571
R36919 DVSS.n6475 DVSS.n6418 0.00658571
R36920 DVSS.n6469 DVSS.n6418 0.00658571
R36921 DVSS.n6469 DVSS.n6468 0.00658571
R36922 DVSS.n6468 DVSS.n6467 0.00658571
R36923 DVSS.n6467 DVSS.n6422 0.00658571
R36924 DVSS.n6461 DVSS.n6422 0.00658571
R36925 DVSS.n6461 DVSS.n6460 0.00658571
R36926 DVSS.n6460 DVSS.n6459 0.00658571
R36927 DVSS.n6459 DVSS.n6426 0.00658571
R36928 DVSS.n6453 DVSS.n6426 0.00658571
R36929 DVSS.n6453 DVSS.n6452 0.00658571
R36930 DVSS.n6452 DVSS.n6451 0.00658571
R36931 DVSS.n6451 DVSS.n6430 0.00658571
R36932 DVSS.n6445 DVSS.n6430 0.00658571
R36933 DVSS.n6445 DVSS.n6444 0.00658571
R36934 DVSS.n6438 DVSS.n6435 0.00658571
R36935 DVSS.n6050 DVSS.n6049 0.00658571
R36936 DVSS.n6050 DVSS.n6041 0.00658571
R36937 DVSS.n6056 DVSS.n6041 0.00658571
R36938 DVSS.n6057 DVSS.n6056 0.00658571
R36939 DVSS.n6058 DVSS.n6057 0.00658571
R36940 DVSS.n6058 DVSS.n6037 0.00658571
R36941 DVSS.n6064 DVSS.n6037 0.00658571
R36942 DVSS.n6065 DVSS.n6064 0.00658571
R36943 DVSS.n6341 DVSS.n6065 0.00658571
R36944 DVSS.n6341 DVSS.n6340 0.00658571
R36945 DVSS.n6340 DVSS.n6339 0.00658571
R36946 DVSS.n6339 DVSS.n6066 0.00658571
R36947 DVSS.n6333 DVSS.n6066 0.00658571
R36948 DVSS.n6333 DVSS.n6332 0.00658571
R36949 DVSS.n6332 DVSS.n6331 0.00658571
R36950 DVSS.n6331 DVSS.n6071 0.00658571
R36951 DVSS.n6325 DVSS.n6071 0.00658571
R36952 DVSS.n6325 DVSS.n6324 0.00658571
R36953 DVSS.n6324 DVSS.n6323 0.00658571
R36954 DVSS.n6323 DVSS.n6075 0.00658571
R36955 DVSS.n6317 DVSS.n6075 0.00658571
R36956 DVSS.n6317 DVSS.n6316 0.00658571
R36957 DVSS.n6316 DVSS.n6315 0.00658571
R36958 DVSS.n6315 DVSS.n6079 0.00658571
R36959 DVSS.n6309 DVSS.n6079 0.00658571
R36960 DVSS.n6309 DVSS.n6308 0.00658571
R36961 DVSS.n6308 DVSS.n6307 0.00658571
R36962 DVSS.n6307 DVSS.n6083 0.00658571
R36963 DVSS.n6301 DVSS.n6083 0.00658571
R36964 DVSS.n6301 DVSS.n6300 0.00658571
R36965 DVSS.n6300 DVSS.n6299 0.00658571
R36966 DVSS.n6299 DVSS.n6087 0.00658571
R36967 DVSS.n6293 DVSS.n6087 0.00658571
R36968 DVSS.n6293 DVSS.n6292 0.00658571
R36969 DVSS.n6292 DVSS.n6291 0.00658571
R36970 DVSS.n6291 DVSS.n6091 0.00658571
R36971 DVSS.n6285 DVSS.n6091 0.00658571
R36972 DVSS.n6285 DVSS.n6284 0.00658571
R36973 DVSS.n6284 DVSS.n6283 0.00658571
R36974 DVSS.n6283 DVSS.n6095 0.00658571
R36975 DVSS.n6277 DVSS.n6095 0.00658571
R36976 DVSS.n6277 DVSS.n6276 0.00658571
R36977 DVSS.n6276 DVSS.n6275 0.00658571
R36978 DVSS.n6275 DVSS.n6099 0.00658571
R36979 DVSS.n6269 DVSS.n6099 0.00658571
R36980 DVSS.n6269 DVSS.n6268 0.00658571
R36981 DVSS.n6268 DVSS.n6267 0.00658571
R36982 DVSS.n6267 DVSS.n6103 0.00658571
R36983 DVSS.n6261 DVSS.n6103 0.00658571
R36984 DVSS.n6261 DVSS.n6260 0.00658571
R36985 DVSS.n6260 DVSS.n6259 0.00658571
R36986 DVSS.n6259 DVSS.n6107 0.00658571
R36987 DVSS.n6253 DVSS.n6107 0.00658571
R36988 DVSS.n6253 DVSS.n6252 0.00658571
R36989 DVSS.n6252 DVSS.n6251 0.00658571
R36990 DVSS.n6251 DVSS.n6111 0.00658571
R36991 DVSS.n6245 DVSS.n6111 0.00658571
R36992 DVSS.n6245 DVSS.n6244 0.00658571
R36993 DVSS.n6244 DVSS.n6243 0.00658571
R36994 DVSS.n6243 DVSS.n6115 0.00658571
R36995 DVSS.n6237 DVSS.n6115 0.00658571
R36996 DVSS.n6237 DVSS.n6236 0.00658571
R36997 DVSS.n6236 DVSS.n6235 0.00658571
R36998 DVSS.n6235 DVSS.n6119 0.00658571
R36999 DVSS.n6229 DVSS.n6119 0.00658571
R37000 DVSS.n6229 DVSS.n6228 0.00658571
R37001 DVSS.n6228 DVSS.n6227 0.00658571
R37002 DVSS.n6227 DVSS.n6123 0.00658571
R37003 DVSS.n6221 DVSS.n6123 0.00658571
R37004 DVSS.n6221 DVSS.n6220 0.00658571
R37005 DVSS.n6220 DVSS.n6219 0.00658571
R37006 DVSS.n6219 DVSS.n6127 0.00658571
R37007 DVSS.n6213 DVSS.n6127 0.00658571
R37008 DVSS.n6213 DVSS.n6212 0.00658571
R37009 DVSS.n6212 DVSS.n6211 0.00658571
R37010 DVSS.n6211 DVSS.n6131 0.00658571
R37011 DVSS.n6205 DVSS.n6131 0.00658571
R37012 DVSS.n6205 DVSS.n6204 0.00658571
R37013 DVSS.n6204 DVSS.n6203 0.00658571
R37014 DVSS.n6203 DVSS.n6135 0.00658571
R37015 DVSS.n6197 DVSS.n6135 0.00658571
R37016 DVSS.n6197 DVSS.n6196 0.00658571
R37017 DVSS.n6196 DVSS.n6195 0.00658571
R37018 DVSS.n6195 DVSS.n6139 0.00658571
R37019 DVSS.n6189 DVSS.n6139 0.00658571
R37020 DVSS.n6189 DVSS.n6188 0.00658571
R37021 DVSS.n6188 DVSS.n6187 0.00658571
R37022 DVSS.n6187 DVSS.n6143 0.00658571
R37023 DVSS.n6181 DVSS.n6143 0.00658571
R37024 DVSS.n6181 DVSS.n6180 0.00658571
R37025 DVSS.n6180 DVSS.n6179 0.00658571
R37026 DVSS.n6179 DVSS.n6147 0.00658571
R37027 DVSS.n6173 DVSS.n6147 0.00658571
R37028 DVSS.n6173 DVSS.n6172 0.00658571
R37029 DVSS.n6172 DVSS.n6171 0.00658571
R37030 DVSS.n6171 DVSS.n6151 0.00658571
R37031 DVSS.n6165 DVSS.n6151 0.00658571
R37032 DVSS.n6164 DVSS.n6163 0.00658571
R37033 DVSS.n9088 DVSS.n9087 0.0065
R37034 DVSS.n9176 DVSS.n237 0.0065
R37035 DVSS.n7032 DVSS.n949 0.0065
R37036 DVSS.n8813 DVSS.n8811 0.0065
R37037 DVSS.n270 DVSS.n162 0.0065
R37038 DVSS.n8813 DVSS.n8812 0.0065
R37039 DVSS.n7033 DVSS.n7032 0.0065
R37040 DVSS.n9180 DVSS.n9179 0.0065
R37041 DVSS.n9180 DVSS.n486 0.0065
R37042 DVSS.n270 DVSS.n269 0.0065
R37043 DVSS.n8600 DVSS.n950 0.0065
R37044 DVSS.n9087 DVSS.n630 0.0065
R37045 DVSS.n9284 DVSS.n237 0.0065
R37046 DVSS.n9868 DVSS.n63 0.0065
R37047 DVSS.n9869 DVSS.n9868 0.0065
R37048 DVSS.n8600 DVSS.n8599 0.0065
R37049 DVSS.n4492 DVSS.n3830 0.00648592
R37050 DVSS.n4519 DVSS.n3811 0.00648592
R37051 DVSS.n4572 DVSS.n3800 0.00648592
R37052 DVSS.n4776 DVSS.n3728 0.00648592
R37053 DVSS.n6744 DVSS.n6736 0.00647857
R37054 DVSS.n6689 DVSS.n6675 0.00647857
R37055 DVSS.n1171 DVSS.n1161 0.00647857
R37056 DVSS.n8435 DVSS.n1334 0.00647857
R37057 DVSS.n1925 DVSS.n1917 0.00647857
R37058 DVSS.n1950 DVSS.n1949 0.00647857
R37059 DVSS.n1976 DVSS.n1975 0.00647857
R37060 DVSS.n2010 DVSS.n2009 0.00647857
R37061 DVSS.n3003 DVSS.n2994 0.00647857
R37062 DVSS.n3117 DVSS.n3105 0.00647857
R37063 DVSS.n3141 DVSS.n3140 0.00647857
R37064 DVSS.n5854 DVSS.n3027 0.00647857
R37065 DVSS.n4172 DVSS.n3887 0.00647857
R37066 DVSS.n3946 DVSS.n3936 0.00647857
R37067 DVSS.n3856 DVSS.n3845 0.00647857
R37068 DVSS.n4252 DVSS.n4223 0.00647857
R37069 DVSS.n4418 DVSS.n4199 0.00647857
R37070 DVSS.n3726 DVSS.n3719 0.00647857
R37071 DVSS.n1270 DVSS.n569 0.00641549
R37072 DVSS.n1279 DVSS.n597 0.00641549
R37073 DVSS.n4937 DVSS 0.00641429
R37074 DVSS.n1741 DVSS 0.00641429
R37075 DVSS.n8393 DVSS.n1398 0.00641429
R37076 DVSS DVSS.n1781 0.00641429
R37077 DVSS.n7901 DVSS.n2068 0.00641429
R37078 DVSS DVSS.n5100 0.00641429
R37079 DVSS.n5196 DVSS.n5016 0.00641429
R37080 DVSS DVSS.n5336 0.00641429
R37081 DVSS.n5238 DVSS.n3474 0.00641429
R37082 DVSS.n4817 DVSS.n3683 0.00641429
R37083 DVSS.n6435 VSS 0.00641429
R37084 VSS DVSS.n6164 0.00641429
R37085 DVSS.n8907 DVSS.n775 0.00634646
R37086 DVSS.n9441 DVSS.n359 0.00634646
R37087 DVSS.n8348 DVSS.n1428 0.00622143
R37088 DVSS.n1667 DVSS.n1427 0.00622143
R37089 DVSS.n8489 DVSS.n1108 0.00622143
R37090 DVSS.n1699 DVSS.n1107 0.00622143
R37091 DVSS.n1724 DVSS.n1601 0.00622143
R37092 DVSS.n1728 DVSS.n1594 0.00622143
R37093 DVSS.n1748 DVSS.n1565 0.00622143
R37094 DVSS.n1586 DVSS.n1564 0.00622143
R37095 DVSS.n7846 DVSS.n7731 0.00622143
R37096 DVSS.n7752 DVSS.n7730 0.00622143
R37097 DVSS.n8121 DVSS.n1816 0.00622143
R37098 DVSS.n8124 DVSS.n1808 0.00622143
R37099 DVSS.n8149 DVSS.n1796 0.00622143
R37100 DVSS.n8153 DVSS.n1788 0.00622143
R37101 DVSS.n8178 DVSS.n1764 0.00622143
R37102 DVSS.n1779 DVSS.n1763 0.00622143
R37103 DVSS.n5047 DVSS.n3326 0.00622143
R37104 DVSS.n3328 DVSS.n3325 0.00622143
R37105 DVSS.n5065 DVSS.n5061 0.00622143
R37106 DVSS.n5074 DVSS.n5073 0.00622143
R37107 DVSS.n5119 DVSS.n3372 0.00622143
R37108 DVSS.n3374 DVSS.n3371 0.00622143
R37109 DVSS.n5912 DVSS.n2943 0.00622143
R37110 DVSS.n5095 DVSS.n2942 0.00622143
R37111 DVSS.n5270 DVSS.n5268 0.00622143
R37112 DVSS.n5272 DVSS.n3446 0.00622143
R37113 DVSS.n5305 DVSS.n5303 0.00622143
R37114 DVSS.n5307 DVSS.n3411 0.00622143
R37115 DVSS.n5353 DVSS.n3380 0.00622143
R37116 DVSS.n3393 DVSS.n3379 0.00622143
R37117 DVSS.n5915 DVSS.n2925 0.00622143
R37118 DVSS.n5331 DVSS.n2924 0.00622143
R37119 DVSS.n4848 DVSS.n3656 0.00622143
R37120 DVSS.n4851 DVSS.n3647 0.00622143
R37121 DVSS.n4886 DVSS.n3627 0.00622143
R37122 DVSS.n4889 DVSS.n3614 0.00622143
R37123 DVSS.n4972 DVSS.n3601 0.00622143
R37124 DVSS.n4955 DVSS.n3600 0.00622143
R37125 DVSS.n4945 DVSS.n4944 0.00622143
R37126 DVSS.n4942 DVSS.n4941 0.00622143
R37127 DVSS.n5551 DVSS.n2292 0.00620423
R37128 DVSS.n7903 DVSS.n7902 0.00620423
R37129 DVSS.n5626 DVSS.n2322 0.00620423
R37130 DVSS.n7935 DVSS.n7934 0.00620423
R37131 DVSS.n6343 DVSS.n6033 0.00609286
R37132 DVSS.n6347 DVSS.n6032 0.00609286
R37133 DVSS.n8915 DVSS.n777 0.00599213
R37134 DVSS.n8950 DVSS.n736 0.00599213
R37135 DVSS.n9449 DVSS.n361 0.00599213
R37136 DVSS.n9484 DVSS.n35 0.00599213
R37137 DVSS.n6854 DVSS.n6850 0.00596429
R37138 DVSS.n6832 DVSS.n6667 0.00596429
R37139 DVSS.n6817 DVSS.n1162 0.00596429
R37140 DVSS.n8428 DVSS.n1326 0.00596429
R37141 DVSS.n8056 DVSS.n8052 0.00596429
R37142 DVSS.n8034 DVSS.n8029 0.00596429
R37143 DVSS.n8011 DVSS.n8006 0.00596429
R37144 DVSS.n7972 DVSS.n7967 0.00596429
R37145 DVSS.n3074 DVSS.n2995 0.00596429
R37146 DVSS.n5811 DVSS.n5808 0.00596429
R37147 DVSS.n5775 DVSS.n5772 0.00596429
R37148 DVSS.n5846 DVSS.n3028 0.00596429
R37149 DVSS.n4164 DVSS.n3888 0.00596429
R37150 DVSS.n3956 DVSS.n3950 0.00596429
R37151 DVSS.n4232 DVSS.n3837 0.00596429
R37152 DVSS.n4260 DVSS.n4211 0.00596429
R37153 DVSS.n4410 DVSS.n4200 0.00596429
R37154 DVSS.n4379 DVSS.n3720 0.00596429
R37155 DVSS.n5938 DVSS.n5936 0.00591803
R37156 DVSS.n4480 DVSS.n4479 0.00591803
R37157 DVSS.n5015 DVSS.n3516 0.00578169
R37158 DVSS.n5571 DVSS.n2301 0.00578169
R37159 DVSS.n515 DVSS.n372 0.00578169
R37160 DVSS.n5204 DVSS.n3180 0.00578169
R37161 DVSS.n5584 DVSS.n2331 0.00578169
R37162 DVSS.n8862 DVSS.n648 0.00578169
R37163 DVSS.n4489 DVSS.n3834 0.00578169
R37164 DVSS.n4516 DVSS.n3815 0.00578169
R37165 DVSS.n4576 DVSS.n3801 0.00578169
R37166 DVSS.n4781 DVSS.n3729 0.00578169
R37167 DVSS.n5831 DVSS.n3056 0.00570714
R37168 DVSS.n5838 DVSS.n5837 0.00570714
R37169 DVSS.n8923 DVSS.n761 0.0056378
R37170 DVSS.n8958 DVSS.n741 0.0056378
R37171 DVSS.n9457 DVSS.n346 0.0056378
R37172 DVSS.n9492 DVSS.n39 0.0056378
R37173 DVSS.n5829 DVSS.n5828 0.00557857
R37174 DVSS.n5834 DVSS.n3054 0.00557857
R37175 DVSS.n6000 DVSS.n2789 0.0055
R37176 DVSS.n6000 DVSS.n5999 0.0055
R37177 DVSS.n5973 DVSS.n2822 0.0055
R37178 DVSS.n5973 DVSS.n5972 0.0055
R37179 DVSS.n5958 DVSS.n2853 0.0055
R37180 DVSS.n5958 DVSS.n5955 0.0055
R37181 DVSS.n5941 DVSS.n2882 0.0055
R37182 DVSS.n5941 DVSS.n5940 0.0055
R37183 DVSS.n4940 DVSS.n4939 0.00548841
R37184 DVSS.n4235 DVSS.n3839 0.00548841
R37185 DVSS.n1742 DVSS.n1587 0.00548841
R37186 DVSS.n6766 DVSS.n6738 0.00548841
R37187 DVSS.n8170 DVSS.n1780 0.00548841
R37188 DVSS.n1938 DVSS.n1919 0.00548841
R37189 DVSS.n5096 DVSS.n5094 0.00548841
R37190 DVSS.n3077 DVSS.n2997 0.00548841
R37191 DVSS.n5332 DVSS.n5330 0.00548841
R37192 DVSS.n5853 DVSS.n3030 0.00548841
R37193 DVSS.n6437 DVSS.n6434 0.00548841
R37194 DVSS.n6639 DVSS.n6018 0.00548841
R37195 DVSS.n6156 DVSS.n6155 0.00548841
R37196 DVSS.n6048 DVSS.n6047 0.00548841
R37197 DVSS.n1259 DVSS.n179 0.00546063
R37198 DVSS.n1264 DVSS.n218 0.00546063
R37199 DVSS.n1284 DVSS.n1075 0.00546063
R37200 DVSS.n1289 DVSS.n1205 0.00546063
R37201 DVSS.n3485 DVSS.n3475 0.00535915
R37202 DVSS.n5574 DVSS.n2282 0.00535915
R37203 DVSS.n3971 DVSS.n3970 0.00535915
R37204 DVSS.n5578 DVSS.n2312 0.00535915
R37205 DVSS.n6767 DVSS.n6737 0.00532143
R37206 DVSS.n6836 DVSS.n6668 0.00532143
R37207 DVSS.n6822 DVSS.n1163 0.00532143
R37208 DVSS.n8434 DVSS.n1327 0.00532143
R37209 DVSS.n1939 DVSS.n1918 0.00532143
R37210 DVSS.n8038 DVSS.n8037 0.00532143
R37211 DVSS.n8015 DVSS.n8014 0.00532143
R37212 DVSS.n7976 DVSS.n7975 0.00532143
R37213 DVSS.n3078 DVSS.n2996 0.00532143
R37214 DVSS.n3122 DVSS.n3112 0.00532143
R37215 DVSS.n5778 DVSS.n5777 0.00532143
R37216 DVSS.n5851 DVSS.n3029 0.00532143
R37217 DVSS.n3896 DVSS.n3889 0.00532143
R37218 DVSS.n4137 DVSS.n3947 0.00532143
R37219 DVSS.n4236 DVSS.n3838 0.00532143
R37220 DVSS.n4222 DVSS.n4215 0.00532143
R37221 DVSS.n4207 DVSS.n4201 0.00532143
R37222 DVSS.n4384 DVSS.n3721 0.00532143
R37223 DVSS.n8899 DVSS.n766 0.00528346
R37224 DVSS.n8997 DVSS.n722 0.00528346
R37225 DVSS.n9433 DVSS.n351 0.00528346
R37226 DVSS.n9530 DVSS.n25 0.00528346
R37227 DVSS.n4493 DVSS.n3834 0.00521831
R37228 DVSS.n4520 DVSS.n3815 0.00521831
R37229 DVSS.n4574 DVSS.n3801 0.00521831
R37230 DVSS.n4778 DVSS.n3729 0.00521831
R37231 DVSS.n1436 DVSS.n1425 0.00506429
R37232 DVSS.n1665 DVSS.n1425 0.00506429
R37233 DVSS.n1114 DVSS.n1105 0.00506429
R37234 DVSS.n1697 DVSS.n1105 0.00506429
R37235 DVSS.n1720 DVSS.n1713 0.00506429
R37236 DVSS.n1720 DVSS.n1719 0.00506429
R37237 DVSS.n1746 DVSS.n1571 0.00506429
R37238 DVSS.n1746 DVSS.n1745 0.00506429
R37239 DVSS.n7844 DVSS.n7737 0.00506429
R37240 DVSS.n7844 DVSS.n7843 0.00506429
R37241 DVSS.n1832 DVSS.n1822 0.00506429
R37242 DVSS.n1832 DVSS.n1831 0.00506429
R37243 DVSS.n8145 DVSS.n8138 0.00506429
R37244 DVSS.n8145 DVSS.n8144 0.00506429
R37245 DVSS.n1770 DVSS.n1762 0.00506429
R37246 DVSS.n8167 DVSS.n1762 0.00506429
R37247 DVSS.n5163 DVSS.n3327 0.00506429
R37248 DVSS.n5161 DVSS.n3327 0.00506429
R37249 DVSS.n5131 DVSS.n5130 0.00506429
R37250 DVSS.n5130 DVSS.n5068 0.00506429
R37251 DVSS.n5088 DVSS.n3373 0.00506429
R37252 DVSS.n5113 DVSS.n3373 0.00506429
R37253 DVSS.n2959 DVSS.n2949 0.00506429
R37254 DVSS.n5097 DVSS.n2959 0.00506429
R37255 DVSS.n5269 DVSS.n3440 0.00506429
R37256 DVSS.n5273 DVSS.n3440 0.00506429
R37257 DVSS.n5304 DVSS.n3405 0.00506429
R37258 DVSS.n5308 DVSS.n3405 0.00506429
R37259 DVSS.n3386 DVSS.n3378 0.00506429
R37260 DVSS.n5324 DVSS.n3378 0.00506429
R37261 DVSS.n2931 DVSS.n2922 0.00506429
R37262 DVSS.n5333 DVSS.n2922 0.00506429
R37263 DVSS.n3666 DVSS.n3660 0.00506429
R37264 DVSS.n3666 DVSS.n3665 0.00506429
R37265 DVSS.n4881 DVSS.n3625 0.00506429
R37266 DVSS.n3625 DVSS.n3624 0.00506429
R37267 DVSS.n4961 DVSS.n3598 0.00506429
R37268 DVSS.n3606 DVSS.n3598 0.00506429
R37269 DVSS.n4922 DVSS.n4912 0.00506429
R37270 DVSS.n4935 DVSS.n4922 0.00506429
R37271 DVSS.n1082 DVSS.n561 0.00493662
R37272 DVSS.n8522 DVSS.n589 0.00493662
R37273 DVSS.n367 DVSS.n268 0.00492913
R37274 DVSS.n421 DVSS.n369 0.00492913
R37275 DVSS.n8861 DVSS.n8860 0.00492913
R37276 DVSS.n6942 DVSS.n796 0.00492913
R37277 DVSS.n8938 DVSS.n752 0.00492913
R37278 DVSS.n8974 DVSS.n731 0.00492913
R37279 DVSS.n9472 DVSS.n337 0.00492913
R37280 DVSS.n9508 DVSS.n30 0.00492913
R37281 DVSS.n2932 DVSS.n2915 0.00492913
R37282 DVSS.n5855 DVSS.n3020 0.00492913
R37283 DVSS.n6762 DVSS.n6737 0.00480714
R37284 DVSS.n6834 DVSS.n6668 0.00480714
R37285 DVSS.n6780 DVSS.n1163 0.00480714
R37286 DVSS.n1345 DVSS.n1327 0.00480714
R37287 DVSS.n1934 DVSS.n1918 0.00480714
R37288 DVSS.n8037 DVSS.n1956 0.00480714
R37289 DVSS.n8014 DVSS.n1982 0.00480714
R37290 DVSS.n7975 DVSS.n2016 0.00480714
R37291 DVSS.n3080 DVSS.n2996 0.00480714
R37292 DVSS.n3118 DVSS.n3112 0.00480714
R37293 DVSS.n5777 DVSS.n3147 0.00480714
R37294 DVSS.n3035 DVSS.n3029 0.00480714
R37295 DVSS.n4166 DVSS.n3889 0.00480714
R37296 DVSS.n4137 DVSS.n4136 0.00480714
R37297 DVSS.n4238 DVSS.n3838 0.00480714
R37298 DVSS.n4261 DVSS.n4215 0.00480714
R37299 DVSS.n4412 DVSS.n4201 0.00480714
R37300 DVSS.n4287 DVSS.n3721 0.00480714
R37301 DVSS.n7382 DVSS.n2529 0.00476
R37302 DVSS.n7382 DVSS.n2527 0.00476
R37303 DVSS.n7386 DVSS.n2527 0.00476
R37304 DVSS.n7386 DVSS.n2525 0.00476
R37305 DVSS.n7390 DVSS.n2525 0.00476
R37306 DVSS.n7390 DVSS.n2523 0.00476
R37307 DVSS.n7394 DVSS.n2523 0.00476
R37308 DVSS.n7394 DVSS.n2472 0.00476
R37309 DVSS.n7401 DVSS.n2472 0.00476
R37310 DVSS.n7401 DVSS.n2470 0.00476
R37311 DVSS.n7405 DVSS.n2470 0.00476
R37312 DVSS.n7405 DVSS.n2468 0.00476
R37313 DVSS.n7409 DVSS.n2468 0.00476
R37314 DVSS.n7409 DVSS.n2466 0.00476
R37315 DVSS.n7413 DVSS.n2466 0.00476
R37316 DVSS.n7413 DVSS.n2416 0.00476
R37317 DVSS.n7421 DVSS.n2416 0.00476
R37318 DVSS.n7421 DVSS.n2414 0.00476
R37319 DVSS.n7425 DVSS.n2414 0.00476
R37320 DVSS.n7425 DVSS.n2412 0.00476
R37321 DVSS.n7429 DVSS.n2412 0.00476
R37322 DVSS.n7429 DVSS.n2410 0.00476
R37323 DVSS.n7433 DVSS.n2410 0.00476
R37324 DVSS.n7433 DVSS.n2408 0.00476
R37325 DVSS.n7437 DVSS.n2408 0.00476
R37326 DVSS.n7437 DVSS.n2406 0.00476
R37327 DVSS.n7441 DVSS.n2406 0.00476
R37328 DVSS.n7441 DVSS.n2404 0.00476
R37329 DVSS.n7445 DVSS.n2404 0.00476
R37330 DVSS.n7445 DVSS.n2402 0.00476
R37331 DVSS.n7449 DVSS.n2402 0.00476
R37332 DVSS.n7449 DVSS.n2351 0.00476
R37333 DVSS.n7456 DVSS.n2351 0.00476
R37334 DVSS.n7456 DVSS.n2349 0.00476
R37335 DVSS.n7460 DVSS.n2349 0.00476
R37336 DVSS.n7460 DVSS.n2347 0.00476
R37337 DVSS.n7464 DVSS.n2347 0.00476
R37338 DVSS.n7464 DVSS.n2345 0.00476
R37339 DVSS.n7468 DVSS.n2345 0.00476
R37340 DVSS.n7468 DVSS.n2343 0.00476
R37341 DVSS.n7472 DVSS.n2343 0.00476
R37342 DVSS.n7472 DVSS.n2341 0.00476
R37343 DVSS.n7476 DVSS.n2341 0.00476
R37344 DVSS.n7476 DVSS.n2339 0.00476
R37345 DVSS.n7480 DVSS.n2339 0.00476
R37346 DVSS.n7480 DVSS.n2337 0.00476
R37347 DVSS.n7484 DVSS.n2337 0.00476
R37348 DVSS.n7484 DVSS.n2309 0.00476
R37349 DVSS.n7491 DVSS.n2309 0.00476
R37350 DVSS.n7491 DVSS.n2307 0.00476
R37351 DVSS.n7495 DVSS.n2307 0.00476
R37352 DVSS.n7495 DVSS.n2279 0.00476
R37353 DVSS.n7502 DVSS.n2279 0.00476
R37354 DVSS.n7502 DVSS.n2277 0.00476
R37355 DVSS.n7506 DVSS.n2277 0.00476
R37356 DVSS.n7506 DVSS.n2275 0.00476
R37357 DVSS.n7510 DVSS.n2275 0.00476
R37358 DVSS.n7510 DVSS.n2273 0.00476
R37359 DVSS.n7514 DVSS.n2273 0.00476
R37360 DVSS.n7514 DVSS.n2271 0.00476
R37361 DVSS.n7518 DVSS.n2271 0.00476
R37362 DVSS.n7518 DVSS.n2269 0.00476
R37363 DVSS.n7522 DVSS.n2269 0.00476
R37364 DVSS.n7522 DVSS.n2267 0.00476
R37365 DVSS.n7526 DVSS.n2267 0.00476
R37366 DVSS.n7526 DVSS.n2265 0.00476
R37367 DVSS.n7530 DVSS.n2265 0.00476
R37368 DVSS.n7530 DVSS.n2237 0.00476
R37369 DVSS.n7560 DVSS.n2237 0.00476
R37370 DVSS.n7560 DVSS.n2235 0.00476
R37371 DVSS.n7564 DVSS.n2235 0.00476
R37372 DVSS.n7564 DVSS.n2233 0.00476
R37373 DVSS.n7568 DVSS.n2233 0.00476
R37374 DVSS.n7568 DVSS.n2231 0.00476
R37375 DVSS.n7572 DVSS.n2231 0.00476
R37376 DVSS.n7572 DVSS.n2229 0.00476
R37377 DVSS.n7576 DVSS.n2229 0.00476
R37378 DVSS.n7576 DVSS.n2227 0.00476
R37379 DVSS.n7580 DVSS.n2227 0.00476
R37380 DVSS.n7580 DVSS.n2225 0.00476
R37381 DVSS.n7584 DVSS.n2225 0.00476
R37382 DVSS.n7584 DVSS.n2223 0.00476
R37383 DVSS.n7588 DVSS.n2223 0.00476
R37384 DVSS.n7588 DVSS.n2195 0.00476
R37385 DVSS.n7618 DVSS.n2195 0.00476
R37386 DVSS.n7618 DVSS.n2193 0.00476
R37387 DVSS.n7622 DVSS.n2193 0.00476
R37388 DVSS.n7622 DVSS.n2191 0.00476
R37389 DVSS.n7626 DVSS.n2191 0.00476
R37390 DVSS.n7626 DVSS.n2189 0.00476
R37391 DVSS.n7630 DVSS.n2189 0.00476
R37392 DVSS.n7630 DVSS.n2161 0.00476
R37393 DVSS.n7660 DVSS.n2161 0.00476
R37394 DVSS.n7660 DVSS.n2159 0.00476
R37395 DVSS.n7665 DVSS.n2159 0.00476
R37396 DVSS.n7665 DVSS.n2156 0.00476
R37397 DVSS.n7669 DVSS.n2156 0.00476
R37398 DVSS.n7670 DVSS.n2155 0.00476
R37399 DVSS.n7677 DVSS.n2155 0.00476
R37400 DVSS.n7677 DVSS.n7676 0.00476
R37401 DVSS.n7388 DVSS.n7387 0.00476
R37402 DVSS.n7389 DVSS.n7388 0.00476
R37403 DVSS.n7389 DVSS.n2522 0.00476
R37404 DVSS.n7395 DVSS.n2522 0.00476
R37405 DVSS.n7407 DVSS.n7406 0.00476
R37406 DVSS.n7408 DVSS.n7407 0.00476
R37407 DVSS.n7408 DVSS.n2465 0.00476
R37408 DVSS.n7414 DVSS.n2465 0.00476
R37409 DVSS.n7427 DVSS.n7426 0.00476
R37410 DVSS.n7428 DVSS.n7427 0.00476
R37411 DVSS.n7428 DVSS.n2409 0.00476
R37412 DVSS.n7434 DVSS.n2409 0.00476
R37413 DVSS.n7435 DVSS.n7434 0.00476
R37414 DVSS.n7436 DVSS.n7435 0.00476
R37415 DVSS.n7436 DVSS.n2405 0.00476
R37416 DVSS.n7442 DVSS.n2405 0.00476
R37417 DVSS.n7443 DVSS.n7442 0.00476
R37418 DVSS.n7444 DVSS.n7443 0.00476
R37419 DVSS.n7444 DVSS.n2401 0.00476
R37420 DVSS.n7450 DVSS.n2401 0.00476
R37421 DVSS.n7462 DVSS.n7461 0.00476
R37422 DVSS.n7463 DVSS.n7462 0.00476
R37423 DVSS.n7463 DVSS.n2344 0.00476
R37424 DVSS.n7469 DVSS.n2344 0.00476
R37425 DVSS.n7470 DVSS.n7469 0.00476
R37426 DVSS.n7471 DVSS.n7470 0.00476
R37427 DVSS.n7471 DVSS.n2340 0.00476
R37428 DVSS.n7477 DVSS.n2340 0.00476
R37429 DVSS.n7478 DVSS.n7477 0.00476
R37430 DVSS.n7479 DVSS.n7478 0.00476
R37431 DVSS.n7479 DVSS.n2336 0.00476
R37432 DVSS.n7485 DVSS.n2336 0.00476
R37433 DVSS.n7496 DVSS.n2306 0.00476
R37434 DVSS.n7507 DVSS.n2276 0.00476
R37435 DVSS.n7508 DVSS.n7507 0.00476
R37436 DVSS.n7509 DVSS.n7508 0.00476
R37437 DVSS.n7509 DVSS.n2272 0.00476
R37438 DVSS.n7515 DVSS.n2272 0.00476
R37439 DVSS.n7516 DVSS.n7515 0.00476
R37440 DVSS.n7517 DVSS.n7516 0.00476
R37441 DVSS.n7517 DVSS.n2268 0.00476
R37442 DVSS.n7523 DVSS.n2268 0.00476
R37443 DVSS.n7524 DVSS.n7523 0.00476
R37444 DVSS.n7525 DVSS.n7524 0.00476
R37445 DVSS.n7525 DVSS.n2253 0.00476
R37446 DVSS.n7565 DVSS.n2234 0.00476
R37447 DVSS.n7566 DVSS.n7565 0.00476
R37448 DVSS.n7567 DVSS.n7566 0.00476
R37449 DVSS.n7567 DVSS.n2230 0.00476
R37450 DVSS.n7573 DVSS.n2230 0.00476
R37451 DVSS.n7574 DVSS.n7573 0.00476
R37452 DVSS.n7575 DVSS.n7574 0.00476
R37453 DVSS.n7575 DVSS.n2226 0.00476
R37454 DVSS.n7581 DVSS.n2226 0.00476
R37455 DVSS.n7582 DVSS.n7581 0.00476
R37456 DVSS.n7583 DVSS.n7582 0.00476
R37457 DVSS.n7583 DVSS.n2211 0.00476
R37458 DVSS.n7623 DVSS.n2192 0.00476
R37459 DVSS.n7624 DVSS.n7623 0.00476
R37460 DVSS.n7625 DVSS.n7624 0.00476
R37461 DVSS.n7625 DVSS.n2177 0.00476
R37462 DVSS.n7666 DVSS.n2158 0.00476
R37463 DVSS.n7667 DVSS.n7666 0.00476
R37464 DVSS.n7668 DVSS.n7667 0.00476
R37465 DVSS.n6921 DVSS.n6730 0.00476
R37466 DVSS.n6922 DVSS.n6921 0.00476
R37467 DVSS.n6923 DVSS.n6922 0.00476
R37468 DVSS.n6923 DVSS.n6693 0.00476
R37469 DVSS.n6930 DVSS.n6929 0.00476
R37470 DVSS.n7035 DVSS.n6930 0.00476
R37471 DVSS.n7035 DVSS.n7034 0.00476
R37472 DVSS.n1042 DVSS.n1039 0.00476
R37473 DVSS.n1043 DVSS.n1042 0.00476
R37474 DVSS.n1044 DVSS.n1043 0.00476
R37475 DVSS.n1045 DVSS.n1044 0.00476
R37476 DVSS.n1048 DVSS.n1045 0.00476
R37477 DVSS.n1049 DVSS.n1048 0.00476
R37478 DVSS.n1050 DVSS.n1049 0.00476
R37479 DVSS.n1051 DVSS.n1050 0.00476
R37480 DVSS.n1054 DVSS.n1051 0.00476
R37481 DVSS.n1055 DVSS.n1054 0.00476
R37482 DVSS.n1056 DVSS.n1055 0.00476
R37483 DVSS.n1057 DVSS.n1056 0.00476
R37484 DVSS.n8564 DVSS.n8562 0.00476
R37485 DVSS.n8564 DVSS.n8563 0.00476
R37486 DVSS.n8563 DVSS.n629 0.00476
R37487 DVSS.n9095 DVSS.n624 0.00476
R37488 DVSS.n9096 DVSS.n9095 0.00476
R37489 DVSS.n9097 DVSS.n9096 0.00476
R37490 DVSS.n9097 DVSS.n620 0.00476
R37491 DVSS.n9103 DVSS.n620 0.00476
R37492 DVSS.n9104 DVSS.n9103 0.00476
R37493 DVSS.n9105 DVSS.n9104 0.00476
R37494 DVSS.n9105 DVSS.n607 0.00476
R37495 DVSS.n9131 DVSS.n575 0.00476
R37496 DVSS.n9161 DVSS.n9160 0.00476
R37497 DVSS.n9161 DVSS.n555 0.00476
R37498 DVSS.n9167 DVSS.n555 0.00476
R37499 DVSS.n9168 DVSS.n9167 0.00476
R37500 DVSS.n9170 DVSS.n9168 0.00476
R37501 DVSS.n9170 DVSS.n9169 0.00476
R37502 DVSS.n9169 DVSS.n551 0.00476
R37503 DVSS.n9178 DVSS.n551 0.00476
R37504 DVSS.n9626 DVSS.n231 0.00476
R37505 DVSS.n9627 DVSS.n9626 0.00476
R37506 DVSS.n9628 DVSS.n9627 0.00476
R37507 DVSS.n9661 DVSS.n200 0.00476
R37508 DVSS.n9667 DVSS.n200 0.00476
R37509 DVSS.n9668 DVSS.n9667 0.00476
R37510 DVSS.n9669 DVSS.n9668 0.00476
R37511 DVSS.n9669 DVSS.n196 0.00476
R37512 DVSS.n9675 DVSS.n196 0.00476
R37513 DVSS.n9676 DVSS.n9675 0.00476
R37514 DVSS.n9677 DVSS.n9676 0.00476
R37515 DVSS.n9677 DVSS.n192 0.00476
R37516 DVSS.n9683 DVSS.n192 0.00476
R37517 DVSS.n9684 DVSS.n9683 0.00476
R37518 DVSS.n9685 DVSS.n9684 0.00476
R37519 DVSS.n9725 DVSS.n9724 0.00476
R37520 DVSS.n9727 DVSS.n9725 0.00476
R37521 DVSS.n9727 DVSS.n9726 0.00476
R37522 DVSS.n9778 DVSS.n139 0.00476
R37523 DVSS.n9779 DVSS.n9778 0.00476
R37524 DVSS.n9780 DVSS.n9779 0.00476
R37525 DVSS.n1018 DVSS.n1017 0.00476
R37526 DVSS.n1019 DVSS.n1018 0.00476
R37527 DVSS.n1020 DVSS.n1019 0.00476
R37528 DVSS.n1020 DVSS.n758 0.00476
R37529 DVSS.n1028 DVSS.n1027 0.00476
R37530 DVSS.n1029 DVSS.n1028 0.00476
R37531 DVSS.n1030 DVSS.n1029 0.00476
R37532 DVSS.n6988 DVSS.n6987 0.00476
R37533 DVSS.n6989 DVSS.n6988 0.00476
R37534 DVSS.n6990 DVSS.n6989 0.00476
R37535 DVSS.n6993 DVSS.n6990 0.00476
R37536 DVSS.n6994 DVSS.n6993 0.00476
R37537 DVSS.n6995 DVSS.n6994 0.00476
R37538 DVSS.n6996 DVSS.n6995 0.00476
R37539 DVSS.n6999 DVSS.n6996 0.00476
R37540 DVSS.n7000 DVSS.n6999 0.00476
R37541 DVSS.n7001 DVSS.n7000 0.00476
R37542 DVSS.n7002 DVSS.n7001 0.00476
R37543 DVSS.n7003 DVSS.n7002 0.00476
R37544 DVSS.n829 DVSS.n810 0.00476
R37545 DVSS.n8815 DVSS.n829 0.00476
R37546 DVSS.n8815 DVSS.n8814 0.00476
R37547 DVSS.n635 DVSS.n632 0.00476
R37548 DVSS.n636 DVSS.n635 0.00476
R37549 DVSS.n637 DVSS.n636 0.00476
R37550 DVSS.n638 DVSS.n637 0.00476
R37551 DVSS.n641 DVSS.n638 0.00476
R37552 DVSS.n642 DVSS.n641 0.00476
R37553 DVSS.n643 DVSS.n642 0.00476
R37554 DVSS.n644 DVSS.n643 0.00476
R37555 DVSS.n9066 DVSS.n503 0.00476
R37556 DVSS.n542 DVSS.n541 0.00476
R37557 DVSS.n543 DVSS.n542 0.00476
R37558 DVSS.n544 DVSS.n543 0.00476
R37559 DVSS.n547 DVSS.n544 0.00476
R37560 DVSS.n548 DVSS.n547 0.00476
R37561 DVSS.n549 DVSS.n548 0.00476
R37562 DVSS.n550 DVSS.n549 0.00476
R37563 DVSS.n9181 DVSS.n550 0.00476
R37564 DVSS.n239 DVSS.n238 0.00476
R37565 DVSS.n240 DVSS.n239 0.00476
R37566 DVSS.n409 DVSS.n240 0.00476
R37567 DVSS.n443 DVSS.n248 0.00476
R37568 DVSS.n249 DVSS.n248 0.00476
R37569 DVSS.n250 DVSS.n249 0.00476
R37570 DVSS.n253 DVSS.n250 0.00476
R37571 DVSS.n254 DVSS.n253 0.00476
R37572 DVSS.n255 DVSS.n254 0.00476
R37573 DVSS.n256 DVSS.n255 0.00476
R37574 DVSS.n259 DVSS.n256 0.00476
R37575 DVSS.n260 DVSS.n259 0.00476
R37576 DVSS.n261 DVSS.n260 0.00476
R37577 DVSS.n262 DVSS.n261 0.00476
R37578 DVSS.n9548 DVSS.n262 0.00476
R37579 DVSS.n68 DVSS.n65 0.00476
R37580 DVSS.n69 DVSS.n68 0.00476
R37581 DVSS.n70 DVSS.n69 0.00476
R37582 DVSS.n76 DVSS.n75 0.00476
R37583 DVSS.n79 DVSS.n76 0.00476
R37584 DVSS.n80 DVSS.n79 0.00476
R37585 DVSS.n81 DVSS.n80 0.00476
R37586 DVSS.n8689 DVSS.n960 0.00476
R37587 DVSS.n8690 DVSS.n8689 0.00476
R37588 DVSS.n8692 DVSS.n8690 0.00476
R37589 DVSS.n8692 DVSS.n8691 0.00476
R37590 DVSS.n8705 DVSS.n738 0.00476
R37591 DVSS.n8706 DVSS.n8705 0.00476
R37592 DVSS.n8707 DVSS.n8706 0.00476
R37593 DVSS.n8725 DVSS.n8724 0.00476
R37594 DVSS.n8726 DVSS.n8725 0.00476
R37595 DVSS.n8726 DVSS.n894 0.00476
R37596 DVSS.n8732 DVSS.n894 0.00476
R37597 DVSS.n8733 DVSS.n8732 0.00476
R37598 DVSS.n8734 DVSS.n8733 0.00476
R37599 DVSS.n8734 DVSS.n890 0.00476
R37600 DVSS.n8740 DVSS.n890 0.00476
R37601 DVSS.n8741 DVSS.n8740 0.00476
R37602 DVSS.n8742 DVSS.n8741 0.00476
R37603 DVSS.n8742 DVSS.n886 0.00476
R37604 DVSS.n8748 DVSS.n886 0.00476
R37605 DVSS.n8761 DVSS.n8760 0.00476
R37606 DVSS.n8762 DVSS.n8761 0.00476
R37607 DVSS.n8762 DVSS.n830 0.00476
R37608 DVSS.n8810 DVSS.n831 0.00476
R37609 DVSS.n8768 DVSS.n831 0.00476
R37610 DVSS.n8769 DVSS.n8768 0.00476
R37611 DVSS.n8770 DVSS.n8769 0.00476
R37612 DVSS.n8773 DVSS.n8770 0.00476
R37613 DVSS.n8774 DVSS.n8773 0.00476
R37614 DVSS.n8775 DVSS.n8774 0.00476
R37615 DVSS.n8775 DVSS.n663 0.00476
R37616 DVSS.n8791 DVSS.n8790 0.00476
R37617 DVSS.n9268 DVSS.n9267 0.00476
R37618 DVSS.n9269 DVSS.n9268 0.00476
R37619 DVSS.n9269 DVSS.n491 0.00476
R37620 DVSS.n9275 DVSS.n491 0.00476
R37621 DVSS.n9276 DVSS.n9275 0.00476
R37622 DVSS.n9278 DVSS.n9276 0.00476
R37623 DVSS.n9278 DVSS.n9277 0.00476
R37624 DVSS.n9277 DVSS.n488 0.00476
R37625 DVSS.n9289 DVSS.n9288 0.00476
R37626 DVSS.n9290 DVSS.n9289 0.00476
R37627 DVSS.n9290 DVSS.n394 0.00476
R37628 DVSS.n9297 DVSS.n9296 0.00476
R37629 DVSS.n9298 DVSS.n9297 0.00476
R37630 DVSS.n9301 DVSS.n9298 0.00476
R37631 DVSS.n9302 DVSS.n9301 0.00476
R37632 DVSS.n9303 DVSS.n9302 0.00476
R37633 DVSS.n9304 DVSS.n9303 0.00476
R37634 DVSS.n9307 DVSS.n9304 0.00476
R37635 DVSS.n9308 DVSS.n9307 0.00476
R37636 DVSS.n9309 DVSS.n9308 0.00476
R37637 DVSS.n9310 DVSS.n9309 0.00476
R37638 DVSS.n9311 DVSS.n9310 0.00476
R37639 DVSS.n9311 DVSS.n288 0.00476
R37640 DVSS.n9876 DVSS.n57 0.00476
R37641 DVSS.n9877 DVSS.n9876 0.00476
R37642 DVSS.n9878 DVSS.n9877 0.00476
R37643 DVSS.n9890 DVSS.n9889 0.00476
R37644 DVSS.n9890 DVSS.n20 0.00476
R37645 DVSS.n9896 DVSS.n20 0.00476
R37646 DVSS.n8654 DVSS.n963 0.00476
R37647 DVSS.n8684 DVSS.n963 0.00476
R37648 DVSS.n8684 DVSS.n961 0.00476
R37649 DVSS.n8688 DVSS.n961 0.00476
R37650 DVSS.n8688 DVSS.n959 0.00476
R37651 DVSS.n8693 DVSS.n959 0.00476
R37652 DVSS.n8693 DVSS.n956 0.00476
R37653 DVSS.n8697 DVSS.n956 0.00476
R37654 DVSS.n8699 DVSS.n8697 0.00476
R37655 DVSS.n8700 DVSS.n8699 0.00476
R37656 DVSS.n8700 DVSS.n954 0.00476
R37657 DVSS.n8704 DVSS.n954 0.00476
R37658 DVSS.n8704 DVSS.n953 0.00476
R37659 DVSS.n8708 DVSS.n953 0.00476
R37660 DVSS.n8712 DVSS.n901 0.00476
R37661 DVSS.n8719 DVSS.n901 0.00476
R37662 DVSS.n8719 DVSS.n899 0.00476
R37663 DVSS.n8723 DVSS.n899 0.00476
R37664 DVSS.n8723 DVSS.n897 0.00476
R37665 DVSS.n8727 DVSS.n897 0.00476
R37666 DVSS.n8727 DVSS.n895 0.00476
R37667 DVSS.n8731 DVSS.n895 0.00476
R37668 DVSS.n8731 DVSS.n893 0.00476
R37669 DVSS.n8735 DVSS.n893 0.00476
R37670 DVSS.n8735 DVSS.n891 0.00476
R37671 DVSS.n8739 DVSS.n891 0.00476
R37672 DVSS.n8739 DVSS.n889 0.00476
R37673 DVSS.n8743 DVSS.n889 0.00476
R37674 DVSS.n8743 DVSS.n887 0.00476
R37675 DVSS.n8747 DVSS.n887 0.00476
R37676 DVSS.n8747 DVSS.n838 0.00476
R37677 DVSS.n8754 DVSS.n838 0.00476
R37678 DVSS.n8754 DVSS.n836 0.00476
R37679 DVSS.n8759 DVSS.n836 0.00476
R37680 DVSS.n8759 DVSS.n834 0.00476
R37681 DVSS.n8763 DVSS.n834 0.00476
R37682 DVSS.n8764 DVSS.n8763 0.00476
R37683 DVSS.n8809 DVSS.n832 0.00476
R37684 DVSS.n8805 DVSS.n832 0.00476
R37685 DVSS.n8805 DVSS.n8804 0.00476
R37686 DVSS.n8804 DVSS.n8803 0.00476
R37687 DVSS.n8803 DVSS.n8771 0.00476
R37688 DVSS.n8799 DVSS.n8771 0.00476
R37689 DVSS.n8799 DVSS.n8798 0.00476
R37690 DVSS.n8798 DVSS.n8797 0.00476
R37691 DVSS.n8797 DVSS.n8776 0.00476
R37692 DVSS.n8793 DVSS.n8776 0.00476
R37693 DVSS.n8793 DVSS.n8792 0.00476
R37694 DVSS.n8792 DVSS.n498 0.00476
R37695 DVSS.n9262 DVSS.n498 0.00476
R37696 DVSS.n9262 DVSS.n496 0.00476
R37697 DVSS.n9266 DVSS.n496 0.00476
R37698 DVSS.n9266 DVSS.n494 0.00476
R37699 DVSS.n9270 DVSS.n494 0.00476
R37700 DVSS.n9270 DVSS.n492 0.00476
R37701 DVSS.n9274 DVSS.n492 0.00476
R37702 DVSS.n9274 DVSS.n490 0.00476
R37703 DVSS.n9279 DVSS.n490 0.00476
R37704 DVSS.n9279 DVSS.n487 0.00476
R37705 DVSS.n9283 DVSS.n487 0.00476
R37706 DVSS.n9287 DVSS.n485 0.00476
R37707 DVSS.n9291 DVSS.n485 0.00476
R37708 DVSS.n9292 DVSS.n9291 0.00476
R37709 DVSS.n9292 DVSS.n481 0.00476
R37710 DVSS.n9351 DVSS.n481 0.00476
R37711 DVSS.n9351 DVSS.n483 0.00476
R37712 DVSS.n9347 DVSS.n483 0.00476
R37713 DVSS.n9347 DVSS.n9346 0.00476
R37714 DVSS.n9346 DVSS.n9345 0.00476
R37715 DVSS.n9345 DVSS.n9299 0.00476
R37716 DVSS.n9341 DVSS.n9299 0.00476
R37717 DVSS.n9341 DVSS.n9340 0.00476
R37718 DVSS.n9340 DVSS.n9339 0.00476
R37719 DVSS.n9339 DVSS.n9305 0.00476
R37720 DVSS.n9335 DVSS.n9305 0.00476
R37721 DVSS.n9335 DVSS.n9334 0.00476
R37722 DVSS.n9334 DVSS.n9333 0.00476
R37723 DVSS.n9333 DVSS.n9312 0.00476
R37724 DVSS.n9329 DVSS.n9312 0.00476
R37725 DVSS.n9329 DVSS.n9328 0.00476
R37726 DVSS.n9328 DVSS.n9327 0.00476
R37727 DVSS.n9327 DVSS.n61 0.00476
R37728 DVSS.n9870 DVSS.n61 0.00476
R37729 DVSS.n9875 DVSS.n58 0.00476
R37730 DVSS.n9875 DVSS.n56 0.00476
R37731 DVSS.n9879 DVSS.n56 0.00476
R37732 DVSS.n9879 DVSS.n53 0.00476
R37733 DVSS.n9884 DVSS.n53 0.00476
R37734 DVSS.n9884 DVSS.n54 0.00476
R37735 DVSS.n54 DVSS.n23 0.00476
R37736 DVSS.n9891 DVSS.n23 0.00476
R37737 DVSS.n9891 DVSS.n21 0.00476
R37738 DVSS.n9895 DVSS.n21 0.00476
R37739 DVSS.n9938 DVSS.n2 0.00476
R37740 DVSS.n9938 DVSS.n9937 0.00476
R37741 DVSS.n9937 DVSS.n9936 0.00476
R37742 DVSS.n8622 DVSS.n1013 0.00476
R37743 DVSS.n8622 DVSS.n1015 0.00476
R37744 DVSS.n8618 DVSS.n1015 0.00476
R37745 DVSS.n8618 DVSS.n8617 0.00476
R37746 DVSS.n8617 DVSS.n8616 0.00476
R37747 DVSS.n8616 DVSS.n1021 0.00476
R37748 DVSS.n8612 DVSS.n1021 0.00476
R37749 DVSS.n8612 DVSS.n8611 0.00476
R37750 DVSS.n8611 DVSS.n8610 0.00476
R37751 DVSS.n8610 DVSS.n1025 0.00476
R37752 DVSS.n8606 DVSS.n1025 0.00476
R37753 DVSS.n8606 DVSS.n8605 0.00476
R37754 DVSS.n8605 DVSS.n8604 0.00476
R37755 DVSS.n8604 DVSS.n8601 0.00476
R37756 DVSS.n6983 DVSS.n1031 0.00476
R37757 DVSS.n6983 DVSS.n6980 0.00476
R37758 DVSS.n7025 DVSS.n6980 0.00476
R37759 DVSS.n7025 DVSS.n6981 0.00476
R37760 DVSS.n7021 DVSS.n6981 0.00476
R37761 DVSS.n7021 DVSS.n7020 0.00476
R37762 DVSS.n7020 DVSS.n7019 0.00476
R37763 DVSS.n7019 DVSS.n6991 0.00476
R37764 DVSS.n7015 DVSS.n6991 0.00476
R37765 DVSS.n7015 DVSS.n7014 0.00476
R37766 DVSS.n7014 DVSS.n7013 0.00476
R37767 DVSS.n7013 DVSS.n6997 0.00476
R37768 DVSS.n7009 DVSS.n6997 0.00476
R37769 DVSS.n7009 DVSS.n7008 0.00476
R37770 DVSS.n7008 DVSS.n7007 0.00476
R37771 DVSS.n7007 DVSS.n7004 0.00476
R37772 DVSS.n7004 DVSS.n825 0.00476
R37773 DVSS.n8824 DVSS.n825 0.00476
R37774 DVSS.n8824 DVSS.n826 0.00476
R37775 DVSS.n8820 DVSS.n826 0.00476
R37776 DVSS.n8820 DVSS.n8819 0.00476
R37777 DVSS.n8819 DVSS.n8818 0.00476
R37778 DVSS.n8818 DVSS.n631 0.00476
R37779 DVSS.n9086 DVSS.n633 0.00476
R37780 DVSS.n9082 DVSS.n633 0.00476
R37781 DVSS.n9082 DVSS.n9081 0.00476
R37782 DVSS.n9081 DVSS.n9080 0.00476
R37783 DVSS.n9080 DVSS.n639 0.00476
R37784 DVSS.n9076 DVSS.n639 0.00476
R37785 DVSS.n9076 DVSS.n9075 0.00476
R37786 DVSS.n9075 DVSS.n9074 0.00476
R37787 DVSS.n9074 DVSS.n645 0.00476
R37788 DVSS.n9070 DVSS.n645 0.00476
R37789 DVSS.n9070 DVSS.n9069 0.00476
R37790 DVSS.n9069 DVSS.n9068 0.00476
R37791 DVSS.n9068 DVSS.n537 0.00476
R37792 DVSS.n9196 DVSS.n537 0.00476
R37793 DVSS.n9196 DVSS.n538 0.00476
R37794 DVSS.n9192 DVSS.n538 0.00476
R37795 DVSS.n9192 DVSS.n9191 0.00476
R37796 DVSS.n9191 DVSS.n9190 0.00476
R37797 DVSS.n9190 DVSS.n545 0.00476
R37798 DVSS.n9186 DVSS.n545 0.00476
R37799 DVSS.n9186 DVSS.n9185 0.00476
R37800 DVSS.n9185 DVSS.n9184 0.00476
R37801 DVSS.n9184 DVSS.n9182 0.00476
R37802 DVSS.n9619 DVSS.n9618 0.00476
R37803 DVSS.n9618 DVSS.n9617 0.00476
R37804 DVSS.n9617 DVSS.n241 0.00476
R37805 DVSS.n9613 DVSS.n241 0.00476
R37806 DVSS.n9613 DVSS.n9612 0.00476
R37807 DVSS.n9612 DVSS.n9611 0.00476
R37808 DVSS.n9611 DVSS.n246 0.00476
R37809 DVSS.n9607 DVSS.n246 0.00476
R37810 DVSS.n9607 DVSS.n9606 0.00476
R37811 DVSS.n9606 DVSS.n9605 0.00476
R37812 DVSS.n9605 DVSS.n251 0.00476
R37813 DVSS.n9601 DVSS.n251 0.00476
R37814 DVSS.n9601 DVSS.n9600 0.00476
R37815 DVSS.n9600 DVSS.n9599 0.00476
R37816 DVSS.n9599 DVSS.n257 0.00476
R37817 DVSS.n9595 DVSS.n257 0.00476
R37818 DVSS.n9595 DVSS.n9594 0.00476
R37819 DVSS.n9594 DVSS.n9593 0.00476
R37820 DVSS.n9593 DVSS.n263 0.00476
R37821 DVSS.n9589 DVSS.n263 0.00476
R37822 DVSS.n9589 DVSS.n9588 0.00476
R37823 DVSS.n9588 DVSS.n9587 0.00476
R37824 DVSS.n9587 DVSS.n64 0.00476
R37825 DVSS.n9867 DVSS.n66 0.00476
R37826 DVSS.n9863 DVSS.n66 0.00476
R37827 DVSS.n9863 DVSS.n9862 0.00476
R37828 DVSS.n9862 DVSS.n9861 0.00476
R37829 DVSS.n9861 DVSS.n72 0.00476
R37830 DVSS.n9857 DVSS.n72 0.00476
R37831 DVSS.n9857 DVSS.n9856 0.00476
R37832 DVSS.n9856 DVSS.n9855 0.00476
R37833 DVSS.n9855 DVSS.n77 0.00476
R37834 DVSS.n9851 DVSS.n77 0.00476
R37835 DVSS.n9851 DVSS.n9850 0.00476
R37836 DVSS.n9849 DVSS.n83 0.00476
R37837 DVSS.n9845 DVSS.n83 0.00476
R37838 DVSS.n6885 DVSS.n6733 0.00476
R37839 DVSS.n6915 DVSS.n6733 0.00476
R37840 DVSS.n6915 DVSS.n6731 0.00476
R37841 DVSS.n6920 DVSS.n6731 0.00476
R37842 DVSS.n6920 DVSS.n6729 0.00476
R37843 DVSS.n6924 DVSS.n6729 0.00476
R37844 DVSS.n6925 DVSS.n6924 0.00476
R37845 DVSS.n6925 DVSS.n6725 0.00476
R37846 DVSS.n7044 DVSS.n6725 0.00476
R37847 DVSS.n7044 DVSS.n6727 0.00476
R37848 DVSS.n7040 DVSS.n6727 0.00476
R37849 DVSS.n7040 DVSS.n7039 0.00476
R37850 DVSS.n7039 DVSS.n7038 0.00476
R37851 DVSS.n7038 DVSS.n1032 0.00476
R37852 DVSS.n8598 DVSS.n1034 0.00476
R37853 DVSS.n8594 DVSS.n1034 0.00476
R37854 DVSS.n8594 DVSS.n8593 0.00476
R37855 DVSS.n8593 DVSS.n8592 0.00476
R37856 DVSS.n8592 DVSS.n1040 0.00476
R37857 DVSS.n8588 DVSS.n1040 0.00476
R37858 DVSS.n8588 DVSS.n8587 0.00476
R37859 DVSS.n8587 DVSS.n8586 0.00476
R37860 DVSS.n8586 DVSS.n1046 0.00476
R37861 DVSS.n8582 DVSS.n1046 0.00476
R37862 DVSS.n8582 DVSS.n8581 0.00476
R37863 DVSS.n8581 DVSS.n8580 0.00476
R37864 DVSS.n8580 DVSS.n1052 0.00476
R37865 DVSS.n8576 DVSS.n1052 0.00476
R37866 DVSS.n8576 DVSS.n8575 0.00476
R37867 DVSS.n8575 DVSS.n8574 0.00476
R37868 DVSS.n8574 DVSS.n1058 0.00476
R37869 DVSS.n8570 DVSS.n1058 0.00476
R37870 DVSS.n8570 DVSS.n8569 0.00476
R37871 DVSS.n8569 DVSS.n8568 0.00476
R37872 DVSS.n8568 DVSS.n8565 0.00476
R37873 DVSS.n8565 DVSS.n628 0.00476
R37874 DVSS.n9089 DVSS.n628 0.00476
R37875 DVSS.n9094 DVSS.n625 0.00476
R37876 DVSS.n9094 DVSS.n623 0.00476
R37877 DVSS.n9098 DVSS.n623 0.00476
R37878 DVSS.n9098 DVSS.n621 0.00476
R37879 DVSS.n9102 DVSS.n621 0.00476
R37880 DVSS.n9102 DVSS.n619 0.00476
R37881 DVSS.n9106 DVSS.n619 0.00476
R37882 DVSS.n9106 DVSS.n617 0.00476
R37883 DVSS.n9110 DVSS.n617 0.00476
R37884 DVSS.n9110 DVSS.n586 0.00476
R37885 DVSS.n9132 DVSS.n586 0.00476
R37886 DVSS.n9132 DVSS.n583 0.00476
R37887 DVSS.n9137 DVSS.n583 0.00476
R37888 DVSS.n9137 DVSS.n584 0.00476
R37889 DVSS.n584 DVSS.n558 0.00476
R37890 DVSS.n9162 DVSS.n558 0.00476
R37891 DVSS.n9162 DVSS.n556 0.00476
R37892 DVSS.n9166 DVSS.n556 0.00476
R37893 DVSS.n9166 DVSS.n554 0.00476
R37894 DVSS.n9171 DVSS.n554 0.00476
R37895 DVSS.n9171 DVSS.n552 0.00476
R37896 DVSS.n9175 DVSS.n552 0.00476
R37897 DVSS.n9177 DVSS.n9175 0.00476
R37898 DVSS.n9625 DVSS.n232 0.00476
R37899 DVSS.n9625 DVSS.n230 0.00476
R37900 DVSS.n9629 DVSS.n230 0.00476
R37901 DVSS.n9629 DVSS.n228 0.00476
R37902 DVSS.n9633 DVSS.n228 0.00476
R37903 DVSS.n9633 DVSS.n203 0.00476
R37904 DVSS.n9662 DVSS.n203 0.00476
R37905 DVSS.n9662 DVSS.n201 0.00476
R37906 DVSS.n9666 DVSS.n201 0.00476
R37907 DVSS.n9666 DVSS.n199 0.00476
R37908 DVSS.n9670 DVSS.n199 0.00476
R37909 DVSS.n9670 DVSS.n197 0.00476
R37910 DVSS.n9674 DVSS.n197 0.00476
R37911 DVSS.n9674 DVSS.n195 0.00476
R37912 DVSS.n9678 DVSS.n195 0.00476
R37913 DVSS.n9678 DVSS.n193 0.00476
R37914 DVSS.n9682 DVSS.n193 0.00476
R37915 DVSS.n9682 DVSS.n191 0.00476
R37916 DVSS.n9686 DVSS.n191 0.00476
R37917 DVSS.n9686 DVSS.n189 0.00476
R37918 DVSS.n9690 DVSS.n189 0.00476
R37919 DVSS.n9690 DVSS.n164 0.00476
R37920 DVSS.n9719 DVSS.n164 0.00476
R37921 DVSS.n9723 DVSS.n161 0.00476
R37922 DVSS.n9728 DVSS.n161 0.00476
R37923 DVSS.n9728 DVSS.n159 0.00476
R37924 DVSS.n9732 DVSS.n159 0.00476
R37925 DVSS.n9732 DVSS.n142 0.00476
R37926 DVSS.n9772 DVSS.n142 0.00476
R37927 DVSS.n9772 DVSS.n140 0.00476
R37928 DVSS.n9777 DVSS.n140 0.00476
R37929 DVSS.n9777 DVSS.n138 0.00476
R37930 DVSS.n9781 DVSS.n138 0.00476
R37931 DVSS.n9782 DVSS.n134 0.00476
R37932 DVSS.n9787 DVSS.n134 0.00476
R37933 DVSS.n9787 DVSS.n136 0.00476
R37934 DVSS.n4627 DVSS.n4624 0.00472535
R37935 DVSS.n4695 DVSS.n3778 0.00472535
R37936 DVSS DVSS.n9896 0.00458
R37937 DVSS.n9895 DVSS 0.00458
R37938 DVSS.n8980 DVSS.n746 0.0045748
R37939 DVSS.n9514 DVSS.n44 0.0045748
R37940 DVSS.n5829 DVSS.n3062 0.00455
R37941 DVSS.n5834 DVSS.n3048 0.00455
R37942 DVSS.n5566 DVSS.n2299 0.00451408
R37943 DVSS.n5594 DVSS.n2329 0.00451408
R37944 DVSS.n4493 DVSS.n4492 0.00451408
R37945 DVSS.n4520 DVSS.n4519 0.00451408
R37946 DVSS.n4574 DVSS.n3800 0.00451408
R37947 DVSS.n4778 DVSS.n3728 0.00451408
R37948 DVSS.n8710 DVSS.n951 0.0045
R37949 DVSS.n8766 DVSS.n626 0.0045
R37950 DVSS.n9721 DVSS.n59 0.0045
R37951 DVSS.n9091 DVSS.n626 0.0045
R37952 DVSS.n1035 DVSS.n951 0.0045
R37953 DVSS.n9622 DVSS.n9621 0.0045
R37954 DVSS.n9621 DVSS.n234 0.0045
R37955 DVSS.n9872 DVSS.n59 0.0045
R37956 DVSS.n7487 DVSS.n7485 0.00446
R37957 DVSS.n9128 DVSS.n607 0.00446
R37958 DVSS.n9063 DVSS.n644 0.00446
R37959 DVSS.n9026 DVSS.n663 0.00446
R37960 DVSS.n5831 DVSS.n3062 0.00442143
R37961 DVSS.n5837 DVSS.n3048 0.00442143
R37962 DVSS.n7500 DVSS.n2276 0.00434
R37963 DVSS.n9160 DVSS.n9159 0.00434
R37964 DVSS.n541 DVSS.n502 0.00434
R37965 DVSS.n9267 DVSS.n495 0.00434
R37966 DVSS.n8391 DVSS.n1405 0.00430282
R37967 DVSS.n8358 DVSS.n1370 0.00430282
R37968 DVSS.n6003 DVSS.n2789 0.00423239
R37969 DVSS.n5999 DVSS.n2782 0.00423239
R37970 DVSS.n5975 DVSS.n2822 0.00423239
R37971 DVSS.n5972 DVSS.n2833 0.00423239
R37972 DVSS.n5960 DVSS.n2853 0.00423239
R37973 DVSS.n5955 DVSS.n2865 0.00423239
R37974 DVSS.n5943 DVSS.n2882 0.00423239
R37975 DVSS.n5940 DVSS.n5930 0.00423239
R37976 DVSS.n8504 DVSS.n188 0.00422047
R37977 DVSS.n8510 DVSS.n227 0.00422047
R37978 DVSS.n8538 DVSS.n1076 0.00422047
R37979 DVSS.n1214 DVSS.n1196 0.00422047
R37980 DVSS.n8893 DVSS.n772 0.00422047
R37981 DVSS.n8990 DVSS.n748 0.00422047
R37982 DVSS.n9427 DVSS.n356 0.00422047
R37983 DVSS.n9524 DVSS.n46 0.00422047
R37984 DVSS.n5377 DVSS.n2954 0.00422047
R37985 DVSS.n5875 DVSS.n3012 0.00422047
R37986 DVSS.n6854 DVSS.n6762 0.00416429
R37987 DVSS.n6834 DVSS.n6667 0.00416429
R37988 DVSS.n6780 DVSS.n1162 0.00416429
R37989 DVSS.n1345 DVSS.n1326 0.00416429
R37990 DVSS.n8056 DVSS.n1934 0.00416429
R37991 DVSS.n8034 DVSS.n1956 0.00416429
R37992 DVSS.n8011 DVSS.n1982 0.00416429
R37993 DVSS.n7972 DVSS.n2016 0.00416429
R37994 DVSS.n3080 DVSS.n2995 0.00416429
R37995 DVSS.n5811 DVSS.n3118 0.00416429
R37996 DVSS.n5775 DVSS.n3147 0.00416429
R37997 DVSS.n3035 DVSS.n3028 0.00416429
R37998 DVSS.n4166 DVSS.n3888 0.00416429
R37999 DVSS.n4136 DVSS.n3950 0.00416429
R38000 DVSS.n4238 DVSS.n3837 0.00416429
R38001 DVSS.n4261 DVSS.n4260 0.00416429
R38002 DVSS.n4412 DVSS.n4200 0.00416429
R38003 DVSS.n4287 DVSS.n3720 0.00416429
R38004 DVSS.n5556 DVSS.n2290 0.00409155
R38005 DVSS.n7888 DVSS.n2072 0.00409155
R38006 DVSS.n5615 DVSS.n2320 0.00409155
R38007 DVSS.n7889 DVSS.n2054 0.00409155
R38008 DVSS.n9724 DVSS.n162 0.00404
R38009 DVSS.n270 DVSS.n65 0.00404
R38010 DVSS.n269 DVSS.n57 0.00404
R38011 DVSS.n9869 DVSS.n58 0.00404
R38012 DVSS.n9868 DVSS.n9867 0.00404
R38013 DVSS.n9723 DVSS.n63 0.00404
R38014 DVSS.n6068 DVSS.n6033 0.00403571
R38015 DVSS.n6617 DVSS.n6347 0.00403571
R38016 DVSS.n4616 DVSS.n4608 0.00402113
R38017 DVSS.n4490 DVSS.n4489 0.0039507
R38018 DVSS.n4517 DVSS.n4516 0.0039507
R38019 DVSS.n4576 DVSS.n3799 0.0039507
R38020 DVSS.n4782 DVSS.n4781 0.0039507
R38021 DVSS DVSS.n7669 0.00392
R38022 DVSS.n7486 DVSS.n2310 0.00392
R38023 DVSS.n7668 DVSS 0.00392
R38024 DVSS.n9111 DVSS.n605 0.00392
R38025 DVSS.n9780 DVSS 0.00392
R38026 DVSS.n9060 DVSS.n9039 0.00392
R38027 DVSS.n8788 DVSS.n675 0.00392
R38028 DVSS DVSS.n9781 0.00392
R38029 DVSS.n8348 DVSS.n1436 0.00390714
R38030 DVSS.n1665 DVSS.n1427 0.00390714
R38031 DVSS.n8489 DVSS.n1114 0.00390714
R38032 DVSS.n1697 DVSS.n1107 0.00390714
R38033 DVSS.n1724 DVSS.n1713 0.00390714
R38034 DVSS.n1719 DVSS.n1594 0.00390714
R38035 DVSS.n1748 DVSS.n1571 0.00390714
R38036 DVSS.n1745 DVSS.n1564 0.00390714
R38037 DVSS.n7846 DVSS.n7737 0.00390714
R38038 DVSS.n7843 DVSS.n7730 0.00390714
R38039 DVSS.n8121 DVSS.n1822 0.00390714
R38040 DVSS.n1831 DVSS.n1808 0.00390714
R38041 DVSS.n8149 DVSS.n8138 0.00390714
R38042 DVSS.n8144 DVSS.n1788 0.00390714
R38043 DVSS.n8178 DVSS.n1770 0.00390714
R38044 DVSS.n8167 DVSS.n1763 0.00390714
R38045 DVSS.n5163 DVSS.n3326 0.00390714
R38046 DVSS.n5161 DVSS.n3325 0.00390714
R38047 DVSS.n5131 DVSS.n5065 0.00390714
R38048 DVSS.n5073 DVSS.n5068 0.00390714
R38049 DVSS.n5088 DVSS.n3372 0.00390714
R38050 DVSS.n5113 DVSS.n3371 0.00390714
R38051 DVSS.n5912 DVSS.n2949 0.00390714
R38052 DVSS.n5097 DVSS.n2942 0.00390714
R38053 DVSS.n5270 DVSS.n5269 0.00390714
R38054 DVSS.n5273 DVSS.n5272 0.00390714
R38055 DVSS.n5305 DVSS.n5304 0.00390714
R38056 DVSS.n5308 DVSS.n5307 0.00390714
R38057 DVSS.n5353 DVSS.n3386 0.00390714
R38058 DVSS.n5324 DVSS.n3379 0.00390714
R38059 DVSS.n5915 DVSS.n2931 0.00390714
R38060 DVSS.n5333 DVSS.n2924 0.00390714
R38061 DVSS.n4848 DVSS.n3660 0.00390714
R38062 DVSS.n3665 DVSS.n3647 0.00390714
R38063 DVSS.n4886 DVSS.n4881 0.00390714
R38064 DVSS.n3624 DVSS.n3614 0.00390714
R38065 DVSS.n4972 DVSS.n4961 0.00390714
R38066 DVSS.n3606 DVSS.n3600 0.00390714
R38067 DVSS.n4944 DVSS.n4912 0.00390714
R38068 DVSS.n4942 DVSS.n4935 0.00390714
R38069 DVSS.n8929 DVSS.n780 0.00386614
R38070 DVSS.n8964 DVSS.n733 0.00386614
R38071 DVSS.n9463 DVSS.n364 0.00386614
R38072 DVSS.n9498 DVSS.n32 0.00386614
R38073 DVSS.n4943 DVSS.n4934 0.00386614
R38074 DVSS.n4450 DVSS.n4449 0.00386614
R38075 DVSS.n7397 DVSS.n7395 0.00383
R38076 DVSS.n7417 DVSS.n7414 0.00383
R38077 DVSS.n7452 DVSS.n7450 0.00383
R38078 DVSS.n7059 DVSS.n6693 0.00383
R38079 DVSS.n1315 DVSS.n1033 0.00383
R38080 DVSS.n8559 DVSS.n1057 0.00383
R38081 DVSS.n8937 DVSS.n758 0.00383
R38082 DVSS.n7031 DVSS.n7030 0.00383
R38083 DVSS.n7003 DVSS.n807 0.00383
R38084 DVSS.n8691 DVSS.n725 0.00383
R38085 DVSS.n8715 DVSS.n8713 0.00383
R38086 DVSS.n8750 DVSS.n8748 0.00383
R38087 DVSS.n7501 DVSS.n2280 0.0038
R38088 DVSS.n9153 DVSS.n559 0.0038
R38089 DVSS.n9179 DVSS.n231 0.0038
R38090 DVSS.n9208 DVSS.n9197 0.0038
R38091 DVSS.n9180 DVSS.n238 0.0038
R38092 DVSS.n9260 DVSS.n500 0.0038
R38093 DVSS.n9288 DVSS.n486 0.0038
R38094 DVSS.n9287 DVSS.n9284 0.0038
R38095 DVSS.n9619 DVSS.n237 0.0038
R38096 DVSS.n9176 DVSS.n232 0.0038
R38097 DVSS.n4755 DVSS.n4754 0.00373944
R38098 DVSS.n1398 DVSS.n1392 0.00371429
R38099 DVSS.n7901 DVSS.n2062 0.00371429
R38100 DVSS.n5196 DVSS.n5011 0.00371429
R38101 DVSS.n3994 DVSS.n3474 0.00371429
R38102 DVSS.n4817 DVSS.n3679 0.00371429
R38103 DVSS.n7558 DVSS.n2234 0.00371
R38104 DVSS.n7616 DVSS.n2192 0.00371
R38105 DVSS.n7658 DVSS.n2158 0.00371
R38106 DVSS.n9661 DVSS.n9660 0.00371
R38107 DVSS.n9718 DVSS.n9717 0.00371
R38108 DVSS.n9770 DVSS.n139 0.00371
R38109 DVSS.n453 DVSS.n443 0.00371
R38110 DVSS.n9583 DVSS.n271 0.00371
R38111 DVSS.n341 DVSS.n75 0.00371
R38112 DVSS.n9296 DVSS.n392 0.00371
R38113 DVSS.n285 DVSS.n62 0.00371
R38114 DVSS.n9889 DVSS.n9888 0.00371
R38115 DVSS.n1121 DVSS.n1098 0.00368898
R38116 DVSS.n8350 DVSS.n1424 0.00368898
R38117 DVSS.n8362 DVSS.n1339 0.00368898
R38118 DVSS.n8454 DVSS.n1160 0.00368898
R38119 DVSS.n5558 DVSS.n2289 0.00366901
R38120 DVSS.n7883 DVSS.n2071 0.00366901
R38121 DVSS.n5612 DVSS.n2319 0.00366901
R38122 DVSS.n7885 DVSS.n2053 0.00366901
R38123 DVSS.n6767 DVSS.n6736 0.00365
R38124 DVSS.n6836 DVSS.n6689 0.00365
R38125 DVSS.n6822 DVSS.n1161 0.00365
R38126 DVSS.n8435 DVSS.n8434 0.00365
R38127 DVSS.n1939 DVSS.n1917 0.00365
R38128 DVSS.n8038 DVSS.n1950 0.00365
R38129 DVSS.n8015 DVSS.n1976 0.00365
R38130 DVSS.n7976 DVSS.n2010 0.00365
R38131 DVSS.n3078 DVSS.n2994 0.00365
R38132 DVSS.n3122 DVSS.n3117 0.00365
R38133 DVSS.n5778 DVSS.n3141 0.00365
R38134 DVSS.n5851 DVSS.n3027 0.00365
R38135 DVSS.n3896 DVSS.n3887 0.00365
R38136 DVSS.n3947 DVSS.n3946 0.00365
R38137 DVSS.n4236 DVSS.n3856 0.00365
R38138 DVSS.n4223 DVSS.n4222 0.00365
R38139 DVSS.n4207 DVSS.n4199 0.00365
R38140 DVSS.n4384 DVSS.n3719 0.00365
R38141 DVSS.n8812 DVSS.n624 0.00356
R38142 DVSS.n8813 DVSS.n632 0.00356
R38143 DVSS.n8811 DVSS.n8810 0.00356
R38144 DVSS.n8809 DVSS.n630 0.00356
R38145 DVSS.n9087 DVSS.n9086 0.00356
R38146 DVSS.n9088 DVSS.n625 0.00356
R38147 DVSS DVSS.n9849 0.00353
R38148 DVSS.n8909 DVSS.n764 0.00351181
R38149 DVSS.n9443 DVSS.n349 0.00351181
R38150 DVSS.n8387 DVSS.n8386 0.00345775
R38151 DVSS.n8377 DVSS.n1371 0.00345775
R38152 DVSS.n8400 DVSS.n8399 0.00345714
R38153 DVSS.n7936 DVSS.n2050 0.00345714
R38154 DVSS.n5741 DVSS.n3181 0.00345714
R38155 DVSS.n4103 DVSS.n3997 0.00345714
R38156 DVSS.n4302 DVSS.n3690 0.00345714
R38157 DVSS.n4677 DVSS 0.003425
R38158 DVSS.n4067 DVSS 0.003425
R38159 DVSS.n5218 DVSS 0.003425
R38160 DVSS DVSS.n3211 0.003425
R38161 DVSS.n5460 DVSS 0.003425
R38162 DVSS.n5599 DVSS 0.003425
R38163 DVSS.n7302 DVSS 0.003425
R38164 DVSS.n7933 DVSS 0.003425
R38165 DVSS.n7214 DVSS 0.003425
R38166 DVSS.n7490 DVSS.n7489 0.00338
R38167 DVSS.n9130 DVSS.n587 0.00338
R38168 DVSS.n9065 DVSS.n647 0.00338
R38169 DVSS.n8789 DVSS.n662 0.00338
R38170 DVSS.n1013 DVSS.n979 0.00334793
R38171 DVSS.n8654 DVSS.n8642 0.00334793
R38172 DVSS.n7384 DVSS.n7383 0.00334
R38173 DVSS.n7385 DVSS.n7384 0.00334
R38174 DVSS.n7385 DVSS.n2524 0.00334
R38175 DVSS.n7391 DVSS.n2524 0.00334
R38176 DVSS.n7392 DVSS.n7391 0.00334
R38177 DVSS.n7393 DVSS.n7392 0.00334
R38178 DVSS.n7393 DVSS.n2471 0.00334
R38179 DVSS.n7402 DVSS.n2471 0.00334
R38180 DVSS.n7403 DVSS.n7402 0.00334
R38181 DVSS.n7404 DVSS.n7403 0.00334
R38182 DVSS.n7404 DVSS.n2467 0.00334
R38183 DVSS.n7410 DVSS.n2467 0.00334
R38184 DVSS.n7411 DVSS.n7410 0.00334
R38185 DVSS.n7412 DVSS.n7411 0.00334
R38186 DVSS.n7412 DVSS.n2415 0.00334
R38187 DVSS.n7422 DVSS.n2415 0.00334
R38188 DVSS.n7423 DVSS.n7422 0.00334
R38189 DVSS.n7424 DVSS.n7423 0.00334
R38190 DVSS.n7424 DVSS.n2411 0.00334
R38191 DVSS.n7430 DVSS.n2411 0.00334
R38192 DVSS.n7431 DVSS.n7430 0.00334
R38193 DVSS.n7432 DVSS.n7431 0.00334
R38194 DVSS.n7432 DVSS.n2407 0.00334
R38195 DVSS.n7438 DVSS.n2407 0.00334
R38196 DVSS.n7439 DVSS.n7438 0.00334
R38197 DVSS.n7440 DVSS.n7439 0.00334
R38198 DVSS.n7440 DVSS.n2403 0.00334
R38199 DVSS.n7446 DVSS.n2403 0.00334
R38200 DVSS.n7447 DVSS.n7446 0.00334
R38201 DVSS.n7448 DVSS.n7447 0.00334
R38202 DVSS.n7448 DVSS.n2350 0.00334
R38203 DVSS.n7457 DVSS.n2350 0.00334
R38204 DVSS.n7458 DVSS.n7457 0.00334
R38205 DVSS.n7459 DVSS.n7458 0.00334
R38206 DVSS.n7459 DVSS.n2346 0.00334
R38207 DVSS.n7465 DVSS.n2346 0.00334
R38208 DVSS.n7466 DVSS.n7465 0.00334
R38209 DVSS.n7467 DVSS.n7466 0.00334
R38210 DVSS.n7467 DVSS.n2342 0.00334
R38211 DVSS.n7473 DVSS.n2342 0.00334
R38212 DVSS.n7474 DVSS.n7473 0.00334
R38213 DVSS.n7475 DVSS.n7474 0.00334
R38214 DVSS.n7475 DVSS.n2338 0.00334
R38215 DVSS.n7481 DVSS.n2338 0.00334
R38216 DVSS.n7482 DVSS.n7481 0.00334
R38217 DVSS.n7483 DVSS.n7482 0.00334
R38218 DVSS.n7483 DVSS.n2308 0.00334
R38219 DVSS.n7492 DVSS.n2308 0.00334
R38220 DVSS.n7493 DVSS.n7492 0.00334
R38221 DVSS.n7494 DVSS.n7493 0.00334
R38222 DVSS.n7494 DVSS.n2278 0.00334
R38223 DVSS.n7503 DVSS.n2278 0.00334
R38224 DVSS.n7504 DVSS.n7503 0.00334
R38225 DVSS.n7505 DVSS.n7504 0.00334
R38226 DVSS.n7505 DVSS.n2274 0.00334
R38227 DVSS.n7511 DVSS.n2274 0.00334
R38228 DVSS.n7512 DVSS.n7511 0.00334
R38229 DVSS.n7513 DVSS.n7512 0.00334
R38230 DVSS.n7513 DVSS.n2270 0.00334
R38231 DVSS.n7519 DVSS.n2270 0.00334
R38232 DVSS.n7520 DVSS.n7519 0.00334
R38233 DVSS.n7521 DVSS.n7520 0.00334
R38234 DVSS.n7521 DVSS.n2266 0.00334
R38235 DVSS.n7527 DVSS.n2266 0.00334
R38236 DVSS.n7528 DVSS.n7527 0.00334
R38237 DVSS.n7529 DVSS.n7528 0.00334
R38238 DVSS.n7529 DVSS.n2236 0.00334
R38239 DVSS.n7561 DVSS.n2236 0.00334
R38240 DVSS.n7562 DVSS.n7561 0.00334
R38241 DVSS.n7563 DVSS.n7562 0.00334
R38242 DVSS.n7563 DVSS.n2232 0.00334
R38243 DVSS.n7569 DVSS.n2232 0.00334
R38244 DVSS.n7570 DVSS.n7569 0.00334
R38245 DVSS.n7571 DVSS.n7570 0.00334
R38246 DVSS.n7571 DVSS.n2228 0.00334
R38247 DVSS.n7577 DVSS.n2228 0.00334
R38248 DVSS.n7578 DVSS.n7577 0.00334
R38249 DVSS.n7579 DVSS.n7578 0.00334
R38250 DVSS.n7579 DVSS.n2224 0.00334
R38251 DVSS.n7585 DVSS.n2224 0.00334
R38252 DVSS.n7586 DVSS.n7585 0.00334
R38253 DVSS.n7587 DVSS.n7586 0.00334
R38254 DVSS.n7587 DVSS.n2194 0.00334
R38255 DVSS.n7619 DVSS.n2194 0.00334
R38256 DVSS.n7620 DVSS.n7619 0.00334
R38257 DVSS.n7621 DVSS.n7620 0.00334
R38258 DVSS.n7621 DVSS.n2190 0.00334
R38259 DVSS.n7627 DVSS.n2190 0.00334
R38260 DVSS.n7628 DVSS.n7627 0.00334
R38261 DVSS.n7629 DVSS.n7628 0.00334
R38262 DVSS.n7629 DVSS.n2160 0.00334
R38263 DVSS.n7661 DVSS.n2160 0.00334
R38264 DVSS.n7662 DVSS.n7661 0.00334
R38265 DVSS.n7664 DVSS.n7662 0.00334
R38266 DVSS.n7664 DVSS.n7663 0.00334
R38267 DVSS.n7663 DVSS.n2157 0.00334
R38268 DVSS.n7673 DVSS.n7672 0.00334
R38269 DVSS.n6916 DVSS.n6732 0.00334
R38270 DVSS.n6917 DVSS.n6916 0.00334
R38271 DVSS.n6919 DVSS.n6917 0.00334
R38272 DVSS.n6919 DVSS.n6918 0.00334
R38273 DVSS.n6918 DVSS.n6728 0.00334
R38274 DVSS.n6926 DVSS.n6728 0.00334
R38275 DVSS.n6927 DVSS.n6926 0.00334
R38276 DVSS.n7043 DVSS.n6927 0.00334
R38277 DVSS.n7043 DVSS.n7042 0.00334
R38278 DVSS.n7042 DVSS.n7041 0.00334
R38279 DVSS.n7041 DVSS.n6928 0.00334
R38280 DVSS.n7037 DVSS.n6928 0.00334
R38281 DVSS.n7037 DVSS.n7036 0.00334
R38282 DVSS.n8597 DVSS.n8596 0.00334
R38283 DVSS.n8596 DVSS.n8595 0.00334
R38284 DVSS.n8595 DVSS.n1036 0.00334
R38285 DVSS.n8591 DVSS.n1036 0.00334
R38286 DVSS.n8591 DVSS.n8590 0.00334
R38287 DVSS.n8590 DVSS.n8589 0.00334
R38288 DVSS.n8589 DVSS.n1041 0.00334
R38289 DVSS.n8585 DVSS.n1041 0.00334
R38290 DVSS.n8585 DVSS.n8584 0.00334
R38291 DVSS.n8584 DVSS.n8583 0.00334
R38292 DVSS.n8583 DVSS.n1047 0.00334
R38293 DVSS.n8579 DVSS.n1047 0.00334
R38294 DVSS.n8579 DVSS.n8578 0.00334
R38295 DVSS.n8578 DVSS.n8577 0.00334
R38296 DVSS.n8577 DVSS.n1053 0.00334
R38297 DVSS.n8573 DVSS.n1053 0.00334
R38298 DVSS.n8573 DVSS.n8572 0.00334
R38299 DVSS.n8572 DVSS.n8571 0.00334
R38300 DVSS.n8571 DVSS.n1059 0.00334
R38301 DVSS.n8567 DVSS.n1059 0.00334
R38302 DVSS.n8567 DVSS.n8566 0.00334
R38303 DVSS.n8566 DVSS.n627 0.00334
R38304 DVSS.n9090 DVSS.n627 0.00334
R38305 DVSS.n9093 DVSS.n9092 0.00334
R38306 DVSS.n9093 DVSS.n622 0.00334
R38307 DVSS.n9099 DVSS.n622 0.00334
R38308 DVSS.n9100 DVSS.n9099 0.00334
R38309 DVSS.n9101 DVSS.n9100 0.00334
R38310 DVSS.n9101 DVSS.n618 0.00334
R38311 DVSS.n9107 DVSS.n618 0.00334
R38312 DVSS.n9108 DVSS.n9107 0.00334
R38313 DVSS.n9109 DVSS.n9108 0.00334
R38314 DVSS.n9109 DVSS.n585 0.00334
R38315 DVSS.n9133 DVSS.n585 0.00334
R38316 DVSS.n9134 DVSS.n9133 0.00334
R38317 DVSS.n9136 DVSS.n9134 0.00334
R38318 DVSS.n9136 DVSS.n9135 0.00334
R38319 DVSS.n9135 DVSS.n557 0.00334
R38320 DVSS.n9163 DVSS.n557 0.00334
R38321 DVSS.n9164 DVSS.n9163 0.00334
R38322 DVSS.n9165 DVSS.n9164 0.00334
R38323 DVSS.n9165 DVSS.n553 0.00334
R38324 DVSS.n9172 DVSS.n553 0.00334
R38325 DVSS.n9173 DVSS.n9172 0.00334
R38326 DVSS.n9174 DVSS.n9173 0.00334
R38327 DVSS.n9174 DVSS.n233 0.00334
R38328 DVSS.n9624 DVSS.n9623 0.00334
R38329 DVSS.n9624 DVSS.n229 0.00334
R38330 DVSS.n9630 DVSS.n229 0.00334
R38331 DVSS.n9631 DVSS.n9630 0.00334
R38332 DVSS.n9632 DVSS.n9631 0.00334
R38333 DVSS.n9632 DVSS.n202 0.00334
R38334 DVSS.n9663 DVSS.n202 0.00334
R38335 DVSS.n9664 DVSS.n9663 0.00334
R38336 DVSS.n9665 DVSS.n9664 0.00334
R38337 DVSS.n9665 DVSS.n198 0.00334
R38338 DVSS.n9671 DVSS.n198 0.00334
R38339 DVSS.n9672 DVSS.n9671 0.00334
R38340 DVSS.n9673 DVSS.n9672 0.00334
R38341 DVSS.n9673 DVSS.n194 0.00334
R38342 DVSS.n9679 DVSS.n194 0.00334
R38343 DVSS.n9680 DVSS.n9679 0.00334
R38344 DVSS.n9681 DVSS.n9680 0.00334
R38345 DVSS.n9681 DVSS.n190 0.00334
R38346 DVSS.n9687 DVSS.n190 0.00334
R38347 DVSS.n9688 DVSS.n9687 0.00334
R38348 DVSS.n9689 DVSS.n9688 0.00334
R38349 DVSS.n9689 DVSS.n163 0.00334
R38350 DVSS.n9720 DVSS.n163 0.00334
R38351 DVSS.n9722 DVSS.n160 0.00334
R38352 DVSS.n9729 DVSS.n160 0.00334
R38353 DVSS.n9730 DVSS.n9729 0.00334
R38354 DVSS.n9731 DVSS.n9730 0.00334
R38355 DVSS.n9731 DVSS.n141 0.00334
R38356 DVSS.n9773 DVSS.n141 0.00334
R38357 DVSS.n9774 DVSS.n9773 0.00334
R38358 DVSS.n9776 DVSS.n9774 0.00334
R38359 DVSS.n9776 DVSS.n9775 0.00334
R38360 DVSS.n9775 DVSS.n137 0.00334
R38361 DVSS.n9783 DVSS.n137 0.00334
R38362 DVSS.n9786 DVSS.n9784 0.00334
R38363 DVSS.n8621 DVSS.n8620 0.00334
R38364 DVSS.n8620 DVSS.n8619 0.00334
R38365 DVSS.n8619 DVSS.n1016 0.00334
R38366 DVSS.n8615 DVSS.n1016 0.00334
R38367 DVSS.n8615 DVSS.n8614 0.00334
R38368 DVSS.n8614 DVSS.n8613 0.00334
R38369 DVSS.n8613 DVSS.n1022 0.00334
R38370 DVSS.n8609 DVSS.n1022 0.00334
R38371 DVSS.n8609 DVSS.n8608 0.00334
R38372 DVSS.n8608 DVSS.n8607 0.00334
R38373 DVSS.n8607 DVSS.n1026 0.00334
R38374 DVSS.n8603 DVSS.n1026 0.00334
R38375 DVSS.n8603 DVSS.n8602 0.00334
R38376 DVSS.n6984 DVSS.n6982 0.00334
R38377 DVSS.n6985 DVSS.n6984 0.00334
R38378 DVSS.n7024 DVSS.n6985 0.00334
R38379 DVSS.n7024 DVSS.n7023 0.00334
R38380 DVSS.n7023 DVSS.n7022 0.00334
R38381 DVSS.n7022 DVSS.n6986 0.00334
R38382 DVSS.n7018 DVSS.n6986 0.00334
R38383 DVSS.n7018 DVSS.n7017 0.00334
R38384 DVSS.n7017 DVSS.n7016 0.00334
R38385 DVSS.n7016 DVSS.n6992 0.00334
R38386 DVSS.n7012 DVSS.n6992 0.00334
R38387 DVSS.n7012 DVSS.n7011 0.00334
R38388 DVSS.n7011 DVSS.n7010 0.00334
R38389 DVSS.n7010 DVSS.n6998 0.00334
R38390 DVSS.n7006 DVSS.n6998 0.00334
R38391 DVSS.n7006 DVSS.n7005 0.00334
R38392 DVSS.n7005 DVSS.n827 0.00334
R38393 DVSS.n8823 DVSS.n827 0.00334
R38394 DVSS.n8823 DVSS.n8822 0.00334
R38395 DVSS.n8822 DVSS.n8821 0.00334
R38396 DVSS.n8821 DVSS.n828 0.00334
R38397 DVSS.n8817 DVSS.n828 0.00334
R38398 DVSS.n8817 DVSS.n8816 0.00334
R38399 DVSS.n9085 DVSS.n9084 0.00334
R38400 DVSS.n9084 DVSS.n9083 0.00334
R38401 DVSS.n9083 DVSS.n634 0.00334
R38402 DVSS.n9079 DVSS.n634 0.00334
R38403 DVSS.n9079 DVSS.n9078 0.00334
R38404 DVSS.n9078 DVSS.n9077 0.00334
R38405 DVSS.n9077 DVSS.n640 0.00334
R38406 DVSS.n9073 DVSS.n640 0.00334
R38407 DVSS.n9073 DVSS.n9072 0.00334
R38408 DVSS.n9072 DVSS.n9071 0.00334
R38409 DVSS.n9071 DVSS.n646 0.00334
R38410 DVSS.n9067 DVSS.n646 0.00334
R38411 DVSS.n9067 DVSS.n539 0.00334
R38412 DVSS.n9195 DVSS.n539 0.00334
R38413 DVSS.n9195 DVSS.n9194 0.00334
R38414 DVSS.n9194 DVSS.n9193 0.00334
R38415 DVSS.n9193 DVSS.n540 0.00334
R38416 DVSS.n9189 DVSS.n540 0.00334
R38417 DVSS.n9189 DVSS.n9188 0.00334
R38418 DVSS.n9188 DVSS.n9187 0.00334
R38419 DVSS.n9187 DVSS.n546 0.00334
R38420 DVSS.n9183 DVSS.n546 0.00334
R38421 DVSS.n9183 DVSS.n235 0.00334
R38422 DVSS.n9620 DVSS.n236 0.00334
R38423 DVSS.n9616 DVSS.n236 0.00334
R38424 DVSS.n9616 DVSS.n9615 0.00334
R38425 DVSS.n9615 DVSS.n9614 0.00334
R38426 DVSS.n9614 DVSS.n242 0.00334
R38427 DVSS.n9610 DVSS.n242 0.00334
R38428 DVSS.n9610 DVSS.n9609 0.00334
R38429 DVSS.n9609 DVSS.n9608 0.00334
R38430 DVSS.n9608 DVSS.n247 0.00334
R38431 DVSS.n9604 DVSS.n247 0.00334
R38432 DVSS.n9604 DVSS.n9603 0.00334
R38433 DVSS.n9603 DVSS.n9602 0.00334
R38434 DVSS.n9602 DVSS.n252 0.00334
R38435 DVSS.n9598 DVSS.n252 0.00334
R38436 DVSS.n9598 DVSS.n9597 0.00334
R38437 DVSS.n9597 DVSS.n9596 0.00334
R38438 DVSS.n9596 DVSS.n258 0.00334
R38439 DVSS.n9592 DVSS.n258 0.00334
R38440 DVSS.n9592 DVSS.n9591 0.00334
R38441 DVSS.n9591 DVSS.n9590 0.00334
R38442 DVSS.n9590 DVSS.n264 0.00334
R38443 DVSS.n9586 DVSS.n264 0.00334
R38444 DVSS.n9586 DVSS.n9585 0.00334
R38445 DVSS.n9866 DVSS.n9865 0.00334
R38446 DVSS.n9865 DVSS.n9864 0.00334
R38447 DVSS.n9864 DVSS.n67 0.00334
R38448 DVSS.n9860 DVSS.n67 0.00334
R38449 DVSS.n9860 DVSS.n9859 0.00334
R38450 DVSS.n9859 DVSS.n9858 0.00334
R38451 DVSS.n9858 DVSS.n73 0.00334
R38452 DVSS.n9854 DVSS.n73 0.00334
R38453 DVSS.n9854 DVSS.n9853 0.00334
R38454 DVSS.n9853 DVSS.n9852 0.00334
R38455 DVSS.n9852 DVSS.n78 0.00334
R38456 DVSS.n9848 DVSS.n9847 0.00334
R38457 DVSS.n8685 DVSS.n962 0.00334
R38458 DVSS.n8686 DVSS.n8685 0.00334
R38459 DVSS.n8687 DVSS.n8686 0.00334
R38460 DVSS.n8687 DVSS.n958 0.00334
R38461 DVSS.n8694 DVSS.n958 0.00334
R38462 DVSS.n8695 DVSS.n8694 0.00334
R38463 DVSS.n8696 DVSS.n8695 0.00334
R38464 DVSS.n8696 DVSS.n955 0.00334
R38465 DVSS.n8701 DVSS.n955 0.00334
R38466 DVSS.n8702 DVSS.n8701 0.00334
R38467 DVSS.n8703 DVSS.n8702 0.00334
R38468 DVSS.n8703 DVSS.n952 0.00334
R38469 DVSS.n8709 DVSS.n952 0.00334
R38470 DVSS.n8711 DVSS.n900 0.00334
R38471 DVSS.n8720 DVSS.n900 0.00334
R38472 DVSS.n8721 DVSS.n8720 0.00334
R38473 DVSS.n8722 DVSS.n8721 0.00334
R38474 DVSS.n8722 DVSS.n896 0.00334
R38475 DVSS.n8728 DVSS.n896 0.00334
R38476 DVSS.n8729 DVSS.n8728 0.00334
R38477 DVSS.n8730 DVSS.n8729 0.00334
R38478 DVSS.n8730 DVSS.n892 0.00334
R38479 DVSS.n8736 DVSS.n892 0.00334
R38480 DVSS.n8737 DVSS.n8736 0.00334
R38481 DVSS.n8738 DVSS.n8737 0.00334
R38482 DVSS.n8738 DVSS.n888 0.00334
R38483 DVSS.n8744 DVSS.n888 0.00334
R38484 DVSS.n8745 DVSS.n8744 0.00334
R38485 DVSS.n8746 DVSS.n8745 0.00334
R38486 DVSS.n8746 DVSS.n837 0.00334
R38487 DVSS.n8755 DVSS.n837 0.00334
R38488 DVSS.n8756 DVSS.n8755 0.00334
R38489 DVSS.n8758 DVSS.n8756 0.00334
R38490 DVSS.n8758 DVSS.n8757 0.00334
R38491 DVSS.n8757 DVSS.n833 0.00334
R38492 DVSS.n8765 DVSS.n833 0.00334
R38493 DVSS.n8808 DVSS.n8807 0.00334
R38494 DVSS.n8807 DVSS.n8806 0.00334
R38495 DVSS.n8806 DVSS.n8767 0.00334
R38496 DVSS.n8802 DVSS.n8767 0.00334
R38497 DVSS.n8802 DVSS.n8801 0.00334
R38498 DVSS.n8801 DVSS.n8800 0.00334
R38499 DVSS.n8800 DVSS.n8772 0.00334
R38500 DVSS.n8796 DVSS.n8772 0.00334
R38501 DVSS.n8796 DVSS.n8795 0.00334
R38502 DVSS.n8795 DVSS.n8794 0.00334
R38503 DVSS.n8794 DVSS.n8777 0.00334
R38504 DVSS.n8777 DVSS.n497 0.00334
R38505 DVSS.n9263 DVSS.n497 0.00334
R38506 DVSS.n9264 DVSS.n9263 0.00334
R38507 DVSS.n9265 DVSS.n9264 0.00334
R38508 DVSS.n9265 DVSS.n493 0.00334
R38509 DVSS.n9271 DVSS.n493 0.00334
R38510 DVSS.n9272 DVSS.n9271 0.00334
R38511 DVSS.n9273 DVSS.n9272 0.00334
R38512 DVSS.n9273 DVSS.n489 0.00334
R38513 DVSS.n9280 DVSS.n489 0.00334
R38514 DVSS.n9281 DVSS.n9280 0.00334
R38515 DVSS.n9282 DVSS.n9281 0.00334
R38516 DVSS.n9286 DVSS.n9285 0.00334
R38517 DVSS.n9285 DVSS.n484 0.00334
R38518 DVSS.n9293 DVSS.n484 0.00334
R38519 DVSS.n9294 DVSS.n9293 0.00334
R38520 DVSS.n9350 DVSS.n9294 0.00334
R38521 DVSS.n9350 DVSS.n9349 0.00334
R38522 DVSS.n9349 DVSS.n9348 0.00334
R38523 DVSS.n9348 DVSS.n9295 0.00334
R38524 DVSS.n9344 DVSS.n9295 0.00334
R38525 DVSS.n9344 DVSS.n9343 0.00334
R38526 DVSS.n9343 DVSS.n9342 0.00334
R38527 DVSS.n9342 DVSS.n9300 0.00334
R38528 DVSS.n9338 DVSS.n9300 0.00334
R38529 DVSS.n9338 DVSS.n9337 0.00334
R38530 DVSS.n9337 DVSS.n9336 0.00334
R38531 DVSS.n9336 DVSS.n9306 0.00334
R38532 DVSS.n9332 DVSS.n9306 0.00334
R38533 DVSS.n9332 DVSS.n9331 0.00334
R38534 DVSS.n9331 DVSS.n9330 0.00334
R38535 DVSS.n9330 DVSS.n9313 0.00334
R38536 DVSS.n9326 DVSS.n9313 0.00334
R38537 DVSS.n9326 DVSS.n60 0.00334
R38538 DVSS.n9871 DVSS.n60 0.00334
R38539 DVSS.n9874 DVSS.n9873 0.00334
R38540 DVSS.n9874 DVSS.n55 0.00334
R38541 DVSS.n9880 DVSS.n55 0.00334
R38542 DVSS.n9881 DVSS.n9880 0.00334
R38543 DVSS.n9883 DVSS.n9881 0.00334
R38544 DVSS.n9883 DVSS.n9882 0.00334
R38545 DVSS.n9882 DVSS.n22 0.00334
R38546 DVSS.n9892 DVSS.n22 0.00334
R38547 DVSS.n9893 DVSS.n9892 0.00334
R38548 DVSS.n9894 DVSS.n9893 0.00334
R38549 DVSS.n9939 DVSS.n1 0.00334
R38550 DVSS.n7033 DVSS.n1033 0.00332
R38551 DVSS.n7032 DVSS.n7031 0.00332
R38552 DVSS.n8713 DVSS.n949 0.00332
R38553 DVSS.n8712 DVSS.n950 0.00332
R38554 DVSS.n8600 DVSS.n1031 0.00332
R38555 DVSS.n8599 DVSS.n8598 0.00332
R38556 DVSS.n7377 DVSS.n2530 0.00329
R38557 DVSS.n7396 DVSS.n2473 0.00329
R38558 DVSS.n7415 DVSS.n2417 0.00329
R38559 DVSS.n7451 DVSS.n2352 0.00329
R38560 DVSS.n6906 DVSS.n6886 0.00329
R38561 DVSS.n7055 DVSS.n6704 0.00329
R38562 DVSS.n1311 DVSS.n1202 0.00329
R38563 DVSS.n8542 DVSS.n1078 0.00329
R38564 DVSS.n8634 DVSS.n992 0.00329
R38565 DVSS.n770 DVSS.n755 0.00329
R38566 DVSS.n6967 DVSS.n6943 0.00329
R38567 DVSS.n824 DVSS.n808 0.00329
R38568 DVSS.n8677 DVSS.n8655 0.00329
R38569 DVSS.n957 DVSS.n724 0.00329
R38570 DVSS.n8714 DVSS.n902 0.00329
R38571 DVSS.n8749 DVSS.n839 0.00329
R38572 DVSS.n7672 DVSS 0.00326
R38573 DVSS.n7498 DVSS.n7497 0.00326
R38574 DVSS.n9156 DVSS.n9138 0.00326
R38575 DVSS.n9212 DVSS.n516 0.00326
R38576 DVSS.n9261 DVSS.n499 0.00326
R38577 DVSS.n9784 DVSS 0.00326
R38578 DVSS.n4656 DVSS.n3684 0.00324648
R38579 DVSS.n5564 DVSS.n2298 0.00324648
R38580 DVSS.n4667 DVSS.n3698 0.00324648
R38581 DVSS.n5598 DVSS.n2328 0.00324648
R38582 DVSS.n9894 DVSS 0.00322
R38583 DVSS.n7556 DVSS.n2253 0.00317
R38584 DVSS.n7559 DVSS.n2238 0.00317
R38585 DVSS.n7614 DVSS.n2211 0.00317
R38586 DVSS.n7617 DVSS.n2196 0.00317
R38587 DVSS.n7656 DVSS.n2177 0.00317
R38588 DVSS.n7659 DVSS.n2162 0.00317
R38589 DVSS.n7693 DVSS.n2121 0.00317
R38590 DVSS.n7675 DVSS.n2120 0.00317
R38591 DVSS.n9628 DVSS.n223 0.00317
R38592 DVSS.n222 DVSS.n204 0.00317
R38593 DVSS.n9685 DVSS.n184 0.00317
R38594 DVSS.n183 DVSS.n165 0.00317
R38595 DVSS.n9726 DVSS.n157 0.00317
R38596 DVSS.n9771 DVSS.n143 0.00317
R38597 DVSS.n9803 DVSS.n100 0.00317
R38598 DVSS.n135 DVSS.n99 0.00317
R38599 DVSS.n457 DVSS.n409 0.00317
R38600 DVSS.n408 DVSS.n245 0.00317
R38601 DVSS.n9580 DVSS.n9548 0.00317
R38602 DVSS.n9584 DVSS.n267 0.00317
R38603 DVSS.n9471 DVSS.n70 0.00317
R38604 DVSS.n343 DVSS.n74 0.00317
R38605 DVSS.n9844 DVSS.n9843 0.00317
R38606 DVSS.n9367 DVSS.n394 0.00317
R38607 DVSS.n482 DVSS.n393 0.00317
R38608 DVSS.n9544 DVSS.n288 0.00317
R38609 DVSS.n287 DVSS.n286 0.00317
R38610 DVSS.n9878 DVSS.n50 0.00317
R38611 DVSS.n49 DVSS.n24 0.00317
R38612 DVSS.n9932 DVSS.n9897 0.00317
R38613 DVSS.n19 DVSS.n5 0.00317
R38614 DVSS.n8884 DVSS.n785 0.00315748
R38615 DVSS.n8913 DVSS.n763 0.00315748
R38616 DVSS.n8948 DVSS.n739 0.00315748
R38617 DVSS.n9769 DVSS.n156 0.00315748
R38618 DVSS.n9447 DVSS.n348 0.00315748
R38619 DVSS.n9482 DVSS.n37 0.00315748
R38620 DVSS.n7676 DVSS.n7674 0.00309529
R38621 DVSS.n2529 DVSS.n2528 0.00309529
R38622 DVSS.n6885 DVSS.n6874 0.00309529
R38623 DVSS.n9785 DVSS.n136 0.00309529
R38624 DVSS.n9846 DVSS.n9845 0.00309529
R38625 DVSS.n9936 DVSS.n9935 0.00309529
R38626 DVSS.n7387 DVSS.n2526 0.00305
R38627 DVSS.n7406 DVSS.n2469 0.00305
R38628 DVSS.n7426 DVSS.n2413 0.00305
R38629 DVSS.n7461 DVSS.n2348 0.00305
R38630 DVSS.n6913 DVSS.n6730 0.00305
R38631 DVSS.n6929 DVSS.n6691 0.00305
R38632 DVSS.n1190 DVSS.n1039 0.00305
R38633 DVSS.n8562 DVSS.n8561 0.00305
R38634 DVSS.n1017 DVSS.n977 0.00305
R38635 DVSS.n1027 DVSS.n756 0.00305
R38636 DVSS.n6987 DVSS.n6979 0.00305
R38637 DVSS.n8859 DVSS.n810 0.00305
R38638 DVSS.n8682 DVSS.n960 0.00305
R38639 DVSS.n8996 DVSS.n738 0.00305
R38640 DVSS.n8724 DVSS.n898 0.00305
R38641 DVSS.n8760 DVSS.n835 0.00305
R38642 DVSS.n1238 DVSS.n566 0.00303521
R38643 DVSS.n1234 DVSS.n594 0.00303521
R38644 DVSS.n8495 DVSS.n1101 0.00298032
R38645 DVSS.n8353 DVSS.n1422 0.00298032
R38646 DVSS.n8371 DVSS.n1341 0.00298032
R38647 DVSS.n8457 DVSS.n1156 0.00298032
R38648 DVSS.n5996 DVSS.n2781 0.00296479
R38649 DVSS.n5969 DVSS.n2830 0.00296479
R38650 DVSS.n5952 DVSS.n2863 0.00296479
R38651 DVSS.n5937 DVSS.n2890 0.00296479
R38652 DVSS.n6344 DVSS.n6343 0.00287857
R38653 DVSS.n6032 DVSS.n6028 0.00287857
R38654 DVSS.n9722 DVSS.n9721 0.00286
R38655 DVSS.n9866 DVSS.n59 0.00286
R38656 DVSS.n9873 DVSS.n9872 0.00286
R38657 DVSS DVSS.n9939 0.00282
R38658 DVSS.n8926 DVSS.n779 0.00280315
R38659 DVSS.n8961 DVSS.n734 0.00280315
R38660 DVSS.n9460 DVSS.n363 0.00280315
R38661 DVSS.n9495 DVSS.n33 0.00280315
R38662 DVSS.n2157 DVSS 0.00278
R38663 DVSS.n4750 DVSS.n4749 0.00275352
R38664 DVSS.n1667 DVSS.n1426 0.00275
R38665 DVSS.n1699 DVSS.n1106 0.00275
R38666 DVSS.n1728 DVSS.n1727 0.00275
R38667 DVSS.n1586 DVSS.n1563 0.00275
R38668 DVSS.n7752 DVSS.n7729 0.00275
R38669 DVSS.n8124 DVSS.n8123 0.00275
R38670 DVSS.n8153 DVSS.n8152 0.00275
R38671 DVSS.n8174 DVSS.n1779 0.00275
R38672 DVSS.n5393 DVSS.n3328 0.00275
R38673 DVSS.n5128 DVSS.n5074 0.00275
R38674 DVSS.n5366 DVSS.n3374 0.00275
R38675 DVSS.n5095 DVSS.n2941 0.00275
R38676 DVSS.n3446 DVSS.n3436 0.00275
R38677 DVSS.n3411 DVSS.n3401 0.00275
R38678 DVSS.n5349 DVSS.n3393 0.00275
R38679 DVSS.n5331 DVSS.n2923 0.00275
R38680 DVSS.n4851 DVSS.n4850 0.00275
R38681 DVSS.n4889 DVSS.n4888 0.00275
R38682 DVSS.n4955 DVSS.n3599 0.00275
R38683 DVSS.n4941 DVSS.n4926 0.00275
R38684 DVSS.n7381 DVSS.n7380 0.00275
R38685 DVSS.n7400 DVSS.n7399 0.00275
R38686 DVSS.n7420 DVSS.n7419 0.00275
R38687 DVSS.n7455 DVSS.n7454 0.00275
R38688 DVSS.n6905 DVSS.n6734 0.00275
R38689 DVSS.n7045 DVSS.n6692 0.00275
R38690 DVSS.n1191 DVSS.n1037 0.00275
R38691 DVSS.n8534 DVSS.n1060 0.00275
R38692 DVSS.n8623 DVSS.n978 0.00275
R38693 DVSS.n1023 DVSS.n757 0.00275
R38694 DVSS.n7028 DVSS.n6968 0.00275
R38695 DVSS.n8856 DVSS.n8825 0.00275
R38696 DVSS.n8666 DVSS.n964 0.00275
R38697 DVSS.n8698 DVSS.n723 0.00275
R38698 DVSS.n8718 DVSS.n8717 0.00275
R38699 DVSS.n8753 DVSS.n8752 0.00275
R38700 DVSS.n9623 DVSS.n9622 0.0027
R38701 DVSS.n9621 DVSS.n9620 0.0027
R38702 DVSS.n9286 DVSS.n234 0.0027
R38703 DVSS.n4481 DVSS.n4461 0.0026831
R38704 DVSS.n4508 DVSS.n3825 0.0026831
R38705 DVSS.n4588 DVSS.n4579 0.0026831
R38706 DVSS.n4784 DVSS.n3735 0.0026831
R38707 DVSS.n7553 DVSS.n7531 0.00263
R38708 DVSS.n7553 DVSS.n7542 0.00263
R38709 DVSS.n7611 DVSS.n7589 0.00263
R38710 DVSS.n7611 DVSS.n7600 0.00263
R38711 DVSS.n7653 DVSS.n7631 0.00263
R38712 DVSS.n7653 DVSS.n7642 0.00263
R38713 DVSS.n7689 DVSS.n2134 0.00263
R38714 DVSS.n7689 DVSS.n7678 0.00263
R38715 DVSS.n9658 DVSS.n225 0.00263
R38716 DVSS.n9658 DVSS.n9634 0.00263
R38717 DVSS.n9715 DVSS.n186 0.00263
R38718 DVSS.n9715 DVSS.n9691 0.00263
R38719 DVSS.n9768 DVSS.n9733 0.00263
R38720 DVSS.n9768 DVSS.n9735 0.00263
R38721 DVSS.n9799 DVSS.n113 0.00263
R38722 DVSS.n9799 DVSS.n9788 0.00263
R38723 DVSS.n407 DVSS.n243 0.00263
R38724 DVSS.n407 DVSS.n244 0.00263
R38725 DVSS.n9576 DVSS.n265 0.00263
R38726 DVSS.n9576 DVSS.n266 0.00263
R38727 DVSS.n340 DVSS.n71 0.00263
R38728 DVSS.n342 DVSS.n340 0.00263
R38729 DVSS.n9839 DVSS.n82 0.00263
R38730 DVSS.n9839 DVSS.n85 0.00263
R38731 DVSS.n9363 DVSS.n460 0.00263
R38732 DVSS.n9363 DVSS.n9352 0.00263
R38733 DVSS.n9324 DVSS.n300 0.00263
R38734 DVSS.n9325 DVSS.n9324 0.00263
R38735 DVSS.n9886 DVSS.n52 0.00263
R38736 DVSS.n9886 DVSS.n9885 0.00263
R38737 DVSS.n9929 DVSS.n3 0.00263
R38738 DVSS.n9929 DVSS.n4 0.00263
R38739 DVSS.n1249 DVSS.n176 0.00262598
R38740 DVSS.n1242 DVSS.n215 0.00262598
R38741 DVSS.n1227 DVSS.n1072 0.00262598
R38742 DVSS.n1220 DVSS.n1201 0.00262598
R38743 DVSS.n8393 DVSS.n8392 0.00255714
R38744 DVSS.n2068 DVSS.n2060 0.00255714
R38745 DVSS.n5194 DVSS.n5016 0.00255714
R38746 DVSS.n5238 DVSS.n5237 0.00255714
R38747 DVSS.n3683 DVSS.n3677 0.00255714
R38748 DVSS.n9092 DVSS.n9091 0.00254
R38749 DVSS.n9085 DVSS.n626 0.00254
R38750 DVSS.n8808 DVSS.n8766 0.00254
R38751 DVSS.n7380 DVSS.n2543 0.00251
R38752 DVSS.n7399 DVSS.n2486 0.00251
R38753 DVSS.n7419 DVSS.n2430 0.00251
R38754 DVSS.n7454 DVSS.n2365 0.00251
R38755 DVSS.n6914 DVSS.n6734 0.00251
R38756 DVSS.n6726 DVSS.n6692 0.00251
R38757 DVSS.n1191 DVSS.n1038 0.00251
R38758 DVSS.n8534 DVSS.n1061 0.00251
R38759 DVSS.n1014 DVSS.n978 0.00251
R38760 DVSS.n1024 DVSS.n757 0.00251
R38761 DVSS.n7028 DVSS.n7026 0.00251
R38762 DVSS.n8856 DVSS.n809 0.00251
R38763 DVSS.n8683 DVSS.n964 0.00251
R38764 DVSS.n726 DVSS.n723 0.00251
R38765 DVSS.n8717 DVSS.n916 0.00251
R38766 DVSS.n8752 DVSS.n853 0.00251
R38767 DVSS.n6858 DVSS.n6744 0.00249286
R38768 DVSS.n7062 DVSS.n6675 0.00249286
R38769 DVSS.n8452 DVSS.n1171 0.00249286
R38770 DVSS.n8439 DVSS.n1334 0.00249286
R38771 DVSS.n8060 DVSS.n1925 0.00249286
R38772 DVSS.n1949 DVSS.n1945 0.00249286
R38773 DVSS.n1975 DVSS.n1971 0.00249286
R38774 DVSS.n2009 DVSS.n2005 0.00249286
R38775 DVSS.n5879 DVSS.n3003 0.00249286
R38776 DVSS.n5813 DVSS.n3105 0.00249286
R38777 DVSS.n3140 DVSS.n3136 0.00249286
R38778 DVSS.n5864 DVSS.n5854 0.00249286
R38779 DVSS.n4186 DVSS.n4172 0.00249286
R38780 DVSS.n4139 DVSS.n3936 0.00249286
R38781 DVSS.n4451 DVSS.n3845 0.00249286
R38782 DVSS.n4258 DVSS.n4252 0.00249286
R38783 DVSS.n4429 DVSS.n4418 0.00249286
R38784 DVSS.n4796 DVSS.n3726 0.00249286
R38785 DVSS DVSS.n5945 0.00247183
R38786 DVSS.n4607 DVSS.n3783 0.00247183
R38787 DVSS.n5944 DVSS 0.00247183
R38788 DVSS.n8897 DVSS.n773 0.00244882
R38789 DVSS.n8995 DVSS.n8994 0.00244882
R38790 DVSS.n9431 DVSS.n357 0.00244882
R38791 DVSS.n9528 DVSS.n47 0.00244882
R38792 DVSS.n5017 DVSS.n3515 0.00240141
R38793 DVSS.n5572 DVSS.n2283 0.00240141
R38794 DVSS.n3512 DVSS.n3182 0.00240141
R38795 DVSS.n5582 DVSS.n2313 0.00240141
R38796 DVSS.n8597 DVSS.n1035 0.00238
R38797 DVSS.n6982 DVSS.n951 0.00238
R38798 DVSS.n8711 DVSS.n8710 0.00238
R38799 DVSS.n4946 DVSS 0.0023
R38800 DVSS.n1739 DVSS 0.0023
R38801 DVSS.n1388 DVSS.n1377 0.0023
R38802 DVSS DVSS.n1565 0.0023
R38803 DVSS.n8165 DVSS 0.0023
R38804 DVSS.n7937 DVSS.n2044 0.0023
R38805 DVSS DVSS.n1764 0.0023
R38806 DVSS DVSS.n5102 0.0023
R38807 DVSS.n5742 DVSS.n3175 0.0023
R38808 DVSS DVSS.n2943 0.0023
R38809 DVSS DVSS.n5338 0.0023
R38810 DVSS.n4105 DVSS.n3976 0.0023
R38811 DVSS DVSS.n2925 0.0023
R38812 DVSS.n4353 DVSS.n3703 0.0023
R38813 DVSS.n4945 DVSS 0.0023
R38814 DVSS.n6443 VSS 0.0023
R38815 DVSS.n6166 VSS 0.0023
R38816 VSS DVSS.n6167 0.0023
R38817 DVSS.n6442 VSS 0.0023
R38818 DVSS.n2543 DVSS.n2526 0.00221
R38819 DVSS.n2486 DVSS.n2469 0.00221
R38820 DVSS.n2430 DVSS.n2413 0.00221
R38821 DVSS.n2365 DVSS.n2348 0.00221
R38822 DVSS.n6914 DVSS.n6913 0.00221
R38823 DVSS.n6726 DVSS.n6691 0.00221
R38824 DVSS.n1190 DVSS.n1038 0.00221
R38825 DVSS.n8561 DVSS.n1061 0.00221
R38826 DVSS.n1014 DVSS.n977 0.00221
R38827 DVSS.n1024 DVSS.n756 0.00221
R38828 DVSS.n7026 DVSS.n6979 0.00221
R38829 DVSS.n8859 DVSS.n809 0.00221
R38830 DVSS.n8683 DVSS.n8682 0.00221
R38831 DVSS.n8996 DVSS.n726 0.00221
R38832 DVSS.n916 DVSS.n898 0.00221
R38833 DVSS.n853 DVSS.n835 0.00221
R38834 DVSS.n8977 DVSS.n745 0.00209449
R38835 DVSS.n9511 DVSS.n43 0.00209449
R38836 DVSS.n7556 DVSS.n7531 0.00209
R38837 DVSS.n7542 DVSS.n2238 0.00209
R38838 DVSS.n7614 DVSS.n7589 0.00209
R38839 DVSS.n7600 DVSS.n2196 0.00209
R38840 DVSS.n7656 DVSS.n7631 0.00209
R38841 DVSS.n7642 DVSS.n2162 0.00209
R38842 DVSS.n7693 DVSS.n2134 0.00209
R38843 DVSS.n7678 DVSS.n2120 0.00209
R38844 DVSS.n225 DVSS.n223 0.00209
R38845 DVSS.n9634 DVSS.n222 0.00209
R38846 DVSS.n186 DVSS.n184 0.00209
R38847 DVSS.n9691 DVSS.n183 0.00209
R38848 DVSS.n9733 DVSS.n157 0.00209
R38849 DVSS.n9735 DVSS.n143 0.00209
R38850 DVSS.n9803 DVSS.n113 0.00209
R38851 DVSS.n9788 DVSS.n99 0.00209
R38852 DVSS.n457 DVSS.n243 0.00209
R38853 DVSS.n408 DVSS.n244 0.00209
R38854 DVSS.n9580 DVSS.n265 0.00209
R38855 DVSS.n267 DVSS.n266 0.00209
R38856 DVSS.n9471 DVSS.n71 0.00209
R38857 DVSS.n343 DVSS.n342 0.00209
R38858 DVSS.n9841 DVSS.n82 0.00209
R38859 DVSS.n9843 DVSS.n85 0.00209
R38860 DVSS.n9367 DVSS.n460 0.00209
R38861 DVSS.n9352 DVSS.n393 0.00209
R38862 DVSS.n9544 DVSS.n300 0.00209
R38863 DVSS.n9325 DVSS.n287 0.00209
R38864 DVSS.n52 DVSS.n50 0.00209
R38865 DVSS.n9885 DVSS.n49 0.00209
R38866 DVSS.n9932 DVSS.n3 0.00209
R38867 DVSS.n19 DVSS.n4 0.00209
R38868 DVSS.n7498 DVSS.n7496 0.002
R38869 DVSS.n9156 DVSS.n575 0.002
R38870 DVSS.n9212 DVSS.n503 0.002
R38871 DVSS.n8790 DVSS.n499 0.002
R38872 DVSS.n5236 DVSS.n5235 0.00197887
R38873 DVSS.n5573 DVSS.n2302 0.00197887
R38874 DVSS.n5233 DVSS.n3489 0.00197887
R38875 DVSS.n5581 DVSS.n2332 0.00197887
R38876 DVSS.n7381 DVSS.n2530 0.00197
R38877 DVSS.n7400 DVSS.n2473 0.00197
R38878 DVSS.n7420 DVSS.n2417 0.00197
R38879 DVSS.n7455 DVSS.n2352 0.00197
R38880 DVSS.n6906 DVSS.n6905 0.00197
R38881 DVSS.n7055 DVSS.n7045 0.00197
R38882 DVSS.n1311 DVSS.n1037 0.00197
R38883 DVSS.n1078 DVSS.n1060 0.00197
R38884 DVSS.n8634 DVSS.n8623 0.00197
R38885 DVSS.n1023 DVSS.n755 0.00197
R38886 DVSS.n6968 DVSS.n6967 0.00197
R38887 DVSS.n8825 DVSS.n808 0.00197
R38888 DVSS.n8677 DVSS.n8666 0.00197
R38889 DVSS.n8698 DVSS.n724 0.00197
R38890 DVSS.n8718 DVSS.n902 0.00197
R38891 DVSS.n8753 DVSS.n839 0.00197
R38892 DVSS DVSS.n78 0.00196
R38893 DVSS.n7034 DVSS.n7033 0.00194
R38894 DVSS.n7032 DVSS.n1030 0.00194
R38895 DVSS.n9841 DVSS 0.00194
R38896 DVSS.n8707 DVSS.n949 0.00194
R38897 DVSS.n8708 DVSS.n950 0.00194
R38898 DVSS.n8601 DVSS.n8600 0.00194
R38899 DVSS.n8599 DVSS.n1032 0.00194
R38900 DVSS.n7489 DVSS.n2306 0.00188
R38901 DVSS.n9131 DVSS.n9130 0.00188
R38902 DVSS.n9066 DVSS.n9065 0.00188
R38903 DVSS.n8791 DVSS.n662 0.00188
R38904 DVSS.n9848 DVSS 0.00188
R38905 DVSS.n8978 DVSS.n730 0.00174016
R38906 DVSS.n9512 DVSS.n29 0.00174016
R38907 DVSS DVSS.n81 0.00173
R38908 DVSS.n9850 DVSS 0.00173
R38909 DVSS.n8812 DVSS.n629 0.0017
R38910 DVSS.n8814 DVSS.n8813 0.0017
R38911 DVSS.n8811 DVSS.n830 0.0017
R38912 DVSS.n8764 DVSS.n630 0.0017
R38913 DVSS.n9087 DVSS.n631 0.0017
R38914 DVSS.n9089 DVSS.n9088 0.0017
R38915 DVSS.n1083 DVSS.n570 0.00155634
R38916 DVSS.n8525 DVSS.n598 0.00155634
R38917 DVSS.n7559 DVSS.n7558 0.00155
R38918 DVSS.n7617 DVSS.n7616 0.00155
R38919 DVSS.n7659 DVSS.n7658 0.00155
R38920 DVSS.n7675 DVSS.n2119 0.00155
R38921 DVSS.n9660 DVSS.n204 0.00155
R38922 DVSS.n9717 DVSS.n165 0.00155
R38923 DVSS.n9771 DVSS.n9770 0.00155
R38924 DVSS.n135 DVSS.n98 0.00155
R38925 DVSS.n453 DVSS.n245 0.00155
R38926 DVSS.n9584 DVSS.n9583 0.00155
R38927 DVSS.n341 DVSS.n74 0.00155
R38928 DVSS.n9844 DVSS.n84 0.00155
R38929 DVSS.n482 DVSS.n392 0.00155
R38930 DVSS.n286 DVSS.n285 0.00155
R38931 DVSS.n9888 DVSS.n24 0.00155
R38932 DVSS.n9934 DVSS.n5 0.00155
R38933 DVSS.n4746 DVSS.n4622 0.00148592
R38934 DVSS.n7497 DVSS.n2280 0.00146
R38935 DVSS.n9153 DVSS.n9138 0.00146
R38936 DVSS.n9179 DVSS.n9178 0.00146
R38937 DVSS.n9208 DVSS.n516 0.00146
R38938 DVSS.n9181 DVSS.n9180 0.00146
R38939 DVSS.n9261 DVSS.n9260 0.00146
R38940 DVSS.n488 DVSS.n486 0.00146
R38941 DVSS.n9284 DVSS.n9283 0.00146
R38942 DVSS.n9182 DVSS.n237 0.00146
R38943 DVSS.n9177 DVSS.n9176 0.00146
R38944 DVSS.n7036 DVSS.n1035 0.00146
R38945 DVSS.n8602 DVSS.n951 0.00146
R38946 DVSS.n8710 DVSS.n8709 0.00146
R38947 DVSS.n7378 DVSS.n7377 0.00143
R38948 DVSS.n7397 DVSS.n7396 0.00143
R38949 DVSS.n7417 DVSS.n7415 0.00143
R38950 DVSS.n7452 DVSS.n7451 0.00143
R38951 DVSS.n6910 DVSS.n6886 0.00143
R38952 DVSS.n7059 DVSS.n6704 0.00143
R38953 DVSS.n1315 DVSS.n1202 0.00143
R38954 DVSS.n8559 DVSS.n8542 0.00143
R38955 DVSS.n8638 DVSS.n992 0.00143
R38956 DVSS.n8937 DVSS.n770 0.00143
R38957 DVSS.n7030 DVSS.n6943 0.00143
R38958 DVSS.n824 DVSS.n807 0.00143
R38959 DVSS.n8680 DVSS.n8655 0.00143
R38960 DVSS.n957 DVSS.n725 0.00143
R38961 DVSS.n8715 DVSS.n8714 0.00143
R38962 DVSS.n8750 DVSS.n8749 0.00143
R38963 DVSS.n8388 DVSS.n1404 0.0014
R38964 DVSS.n7770 DVSS.n2061 0.0014
R38965 DVSS.n5193 DVSS.n5010 0.0014
R38966 DVSS.n3480 DVSS.n3470 0.0014
R38967 DVSS.n4346 DVSS.n3678 0.0014
R38968 DVSS.n8507 DVSS.n180 0.00138583
R38969 DVSS.n8513 DVSS.n219 0.00138583
R38970 DVSS.n8560 DVSS.n8532 0.00138583
R38971 DVSS.n1297 DVSS.n1296 0.00138583
R38972 DVSS.n8896 DVSS.n767 0.00138583
R38973 DVSS.n749 DVSS.n727 0.00138583
R38974 DVSS.n9430 DVSS.n352 0.00138583
R38975 DVSS.n9527 DVSS.n26 0.00138583
R38976 DVSS.n4628 DVSS.n4617 0.00134507
R38977 DVSS.n1267 DVSS.n568 0.00134507
R38978 DVSS.n4693 DVSS.n3771 0.00134507
R38979 DVSS.n1276 DVSS.n596 0.00134507
R38980 DVSS.n7670 DVSS 0.00134
R38981 DVSS.n7490 DVSS.n2310 0.00134
R38982 DVSS DVSS.n2121 0.00134
R38983 DVSS.n605 DVSS.n587 0.00134
R38984 DVSS DVSS.n100 0.00134
R38985 DVSS.n9060 DVSS.n647 0.00134
R38986 DVSS.n8789 DVSS.n8788 0.00134
R38987 DVSS.n9782 DVSS 0.00134
R38988 DVSS.n9091 DVSS.n9090 0.0013
R38989 DVSS.n8816 DVSS.n626 0.0013
R38990 DVSS.n8766 DVSS.n8765 0.0013
R38991 DVSS.n9718 DVSS.n162 0.00122
R38992 DVSS.n271 DVSS.n270 0.00122
R38993 DVSS.n269 DVSS.n62 0.00122
R38994 DVSS.n9870 DVSS.n9869 0.00122
R38995 DVSS.n9868 DVSS.n64 0.00122
R38996 DVSS.n9719 DVSS.n63 0.00122
R38997 DVSS.n1257 DVSS.n178 0.00120866
R38998 DVSS.n1262 DVSS.n217 0.00120866
R38999 DVSS.n1282 DVSS.n1074 0.00120866
R39000 DVSS.n1287 DVSS.n1203 0.00120866
R39001 DVSS.n4757 DVSS.n3775 0.00120422
R39002 DVSS.n8403 DVSS.n1367 0.00114286
R39003 DVSS.n2043 DVSS.n2039 0.00114286
R39004 DVSS.n3174 DVSS.n3170 0.00114286
R39005 DVSS.n4106 DVSS.n3969 0.00114286
R39006 DVSS.n4809 DVSS.n3697 0.00114286
R39007 DVSS.n9622 DVSS.n233 0.00114
R39008 DVSS.n9621 DVSS.n235 0.00114
R39009 DVSS.n9282 DVSS.n234 0.00114
R39010 DVSS.n5565 DVSS.n2286 0.0011338
R39011 DVSS.n5597 DVSS.n2316 0.0011338
R39012 DVSS.n7671 DVSS 0.00106
R39013 DVSS.n8927 DVSS.n760 0.0010315
R39014 DVSS.n8962 DVSS.n742 0.0010315
R39015 DVSS.n9461 DVSS.n345 0.0010315
R39016 DVSS.n9496 DVSS.n40 0.0010315
R39017 DVSS DVSS.n0 0.00102
R39018 DVSS.n9721 DVSS.n9720 0.00098
R39019 DVSS.n9585 DVSS.n59 0.00098
R39020 DVSS.n9872 DVSS.n9871 0.00098
R39021 DVSS.n8382 DVSS.n1401 0.000922535
R39022 DVSS.n8373 DVSS.n1364 0.000922535
R39023 DVSS.n7501 DVSS.n7500 0.00092
R39024 DVSS.n9159 DVSS.n559 0.00092
R39025 DVSS.n9197 DVSS.n502 0.00092
R39026 DVSS.n500 DVSS.n495 0.00092
R39027 DVSS.n8491 DVSS.n8490 0.000854331
R39028 DVSS.n8349 DVSS.n1417 0.000854331
R39029 DVSS.n8367 DVSS.n1331 0.000854331
R39030 DVSS.n8453 DVSS.n1152 0.000854331
R39031 DVSS.n7487 DVSS.n7486 0.0008
R39032 DVSS.n9128 DVSS.n9111 0.0008
R39033 DVSS.n9063 DVSS.n9039 0.0008
R39034 DVSS.n9026 DVSS.n675 0.0008
R39035 DVSS.n5557 DVSS.n2295 0.000711268
R39036 DVSS.n7884 DVSS.n2065 0.000711268
R39037 DVSS.n5613 DVSS.n2325 0.000711268
R39038 DVSS.n7886 DVSS.n2047 0.000711268
R39039 DVSS DVSS.n2875 0.000687793
R39040 DVSS.n9897 DVSS 0.00068
R39041 DVSS DVSS.n2 0.00068
R39042 DVSS.n8912 DVSS.n776 0.000677165
R39043 DVSS.n8947 DVSS.n737 0.000677165
R39044 DVSS.n9446 DVSS.n360 0.000677165
R39045 DVSS.n9481 DVSS.n36 0.000677165
R39046 DVSS.n4947 DVSS 0.000671429
R39047 DVSS DVSS.n1740 0.000671429
R39048 DVSS.n8164 DVSS 0.000671429
R39049 DVSS.n5101 DVSS 0.000671429
R39050 DVSS.n5337 DVSS 0.000671429
R39051 DVSS.n6444 VSS 0.000671429
R39052 DVSS.n6165 VSS 0.000671429
R39053 DVSS DVSS.n0 0.00062
R39054 DVSS DVSS.n7671 0.00058
R39055 DVSS DVSS.n9783 0.00058
R39056 ASIG5V.n3081 ASIG5V 7.63331
R39057 ASIG5V.n3087 ASIG5V 7.63331
R39058 ASIG5V.n3094 ASIG5V 7.63331
R39059 ASIG5V.n3101 ASIG5V 7.63331
R39060 ASIG5V.n3108 ASIG5V 7.63331
R39061 ASIG5V.n3122 ASIG5V 7.63331
R39062 ASIG5V.n9901 ASIG5V 7.63331
R39063 ASIG5V.n3115 ASIG5V 7.63331
R39064 ASIG5V.n3083 ASIG5V.n3067 4.5005
R39065 ASIG5V.n7472 ASIG5V.n7469 4.5005
R39066 ASIG5V.n7472 ASIG5V.n3067 4.5005
R39067 ASIG5V.n7470 ASIG5V.n3067 4.5005
R39068 ASIG5V.n8105 ASIG5V.n7470 4.5005
R39069 ASIG5V.n8107 ASIG5V.n3067 4.5005
R39070 ASIG5V.n9892 ASIG5V.n3081 4.5005
R39071 ASIG5V.n9887 ASIG5V.n3080 4.5005
R39072 ASIG5V.n9892 ASIG5V.n3080 4.5005
R39073 ASIG5V.n9892 ASIG5V.n3079 4.5005
R39074 ASIG5V.n9889 ASIG5V.n3079 4.5005
R39075 ASIG5V.n9892 ASIG5V.n9891 4.5005
R39076 ASIG5V.n8115 ASIG5V.n8109 4.5005
R39077 ASIG5V.n8115 ASIG5V.n7466 4.5005
R39078 ASIG5V.n7466 ASIG5V.n3056 4.5005
R39079 ASIG5V.n8114 ASIG5V.n3056 4.5005
R39080 ASIG5V.n8115 ASIG5V.n8114 4.5005
R39081 ASIG5V.n8111 ASIG5V.n7465 4.5005
R39082 ASIG5V.n8115 ASIG5V.n7465 4.5005
R39083 ASIG5V.n8116 ASIG5V.n8115 4.5005
R39084 ASIG5V.n7633 ASIG5V.n7464 4.5005
R39085 ASIG5V.n7631 ASIG5V.n7623 4.5005
R39086 ASIG5V.n7631 ASIG5V.n7464 4.5005
R39087 ASIG5V.n7626 ASIG5V.n7464 4.5005
R39088 ASIG5V.n7630 ASIG5V.n7626 4.5005
R39089 ASIG5V.n7624 ASIG5V.n7464 4.5005
R39090 ASIG5V.n8098 ASIG5V.n7475 4.5005
R39091 ASIG5V.n8091 ASIG5V.n7474 4.5005
R39092 ASIG5V.n8098 ASIG5V.n7474 4.5005
R39093 ASIG5V.n8096 ASIG5V.n7479 4.5005
R39094 ASIG5V.n8096 ASIG5V.n8095 4.5005
R39095 ASIG5V.n8095 ASIG5V.n7476 4.5005
R39096 ASIG5V.n9882 ASIG5V.n3087 4.5005
R39097 ASIG5V.n9875 ASIG5V.n3086 4.5005
R39098 ASIG5V.n9882 ASIG5V.n3086 4.5005
R39099 ASIG5V.n9880 ASIG5V.n3091 4.5005
R39100 ASIG5V.n9880 ASIG5V.n9879 4.5005
R39101 ASIG5V.n9879 ASIG5V.n3088 4.5005
R39102 ASIG5V.n8128 ASIG5V.n7315 4.5005
R39103 ASIG5V.n8117 ASIG5V.n3045 4.5005
R39104 ASIG5V.n8128 ASIG5V.n7312 4.5005
R39105 ASIG5V.n8126 ASIG5V.n7312 4.5005
R39106 ASIG5V.n7461 ASIG5V.n7460 4.5005
R39107 ASIG5V.n7461 ASIG5V.n3045 4.5005
R39108 ASIG5V.n8127 ASIG5V.n8126 4.5005
R39109 ASIG5V.n8128 ASIG5V.n8127 4.5005
R39110 ASIG5V.n8122 ASIG5V.n7320 4.5005
R39111 ASIG5V.n8125 ASIG5V.n7320 4.5005
R39112 ASIG5V.n7318 ASIG5V.n7311 4.5005
R39113 ASIG5V.n8128 ASIG5V.n7311 4.5005
R39114 ASIG5V.n8125 ASIG5V.n8124 4.5005
R39115 ASIG5V.n8129 ASIG5V.n8128 4.5005
R39116 ASIG5V.n7617 ASIG5V.n7310 4.5005
R39117 ASIG5V.n7613 ASIG5V.n7575 4.5005
R39118 ASIG5V.n7613 ASIG5V.n7310 4.5005
R39119 ASIG5V.n7609 ASIG5V.n7310 4.5005
R39120 ASIG5V.n7610 ASIG5V.n7609 4.5005
R39121 ASIG5V.n7607 ASIG5V.n7310 4.5005
R39122 ASIG5V.n7637 ASIG5V.n7636 4.5005
R39123 ASIG5V.n7620 ASIG5V.n7618 4.5005
R39124 ASIG5V.n7637 ASIG5V.n7620 4.5005
R39125 ASIG5V.n7641 ASIG5V.n7570 4.5005
R39126 ASIG5V.n7644 ASIG5V.n7570 4.5005
R39127 ASIG5V.n7644 ASIG5V.n7643 4.5005
R39128 ASIG5V.n8089 ASIG5V.n7482 4.5005
R39129 ASIG5V.n8082 ASIG5V.n7481 4.5005
R39130 ASIG5V.n8089 ASIG5V.n7481 4.5005
R39131 ASIG5V.n8087 ASIG5V.n7486 4.5005
R39132 ASIG5V.n8087 ASIG5V.n8086 4.5005
R39133 ASIG5V.n8086 ASIG5V.n7483 4.5005
R39134 ASIG5V.n9873 ASIG5V.n3094 4.5005
R39135 ASIG5V.n9866 ASIG5V.n3093 4.5005
R39136 ASIG5V.n9873 ASIG5V.n3093 4.5005
R39137 ASIG5V.n9871 ASIG5V.n3098 4.5005
R39138 ASIG5V.n9871 ASIG5V.n9870 4.5005
R39139 ASIG5V.n9870 ASIG5V.n3095 4.5005
R39140 ASIG5V.n8141 ASIG5V.n7294 4.5005
R39141 ASIG5V.n8131 ASIG5V.n8130 4.5005
R39142 ASIG5V.n7459 ASIG5V.n3034 4.5005
R39143 ASIG5V.n8141 ASIG5V.n7291 4.5005
R39144 ASIG5V.n8139 ASIG5V.n7291 4.5005
R39145 ASIG5V.n7306 ASIG5V.n7304 4.5005
R39146 ASIG5V.n8131 ASIG5V.n7306 4.5005
R39147 ASIG5V.n7457 ASIG5V.n7326 4.5005
R39148 ASIG5V.n7326 ASIG5V.n3034 4.5005
R39149 ASIG5V.n8140 ASIG5V.n8139 4.5005
R39150 ASIG5V.n8141 ASIG5V.n8140 4.5005
R39151 ASIG5V.n7455 ASIG5V.n7451 4.5005
R39152 ASIG5V.n7451 ASIG5V.n7307 4.5005
R39153 ASIG5V.n8135 ASIG5V.n7299 4.5005
R39154 ASIG5V.n8138 ASIG5V.n7299 4.5005
R39155 ASIG5V.n7297 ASIG5V.n7290 4.5005
R39156 ASIG5V.n8141 ASIG5V.n7290 4.5005
R39157 ASIG5V.n7449 ASIG5V.n7307 4.5005
R39158 ASIG5V.n8138 ASIG5V.n8137 4.5005
R39159 ASIG5V.n8142 ASIG5V.n8141 4.5005
R39160 ASIG5V.n7592 ASIG5V.n7591 4.5005
R39161 ASIG5V.n7587 ASIG5V.n7582 4.5005
R39162 ASIG5V.n7591 ASIG5V.n7582 4.5005
R39163 ASIG5V.n7591 ASIG5V.n7581 4.5005
R39164 ASIG5V.n7588 ASIG5V.n7581 4.5005
R39165 ASIG5V.n7591 ASIG5V.n7590 4.5005
R39166 ASIG5V.n7604 ASIG5V.n7566 4.5005
R39167 ASIG5V.n7598 ASIG5V.n7577 4.5005
R39168 ASIG5V.n7604 ASIG5V.n7577 4.5005
R39169 ASIG5V.n7602 ASIG5V.n7601 4.5005
R39170 ASIG5V.n7602 ASIG5V.n7557 4.5005
R39171 ASIG5V.n7593 ASIG5V.n7557 4.5005
R39172 ASIG5V.n7646 ASIG5V.n7645 4.5005
R39173 ASIG5V.n7569 ASIG5V.n7567 4.5005
R39174 ASIG5V.n7646 ASIG5V.n7569 4.5005
R39175 ASIG5V.n7650 ASIG5V.n7562 4.5005
R39176 ASIG5V.n7653 ASIG5V.n7562 4.5005
R39177 ASIG5V.n7653 ASIG5V.n7652 4.5005
R39178 ASIG5V.n8080 ASIG5V.n7489 4.5005
R39179 ASIG5V.n8073 ASIG5V.n7488 4.5005
R39180 ASIG5V.n8080 ASIG5V.n7488 4.5005
R39181 ASIG5V.n8078 ASIG5V.n7493 4.5005
R39182 ASIG5V.n8078 ASIG5V.n8077 4.5005
R39183 ASIG5V.n8077 ASIG5V.n7490 4.5005
R39184 ASIG5V.n9864 ASIG5V.n3101 4.5005
R39185 ASIG5V.n9857 ASIG5V.n3100 4.5005
R39186 ASIG5V.n9864 ASIG5V.n3100 4.5005
R39187 ASIG5V.n9862 ASIG5V.n3105 4.5005
R39188 ASIG5V.n9862 ASIG5V.n9861 4.5005
R39189 ASIG5V.n9861 ASIG5V.n3102 4.5005
R39190 ASIG5V.n8154 ASIG5V.n7274 4.5005
R39191 ASIG5V.n8144 ASIG5V.n8143 4.5005
R39192 ASIG5V.n7369 ASIG5V.n7303 4.5005
R39193 ASIG5V.n7448 ASIG5V.n3023 4.5005
R39194 ASIG5V.n8154 ASIG5V.n7271 4.5005
R39195 ASIG5V.n8152 ASIG5V.n7271 4.5005
R39196 ASIG5V.n7286 ASIG5V.n7284 4.5005
R39197 ASIG5V.n8144 ASIG5V.n7286 4.5005
R39198 ASIG5V.n7370 ASIG5V.n7366 4.5005
R39199 ASIG5V.n7370 ASIG5V.n7369 4.5005
R39200 ASIG5V.n7446 ASIG5V.n7330 4.5005
R39201 ASIG5V.n7330 ASIG5V.n3023 4.5005
R39202 ASIG5V.n8153 ASIG5V.n8152 4.5005
R39203 ASIG5V.n8154 ASIG5V.n8153 4.5005
R39204 ASIG5V.n7444 ASIG5V.n7440 4.5005
R39205 ASIG5V.n7440 ASIG5V.n7328 4.5005
R39206 ASIG5V.n7375 ASIG5V.n7367 4.5005
R39207 ASIG5V.n7367 ASIG5V.n7287 4.5005
R39208 ASIG5V.n8148 ASIG5V.n7279 4.5005
R39209 ASIG5V.n8151 ASIG5V.n7279 4.5005
R39210 ASIG5V.n7277 ASIG5V.n7270 4.5005
R39211 ASIG5V.n8154 ASIG5V.n7270 4.5005
R39212 ASIG5V.n7438 ASIG5V.n7328 4.5005
R39213 ASIG5V.n7377 ASIG5V.n7287 4.5005
R39214 ASIG5V.n8151 ASIG5V.n8150 4.5005
R39215 ASIG5V.n8155 ASIG5V.n8154 4.5005
R39216 ASIG5V.n7688 ASIG5V.n7269 4.5005
R39217 ASIG5V.n7690 ASIG5V.n7546 4.5005
R39218 ASIG5V.n7690 ASIG5V.n7269 4.5005
R39219 ASIG5V.n7547 ASIG5V.n7269 4.5005
R39220 ASIG5V.n7695 ASIG5V.n7547 4.5005
R39221 ASIG5V.n7697 ASIG5V.n7269 4.5005
R39222 ASIG5V.n7678 ASIG5V.n7677 4.5005
R39223 ASIG5V.n7679 ASIG5V.n7549 4.5005
R39224 ASIG5V.n7679 ASIG5V.n7678 4.5005
R39225 ASIG5V.n7684 ASIG5V.n7550 4.5005
R39226 ASIG5V.n7550 ASIG5V.n7518 4.5005
R39227 ASIG5V.n7686 ASIG5V.n7518 4.5005
R39228 ASIG5V.n7667 ASIG5V.n7666 4.5005
R39229 ASIG5V.n7668 ASIG5V.n7554 4.5005
R39230 ASIG5V.n7668 ASIG5V.n7667 4.5005
R39231 ASIG5V.n7673 ASIG5V.n7555 4.5005
R39232 ASIG5V.n7555 ASIG5V.n7513 4.5005
R39233 ASIG5V.n7675 ASIG5V.n7513 4.5005
R39234 ASIG5V.n7656 ASIG5V.n7655 4.5005
R39235 ASIG5V.n7657 ASIG5V.n7559 4.5005
R39236 ASIG5V.n7657 ASIG5V.n7656 4.5005
R39237 ASIG5V.n7662 ASIG5V.n7560 4.5005
R39238 ASIG5V.n7560 ASIG5V.n7508 4.5005
R39239 ASIG5V.n7664 ASIG5V.n7508 4.5005
R39240 ASIG5V.n8071 ASIG5V.n7496 4.5005
R39241 ASIG5V.n8064 ASIG5V.n7495 4.5005
R39242 ASIG5V.n8071 ASIG5V.n7495 4.5005
R39243 ASIG5V.n8069 ASIG5V.n7500 4.5005
R39244 ASIG5V.n8069 ASIG5V.n8068 4.5005
R39245 ASIG5V.n8068 ASIG5V.n7497 4.5005
R39246 ASIG5V.n9855 ASIG5V.n3108 4.5005
R39247 ASIG5V.n9848 ASIG5V.n3107 4.5005
R39248 ASIG5V.n9855 ASIG5V.n3107 4.5005
R39249 ASIG5V.n9853 ASIG5V.n3112 4.5005
R39250 ASIG5V.n9853 ASIG5V.n9852 4.5005
R39251 ASIG5V.n9852 ASIG5V.n3109 4.5005
R39252 ASIG5V.n7698 ASIG5V.n7528 4.5005
R39253 ASIG5V.n8157 ASIG5V.n8156 4.5005
R39254 ASIG5V.n7387 ASIG5V.n7283 4.5005
R39255 ASIG5V.n7379 ASIG5V.n7378 4.5005
R39256 ASIG5V.n7437 ASIG5V.n3012 4.5005
R39257 ASIG5V.n7700 ASIG5V.n7528 4.5005
R39258 ASIG5V.n7700 ASIG5V.n7258 4.5005
R39259 ASIG5V.n8158 ASIG5V.n7264 4.5005
R39260 ASIG5V.n8158 ASIG5V.n8157 4.5005
R39261 ASIG5V.n7388 ASIG5V.n7354 4.5005
R39262 ASIG5V.n7388 ASIG5V.n7387 4.5005
R39263 ASIG5V.n7363 ASIG5V.n7361 4.5005
R39264 ASIG5V.n7379 ASIG5V.n7363 4.5005
R39265 ASIG5V.n7435 ASIG5V.n7334 4.5005
R39266 ASIG5V.n7334 ASIG5V.n3012 4.5005
R39267 ASIG5V.n7544 ASIG5V.n7258 4.5005
R39268 ASIG5V.n7544 ASIG5V.n7528 4.5005
R39269 ASIG5V.n7433 ASIG5V.n7429 4.5005
R39270 ASIG5V.n7429 ASIG5V.n7332 4.5005
R39271 ASIG5V.n7383 ASIG5V.n7357 4.5005
R39272 ASIG5V.n7386 ASIG5V.n7357 4.5005
R39273 ASIG5V.n7355 ASIG5V.n7349 4.5005
R39274 ASIG5V.n7390 ASIG5V.n7349 4.5005
R39275 ASIG5V.n7265 ASIG5V.n7259 4.5005
R39276 ASIG5V.n8160 ASIG5V.n7259 4.5005
R39277 ASIG5V.n7702 ASIG5V.n7541 4.5005
R39278 ASIG5V.n7541 ASIG5V.n7528 4.5005
R39279 ASIG5V.n7427 ASIG5V.n7332 4.5005
R39280 ASIG5V.n7386 ASIG5V.n7385 4.5005
R39281 ASIG5V.n7391 ASIG5V.n7390 4.5005
R39282 ASIG5V.n8161 ASIG5V.n8160 4.5005
R39283 ASIG5V.n7704 ASIG5V.n7528 4.5005
R39284 ASIG5V.n9764 ASIG5V.n9763 4.5005
R39285 ASIG5V.n9759 ASIG5V.n3152 4.5005
R39286 ASIG5V.n9763 ASIG5V.n3152 4.5005
R39287 ASIG5V.n9763 ASIG5V.n3151 4.5005
R39288 ASIG5V.n9760 ASIG5V.n3151 4.5005
R39289 ASIG5V.n9763 ASIG5V.n9762 4.5005
R39290 ASIG5V.n9776 ASIG5V.n9775 4.5005
R39291 ASIG5V.n9767 ASIG5V.n3146 4.5005
R39292 ASIG5V.n9775 ASIG5V.n3146 4.5005
R39293 ASIG5V.n9773 ASIG5V.n9769 4.5005
R39294 ASIG5V.n9773 ASIG5V.n9772 4.5005
R39295 ASIG5V.n9772 ASIG5V.n9765 4.5005
R39296 ASIG5V.n9788 ASIG5V.n9787 4.5005
R39297 ASIG5V.n9779 ASIG5V.n3141 4.5005
R39298 ASIG5V.n9787 ASIG5V.n3141 4.5005
R39299 ASIG5V.n9785 ASIG5V.n9781 4.5005
R39300 ASIG5V.n9785 ASIG5V.n9784 4.5005
R39301 ASIG5V.n9784 ASIG5V.n9777 4.5005
R39302 ASIG5V.n9800 ASIG5V.n9799 4.5005
R39303 ASIG5V.n9791 ASIG5V.n3136 4.5005
R39304 ASIG5V.n9799 ASIG5V.n3136 4.5005
R39305 ASIG5V.n9797 ASIG5V.n9793 4.5005
R39306 ASIG5V.n9797 ASIG5V.n9796 4.5005
R39307 ASIG5V.n9796 ASIG5V.n9789 4.5005
R39308 ASIG5V.n9812 ASIG5V.n9811 4.5005
R39309 ASIG5V.n9803 ASIG5V.n3131 4.5005
R39310 ASIG5V.n9811 ASIG5V.n3131 4.5005
R39311 ASIG5V.n9809 ASIG5V.n9805 4.5005
R39312 ASIG5V.n9809 ASIG5V.n9808 4.5005
R39313 ASIG5V.n9808 ASIG5V.n9801 4.5005
R39314 ASIG5V.n9824 ASIG5V.n9823 4.5005
R39315 ASIG5V.n9815 ASIG5V.n3126 4.5005
R39316 ASIG5V.n9823 ASIG5V.n3126 4.5005
R39317 ASIG5V.n9821 ASIG5V.n9817 4.5005
R39318 ASIG5V.n9821 ASIG5V.n9820 4.5005
R39319 ASIG5V.n9820 ASIG5V.n9813 4.5005
R39320 ASIG5V.n9837 ASIG5V.n3122 4.5005
R39321 ASIG5V.n9830 ASIG5V.n3121 4.5005
R39322 ASIG5V.n9837 ASIG5V.n3121 4.5005
R39323 ASIG5V.n9835 ASIG5V.n9828 4.5005
R39324 ASIG5V.n9835 ASIG5V.n9834 4.5005
R39325 ASIG5V.n9834 ASIG5V.n9825 4.5005
R39326 ASIG5V.n9754 ASIG5V.n9753 4.5005
R39327 ASIG5V.n7705 ASIG5V.n7247 4.5005
R39328 ASIG5V.n8163 ASIG5V.n8162 4.5005
R39329 ASIG5V.n7404 ASIG5V.n7392 4.5005
R39330 ASIG5V.n7413 ASIG5V.n7338 4.5005
R39331 ASIG5V.n7426 ASIG5V.n3009 4.5005
R39332 ASIG5V.n9753 ASIG5V.n3158 4.5005
R39333 ASIG5V.n7988 ASIG5V.n3158 4.5005
R39334 ASIG5V.n7538 ASIG5V.n7537 4.5005
R39335 ASIG5V.n7538 ASIG5V.n7247 4.5005
R39336 ASIG5V.n8164 ASIG5V.n7253 4.5005
R39337 ASIG5V.n8164 ASIG5V.n8163 4.5005
R39338 ASIG5V.n7397 ASIG5V.n7346 4.5005
R39339 ASIG5V.n7404 ASIG5V.n7346 4.5005
R39340 ASIG5V.n7406 ASIG5V.n7337 4.5005
R39341 ASIG5V.n7413 ASIG5V.n7337 4.5005
R39342 ASIG5V.n7424 ASIG5V.n7416 4.5005
R39343 ASIG5V.n7416 ASIG5V.n3009 4.5005
R39344 ASIG5V.n7988 ASIG5V.n3161 4.5005
R39345 ASIG5V.n9753 ASIG5V.n3161 4.5005
R39346 ASIG5V.n7422 ASIG5V.n7418 4.5005
R39347 ASIG5V.n7418 ASIG5V.n7414 4.5005
R39348 ASIG5V.n7411 ASIG5V.n7344 4.5005
R39349 ASIG5V.n7411 ASIG5V.n7410 4.5005
R39350 ASIG5V.n7402 ASIG5V.n7395 4.5005
R39351 ASIG5V.n7402 ASIG5V.n7401 4.5005
R39352 ASIG5V.n7254 ASIG5V.n7248 4.5005
R39353 ASIG5V.n8166 ASIG5V.n7248 4.5005
R39354 ASIG5V.n7710 ASIG5V.n7533 4.5005
R39355 ASIG5V.n7713 ASIG5V.n7533 4.5005
R39356 ASIG5V.n9750 ASIG5V.n3157 4.5005
R39357 ASIG5V.n9753 ASIG5V.n3157 4.5005
R39358 ASIG5V.n7414 ASIG5V.n1841 4.5005
R39359 ASIG5V.n7410 ASIG5V.n7341 4.5005
R39360 ASIG5V.n7401 ASIG5V.n169 4.5005
R39361 ASIG5V.n8167 ASIG5V.n8166 4.5005
R39362 ASIG5V.n7713 ASIG5V.n7712 4.5005
R39363 ASIG5V.n9753 ASIG5V.n9752 4.5005
R39364 ASIG5V.n9943 ASIG5V.n3004 4.5005
R39365 ASIG5V.n3008 ASIG5V.n3005 4.5005
R39366 ASIG5V.n3008 ASIG5V.n3004 4.5005
R39367 ASIG5V.n3006 ASIG5V.n3004 4.5005
R39368 ASIG5V.n9950 ASIG5V.n3006 4.5005
R39369 ASIG5V.n9952 ASIG5V.n3004 4.5005
R39370 ASIG5V.n9938 ASIG5V.n9937 4.5005
R39371 ASIG5V.n9939 ASIG5V.n3018 4.5005
R39372 ASIG5V.n9939 ASIG5V.n9938 4.5005
R39373 ASIG5V.n3019 ASIG5V.n3013 4.5005
R39374 ASIG5V.n9941 ASIG5V.n3013 4.5005
R39375 ASIG5V.n9942 ASIG5V.n9941 4.5005
R39376 ASIG5V.n9932 ASIG5V.n9931 4.5005
R39377 ASIG5V.n9933 ASIG5V.n3029 4.5005
R39378 ASIG5V.n9933 ASIG5V.n9932 4.5005
R39379 ASIG5V.n3030 ASIG5V.n3024 4.5005
R39380 ASIG5V.n9935 ASIG5V.n3024 4.5005
R39381 ASIG5V.n9936 ASIG5V.n9935 4.5005
R39382 ASIG5V.n9926 ASIG5V.n9925 4.5005
R39383 ASIG5V.n9927 ASIG5V.n3040 4.5005
R39384 ASIG5V.n9927 ASIG5V.n9926 4.5005
R39385 ASIG5V.n3041 ASIG5V.n3035 4.5005
R39386 ASIG5V.n9929 ASIG5V.n3035 4.5005
R39387 ASIG5V.n9930 ASIG5V.n9929 4.5005
R39388 ASIG5V.n9920 ASIG5V.n9919 4.5005
R39389 ASIG5V.n9921 ASIG5V.n3051 4.5005
R39390 ASIG5V.n9921 ASIG5V.n9920 4.5005
R39391 ASIG5V.n3052 ASIG5V.n3046 4.5005
R39392 ASIG5V.n9923 ASIG5V.n3046 4.5005
R39393 ASIG5V.n9924 ASIG5V.n9923 4.5005
R39394 ASIG5V.n9914 ASIG5V.n9913 4.5005
R39395 ASIG5V.n9915 ASIG5V.n3062 4.5005
R39396 ASIG5V.n9915 ASIG5V.n9914 4.5005
R39397 ASIG5V.n3063 ASIG5V.n3057 4.5005
R39398 ASIG5V.n9917 ASIG5V.n3057 4.5005
R39399 ASIG5V.n9918 ASIG5V.n9917 4.5005
R39400 ASIG5V.n9908 ASIG5V.n9907 4.5005
R39401 ASIG5V.n9909 ASIG5V.n3073 4.5005
R39402 ASIG5V.n9909 ASIG5V.n9908 4.5005
R39403 ASIG5V.n3074 ASIG5V.n3068 4.5005
R39404 ASIG5V.n9911 ASIG5V.n3068 4.5005
R39405 ASIG5V.n9912 ASIG5V.n9911 4.5005
R39406 ASIG5V.n9902 ASIG5V.n9901 4.5005
R39407 ASIG5V.n9903 ASIG5V.n9898 4.5005
R39408 ASIG5V.n9903 ASIG5V.n9902 4.5005
R39409 ASIG5V.n9899 ASIG5V.n9893 4.5005
R39410 ASIG5V.n9905 ASIG5V.n9893 4.5005
R39411 ASIG5V.n9906 ASIG5V.n9905 4.5005
R39412 ASIG5V.n4255 ASIG5V.n3909 4.5005
R39413 ASIG5V.n4051 ASIG5V.n3909 4.5005
R39414 ASIG5V.n3909 ASIG5V.n3858 4.5005
R39415 ASIG5V.n3909 ASIG5V.n3855 4.5005
R39416 ASIG5V.n10911 ASIG5V.n10548 4.5005
R39417 ASIG5V.n10548 ASIG5V.n10492 4.5005
R39418 ASIG5V.n10548 ASIG5V.n10495 4.5005
R39419 ASIG5V.n10548 ASIG5V.n10493 4.5005
R39420 ASIG5V.n4255 ASIG5V.n3908 4.5005
R39421 ASIG5V.n3908 ASIG5V.n3858 4.5005
R39422 ASIG5V.n3908 ASIG5V.n3857 4.5005
R39423 ASIG5V.n10911 ASIG5V.n10545 4.5005
R39424 ASIG5V.n10545 ASIG5V.n10492 4.5005
R39425 ASIG5V.n10545 ASIG5V.n10495 4.5005
R39426 ASIG5V.n10911 ASIG5V.n10551 4.5005
R39427 ASIG5V.n10551 ASIG5V.n10495 4.5005
R39428 ASIG5V.n10551 ASIG5V.n10494 4.5005
R39429 ASIG5V.n10911 ASIG5V.n10544 4.5005
R39430 ASIG5V.n10544 ASIG5V.n10495 4.5005
R39431 ASIG5V.n10544 ASIG5V.n10494 4.5005
R39432 ASIG5V.n10911 ASIG5V.n10554 4.5005
R39433 ASIG5V.n10554 ASIG5V.n10495 4.5005
R39434 ASIG5V.n10554 ASIG5V.n10494 4.5005
R39435 ASIG5V.n10911 ASIG5V.n10543 4.5005
R39436 ASIG5V.n10543 ASIG5V.n10495 4.5005
R39437 ASIG5V.n10543 ASIG5V.n10494 4.5005
R39438 ASIG5V.n10911 ASIG5V.n10557 4.5005
R39439 ASIG5V.n10557 ASIG5V.n10495 4.5005
R39440 ASIG5V.n10557 ASIG5V.n10494 4.5005
R39441 ASIG5V.n10911 ASIG5V.n10542 4.5005
R39442 ASIG5V.n10542 ASIG5V.n10495 4.5005
R39443 ASIG5V.n10542 ASIG5V.n10494 4.5005
R39444 ASIG5V.n10911 ASIG5V.n10560 4.5005
R39445 ASIG5V.n10560 ASIG5V.n10495 4.5005
R39446 ASIG5V.n10560 ASIG5V.n10494 4.5005
R39447 ASIG5V.n10911 ASIG5V.n10541 4.5005
R39448 ASIG5V.n10541 ASIG5V.n10495 4.5005
R39449 ASIG5V.n10541 ASIG5V.n10494 4.5005
R39450 ASIG5V.n10911 ASIG5V.n10563 4.5005
R39451 ASIG5V.n10563 ASIG5V.n10495 4.5005
R39452 ASIG5V.n10563 ASIG5V.n10494 4.5005
R39453 ASIG5V.n10911 ASIG5V.n10540 4.5005
R39454 ASIG5V.n10540 ASIG5V.n10495 4.5005
R39455 ASIG5V.n10540 ASIG5V.n10494 4.5005
R39456 ASIG5V.n10911 ASIG5V.n10566 4.5005
R39457 ASIG5V.n10566 ASIG5V.n10495 4.5005
R39458 ASIG5V.n10566 ASIG5V.n10494 4.5005
R39459 ASIG5V.n10911 ASIG5V.n10539 4.5005
R39460 ASIG5V.n10539 ASIG5V.n10495 4.5005
R39461 ASIG5V.n10539 ASIG5V.n10494 4.5005
R39462 ASIG5V.n10911 ASIG5V.n10569 4.5005
R39463 ASIG5V.n10569 ASIG5V.n10495 4.5005
R39464 ASIG5V.n10569 ASIG5V.n10494 4.5005
R39465 ASIG5V.n10911 ASIG5V.n10538 4.5005
R39466 ASIG5V.n10538 ASIG5V.n10495 4.5005
R39467 ASIG5V.n10538 ASIG5V.n10494 4.5005
R39468 ASIG5V.n10911 ASIG5V.n10572 4.5005
R39469 ASIG5V.n10572 ASIG5V.n10495 4.5005
R39470 ASIG5V.n10572 ASIG5V.n10494 4.5005
R39471 ASIG5V.n10911 ASIG5V.n10537 4.5005
R39472 ASIG5V.n10537 ASIG5V.n10495 4.5005
R39473 ASIG5V.n10537 ASIG5V.n10494 4.5005
R39474 ASIG5V.n10911 ASIG5V.n10575 4.5005
R39475 ASIG5V.n10575 ASIG5V.n10495 4.5005
R39476 ASIG5V.n10575 ASIG5V.n10494 4.5005
R39477 ASIG5V.n10911 ASIG5V.n10536 4.5005
R39478 ASIG5V.n10536 ASIG5V.n10495 4.5005
R39479 ASIG5V.n10536 ASIG5V.n10494 4.5005
R39480 ASIG5V.n10911 ASIG5V.n10578 4.5005
R39481 ASIG5V.n10578 ASIG5V.n10495 4.5005
R39482 ASIG5V.n10578 ASIG5V.n10494 4.5005
R39483 ASIG5V.n10911 ASIG5V.n10535 4.5005
R39484 ASIG5V.n10535 ASIG5V.n10495 4.5005
R39485 ASIG5V.n10535 ASIG5V.n10494 4.5005
R39486 ASIG5V.n10911 ASIG5V.n10581 4.5005
R39487 ASIG5V.n10581 ASIG5V.n10495 4.5005
R39488 ASIG5V.n10581 ASIG5V.n10494 4.5005
R39489 ASIG5V.n10911 ASIG5V.n10534 4.5005
R39490 ASIG5V.n10534 ASIG5V.n10495 4.5005
R39491 ASIG5V.n10534 ASIG5V.n10494 4.5005
R39492 ASIG5V.n10911 ASIG5V.n10584 4.5005
R39493 ASIG5V.n10584 ASIG5V.n10495 4.5005
R39494 ASIG5V.n10584 ASIG5V.n10494 4.5005
R39495 ASIG5V.n10911 ASIG5V.n10533 4.5005
R39496 ASIG5V.n10533 ASIG5V.n10495 4.5005
R39497 ASIG5V.n10533 ASIG5V.n10494 4.5005
R39498 ASIG5V.n10911 ASIG5V.n10587 4.5005
R39499 ASIG5V.n10587 ASIG5V.n10495 4.5005
R39500 ASIG5V.n10587 ASIG5V.n10494 4.5005
R39501 ASIG5V.n10911 ASIG5V.n10532 4.5005
R39502 ASIG5V.n10532 ASIG5V.n10495 4.5005
R39503 ASIG5V.n10532 ASIG5V.n10494 4.5005
R39504 ASIG5V.n10911 ASIG5V.n10590 4.5005
R39505 ASIG5V.n10590 ASIG5V.n10495 4.5005
R39506 ASIG5V.n10590 ASIG5V.n10494 4.5005
R39507 ASIG5V.n10911 ASIG5V.n10531 4.5005
R39508 ASIG5V.n10531 ASIG5V.n10495 4.5005
R39509 ASIG5V.n10531 ASIG5V.n10494 4.5005
R39510 ASIG5V.n10911 ASIG5V.n10593 4.5005
R39511 ASIG5V.n10593 ASIG5V.n10495 4.5005
R39512 ASIG5V.n10593 ASIG5V.n10494 4.5005
R39513 ASIG5V.n10911 ASIG5V.n10530 4.5005
R39514 ASIG5V.n10530 ASIG5V.n10495 4.5005
R39515 ASIG5V.n10530 ASIG5V.n10494 4.5005
R39516 ASIG5V.n10911 ASIG5V.n10596 4.5005
R39517 ASIG5V.n10596 ASIG5V.n10495 4.5005
R39518 ASIG5V.n10596 ASIG5V.n10494 4.5005
R39519 ASIG5V.n10911 ASIG5V.n10529 4.5005
R39520 ASIG5V.n10529 ASIG5V.n10495 4.5005
R39521 ASIG5V.n10529 ASIG5V.n10494 4.5005
R39522 ASIG5V.n10911 ASIG5V.n10599 4.5005
R39523 ASIG5V.n10599 ASIG5V.n10495 4.5005
R39524 ASIG5V.n10599 ASIG5V.n10494 4.5005
R39525 ASIG5V.n10911 ASIG5V.n10528 4.5005
R39526 ASIG5V.n10528 ASIG5V.n10495 4.5005
R39527 ASIG5V.n10528 ASIG5V.n10494 4.5005
R39528 ASIG5V.n10911 ASIG5V.n10602 4.5005
R39529 ASIG5V.n10602 ASIG5V.n10495 4.5005
R39530 ASIG5V.n10602 ASIG5V.n10494 4.5005
R39531 ASIG5V.n10911 ASIG5V.n10527 4.5005
R39532 ASIG5V.n10527 ASIG5V.n10495 4.5005
R39533 ASIG5V.n10527 ASIG5V.n10494 4.5005
R39534 ASIG5V.n10911 ASIG5V.n10605 4.5005
R39535 ASIG5V.n10605 ASIG5V.n10495 4.5005
R39536 ASIG5V.n10605 ASIG5V.n10494 4.5005
R39537 ASIG5V.n10911 ASIG5V.n10526 4.5005
R39538 ASIG5V.n10526 ASIG5V.n10495 4.5005
R39539 ASIG5V.n10526 ASIG5V.n10494 4.5005
R39540 ASIG5V.n10911 ASIG5V.n10608 4.5005
R39541 ASIG5V.n10608 ASIG5V.n10495 4.5005
R39542 ASIG5V.n10608 ASIG5V.n10494 4.5005
R39543 ASIG5V.n10911 ASIG5V.n10525 4.5005
R39544 ASIG5V.n10525 ASIG5V.n10495 4.5005
R39545 ASIG5V.n10525 ASIG5V.n10494 4.5005
R39546 ASIG5V.n10911 ASIG5V.n10611 4.5005
R39547 ASIG5V.n10611 ASIG5V.n10495 4.5005
R39548 ASIG5V.n10611 ASIG5V.n10494 4.5005
R39549 ASIG5V.n10911 ASIG5V.n10524 4.5005
R39550 ASIG5V.n10524 ASIG5V.n10495 4.5005
R39551 ASIG5V.n10524 ASIG5V.n10494 4.5005
R39552 ASIG5V.n10911 ASIG5V.n10614 4.5005
R39553 ASIG5V.n10614 ASIG5V.n10495 4.5005
R39554 ASIG5V.n10614 ASIG5V.n10494 4.5005
R39555 ASIG5V.n10911 ASIG5V.n10523 4.5005
R39556 ASIG5V.n10523 ASIG5V.n10495 4.5005
R39557 ASIG5V.n10523 ASIG5V.n10494 4.5005
R39558 ASIG5V.n10911 ASIG5V.n10617 4.5005
R39559 ASIG5V.n10617 ASIG5V.n10495 4.5005
R39560 ASIG5V.n10617 ASIG5V.n10494 4.5005
R39561 ASIG5V.n10911 ASIG5V.n10522 4.5005
R39562 ASIG5V.n10522 ASIG5V.n10495 4.5005
R39563 ASIG5V.n10522 ASIG5V.n10494 4.5005
R39564 ASIG5V.n10911 ASIG5V.n10620 4.5005
R39565 ASIG5V.n10620 ASIG5V.n10495 4.5005
R39566 ASIG5V.n10620 ASIG5V.n10494 4.5005
R39567 ASIG5V.n10911 ASIG5V.n10521 4.5005
R39568 ASIG5V.n10521 ASIG5V.n10495 4.5005
R39569 ASIG5V.n10521 ASIG5V.n10494 4.5005
R39570 ASIG5V.n10911 ASIG5V.n10623 4.5005
R39571 ASIG5V.n10623 ASIG5V.n10495 4.5005
R39572 ASIG5V.n10623 ASIG5V.n10494 4.5005
R39573 ASIG5V.n10911 ASIG5V.n10520 4.5005
R39574 ASIG5V.n10520 ASIG5V.n10495 4.5005
R39575 ASIG5V.n10520 ASIG5V.n10494 4.5005
R39576 ASIG5V.n10911 ASIG5V.n10626 4.5005
R39577 ASIG5V.n10626 ASIG5V.n10495 4.5005
R39578 ASIG5V.n10626 ASIG5V.n10494 4.5005
R39579 ASIG5V.n10911 ASIG5V.n10519 4.5005
R39580 ASIG5V.n10519 ASIG5V.n10495 4.5005
R39581 ASIG5V.n10519 ASIG5V.n10494 4.5005
R39582 ASIG5V.n10911 ASIG5V.n10629 4.5005
R39583 ASIG5V.n10629 ASIG5V.n10495 4.5005
R39584 ASIG5V.n10629 ASIG5V.n10494 4.5005
R39585 ASIG5V.n10911 ASIG5V.n10518 4.5005
R39586 ASIG5V.n10518 ASIG5V.n10495 4.5005
R39587 ASIG5V.n10518 ASIG5V.n10494 4.5005
R39588 ASIG5V.n10911 ASIG5V.n10632 4.5005
R39589 ASIG5V.n10632 ASIG5V.n10495 4.5005
R39590 ASIG5V.n10632 ASIG5V.n10494 4.5005
R39591 ASIG5V.n10911 ASIG5V.n10517 4.5005
R39592 ASIG5V.n10517 ASIG5V.n10495 4.5005
R39593 ASIG5V.n10517 ASIG5V.n10494 4.5005
R39594 ASIG5V.n10911 ASIG5V.n10635 4.5005
R39595 ASIG5V.n10635 ASIG5V.n10495 4.5005
R39596 ASIG5V.n10635 ASIG5V.n10494 4.5005
R39597 ASIG5V.n10911 ASIG5V.n10516 4.5005
R39598 ASIG5V.n10516 ASIG5V.n10495 4.5005
R39599 ASIG5V.n10516 ASIG5V.n10494 4.5005
R39600 ASIG5V.n10911 ASIG5V.n10638 4.5005
R39601 ASIG5V.n10638 ASIG5V.n10495 4.5005
R39602 ASIG5V.n10638 ASIG5V.n10494 4.5005
R39603 ASIG5V.n10911 ASIG5V.n10515 4.5005
R39604 ASIG5V.n10515 ASIG5V.n10495 4.5005
R39605 ASIG5V.n10515 ASIG5V.n10494 4.5005
R39606 ASIG5V.n10911 ASIG5V.n10641 4.5005
R39607 ASIG5V.n10641 ASIG5V.n10495 4.5005
R39608 ASIG5V.n10641 ASIG5V.n10494 4.5005
R39609 ASIG5V.n10911 ASIG5V.n10514 4.5005
R39610 ASIG5V.n10514 ASIG5V.n10495 4.5005
R39611 ASIG5V.n10514 ASIG5V.n10494 4.5005
R39612 ASIG5V.n10911 ASIG5V.n10644 4.5005
R39613 ASIG5V.n10644 ASIG5V.n10495 4.5005
R39614 ASIG5V.n10644 ASIG5V.n10494 4.5005
R39615 ASIG5V.n10911 ASIG5V.n10513 4.5005
R39616 ASIG5V.n10513 ASIG5V.n10495 4.5005
R39617 ASIG5V.n10513 ASIG5V.n10494 4.5005
R39618 ASIG5V.n10911 ASIG5V.n10647 4.5005
R39619 ASIG5V.n10647 ASIG5V.n10495 4.5005
R39620 ASIG5V.n10647 ASIG5V.n10494 4.5005
R39621 ASIG5V.n10911 ASIG5V.n10512 4.5005
R39622 ASIG5V.n10512 ASIG5V.n10495 4.5005
R39623 ASIG5V.n10512 ASIG5V.n10494 4.5005
R39624 ASIG5V.n10911 ASIG5V.n10650 4.5005
R39625 ASIG5V.n10650 ASIG5V.n10495 4.5005
R39626 ASIG5V.n10650 ASIG5V.n10494 4.5005
R39627 ASIG5V.n10911 ASIG5V.n10511 4.5005
R39628 ASIG5V.n10511 ASIG5V.n10495 4.5005
R39629 ASIG5V.n10511 ASIG5V.n10494 4.5005
R39630 ASIG5V.n10911 ASIG5V.n10653 4.5005
R39631 ASIG5V.n10653 ASIG5V.n10495 4.5005
R39632 ASIG5V.n10653 ASIG5V.n10494 4.5005
R39633 ASIG5V.n10911 ASIG5V.n10510 4.5005
R39634 ASIG5V.n10510 ASIG5V.n10495 4.5005
R39635 ASIG5V.n10510 ASIG5V.n10494 4.5005
R39636 ASIG5V.n10911 ASIG5V.n10656 4.5005
R39637 ASIG5V.n10656 ASIG5V.n10495 4.5005
R39638 ASIG5V.n10656 ASIG5V.n10494 4.5005
R39639 ASIG5V.n10911 ASIG5V.n10509 4.5005
R39640 ASIG5V.n10509 ASIG5V.n10495 4.5005
R39641 ASIG5V.n10509 ASIG5V.n10494 4.5005
R39642 ASIG5V.n10911 ASIG5V.n10659 4.5005
R39643 ASIG5V.n10659 ASIG5V.n10495 4.5005
R39644 ASIG5V.n10659 ASIG5V.n10494 4.5005
R39645 ASIG5V.n10911 ASIG5V.n10508 4.5005
R39646 ASIG5V.n10508 ASIG5V.n10495 4.5005
R39647 ASIG5V.n10508 ASIG5V.n10494 4.5005
R39648 ASIG5V.n10911 ASIG5V.n10662 4.5005
R39649 ASIG5V.n10662 ASIG5V.n10495 4.5005
R39650 ASIG5V.n10662 ASIG5V.n10494 4.5005
R39651 ASIG5V.n10911 ASIG5V.n10507 4.5005
R39652 ASIG5V.n10507 ASIG5V.n10495 4.5005
R39653 ASIG5V.n10507 ASIG5V.n10494 4.5005
R39654 ASIG5V.n10911 ASIG5V.n10665 4.5005
R39655 ASIG5V.n10665 ASIG5V.n10495 4.5005
R39656 ASIG5V.n10665 ASIG5V.n10494 4.5005
R39657 ASIG5V.n10911 ASIG5V.n10506 4.5005
R39658 ASIG5V.n10506 ASIG5V.n10495 4.5005
R39659 ASIG5V.n10506 ASIG5V.n10494 4.5005
R39660 ASIG5V.n10911 ASIG5V.n10668 4.5005
R39661 ASIG5V.n10668 ASIG5V.n10495 4.5005
R39662 ASIG5V.n10668 ASIG5V.n10494 4.5005
R39663 ASIG5V.n10911 ASIG5V.n10505 4.5005
R39664 ASIG5V.n10505 ASIG5V.n10495 4.5005
R39665 ASIG5V.n10505 ASIG5V.n10494 4.5005
R39666 ASIG5V.n10911 ASIG5V.n10671 4.5005
R39667 ASIG5V.n10671 ASIG5V.n10495 4.5005
R39668 ASIG5V.n10671 ASIG5V.n10494 4.5005
R39669 ASIG5V.n10911 ASIG5V.n10504 4.5005
R39670 ASIG5V.n10504 ASIG5V.n10495 4.5005
R39671 ASIG5V.n10504 ASIG5V.n10494 4.5005
R39672 ASIG5V.n10911 ASIG5V.n10674 4.5005
R39673 ASIG5V.n10674 ASIG5V.n10495 4.5005
R39674 ASIG5V.n10674 ASIG5V.n10494 4.5005
R39675 ASIG5V.n10911 ASIG5V.n10503 4.5005
R39676 ASIG5V.n10503 ASIG5V.n10495 4.5005
R39677 ASIG5V.n10503 ASIG5V.n10494 4.5005
R39678 ASIG5V.n10911 ASIG5V.n10677 4.5005
R39679 ASIG5V.n10677 ASIG5V.n10495 4.5005
R39680 ASIG5V.n10677 ASIG5V.n10494 4.5005
R39681 ASIG5V.n10911 ASIG5V.n10502 4.5005
R39682 ASIG5V.n10502 ASIG5V.n10495 4.5005
R39683 ASIG5V.n10502 ASIG5V.n10494 4.5005
R39684 ASIG5V.n10911 ASIG5V.n10680 4.5005
R39685 ASIG5V.n10680 ASIG5V.n10495 4.5005
R39686 ASIG5V.n10680 ASIG5V.n10494 4.5005
R39687 ASIG5V.n10911 ASIG5V.n10501 4.5005
R39688 ASIG5V.n10501 ASIG5V.n10495 4.5005
R39689 ASIG5V.n10501 ASIG5V.n10494 4.5005
R39690 ASIG5V.n10911 ASIG5V.n10683 4.5005
R39691 ASIG5V.n10683 ASIG5V.n10495 4.5005
R39692 ASIG5V.n10683 ASIG5V.n10494 4.5005
R39693 ASIG5V.n10911 ASIG5V.n10500 4.5005
R39694 ASIG5V.n10500 ASIG5V.n10495 4.5005
R39695 ASIG5V.n10500 ASIG5V.n10494 4.5005
R39696 ASIG5V.n10911 ASIG5V.n10686 4.5005
R39697 ASIG5V.n10686 ASIG5V.n10495 4.5005
R39698 ASIG5V.n10686 ASIG5V.n10494 4.5005
R39699 ASIG5V.n10911 ASIG5V.n10499 4.5005
R39700 ASIG5V.n10499 ASIG5V.n10495 4.5005
R39701 ASIG5V.n10499 ASIG5V.n10494 4.5005
R39702 ASIG5V.n10911 ASIG5V.n10689 4.5005
R39703 ASIG5V.n10689 ASIG5V.n10495 4.5005
R39704 ASIG5V.n10689 ASIG5V.n10494 4.5005
R39705 ASIG5V.n10911 ASIG5V.n10498 4.5005
R39706 ASIG5V.n10498 ASIG5V.n10495 4.5005
R39707 ASIG5V.n10498 ASIG5V.n10494 4.5005
R39708 ASIG5V.n10911 ASIG5V.n10910 4.5005
R39709 ASIG5V.n10910 ASIG5V.n10495 4.5005
R39710 ASIG5V.n10910 ASIG5V.n10494 4.5005
R39711 ASIG5V.n10911 ASIG5V.n10497 4.5005
R39712 ASIG5V.n10497 ASIG5V.n10495 4.5005
R39713 ASIG5V.n10497 ASIG5V.n10493 4.5005
R39714 ASIG5V.n10497 ASIG5V.n10494 4.5005
R39715 ASIG5V.n4257 ASIG5V.n3848 4.5005
R39716 ASIG5V.n4257 ASIG5V.n3849 4.5005
R39717 ASIG5V.n4257 ASIG5V.n3847 4.5005
R39718 ASIG5V.n4257 ASIG5V.n3850 4.5005
R39719 ASIG5V.n4260 ASIG5V.n4257 4.5005
R39720 ASIG5V.n10713 ASIG5V.n10546 4.5005
R39721 ASIG5V.n10713 ASIG5V.n10697 4.5005
R39722 ASIG5V.n10713 ASIG5V.n10712 4.5005
R39723 ASIG5V.n4261 ASIG5V.n3848 4.5005
R39724 ASIG5V.n4261 ASIG5V.n3849 4.5005
R39725 ASIG5V.n4261 ASIG5V.n3847 4.5005
R39726 ASIG5V.n4261 ASIG5V.n3850 4.5005
R39727 ASIG5V.n4261 ASIG5V.n4260 4.5005
R39728 ASIG5V.n10704 ASIG5V.n10700 4.5005
R39729 ASIG5V.n10700 ASIG5V.n10496 4.5005
R39730 ASIG5V.n10700 ASIG5V.n10546 4.5005
R39731 ASIG5V.n10700 ASIG5V.n10697 4.5005
R39732 ASIG5V.n10712 ASIG5V.n10700 4.5005
R39733 ASIG5V.n3853 ASIG5V.n3848 4.5005
R39734 ASIG5V.n3853 ASIG5V.n3849 4.5005
R39735 ASIG5V.n3853 ASIG5V.n3847 4.5005
R39736 ASIG5V.n3853 ASIG5V.n3850 4.5005
R39737 ASIG5V.n4260 ASIG5V.n3853 4.5005
R39738 ASIG5V.n10704 ASIG5V.n10698 4.5005
R39739 ASIG5V.n10698 ASIG5V.n10496 4.5005
R39740 ASIG5V.n10698 ASIG5V.n10546 4.5005
R39741 ASIG5V.n10698 ASIG5V.n10697 4.5005
R39742 ASIG5V.n10712 ASIG5V.n10698 4.5005
R39743 ASIG5V.n4259 ASIG5V.n3848 4.5005
R39744 ASIG5V.n4259 ASIG5V.n3849 4.5005
R39745 ASIG5V.n4259 ASIG5V.n3847 4.5005
R39746 ASIG5V.n4259 ASIG5V.n3850 4.5005
R39747 ASIG5V.n4260 ASIG5V.n4259 4.5005
R39748 ASIG5V.n10711 ASIG5V.n10704 4.5005
R39749 ASIG5V.n10711 ASIG5V.n10496 4.5005
R39750 ASIG5V.n10711 ASIG5V.n10546 4.5005
R39751 ASIG5V.n10711 ASIG5V.n10697 4.5005
R39752 ASIG5V.n10712 ASIG5V.n10711 4.5005
R39753 ASIG5V.n11183 ASIG5V.n10067 4.5005
R39754 ASIG5V.n11183 ASIG5V.n11182 4.5005
R39755 ASIG5V.n11485 ASIG5V.n10015 4.5005
R39756 ASIG5V.n11485 ASIG5V.n11484 4.5005
R39757 ASIG5V.n11751 ASIG5V.n2955 4.5005
R39758 ASIG5V.n11751 ASIG5V.n11750 4.5005
R39759 ASIG5V.n11771 ASIG5V.n2611 4.5005
R39760 ASIG5V.n11771 ASIG5V.n11770 4.5005
R39761 ASIG5V.n2555 ASIG5V.n2263 4.5005
R39762 ASIG5V.n2555 ASIG5V.n2554 4.5005
R39763 ASIG5V.n2198 ASIG5V.n1906 4.5005
R39764 ASIG5V.n2198 ASIG5V.n2197 4.5005
R39765 ASIG5V.n11995 ASIG5V.n11994 4.5005
R39766 ASIG5V.n11994 ASIG5V.n11993 4.5005
R39767 ASIG5V.n12009 ASIG5V.n12008 4.5005
R39768 ASIG5V.n12008 ASIG5V.n12007 4.5005
R39769 ASIG5V.n12268 ASIG5V.n1268 4.5005
R39770 ASIG5V.n12268 ASIG5V.n12267 4.5005
R39771 ASIG5V.n967 ASIG5V.n877 4.5005
R39772 ASIG5V.n1214 ASIG5V.n877 4.5005
R39773 ASIG5V.n12301 ASIG5V.n570 4.5005
R39774 ASIG5V.n12301 ASIG5V.n12300 4.5005
R39775 ASIG5V.n12323 ASIG5V.n215 4.5005
R39776 ASIG5V.n12323 ASIG5V.n12322 4.5005
R39777 ASIG5V.n12526 ASIG5V.n12525 4.5005
R39778 ASIG5V.n12525 ASIG5V.n12524 4.5005
R39779 ASIG5V.n8879 ASIG5V.n1 4.5005
R39780 ASIG5V.n8632 ASIG5V.n1 4.5005
R39781 ASIG5V.n8893 ASIG5V.n8892 4.5005
R39782 ASIG5V.n8892 ASIG5V.n8891 4.5005
R39783 ASIG5V.n7229 ASIG5V.n6892 4.5005
R39784 ASIG5V.n7020 ASIG5V.n6892 4.5005
R39785 ASIG5V.n8917 ASIG5V.n8916 4.5005
R39786 ASIG5V.n8916 ASIG5V.n8915 4.5005
R39787 ASIG5V.n9176 ASIG5V.n6487 4.5005
R39788 ASIG5V.n9176 ASIG5V.n9175 4.5005
R39789 ASIG5V.n9380 ASIG5V.n9379 4.5005
R39790 ASIG5V.n9379 ASIG5V.n9378 4.5005
R39791 ASIG5V.n9394 ASIG5V.n9393 4.5005
R39792 ASIG5V.n9393 ASIG5V.n9392 4.5005
R39793 ASIG5V.n5905 ASIG5V.n5568 4.5005
R39794 ASIG5V.n5696 ASIG5V.n5568 4.5005
R39795 ASIG5V.n9417 ASIG5V.n9416 4.5005
R39796 ASIG5V.n9416 ASIG5V.n9415 4.5005
R39797 ASIG5V.n9432 ASIG5V.n5165 4.5005
R39798 ASIG5V.n9432 ASIG5V.n9431 4.5005
R39799 ASIG5V.n9734 ASIG5V.n5116 4.5005
R39800 ASIG5V.n9734 ASIG5V.n9733 4.5005
R39801 ASIG5V.n5064 ASIG5V.n3220 4.5005
R39802 ASIG5V.n5064 ASIG5V.n5063 4.5005
R39803 ASIG5V.n3614 ASIG5V.n3278 4.5005
R39804 ASIG5V.n3405 ASIG5V.n3278 4.5005
R39805 ASIG5V.n4256 ASIG5V.n3857 4.5005
R39806 ASIG5V.n4256 ASIG5V.n3855 4.5005
R39807 ASIG5V.n4256 ASIG5V.n3858 4.5005
R39808 ASIG5V.n4256 ASIG5V.n4255 4.5005
R39809 ASIG5V.n3906 ASIG5V.n3857 4.5005
R39810 ASIG5V.n3906 ASIG5V.n3858 4.5005
R39811 ASIG5V.n4255 ASIG5V.n3906 4.5005
R39812 ASIG5V.n3911 ASIG5V.n3857 4.5005
R39813 ASIG5V.n3911 ASIG5V.n3858 4.5005
R39814 ASIG5V.n4255 ASIG5V.n3911 4.5005
R39815 ASIG5V.n3905 ASIG5V.n3857 4.5005
R39816 ASIG5V.n3905 ASIG5V.n3858 4.5005
R39817 ASIG5V.n4255 ASIG5V.n3905 4.5005
R39818 ASIG5V.n3913 ASIG5V.n3857 4.5005
R39819 ASIG5V.n3913 ASIG5V.n3858 4.5005
R39820 ASIG5V.n4255 ASIG5V.n3913 4.5005
R39821 ASIG5V.n3904 ASIG5V.n3857 4.5005
R39822 ASIG5V.n3904 ASIG5V.n3858 4.5005
R39823 ASIG5V.n4255 ASIG5V.n3904 4.5005
R39824 ASIG5V.n3915 ASIG5V.n3857 4.5005
R39825 ASIG5V.n3915 ASIG5V.n3858 4.5005
R39826 ASIG5V.n4255 ASIG5V.n3915 4.5005
R39827 ASIG5V.n3903 ASIG5V.n3857 4.5005
R39828 ASIG5V.n3903 ASIG5V.n3858 4.5005
R39829 ASIG5V.n4255 ASIG5V.n3903 4.5005
R39830 ASIG5V.n3917 ASIG5V.n3857 4.5005
R39831 ASIG5V.n3917 ASIG5V.n3858 4.5005
R39832 ASIG5V.n4255 ASIG5V.n3917 4.5005
R39833 ASIG5V.n3902 ASIG5V.n3857 4.5005
R39834 ASIG5V.n3902 ASIG5V.n3858 4.5005
R39835 ASIG5V.n4255 ASIG5V.n3902 4.5005
R39836 ASIG5V.n3919 ASIG5V.n3857 4.5005
R39837 ASIG5V.n3919 ASIG5V.n3858 4.5005
R39838 ASIG5V.n4255 ASIG5V.n3919 4.5005
R39839 ASIG5V.n3901 ASIG5V.n3857 4.5005
R39840 ASIG5V.n3901 ASIG5V.n3858 4.5005
R39841 ASIG5V.n4255 ASIG5V.n3901 4.5005
R39842 ASIG5V.n3921 ASIG5V.n3857 4.5005
R39843 ASIG5V.n3921 ASIG5V.n3858 4.5005
R39844 ASIG5V.n4255 ASIG5V.n3921 4.5005
R39845 ASIG5V.n3900 ASIG5V.n3857 4.5005
R39846 ASIG5V.n3900 ASIG5V.n3858 4.5005
R39847 ASIG5V.n4255 ASIG5V.n3900 4.5005
R39848 ASIG5V.n3923 ASIG5V.n3857 4.5005
R39849 ASIG5V.n3923 ASIG5V.n3858 4.5005
R39850 ASIG5V.n4255 ASIG5V.n3923 4.5005
R39851 ASIG5V.n3899 ASIG5V.n3857 4.5005
R39852 ASIG5V.n3899 ASIG5V.n3858 4.5005
R39853 ASIG5V.n4255 ASIG5V.n3899 4.5005
R39854 ASIG5V.n3925 ASIG5V.n3857 4.5005
R39855 ASIG5V.n3925 ASIG5V.n3858 4.5005
R39856 ASIG5V.n4255 ASIG5V.n3925 4.5005
R39857 ASIG5V.n3898 ASIG5V.n3857 4.5005
R39858 ASIG5V.n3898 ASIG5V.n3858 4.5005
R39859 ASIG5V.n4255 ASIG5V.n3898 4.5005
R39860 ASIG5V.n3927 ASIG5V.n3857 4.5005
R39861 ASIG5V.n3927 ASIG5V.n3858 4.5005
R39862 ASIG5V.n4255 ASIG5V.n3927 4.5005
R39863 ASIG5V.n3897 ASIG5V.n3857 4.5005
R39864 ASIG5V.n3897 ASIG5V.n3858 4.5005
R39865 ASIG5V.n4255 ASIG5V.n3897 4.5005
R39866 ASIG5V.n3929 ASIG5V.n3857 4.5005
R39867 ASIG5V.n3929 ASIG5V.n3858 4.5005
R39868 ASIG5V.n4255 ASIG5V.n3929 4.5005
R39869 ASIG5V.n3896 ASIG5V.n3857 4.5005
R39870 ASIG5V.n3896 ASIG5V.n3858 4.5005
R39871 ASIG5V.n4255 ASIG5V.n3896 4.5005
R39872 ASIG5V.n3931 ASIG5V.n3857 4.5005
R39873 ASIG5V.n3931 ASIG5V.n3858 4.5005
R39874 ASIG5V.n4255 ASIG5V.n3931 4.5005
R39875 ASIG5V.n3895 ASIG5V.n3857 4.5005
R39876 ASIG5V.n3895 ASIG5V.n3858 4.5005
R39877 ASIG5V.n4255 ASIG5V.n3895 4.5005
R39878 ASIG5V.n3933 ASIG5V.n3857 4.5005
R39879 ASIG5V.n3933 ASIG5V.n3858 4.5005
R39880 ASIG5V.n4255 ASIG5V.n3933 4.5005
R39881 ASIG5V.n3894 ASIG5V.n3857 4.5005
R39882 ASIG5V.n3894 ASIG5V.n3858 4.5005
R39883 ASIG5V.n4255 ASIG5V.n3894 4.5005
R39884 ASIG5V.n3935 ASIG5V.n3857 4.5005
R39885 ASIG5V.n3935 ASIG5V.n3858 4.5005
R39886 ASIG5V.n4255 ASIG5V.n3935 4.5005
R39887 ASIG5V.n3893 ASIG5V.n3857 4.5005
R39888 ASIG5V.n3893 ASIG5V.n3858 4.5005
R39889 ASIG5V.n4255 ASIG5V.n3893 4.5005
R39890 ASIG5V.n3937 ASIG5V.n3857 4.5005
R39891 ASIG5V.n3937 ASIG5V.n3858 4.5005
R39892 ASIG5V.n4255 ASIG5V.n3937 4.5005
R39893 ASIG5V.n3892 ASIG5V.n3857 4.5005
R39894 ASIG5V.n3892 ASIG5V.n3858 4.5005
R39895 ASIG5V.n4255 ASIG5V.n3892 4.5005
R39896 ASIG5V.n3939 ASIG5V.n3857 4.5005
R39897 ASIG5V.n3939 ASIG5V.n3858 4.5005
R39898 ASIG5V.n4255 ASIG5V.n3939 4.5005
R39899 ASIG5V.n3891 ASIG5V.n3857 4.5005
R39900 ASIG5V.n3891 ASIG5V.n3858 4.5005
R39901 ASIG5V.n4255 ASIG5V.n3891 4.5005
R39902 ASIG5V.n3941 ASIG5V.n3857 4.5005
R39903 ASIG5V.n3941 ASIG5V.n3858 4.5005
R39904 ASIG5V.n4255 ASIG5V.n3941 4.5005
R39905 ASIG5V.n3890 ASIG5V.n3857 4.5005
R39906 ASIG5V.n3890 ASIG5V.n3858 4.5005
R39907 ASIG5V.n4255 ASIG5V.n3890 4.5005
R39908 ASIG5V.n3943 ASIG5V.n3857 4.5005
R39909 ASIG5V.n3943 ASIG5V.n3858 4.5005
R39910 ASIG5V.n4255 ASIG5V.n3943 4.5005
R39911 ASIG5V.n3889 ASIG5V.n3857 4.5005
R39912 ASIG5V.n3889 ASIG5V.n3858 4.5005
R39913 ASIG5V.n4255 ASIG5V.n3889 4.5005
R39914 ASIG5V.n3945 ASIG5V.n3857 4.5005
R39915 ASIG5V.n3945 ASIG5V.n3858 4.5005
R39916 ASIG5V.n4255 ASIG5V.n3945 4.5005
R39917 ASIG5V.n3888 ASIG5V.n3857 4.5005
R39918 ASIG5V.n3888 ASIG5V.n3858 4.5005
R39919 ASIG5V.n4255 ASIG5V.n3888 4.5005
R39920 ASIG5V.n3947 ASIG5V.n3857 4.5005
R39921 ASIG5V.n3947 ASIG5V.n3858 4.5005
R39922 ASIG5V.n4255 ASIG5V.n3947 4.5005
R39923 ASIG5V.n3887 ASIG5V.n3857 4.5005
R39924 ASIG5V.n3887 ASIG5V.n3858 4.5005
R39925 ASIG5V.n4255 ASIG5V.n3887 4.5005
R39926 ASIG5V.n3949 ASIG5V.n3857 4.5005
R39927 ASIG5V.n3949 ASIG5V.n3858 4.5005
R39928 ASIG5V.n4255 ASIG5V.n3949 4.5005
R39929 ASIG5V.n3886 ASIG5V.n3857 4.5005
R39930 ASIG5V.n3886 ASIG5V.n3858 4.5005
R39931 ASIG5V.n4255 ASIG5V.n3886 4.5005
R39932 ASIG5V.n3951 ASIG5V.n3857 4.5005
R39933 ASIG5V.n3951 ASIG5V.n3858 4.5005
R39934 ASIG5V.n4255 ASIG5V.n3951 4.5005
R39935 ASIG5V.n3885 ASIG5V.n3857 4.5005
R39936 ASIG5V.n3885 ASIG5V.n3858 4.5005
R39937 ASIG5V.n4255 ASIG5V.n3885 4.5005
R39938 ASIG5V.n3953 ASIG5V.n3857 4.5005
R39939 ASIG5V.n3953 ASIG5V.n3858 4.5005
R39940 ASIG5V.n4255 ASIG5V.n3953 4.5005
R39941 ASIG5V.n3884 ASIG5V.n3857 4.5005
R39942 ASIG5V.n3884 ASIG5V.n3858 4.5005
R39943 ASIG5V.n4255 ASIG5V.n3884 4.5005
R39944 ASIG5V.n3955 ASIG5V.n3857 4.5005
R39945 ASIG5V.n3955 ASIG5V.n3858 4.5005
R39946 ASIG5V.n4255 ASIG5V.n3955 4.5005
R39947 ASIG5V.n3883 ASIG5V.n3857 4.5005
R39948 ASIG5V.n3883 ASIG5V.n3858 4.5005
R39949 ASIG5V.n4255 ASIG5V.n3883 4.5005
R39950 ASIG5V.n3957 ASIG5V.n3857 4.5005
R39951 ASIG5V.n3957 ASIG5V.n3858 4.5005
R39952 ASIG5V.n4255 ASIG5V.n3957 4.5005
R39953 ASIG5V.n3882 ASIG5V.n3857 4.5005
R39954 ASIG5V.n3882 ASIG5V.n3858 4.5005
R39955 ASIG5V.n4255 ASIG5V.n3882 4.5005
R39956 ASIG5V.n3959 ASIG5V.n3857 4.5005
R39957 ASIG5V.n3959 ASIG5V.n3858 4.5005
R39958 ASIG5V.n4255 ASIG5V.n3959 4.5005
R39959 ASIG5V.n3881 ASIG5V.n3857 4.5005
R39960 ASIG5V.n3881 ASIG5V.n3858 4.5005
R39961 ASIG5V.n4255 ASIG5V.n3881 4.5005
R39962 ASIG5V.n3961 ASIG5V.n3857 4.5005
R39963 ASIG5V.n3961 ASIG5V.n3858 4.5005
R39964 ASIG5V.n4255 ASIG5V.n3961 4.5005
R39965 ASIG5V.n3880 ASIG5V.n3857 4.5005
R39966 ASIG5V.n3880 ASIG5V.n3858 4.5005
R39967 ASIG5V.n4255 ASIG5V.n3880 4.5005
R39968 ASIG5V.n3963 ASIG5V.n3857 4.5005
R39969 ASIG5V.n3963 ASIG5V.n3858 4.5005
R39970 ASIG5V.n4255 ASIG5V.n3963 4.5005
R39971 ASIG5V.n3879 ASIG5V.n3857 4.5005
R39972 ASIG5V.n3879 ASIG5V.n3858 4.5005
R39973 ASIG5V.n4255 ASIG5V.n3879 4.5005
R39974 ASIG5V.n3965 ASIG5V.n3857 4.5005
R39975 ASIG5V.n3965 ASIG5V.n3858 4.5005
R39976 ASIG5V.n4255 ASIG5V.n3965 4.5005
R39977 ASIG5V.n3878 ASIG5V.n3857 4.5005
R39978 ASIG5V.n3878 ASIG5V.n3858 4.5005
R39979 ASIG5V.n4255 ASIG5V.n3878 4.5005
R39980 ASIG5V.n3967 ASIG5V.n3857 4.5005
R39981 ASIG5V.n3967 ASIG5V.n3858 4.5005
R39982 ASIG5V.n4255 ASIG5V.n3967 4.5005
R39983 ASIG5V.n3877 ASIG5V.n3857 4.5005
R39984 ASIG5V.n3877 ASIG5V.n3858 4.5005
R39985 ASIG5V.n4255 ASIG5V.n3877 4.5005
R39986 ASIG5V.n3969 ASIG5V.n3857 4.5005
R39987 ASIG5V.n3969 ASIG5V.n3858 4.5005
R39988 ASIG5V.n4255 ASIG5V.n3969 4.5005
R39989 ASIG5V.n3876 ASIG5V.n3857 4.5005
R39990 ASIG5V.n3876 ASIG5V.n3858 4.5005
R39991 ASIG5V.n4255 ASIG5V.n3876 4.5005
R39992 ASIG5V.n3971 ASIG5V.n3857 4.5005
R39993 ASIG5V.n3971 ASIG5V.n3858 4.5005
R39994 ASIG5V.n4255 ASIG5V.n3971 4.5005
R39995 ASIG5V.n3875 ASIG5V.n3857 4.5005
R39996 ASIG5V.n3875 ASIG5V.n3858 4.5005
R39997 ASIG5V.n4255 ASIG5V.n3875 4.5005
R39998 ASIG5V.n3973 ASIG5V.n3857 4.5005
R39999 ASIG5V.n3973 ASIG5V.n3858 4.5005
R40000 ASIG5V.n4255 ASIG5V.n3973 4.5005
R40001 ASIG5V.n3874 ASIG5V.n3857 4.5005
R40002 ASIG5V.n3874 ASIG5V.n3858 4.5005
R40003 ASIG5V.n4255 ASIG5V.n3874 4.5005
R40004 ASIG5V.n3975 ASIG5V.n3857 4.5005
R40005 ASIG5V.n3975 ASIG5V.n3858 4.5005
R40006 ASIG5V.n4255 ASIG5V.n3975 4.5005
R40007 ASIG5V.n3873 ASIG5V.n3857 4.5005
R40008 ASIG5V.n3873 ASIG5V.n3858 4.5005
R40009 ASIG5V.n4255 ASIG5V.n3873 4.5005
R40010 ASIG5V.n3977 ASIG5V.n3857 4.5005
R40011 ASIG5V.n3977 ASIG5V.n3858 4.5005
R40012 ASIG5V.n4255 ASIG5V.n3977 4.5005
R40013 ASIG5V.n3872 ASIG5V.n3857 4.5005
R40014 ASIG5V.n3872 ASIG5V.n3858 4.5005
R40015 ASIG5V.n4255 ASIG5V.n3872 4.5005
R40016 ASIG5V.n3979 ASIG5V.n3857 4.5005
R40017 ASIG5V.n3979 ASIG5V.n3858 4.5005
R40018 ASIG5V.n4255 ASIG5V.n3979 4.5005
R40019 ASIG5V.n3871 ASIG5V.n3857 4.5005
R40020 ASIG5V.n3871 ASIG5V.n3858 4.5005
R40021 ASIG5V.n4255 ASIG5V.n3871 4.5005
R40022 ASIG5V.n3981 ASIG5V.n3857 4.5005
R40023 ASIG5V.n3981 ASIG5V.n3858 4.5005
R40024 ASIG5V.n4255 ASIG5V.n3981 4.5005
R40025 ASIG5V.n3870 ASIG5V.n3857 4.5005
R40026 ASIG5V.n3870 ASIG5V.n3858 4.5005
R40027 ASIG5V.n4255 ASIG5V.n3870 4.5005
R40028 ASIG5V.n3983 ASIG5V.n3857 4.5005
R40029 ASIG5V.n3983 ASIG5V.n3858 4.5005
R40030 ASIG5V.n4255 ASIG5V.n3983 4.5005
R40031 ASIG5V.n3869 ASIG5V.n3857 4.5005
R40032 ASIG5V.n3869 ASIG5V.n3858 4.5005
R40033 ASIG5V.n4255 ASIG5V.n3869 4.5005
R40034 ASIG5V.n3985 ASIG5V.n3857 4.5005
R40035 ASIG5V.n3985 ASIG5V.n3858 4.5005
R40036 ASIG5V.n4255 ASIG5V.n3985 4.5005
R40037 ASIG5V.n3868 ASIG5V.n3857 4.5005
R40038 ASIG5V.n3868 ASIG5V.n3858 4.5005
R40039 ASIG5V.n4255 ASIG5V.n3868 4.5005
R40040 ASIG5V.n3987 ASIG5V.n3857 4.5005
R40041 ASIG5V.n3987 ASIG5V.n3858 4.5005
R40042 ASIG5V.n4255 ASIG5V.n3987 4.5005
R40043 ASIG5V.n3867 ASIG5V.n3857 4.5005
R40044 ASIG5V.n3867 ASIG5V.n3858 4.5005
R40045 ASIG5V.n4255 ASIG5V.n3867 4.5005
R40046 ASIG5V.n3989 ASIG5V.n3857 4.5005
R40047 ASIG5V.n3989 ASIG5V.n3858 4.5005
R40048 ASIG5V.n4255 ASIG5V.n3989 4.5005
R40049 ASIG5V.n3866 ASIG5V.n3857 4.5005
R40050 ASIG5V.n3866 ASIG5V.n3858 4.5005
R40051 ASIG5V.n4255 ASIG5V.n3866 4.5005
R40052 ASIG5V.n3991 ASIG5V.n3857 4.5005
R40053 ASIG5V.n3991 ASIG5V.n3858 4.5005
R40054 ASIG5V.n4255 ASIG5V.n3991 4.5005
R40055 ASIG5V.n3865 ASIG5V.n3857 4.5005
R40056 ASIG5V.n3865 ASIG5V.n3858 4.5005
R40057 ASIG5V.n4255 ASIG5V.n3865 4.5005
R40058 ASIG5V.n3993 ASIG5V.n3857 4.5005
R40059 ASIG5V.n3993 ASIG5V.n3858 4.5005
R40060 ASIG5V.n4255 ASIG5V.n3993 4.5005
R40061 ASIG5V.n3864 ASIG5V.n3857 4.5005
R40062 ASIG5V.n3864 ASIG5V.n3858 4.5005
R40063 ASIG5V.n4255 ASIG5V.n3864 4.5005
R40064 ASIG5V.n3995 ASIG5V.n3857 4.5005
R40065 ASIG5V.n3995 ASIG5V.n3858 4.5005
R40066 ASIG5V.n4255 ASIG5V.n3995 4.5005
R40067 ASIG5V.n3863 ASIG5V.n3857 4.5005
R40068 ASIG5V.n3863 ASIG5V.n3858 4.5005
R40069 ASIG5V.n4255 ASIG5V.n3863 4.5005
R40070 ASIG5V.n3997 ASIG5V.n3857 4.5005
R40071 ASIG5V.n3997 ASIG5V.n3858 4.5005
R40072 ASIG5V.n4255 ASIG5V.n3997 4.5005
R40073 ASIG5V.n3862 ASIG5V.n3857 4.5005
R40074 ASIG5V.n3862 ASIG5V.n3858 4.5005
R40075 ASIG5V.n4255 ASIG5V.n3862 4.5005
R40076 ASIG5V.n3999 ASIG5V.n3857 4.5005
R40077 ASIG5V.n3999 ASIG5V.n3858 4.5005
R40078 ASIG5V.n4255 ASIG5V.n3999 4.5005
R40079 ASIG5V.n3861 ASIG5V.n3857 4.5005
R40080 ASIG5V.n3861 ASIG5V.n3858 4.5005
R40081 ASIG5V.n4255 ASIG5V.n3861 4.5005
R40082 ASIG5V.n4001 ASIG5V.n3857 4.5005
R40083 ASIG5V.n4001 ASIG5V.n3858 4.5005
R40084 ASIG5V.n4255 ASIG5V.n4001 4.5005
R40085 ASIG5V.n3860 ASIG5V.n3857 4.5005
R40086 ASIG5V.n3860 ASIG5V.n3858 4.5005
R40087 ASIG5V.n4255 ASIG5V.n3860 4.5005
R40088 ASIG5V.n4003 ASIG5V.n3857 4.5005
R40089 ASIG5V.n4003 ASIG5V.n3858 4.5005
R40090 ASIG5V.n4255 ASIG5V.n4003 4.5005
R40091 ASIG5V.n3859 ASIG5V.n3857 4.5005
R40092 ASIG5V.n3859 ASIG5V.n3858 4.5005
R40093 ASIG5V.n4255 ASIG5V.n3859 4.5005
R40094 ASIG5V.n4254 ASIG5V.n3857 4.5005
R40095 ASIG5V.n4254 ASIG5V.n3855 4.5005
R40096 ASIG5V.n4254 ASIG5V.n3858 4.5005
R40097 ASIG5V.n4255 ASIG5V.n4254 4.5005
R40098 ASIG5V.n10912 ASIG5V.n10494 4.5005
R40099 ASIG5V.n10912 ASIG5V.n10493 4.5005
R40100 ASIG5V.n10912 ASIG5V.n10495 4.5005
R40101 ASIG5V.n10912 ASIG5V.n10492 4.5005
R40102 ASIG5V.n10912 ASIG5V.n10911 4.5005
R40103 ASIG5V.n3909 ASIG5V.n3857 4.5005
R40104 ASIG5V.n4773 ASIG5V.n4772 4.5005
R40105 ASIG5V.n4772 ASIG5V.n4771 4.5005
R40106 ASIG5V.n11172 ASIG5V.n10415 4.5005
R40107 ASIG5V.n11172 ASIG5V.n11171 4.5005
R40108 ASIG5V.n4568 ASIG5V.n3829 4.5005
R40109 ASIG5V.n4568 ASIG5V.n4567 4.5005
R40110 ASIG5V.n7995 ASIG5V.n7994 4.5005
R40111 ASIG5V.n7985 ASIG5V.n7532 4.5005
R40112 ASIG5V.n7994 ASIG5V.n7532 4.5005
R40113 ASIG5V.n7992 ASIG5V.n7987 4.5005
R40114 ASIG5V.n7992 ASIG5V.n7991 4.5005
R40115 ASIG5V.n7991 ASIG5V.n7983 4.5005
R40116 ASIG5V.n8006 ASIG5V.n8005 4.5005
R40117 ASIG5V.n8000 ASIG5V.n7527 4.5005
R40118 ASIG5V.n8005 ASIG5V.n7527 4.5005
R40119 ASIG5V.n8003 ASIG5V.n8002 4.5005
R40120 ASIG5V.n8003 ASIG5V.n3153 4.5005
R40121 ASIG5V.n7996 ASIG5V.n3153 4.5005
R40122 ASIG5V.n8017 ASIG5V.n8016 4.5005
R40123 ASIG5V.n8011 ASIG5V.n7522 4.5005
R40124 ASIG5V.n8016 ASIG5V.n7522 4.5005
R40125 ASIG5V.n8014 ASIG5V.n8013 4.5005
R40126 ASIG5V.n8014 ASIG5V.n3147 4.5005
R40127 ASIG5V.n8007 ASIG5V.n3147 4.5005
R40128 ASIG5V.n8028 ASIG5V.n8027 4.5005
R40129 ASIG5V.n8022 ASIG5V.n7517 4.5005
R40130 ASIG5V.n8027 ASIG5V.n7517 4.5005
R40131 ASIG5V.n8025 ASIG5V.n8024 4.5005
R40132 ASIG5V.n8025 ASIG5V.n3142 4.5005
R40133 ASIG5V.n8018 ASIG5V.n3142 4.5005
R40134 ASIG5V.n8039 ASIG5V.n8038 4.5005
R40135 ASIG5V.n8033 ASIG5V.n7512 4.5005
R40136 ASIG5V.n8038 ASIG5V.n7512 4.5005
R40137 ASIG5V.n8036 ASIG5V.n8035 4.5005
R40138 ASIG5V.n8036 ASIG5V.n3137 4.5005
R40139 ASIG5V.n8029 ASIG5V.n3137 4.5005
R40140 ASIG5V.n8050 ASIG5V.n8049 4.5005
R40141 ASIG5V.n8044 ASIG5V.n7507 4.5005
R40142 ASIG5V.n8049 ASIG5V.n7507 4.5005
R40143 ASIG5V.n8047 ASIG5V.n8046 4.5005
R40144 ASIG5V.n8047 ASIG5V.n3132 4.5005
R40145 ASIG5V.n8040 ASIG5V.n3132 4.5005
R40146 ASIG5V.n8062 ASIG5V.n7503 4.5005
R40147 ASIG5V.n8056 ASIG5V.n7502 4.5005
R40148 ASIG5V.n8062 ASIG5V.n7502 4.5005
R40149 ASIG5V.n8060 ASIG5V.n8059 4.5005
R40150 ASIG5V.n8060 ASIG5V.n3127 4.5005
R40151 ASIG5V.n8051 ASIG5V.n3127 4.5005
R40152 ASIG5V.n9846 ASIG5V.n3115 4.5005
R40153 ASIG5V.n9839 ASIG5V.n3114 4.5005
R40154 ASIG5V.n9846 ASIG5V.n3114 4.5005
R40155 ASIG5V.n9844 ASIG5V.n3119 4.5005
R40156 ASIG5V.n9844 ASIG5V.n9843 4.5005
R40157 ASIG5V.n9843 ASIG5V.n3116 4.5005
R40158 ASIG5V.n10713 ASIG5V.n10696 2.25086
R40159 ASIG5V.n3407 ASIG5V.n3406 2.2505
R40160 ASIG5V.n3409 ASIG5V.n3408 2.2505
R40161 ASIG5V.n3401 ASIG5V.n3400 2.2505
R40162 ASIG5V.n3416 ASIG5V.n3415 2.2505
R40163 ASIG5V.n3417 ASIG5V.n3399 2.2505
R40164 ASIG5V.n3419 ASIG5V.n3418 2.2505
R40165 ASIG5V.n3395 ASIG5V.n3394 2.2505
R40166 ASIG5V.n3426 ASIG5V.n3425 2.2505
R40167 ASIG5V.n3427 ASIG5V.n3393 2.2505
R40168 ASIG5V.n3429 ASIG5V.n3428 2.2505
R40169 ASIG5V.n3389 ASIG5V.n3388 2.2505
R40170 ASIG5V.n3436 ASIG5V.n3435 2.2505
R40171 ASIG5V.n3437 ASIG5V.n3387 2.2505
R40172 ASIG5V.n3439 ASIG5V.n3438 2.2505
R40173 ASIG5V.n3383 ASIG5V.n3382 2.2505
R40174 ASIG5V.n3446 ASIG5V.n3445 2.2505
R40175 ASIG5V.n3447 ASIG5V.n3381 2.2505
R40176 ASIG5V.n3449 ASIG5V.n3448 2.2505
R40177 ASIG5V.n3377 ASIG5V.n3376 2.2505
R40178 ASIG5V.n3456 ASIG5V.n3455 2.2505
R40179 ASIG5V.n3457 ASIG5V.n3375 2.2505
R40180 ASIG5V.n3459 ASIG5V.n3458 2.2505
R40181 ASIG5V.n3371 ASIG5V.n3370 2.2505
R40182 ASIG5V.n3466 ASIG5V.n3465 2.2505
R40183 ASIG5V.n3467 ASIG5V.n3369 2.2505
R40184 ASIG5V.n3469 ASIG5V.n3468 2.2505
R40185 ASIG5V.n3365 ASIG5V.n3364 2.2505
R40186 ASIG5V.n3476 ASIG5V.n3475 2.2505
R40187 ASIG5V.n3477 ASIG5V.n3363 2.2505
R40188 ASIG5V.n3479 ASIG5V.n3478 2.2505
R40189 ASIG5V.n3359 ASIG5V.n3358 2.2505
R40190 ASIG5V.n3486 ASIG5V.n3485 2.2505
R40191 ASIG5V.n3487 ASIG5V.n3357 2.2505
R40192 ASIG5V.n3489 ASIG5V.n3488 2.2505
R40193 ASIG5V.n3353 ASIG5V.n3352 2.2505
R40194 ASIG5V.n3496 ASIG5V.n3495 2.2505
R40195 ASIG5V.n3497 ASIG5V.n3351 2.2505
R40196 ASIG5V.n3499 ASIG5V.n3498 2.2505
R40197 ASIG5V.n3347 ASIG5V.n3346 2.2505
R40198 ASIG5V.n3506 ASIG5V.n3505 2.2505
R40199 ASIG5V.n3507 ASIG5V.n3345 2.2505
R40200 ASIG5V.n3509 ASIG5V.n3508 2.2505
R40201 ASIG5V.n3341 ASIG5V.n3340 2.2505
R40202 ASIG5V.n3516 ASIG5V.n3515 2.2505
R40203 ASIG5V.n3517 ASIG5V.n3339 2.2505
R40204 ASIG5V.n3519 ASIG5V.n3518 2.2505
R40205 ASIG5V.n3335 ASIG5V.n3334 2.2505
R40206 ASIG5V.n3526 ASIG5V.n3525 2.2505
R40207 ASIG5V.n3527 ASIG5V.n3333 2.2505
R40208 ASIG5V.n3529 ASIG5V.n3528 2.2505
R40209 ASIG5V.n3329 ASIG5V.n3328 2.2505
R40210 ASIG5V.n3536 ASIG5V.n3535 2.2505
R40211 ASIG5V.n3537 ASIG5V.n3327 2.2505
R40212 ASIG5V.n3539 ASIG5V.n3538 2.2505
R40213 ASIG5V.n3323 ASIG5V.n3322 2.2505
R40214 ASIG5V.n3546 ASIG5V.n3545 2.2505
R40215 ASIG5V.n3547 ASIG5V.n3321 2.2505
R40216 ASIG5V.n3549 ASIG5V.n3548 2.2505
R40217 ASIG5V.n3317 ASIG5V.n3316 2.2505
R40218 ASIG5V.n3556 ASIG5V.n3555 2.2505
R40219 ASIG5V.n3557 ASIG5V.n3315 2.2505
R40220 ASIG5V.n3559 ASIG5V.n3558 2.2505
R40221 ASIG5V.n3311 ASIG5V.n3310 2.2505
R40222 ASIG5V.n3566 ASIG5V.n3565 2.2505
R40223 ASIG5V.n3567 ASIG5V.n3309 2.2505
R40224 ASIG5V.n3569 ASIG5V.n3568 2.2505
R40225 ASIG5V.n3305 ASIG5V.n3304 2.2505
R40226 ASIG5V.n3576 ASIG5V.n3575 2.2505
R40227 ASIG5V.n3577 ASIG5V.n3303 2.2505
R40228 ASIG5V.n3579 ASIG5V.n3578 2.2505
R40229 ASIG5V.n3299 ASIG5V.n3298 2.2505
R40230 ASIG5V.n3586 ASIG5V.n3585 2.2505
R40231 ASIG5V.n3587 ASIG5V.n3297 2.2505
R40232 ASIG5V.n3589 ASIG5V.n3588 2.2505
R40233 ASIG5V.n3293 ASIG5V.n3292 2.2505
R40234 ASIG5V.n3596 ASIG5V.n3595 2.2505
R40235 ASIG5V.n3597 ASIG5V.n3291 2.2505
R40236 ASIG5V.n3599 ASIG5V.n3598 2.2505
R40237 ASIG5V.n3287 ASIG5V.n3286 2.2505
R40238 ASIG5V.n3606 ASIG5V.n3605 2.2505
R40239 ASIG5V.n3607 ASIG5V.n3285 2.2505
R40240 ASIG5V.n3609 ASIG5V.n3608 2.2505
R40241 ASIG5V.n3283 ASIG5V.n3282 2.2505
R40242 ASIG5V.n3616 ASIG5V.n3615 2.2505
R40243 ASIG5V.n3615 ASIG5V.n3614 2.2505
R40244 ASIG5V.n3612 ASIG5V.n3283 2.2505
R40245 ASIG5V.n3610 ASIG5V.n3609 2.2505
R40246 ASIG5V.n3288 ASIG5V.n3285 2.2505
R40247 ASIG5V.n3605 ASIG5V.n3604 2.2505
R40248 ASIG5V.n3602 ASIG5V.n3287 2.2505
R40249 ASIG5V.n3600 ASIG5V.n3599 2.2505
R40250 ASIG5V.n3294 ASIG5V.n3291 2.2505
R40251 ASIG5V.n3595 ASIG5V.n3594 2.2505
R40252 ASIG5V.n3592 ASIG5V.n3293 2.2505
R40253 ASIG5V.n3590 ASIG5V.n3589 2.2505
R40254 ASIG5V.n3300 ASIG5V.n3297 2.2505
R40255 ASIG5V.n3585 ASIG5V.n3584 2.2505
R40256 ASIG5V.n3582 ASIG5V.n3299 2.2505
R40257 ASIG5V.n3580 ASIG5V.n3579 2.2505
R40258 ASIG5V.n3306 ASIG5V.n3303 2.2505
R40259 ASIG5V.n3575 ASIG5V.n3574 2.2505
R40260 ASIG5V.n3572 ASIG5V.n3305 2.2505
R40261 ASIG5V.n3570 ASIG5V.n3569 2.2505
R40262 ASIG5V.n3312 ASIG5V.n3309 2.2505
R40263 ASIG5V.n3565 ASIG5V.n3564 2.2505
R40264 ASIG5V.n3562 ASIG5V.n3311 2.2505
R40265 ASIG5V.n3560 ASIG5V.n3559 2.2505
R40266 ASIG5V.n3318 ASIG5V.n3315 2.2505
R40267 ASIG5V.n3555 ASIG5V.n3554 2.2505
R40268 ASIG5V.n3552 ASIG5V.n3317 2.2505
R40269 ASIG5V.n3550 ASIG5V.n3549 2.2505
R40270 ASIG5V.n3324 ASIG5V.n3321 2.2505
R40271 ASIG5V.n3545 ASIG5V.n3544 2.2505
R40272 ASIG5V.n3542 ASIG5V.n3323 2.2505
R40273 ASIG5V.n3540 ASIG5V.n3539 2.2505
R40274 ASIG5V.n3330 ASIG5V.n3327 2.2505
R40275 ASIG5V.n3535 ASIG5V.n3534 2.2505
R40276 ASIG5V.n3532 ASIG5V.n3329 2.2505
R40277 ASIG5V.n3530 ASIG5V.n3529 2.2505
R40278 ASIG5V.n3336 ASIG5V.n3333 2.2505
R40279 ASIG5V.n3525 ASIG5V.n3524 2.2505
R40280 ASIG5V.n3522 ASIG5V.n3335 2.2505
R40281 ASIG5V.n3520 ASIG5V.n3519 2.2505
R40282 ASIG5V.n3342 ASIG5V.n3339 2.2505
R40283 ASIG5V.n3515 ASIG5V.n3514 2.2505
R40284 ASIG5V.n3512 ASIG5V.n3341 2.2505
R40285 ASIG5V.n3510 ASIG5V.n3509 2.2505
R40286 ASIG5V.n3348 ASIG5V.n3345 2.2505
R40287 ASIG5V.n3505 ASIG5V.n3504 2.2505
R40288 ASIG5V.n3502 ASIG5V.n3347 2.2505
R40289 ASIG5V.n3500 ASIG5V.n3499 2.2505
R40290 ASIG5V.n3354 ASIG5V.n3351 2.2505
R40291 ASIG5V.n3495 ASIG5V.n3494 2.2505
R40292 ASIG5V.n3492 ASIG5V.n3353 2.2505
R40293 ASIG5V.n3490 ASIG5V.n3489 2.2505
R40294 ASIG5V.n3360 ASIG5V.n3357 2.2505
R40295 ASIG5V.n3485 ASIG5V.n3484 2.2505
R40296 ASIG5V.n3482 ASIG5V.n3359 2.2505
R40297 ASIG5V.n3480 ASIG5V.n3479 2.2505
R40298 ASIG5V.n3366 ASIG5V.n3363 2.2505
R40299 ASIG5V.n3475 ASIG5V.n3474 2.2505
R40300 ASIG5V.n3472 ASIG5V.n3365 2.2505
R40301 ASIG5V.n3470 ASIG5V.n3469 2.2505
R40302 ASIG5V.n3372 ASIG5V.n3369 2.2505
R40303 ASIG5V.n3465 ASIG5V.n3464 2.2505
R40304 ASIG5V.n3462 ASIG5V.n3371 2.2505
R40305 ASIG5V.n3460 ASIG5V.n3459 2.2505
R40306 ASIG5V.n3378 ASIG5V.n3375 2.2505
R40307 ASIG5V.n3455 ASIG5V.n3454 2.2505
R40308 ASIG5V.n3452 ASIG5V.n3377 2.2505
R40309 ASIG5V.n3450 ASIG5V.n3449 2.2505
R40310 ASIG5V.n3384 ASIG5V.n3381 2.2505
R40311 ASIG5V.n3445 ASIG5V.n3444 2.2505
R40312 ASIG5V.n3442 ASIG5V.n3383 2.2505
R40313 ASIG5V.n3440 ASIG5V.n3439 2.2505
R40314 ASIG5V.n3390 ASIG5V.n3387 2.2505
R40315 ASIG5V.n3435 ASIG5V.n3434 2.2505
R40316 ASIG5V.n3432 ASIG5V.n3389 2.2505
R40317 ASIG5V.n3430 ASIG5V.n3429 2.2505
R40318 ASIG5V.n3396 ASIG5V.n3393 2.2505
R40319 ASIG5V.n3425 ASIG5V.n3424 2.2505
R40320 ASIG5V.n3422 ASIG5V.n3395 2.2505
R40321 ASIG5V.n3420 ASIG5V.n3419 2.2505
R40322 ASIG5V.n3402 ASIG5V.n3399 2.2505
R40323 ASIG5V.n3415 ASIG5V.n3414 2.2505
R40324 ASIG5V.n3412 ASIG5V.n3401 2.2505
R40325 ASIG5V.n3410 ASIG5V.n3409 2.2505
R40326 ASIG5V.n3406 ASIG5V.n3405 2.2505
R40327 ASIG5V.n5058 ASIG5V.n3222 2.2505
R40328 ASIG5V.n5060 ASIG5V.n5059 2.2505
R40329 ASIG5V.n5057 ASIG5V.n3224 2.2505
R40330 ASIG5V.n5056 ASIG5V.n5055 2.2505
R40331 ASIG5V.n5051 ASIG5V.n3225 2.2505
R40332 ASIG5V.n5047 ASIG5V.n5046 2.2505
R40333 ASIG5V.n5045 ASIG5V.n3226 2.2505
R40334 ASIG5V.n5044 ASIG5V.n5043 2.2505
R40335 ASIG5V.n5039 ASIG5V.n3227 2.2505
R40336 ASIG5V.n5035 ASIG5V.n5034 2.2505
R40337 ASIG5V.n5033 ASIG5V.n3228 2.2505
R40338 ASIG5V.n5032 ASIG5V.n5031 2.2505
R40339 ASIG5V.n5027 ASIG5V.n3229 2.2505
R40340 ASIG5V.n5023 ASIG5V.n5022 2.2505
R40341 ASIG5V.n5021 ASIG5V.n3230 2.2505
R40342 ASIG5V.n5020 ASIG5V.n5019 2.2505
R40343 ASIG5V.n5015 ASIG5V.n3231 2.2505
R40344 ASIG5V.n5011 ASIG5V.n5010 2.2505
R40345 ASIG5V.n5009 ASIG5V.n3232 2.2505
R40346 ASIG5V.n5008 ASIG5V.n5007 2.2505
R40347 ASIG5V.n5003 ASIG5V.n3233 2.2505
R40348 ASIG5V.n4999 ASIG5V.n4998 2.2505
R40349 ASIG5V.n4997 ASIG5V.n3234 2.2505
R40350 ASIG5V.n4996 ASIG5V.n4995 2.2505
R40351 ASIG5V.n4991 ASIG5V.n3235 2.2505
R40352 ASIG5V.n4987 ASIG5V.n4986 2.2505
R40353 ASIG5V.n4985 ASIG5V.n3236 2.2505
R40354 ASIG5V.n4984 ASIG5V.n4983 2.2505
R40355 ASIG5V.n4979 ASIG5V.n3237 2.2505
R40356 ASIG5V.n4975 ASIG5V.n4974 2.2505
R40357 ASIG5V.n4973 ASIG5V.n3238 2.2505
R40358 ASIG5V.n4972 ASIG5V.n4971 2.2505
R40359 ASIG5V.n4967 ASIG5V.n3239 2.2505
R40360 ASIG5V.n4963 ASIG5V.n4962 2.2505
R40361 ASIG5V.n4961 ASIG5V.n3240 2.2505
R40362 ASIG5V.n4960 ASIG5V.n4959 2.2505
R40363 ASIG5V.n4955 ASIG5V.n3241 2.2505
R40364 ASIG5V.n4951 ASIG5V.n4950 2.2505
R40365 ASIG5V.n4949 ASIG5V.n3242 2.2505
R40366 ASIG5V.n4948 ASIG5V.n4947 2.2505
R40367 ASIG5V.n4943 ASIG5V.n3243 2.2505
R40368 ASIG5V.n4939 ASIG5V.n4938 2.2505
R40369 ASIG5V.n4937 ASIG5V.n3244 2.2505
R40370 ASIG5V.n4936 ASIG5V.n4935 2.2505
R40371 ASIG5V.n4931 ASIG5V.n3245 2.2505
R40372 ASIG5V.n4927 ASIG5V.n4926 2.2505
R40373 ASIG5V.n4925 ASIG5V.n3246 2.2505
R40374 ASIG5V.n4924 ASIG5V.n4923 2.2505
R40375 ASIG5V.n4919 ASIG5V.n3247 2.2505
R40376 ASIG5V.n4915 ASIG5V.n4914 2.2505
R40377 ASIG5V.n4913 ASIG5V.n3248 2.2505
R40378 ASIG5V.n4912 ASIG5V.n4911 2.2505
R40379 ASIG5V.n4907 ASIG5V.n3249 2.2505
R40380 ASIG5V.n4903 ASIG5V.n4902 2.2505
R40381 ASIG5V.n4901 ASIG5V.n3250 2.2505
R40382 ASIG5V.n4900 ASIG5V.n4899 2.2505
R40383 ASIG5V.n4895 ASIG5V.n3251 2.2505
R40384 ASIG5V.n4891 ASIG5V.n4890 2.2505
R40385 ASIG5V.n4889 ASIG5V.n3252 2.2505
R40386 ASIG5V.n4888 ASIG5V.n4887 2.2505
R40387 ASIG5V.n4883 ASIG5V.n3253 2.2505
R40388 ASIG5V.n4879 ASIG5V.n4878 2.2505
R40389 ASIG5V.n4877 ASIG5V.n3254 2.2505
R40390 ASIG5V.n4876 ASIG5V.n4875 2.2505
R40391 ASIG5V.n4871 ASIG5V.n3255 2.2505
R40392 ASIG5V.n4867 ASIG5V.n4866 2.2505
R40393 ASIG5V.n4865 ASIG5V.n3256 2.2505
R40394 ASIG5V.n4864 ASIG5V.n4863 2.2505
R40395 ASIG5V.n4859 ASIG5V.n3257 2.2505
R40396 ASIG5V.n4855 ASIG5V.n4854 2.2505
R40397 ASIG5V.n4853 ASIG5V.n3258 2.2505
R40398 ASIG5V.n4852 ASIG5V.n4851 2.2505
R40399 ASIG5V.n4847 ASIG5V.n3259 2.2505
R40400 ASIG5V.n4843 ASIG5V.n4842 2.2505
R40401 ASIG5V.n4841 ASIG5V.n3260 2.2505
R40402 ASIG5V.n4840 ASIG5V.n4839 2.2505
R40403 ASIG5V.n4835 ASIG5V.n3261 2.2505
R40404 ASIG5V.n4831 ASIG5V.n4830 2.2505
R40405 ASIG5V.n4829 ASIG5V.n3262 2.2505
R40406 ASIG5V.n4828 ASIG5V.n4827 2.2505
R40407 ASIG5V.n4823 ASIG5V.n3263 2.2505
R40408 ASIG5V.n4819 ASIG5V.n4818 2.2505
R40409 ASIG5V.n4817 ASIG5V.n3266 2.2505
R40410 ASIG5V.n4816 ASIG5V.n4815 2.2505
R40411 ASIG5V.n4815 ASIG5V.n3220 2.2505
R40412 ASIG5V.n3266 ASIG5V.n3265 2.2505
R40413 ASIG5V.n4820 ASIG5V.n4819 2.2505
R40414 ASIG5V.n4823 ASIG5V.n4822 2.2505
R40415 ASIG5V.n4827 ASIG5V.n4826 2.2505
R40416 ASIG5V.n4824 ASIG5V.n3262 2.2505
R40417 ASIG5V.n4832 ASIG5V.n4831 2.2505
R40418 ASIG5V.n4835 ASIG5V.n4834 2.2505
R40419 ASIG5V.n4839 ASIG5V.n4838 2.2505
R40420 ASIG5V.n4836 ASIG5V.n3260 2.2505
R40421 ASIG5V.n4844 ASIG5V.n4843 2.2505
R40422 ASIG5V.n4847 ASIG5V.n4846 2.2505
R40423 ASIG5V.n4851 ASIG5V.n4850 2.2505
R40424 ASIG5V.n4848 ASIG5V.n3258 2.2505
R40425 ASIG5V.n4856 ASIG5V.n4855 2.2505
R40426 ASIG5V.n4859 ASIG5V.n4858 2.2505
R40427 ASIG5V.n4863 ASIG5V.n4862 2.2505
R40428 ASIG5V.n4860 ASIG5V.n3256 2.2505
R40429 ASIG5V.n4868 ASIG5V.n4867 2.2505
R40430 ASIG5V.n4871 ASIG5V.n4870 2.2505
R40431 ASIG5V.n4875 ASIG5V.n4874 2.2505
R40432 ASIG5V.n4872 ASIG5V.n3254 2.2505
R40433 ASIG5V.n4880 ASIG5V.n4879 2.2505
R40434 ASIG5V.n4883 ASIG5V.n4882 2.2505
R40435 ASIG5V.n4887 ASIG5V.n4886 2.2505
R40436 ASIG5V.n4884 ASIG5V.n3252 2.2505
R40437 ASIG5V.n4892 ASIG5V.n4891 2.2505
R40438 ASIG5V.n4895 ASIG5V.n4894 2.2505
R40439 ASIG5V.n4899 ASIG5V.n4898 2.2505
R40440 ASIG5V.n4896 ASIG5V.n3250 2.2505
R40441 ASIG5V.n4904 ASIG5V.n4903 2.2505
R40442 ASIG5V.n4907 ASIG5V.n4906 2.2505
R40443 ASIG5V.n4911 ASIG5V.n4910 2.2505
R40444 ASIG5V.n4908 ASIG5V.n3248 2.2505
R40445 ASIG5V.n4916 ASIG5V.n4915 2.2505
R40446 ASIG5V.n4919 ASIG5V.n4918 2.2505
R40447 ASIG5V.n4923 ASIG5V.n4922 2.2505
R40448 ASIG5V.n4920 ASIG5V.n3246 2.2505
R40449 ASIG5V.n4928 ASIG5V.n4927 2.2505
R40450 ASIG5V.n4931 ASIG5V.n4930 2.2505
R40451 ASIG5V.n4935 ASIG5V.n4934 2.2505
R40452 ASIG5V.n4932 ASIG5V.n3244 2.2505
R40453 ASIG5V.n4940 ASIG5V.n4939 2.2505
R40454 ASIG5V.n4943 ASIG5V.n4942 2.2505
R40455 ASIG5V.n4947 ASIG5V.n4946 2.2505
R40456 ASIG5V.n4944 ASIG5V.n3242 2.2505
R40457 ASIG5V.n4952 ASIG5V.n4951 2.2505
R40458 ASIG5V.n4955 ASIG5V.n4954 2.2505
R40459 ASIG5V.n4959 ASIG5V.n4958 2.2505
R40460 ASIG5V.n4956 ASIG5V.n3240 2.2505
R40461 ASIG5V.n4964 ASIG5V.n4963 2.2505
R40462 ASIG5V.n4967 ASIG5V.n4966 2.2505
R40463 ASIG5V.n4971 ASIG5V.n4970 2.2505
R40464 ASIG5V.n4968 ASIG5V.n3238 2.2505
R40465 ASIG5V.n4976 ASIG5V.n4975 2.2505
R40466 ASIG5V.n4979 ASIG5V.n4978 2.2505
R40467 ASIG5V.n4983 ASIG5V.n4982 2.2505
R40468 ASIG5V.n4980 ASIG5V.n3236 2.2505
R40469 ASIG5V.n4988 ASIG5V.n4987 2.2505
R40470 ASIG5V.n4991 ASIG5V.n4990 2.2505
R40471 ASIG5V.n4995 ASIG5V.n4994 2.2505
R40472 ASIG5V.n4992 ASIG5V.n3234 2.2505
R40473 ASIG5V.n5000 ASIG5V.n4999 2.2505
R40474 ASIG5V.n5003 ASIG5V.n5002 2.2505
R40475 ASIG5V.n5007 ASIG5V.n5006 2.2505
R40476 ASIG5V.n5004 ASIG5V.n3232 2.2505
R40477 ASIG5V.n5012 ASIG5V.n5011 2.2505
R40478 ASIG5V.n5015 ASIG5V.n5014 2.2505
R40479 ASIG5V.n5019 ASIG5V.n5018 2.2505
R40480 ASIG5V.n5016 ASIG5V.n3230 2.2505
R40481 ASIG5V.n5024 ASIG5V.n5023 2.2505
R40482 ASIG5V.n5027 ASIG5V.n5026 2.2505
R40483 ASIG5V.n5031 ASIG5V.n5030 2.2505
R40484 ASIG5V.n5028 ASIG5V.n3228 2.2505
R40485 ASIG5V.n5036 ASIG5V.n5035 2.2505
R40486 ASIG5V.n5039 ASIG5V.n5038 2.2505
R40487 ASIG5V.n5043 ASIG5V.n5042 2.2505
R40488 ASIG5V.n5040 ASIG5V.n3226 2.2505
R40489 ASIG5V.n5048 ASIG5V.n5047 2.2505
R40490 ASIG5V.n5051 ASIG5V.n5050 2.2505
R40491 ASIG5V.n5055 ASIG5V.n5054 2.2505
R40492 ASIG5V.n5052 ASIG5V.n3224 2.2505
R40493 ASIG5V.n5061 ASIG5V.n5060 2.2505
R40494 ASIG5V.n5063 ASIG5V.n3222 2.2505
R40495 ASIG5V.n9442 ASIG5V.n5070 2.2505
R40496 ASIG5V.n9730 ASIG5V.n9729 2.2505
R40497 ASIG5V.n9728 ASIG5V.n9443 2.2505
R40498 ASIG5V.n9727 ASIG5V.n9726 2.2505
R40499 ASIG5V.n9722 ASIG5V.n9444 2.2505
R40500 ASIG5V.n9718 ASIG5V.n9717 2.2505
R40501 ASIG5V.n9716 ASIG5V.n9445 2.2505
R40502 ASIG5V.n9715 ASIG5V.n9714 2.2505
R40503 ASIG5V.n9710 ASIG5V.n9446 2.2505
R40504 ASIG5V.n9706 ASIG5V.n9705 2.2505
R40505 ASIG5V.n9704 ASIG5V.n9447 2.2505
R40506 ASIG5V.n9703 ASIG5V.n9702 2.2505
R40507 ASIG5V.n9698 ASIG5V.n9448 2.2505
R40508 ASIG5V.n9694 ASIG5V.n9693 2.2505
R40509 ASIG5V.n9692 ASIG5V.n9449 2.2505
R40510 ASIG5V.n9691 ASIG5V.n9690 2.2505
R40511 ASIG5V.n9686 ASIG5V.n9450 2.2505
R40512 ASIG5V.n9682 ASIG5V.n9681 2.2505
R40513 ASIG5V.n9680 ASIG5V.n9451 2.2505
R40514 ASIG5V.n9679 ASIG5V.n9678 2.2505
R40515 ASIG5V.n9674 ASIG5V.n9452 2.2505
R40516 ASIG5V.n9670 ASIG5V.n9669 2.2505
R40517 ASIG5V.n9668 ASIG5V.n9453 2.2505
R40518 ASIG5V.n9667 ASIG5V.n9666 2.2505
R40519 ASIG5V.n9662 ASIG5V.n9454 2.2505
R40520 ASIG5V.n9658 ASIG5V.n9657 2.2505
R40521 ASIG5V.n9656 ASIG5V.n9455 2.2505
R40522 ASIG5V.n9655 ASIG5V.n9654 2.2505
R40523 ASIG5V.n9650 ASIG5V.n9456 2.2505
R40524 ASIG5V.n9646 ASIG5V.n9645 2.2505
R40525 ASIG5V.n9644 ASIG5V.n9457 2.2505
R40526 ASIG5V.n9643 ASIG5V.n9642 2.2505
R40527 ASIG5V.n9638 ASIG5V.n9458 2.2505
R40528 ASIG5V.n9634 ASIG5V.n9633 2.2505
R40529 ASIG5V.n9632 ASIG5V.n9459 2.2505
R40530 ASIG5V.n9631 ASIG5V.n9630 2.2505
R40531 ASIG5V.n9626 ASIG5V.n9460 2.2505
R40532 ASIG5V.n9622 ASIG5V.n9621 2.2505
R40533 ASIG5V.n9620 ASIG5V.n9461 2.2505
R40534 ASIG5V.n9619 ASIG5V.n9618 2.2505
R40535 ASIG5V.n9614 ASIG5V.n9462 2.2505
R40536 ASIG5V.n9610 ASIG5V.n9609 2.2505
R40537 ASIG5V.n9608 ASIG5V.n9463 2.2505
R40538 ASIG5V.n9607 ASIG5V.n9606 2.2505
R40539 ASIG5V.n9602 ASIG5V.n9464 2.2505
R40540 ASIG5V.n9598 ASIG5V.n9597 2.2505
R40541 ASIG5V.n9596 ASIG5V.n9465 2.2505
R40542 ASIG5V.n9595 ASIG5V.n9594 2.2505
R40543 ASIG5V.n9590 ASIG5V.n9466 2.2505
R40544 ASIG5V.n9586 ASIG5V.n9585 2.2505
R40545 ASIG5V.n9584 ASIG5V.n9467 2.2505
R40546 ASIG5V.n9583 ASIG5V.n9582 2.2505
R40547 ASIG5V.n9578 ASIG5V.n9468 2.2505
R40548 ASIG5V.n9574 ASIG5V.n9573 2.2505
R40549 ASIG5V.n9572 ASIG5V.n9469 2.2505
R40550 ASIG5V.n9571 ASIG5V.n9570 2.2505
R40551 ASIG5V.n9566 ASIG5V.n9470 2.2505
R40552 ASIG5V.n9562 ASIG5V.n9561 2.2505
R40553 ASIG5V.n9560 ASIG5V.n9471 2.2505
R40554 ASIG5V.n9559 ASIG5V.n9558 2.2505
R40555 ASIG5V.n9554 ASIG5V.n9472 2.2505
R40556 ASIG5V.n9550 ASIG5V.n9549 2.2505
R40557 ASIG5V.n9548 ASIG5V.n9473 2.2505
R40558 ASIG5V.n9547 ASIG5V.n9546 2.2505
R40559 ASIG5V.n9542 ASIG5V.n9474 2.2505
R40560 ASIG5V.n9538 ASIG5V.n9537 2.2505
R40561 ASIG5V.n9536 ASIG5V.n9475 2.2505
R40562 ASIG5V.n9535 ASIG5V.n9534 2.2505
R40563 ASIG5V.n9530 ASIG5V.n9476 2.2505
R40564 ASIG5V.n9526 ASIG5V.n9525 2.2505
R40565 ASIG5V.n9524 ASIG5V.n9477 2.2505
R40566 ASIG5V.n9523 ASIG5V.n9522 2.2505
R40567 ASIG5V.n9518 ASIG5V.n9478 2.2505
R40568 ASIG5V.n9514 ASIG5V.n9513 2.2505
R40569 ASIG5V.n9512 ASIG5V.n9479 2.2505
R40570 ASIG5V.n9511 ASIG5V.n9510 2.2505
R40571 ASIG5V.n9506 ASIG5V.n9480 2.2505
R40572 ASIG5V.n9502 ASIG5V.n9501 2.2505
R40573 ASIG5V.n9500 ASIG5V.n9481 2.2505
R40574 ASIG5V.n9499 ASIG5V.n9498 2.2505
R40575 ASIG5V.n9494 ASIG5V.n9482 2.2505
R40576 ASIG5V.n9490 ASIG5V.n9489 2.2505
R40577 ASIG5V.n9488 ASIG5V.n9485 2.2505
R40578 ASIG5V.n9487 ASIG5V.n9486 2.2505
R40579 ASIG5V.n9486 ASIG5V.n5116 2.2505
R40580 ASIG5V.n9485 ASIG5V.n9484 2.2505
R40581 ASIG5V.n9491 ASIG5V.n9490 2.2505
R40582 ASIG5V.n9494 ASIG5V.n9493 2.2505
R40583 ASIG5V.n9498 ASIG5V.n9497 2.2505
R40584 ASIG5V.n9495 ASIG5V.n9481 2.2505
R40585 ASIG5V.n9503 ASIG5V.n9502 2.2505
R40586 ASIG5V.n9506 ASIG5V.n9505 2.2505
R40587 ASIG5V.n9510 ASIG5V.n9509 2.2505
R40588 ASIG5V.n9507 ASIG5V.n9479 2.2505
R40589 ASIG5V.n9515 ASIG5V.n9514 2.2505
R40590 ASIG5V.n9518 ASIG5V.n9517 2.2505
R40591 ASIG5V.n9522 ASIG5V.n9521 2.2505
R40592 ASIG5V.n9519 ASIG5V.n9477 2.2505
R40593 ASIG5V.n9527 ASIG5V.n9526 2.2505
R40594 ASIG5V.n9530 ASIG5V.n9529 2.2505
R40595 ASIG5V.n9534 ASIG5V.n9533 2.2505
R40596 ASIG5V.n9531 ASIG5V.n9475 2.2505
R40597 ASIG5V.n9539 ASIG5V.n9538 2.2505
R40598 ASIG5V.n9542 ASIG5V.n9541 2.2505
R40599 ASIG5V.n9546 ASIG5V.n9545 2.2505
R40600 ASIG5V.n9543 ASIG5V.n9473 2.2505
R40601 ASIG5V.n9551 ASIG5V.n9550 2.2505
R40602 ASIG5V.n9554 ASIG5V.n9553 2.2505
R40603 ASIG5V.n9558 ASIG5V.n9557 2.2505
R40604 ASIG5V.n9555 ASIG5V.n9471 2.2505
R40605 ASIG5V.n9563 ASIG5V.n9562 2.2505
R40606 ASIG5V.n9566 ASIG5V.n9565 2.2505
R40607 ASIG5V.n9570 ASIG5V.n9569 2.2505
R40608 ASIG5V.n9567 ASIG5V.n9469 2.2505
R40609 ASIG5V.n9575 ASIG5V.n9574 2.2505
R40610 ASIG5V.n9578 ASIG5V.n9577 2.2505
R40611 ASIG5V.n9582 ASIG5V.n9581 2.2505
R40612 ASIG5V.n9579 ASIG5V.n9467 2.2505
R40613 ASIG5V.n9587 ASIG5V.n9586 2.2505
R40614 ASIG5V.n9590 ASIG5V.n9589 2.2505
R40615 ASIG5V.n9594 ASIG5V.n9593 2.2505
R40616 ASIG5V.n9591 ASIG5V.n9465 2.2505
R40617 ASIG5V.n9599 ASIG5V.n9598 2.2505
R40618 ASIG5V.n9602 ASIG5V.n9601 2.2505
R40619 ASIG5V.n9606 ASIG5V.n9605 2.2505
R40620 ASIG5V.n9603 ASIG5V.n9463 2.2505
R40621 ASIG5V.n9611 ASIG5V.n9610 2.2505
R40622 ASIG5V.n9614 ASIG5V.n9613 2.2505
R40623 ASIG5V.n9618 ASIG5V.n9617 2.2505
R40624 ASIG5V.n9615 ASIG5V.n9461 2.2505
R40625 ASIG5V.n9623 ASIG5V.n9622 2.2505
R40626 ASIG5V.n9626 ASIG5V.n9625 2.2505
R40627 ASIG5V.n9630 ASIG5V.n9629 2.2505
R40628 ASIG5V.n9627 ASIG5V.n9459 2.2505
R40629 ASIG5V.n9635 ASIG5V.n9634 2.2505
R40630 ASIG5V.n9638 ASIG5V.n9637 2.2505
R40631 ASIG5V.n9642 ASIG5V.n9641 2.2505
R40632 ASIG5V.n9639 ASIG5V.n9457 2.2505
R40633 ASIG5V.n9647 ASIG5V.n9646 2.2505
R40634 ASIG5V.n9650 ASIG5V.n9649 2.2505
R40635 ASIG5V.n9654 ASIG5V.n9653 2.2505
R40636 ASIG5V.n9651 ASIG5V.n9455 2.2505
R40637 ASIG5V.n9659 ASIG5V.n9658 2.2505
R40638 ASIG5V.n9662 ASIG5V.n9661 2.2505
R40639 ASIG5V.n9666 ASIG5V.n9665 2.2505
R40640 ASIG5V.n9663 ASIG5V.n9453 2.2505
R40641 ASIG5V.n9671 ASIG5V.n9670 2.2505
R40642 ASIG5V.n9674 ASIG5V.n9673 2.2505
R40643 ASIG5V.n9678 ASIG5V.n9677 2.2505
R40644 ASIG5V.n9675 ASIG5V.n9451 2.2505
R40645 ASIG5V.n9683 ASIG5V.n9682 2.2505
R40646 ASIG5V.n9686 ASIG5V.n9685 2.2505
R40647 ASIG5V.n9690 ASIG5V.n9689 2.2505
R40648 ASIG5V.n9687 ASIG5V.n9449 2.2505
R40649 ASIG5V.n9695 ASIG5V.n9694 2.2505
R40650 ASIG5V.n9698 ASIG5V.n9697 2.2505
R40651 ASIG5V.n9702 ASIG5V.n9701 2.2505
R40652 ASIG5V.n9699 ASIG5V.n9447 2.2505
R40653 ASIG5V.n9707 ASIG5V.n9706 2.2505
R40654 ASIG5V.n9710 ASIG5V.n9709 2.2505
R40655 ASIG5V.n9714 ASIG5V.n9713 2.2505
R40656 ASIG5V.n9711 ASIG5V.n9445 2.2505
R40657 ASIG5V.n9719 ASIG5V.n9718 2.2505
R40658 ASIG5V.n9722 ASIG5V.n9721 2.2505
R40659 ASIG5V.n9726 ASIG5V.n9725 2.2505
R40660 ASIG5V.n9723 ASIG5V.n9443 2.2505
R40661 ASIG5V.n9731 ASIG5V.n9730 2.2505
R40662 ASIG5V.n9733 ASIG5V.n9442 2.2505
R40663 ASIG5V.n9426 ASIG5V.n5168 2.2505
R40664 ASIG5V.n9428 ASIG5V.n9427 2.2505
R40665 ASIG5V.n5456 ASIG5V.n5171 2.2505
R40666 ASIG5V.n5455 ASIG5V.n5454 2.2505
R40667 ASIG5V.n5450 ASIG5V.n5172 2.2505
R40668 ASIG5V.n5446 ASIG5V.n5445 2.2505
R40669 ASIG5V.n5444 ASIG5V.n5173 2.2505
R40670 ASIG5V.n5443 ASIG5V.n5442 2.2505
R40671 ASIG5V.n5438 ASIG5V.n5174 2.2505
R40672 ASIG5V.n5434 ASIG5V.n5433 2.2505
R40673 ASIG5V.n5432 ASIG5V.n5175 2.2505
R40674 ASIG5V.n5431 ASIG5V.n5430 2.2505
R40675 ASIG5V.n5426 ASIG5V.n5176 2.2505
R40676 ASIG5V.n5422 ASIG5V.n5421 2.2505
R40677 ASIG5V.n5420 ASIG5V.n5177 2.2505
R40678 ASIG5V.n5419 ASIG5V.n5418 2.2505
R40679 ASIG5V.n5414 ASIG5V.n5178 2.2505
R40680 ASIG5V.n5410 ASIG5V.n5409 2.2505
R40681 ASIG5V.n5408 ASIG5V.n5179 2.2505
R40682 ASIG5V.n5407 ASIG5V.n5406 2.2505
R40683 ASIG5V.n5402 ASIG5V.n5180 2.2505
R40684 ASIG5V.n5398 ASIG5V.n5397 2.2505
R40685 ASIG5V.n5396 ASIG5V.n5181 2.2505
R40686 ASIG5V.n5395 ASIG5V.n5394 2.2505
R40687 ASIG5V.n5390 ASIG5V.n5182 2.2505
R40688 ASIG5V.n5386 ASIG5V.n5385 2.2505
R40689 ASIG5V.n5384 ASIG5V.n5183 2.2505
R40690 ASIG5V.n5383 ASIG5V.n5382 2.2505
R40691 ASIG5V.n5378 ASIG5V.n5184 2.2505
R40692 ASIG5V.n5374 ASIG5V.n5373 2.2505
R40693 ASIG5V.n5372 ASIG5V.n5185 2.2505
R40694 ASIG5V.n5371 ASIG5V.n5370 2.2505
R40695 ASIG5V.n5366 ASIG5V.n5186 2.2505
R40696 ASIG5V.n5362 ASIG5V.n5361 2.2505
R40697 ASIG5V.n5360 ASIG5V.n5187 2.2505
R40698 ASIG5V.n5359 ASIG5V.n5358 2.2505
R40699 ASIG5V.n5354 ASIG5V.n5188 2.2505
R40700 ASIG5V.n5350 ASIG5V.n5349 2.2505
R40701 ASIG5V.n5348 ASIG5V.n5189 2.2505
R40702 ASIG5V.n5347 ASIG5V.n5346 2.2505
R40703 ASIG5V.n5342 ASIG5V.n5190 2.2505
R40704 ASIG5V.n5338 ASIG5V.n5337 2.2505
R40705 ASIG5V.n5336 ASIG5V.n5191 2.2505
R40706 ASIG5V.n5335 ASIG5V.n5334 2.2505
R40707 ASIG5V.n5330 ASIG5V.n5192 2.2505
R40708 ASIG5V.n5326 ASIG5V.n5325 2.2505
R40709 ASIG5V.n5324 ASIG5V.n5193 2.2505
R40710 ASIG5V.n5323 ASIG5V.n5322 2.2505
R40711 ASIG5V.n5318 ASIG5V.n5194 2.2505
R40712 ASIG5V.n5314 ASIG5V.n5313 2.2505
R40713 ASIG5V.n5312 ASIG5V.n5195 2.2505
R40714 ASIG5V.n5311 ASIG5V.n5310 2.2505
R40715 ASIG5V.n5306 ASIG5V.n5196 2.2505
R40716 ASIG5V.n5302 ASIG5V.n5301 2.2505
R40717 ASIG5V.n5300 ASIG5V.n5197 2.2505
R40718 ASIG5V.n5299 ASIG5V.n5298 2.2505
R40719 ASIG5V.n5294 ASIG5V.n5198 2.2505
R40720 ASIG5V.n5290 ASIG5V.n5289 2.2505
R40721 ASIG5V.n5288 ASIG5V.n5199 2.2505
R40722 ASIG5V.n5287 ASIG5V.n5286 2.2505
R40723 ASIG5V.n5282 ASIG5V.n5200 2.2505
R40724 ASIG5V.n5278 ASIG5V.n5277 2.2505
R40725 ASIG5V.n5276 ASIG5V.n5201 2.2505
R40726 ASIG5V.n5275 ASIG5V.n5274 2.2505
R40727 ASIG5V.n5270 ASIG5V.n5202 2.2505
R40728 ASIG5V.n5266 ASIG5V.n5265 2.2505
R40729 ASIG5V.n5264 ASIG5V.n5203 2.2505
R40730 ASIG5V.n5263 ASIG5V.n5262 2.2505
R40731 ASIG5V.n5258 ASIG5V.n5204 2.2505
R40732 ASIG5V.n5254 ASIG5V.n5253 2.2505
R40733 ASIG5V.n5252 ASIG5V.n5205 2.2505
R40734 ASIG5V.n5251 ASIG5V.n5250 2.2505
R40735 ASIG5V.n5246 ASIG5V.n5206 2.2505
R40736 ASIG5V.n5242 ASIG5V.n5241 2.2505
R40737 ASIG5V.n5240 ASIG5V.n5207 2.2505
R40738 ASIG5V.n5239 ASIG5V.n5238 2.2505
R40739 ASIG5V.n5234 ASIG5V.n5208 2.2505
R40740 ASIG5V.n5230 ASIG5V.n5229 2.2505
R40741 ASIG5V.n5228 ASIG5V.n5209 2.2505
R40742 ASIG5V.n5227 ASIG5V.n5226 2.2505
R40743 ASIG5V.n5222 ASIG5V.n5210 2.2505
R40744 ASIG5V.n5218 ASIG5V.n5217 2.2505
R40745 ASIG5V.n5216 ASIG5V.n5213 2.2505
R40746 ASIG5V.n5215 ASIG5V.n5214 2.2505
R40747 ASIG5V.n5214 ASIG5V.n5165 2.2505
R40748 ASIG5V.n5213 ASIG5V.n5212 2.2505
R40749 ASIG5V.n5219 ASIG5V.n5218 2.2505
R40750 ASIG5V.n5222 ASIG5V.n5221 2.2505
R40751 ASIG5V.n5226 ASIG5V.n5225 2.2505
R40752 ASIG5V.n5223 ASIG5V.n5209 2.2505
R40753 ASIG5V.n5231 ASIG5V.n5230 2.2505
R40754 ASIG5V.n5234 ASIG5V.n5233 2.2505
R40755 ASIG5V.n5238 ASIG5V.n5237 2.2505
R40756 ASIG5V.n5235 ASIG5V.n5207 2.2505
R40757 ASIG5V.n5243 ASIG5V.n5242 2.2505
R40758 ASIG5V.n5246 ASIG5V.n5245 2.2505
R40759 ASIG5V.n5250 ASIG5V.n5249 2.2505
R40760 ASIG5V.n5247 ASIG5V.n5205 2.2505
R40761 ASIG5V.n5255 ASIG5V.n5254 2.2505
R40762 ASIG5V.n5258 ASIG5V.n5257 2.2505
R40763 ASIG5V.n5262 ASIG5V.n5261 2.2505
R40764 ASIG5V.n5259 ASIG5V.n5203 2.2505
R40765 ASIG5V.n5267 ASIG5V.n5266 2.2505
R40766 ASIG5V.n5270 ASIG5V.n5269 2.2505
R40767 ASIG5V.n5274 ASIG5V.n5273 2.2505
R40768 ASIG5V.n5271 ASIG5V.n5201 2.2505
R40769 ASIG5V.n5279 ASIG5V.n5278 2.2505
R40770 ASIG5V.n5282 ASIG5V.n5281 2.2505
R40771 ASIG5V.n5286 ASIG5V.n5285 2.2505
R40772 ASIG5V.n5283 ASIG5V.n5199 2.2505
R40773 ASIG5V.n5291 ASIG5V.n5290 2.2505
R40774 ASIG5V.n5294 ASIG5V.n5293 2.2505
R40775 ASIG5V.n5298 ASIG5V.n5297 2.2505
R40776 ASIG5V.n5295 ASIG5V.n5197 2.2505
R40777 ASIG5V.n5303 ASIG5V.n5302 2.2505
R40778 ASIG5V.n5306 ASIG5V.n5305 2.2505
R40779 ASIG5V.n5310 ASIG5V.n5309 2.2505
R40780 ASIG5V.n5307 ASIG5V.n5195 2.2505
R40781 ASIG5V.n5315 ASIG5V.n5314 2.2505
R40782 ASIG5V.n5318 ASIG5V.n5317 2.2505
R40783 ASIG5V.n5322 ASIG5V.n5321 2.2505
R40784 ASIG5V.n5319 ASIG5V.n5193 2.2505
R40785 ASIG5V.n5327 ASIG5V.n5326 2.2505
R40786 ASIG5V.n5330 ASIG5V.n5329 2.2505
R40787 ASIG5V.n5334 ASIG5V.n5333 2.2505
R40788 ASIG5V.n5331 ASIG5V.n5191 2.2505
R40789 ASIG5V.n5339 ASIG5V.n5338 2.2505
R40790 ASIG5V.n5342 ASIG5V.n5341 2.2505
R40791 ASIG5V.n5346 ASIG5V.n5345 2.2505
R40792 ASIG5V.n5343 ASIG5V.n5189 2.2505
R40793 ASIG5V.n5351 ASIG5V.n5350 2.2505
R40794 ASIG5V.n5354 ASIG5V.n5353 2.2505
R40795 ASIG5V.n5358 ASIG5V.n5357 2.2505
R40796 ASIG5V.n5355 ASIG5V.n5187 2.2505
R40797 ASIG5V.n5363 ASIG5V.n5362 2.2505
R40798 ASIG5V.n5366 ASIG5V.n5365 2.2505
R40799 ASIG5V.n5370 ASIG5V.n5369 2.2505
R40800 ASIG5V.n5367 ASIG5V.n5185 2.2505
R40801 ASIG5V.n5375 ASIG5V.n5374 2.2505
R40802 ASIG5V.n5378 ASIG5V.n5377 2.2505
R40803 ASIG5V.n5382 ASIG5V.n5381 2.2505
R40804 ASIG5V.n5379 ASIG5V.n5183 2.2505
R40805 ASIG5V.n5387 ASIG5V.n5386 2.2505
R40806 ASIG5V.n5390 ASIG5V.n5389 2.2505
R40807 ASIG5V.n5394 ASIG5V.n5393 2.2505
R40808 ASIG5V.n5391 ASIG5V.n5181 2.2505
R40809 ASIG5V.n5399 ASIG5V.n5398 2.2505
R40810 ASIG5V.n5402 ASIG5V.n5401 2.2505
R40811 ASIG5V.n5406 ASIG5V.n5405 2.2505
R40812 ASIG5V.n5403 ASIG5V.n5179 2.2505
R40813 ASIG5V.n5411 ASIG5V.n5410 2.2505
R40814 ASIG5V.n5414 ASIG5V.n5413 2.2505
R40815 ASIG5V.n5418 ASIG5V.n5417 2.2505
R40816 ASIG5V.n5415 ASIG5V.n5177 2.2505
R40817 ASIG5V.n5423 ASIG5V.n5422 2.2505
R40818 ASIG5V.n5426 ASIG5V.n5425 2.2505
R40819 ASIG5V.n5430 ASIG5V.n5429 2.2505
R40820 ASIG5V.n5427 ASIG5V.n5175 2.2505
R40821 ASIG5V.n5435 ASIG5V.n5434 2.2505
R40822 ASIG5V.n5438 ASIG5V.n5437 2.2505
R40823 ASIG5V.n5442 ASIG5V.n5441 2.2505
R40824 ASIG5V.n5439 ASIG5V.n5173 2.2505
R40825 ASIG5V.n5447 ASIG5V.n5446 2.2505
R40826 ASIG5V.n5450 ASIG5V.n5449 2.2505
R40827 ASIG5V.n5454 ASIG5V.n5453 2.2505
R40828 ASIG5V.n5451 ASIG5V.n5171 2.2505
R40829 ASIG5V.n9429 ASIG5V.n9428 2.2505
R40830 ASIG5V.n9431 ASIG5V.n5168 2.2505
R40831 ASIG5V.n9414 ASIG5V.n5557 2.2505
R40832 ASIG5V.n7777 ASIG5V.n5556 2.2505
R40833 ASIG5V.n7780 ASIG5V.n7779 2.2505
R40834 ASIG5V.n7781 ASIG5V.n7776 2.2505
R40835 ASIG5V.n7784 ASIG5V.n7782 2.2505
R40836 ASIG5V.n7786 ASIG5V.n7774 2.2505
R40837 ASIG5V.n7789 ASIG5V.n7788 2.2505
R40838 ASIG5V.n7790 ASIG5V.n7773 2.2505
R40839 ASIG5V.n7793 ASIG5V.n7791 2.2505
R40840 ASIG5V.n7795 ASIG5V.n7771 2.2505
R40841 ASIG5V.n7798 ASIG5V.n7797 2.2505
R40842 ASIG5V.n7799 ASIG5V.n7770 2.2505
R40843 ASIG5V.n7802 ASIG5V.n7800 2.2505
R40844 ASIG5V.n7804 ASIG5V.n7768 2.2505
R40845 ASIG5V.n7807 ASIG5V.n7806 2.2505
R40846 ASIG5V.n7808 ASIG5V.n7767 2.2505
R40847 ASIG5V.n7811 ASIG5V.n7809 2.2505
R40848 ASIG5V.n7813 ASIG5V.n7765 2.2505
R40849 ASIG5V.n7816 ASIG5V.n7815 2.2505
R40850 ASIG5V.n7817 ASIG5V.n7764 2.2505
R40851 ASIG5V.n7820 ASIG5V.n7818 2.2505
R40852 ASIG5V.n7822 ASIG5V.n7762 2.2505
R40853 ASIG5V.n7825 ASIG5V.n7824 2.2505
R40854 ASIG5V.n7826 ASIG5V.n7761 2.2505
R40855 ASIG5V.n7829 ASIG5V.n7827 2.2505
R40856 ASIG5V.n7831 ASIG5V.n7759 2.2505
R40857 ASIG5V.n7834 ASIG5V.n7833 2.2505
R40858 ASIG5V.n7835 ASIG5V.n7758 2.2505
R40859 ASIG5V.n7838 ASIG5V.n7836 2.2505
R40860 ASIG5V.n7840 ASIG5V.n7756 2.2505
R40861 ASIG5V.n7843 ASIG5V.n7842 2.2505
R40862 ASIG5V.n7844 ASIG5V.n7755 2.2505
R40863 ASIG5V.n7847 ASIG5V.n7845 2.2505
R40864 ASIG5V.n7849 ASIG5V.n7753 2.2505
R40865 ASIG5V.n7852 ASIG5V.n7851 2.2505
R40866 ASIG5V.n7853 ASIG5V.n7752 2.2505
R40867 ASIG5V.n7856 ASIG5V.n7854 2.2505
R40868 ASIG5V.n7858 ASIG5V.n7750 2.2505
R40869 ASIG5V.n7861 ASIG5V.n7860 2.2505
R40870 ASIG5V.n7862 ASIG5V.n7749 2.2505
R40871 ASIG5V.n7865 ASIG5V.n7863 2.2505
R40872 ASIG5V.n7867 ASIG5V.n7747 2.2505
R40873 ASIG5V.n7870 ASIG5V.n7869 2.2505
R40874 ASIG5V.n7871 ASIG5V.n7746 2.2505
R40875 ASIG5V.n7874 ASIG5V.n7872 2.2505
R40876 ASIG5V.n7876 ASIG5V.n7744 2.2505
R40877 ASIG5V.n7879 ASIG5V.n7878 2.2505
R40878 ASIG5V.n7880 ASIG5V.n7743 2.2505
R40879 ASIG5V.n7883 ASIG5V.n7881 2.2505
R40880 ASIG5V.n7885 ASIG5V.n7741 2.2505
R40881 ASIG5V.n7888 ASIG5V.n7887 2.2505
R40882 ASIG5V.n7889 ASIG5V.n7740 2.2505
R40883 ASIG5V.n7892 ASIG5V.n7890 2.2505
R40884 ASIG5V.n7894 ASIG5V.n7738 2.2505
R40885 ASIG5V.n7897 ASIG5V.n7896 2.2505
R40886 ASIG5V.n7898 ASIG5V.n7737 2.2505
R40887 ASIG5V.n7901 ASIG5V.n7899 2.2505
R40888 ASIG5V.n7903 ASIG5V.n7735 2.2505
R40889 ASIG5V.n7906 ASIG5V.n7905 2.2505
R40890 ASIG5V.n7907 ASIG5V.n7734 2.2505
R40891 ASIG5V.n7910 ASIG5V.n7908 2.2505
R40892 ASIG5V.n7912 ASIG5V.n7732 2.2505
R40893 ASIG5V.n7915 ASIG5V.n7914 2.2505
R40894 ASIG5V.n7916 ASIG5V.n7731 2.2505
R40895 ASIG5V.n7919 ASIG5V.n7917 2.2505
R40896 ASIG5V.n7921 ASIG5V.n7729 2.2505
R40897 ASIG5V.n7924 ASIG5V.n7923 2.2505
R40898 ASIG5V.n7925 ASIG5V.n7728 2.2505
R40899 ASIG5V.n7928 ASIG5V.n7926 2.2505
R40900 ASIG5V.n7930 ASIG5V.n7726 2.2505
R40901 ASIG5V.n7933 ASIG5V.n7932 2.2505
R40902 ASIG5V.n7934 ASIG5V.n7725 2.2505
R40903 ASIG5V.n7937 ASIG5V.n7935 2.2505
R40904 ASIG5V.n7939 ASIG5V.n7723 2.2505
R40905 ASIG5V.n7942 ASIG5V.n7941 2.2505
R40906 ASIG5V.n7943 ASIG5V.n7722 2.2505
R40907 ASIG5V.n7946 ASIG5V.n7944 2.2505
R40908 ASIG5V.n7948 ASIG5V.n7720 2.2505
R40909 ASIG5V.n7951 ASIG5V.n7950 2.2505
R40910 ASIG5V.n7952 ASIG5V.n7719 2.2505
R40911 ASIG5V.n7955 ASIG5V.n7953 2.2505
R40912 ASIG5V.n7957 ASIG5V.n7717 2.2505
R40913 ASIG5V.n7959 ASIG5V.n7958 2.2505
R40914 ASIG5V.n7960 ASIG5V.n5509 2.2505
R40915 ASIG5V.n9417 ASIG5V.n5509 2.2505
R40916 ASIG5V.n7958 ASIG5V.n5507 2.2505
R40917 ASIG5V.n7957 ASIG5V.n7956 2.2505
R40918 ASIG5V.n7955 ASIG5V.n7954 2.2505
R40919 ASIG5V.n7719 ASIG5V.n7718 2.2505
R40920 ASIG5V.n7950 ASIG5V.n7949 2.2505
R40921 ASIG5V.n7948 ASIG5V.n7947 2.2505
R40922 ASIG5V.n7946 ASIG5V.n7945 2.2505
R40923 ASIG5V.n7722 ASIG5V.n7721 2.2505
R40924 ASIG5V.n7941 ASIG5V.n7940 2.2505
R40925 ASIG5V.n7939 ASIG5V.n7938 2.2505
R40926 ASIG5V.n7937 ASIG5V.n7936 2.2505
R40927 ASIG5V.n7725 ASIG5V.n7724 2.2505
R40928 ASIG5V.n7932 ASIG5V.n7931 2.2505
R40929 ASIG5V.n7930 ASIG5V.n7929 2.2505
R40930 ASIG5V.n7928 ASIG5V.n7927 2.2505
R40931 ASIG5V.n7728 ASIG5V.n7727 2.2505
R40932 ASIG5V.n7923 ASIG5V.n7922 2.2505
R40933 ASIG5V.n7921 ASIG5V.n7920 2.2505
R40934 ASIG5V.n7919 ASIG5V.n7918 2.2505
R40935 ASIG5V.n7731 ASIG5V.n7730 2.2505
R40936 ASIG5V.n7914 ASIG5V.n7913 2.2505
R40937 ASIG5V.n7912 ASIG5V.n7911 2.2505
R40938 ASIG5V.n7910 ASIG5V.n7909 2.2505
R40939 ASIG5V.n7734 ASIG5V.n7733 2.2505
R40940 ASIG5V.n7905 ASIG5V.n7904 2.2505
R40941 ASIG5V.n7903 ASIG5V.n7902 2.2505
R40942 ASIG5V.n7901 ASIG5V.n7900 2.2505
R40943 ASIG5V.n7737 ASIG5V.n7736 2.2505
R40944 ASIG5V.n7896 ASIG5V.n7895 2.2505
R40945 ASIG5V.n7894 ASIG5V.n7893 2.2505
R40946 ASIG5V.n7892 ASIG5V.n7891 2.2505
R40947 ASIG5V.n7740 ASIG5V.n7739 2.2505
R40948 ASIG5V.n7887 ASIG5V.n7886 2.2505
R40949 ASIG5V.n7885 ASIG5V.n7884 2.2505
R40950 ASIG5V.n7883 ASIG5V.n7882 2.2505
R40951 ASIG5V.n7743 ASIG5V.n7742 2.2505
R40952 ASIG5V.n7878 ASIG5V.n7877 2.2505
R40953 ASIG5V.n7876 ASIG5V.n7875 2.2505
R40954 ASIG5V.n7874 ASIG5V.n7873 2.2505
R40955 ASIG5V.n7746 ASIG5V.n7745 2.2505
R40956 ASIG5V.n7869 ASIG5V.n7868 2.2505
R40957 ASIG5V.n7867 ASIG5V.n7866 2.2505
R40958 ASIG5V.n7865 ASIG5V.n7864 2.2505
R40959 ASIG5V.n7749 ASIG5V.n7748 2.2505
R40960 ASIG5V.n7860 ASIG5V.n7859 2.2505
R40961 ASIG5V.n7858 ASIG5V.n7857 2.2505
R40962 ASIG5V.n7856 ASIG5V.n7855 2.2505
R40963 ASIG5V.n7752 ASIG5V.n7751 2.2505
R40964 ASIG5V.n7851 ASIG5V.n7850 2.2505
R40965 ASIG5V.n7849 ASIG5V.n7848 2.2505
R40966 ASIG5V.n7847 ASIG5V.n7846 2.2505
R40967 ASIG5V.n7755 ASIG5V.n7754 2.2505
R40968 ASIG5V.n7842 ASIG5V.n7841 2.2505
R40969 ASIG5V.n7840 ASIG5V.n7839 2.2505
R40970 ASIG5V.n7838 ASIG5V.n7837 2.2505
R40971 ASIG5V.n7758 ASIG5V.n7757 2.2505
R40972 ASIG5V.n7833 ASIG5V.n7832 2.2505
R40973 ASIG5V.n7831 ASIG5V.n7830 2.2505
R40974 ASIG5V.n7829 ASIG5V.n7828 2.2505
R40975 ASIG5V.n7761 ASIG5V.n7760 2.2505
R40976 ASIG5V.n7824 ASIG5V.n7823 2.2505
R40977 ASIG5V.n7822 ASIG5V.n7821 2.2505
R40978 ASIG5V.n7820 ASIG5V.n7819 2.2505
R40979 ASIG5V.n7764 ASIG5V.n7763 2.2505
R40980 ASIG5V.n7815 ASIG5V.n7814 2.2505
R40981 ASIG5V.n7813 ASIG5V.n7812 2.2505
R40982 ASIG5V.n7811 ASIG5V.n7810 2.2505
R40983 ASIG5V.n7767 ASIG5V.n7766 2.2505
R40984 ASIG5V.n7806 ASIG5V.n7805 2.2505
R40985 ASIG5V.n7804 ASIG5V.n7803 2.2505
R40986 ASIG5V.n7802 ASIG5V.n7801 2.2505
R40987 ASIG5V.n7770 ASIG5V.n7769 2.2505
R40988 ASIG5V.n7797 ASIG5V.n7796 2.2505
R40989 ASIG5V.n7795 ASIG5V.n7794 2.2505
R40990 ASIG5V.n7793 ASIG5V.n7792 2.2505
R40991 ASIG5V.n7773 ASIG5V.n7772 2.2505
R40992 ASIG5V.n7788 ASIG5V.n7787 2.2505
R40993 ASIG5V.n7786 ASIG5V.n7785 2.2505
R40994 ASIG5V.n7784 ASIG5V.n7783 2.2505
R40995 ASIG5V.n7776 ASIG5V.n7775 2.2505
R40996 ASIG5V.n7779 ASIG5V.n7778 2.2505
R40997 ASIG5V.n5556 ASIG5V.n5555 2.2505
R40998 ASIG5V.n9415 ASIG5V.n9414 2.2505
R40999 ASIG5V.n5698 ASIG5V.n5697 2.2505
R41000 ASIG5V.n5700 ASIG5V.n5699 2.2505
R41001 ASIG5V.n5692 ASIG5V.n5691 2.2505
R41002 ASIG5V.n5707 ASIG5V.n5706 2.2505
R41003 ASIG5V.n5708 ASIG5V.n5690 2.2505
R41004 ASIG5V.n5710 ASIG5V.n5709 2.2505
R41005 ASIG5V.n5686 ASIG5V.n5685 2.2505
R41006 ASIG5V.n5717 ASIG5V.n5716 2.2505
R41007 ASIG5V.n5718 ASIG5V.n5684 2.2505
R41008 ASIG5V.n5720 ASIG5V.n5719 2.2505
R41009 ASIG5V.n5680 ASIG5V.n5679 2.2505
R41010 ASIG5V.n5727 ASIG5V.n5726 2.2505
R41011 ASIG5V.n5728 ASIG5V.n5678 2.2505
R41012 ASIG5V.n5730 ASIG5V.n5729 2.2505
R41013 ASIG5V.n5674 ASIG5V.n5673 2.2505
R41014 ASIG5V.n5737 ASIG5V.n5736 2.2505
R41015 ASIG5V.n5738 ASIG5V.n5672 2.2505
R41016 ASIG5V.n5740 ASIG5V.n5739 2.2505
R41017 ASIG5V.n5668 ASIG5V.n5667 2.2505
R41018 ASIG5V.n5747 ASIG5V.n5746 2.2505
R41019 ASIG5V.n5748 ASIG5V.n5666 2.2505
R41020 ASIG5V.n5750 ASIG5V.n5749 2.2505
R41021 ASIG5V.n5662 ASIG5V.n5661 2.2505
R41022 ASIG5V.n5757 ASIG5V.n5756 2.2505
R41023 ASIG5V.n5758 ASIG5V.n5660 2.2505
R41024 ASIG5V.n5760 ASIG5V.n5759 2.2505
R41025 ASIG5V.n5656 ASIG5V.n5655 2.2505
R41026 ASIG5V.n5767 ASIG5V.n5766 2.2505
R41027 ASIG5V.n5768 ASIG5V.n5654 2.2505
R41028 ASIG5V.n5770 ASIG5V.n5769 2.2505
R41029 ASIG5V.n5650 ASIG5V.n5649 2.2505
R41030 ASIG5V.n5777 ASIG5V.n5776 2.2505
R41031 ASIG5V.n5778 ASIG5V.n5648 2.2505
R41032 ASIG5V.n5780 ASIG5V.n5779 2.2505
R41033 ASIG5V.n5644 ASIG5V.n5643 2.2505
R41034 ASIG5V.n5787 ASIG5V.n5786 2.2505
R41035 ASIG5V.n5788 ASIG5V.n5642 2.2505
R41036 ASIG5V.n5790 ASIG5V.n5789 2.2505
R41037 ASIG5V.n5638 ASIG5V.n5637 2.2505
R41038 ASIG5V.n5797 ASIG5V.n5796 2.2505
R41039 ASIG5V.n5798 ASIG5V.n5636 2.2505
R41040 ASIG5V.n5800 ASIG5V.n5799 2.2505
R41041 ASIG5V.n5632 ASIG5V.n5631 2.2505
R41042 ASIG5V.n5807 ASIG5V.n5806 2.2505
R41043 ASIG5V.n5808 ASIG5V.n5630 2.2505
R41044 ASIG5V.n5810 ASIG5V.n5809 2.2505
R41045 ASIG5V.n5626 ASIG5V.n5625 2.2505
R41046 ASIG5V.n5817 ASIG5V.n5816 2.2505
R41047 ASIG5V.n5818 ASIG5V.n5624 2.2505
R41048 ASIG5V.n5820 ASIG5V.n5819 2.2505
R41049 ASIG5V.n5620 ASIG5V.n5619 2.2505
R41050 ASIG5V.n5827 ASIG5V.n5826 2.2505
R41051 ASIG5V.n5828 ASIG5V.n5618 2.2505
R41052 ASIG5V.n5830 ASIG5V.n5829 2.2505
R41053 ASIG5V.n5614 ASIG5V.n5613 2.2505
R41054 ASIG5V.n5837 ASIG5V.n5836 2.2505
R41055 ASIG5V.n5838 ASIG5V.n5612 2.2505
R41056 ASIG5V.n5840 ASIG5V.n5839 2.2505
R41057 ASIG5V.n5608 ASIG5V.n5607 2.2505
R41058 ASIG5V.n5847 ASIG5V.n5846 2.2505
R41059 ASIG5V.n5848 ASIG5V.n5606 2.2505
R41060 ASIG5V.n5850 ASIG5V.n5849 2.2505
R41061 ASIG5V.n5602 ASIG5V.n5601 2.2505
R41062 ASIG5V.n5857 ASIG5V.n5856 2.2505
R41063 ASIG5V.n5858 ASIG5V.n5600 2.2505
R41064 ASIG5V.n5860 ASIG5V.n5859 2.2505
R41065 ASIG5V.n5596 ASIG5V.n5595 2.2505
R41066 ASIG5V.n5867 ASIG5V.n5866 2.2505
R41067 ASIG5V.n5868 ASIG5V.n5594 2.2505
R41068 ASIG5V.n5870 ASIG5V.n5869 2.2505
R41069 ASIG5V.n5590 ASIG5V.n5589 2.2505
R41070 ASIG5V.n5877 ASIG5V.n5876 2.2505
R41071 ASIG5V.n5878 ASIG5V.n5588 2.2505
R41072 ASIG5V.n5880 ASIG5V.n5879 2.2505
R41073 ASIG5V.n5584 ASIG5V.n5583 2.2505
R41074 ASIG5V.n5887 ASIG5V.n5886 2.2505
R41075 ASIG5V.n5888 ASIG5V.n5582 2.2505
R41076 ASIG5V.n5890 ASIG5V.n5889 2.2505
R41077 ASIG5V.n5578 ASIG5V.n5577 2.2505
R41078 ASIG5V.n5897 ASIG5V.n5896 2.2505
R41079 ASIG5V.n5898 ASIG5V.n5576 2.2505
R41080 ASIG5V.n5900 ASIG5V.n5899 2.2505
R41081 ASIG5V.n5574 ASIG5V.n5573 2.2505
R41082 ASIG5V.n5907 ASIG5V.n5906 2.2505
R41083 ASIG5V.n5906 ASIG5V.n5905 2.2505
R41084 ASIG5V.n5903 ASIG5V.n5574 2.2505
R41085 ASIG5V.n5901 ASIG5V.n5900 2.2505
R41086 ASIG5V.n5579 ASIG5V.n5576 2.2505
R41087 ASIG5V.n5896 ASIG5V.n5895 2.2505
R41088 ASIG5V.n5893 ASIG5V.n5578 2.2505
R41089 ASIG5V.n5891 ASIG5V.n5890 2.2505
R41090 ASIG5V.n5585 ASIG5V.n5582 2.2505
R41091 ASIG5V.n5886 ASIG5V.n5885 2.2505
R41092 ASIG5V.n5883 ASIG5V.n5584 2.2505
R41093 ASIG5V.n5881 ASIG5V.n5880 2.2505
R41094 ASIG5V.n5591 ASIG5V.n5588 2.2505
R41095 ASIG5V.n5876 ASIG5V.n5875 2.2505
R41096 ASIG5V.n5873 ASIG5V.n5590 2.2505
R41097 ASIG5V.n5871 ASIG5V.n5870 2.2505
R41098 ASIG5V.n5597 ASIG5V.n5594 2.2505
R41099 ASIG5V.n5866 ASIG5V.n5865 2.2505
R41100 ASIG5V.n5863 ASIG5V.n5596 2.2505
R41101 ASIG5V.n5861 ASIG5V.n5860 2.2505
R41102 ASIG5V.n5603 ASIG5V.n5600 2.2505
R41103 ASIG5V.n5856 ASIG5V.n5855 2.2505
R41104 ASIG5V.n5853 ASIG5V.n5602 2.2505
R41105 ASIG5V.n5851 ASIG5V.n5850 2.2505
R41106 ASIG5V.n5609 ASIG5V.n5606 2.2505
R41107 ASIG5V.n5846 ASIG5V.n5845 2.2505
R41108 ASIG5V.n5843 ASIG5V.n5608 2.2505
R41109 ASIG5V.n5841 ASIG5V.n5840 2.2505
R41110 ASIG5V.n5615 ASIG5V.n5612 2.2505
R41111 ASIG5V.n5836 ASIG5V.n5835 2.2505
R41112 ASIG5V.n5833 ASIG5V.n5614 2.2505
R41113 ASIG5V.n5831 ASIG5V.n5830 2.2505
R41114 ASIG5V.n5621 ASIG5V.n5618 2.2505
R41115 ASIG5V.n5826 ASIG5V.n5825 2.2505
R41116 ASIG5V.n5823 ASIG5V.n5620 2.2505
R41117 ASIG5V.n5821 ASIG5V.n5820 2.2505
R41118 ASIG5V.n5627 ASIG5V.n5624 2.2505
R41119 ASIG5V.n5816 ASIG5V.n5815 2.2505
R41120 ASIG5V.n5813 ASIG5V.n5626 2.2505
R41121 ASIG5V.n5811 ASIG5V.n5810 2.2505
R41122 ASIG5V.n5633 ASIG5V.n5630 2.2505
R41123 ASIG5V.n5806 ASIG5V.n5805 2.2505
R41124 ASIG5V.n5803 ASIG5V.n5632 2.2505
R41125 ASIG5V.n5801 ASIG5V.n5800 2.2505
R41126 ASIG5V.n5639 ASIG5V.n5636 2.2505
R41127 ASIG5V.n5796 ASIG5V.n5795 2.2505
R41128 ASIG5V.n5793 ASIG5V.n5638 2.2505
R41129 ASIG5V.n5791 ASIG5V.n5790 2.2505
R41130 ASIG5V.n5645 ASIG5V.n5642 2.2505
R41131 ASIG5V.n5786 ASIG5V.n5785 2.2505
R41132 ASIG5V.n5783 ASIG5V.n5644 2.2505
R41133 ASIG5V.n5781 ASIG5V.n5780 2.2505
R41134 ASIG5V.n5651 ASIG5V.n5648 2.2505
R41135 ASIG5V.n5776 ASIG5V.n5775 2.2505
R41136 ASIG5V.n5773 ASIG5V.n5650 2.2505
R41137 ASIG5V.n5771 ASIG5V.n5770 2.2505
R41138 ASIG5V.n5657 ASIG5V.n5654 2.2505
R41139 ASIG5V.n5766 ASIG5V.n5765 2.2505
R41140 ASIG5V.n5763 ASIG5V.n5656 2.2505
R41141 ASIG5V.n5761 ASIG5V.n5760 2.2505
R41142 ASIG5V.n5663 ASIG5V.n5660 2.2505
R41143 ASIG5V.n5756 ASIG5V.n5755 2.2505
R41144 ASIG5V.n5753 ASIG5V.n5662 2.2505
R41145 ASIG5V.n5751 ASIG5V.n5750 2.2505
R41146 ASIG5V.n5669 ASIG5V.n5666 2.2505
R41147 ASIG5V.n5746 ASIG5V.n5745 2.2505
R41148 ASIG5V.n5743 ASIG5V.n5668 2.2505
R41149 ASIG5V.n5741 ASIG5V.n5740 2.2505
R41150 ASIG5V.n5675 ASIG5V.n5672 2.2505
R41151 ASIG5V.n5736 ASIG5V.n5735 2.2505
R41152 ASIG5V.n5733 ASIG5V.n5674 2.2505
R41153 ASIG5V.n5731 ASIG5V.n5730 2.2505
R41154 ASIG5V.n5681 ASIG5V.n5678 2.2505
R41155 ASIG5V.n5726 ASIG5V.n5725 2.2505
R41156 ASIG5V.n5723 ASIG5V.n5680 2.2505
R41157 ASIG5V.n5721 ASIG5V.n5720 2.2505
R41158 ASIG5V.n5687 ASIG5V.n5684 2.2505
R41159 ASIG5V.n5716 ASIG5V.n5715 2.2505
R41160 ASIG5V.n5713 ASIG5V.n5686 2.2505
R41161 ASIG5V.n5711 ASIG5V.n5710 2.2505
R41162 ASIG5V.n5693 ASIG5V.n5690 2.2505
R41163 ASIG5V.n5706 ASIG5V.n5705 2.2505
R41164 ASIG5V.n5703 ASIG5V.n5692 2.2505
R41165 ASIG5V.n5701 ASIG5V.n5700 2.2505
R41166 ASIG5V.n5697 ASIG5V.n5696 2.2505
R41167 ASIG5V.n9391 ASIG5V.n6247 2.2505
R41168 ASIG5V.n6246 ASIG5V.n6002 2.2505
R41169 ASIG5V.n6245 ASIG5V.n6244 2.2505
R41170 ASIG5V.n6242 ASIG5V.n6003 2.2505
R41171 ASIG5V.n6240 ASIG5V.n6238 2.2505
R41172 ASIG5V.n6237 ASIG5V.n6005 2.2505
R41173 ASIG5V.n6236 ASIG5V.n6235 2.2505
R41174 ASIG5V.n6233 ASIG5V.n6006 2.2505
R41175 ASIG5V.n6231 ASIG5V.n6229 2.2505
R41176 ASIG5V.n6228 ASIG5V.n6008 2.2505
R41177 ASIG5V.n6227 ASIG5V.n6226 2.2505
R41178 ASIG5V.n6224 ASIG5V.n6009 2.2505
R41179 ASIG5V.n6222 ASIG5V.n6220 2.2505
R41180 ASIG5V.n6219 ASIG5V.n6011 2.2505
R41181 ASIG5V.n6218 ASIG5V.n6217 2.2505
R41182 ASIG5V.n6215 ASIG5V.n6012 2.2505
R41183 ASIG5V.n6213 ASIG5V.n6211 2.2505
R41184 ASIG5V.n6210 ASIG5V.n6014 2.2505
R41185 ASIG5V.n6209 ASIG5V.n6208 2.2505
R41186 ASIG5V.n6206 ASIG5V.n6015 2.2505
R41187 ASIG5V.n6204 ASIG5V.n6202 2.2505
R41188 ASIG5V.n6201 ASIG5V.n6017 2.2505
R41189 ASIG5V.n6200 ASIG5V.n6199 2.2505
R41190 ASIG5V.n6197 ASIG5V.n6018 2.2505
R41191 ASIG5V.n6195 ASIG5V.n6193 2.2505
R41192 ASIG5V.n6192 ASIG5V.n6020 2.2505
R41193 ASIG5V.n6191 ASIG5V.n6190 2.2505
R41194 ASIG5V.n6188 ASIG5V.n6021 2.2505
R41195 ASIG5V.n6186 ASIG5V.n6184 2.2505
R41196 ASIG5V.n6183 ASIG5V.n6023 2.2505
R41197 ASIG5V.n6182 ASIG5V.n6181 2.2505
R41198 ASIG5V.n6179 ASIG5V.n6024 2.2505
R41199 ASIG5V.n6177 ASIG5V.n6175 2.2505
R41200 ASIG5V.n6174 ASIG5V.n6026 2.2505
R41201 ASIG5V.n6173 ASIG5V.n6172 2.2505
R41202 ASIG5V.n6170 ASIG5V.n6027 2.2505
R41203 ASIG5V.n6168 ASIG5V.n6166 2.2505
R41204 ASIG5V.n6165 ASIG5V.n6029 2.2505
R41205 ASIG5V.n6164 ASIG5V.n6163 2.2505
R41206 ASIG5V.n6161 ASIG5V.n6030 2.2505
R41207 ASIG5V.n6159 ASIG5V.n6157 2.2505
R41208 ASIG5V.n6156 ASIG5V.n6032 2.2505
R41209 ASIG5V.n6155 ASIG5V.n6154 2.2505
R41210 ASIG5V.n6152 ASIG5V.n6033 2.2505
R41211 ASIG5V.n6150 ASIG5V.n6148 2.2505
R41212 ASIG5V.n6147 ASIG5V.n6035 2.2505
R41213 ASIG5V.n6146 ASIG5V.n6145 2.2505
R41214 ASIG5V.n6143 ASIG5V.n6036 2.2505
R41215 ASIG5V.n6141 ASIG5V.n6139 2.2505
R41216 ASIG5V.n6138 ASIG5V.n6038 2.2505
R41217 ASIG5V.n6137 ASIG5V.n6136 2.2505
R41218 ASIG5V.n6134 ASIG5V.n6039 2.2505
R41219 ASIG5V.n6132 ASIG5V.n6130 2.2505
R41220 ASIG5V.n6129 ASIG5V.n6041 2.2505
R41221 ASIG5V.n6128 ASIG5V.n6127 2.2505
R41222 ASIG5V.n6125 ASIG5V.n6042 2.2505
R41223 ASIG5V.n6123 ASIG5V.n6121 2.2505
R41224 ASIG5V.n6120 ASIG5V.n6044 2.2505
R41225 ASIG5V.n6119 ASIG5V.n6118 2.2505
R41226 ASIG5V.n6116 ASIG5V.n6045 2.2505
R41227 ASIG5V.n6114 ASIG5V.n6112 2.2505
R41228 ASIG5V.n6111 ASIG5V.n6047 2.2505
R41229 ASIG5V.n6110 ASIG5V.n6109 2.2505
R41230 ASIG5V.n6107 ASIG5V.n6048 2.2505
R41231 ASIG5V.n6105 ASIG5V.n6103 2.2505
R41232 ASIG5V.n6102 ASIG5V.n6050 2.2505
R41233 ASIG5V.n6101 ASIG5V.n6100 2.2505
R41234 ASIG5V.n6098 ASIG5V.n6051 2.2505
R41235 ASIG5V.n6096 ASIG5V.n6094 2.2505
R41236 ASIG5V.n6093 ASIG5V.n6053 2.2505
R41237 ASIG5V.n6092 ASIG5V.n6091 2.2505
R41238 ASIG5V.n6089 ASIG5V.n6054 2.2505
R41239 ASIG5V.n6087 ASIG5V.n6085 2.2505
R41240 ASIG5V.n6084 ASIG5V.n6056 2.2505
R41241 ASIG5V.n6083 ASIG5V.n6082 2.2505
R41242 ASIG5V.n6080 ASIG5V.n6057 2.2505
R41243 ASIG5V.n6078 ASIG5V.n6076 2.2505
R41244 ASIG5V.n6075 ASIG5V.n6059 2.2505
R41245 ASIG5V.n6074 ASIG5V.n6073 2.2505
R41246 ASIG5V.n6071 ASIG5V.n6060 2.2505
R41247 ASIG5V.n6069 ASIG5V.n6067 2.2505
R41248 ASIG5V.n6066 ASIG5V.n6062 2.2505
R41249 ASIG5V.n6065 ASIG5V.n6064 2.2505
R41250 ASIG5V.n6063 ASIG5V.n5956 2.2505
R41251 ASIG5V.n9394 ASIG5V.n5956 2.2505
R41252 ASIG5V.n6064 ASIG5V.n5955 2.2505
R41253 ASIG5V.n6062 ASIG5V.n6061 2.2505
R41254 ASIG5V.n6069 ASIG5V.n6068 2.2505
R41255 ASIG5V.n6071 ASIG5V.n6070 2.2505
R41256 ASIG5V.n6073 ASIG5V.n6072 2.2505
R41257 ASIG5V.n6059 ASIG5V.n6058 2.2505
R41258 ASIG5V.n6078 ASIG5V.n6077 2.2505
R41259 ASIG5V.n6080 ASIG5V.n6079 2.2505
R41260 ASIG5V.n6082 ASIG5V.n6081 2.2505
R41261 ASIG5V.n6056 ASIG5V.n6055 2.2505
R41262 ASIG5V.n6087 ASIG5V.n6086 2.2505
R41263 ASIG5V.n6089 ASIG5V.n6088 2.2505
R41264 ASIG5V.n6091 ASIG5V.n6090 2.2505
R41265 ASIG5V.n6053 ASIG5V.n6052 2.2505
R41266 ASIG5V.n6096 ASIG5V.n6095 2.2505
R41267 ASIG5V.n6098 ASIG5V.n6097 2.2505
R41268 ASIG5V.n6100 ASIG5V.n6099 2.2505
R41269 ASIG5V.n6050 ASIG5V.n6049 2.2505
R41270 ASIG5V.n6105 ASIG5V.n6104 2.2505
R41271 ASIG5V.n6107 ASIG5V.n6106 2.2505
R41272 ASIG5V.n6109 ASIG5V.n6108 2.2505
R41273 ASIG5V.n6047 ASIG5V.n6046 2.2505
R41274 ASIG5V.n6114 ASIG5V.n6113 2.2505
R41275 ASIG5V.n6116 ASIG5V.n6115 2.2505
R41276 ASIG5V.n6118 ASIG5V.n6117 2.2505
R41277 ASIG5V.n6044 ASIG5V.n6043 2.2505
R41278 ASIG5V.n6123 ASIG5V.n6122 2.2505
R41279 ASIG5V.n6125 ASIG5V.n6124 2.2505
R41280 ASIG5V.n6127 ASIG5V.n6126 2.2505
R41281 ASIG5V.n6041 ASIG5V.n6040 2.2505
R41282 ASIG5V.n6132 ASIG5V.n6131 2.2505
R41283 ASIG5V.n6134 ASIG5V.n6133 2.2505
R41284 ASIG5V.n6136 ASIG5V.n6135 2.2505
R41285 ASIG5V.n6038 ASIG5V.n6037 2.2505
R41286 ASIG5V.n6141 ASIG5V.n6140 2.2505
R41287 ASIG5V.n6143 ASIG5V.n6142 2.2505
R41288 ASIG5V.n6145 ASIG5V.n6144 2.2505
R41289 ASIG5V.n6035 ASIG5V.n6034 2.2505
R41290 ASIG5V.n6150 ASIG5V.n6149 2.2505
R41291 ASIG5V.n6152 ASIG5V.n6151 2.2505
R41292 ASIG5V.n6154 ASIG5V.n6153 2.2505
R41293 ASIG5V.n6032 ASIG5V.n6031 2.2505
R41294 ASIG5V.n6159 ASIG5V.n6158 2.2505
R41295 ASIG5V.n6161 ASIG5V.n6160 2.2505
R41296 ASIG5V.n6163 ASIG5V.n6162 2.2505
R41297 ASIG5V.n6029 ASIG5V.n6028 2.2505
R41298 ASIG5V.n6168 ASIG5V.n6167 2.2505
R41299 ASIG5V.n6170 ASIG5V.n6169 2.2505
R41300 ASIG5V.n6172 ASIG5V.n6171 2.2505
R41301 ASIG5V.n6026 ASIG5V.n6025 2.2505
R41302 ASIG5V.n6177 ASIG5V.n6176 2.2505
R41303 ASIG5V.n6179 ASIG5V.n6178 2.2505
R41304 ASIG5V.n6181 ASIG5V.n6180 2.2505
R41305 ASIG5V.n6023 ASIG5V.n6022 2.2505
R41306 ASIG5V.n6186 ASIG5V.n6185 2.2505
R41307 ASIG5V.n6188 ASIG5V.n6187 2.2505
R41308 ASIG5V.n6190 ASIG5V.n6189 2.2505
R41309 ASIG5V.n6020 ASIG5V.n6019 2.2505
R41310 ASIG5V.n6195 ASIG5V.n6194 2.2505
R41311 ASIG5V.n6197 ASIG5V.n6196 2.2505
R41312 ASIG5V.n6199 ASIG5V.n6198 2.2505
R41313 ASIG5V.n6017 ASIG5V.n6016 2.2505
R41314 ASIG5V.n6204 ASIG5V.n6203 2.2505
R41315 ASIG5V.n6206 ASIG5V.n6205 2.2505
R41316 ASIG5V.n6208 ASIG5V.n6207 2.2505
R41317 ASIG5V.n6014 ASIG5V.n6013 2.2505
R41318 ASIG5V.n6213 ASIG5V.n6212 2.2505
R41319 ASIG5V.n6215 ASIG5V.n6214 2.2505
R41320 ASIG5V.n6217 ASIG5V.n6216 2.2505
R41321 ASIG5V.n6011 ASIG5V.n6010 2.2505
R41322 ASIG5V.n6222 ASIG5V.n6221 2.2505
R41323 ASIG5V.n6224 ASIG5V.n6223 2.2505
R41324 ASIG5V.n6226 ASIG5V.n6225 2.2505
R41325 ASIG5V.n6008 ASIG5V.n6007 2.2505
R41326 ASIG5V.n6231 ASIG5V.n6230 2.2505
R41327 ASIG5V.n6233 ASIG5V.n6232 2.2505
R41328 ASIG5V.n6235 ASIG5V.n6234 2.2505
R41329 ASIG5V.n6005 ASIG5V.n6004 2.2505
R41330 ASIG5V.n6240 ASIG5V.n6239 2.2505
R41331 ASIG5V.n6242 ASIG5V.n6241 2.2505
R41332 ASIG5V.n6244 ASIG5V.n6243 2.2505
R41333 ASIG5V.n6002 ASIG5V.n6001 2.2505
R41334 ASIG5V.n9392 ASIG5V.n9391 2.2505
R41335 ASIG5V.n9377 ASIG5V.n9376 2.2505
R41336 ASIG5V.n9375 ASIG5V.n6354 2.2505
R41337 ASIG5V.n9374 ASIG5V.n9373 2.2505
R41338 ASIG5V.n9371 ASIG5V.n6355 2.2505
R41339 ASIG5V.n9369 ASIG5V.n9367 2.2505
R41340 ASIG5V.n9366 ASIG5V.n6357 2.2505
R41341 ASIG5V.n9365 ASIG5V.n9364 2.2505
R41342 ASIG5V.n9362 ASIG5V.n6358 2.2505
R41343 ASIG5V.n9360 ASIG5V.n9358 2.2505
R41344 ASIG5V.n9357 ASIG5V.n6360 2.2505
R41345 ASIG5V.n9356 ASIG5V.n9355 2.2505
R41346 ASIG5V.n9353 ASIG5V.n6361 2.2505
R41347 ASIG5V.n9351 ASIG5V.n9349 2.2505
R41348 ASIG5V.n9348 ASIG5V.n6363 2.2505
R41349 ASIG5V.n9347 ASIG5V.n9346 2.2505
R41350 ASIG5V.n9344 ASIG5V.n6364 2.2505
R41351 ASIG5V.n9342 ASIG5V.n9340 2.2505
R41352 ASIG5V.n9339 ASIG5V.n6366 2.2505
R41353 ASIG5V.n9338 ASIG5V.n9337 2.2505
R41354 ASIG5V.n9335 ASIG5V.n6367 2.2505
R41355 ASIG5V.n9333 ASIG5V.n9331 2.2505
R41356 ASIG5V.n9330 ASIG5V.n6369 2.2505
R41357 ASIG5V.n9329 ASIG5V.n9328 2.2505
R41358 ASIG5V.n9326 ASIG5V.n6370 2.2505
R41359 ASIG5V.n9324 ASIG5V.n9322 2.2505
R41360 ASIG5V.n9321 ASIG5V.n6372 2.2505
R41361 ASIG5V.n9320 ASIG5V.n9319 2.2505
R41362 ASIG5V.n9317 ASIG5V.n6373 2.2505
R41363 ASIG5V.n9315 ASIG5V.n9313 2.2505
R41364 ASIG5V.n9312 ASIG5V.n6375 2.2505
R41365 ASIG5V.n9311 ASIG5V.n9310 2.2505
R41366 ASIG5V.n9308 ASIG5V.n6376 2.2505
R41367 ASIG5V.n9306 ASIG5V.n9304 2.2505
R41368 ASIG5V.n9303 ASIG5V.n6378 2.2505
R41369 ASIG5V.n9302 ASIG5V.n9301 2.2505
R41370 ASIG5V.n9299 ASIG5V.n6379 2.2505
R41371 ASIG5V.n9297 ASIG5V.n9295 2.2505
R41372 ASIG5V.n9294 ASIG5V.n6381 2.2505
R41373 ASIG5V.n9293 ASIG5V.n9292 2.2505
R41374 ASIG5V.n9290 ASIG5V.n6382 2.2505
R41375 ASIG5V.n9288 ASIG5V.n9286 2.2505
R41376 ASIG5V.n9285 ASIG5V.n6384 2.2505
R41377 ASIG5V.n9284 ASIG5V.n9283 2.2505
R41378 ASIG5V.n9281 ASIG5V.n6385 2.2505
R41379 ASIG5V.n9279 ASIG5V.n9277 2.2505
R41380 ASIG5V.n9276 ASIG5V.n6387 2.2505
R41381 ASIG5V.n9275 ASIG5V.n9274 2.2505
R41382 ASIG5V.n9272 ASIG5V.n6388 2.2505
R41383 ASIG5V.n9270 ASIG5V.n9268 2.2505
R41384 ASIG5V.n9267 ASIG5V.n6390 2.2505
R41385 ASIG5V.n9266 ASIG5V.n9265 2.2505
R41386 ASIG5V.n9263 ASIG5V.n6391 2.2505
R41387 ASIG5V.n9261 ASIG5V.n9259 2.2505
R41388 ASIG5V.n9258 ASIG5V.n6393 2.2505
R41389 ASIG5V.n9257 ASIG5V.n9256 2.2505
R41390 ASIG5V.n9254 ASIG5V.n6394 2.2505
R41391 ASIG5V.n9252 ASIG5V.n9250 2.2505
R41392 ASIG5V.n9249 ASIG5V.n6396 2.2505
R41393 ASIG5V.n9248 ASIG5V.n9247 2.2505
R41394 ASIG5V.n9245 ASIG5V.n6397 2.2505
R41395 ASIG5V.n9243 ASIG5V.n9241 2.2505
R41396 ASIG5V.n9240 ASIG5V.n6399 2.2505
R41397 ASIG5V.n9239 ASIG5V.n9238 2.2505
R41398 ASIG5V.n9236 ASIG5V.n6400 2.2505
R41399 ASIG5V.n9234 ASIG5V.n9232 2.2505
R41400 ASIG5V.n9231 ASIG5V.n6402 2.2505
R41401 ASIG5V.n9230 ASIG5V.n9229 2.2505
R41402 ASIG5V.n9227 ASIG5V.n6403 2.2505
R41403 ASIG5V.n9225 ASIG5V.n9223 2.2505
R41404 ASIG5V.n9222 ASIG5V.n6405 2.2505
R41405 ASIG5V.n9221 ASIG5V.n9220 2.2505
R41406 ASIG5V.n9218 ASIG5V.n6406 2.2505
R41407 ASIG5V.n9216 ASIG5V.n9214 2.2505
R41408 ASIG5V.n9213 ASIG5V.n6408 2.2505
R41409 ASIG5V.n9212 ASIG5V.n9211 2.2505
R41410 ASIG5V.n9209 ASIG5V.n6409 2.2505
R41411 ASIG5V.n9207 ASIG5V.n9205 2.2505
R41412 ASIG5V.n9204 ASIG5V.n6411 2.2505
R41413 ASIG5V.n9203 ASIG5V.n9202 2.2505
R41414 ASIG5V.n9200 ASIG5V.n6412 2.2505
R41415 ASIG5V.n9198 ASIG5V.n9196 2.2505
R41416 ASIG5V.n9195 ASIG5V.n6414 2.2505
R41417 ASIG5V.n9194 ASIG5V.n9193 2.2505
R41418 ASIG5V.n9192 ASIG5V.n6309 2.2505
R41419 ASIG5V.n9380 ASIG5V.n6309 2.2505
R41420 ASIG5V.n9193 ASIG5V.n6307 2.2505
R41421 ASIG5V.n6414 ASIG5V.n6413 2.2505
R41422 ASIG5V.n9198 ASIG5V.n9197 2.2505
R41423 ASIG5V.n9200 ASIG5V.n9199 2.2505
R41424 ASIG5V.n9202 ASIG5V.n9201 2.2505
R41425 ASIG5V.n6411 ASIG5V.n6410 2.2505
R41426 ASIG5V.n9207 ASIG5V.n9206 2.2505
R41427 ASIG5V.n9209 ASIG5V.n9208 2.2505
R41428 ASIG5V.n9211 ASIG5V.n9210 2.2505
R41429 ASIG5V.n6408 ASIG5V.n6407 2.2505
R41430 ASIG5V.n9216 ASIG5V.n9215 2.2505
R41431 ASIG5V.n9218 ASIG5V.n9217 2.2505
R41432 ASIG5V.n9220 ASIG5V.n9219 2.2505
R41433 ASIG5V.n6405 ASIG5V.n6404 2.2505
R41434 ASIG5V.n9225 ASIG5V.n9224 2.2505
R41435 ASIG5V.n9227 ASIG5V.n9226 2.2505
R41436 ASIG5V.n9229 ASIG5V.n9228 2.2505
R41437 ASIG5V.n6402 ASIG5V.n6401 2.2505
R41438 ASIG5V.n9234 ASIG5V.n9233 2.2505
R41439 ASIG5V.n9236 ASIG5V.n9235 2.2505
R41440 ASIG5V.n9238 ASIG5V.n9237 2.2505
R41441 ASIG5V.n6399 ASIG5V.n6398 2.2505
R41442 ASIG5V.n9243 ASIG5V.n9242 2.2505
R41443 ASIG5V.n9245 ASIG5V.n9244 2.2505
R41444 ASIG5V.n9247 ASIG5V.n9246 2.2505
R41445 ASIG5V.n6396 ASIG5V.n6395 2.2505
R41446 ASIG5V.n9252 ASIG5V.n9251 2.2505
R41447 ASIG5V.n9254 ASIG5V.n9253 2.2505
R41448 ASIG5V.n9256 ASIG5V.n9255 2.2505
R41449 ASIG5V.n6393 ASIG5V.n6392 2.2505
R41450 ASIG5V.n9261 ASIG5V.n9260 2.2505
R41451 ASIG5V.n9263 ASIG5V.n9262 2.2505
R41452 ASIG5V.n9265 ASIG5V.n9264 2.2505
R41453 ASIG5V.n6390 ASIG5V.n6389 2.2505
R41454 ASIG5V.n9270 ASIG5V.n9269 2.2505
R41455 ASIG5V.n9272 ASIG5V.n9271 2.2505
R41456 ASIG5V.n9274 ASIG5V.n9273 2.2505
R41457 ASIG5V.n6387 ASIG5V.n6386 2.2505
R41458 ASIG5V.n9279 ASIG5V.n9278 2.2505
R41459 ASIG5V.n9281 ASIG5V.n9280 2.2505
R41460 ASIG5V.n9283 ASIG5V.n9282 2.2505
R41461 ASIG5V.n6384 ASIG5V.n6383 2.2505
R41462 ASIG5V.n9288 ASIG5V.n9287 2.2505
R41463 ASIG5V.n9290 ASIG5V.n9289 2.2505
R41464 ASIG5V.n9292 ASIG5V.n9291 2.2505
R41465 ASIG5V.n6381 ASIG5V.n6380 2.2505
R41466 ASIG5V.n9297 ASIG5V.n9296 2.2505
R41467 ASIG5V.n9299 ASIG5V.n9298 2.2505
R41468 ASIG5V.n9301 ASIG5V.n9300 2.2505
R41469 ASIG5V.n6378 ASIG5V.n6377 2.2505
R41470 ASIG5V.n9306 ASIG5V.n9305 2.2505
R41471 ASIG5V.n9308 ASIG5V.n9307 2.2505
R41472 ASIG5V.n9310 ASIG5V.n9309 2.2505
R41473 ASIG5V.n6375 ASIG5V.n6374 2.2505
R41474 ASIG5V.n9315 ASIG5V.n9314 2.2505
R41475 ASIG5V.n9317 ASIG5V.n9316 2.2505
R41476 ASIG5V.n9319 ASIG5V.n9318 2.2505
R41477 ASIG5V.n6372 ASIG5V.n6371 2.2505
R41478 ASIG5V.n9324 ASIG5V.n9323 2.2505
R41479 ASIG5V.n9326 ASIG5V.n9325 2.2505
R41480 ASIG5V.n9328 ASIG5V.n9327 2.2505
R41481 ASIG5V.n6369 ASIG5V.n6368 2.2505
R41482 ASIG5V.n9333 ASIG5V.n9332 2.2505
R41483 ASIG5V.n9335 ASIG5V.n9334 2.2505
R41484 ASIG5V.n9337 ASIG5V.n9336 2.2505
R41485 ASIG5V.n6366 ASIG5V.n6365 2.2505
R41486 ASIG5V.n9342 ASIG5V.n9341 2.2505
R41487 ASIG5V.n9344 ASIG5V.n9343 2.2505
R41488 ASIG5V.n9346 ASIG5V.n9345 2.2505
R41489 ASIG5V.n6363 ASIG5V.n6362 2.2505
R41490 ASIG5V.n9351 ASIG5V.n9350 2.2505
R41491 ASIG5V.n9353 ASIG5V.n9352 2.2505
R41492 ASIG5V.n9355 ASIG5V.n9354 2.2505
R41493 ASIG5V.n6360 ASIG5V.n6359 2.2505
R41494 ASIG5V.n9360 ASIG5V.n9359 2.2505
R41495 ASIG5V.n9362 ASIG5V.n9361 2.2505
R41496 ASIG5V.n9364 ASIG5V.n9363 2.2505
R41497 ASIG5V.n6357 ASIG5V.n6356 2.2505
R41498 ASIG5V.n9369 ASIG5V.n9368 2.2505
R41499 ASIG5V.n9371 ASIG5V.n9370 2.2505
R41500 ASIG5V.n9373 ASIG5V.n9372 2.2505
R41501 ASIG5V.n6354 ASIG5V.n6353 2.2505
R41502 ASIG5V.n9378 ASIG5V.n9377 2.2505
R41503 ASIG5V.n6489 ASIG5V.n6441 2.2505
R41504 ASIG5V.n9172 ASIG5V.n9171 2.2505
R41505 ASIG5V.n9170 ASIG5V.n6490 2.2505
R41506 ASIG5V.n9169 ASIG5V.n9168 2.2505
R41507 ASIG5V.n9164 ASIG5V.n6491 2.2505
R41508 ASIG5V.n9160 ASIG5V.n9159 2.2505
R41509 ASIG5V.n9158 ASIG5V.n6492 2.2505
R41510 ASIG5V.n9157 ASIG5V.n9156 2.2505
R41511 ASIG5V.n9152 ASIG5V.n6493 2.2505
R41512 ASIG5V.n9148 ASIG5V.n9147 2.2505
R41513 ASIG5V.n9146 ASIG5V.n6494 2.2505
R41514 ASIG5V.n9145 ASIG5V.n9144 2.2505
R41515 ASIG5V.n9140 ASIG5V.n6495 2.2505
R41516 ASIG5V.n9136 ASIG5V.n9135 2.2505
R41517 ASIG5V.n9134 ASIG5V.n6496 2.2505
R41518 ASIG5V.n9133 ASIG5V.n9132 2.2505
R41519 ASIG5V.n9128 ASIG5V.n6497 2.2505
R41520 ASIG5V.n9124 ASIG5V.n9123 2.2505
R41521 ASIG5V.n9122 ASIG5V.n6498 2.2505
R41522 ASIG5V.n9121 ASIG5V.n9120 2.2505
R41523 ASIG5V.n9116 ASIG5V.n6499 2.2505
R41524 ASIG5V.n9112 ASIG5V.n9111 2.2505
R41525 ASIG5V.n9110 ASIG5V.n6500 2.2505
R41526 ASIG5V.n9109 ASIG5V.n9108 2.2505
R41527 ASIG5V.n9104 ASIG5V.n6501 2.2505
R41528 ASIG5V.n9100 ASIG5V.n9099 2.2505
R41529 ASIG5V.n9098 ASIG5V.n6502 2.2505
R41530 ASIG5V.n9097 ASIG5V.n9096 2.2505
R41531 ASIG5V.n9092 ASIG5V.n6503 2.2505
R41532 ASIG5V.n9088 ASIG5V.n9087 2.2505
R41533 ASIG5V.n9086 ASIG5V.n6504 2.2505
R41534 ASIG5V.n9085 ASIG5V.n9084 2.2505
R41535 ASIG5V.n9080 ASIG5V.n6505 2.2505
R41536 ASIG5V.n9076 ASIG5V.n9075 2.2505
R41537 ASIG5V.n9074 ASIG5V.n6506 2.2505
R41538 ASIG5V.n9073 ASIG5V.n9072 2.2505
R41539 ASIG5V.n9068 ASIG5V.n6507 2.2505
R41540 ASIG5V.n9064 ASIG5V.n9063 2.2505
R41541 ASIG5V.n9062 ASIG5V.n6508 2.2505
R41542 ASIG5V.n9061 ASIG5V.n9060 2.2505
R41543 ASIG5V.n9056 ASIG5V.n6509 2.2505
R41544 ASIG5V.n9052 ASIG5V.n9051 2.2505
R41545 ASIG5V.n9050 ASIG5V.n6510 2.2505
R41546 ASIG5V.n9049 ASIG5V.n9048 2.2505
R41547 ASIG5V.n9044 ASIG5V.n6511 2.2505
R41548 ASIG5V.n9040 ASIG5V.n9039 2.2505
R41549 ASIG5V.n9038 ASIG5V.n6512 2.2505
R41550 ASIG5V.n9037 ASIG5V.n9036 2.2505
R41551 ASIG5V.n9032 ASIG5V.n6513 2.2505
R41552 ASIG5V.n9028 ASIG5V.n9027 2.2505
R41553 ASIG5V.n9026 ASIG5V.n6514 2.2505
R41554 ASIG5V.n9025 ASIG5V.n9024 2.2505
R41555 ASIG5V.n9020 ASIG5V.n6515 2.2505
R41556 ASIG5V.n9016 ASIG5V.n9015 2.2505
R41557 ASIG5V.n9014 ASIG5V.n6516 2.2505
R41558 ASIG5V.n9013 ASIG5V.n9012 2.2505
R41559 ASIG5V.n9008 ASIG5V.n6517 2.2505
R41560 ASIG5V.n9004 ASIG5V.n9003 2.2505
R41561 ASIG5V.n9002 ASIG5V.n6518 2.2505
R41562 ASIG5V.n9001 ASIG5V.n9000 2.2505
R41563 ASIG5V.n8996 ASIG5V.n6519 2.2505
R41564 ASIG5V.n8992 ASIG5V.n8991 2.2505
R41565 ASIG5V.n8990 ASIG5V.n6520 2.2505
R41566 ASIG5V.n8989 ASIG5V.n8988 2.2505
R41567 ASIG5V.n8984 ASIG5V.n6521 2.2505
R41568 ASIG5V.n8980 ASIG5V.n8979 2.2505
R41569 ASIG5V.n8978 ASIG5V.n6522 2.2505
R41570 ASIG5V.n8977 ASIG5V.n8976 2.2505
R41571 ASIG5V.n8972 ASIG5V.n6523 2.2505
R41572 ASIG5V.n8968 ASIG5V.n8967 2.2505
R41573 ASIG5V.n8966 ASIG5V.n6524 2.2505
R41574 ASIG5V.n8965 ASIG5V.n8964 2.2505
R41575 ASIG5V.n8960 ASIG5V.n6525 2.2505
R41576 ASIG5V.n8956 ASIG5V.n8955 2.2505
R41577 ASIG5V.n8954 ASIG5V.n6526 2.2505
R41578 ASIG5V.n8953 ASIG5V.n8952 2.2505
R41579 ASIG5V.n8948 ASIG5V.n6527 2.2505
R41580 ASIG5V.n8944 ASIG5V.n8943 2.2505
R41581 ASIG5V.n8942 ASIG5V.n6528 2.2505
R41582 ASIG5V.n8941 ASIG5V.n8940 2.2505
R41583 ASIG5V.n8936 ASIG5V.n6529 2.2505
R41584 ASIG5V.n8932 ASIG5V.n8931 2.2505
R41585 ASIG5V.n8930 ASIG5V.n6532 2.2505
R41586 ASIG5V.n8929 ASIG5V.n8928 2.2505
R41587 ASIG5V.n8928 ASIG5V.n6487 2.2505
R41588 ASIG5V.n6532 ASIG5V.n6531 2.2505
R41589 ASIG5V.n8933 ASIG5V.n8932 2.2505
R41590 ASIG5V.n8936 ASIG5V.n8935 2.2505
R41591 ASIG5V.n8940 ASIG5V.n8939 2.2505
R41592 ASIG5V.n8937 ASIG5V.n6528 2.2505
R41593 ASIG5V.n8945 ASIG5V.n8944 2.2505
R41594 ASIG5V.n8948 ASIG5V.n8947 2.2505
R41595 ASIG5V.n8952 ASIG5V.n8951 2.2505
R41596 ASIG5V.n8949 ASIG5V.n6526 2.2505
R41597 ASIG5V.n8957 ASIG5V.n8956 2.2505
R41598 ASIG5V.n8960 ASIG5V.n8959 2.2505
R41599 ASIG5V.n8964 ASIG5V.n8963 2.2505
R41600 ASIG5V.n8961 ASIG5V.n6524 2.2505
R41601 ASIG5V.n8969 ASIG5V.n8968 2.2505
R41602 ASIG5V.n8972 ASIG5V.n8971 2.2505
R41603 ASIG5V.n8976 ASIG5V.n8975 2.2505
R41604 ASIG5V.n8973 ASIG5V.n6522 2.2505
R41605 ASIG5V.n8981 ASIG5V.n8980 2.2505
R41606 ASIG5V.n8984 ASIG5V.n8983 2.2505
R41607 ASIG5V.n8988 ASIG5V.n8987 2.2505
R41608 ASIG5V.n8985 ASIG5V.n6520 2.2505
R41609 ASIG5V.n8993 ASIG5V.n8992 2.2505
R41610 ASIG5V.n8996 ASIG5V.n8995 2.2505
R41611 ASIG5V.n9000 ASIG5V.n8999 2.2505
R41612 ASIG5V.n8997 ASIG5V.n6518 2.2505
R41613 ASIG5V.n9005 ASIG5V.n9004 2.2505
R41614 ASIG5V.n9008 ASIG5V.n9007 2.2505
R41615 ASIG5V.n9012 ASIG5V.n9011 2.2505
R41616 ASIG5V.n9009 ASIG5V.n6516 2.2505
R41617 ASIG5V.n9017 ASIG5V.n9016 2.2505
R41618 ASIG5V.n9020 ASIG5V.n9019 2.2505
R41619 ASIG5V.n9024 ASIG5V.n9023 2.2505
R41620 ASIG5V.n9021 ASIG5V.n6514 2.2505
R41621 ASIG5V.n9029 ASIG5V.n9028 2.2505
R41622 ASIG5V.n9032 ASIG5V.n9031 2.2505
R41623 ASIG5V.n9036 ASIG5V.n9035 2.2505
R41624 ASIG5V.n9033 ASIG5V.n6512 2.2505
R41625 ASIG5V.n9041 ASIG5V.n9040 2.2505
R41626 ASIG5V.n9044 ASIG5V.n9043 2.2505
R41627 ASIG5V.n9048 ASIG5V.n9047 2.2505
R41628 ASIG5V.n9045 ASIG5V.n6510 2.2505
R41629 ASIG5V.n9053 ASIG5V.n9052 2.2505
R41630 ASIG5V.n9056 ASIG5V.n9055 2.2505
R41631 ASIG5V.n9060 ASIG5V.n9059 2.2505
R41632 ASIG5V.n9057 ASIG5V.n6508 2.2505
R41633 ASIG5V.n9065 ASIG5V.n9064 2.2505
R41634 ASIG5V.n9068 ASIG5V.n9067 2.2505
R41635 ASIG5V.n9072 ASIG5V.n9071 2.2505
R41636 ASIG5V.n9069 ASIG5V.n6506 2.2505
R41637 ASIG5V.n9077 ASIG5V.n9076 2.2505
R41638 ASIG5V.n9080 ASIG5V.n9079 2.2505
R41639 ASIG5V.n9084 ASIG5V.n9083 2.2505
R41640 ASIG5V.n9081 ASIG5V.n6504 2.2505
R41641 ASIG5V.n9089 ASIG5V.n9088 2.2505
R41642 ASIG5V.n9092 ASIG5V.n9091 2.2505
R41643 ASIG5V.n9096 ASIG5V.n9095 2.2505
R41644 ASIG5V.n9093 ASIG5V.n6502 2.2505
R41645 ASIG5V.n9101 ASIG5V.n9100 2.2505
R41646 ASIG5V.n9104 ASIG5V.n9103 2.2505
R41647 ASIG5V.n9108 ASIG5V.n9107 2.2505
R41648 ASIG5V.n9105 ASIG5V.n6500 2.2505
R41649 ASIG5V.n9113 ASIG5V.n9112 2.2505
R41650 ASIG5V.n9116 ASIG5V.n9115 2.2505
R41651 ASIG5V.n9120 ASIG5V.n9119 2.2505
R41652 ASIG5V.n9117 ASIG5V.n6498 2.2505
R41653 ASIG5V.n9125 ASIG5V.n9124 2.2505
R41654 ASIG5V.n9128 ASIG5V.n9127 2.2505
R41655 ASIG5V.n9132 ASIG5V.n9131 2.2505
R41656 ASIG5V.n9129 ASIG5V.n6496 2.2505
R41657 ASIG5V.n9137 ASIG5V.n9136 2.2505
R41658 ASIG5V.n9140 ASIG5V.n9139 2.2505
R41659 ASIG5V.n9144 ASIG5V.n9143 2.2505
R41660 ASIG5V.n9141 ASIG5V.n6494 2.2505
R41661 ASIG5V.n9149 ASIG5V.n9148 2.2505
R41662 ASIG5V.n9152 ASIG5V.n9151 2.2505
R41663 ASIG5V.n9156 ASIG5V.n9155 2.2505
R41664 ASIG5V.n9153 ASIG5V.n6492 2.2505
R41665 ASIG5V.n9161 ASIG5V.n9160 2.2505
R41666 ASIG5V.n9164 ASIG5V.n9163 2.2505
R41667 ASIG5V.n9168 ASIG5V.n9167 2.2505
R41668 ASIG5V.n9165 ASIG5V.n6490 2.2505
R41669 ASIG5V.n9173 ASIG5V.n9172 2.2505
R41670 ASIG5V.n9175 ASIG5V.n6489 2.2505
R41671 ASIG5V.n8914 ASIG5V.n6880 2.2505
R41672 ASIG5V.n6879 ASIG5V.n6635 2.2505
R41673 ASIG5V.n6878 ASIG5V.n6877 2.2505
R41674 ASIG5V.n6875 ASIG5V.n6636 2.2505
R41675 ASIG5V.n6873 ASIG5V.n6871 2.2505
R41676 ASIG5V.n6870 ASIG5V.n6638 2.2505
R41677 ASIG5V.n6869 ASIG5V.n6868 2.2505
R41678 ASIG5V.n6866 ASIG5V.n6639 2.2505
R41679 ASIG5V.n6864 ASIG5V.n6862 2.2505
R41680 ASIG5V.n6861 ASIG5V.n6641 2.2505
R41681 ASIG5V.n6860 ASIG5V.n6859 2.2505
R41682 ASIG5V.n6857 ASIG5V.n6642 2.2505
R41683 ASIG5V.n6855 ASIG5V.n6853 2.2505
R41684 ASIG5V.n6852 ASIG5V.n6644 2.2505
R41685 ASIG5V.n6851 ASIG5V.n6850 2.2505
R41686 ASIG5V.n6848 ASIG5V.n6645 2.2505
R41687 ASIG5V.n6846 ASIG5V.n6844 2.2505
R41688 ASIG5V.n6843 ASIG5V.n6647 2.2505
R41689 ASIG5V.n6842 ASIG5V.n6841 2.2505
R41690 ASIG5V.n6839 ASIG5V.n6648 2.2505
R41691 ASIG5V.n6837 ASIG5V.n6835 2.2505
R41692 ASIG5V.n6834 ASIG5V.n6650 2.2505
R41693 ASIG5V.n6833 ASIG5V.n6832 2.2505
R41694 ASIG5V.n6830 ASIG5V.n6651 2.2505
R41695 ASIG5V.n6828 ASIG5V.n6826 2.2505
R41696 ASIG5V.n6825 ASIG5V.n6653 2.2505
R41697 ASIG5V.n6824 ASIG5V.n6823 2.2505
R41698 ASIG5V.n6821 ASIG5V.n6654 2.2505
R41699 ASIG5V.n6819 ASIG5V.n6817 2.2505
R41700 ASIG5V.n6816 ASIG5V.n6656 2.2505
R41701 ASIG5V.n6815 ASIG5V.n6814 2.2505
R41702 ASIG5V.n6812 ASIG5V.n6657 2.2505
R41703 ASIG5V.n6810 ASIG5V.n6808 2.2505
R41704 ASIG5V.n6807 ASIG5V.n6659 2.2505
R41705 ASIG5V.n6806 ASIG5V.n6805 2.2505
R41706 ASIG5V.n6803 ASIG5V.n6660 2.2505
R41707 ASIG5V.n6801 ASIG5V.n6799 2.2505
R41708 ASIG5V.n6798 ASIG5V.n6662 2.2505
R41709 ASIG5V.n6797 ASIG5V.n6796 2.2505
R41710 ASIG5V.n6794 ASIG5V.n6663 2.2505
R41711 ASIG5V.n6792 ASIG5V.n6790 2.2505
R41712 ASIG5V.n6789 ASIG5V.n6665 2.2505
R41713 ASIG5V.n6788 ASIG5V.n6787 2.2505
R41714 ASIG5V.n6785 ASIG5V.n6666 2.2505
R41715 ASIG5V.n6783 ASIG5V.n6781 2.2505
R41716 ASIG5V.n6780 ASIG5V.n6668 2.2505
R41717 ASIG5V.n6779 ASIG5V.n6778 2.2505
R41718 ASIG5V.n6776 ASIG5V.n6669 2.2505
R41719 ASIG5V.n6774 ASIG5V.n6772 2.2505
R41720 ASIG5V.n6771 ASIG5V.n6671 2.2505
R41721 ASIG5V.n6770 ASIG5V.n6769 2.2505
R41722 ASIG5V.n6767 ASIG5V.n6672 2.2505
R41723 ASIG5V.n6765 ASIG5V.n6763 2.2505
R41724 ASIG5V.n6762 ASIG5V.n6674 2.2505
R41725 ASIG5V.n6761 ASIG5V.n6760 2.2505
R41726 ASIG5V.n6758 ASIG5V.n6675 2.2505
R41727 ASIG5V.n6756 ASIG5V.n6754 2.2505
R41728 ASIG5V.n6753 ASIG5V.n6677 2.2505
R41729 ASIG5V.n6752 ASIG5V.n6751 2.2505
R41730 ASIG5V.n6749 ASIG5V.n6678 2.2505
R41731 ASIG5V.n6747 ASIG5V.n6745 2.2505
R41732 ASIG5V.n6744 ASIG5V.n6680 2.2505
R41733 ASIG5V.n6743 ASIG5V.n6742 2.2505
R41734 ASIG5V.n6740 ASIG5V.n6681 2.2505
R41735 ASIG5V.n6738 ASIG5V.n6736 2.2505
R41736 ASIG5V.n6735 ASIG5V.n6683 2.2505
R41737 ASIG5V.n6734 ASIG5V.n6733 2.2505
R41738 ASIG5V.n6731 ASIG5V.n6684 2.2505
R41739 ASIG5V.n6729 ASIG5V.n6727 2.2505
R41740 ASIG5V.n6726 ASIG5V.n6686 2.2505
R41741 ASIG5V.n6725 ASIG5V.n6724 2.2505
R41742 ASIG5V.n6722 ASIG5V.n6687 2.2505
R41743 ASIG5V.n6720 ASIG5V.n6718 2.2505
R41744 ASIG5V.n6717 ASIG5V.n6689 2.2505
R41745 ASIG5V.n6716 ASIG5V.n6715 2.2505
R41746 ASIG5V.n6713 ASIG5V.n6690 2.2505
R41747 ASIG5V.n6711 ASIG5V.n6709 2.2505
R41748 ASIG5V.n6708 ASIG5V.n6692 2.2505
R41749 ASIG5V.n6707 ASIG5V.n6706 2.2505
R41750 ASIG5V.n6704 ASIG5V.n6693 2.2505
R41751 ASIG5V.n6702 ASIG5V.n6700 2.2505
R41752 ASIG5V.n6699 ASIG5V.n6695 2.2505
R41753 ASIG5V.n6698 ASIG5V.n6697 2.2505
R41754 ASIG5V.n6696 ASIG5V.n6589 2.2505
R41755 ASIG5V.n8917 ASIG5V.n6589 2.2505
R41756 ASIG5V.n6697 ASIG5V.n6588 2.2505
R41757 ASIG5V.n6695 ASIG5V.n6694 2.2505
R41758 ASIG5V.n6702 ASIG5V.n6701 2.2505
R41759 ASIG5V.n6704 ASIG5V.n6703 2.2505
R41760 ASIG5V.n6706 ASIG5V.n6705 2.2505
R41761 ASIG5V.n6692 ASIG5V.n6691 2.2505
R41762 ASIG5V.n6711 ASIG5V.n6710 2.2505
R41763 ASIG5V.n6713 ASIG5V.n6712 2.2505
R41764 ASIG5V.n6715 ASIG5V.n6714 2.2505
R41765 ASIG5V.n6689 ASIG5V.n6688 2.2505
R41766 ASIG5V.n6720 ASIG5V.n6719 2.2505
R41767 ASIG5V.n6722 ASIG5V.n6721 2.2505
R41768 ASIG5V.n6724 ASIG5V.n6723 2.2505
R41769 ASIG5V.n6686 ASIG5V.n6685 2.2505
R41770 ASIG5V.n6729 ASIG5V.n6728 2.2505
R41771 ASIG5V.n6731 ASIG5V.n6730 2.2505
R41772 ASIG5V.n6733 ASIG5V.n6732 2.2505
R41773 ASIG5V.n6683 ASIG5V.n6682 2.2505
R41774 ASIG5V.n6738 ASIG5V.n6737 2.2505
R41775 ASIG5V.n6740 ASIG5V.n6739 2.2505
R41776 ASIG5V.n6742 ASIG5V.n6741 2.2505
R41777 ASIG5V.n6680 ASIG5V.n6679 2.2505
R41778 ASIG5V.n6747 ASIG5V.n6746 2.2505
R41779 ASIG5V.n6749 ASIG5V.n6748 2.2505
R41780 ASIG5V.n6751 ASIG5V.n6750 2.2505
R41781 ASIG5V.n6677 ASIG5V.n6676 2.2505
R41782 ASIG5V.n6756 ASIG5V.n6755 2.2505
R41783 ASIG5V.n6758 ASIG5V.n6757 2.2505
R41784 ASIG5V.n6760 ASIG5V.n6759 2.2505
R41785 ASIG5V.n6674 ASIG5V.n6673 2.2505
R41786 ASIG5V.n6765 ASIG5V.n6764 2.2505
R41787 ASIG5V.n6767 ASIG5V.n6766 2.2505
R41788 ASIG5V.n6769 ASIG5V.n6768 2.2505
R41789 ASIG5V.n6671 ASIG5V.n6670 2.2505
R41790 ASIG5V.n6774 ASIG5V.n6773 2.2505
R41791 ASIG5V.n6776 ASIG5V.n6775 2.2505
R41792 ASIG5V.n6778 ASIG5V.n6777 2.2505
R41793 ASIG5V.n6668 ASIG5V.n6667 2.2505
R41794 ASIG5V.n6783 ASIG5V.n6782 2.2505
R41795 ASIG5V.n6785 ASIG5V.n6784 2.2505
R41796 ASIG5V.n6787 ASIG5V.n6786 2.2505
R41797 ASIG5V.n6665 ASIG5V.n6664 2.2505
R41798 ASIG5V.n6792 ASIG5V.n6791 2.2505
R41799 ASIG5V.n6794 ASIG5V.n6793 2.2505
R41800 ASIG5V.n6796 ASIG5V.n6795 2.2505
R41801 ASIG5V.n6662 ASIG5V.n6661 2.2505
R41802 ASIG5V.n6801 ASIG5V.n6800 2.2505
R41803 ASIG5V.n6803 ASIG5V.n6802 2.2505
R41804 ASIG5V.n6805 ASIG5V.n6804 2.2505
R41805 ASIG5V.n6659 ASIG5V.n6658 2.2505
R41806 ASIG5V.n6810 ASIG5V.n6809 2.2505
R41807 ASIG5V.n6812 ASIG5V.n6811 2.2505
R41808 ASIG5V.n6814 ASIG5V.n6813 2.2505
R41809 ASIG5V.n6656 ASIG5V.n6655 2.2505
R41810 ASIG5V.n6819 ASIG5V.n6818 2.2505
R41811 ASIG5V.n6821 ASIG5V.n6820 2.2505
R41812 ASIG5V.n6823 ASIG5V.n6822 2.2505
R41813 ASIG5V.n6653 ASIG5V.n6652 2.2505
R41814 ASIG5V.n6828 ASIG5V.n6827 2.2505
R41815 ASIG5V.n6830 ASIG5V.n6829 2.2505
R41816 ASIG5V.n6832 ASIG5V.n6831 2.2505
R41817 ASIG5V.n6650 ASIG5V.n6649 2.2505
R41818 ASIG5V.n6837 ASIG5V.n6836 2.2505
R41819 ASIG5V.n6839 ASIG5V.n6838 2.2505
R41820 ASIG5V.n6841 ASIG5V.n6840 2.2505
R41821 ASIG5V.n6647 ASIG5V.n6646 2.2505
R41822 ASIG5V.n6846 ASIG5V.n6845 2.2505
R41823 ASIG5V.n6848 ASIG5V.n6847 2.2505
R41824 ASIG5V.n6850 ASIG5V.n6849 2.2505
R41825 ASIG5V.n6644 ASIG5V.n6643 2.2505
R41826 ASIG5V.n6855 ASIG5V.n6854 2.2505
R41827 ASIG5V.n6857 ASIG5V.n6856 2.2505
R41828 ASIG5V.n6859 ASIG5V.n6858 2.2505
R41829 ASIG5V.n6641 ASIG5V.n6640 2.2505
R41830 ASIG5V.n6864 ASIG5V.n6863 2.2505
R41831 ASIG5V.n6866 ASIG5V.n6865 2.2505
R41832 ASIG5V.n6868 ASIG5V.n6867 2.2505
R41833 ASIG5V.n6638 ASIG5V.n6637 2.2505
R41834 ASIG5V.n6873 ASIG5V.n6872 2.2505
R41835 ASIG5V.n6875 ASIG5V.n6874 2.2505
R41836 ASIG5V.n6877 ASIG5V.n6876 2.2505
R41837 ASIG5V.n6635 ASIG5V.n6634 2.2505
R41838 ASIG5V.n8915 ASIG5V.n8914 2.2505
R41839 ASIG5V.n7022 ASIG5V.n7021 2.2505
R41840 ASIG5V.n7024 ASIG5V.n7023 2.2505
R41841 ASIG5V.n7016 ASIG5V.n7015 2.2505
R41842 ASIG5V.n7031 ASIG5V.n7030 2.2505
R41843 ASIG5V.n7032 ASIG5V.n7014 2.2505
R41844 ASIG5V.n7034 ASIG5V.n7033 2.2505
R41845 ASIG5V.n7010 ASIG5V.n7009 2.2505
R41846 ASIG5V.n7041 ASIG5V.n7040 2.2505
R41847 ASIG5V.n7042 ASIG5V.n7008 2.2505
R41848 ASIG5V.n7044 ASIG5V.n7043 2.2505
R41849 ASIG5V.n7004 ASIG5V.n7003 2.2505
R41850 ASIG5V.n7051 ASIG5V.n7050 2.2505
R41851 ASIG5V.n7052 ASIG5V.n7002 2.2505
R41852 ASIG5V.n7054 ASIG5V.n7053 2.2505
R41853 ASIG5V.n6998 ASIG5V.n6997 2.2505
R41854 ASIG5V.n7061 ASIG5V.n7060 2.2505
R41855 ASIG5V.n7062 ASIG5V.n6996 2.2505
R41856 ASIG5V.n7064 ASIG5V.n7063 2.2505
R41857 ASIG5V.n6992 ASIG5V.n6991 2.2505
R41858 ASIG5V.n7071 ASIG5V.n7070 2.2505
R41859 ASIG5V.n7072 ASIG5V.n6990 2.2505
R41860 ASIG5V.n7074 ASIG5V.n7073 2.2505
R41861 ASIG5V.n6986 ASIG5V.n6985 2.2505
R41862 ASIG5V.n7081 ASIG5V.n7080 2.2505
R41863 ASIG5V.n7082 ASIG5V.n6984 2.2505
R41864 ASIG5V.n7084 ASIG5V.n7083 2.2505
R41865 ASIG5V.n6980 ASIG5V.n6979 2.2505
R41866 ASIG5V.n7091 ASIG5V.n7090 2.2505
R41867 ASIG5V.n7092 ASIG5V.n6978 2.2505
R41868 ASIG5V.n7094 ASIG5V.n7093 2.2505
R41869 ASIG5V.n6974 ASIG5V.n6973 2.2505
R41870 ASIG5V.n7101 ASIG5V.n7100 2.2505
R41871 ASIG5V.n7102 ASIG5V.n6972 2.2505
R41872 ASIG5V.n7104 ASIG5V.n7103 2.2505
R41873 ASIG5V.n6968 ASIG5V.n6967 2.2505
R41874 ASIG5V.n7111 ASIG5V.n7110 2.2505
R41875 ASIG5V.n7112 ASIG5V.n6966 2.2505
R41876 ASIG5V.n7114 ASIG5V.n7113 2.2505
R41877 ASIG5V.n6962 ASIG5V.n6961 2.2505
R41878 ASIG5V.n7121 ASIG5V.n7120 2.2505
R41879 ASIG5V.n7122 ASIG5V.n6960 2.2505
R41880 ASIG5V.n7124 ASIG5V.n7123 2.2505
R41881 ASIG5V.n6956 ASIG5V.n6955 2.2505
R41882 ASIG5V.n7131 ASIG5V.n7130 2.2505
R41883 ASIG5V.n7132 ASIG5V.n6954 2.2505
R41884 ASIG5V.n7134 ASIG5V.n7133 2.2505
R41885 ASIG5V.n6950 ASIG5V.n6949 2.2505
R41886 ASIG5V.n7141 ASIG5V.n7140 2.2505
R41887 ASIG5V.n7142 ASIG5V.n6948 2.2505
R41888 ASIG5V.n7144 ASIG5V.n7143 2.2505
R41889 ASIG5V.n6944 ASIG5V.n6943 2.2505
R41890 ASIG5V.n7151 ASIG5V.n7150 2.2505
R41891 ASIG5V.n7152 ASIG5V.n6942 2.2505
R41892 ASIG5V.n7154 ASIG5V.n7153 2.2505
R41893 ASIG5V.n6938 ASIG5V.n6937 2.2505
R41894 ASIG5V.n7161 ASIG5V.n7160 2.2505
R41895 ASIG5V.n7162 ASIG5V.n6936 2.2505
R41896 ASIG5V.n7164 ASIG5V.n7163 2.2505
R41897 ASIG5V.n6932 ASIG5V.n6931 2.2505
R41898 ASIG5V.n7171 ASIG5V.n7170 2.2505
R41899 ASIG5V.n7172 ASIG5V.n6930 2.2505
R41900 ASIG5V.n7174 ASIG5V.n7173 2.2505
R41901 ASIG5V.n6926 ASIG5V.n6925 2.2505
R41902 ASIG5V.n7181 ASIG5V.n7180 2.2505
R41903 ASIG5V.n7182 ASIG5V.n6924 2.2505
R41904 ASIG5V.n7184 ASIG5V.n7183 2.2505
R41905 ASIG5V.n6920 ASIG5V.n6919 2.2505
R41906 ASIG5V.n7191 ASIG5V.n7190 2.2505
R41907 ASIG5V.n7192 ASIG5V.n6918 2.2505
R41908 ASIG5V.n7194 ASIG5V.n7193 2.2505
R41909 ASIG5V.n6914 ASIG5V.n6913 2.2505
R41910 ASIG5V.n7201 ASIG5V.n7200 2.2505
R41911 ASIG5V.n7202 ASIG5V.n6912 2.2505
R41912 ASIG5V.n7204 ASIG5V.n7203 2.2505
R41913 ASIG5V.n6908 ASIG5V.n6907 2.2505
R41914 ASIG5V.n7211 ASIG5V.n7210 2.2505
R41915 ASIG5V.n7212 ASIG5V.n6906 2.2505
R41916 ASIG5V.n7214 ASIG5V.n7213 2.2505
R41917 ASIG5V.n6902 ASIG5V.n6901 2.2505
R41918 ASIG5V.n7221 ASIG5V.n7220 2.2505
R41919 ASIG5V.n7222 ASIG5V.n6900 2.2505
R41920 ASIG5V.n7224 ASIG5V.n7223 2.2505
R41921 ASIG5V.n6898 ASIG5V.n6897 2.2505
R41922 ASIG5V.n7231 ASIG5V.n7230 2.2505
R41923 ASIG5V.n7230 ASIG5V.n7229 2.2505
R41924 ASIG5V.n7227 ASIG5V.n6898 2.2505
R41925 ASIG5V.n7225 ASIG5V.n7224 2.2505
R41926 ASIG5V.n6903 ASIG5V.n6900 2.2505
R41927 ASIG5V.n7220 ASIG5V.n7219 2.2505
R41928 ASIG5V.n7217 ASIG5V.n6902 2.2505
R41929 ASIG5V.n7215 ASIG5V.n7214 2.2505
R41930 ASIG5V.n6909 ASIG5V.n6906 2.2505
R41931 ASIG5V.n7210 ASIG5V.n7209 2.2505
R41932 ASIG5V.n7207 ASIG5V.n6908 2.2505
R41933 ASIG5V.n7205 ASIG5V.n7204 2.2505
R41934 ASIG5V.n6915 ASIG5V.n6912 2.2505
R41935 ASIG5V.n7200 ASIG5V.n7199 2.2505
R41936 ASIG5V.n7197 ASIG5V.n6914 2.2505
R41937 ASIG5V.n7195 ASIG5V.n7194 2.2505
R41938 ASIG5V.n6921 ASIG5V.n6918 2.2505
R41939 ASIG5V.n7190 ASIG5V.n7189 2.2505
R41940 ASIG5V.n7187 ASIG5V.n6920 2.2505
R41941 ASIG5V.n7185 ASIG5V.n7184 2.2505
R41942 ASIG5V.n6927 ASIG5V.n6924 2.2505
R41943 ASIG5V.n7180 ASIG5V.n7179 2.2505
R41944 ASIG5V.n7177 ASIG5V.n6926 2.2505
R41945 ASIG5V.n7175 ASIG5V.n7174 2.2505
R41946 ASIG5V.n6933 ASIG5V.n6930 2.2505
R41947 ASIG5V.n7170 ASIG5V.n7169 2.2505
R41948 ASIG5V.n7167 ASIG5V.n6932 2.2505
R41949 ASIG5V.n7165 ASIG5V.n7164 2.2505
R41950 ASIG5V.n6939 ASIG5V.n6936 2.2505
R41951 ASIG5V.n7160 ASIG5V.n7159 2.2505
R41952 ASIG5V.n7157 ASIG5V.n6938 2.2505
R41953 ASIG5V.n7155 ASIG5V.n7154 2.2505
R41954 ASIG5V.n6945 ASIG5V.n6942 2.2505
R41955 ASIG5V.n7150 ASIG5V.n7149 2.2505
R41956 ASIG5V.n7147 ASIG5V.n6944 2.2505
R41957 ASIG5V.n7145 ASIG5V.n7144 2.2505
R41958 ASIG5V.n6951 ASIG5V.n6948 2.2505
R41959 ASIG5V.n7140 ASIG5V.n7139 2.2505
R41960 ASIG5V.n7137 ASIG5V.n6950 2.2505
R41961 ASIG5V.n7135 ASIG5V.n7134 2.2505
R41962 ASIG5V.n6957 ASIG5V.n6954 2.2505
R41963 ASIG5V.n7130 ASIG5V.n7129 2.2505
R41964 ASIG5V.n7127 ASIG5V.n6956 2.2505
R41965 ASIG5V.n7125 ASIG5V.n7124 2.2505
R41966 ASIG5V.n6963 ASIG5V.n6960 2.2505
R41967 ASIG5V.n7120 ASIG5V.n7119 2.2505
R41968 ASIG5V.n7117 ASIG5V.n6962 2.2505
R41969 ASIG5V.n7115 ASIG5V.n7114 2.2505
R41970 ASIG5V.n6969 ASIG5V.n6966 2.2505
R41971 ASIG5V.n7110 ASIG5V.n7109 2.2505
R41972 ASIG5V.n7107 ASIG5V.n6968 2.2505
R41973 ASIG5V.n7105 ASIG5V.n7104 2.2505
R41974 ASIG5V.n6975 ASIG5V.n6972 2.2505
R41975 ASIG5V.n7100 ASIG5V.n7099 2.2505
R41976 ASIG5V.n7097 ASIG5V.n6974 2.2505
R41977 ASIG5V.n7095 ASIG5V.n7094 2.2505
R41978 ASIG5V.n6981 ASIG5V.n6978 2.2505
R41979 ASIG5V.n7090 ASIG5V.n7089 2.2505
R41980 ASIG5V.n7087 ASIG5V.n6980 2.2505
R41981 ASIG5V.n7085 ASIG5V.n7084 2.2505
R41982 ASIG5V.n6987 ASIG5V.n6984 2.2505
R41983 ASIG5V.n7080 ASIG5V.n7079 2.2505
R41984 ASIG5V.n7077 ASIG5V.n6986 2.2505
R41985 ASIG5V.n7075 ASIG5V.n7074 2.2505
R41986 ASIG5V.n6993 ASIG5V.n6990 2.2505
R41987 ASIG5V.n7070 ASIG5V.n7069 2.2505
R41988 ASIG5V.n7067 ASIG5V.n6992 2.2505
R41989 ASIG5V.n7065 ASIG5V.n7064 2.2505
R41990 ASIG5V.n6999 ASIG5V.n6996 2.2505
R41991 ASIG5V.n7060 ASIG5V.n7059 2.2505
R41992 ASIG5V.n7057 ASIG5V.n6998 2.2505
R41993 ASIG5V.n7055 ASIG5V.n7054 2.2505
R41994 ASIG5V.n7005 ASIG5V.n7002 2.2505
R41995 ASIG5V.n7050 ASIG5V.n7049 2.2505
R41996 ASIG5V.n7047 ASIG5V.n7004 2.2505
R41997 ASIG5V.n7045 ASIG5V.n7044 2.2505
R41998 ASIG5V.n7011 ASIG5V.n7008 2.2505
R41999 ASIG5V.n7040 ASIG5V.n7039 2.2505
R42000 ASIG5V.n7037 ASIG5V.n7010 2.2505
R42001 ASIG5V.n7035 ASIG5V.n7034 2.2505
R42002 ASIG5V.n7017 ASIG5V.n7014 2.2505
R42003 ASIG5V.n7030 ASIG5V.n7029 2.2505
R42004 ASIG5V.n7027 ASIG5V.n7016 2.2505
R42005 ASIG5V.n7025 ASIG5V.n7024 2.2505
R42006 ASIG5V.n7021 ASIG5V.n7020 2.2505
R42007 ASIG5V.n8890 ASIG5V.n8263 2.2505
R42008 ASIG5V.n8385 ASIG5V.n8262 2.2505
R42009 ASIG5V.n8388 ASIG5V.n8387 2.2505
R42010 ASIG5V.n8389 ASIG5V.n8384 2.2505
R42011 ASIG5V.n8392 ASIG5V.n8390 2.2505
R42012 ASIG5V.n8394 ASIG5V.n8382 2.2505
R42013 ASIG5V.n8397 ASIG5V.n8396 2.2505
R42014 ASIG5V.n8398 ASIG5V.n8381 2.2505
R42015 ASIG5V.n8401 ASIG5V.n8399 2.2505
R42016 ASIG5V.n8403 ASIG5V.n8379 2.2505
R42017 ASIG5V.n8406 ASIG5V.n8405 2.2505
R42018 ASIG5V.n8407 ASIG5V.n8378 2.2505
R42019 ASIG5V.n8410 ASIG5V.n8408 2.2505
R42020 ASIG5V.n8412 ASIG5V.n8376 2.2505
R42021 ASIG5V.n8415 ASIG5V.n8414 2.2505
R42022 ASIG5V.n8416 ASIG5V.n8375 2.2505
R42023 ASIG5V.n8419 ASIG5V.n8417 2.2505
R42024 ASIG5V.n8421 ASIG5V.n8373 2.2505
R42025 ASIG5V.n8424 ASIG5V.n8423 2.2505
R42026 ASIG5V.n8425 ASIG5V.n8372 2.2505
R42027 ASIG5V.n8428 ASIG5V.n8426 2.2505
R42028 ASIG5V.n8430 ASIG5V.n8370 2.2505
R42029 ASIG5V.n8433 ASIG5V.n8432 2.2505
R42030 ASIG5V.n8434 ASIG5V.n8369 2.2505
R42031 ASIG5V.n8437 ASIG5V.n8435 2.2505
R42032 ASIG5V.n8439 ASIG5V.n8367 2.2505
R42033 ASIG5V.n8442 ASIG5V.n8441 2.2505
R42034 ASIG5V.n8443 ASIG5V.n8366 2.2505
R42035 ASIG5V.n8446 ASIG5V.n8444 2.2505
R42036 ASIG5V.n8448 ASIG5V.n8364 2.2505
R42037 ASIG5V.n8451 ASIG5V.n8450 2.2505
R42038 ASIG5V.n8452 ASIG5V.n8363 2.2505
R42039 ASIG5V.n8455 ASIG5V.n8453 2.2505
R42040 ASIG5V.n8457 ASIG5V.n8361 2.2505
R42041 ASIG5V.n8460 ASIG5V.n8459 2.2505
R42042 ASIG5V.n8461 ASIG5V.n8360 2.2505
R42043 ASIG5V.n8464 ASIG5V.n8462 2.2505
R42044 ASIG5V.n8466 ASIG5V.n8358 2.2505
R42045 ASIG5V.n8469 ASIG5V.n8468 2.2505
R42046 ASIG5V.n8470 ASIG5V.n8357 2.2505
R42047 ASIG5V.n8473 ASIG5V.n8471 2.2505
R42048 ASIG5V.n8475 ASIG5V.n8355 2.2505
R42049 ASIG5V.n8478 ASIG5V.n8477 2.2505
R42050 ASIG5V.n8479 ASIG5V.n8354 2.2505
R42051 ASIG5V.n8482 ASIG5V.n8480 2.2505
R42052 ASIG5V.n8484 ASIG5V.n8352 2.2505
R42053 ASIG5V.n8487 ASIG5V.n8486 2.2505
R42054 ASIG5V.n8488 ASIG5V.n8351 2.2505
R42055 ASIG5V.n8491 ASIG5V.n8489 2.2505
R42056 ASIG5V.n8493 ASIG5V.n8349 2.2505
R42057 ASIG5V.n8496 ASIG5V.n8495 2.2505
R42058 ASIG5V.n8497 ASIG5V.n8348 2.2505
R42059 ASIG5V.n8500 ASIG5V.n8498 2.2505
R42060 ASIG5V.n8502 ASIG5V.n8346 2.2505
R42061 ASIG5V.n8505 ASIG5V.n8504 2.2505
R42062 ASIG5V.n8506 ASIG5V.n8345 2.2505
R42063 ASIG5V.n8509 ASIG5V.n8507 2.2505
R42064 ASIG5V.n8511 ASIG5V.n8343 2.2505
R42065 ASIG5V.n8514 ASIG5V.n8513 2.2505
R42066 ASIG5V.n8515 ASIG5V.n8342 2.2505
R42067 ASIG5V.n8518 ASIG5V.n8516 2.2505
R42068 ASIG5V.n8520 ASIG5V.n8340 2.2505
R42069 ASIG5V.n8523 ASIG5V.n8522 2.2505
R42070 ASIG5V.n8524 ASIG5V.n8339 2.2505
R42071 ASIG5V.n8527 ASIG5V.n8525 2.2505
R42072 ASIG5V.n8529 ASIG5V.n8337 2.2505
R42073 ASIG5V.n8532 ASIG5V.n8531 2.2505
R42074 ASIG5V.n8533 ASIG5V.n8336 2.2505
R42075 ASIG5V.n8536 ASIG5V.n8534 2.2505
R42076 ASIG5V.n8538 ASIG5V.n8334 2.2505
R42077 ASIG5V.n8541 ASIG5V.n8540 2.2505
R42078 ASIG5V.n8542 ASIG5V.n8333 2.2505
R42079 ASIG5V.n8545 ASIG5V.n8543 2.2505
R42080 ASIG5V.n8547 ASIG5V.n8331 2.2505
R42081 ASIG5V.n8550 ASIG5V.n8549 2.2505
R42082 ASIG5V.n8551 ASIG5V.n8330 2.2505
R42083 ASIG5V.n8554 ASIG5V.n8552 2.2505
R42084 ASIG5V.n8556 ASIG5V.n8328 2.2505
R42085 ASIG5V.n8559 ASIG5V.n8558 2.2505
R42086 ASIG5V.n8560 ASIG5V.n8327 2.2505
R42087 ASIG5V.n8563 ASIG5V.n8561 2.2505
R42088 ASIG5V.n8565 ASIG5V.n8325 2.2505
R42089 ASIG5V.n8567 ASIG5V.n8566 2.2505
R42090 ASIG5V.n8568 ASIG5V.n8216 2.2505
R42091 ASIG5V.n8893 ASIG5V.n8216 2.2505
R42092 ASIG5V.n8566 ASIG5V.n8214 2.2505
R42093 ASIG5V.n8565 ASIG5V.n8564 2.2505
R42094 ASIG5V.n8563 ASIG5V.n8562 2.2505
R42095 ASIG5V.n8327 ASIG5V.n8326 2.2505
R42096 ASIG5V.n8558 ASIG5V.n8557 2.2505
R42097 ASIG5V.n8556 ASIG5V.n8555 2.2505
R42098 ASIG5V.n8554 ASIG5V.n8553 2.2505
R42099 ASIG5V.n8330 ASIG5V.n8329 2.2505
R42100 ASIG5V.n8549 ASIG5V.n8548 2.2505
R42101 ASIG5V.n8547 ASIG5V.n8546 2.2505
R42102 ASIG5V.n8545 ASIG5V.n8544 2.2505
R42103 ASIG5V.n8333 ASIG5V.n8332 2.2505
R42104 ASIG5V.n8540 ASIG5V.n8539 2.2505
R42105 ASIG5V.n8538 ASIG5V.n8537 2.2505
R42106 ASIG5V.n8536 ASIG5V.n8535 2.2505
R42107 ASIG5V.n8336 ASIG5V.n8335 2.2505
R42108 ASIG5V.n8531 ASIG5V.n8530 2.2505
R42109 ASIG5V.n8529 ASIG5V.n8528 2.2505
R42110 ASIG5V.n8527 ASIG5V.n8526 2.2505
R42111 ASIG5V.n8339 ASIG5V.n8338 2.2505
R42112 ASIG5V.n8522 ASIG5V.n8521 2.2505
R42113 ASIG5V.n8520 ASIG5V.n8519 2.2505
R42114 ASIG5V.n8518 ASIG5V.n8517 2.2505
R42115 ASIG5V.n8342 ASIG5V.n8341 2.2505
R42116 ASIG5V.n8513 ASIG5V.n8512 2.2505
R42117 ASIG5V.n8511 ASIG5V.n8510 2.2505
R42118 ASIG5V.n8509 ASIG5V.n8508 2.2505
R42119 ASIG5V.n8345 ASIG5V.n8344 2.2505
R42120 ASIG5V.n8504 ASIG5V.n8503 2.2505
R42121 ASIG5V.n8502 ASIG5V.n8501 2.2505
R42122 ASIG5V.n8500 ASIG5V.n8499 2.2505
R42123 ASIG5V.n8348 ASIG5V.n8347 2.2505
R42124 ASIG5V.n8495 ASIG5V.n8494 2.2505
R42125 ASIG5V.n8493 ASIG5V.n8492 2.2505
R42126 ASIG5V.n8491 ASIG5V.n8490 2.2505
R42127 ASIG5V.n8351 ASIG5V.n8350 2.2505
R42128 ASIG5V.n8486 ASIG5V.n8485 2.2505
R42129 ASIG5V.n8484 ASIG5V.n8483 2.2505
R42130 ASIG5V.n8482 ASIG5V.n8481 2.2505
R42131 ASIG5V.n8354 ASIG5V.n8353 2.2505
R42132 ASIG5V.n8477 ASIG5V.n8476 2.2505
R42133 ASIG5V.n8475 ASIG5V.n8474 2.2505
R42134 ASIG5V.n8473 ASIG5V.n8472 2.2505
R42135 ASIG5V.n8357 ASIG5V.n8356 2.2505
R42136 ASIG5V.n8468 ASIG5V.n8467 2.2505
R42137 ASIG5V.n8466 ASIG5V.n8465 2.2505
R42138 ASIG5V.n8464 ASIG5V.n8463 2.2505
R42139 ASIG5V.n8360 ASIG5V.n8359 2.2505
R42140 ASIG5V.n8459 ASIG5V.n8458 2.2505
R42141 ASIG5V.n8457 ASIG5V.n8456 2.2505
R42142 ASIG5V.n8455 ASIG5V.n8454 2.2505
R42143 ASIG5V.n8363 ASIG5V.n8362 2.2505
R42144 ASIG5V.n8450 ASIG5V.n8449 2.2505
R42145 ASIG5V.n8448 ASIG5V.n8447 2.2505
R42146 ASIG5V.n8446 ASIG5V.n8445 2.2505
R42147 ASIG5V.n8366 ASIG5V.n8365 2.2505
R42148 ASIG5V.n8441 ASIG5V.n8440 2.2505
R42149 ASIG5V.n8439 ASIG5V.n8438 2.2505
R42150 ASIG5V.n8437 ASIG5V.n8436 2.2505
R42151 ASIG5V.n8369 ASIG5V.n8368 2.2505
R42152 ASIG5V.n8432 ASIG5V.n8431 2.2505
R42153 ASIG5V.n8430 ASIG5V.n8429 2.2505
R42154 ASIG5V.n8428 ASIG5V.n8427 2.2505
R42155 ASIG5V.n8372 ASIG5V.n8371 2.2505
R42156 ASIG5V.n8423 ASIG5V.n8422 2.2505
R42157 ASIG5V.n8421 ASIG5V.n8420 2.2505
R42158 ASIG5V.n8419 ASIG5V.n8418 2.2505
R42159 ASIG5V.n8375 ASIG5V.n8374 2.2505
R42160 ASIG5V.n8414 ASIG5V.n8413 2.2505
R42161 ASIG5V.n8412 ASIG5V.n8411 2.2505
R42162 ASIG5V.n8410 ASIG5V.n8409 2.2505
R42163 ASIG5V.n8378 ASIG5V.n8377 2.2505
R42164 ASIG5V.n8405 ASIG5V.n8404 2.2505
R42165 ASIG5V.n8403 ASIG5V.n8402 2.2505
R42166 ASIG5V.n8401 ASIG5V.n8400 2.2505
R42167 ASIG5V.n8381 ASIG5V.n8380 2.2505
R42168 ASIG5V.n8396 ASIG5V.n8395 2.2505
R42169 ASIG5V.n8394 ASIG5V.n8393 2.2505
R42170 ASIG5V.n8392 ASIG5V.n8391 2.2505
R42171 ASIG5V.n8384 ASIG5V.n8383 2.2505
R42172 ASIG5V.n8387 ASIG5V.n8386 2.2505
R42173 ASIG5V.n8262 ASIG5V.n8261 2.2505
R42174 ASIG5V.n8891 ASIG5V.n8890 2.2505
R42175 ASIG5V.n8634 ASIG5V.n8633 2.2505
R42176 ASIG5V.n8635 ASIG5V.n8631 2.2505
R42177 ASIG5V.n8640 ASIG5V.n8636 2.2505
R42178 ASIG5V.n8641 ASIG5V.n8630 2.2505
R42179 ASIG5V.n8646 ASIG5V.n8645 2.2505
R42180 ASIG5V.n8647 ASIG5V.n8629 2.2505
R42181 ASIG5V.n8652 ASIG5V.n8648 2.2505
R42182 ASIG5V.n8653 ASIG5V.n8628 2.2505
R42183 ASIG5V.n8658 ASIG5V.n8657 2.2505
R42184 ASIG5V.n8659 ASIG5V.n8627 2.2505
R42185 ASIG5V.n8664 ASIG5V.n8660 2.2505
R42186 ASIG5V.n8665 ASIG5V.n8626 2.2505
R42187 ASIG5V.n8670 ASIG5V.n8669 2.2505
R42188 ASIG5V.n8671 ASIG5V.n8625 2.2505
R42189 ASIG5V.n8676 ASIG5V.n8672 2.2505
R42190 ASIG5V.n8677 ASIG5V.n8624 2.2505
R42191 ASIG5V.n8682 ASIG5V.n8681 2.2505
R42192 ASIG5V.n8683 ASIG5V.n8623 2.2505
R42193 ASIG5V.n8688 ASIG5V.n8684 2.2505
R42194 ASIG5V.n8689 ASIG5V.n8622 2.2505
R42195 ASIG5V.n8694 ASIG5V.n8693 2.2505
R42196 ASIG5V.n8695 ASIG5V.n8621 2.2505
R42197 ASIG5V.n8700 ASIG5V.n8696 2.2505
R42198 ASIG5V.n8701 ASIG5V.n8620 2.2505
R42199 ASIG5V.n8706 ASIG5V.n8705 2.2505
R42200 ASIG5V.n8707 ASIG5V.n8619 2.2505
R42201 ASIG5V.n8712 ASIG5V.n8708 2.2505
R42202 ASIG5V.n8713 ASIG5V.n8618 2.2505
R42203 ASIG5V.n8718 ASIG5V.n8717 2.2505
R42204 ASIG5V.n8719 ASIG5V.n8617 2.2505
R42205 ASIG5V.n8724 ASIG5V.n8720 2.2505
R42206 ASIG5V.n8725 ASIG5V.n8616 2.2505
R42207 ASIG5V.n8730 ASIG5V.n8729 2.2505
R42208 ASIG5V.n8731 ASIG5V.n8615 2.2505
R42209 ASIG5V.n8736 ASIG5V.n8732 2.2505
R42210 ASIG5V.n8737 ASIG5V.n8614 2.2505
R42211 ASIG5V.n8742 ASIG5V.n8741 2.2505
R42212 ASIG5V.n8743 ASIG5V.n8613 2.2505
R42213 ASIG5V.n8748 ASIG5V.n8744 2.2505
R42214 ASIG5V.n8749 ASIG5V.n8612 2.2505
R42215 ASIG5V.n8754 ASIG5V.n8753 2.2505
R42216 ASIG5V.n8755 ASIG5V.n8611 2.2505
R42217 ASIG5V.n8760 ASIG5V.n8756 2.2505
R42218 ASIG5V.n8761 ASIG5V.n8610 2.2505
R42219 ASIG5V.n8766 ASIG5V.n8765 2.2505
R42220 ASIG5V.n8767 ASIG5V.n8609 2.2505
R42221 ASIG5V.n8772 ASIG5V.n8768 2.2505
R42222 ASIG5V.n8773 ASIG5V.n8608 2.2505
R42223 ASIG5V.n8778 ASIG5V.n8777 2.2505
R42224 ASIG5V.n8779 ASIG5V.n8607 2.2505
R42225 ASIG5V.n8784 ASIG5V.n8780 2.2505
R42226 ASIG5V.n8785 ASIG5V.n8606 2.2505
R42227 ASIG5V.n8790 ASIG5V.n8789 2.2505
R42228 ASIG5V.n8791 ASIG5V.n8605 2.2505
R42229 ASIG5V.n8796 ASIG5V.n8792 2.2505
R42230 ASIG5V.n8797 ASIG5V.n8604 2.2505
R42231 ASIG5V.n8802 ASIG5V.n8801 2.2505
R42232 ASIG5V.n8803 ASIG5V.n8603 2.2505
R42233 ASIG5V.n8808 ASIG5V.n8804 2.2505
R42234 ASIG5V.n8809 ASIG5V.n8602 2.2505
R42235 ASIG5V.n8814 ASIG5V.n8813 2.2505
R42236 ASIG5V.n8815 ASIG5V.n8601 2.2505
R42237 ASIG5V.n8820 ASIG5V.n8816 2.2505
R42238 ASIG5V.n8821 ASIG5V.n8600 2.2505
R42239 ASIG5V.n8826 ASIG5V.n8825 2.2505
R42240 ASIG5V.n8827 ASIG5V.n8599 2.2505
R42241 ASIG5V.n8832 ASIG5V.n8828 2.2505
R42242 ASIG5V.n8833 ASIG5V.n8598 2.2505
R42243 ASIG5V.n8838 ASIG5V.n8837 2.2505
R42244 ASIG5V.n8839 ASIG5V.n8597 2.2505
R42245 ASIG5V.n8844 ASIG5V.n8840 2.2505
R42246 ASIG5V.n8845 ASIG5V.n8596 2.2505
R42247 ASIG5V.n8850 ASIG5V.n8849 2.2505
R42248 ASIG5V.n8851 ASIG5V.n8595 2.2505
R42249 ASIG5V.n8856 ASIG5V.n8852 2.2505
R42250 ASIG5V.n8857 ASIG5V.n8594 2.2505
R42251 ASIG5V.n8862 ASIG5V.n8861 2.2505
R42252 ASIG5V.n8863 ASIG5V.n8593 2.2505
R42253 ASIG5V.n8868 ASIG5V.n8864 2.2505
R42254 ASIG5V.n8869 ASIG5V.n8592 2.2505
R42255 ASIG5V.n8874 ASIG5V.n8873 2.2505
R42256 ASIG5V.n8875 ASIG5V.n8591 2.2505
R42257 ASIG5V.n8877 ASIG5V.n8876 2.2505
R42258 ASIG5V.n8878 ASIG5V.n8588 2.2505
R42259 ASIG5V.n8879 ASIG5V.n8878 2.2505
R42260 ASIG5V.n8877 ASIG5V.n8319 2.2505
R42261 ASIG5V.n8591 ASIG5V.n8590 2.2505
R42262 ASIG5V.n8873 ASIG5V.n8872 2.2505
R42263 ASIG5V.n8870 ASIG5V.n8869 2.2505
R42264 ASIG5V.n8868 ASIG5V.n8867 2.2505
R42265 ASIG5V.n8865 ASIG5V.n8593 2.2505
R42266 ASIG5V.n8861 ASIG5V.n8860 2.2505
R42267 ASIG5V.n8858 ASIG5V.n8857 2.2505
R42268 ASIG5V.n8856 ASIG5V.n8855 2.2505
R42269 ASIG5V.n8853 ASIG5V.n8595 2.2505
R42270 ASIG5V.n8849 ASIG5V.n8848 2.2505
R42271 ASIG5V.n8846 ASIG5V.n8845 2.2505
R42272 ASIG5V.n8844 ASIG5V.n8843 2.2505
R42273 ASIG5V.n8841 ASIG5V.n8597 2.2505
R42274 ASIG5V.n8837 ASIG5V.n8836 2.2505
R42275 ASIG5V.n8834 ASIG5V.n8833 2.2505
R42276 ASIG5V.n8832 ASIG5V.n8831 2.2505
R42277 ASIG5V.n8829 ASIG5V.n8599 2.2505
R42278 ASIG5V.n8825 ASIG5V.n8824 2.2505
R42279 ASIG5V.n8822 ASIG5V.n8821 2.2505
R42280 ASIG5V.n8820 ASIG5V.n8819 2.2505
R42281 ASIG5V.n8817 ASIG5V.n8601 2.2505
R42282 ASIG5V.n8813 ASIG5V.n8812 2.2505
R42283 ASIG5V.n8810 ASIG5V.n8809 2.2505
R42284 ASIG5V.n8808 ASIG5V.n8807 2.2505
R42285 ASIG5V.n8805 ASIG5V.n8603 2.2505
R42286 ASIG5V.n8801 ASIG5V.n8800 2.2505
R42287 ASIG5V.n8798 ASIG5V.n8797 2.2505
R42288 ASIG5V.n8796 ASIG5V.n8795 2.2505
R42289 ASIG5V.n8793 ASIG5V.n8605 2.2505
R42290 ASIG5V.n8789 ASIG5V.n8788 2.2505
R42291 ASIG5V.n8786 ASIG5V.n8785 2.2505
R42292 ASIG5V.n8784 ASIG5V.n8783 2.2505
R42293 ASIG5V.n8781 ASIG5V.n8607 2.2505
R42294 ASIG5V.n8777 ASIG5V.n8776 2.2505
R42295 ASIG5V.n8774 ASIG5V.n8773 2.2505
R42296 ASIG5V.n8772 ASIG5V.n8771 2.2505
R42297 ASIG5V.n8769 ASIG5V.n8609 2.2505
R42298 ASIG5V.n8765 ASIG5V.n8764 2.2505
R42299 ASIG5V.n8762 ASIG5V.n8761 2.2505
R42300 ASIG5V.n8760 ASIG5V.n8759 2.2505
R42301 ASIG5V.n8757 ASIG5V.n8611 2.2505
R42302 ASIG5V.n8753 ASIG5V.n8752 2.2505
R42303 ASIG5V.n8750 ASIG5V.n8749 2.2505
R42304 ASIG5V.n8748 ASIG5V.n8747 2.2505
R42305 ASIG5V.n8745 ASIG5V.n8613 2.2505
R42306 ASIG5V.n8741 ASIG5V.n8740 2.2505
R42307 ASIG5V.n8738 ASIG5V.n8737 2.2505
R42308 ASIG5V.n8736 ASIG5V.n8735 2.2505
R42309 ASIG5V.n8733 ASIG5V.n8615 2.2505
R42310 ASIG5V.n8729 ASIG5V.n8728 2.2505
R42311 ASIG5V.n8726 ASIG5V.n8725 2.2505
R42312 ASIG5V.n8724 ASIG5V.n8723 2.2505
R42313 ASIG5V.n8721 ASIG5V.n8617 2.2505
R42314 ASIG5V.n8717 ASIG5V.n8716 2.2505
R42315 ASIG5V.n8714 ASIG5V.n8713 2.2505
R42316 ASIG5V.n8712 ASIG5V.n8711 2.2505
R42317 ASIG5V.n8709 ASIG5V.n8619 2.2505
R42318 ASIG5V.n8705 ASIG5V.n8704 2.2505
R42319 ASIG5V.n8702 ASIG5V.n8701 2.2505
R42320 ASIG5V.n8700 ASIG5V.n8699 2.2505
R42321 ASIG5V.n8697 ASIG5V.n8621 2.2505
R42322 ASIG5V.n8693 ASIG5V.n8692 2.2505
R42323 ASIG5V.n8690 ASIG5V.n8689 2.2505
R42324 ASIG5V.n8688 ASIG5V.n8687 2.2505
R42325 ASIG5V.n8685 ASIG5V.n8623 2.2505
R42326 ASIG5V.n8681 ASIG5V.n8680 2.2505
R42327 ASIG5V.n8678 ASIG5V.n8677 2.2505
R42328 ASIG5V.n8676 ASIG5V.n8675 2.2505
R42329 ASIG5V.n8673 ASIG5V.n8625 2.2505
R42330 ASIG5V.n8669 ASIG5V.n8668 2.2505
R42331 ASIG5V.n8666 ASIG5V.n8665 2.2505
R42332 ASIG5V.n8664 ASIG5V.n8663 2.2505
R42333 ASIG5V.n8661 ASIG5V.n8627 2.2505
R42334 ASIG5V.n8657 ASIG5V.n8656 2.2505
R42335 ASIG5V.n8654 ASIG5V.n8653 2.2505
R42336 ASIG5V.n8652 ASIG5V.n8651 2.2505
R42337 ASIG5V.n8649 ASIG5V.n8629 2.2505
R42338 ASIG5V.n8645 ASIG5V.n8644 2.2505
R42339 ASIG5V.n8642 ASIG5V.n8641 2.2505
R42340 ASIG5V.n8640 ASIG5V.n8639 2.2505
R42341 ASIG5V.n8637 ASIG5V.n8631 2.2505
R42342 ASIG5V.n8633 ASIG5V.n8632 2.2505
R42343 ASIG5V.n12523 ASIG5V.n12522 2.2505
R42344 ASIG5V.n12521 ASIG5V.n100 2.2505
R42345 ASIG5V.n12520 ASIG5V.n12519 2.2505
R42346 ASIG5V.n12517 ASIG5V.n101 2.2505
R42347 ASIG5V.n12515 ASIG5V.n12513 2.2505
R42348 ASIG5V.n12512 ASIG5V.n103 2.2505
R42349 ASIG5V.n12511 ASIG5V.n12510 2.2505
R42350 ASIG5V.n12508 ASIG5V.n104 2.2505
R42351 ASIG5V.n12506 ASIG5V.n12504 2.2505
R42352 ASIG5V.n12503 ASIG5V.n106 2.2505
R42353 ASIG5V.n12502 ASIG5V.n12501 2.2505
R42354 ASIG5V.n12499 ASIG5V.n107 2.2505
R42355 ASIG5V.n12497 ASIG5V.n12495 2.2505
R42356 ASIG5V.n12494 ASIG5V.n109 2.2505
R42357 ASIG5V.n12493 ASIG5V.n12492 2.2505
R42358 ASIG5V.n12490 ASIG5V.n110 2.2505
R42359 ASIG5V.n12488 ASIG5V.n12486 2.2505
R42360 ASIG5V.n12485 ASIG5V.n112 2.2505
R42361 ASIG5V.n12484 ASIG5V.n12483 2.2505
R42362 ASIG5V.n12481 ASIG5V.n113 2.2505
R42363 ASIG5V.n12479 ASIG5V.n12477 2.2505
R42364 ASIG5V.n12476 ASIG5V.n115 2.2505
R42365 ASIG5V.n12475 ASIG5V.n12474 2.2505
R42366 ASIG5V.n12472 ASIG5V.n116 2.2505
R42367 ASIG5V.n12470 ASIG5V.n12468 2.2505
R42368 ASIG5V.n12467 ASIG5V.n118 2.2505
R42369 ASIG5V.n12466 ASIG5V.n12465 2.2505
R42370 ASIG5V.n12463 ASIG5V.n119 2.2505
R42371 ASIG5V.n12461 ASIG5V.n12459 2.2505
R42372 ASIG5V.n12458 ASIG5V.n121 2.2505
R42373 ASIG5V.n12457 ASIG5V.n12456 2.2505
R42374 ASIG5V.n12454 ASIG5V.n122 2.2505
R42375 ASIG5V.n12452 ASIG5V.n12450 2.2505
R42376 ASIG5V.n12449 ASIG5V.n124 2.2505
R42377 ASIG5V.n12448 ASIG5V.n12447 2.2505
R42378 ASIG5V.n12445 ASIG5V.n125 2.2505
R42379 ASIG5V.n12443 ASIG5V.n12441 2.2505
R42380 ASIG5V.n12440 ASIG5V.n127 2.2505
R42381 ASIG5V.n12439 ASIG5V.n12438 2.2505
R42382 ASIG5V.n12436 ASIG5V.n128 2.2505
R42383 ASIG5V.n12434 ASIG5V.n12432 2.2505
R42384 ASIG5V.n12431 ASIG5V.n130 2.2505
R42385 ASIG5V.n12430 ASIG5V.n12429 2.2505
R42386 ASIG5V.n12427 ASIG5V.n131 2.2505
R42387 ASIG5V.n12425 ASIG5V.n12423 2.2505
R42388 ASIG5V.n12422 ASIG5V.n133 2.2505
R42389 ASIG5V.n12421 ASIG5V.n12420 2.2505
R42390 ASIG5V.n12418 ASIG5V.n134 2.2505
R42391 ASIG5V.n12416 ASIG5V.n12414 2.2505
R42392 ASIG5V.n12413 ASIG5V.n136 2.2505
R42393 ASIG5V.n12412 ASIG5V.n12411 2.2505
R42394 ASIG5V.n12409 ASIG5V.n137 2.2505
R42395 ASIG5V.n12407 ASIG5V.n12405 2.2505
R42396 ASIG5V.n12404 ASIG5V.n139 2.2505
R42397 ASIG5V.n12403 ASIG5V.n12402 2.2505
R42398 ASIG5V.n12400 ASIG5V.n140 2.2505
R42399 ASIG5V.n12398 ASIG5V.n12396 2.2505
R42400 ASIG5V.n12395 ASIG5V.n142 2.2505
R42401 ASIG5V.n12394 ASIG5V.n12393 2.2505
R42402 ASIG5V.n12391 ASIG5V.n143 2.2505
R42403 ASIG5V.n12389 ASIG5V.n12387 2.2505
R42404 ASIG5V.n12386 ASIG5V.n145 2.2505
R42405 ASIG5V.n12385 ASIG5V.n12384 2.2505
R42406 ASIG5V.n12382 ASIG5V.n146 2.2505
R42407 ASIG5V.n12380 ASIG5V.n12378 2.2505
R42408 ASIG5V.n12377 ASIG5V.n148 2.2505
R42409 ASIG5V.n12376 ASIG5V.n12375 2.2505
R42410 ASIG5V.n12373 ASIG5V.n149 2.2505
R42411 ASIG5V.n12371 ASIG5V.n12369 2.2505
R42412 ASIG5V.n12368 ASIG5V.n151 2.2505
R42413 ASIG5V.n12367 ASIG5V.n12366 2.2505
R42414 ASIG5V.n12364 ASIG5V.n152 2.2505
R42415 ASIG5V.n12362 ASIG5V.n12360 2.2505
R42416 ASIG5V.n12359 ASIG5V.n154 2.2505
R42417 ASIG5V.n12358 ASIG5V.n12357 2.2505
R42418 ASIG5V.n12355 ASIG5V.n155 2.2505
R42419 ASIG5V.n12353 ASIG5V.n12351 2.2505
R42420 ASIG5V.n12350 ASIG5V.n157 2.2505
R42421 ASIG5V.n12349 ASIG5V.n12348 2.2505
R42422 ASIG5V.n12346 ASIG5V.n158 2.2505
R42423 ASIG5V.n12344 ASIG5V.n12342 2.2505
R42424 ASIG5V.n12341 ASIG5V.n160 2.2505
R42425 ASIG5V.n12340 ASIG5V.n12339 2.2505
R42426 ASIG5V.n12338 ASIG5V.n55 2.2505
R42427 ASIG5V.n12526 ASIG5V.n55 2.2505
R42428 ASIG5V.n12339 ASIG5V.n53 2.2505
R42429 ASIG5V.n160 ASIG5V.n159 2.2505
R42430 ASIG5V.n12344 ASIG5V.n12343 2.2505
R42431 ASIG5V.n12346 ASIG5V.n12345 2.2505
R42432 ASIG5V.n12348 ASIG5V.n12347 2.2505
R42433 ASIG5V.n157 ASIG5V.n156 2.2505
R42434 ASIG5V.n12353 ASIG5V.n12352 2.2505
R42435 ASIG5V.n12355 ASIG5V.n12354 2.2505
R42436 ASIG5V.n12357 ASIG5V.n12356 2.2505
R42437 ASIG5V.n154 ASIG5V.n153 2.2505
R42438 ASIG5V.n12362 ASIG5V.n12361 2.2505
R42439 ASIG5V.n12364 ASIG5V.n12363 2.2505
R42440 ASIG5V.n12366 ASIG5V.n12365 2.2505
R42441 ASIG5V.n151 ASIG5V.n150 2.2505
R42442 ASIG5V.n12371 ASIG5V.n12370 2.2505
R42443 ASIG5V.n12373 ASIG5V.n12372 2.2505
R42444 ASIG5V.n12375 ASIG5V.n12374 2.2505
R42445 ASIG5V.n148 ASIG5V.n147 2.2505
R42446 ASIG5V.n12380 ASIG5V.n12379 2.2505
R42447 ASIG5V.n12382 ASIG5V.n12381 2.2505
R42448 ASIG5V.n12384 ASIG5V.n12383 2.2505
R42449 ASIG5V.n145 ASIG5V.n144 2.2505
R42450 ASIG5V.n12389 ASIG5V.n12388 2.2505
R42451 ASIG5V.n12391 ASIG5V.n12390 2.2505
R42452 ASIG5V.n12393 ASIG5V.n12392 2.2505
R42453 ASIG5V.n142 ASIG5V.n141 2.2505
R42454 ASIG5V.n12398 ASIG5V.n12397 2.2505
R42455 ASIG5V.n12400 ASIG5V.n12399 2.2505
R42456 ASIG5V.n12402 ASIG5V.n12401 2.2505
R42457 ASIG5V.n139 ASIG5V.n138 2.2505
R42458 ASIG5V.n12407 ASIG5V.n12406 2.2505
R42459 ASIG5V.n12409 ASIG5V.n12408 2.2505
R42460 ASIG5V.n12411 ASIG5V.n12410 2.2505
R42461 ASIG5V.n136 ASIG5V.n135 2.2505
R42462 ASIG5V.n12416 ASIG5V.n12415 2.2505
R42463 ASIG5V.n12418 ASIG5V.n12417 2.2505
R42464 ASIG5V.n12420 ASIG5V.n12419 2.2505
R42465 ASIG5V.n133 ASIG5V.n132 2.2505
R42466 ASIG5V.n12425 ASIG5V.n12424 2.2505
R42467 ASIG5V.n12427 ASIG5V.n12426 2.2505
R42468 ASIG5V.n12429 ASIG5V.n12428 2.2505
R42469 ASIG5V.n130 ASIG5V.n129 2.2505
R42470 ASIG5V.n12434 ASIG5V.n12433 2.2505
R42471 ASIG5V.n12436 ASIG5V.n12435 2.2505
R42472 ASIG5V.n12438 ASIG5V.n12437 2.2505
R42473 ASIG5V.n127 ASIG5V.n126 2.2505
R42474 ASIG5V.n12443 ASIG5V.n12442 2.2505
R42475 ASIG5V.n12445 ASIG5V.n12444 2.2505
R42476 ASIG5V.n12447 ASIG5V.n12446 2.2505
R42477 ASIG5V.n124 ASIG5V.n123 2.2505
R42478 ASIG5V.n12452 ASIG5V.n12451 2.2505
R42479 ASIG5V.n12454 ASIG5V.n12453 2.2505
R42480 ASIG5V.n12456 ASIG5V.n12455 2.2505
R42481 ASIG5V.n121 ASIG5V.n120 2.2505
R42482 ASIG5V.n12461 ASIG5V.n12460 2.2505
R42483 ASIG5V.n12463 ASIG5V.n12462 2.2505
R42484 ASIG5V.n12465 ASIG5V.n12464 2.2505
R42485 ASIG5V.n118 ASIG5V.n117 2.2505
R42486 ASIG5V.n12470 ASIG5V.n12469 2.2505
R42487 ASIG5V.n12472 ASIG5V.n12471 2.2505
R42488 ASIG5V.n12474 ASIG5V.n12473 2.2505
R42489 ASIG5V.n115 ASIG5V.n114 2.2505
R42490 ASIG5V.n12479 ASIG5V.n12478 2.2505
R42491 ASIG5V.n12481 ASIG5V.n12480 2.2505
R42492 ASIG5V.n12483 ASIG5V.n12482 2.2505
R42493 ASIG5V.n112 ASIG5V.n111 2.2505
R42494 ASIG5V.n12488 ASIG5V.n12487 2.2505
R42495 ASIG5V.n12490 ASIG5V.n12489 2.2505
R42496 ASIG5V.n12492 ASIG5V.n12491 2.2505
R42497 ASIG5V.n109 ASIG5V.n108 2.2505
R42498 ASIG5V.n12497 ASIG5V.n12496 2.2505
R42499 ASIG5V.n12499 ASIG5V.n12498 2.2505
R42500 ASIG5V.n12501 ASIG5V.n12500 2.2505
R42501 ASIG5V.n106 ASIG5V.n105 2.2505
R42502 ASIG5V.n12506 ASIG5V.n12505 2.2505
R42503 ASIG5V.n12508 ASIG5V.n12507 2.2505
R42504 ASIG5V.n12510 ASIG5V.n12509 2.2505
R42505 ASIG5V.n103 ASIG5V.n102 2.2505
R42506 ASIG5V.n12515 ASIG5V.n12514 2.2505
R42507 ASIG5V.n12517 ASIG5V.n12516 2.2505
R42508 ASIG5V.n12519 ASIG5V.n12518 2.2505
R42509 ASIG5V.n100 ASIG5V.n99 2.2505
R42510 ASIG5V.n12524 ASIG5V.n12523 2.2505
R42511 ASIG5V.n12317 ASIG5V.n218 2.2505
R42512 ASIG5V.n12319 ASIG5V.n12318 2.2505
R42513 ASIG5V.n504 ASIG5V.n220 2.2505
R42514 ASIG5V.n503 ASIG5V.n502 2.2505
R42515 ASIG5V.n498 ASIG5V.n221 2.2505
R42516 ASIG5V.n494 ASIG5V.n493 2.2505
R42517 ASIG5V.n492 ASIG5V.n222 2.2505
R42518 ASIG5V.n491 ASIG5V.n490 2.2505
R42519 ASIG5V.n486 ASIG5V.n223 2.2505
R42520 ASIG5V.n482 ASIG5V.n481 2.2505
R42521 ASIG5V.n480 ASIG5V.n224 2.2505
R42522 ASIG5V.n479 ASIG5V.n478 2.2505
R42523 ASIG5V.n474 ASIG5V.n225 2.2505
R42524 ASIG5V.n470 ASIG5V.n469 2.2505
R42525 ASIG5V.n468 ASIG5V.n226 2.2505
R42526 ASIG5V.n467 ASIG5V.n466 2.2505
R42527 ASIG5V.n462 ASIG5V.n227 2.2505
R42528 ASIG5V.n458 ASIG5V.n457 2.2505
R42529 ASIG5V.n456 ASIG5V.n228 2.2505
R42530 ASIG5V.n455 ASIG5V.n454 2.2505
R42531 ASIG5V.n450 ASIG5V.n229 2.2505
R42532 ASIG5V.n446 ASIG5V.n445 2.2505
R42533 ASIG5V.n444 ASIG5V.n230 2.2505
R42534 ASIG5V.n443 ASIG5V.n442 2.2505
R42535 ASIG5V.n438 ASIG5V.n231 2.2505
R42536 ASIG5V.n434 ASIG5V.n433 2.2505
R42537 ASIG5V.n432 ASIG5V.n232 2.2505
R42538 ASIG5V.n431 ASIG5V.n430 2.2505
R42539 ASIG5V.n426 ASIG5V.n233 2.2505
R42540 ASIG5V.n422 ASIG5V.n421 2.2505
R42541 ASIG5V.n420 ASIG5V.n234 2.2505
R42542 ASIG5V.n419 ASIG5V.n418 2.2505
R42543 ASIG5V.n414 ASIG5V.n235 2.2505
R42544 ASIG5V.n410 ASIG5V.n409 2.2505
R42545 ASIG5V.n408 ASIG5V.n236 2.2505
R42546 ASIG5V.n407 ASIG5V.n406 2.2505
R42547 ASIG5V.n402 ASIG5V.n237 2.2505
R42548 ASIG5V.n398 ASIG5V.n397 2.2505
R42549 ASIG5V.n396 ASIG5V.n238 2.2505
R42550 ASIG5V.n395 ASIG5V.n394 2.2505
R42551 ASIG5V.n390 ASIG5V.n239 2.2505
R42552 ASIG5V.n386 ASIG5V.n385 2.2505
R42553 ASIG5V.n384 ASIG5V.n240 2.2505
R42554 ASIG5V.n383 ASIG5V.n382 2.2505
R42555 ASIG5V.n378 ASIG5V.n241 2.2505
R42556 ASIG5V.n374 ASIG5V.n373 2.2505
R42557 ASIG5V.n372 ASIG5V.n242 2.2505
R42558 ASIG5V.n371 ASIG5V.n370 2.2505
R42559 ASIG5V.n366 ASIG5V.n243 2.2505
R42560 ASIG5V.n362 ASIG5V.n361 2.2505
R42561 ASIG5V.n360 ASIG5V.n244 2.2505
R42562 ASIG5V.n359 ASIG5V.n358 2.2505
R42563 ASIG5V.n354 ASIG5V.n245 2.2505
R42564 ASIG5V.n350 ASIG5V.n349 2.2505
R42565 ASIG5V.n348 ASIG5V.n246 2.2505
R42566 ASIG5V.n347 ASIG5V.n346 2.2505
R42567 ASIG5V.n342 ASIG5V.n247 2.2505
R42568 ASIG5V.n338 ASIG5V.n337 2.2505
R42569 ASIG5V.n336 ASIG5V.n248 2.2505
R42570 ASIG5V.n335 ASIG5V.n334 2.2505
R42571 ASIG5V.n330 ASIG5V.n249 2.2505
R42572 ASIG5V.n326 ASIG5V.n325 2.2505
R42573 ASIG5V.n324 ASIG5V.n250 2.2505
R42574 ASIG5V.n323 ASIG5V.n322 2.2505
R42575 ASIG5V.n318 ASIG5V.n251 2.2505
R42576 ASIG5V.n314 ASIG5V.n313 2.2505
R42577 ASIG5V.n312 ASIG5V.n252 2.2505
R42578 ASIG5V.n311 ASIG5V.n310 2.2505
R42579 ASIG5V.n306 ASIG5V.n253 2.2505
R42580 ASIG5V.n302 ASIG5V.n301 2.2505
R42581 ASIG5V.n300 ASIG5V.n254 2.2505
R42582 ASIG5V.n299 ASIG5V.n298 2.2505
R42583 ASIG5V.n294 ASIG5V.n255 2.2505
R42584 ASIG5V.n290 ASIG5V.n289 2.2505
R42585 ASIG5V.n288 ASIG5V.n256 2.2505
R42586 ASIG5V.n287 ASIG5V.n286 2.2505
R42587 ASIG5V.n282 ASIG5V.n257 2.2505
R42588 ASIG5V.n278 ASIG5V.n277 2.2505
R42589 ASIG5V.n276 ASIG5V.n258 2.2505
R42590 ASIG5V.n275 ASIG5V.n274 2.2505
R42591 ASIG5V.n270 ASIG5V.n259 2.2505
R42592 ASIG5V.n266 ASIG5V.n265 2.2505
R42593 ASIG5V.n264 ASIG5V.n263 2.2505
R42594 ASIG5V.n260 ASIG5V.n168 2.2505
R42595 ASIG5V.n260 ASIG5V.n215 2.2505
R42596 ASIG5V.n263 ASIG5V.n262 2.2505
R42597 ASIG5V.n267 ASIG5V.n266 2.2505
R42598 ASIG5V.n270 ASIG5V.n269 2.2505
R42599 ASIG5V.n274 ASIG5V.n273 2.2505
R42600 ASIG5V.n271 ASIG5V.n258 2.2505
R42601 ASIG5V.n279 ASIG5V.n278 2.2505
R42602 ASIG5V.n282 ASIG5V.n281 2.2505
R42603 ASIG5V.n286 ASIG5V.n285 2.2505
R42604 ASIG5V.n283 ASIG5V.n256 2.2505
R42605 ASIG5V.n291 ASIG5V.n290 2.2505
R42606 ASIG5V.n294 ASIG5V.n293 2.2505
R42607 ASIG5V.n298 ASIG5V.n297 2.2505
R42608 ASIG5V.n295 ASIG5V.n254 2.2505
R42609 ASIG5V.n303 ASIG5V.n302 2.2505
R42610 ASIG5V.n306 ASIG5V.n305 2.2505
R42611 ASIG5V.n310 ASIG5V.n309 2.2505
R42612 ASIG5V.n307 ASIG5V.n252 2.2505
R42613 ASIG5V.n315 ASIG5V.n314 2.2505
R42614 ASIG5V.n318 ASIG5V.n317 2.2505
R42615 ASIG5V.n322 ASIG5V.n321 2.2505
R42616 ASIG5V.n319 ASIG5V.n250 2.2505
R42617 ASIG5V.n327 ASIG5V.n326 2.2505
R42618 ASIG5V.n330 ASIG5V.n329 2.2505
R42619 ASIG5V.n334 ASIG5V.n333 2.2505
R42620 ASIG5V.n331 ASIG5V.n248 2.2505
R42621 ASIG5V.n339 ASIG5V.n338 2.2505
R42622 ASIG5V.n342 ASIG5V.n341 2.2505
R42623 ASIG5V.n346 ASIG5V.n345 2.2505
R42624 ASIG5V.n343 ASIG5V.n246 2.2505
R42625 ASIG5V.n351 ASIG5V.n350 2.2505
R42626 ASIG5V.n354 ASIG5V.n353 2.2505
R42627 ASIG5V.n358 ASIG5V.n357 2.2505
R42628 ASIG5V.n355 ASIG5V.n244 2.2505
R42629 ASIG5V.n363 ASIG5V.n362 2.2505
R42630 ASIG5V.n366 ASIG5V.n365 2.2505
R42631 ASIG5V.n370 ASIG5V.n369 2.2505
R42632 ASIG5V.n367 ASIG5V.n242 2.2505
R42633 ASIG5V.n375 ASIG5V.n374 2.2505
R42634 ASIG5V.n378 ASIG5V.n377 2.2505
R42635 ASIG5V.n382 ASIG5V.n381 2.2505
R42636 ASIG5V.n379 ASIG5V.n240 2.2505
R42637 ASIG5V.n387 ASIG5V.n386 2.2505
R42638 ASIG5V.n390 ASIG5V.n389 2.2505
R42639 ASIG5V.n394 ASIG5V.n393 2.2505
R42640 ASIG5V.n391 ASIG5V.n238 2.2505
R42641 ASIG5V.n399 ASIG5V.n398 2.2505
R42642 ASIG5V.n402 ASIG5V.n401 2.2505
R42643 ASIG5V.n406 ASIG5V.n405 2.2505
R42644 ASIG5V.n403 ASIG5V.n236 2.2505
R42645 ASIG5V.n411 ASIG5V.n410 2.2505
R42646 ASIG5V.n414 ASIG5V.n413 2.2505
R42647 ASIG5V.n418 ASIG5V.n417 2.2505
R42648 ASIG5V.n415 ASIG5V.n234 2.2505
R42649 ASIG5V.n423 ASIG5V.n422 2.2505
R42650 ASIG5V.n426 ASIG5V.n425 2.2505
R42651 ASIG5V.n430 ASIG5V.n429 2.2505
R42652 ASIG5V.n427 ASIG5V.n232 2.2505
R42653 ASIG5V.n435 ASIG5V.n434 2.2505
R42654 ASIG5V.n438 ASIG5V.n437 2.2505
R42655 ASIG5V.n442 ASIG5V.n441 2.2505
R42656 ASIG5V.n439 ASIG5V.n230 2.2505
R42657 ASIG5V.n447 ASIG5V.n446 2.2505
R42658 ASIG5V.n450 ASIG5V.n449 2.2505
R42659 ASIG5V.n454 ASIG5V.n453 2.2505
R42660 ASIG5V.n451 ASIG5V.n228 2.2505
R42661 ASIG5V.n459 ASIG5V.n458 2.2505
R42662 ASIG5V.n462 ASIG5V.n461 2.2505
R42663 ASIG5V.n466 ASIG5V.n465 2.2505
R42664 ASIG5V.n463 ASIG5V.n226 2.2505
R42665 ASIG5V.n471 ASIG5V.n470 2.2505
R42666 ASIG5V.n474 ASIG5V.n473 2.2505
R42667 ASIG5V.n478 ASIG5V.n477 2.2505
R42668 ASIG5V.n475 ASIG5V.n224 2.2505
R42669 ASIG5V.n483 ASIG5V.n482 2.2505
R42670 ASIG5V.n486 ASIG5V.n485 2.2505
R42671 ASIG5V.n490 ASIG5V.n489 2.2505
R42672 ASIG5V.n487 ASIG5V.n222 2.2505
R42673 ASIG5V.n495 ASIG5V.n494 2.2505
R42674 ASIG5V.n498 ASIG5V.n497 2.2505
R42675 ASIG5V.n502 ASIG5V.n501 2.2505
R42676 ASIG5V.n499 ASIG5V.n220 2.2505
R42677 ASIG5V.n12320 ASIG5V.n12319 2.2505
R42678 ASIG5V.n12322 ASIG5V.n218 2.2505
R42679 ASIG5V.n12295 ASIG5V.n573 2.2505
R42680 ASIG5V.n12297 ASIG5V.n12296 2.2505
R42681 ASIG5V.n858 ASIG5V.n574 2.2505
R42682 ASIG5V.n857 ASIG5V.n856 2.2505
R42683 ASIG5V.n852 ASIG5V.n575 2.2505
R42684 ASIG5V.n848 ASIG5V.n847 2.2505
R42685 ASIG5V.n846 ASIG5V.n576 2.2505
R42686 ASIG5V.n845 ASIG5V.n844 2.2505
R42687 ASIG5V.n840 ASIG5V.n577 2.2505
R42688 ASIG5V.n836 ASIG5V.n835 2.2505
R42689 ASIG5V.n834 ASIG5V.n578 2.2505
R42690 ASIG5V.n833 ASIG5V.n832 2.2505
R42691 ASIG5V.n828 ASIG5V.n579 2.2505
R42692 ASIG5V.n824 ASIG5V.n823 2.2505
R42693 ASIG5V.n822 ASIG5V.n580 2.2505
R42694 ASIG5V.n821 ASIG5V.n820 2.2505
R42695 ASIG5V.n816 ASIG5V.n581 2.2505
R42696 ASIG5V.n812 ASIG5V.n811 2.2505
R42697 ASIG5V.n810 ASIG5V.n582 2.2505
R42698 ASIG5V.n809 ASIG5V.n808 2.2505
R42699 ASIG5V.n804 ASIG5V.n583 2.2505
R42700 ASIG5V.n800 ASIG5V.n799 2.2505
R42701 ASIG5V.n798 ASIG5V.n584 2.2505
R42702 ASIG5V.n797 ASIG5V.n796 2.2505
R42703 ASIG5V.n792 ASIG5V.n585 2.2505
R42704 ASIG5V.n788 ASIG5V.n787 2.2505
R42705 ASIG5V.n786 ASIG5V.n586 2.2505
R42706 ASIG5V.n785 ASIG5V.n784 2.2505
R42707 ASIG5V.n780 ASIG5V.n587 2.2505
R42708 ASIG5V.n776 ASIG5V.n775 2.2505
R42709 ASIG5V.n774 ASIG5V.n588 2.2505
R42710 ASIG5V.n773 ASIG5V.n772 2.2505
R42711 ASIG5V.n768 ASIG5V.n589 2.2505
R42712 ASIG5V.n764 ASIG5V.n763 2.2505
R42713 ASIG5V.n762 ASIG5V.n590 2.2505
R42714 ASIG5V.n761 ASIG5V.n760 2.2505
R42715 ASIG5V.n756 ASIG5V.n591 2.2505
R42716 ASIG5V.n752 ASIG5V.n751 2.2505
R42717 ASIG5V.n750 ASIG5V.n592 2.2505
R42718 ASIG5V.n749 ASIG5V.n748 2.2505
R42719 ASIG5V.n744 ASIG5V.n593 2.2505
R42720 ASIG5V.n740 ASIG5V.n739 2.2505
R42721 ASIG5V.n738 ASIG5V.n594 2.2505
R42722 ASIG5V.n737 ASIG5V.n736 2.2505
R42723 ASIG5V.n732 ASIG5V.n595 2.2505
R42724 ASIG5V.n728 ASIG5V.n727 2.2505
R42725 ASIG5V.n726 ASIG5V.n596 2.2505
R42726 ASIG5V.n725 ASIG5V.n724 2.2505
R42727 ASIG5V.n720 ASIG5V.n597 2.2505
R42728 ASIG5V.n716 ASIG5V.n715 2.2505
R42729 ASIG5V.n714 ASIG5V.n598 2.2505
R42730 ASIG5V.n713 ASIG5V.n712 2.2505
R42731 ASIG5V.n708 ASIG5V.n599 2.2505
R42732 ASIG5V.n704 ASIG5V.n703 2.2505
R42733 ASIG5V.n702 ASIG5V.n600 2.2505
R42734 ASIG5V.n701 ASIG5V.n700 2.2505
R42735 ASIG5V.n696 ASIG5V.n601 2.2505
R42736 ASIG5V.n692 ASIG5V.n691 2.2505
R42737 ASIG5V.n690 ASIG5V.n602 2.2505
R42738 ASIG5V.n689 ASIG5V.n688 2.2505
R42739 ASIG5V.n684 ASIG5V.n603 2.2505
R42740 ASIG5V.n680 ASIG5V.n679 2.2505
R42741 ASIG5V.n678 ASIG5V.n604 2.2505
R42742 ASIG5V.n677 ASIG5V.n676 2.2505
R42743 ASIG5V.n672 ASIG5V.n605 2.2505
R42744 ASIG5V.n668 ASIG5V.n667 2.2505
R42745 ASIG5V.n666 ASIG5V.n606 2.2505
R42746 ASIG5V.n665 ASIG5V.n664 2.2505
R42747 ASIG5V.n660 ASIG5V.n607 2.2505
R42748 ASIG5V.n656 ASIG5V.n655 2.2505
R42749 ASIG5V.n654 ASIG5V.n608 2.2505
R42750 ASIG5V.n653 ASIG5V.n652 2.2505
R42751 ASIG5V.n648 ASIG5V.n609 2.2505
R42752 ASIG5V.n644 ASIG5V.n643 2.2505
R42753 ASIG5V.n642 ASIG5V.n610 2.2505
R42754 ASIG5V.n641 ASIG5V.n640 2.2505
R42755 ASIG5V.n636 ASIG5V.n611 2.2505
R42756 ASIG5V.n632 ASIG5V.n631 2.2505
R42757 ASIG5V.n630 ASIG5V.n612 2.2505
R42758 ASIG5V.n629 ASIG5V.n628 2.2505
R42759 ASIG5V.n624 ASIG5V.n613 2.2505
R42760 ASIG5V.n620 ASIG5V.n619 2.2505
R42761 ASIG5V.n618 ASIG5V.n617 2.2505
R42762 ASIG5V.n614 ASIG5V.n524 2.2505
R42763 ASIG5V.n614 ASIG5V.n570 2.2505
R42764 ASIG5V.n617 ASIG5V.n616 2.2505
R42765 ASIG5V.n621 ASIG5V.n620 2.2505
R42766 ASIG5V.n624 ASIG5V.n623 2.2505
R42767 ASIG5V.n628 ASIG5V.n627 2.2505
R42768 ASIG5V.n625 ASIG5V.n612 2.2505
R42769 ASIG5V.n633 ASIG5V.n632 2.2505
R42770 ASIG5V.n636 ASIG5V.n635 2.2505
R42771 ASIG5V.n640 ASIG5V.n639 2.2505
R42772 ASIG5V.n637 ASIG5V.n610 2.2505
R42773 ASIG5V.n645 ASIG5V.n644 2.2505
R42774 ASIG5V.n648 ASIG5V.n647 2.2505
R42775 ASIG5V.n652 ASIG5V.n651 2.2505
R42776 ASIG5V.n649 ASIG5V.n608 2.2505
R42777 ASIG5V.n657 ASIG5V.n656 2.2505
R42778 ASIG5V.n660 ASIG5V.n659 2.2505
R42779 ASIG5V.n664 ASIG5V.n663 2.2505
R42780 ASIG5V.n661 ASIG5V.n606 2.2505
R42781 ASIG5V.n669 ASIG5V.n668 2.2505
R42782 ASIG5V.n672 ASIG5V.n671 2.2505
R42783 ASIG5V.n676 ASIG5V.n675 2.2505
R42784 ASIG5V.n673 ASIG5V.n604 2.2505
R42785 ASIG5V.n681 ASIG5V.n680 2.2505
R42786 ASIG5V.n684 ASIG5V.n683 2.2505
R42787 ASIG5V.n688 ASIG5V.n687 2.2505
R42788 ASIG5V.n685 ASIG5V.n602 2.2505
R42789 ASIG5V.n693 ASIG5V.n692 2.2505
R42790 ASIG5V.n696 ASIG5V.n695 2.2505
R42791 ASIG5V.n700 ASIG5V.n699 2.2505
R42792 ASIG5V.n697 ASIG5V.n600 2.2505
R42793 ASIG5V.n705 ASIG5V.n704 2.2505
R42794 ASIG5V.n708 ASIG5V.n707 2.2505
R42795 ASIG5V.n712 ASIG5V.n711 2.2505
R42796 ASIG5V.n709 ASIG5V.n598 2.2505
R42797 ASIG5V.n717 ASIG5V.n716 2.2505
R42798 ASIG5V.n720 ASIG5V.n719 2.2505
R42799 ASIG5V.n724 ASIG5V.n723 2.2505
R42800 ASIG5V.n721 ASIG5V.n596 2.2505
R42801 ASIG5V.n729 ASIG5V.n728 2.2505
R42802 ASIG5V.n732 ASIG5V.n731 2.2505
R42803 ASIG5V.n736 ASIG5V.n735 2.2505
R42804 ASIG5V.n733 ASIG5V.n594 2.2505
R42805 ASIG5V.n741 ASIG5V.n740 2.2505
R42806 ASIG5V.n744 ASIG5V.n743 2.2505
R42807 ASIG5V.n748 ASIG5V.n747 2.2505
R42808 ASIG5V.n745 ASIG5V.n592 2.2505
R42809 ASIG5V.n753 ASIG5V.n752 2.2505
R42810 ASIG5V.n756 ASIG5V.n755 2.2505
R42811 ASIG5V.n760 ASIG5V.n759 2.2505
R42812 ASIG5V.n757 ASIG5V.n590 2.2505
R42813 ASIG5V.n765 ASIG5V.n764 2.2505
R42814 ASIG5V.n768 ASIG5V.n767 2.2505
R42815 ASIG5V.n772 ASIG5V.n771 2.2505
R42816 ASIG5V.n769 ASIG5V.n588 2.2505
R42817 ASIG5V.n777 ASIG5V.n776 2.2505
R42818 ASIG5V.n780 ASIG5V.n779 2.2505
R42819 ASIG5V.n784 ASIG5V.n783 2.2505
R42820 ASIG5V.n781 ASIG5V.n586 2.2505
R42821 ASIG5V.n789 ASIG5V.n788 2.2505
R42822 ASIG5V.n792 ASIG5V.n791 2.2505
R42823 ASIG5V.n796 ASIG5V.n795 2.2505
R42824 ASIG5V.n793 ASIG5V.n584 2.2505
R42825 ASIG5V.n801 ASIG5V.n800 2.2505
R42826 ASIG5V.n804 ASIG5V.n803 2.2505
R42827 ASIG5V.n808 ASIG5V.n807 2.2505
R42828 ASIG5V.n805 ASIG5V.n582 2.2505
R42829 ASIG5V.n813 ASIG5V.n812 2.2505
R42830 ASIG5V.n816 ASIG5V.n815 2.2505
R42831 ASIG5V.n820 ASIG5V.n819 2.2505
R42832 ASIG5V.n817 ASIG5V.n580 2.2505
R42833 ASIG5V.n825 ASIG5V.n824 2.2505
R42834 ASIG5V.n828 ASIG5V.n827 2.2505
R42835 ASIG5V.n832 ASIG5V.n831 2.2505
R42836 ASIG5V.n829 ASIG5V.n578 2.2505
R42837 ASIG5V.n837 ASIG5V.n836 2.2505
R42838 ASIG5V.n840 ASIG5V.n839 2.2505
R42839 ASIG5V.n844 ASIG5V.n843 2.2505
R42840 ASIG5V.n841 ASIG5V.n576 2.2505
R42841 ASIG5V.n849 ASIG5V.n848 2.2505
R42842 ASIG5V.n852 ASIG5V.n851 2.2505
R42843 ASIG5V.n856 ASIG5V.n855 2.2505
R42844 ASIG5V.n853 ASIG5V.n574 2.2505
R42845 ASIG5V.n12298 ASIG5V.n12297 2.2505
R42846 ASIG5V.n12300 ASIG5V.n573 2.2505
R42847 ASIG5V.n1216 ASIG5V.n1215 2.2505
R42848 ASIG5V.n884 ASIG5V.n883 2.2505
R42849 ASIG5V.n1205 ASIG5V.n885 2.2505
R42850 ASIG5V.n1207 ASIG5V.n1206 2.2505
R42851 ASIG5V.n1204 ASIG5V.n887 2.2505
R42852 ASIG5V.n1203 ASIG5V.n1202 2.2505
R42853 ASIG5V.n889 ASIG5V.n888 2.2505
R42854 ASIG5V.n1194 ASIG5V.n1193 2.2505
R42855 ASIG5V.n1192 ASIG5V.n891 2.2505
R42856 ASIG5V.n1191 ASIG5V.n1190 2.2505
R42857 ASIG5V.n893 ASIG5V.n892 2.2505
R42858 ASIG5V.n1182 ASIG5V.n1181 2.2505
R42859 ASIG5V.n1180 ASIG5V.n895 2.2505
R42860 ASIG5V.n1179 ASIG5V.n1178 2.2505
R42861 ASIG5V.n897 ASIG5V.n896 2.2505
R42862 ASIG5V.n1170 ASIG5V.n1169 2.2505
R42863 ASIG5V.n1168 ASIG5V.n899 2.2505
R42864 ASIG5V.n1167 ASIG5V.n1166 2.2505
R42865 ASIG5V.n901 ASIG5V.n900 2.2505
R42866 ASIG5V.n1158 ASIG5V.n1157 2.2505
R42867 ASIG5V.n1156 ASIG5V.n903 2.2505
R42868 ASIG5V.n1155 ASIG5V.n1154 2.2505
R42869 ASIG5V.n905 ASIG5V.n904 2.2505
R42870 ASIG5V.n1146 ASIG5V.n1145 2.2505
R42871 ASIG5V.n1144 ASIG5V.n907 2.2505
R42872 ASIG5V.n1143 ASIG5V.n1142 2.2505
R42873 ASIG5V.n909 ASIG5V.n908 2.2505
R42874 ASIG5V.n1134 ASIG5V.n1133 2.2505
R42875 ASIG5V.n1132 ASIG5V.n911 2.2505
R42876 ASIG5V.n1131 ASIG5V.n1130 2.2505
R42877 ASIG5V.n913 ASIG5V.n912 2.2505
R42878 ASIG5V.n1122 ASIG5V.n1121 2.2505
R42879 ASIG5V.n1120 ASIG5V.n915 2.2505
R42880 ASIG5V.n1119 ASIG5V.n1118 2.2505
R42881 ASIG5V.n917 ASIG5V.n916 2.2505
R42882 ASIG5V.n1110 ASIG5V.n1109 2.2505
R42883 ASIG5V.n1108 ASIG5V.n919 2.2505
R42884 ASIG5V.n1107 ASIG5V.n1106 2.2505
R42885 ASIG5V.n921 ASIG5V.n920 2.2505
R42886 ASIG5V.n1098 ASIG5V.n1097 2.2505
R42887 ASIG5V.n1096 ASIG5V.n923 2.2505
R42888 ASIG5V.n1095 ASIG5V.n1094 2.2505
R42889 ASIG5V.n925 ASIG5V.n924 2.2505
R42890 ASIG5V.n1086 ASIG5V.n1085 2.2505
R42891 ASIG5V.n1084 ASIG5V.n927 2.2505
R42892 ASIG5V.n1083 ASIG5V.n1082 2.2505
R42893 ASIG5V.n929 ASIG5V.n928 2.2505
R42894 ASIG5V.n1074 ASIG5V.n1073 2.2505
R42895 ASIG5V.n1072 ASIG5V.n931 2.2505
R42896 ASIG5V.n1071 ASIG5V.n1070 2.2505
R42897 ASIG5V.n933 ASIG5V.n932 2.2505
R42898 ASIG5V.n1062 ASIG5V.n1061 2.2505
R42899 ASIG5V.n1060 ASIG5V.n935 2.2505
R42900 ASIG5V.n1059 ASIG5V.n1058 2.2505
R42901 ASIG5V.n937 ASIG5V.n936 2.2505
R42902 ASIG5V.n1050 ASIG5V.n1049 2.2505
R42903 ASIG5V.n1048 ASIG5V.n939 2.2505
R42904 ASIG5V.n1047 ASIG5V.n1046 2.2505
R42905 ASIG5V.n941 ASIG5V.n940 2.2505
R42906 ASIG5V.n1038 ASIG5V.n1037 2.2505
R42907 ASIG5V.n1036 ASIG5V.n943 2.2505
R42908 ASIG5V.n1035 ASIG5V.n1034 2.2505
R42909 ASIG5V.n945 ASIG5V.n944 2.2505
R42910 ASIG5V.n1026 ASIG5V.n1025 2.2505
R42911 ASIG5V.n1024 ASIG5V.n947 2.2505
R42912 ASIG5V.n1023 ASIG5V.n1022 2.2505
R42913 ASIG5V.n949 ASIG5V.n948 2.2505
R42914 ASIG5V.n1014 ASIG5V.n1013 2.2505
R42915 ASIG5V.n1012 ASIG5V.n951 2.2505
R42916 ASIG5V.n1011 ASIG5V.n1010 2.2505
R42917 ASIG5V.n953 ASIG5V.n952 2.2505
R42918 ASIG5V.n1002 ASIG5V.n1001 2.2505
R42919 ASIG5V.n1000 ASIG5V.n955 2.2505
R42920 ASIG5V.n999 ASIG5V.n998 2.2505
R42921 ASIG5V.n957 ASIG5V.n956 2.2505
R42922 ASIG5V.n990 ASIG5V.n989 2.2505
R42923 ASIG5V.n988 ASIG5V.n959 2.2505
R42924 ASIG5V.n987 ASIG5V.n986 2.2505
R42925 ASIG5V.n961 ASIG5V.n960 2.2505
R42926 ASIG5V.n978 ASIG5V.n977 2.2505
R42927 ASIG5V.n976 ASIG5V.n963 2.2505
R42928 ASIG5V.n975 ASIG5V.n974 2.2505
R42929 ASIG5V.n965 ASIG5V.n964 2.2505
R42930 ASIG5V.n966 ASIG5V.n869 2.2505
R42931 ASIG5V.n967 ASIG5V.n966 2.2505
R42932 ASIG5V.n969 ASIG5V.n965 2.2505
R42933 ASIG5V.n974 ASIG5V.n973 2.2505
R42934 ASIG5V.n971 ASIG5V.n963 2.2505
R42935 ASIG5V.n979 ASIG5V.n978 2.2505
R42936 ASIG5V.n981 ASIG5V.n961 2.2505
R42937 ASIG5V.n986 ASIG5V.n985 2.2505
R42938 ASIG5V.n983 ASIG5V.n959 2.2505
R42939 ASIG5V.n991 ASIG5V.n990 2.2505
R42940 ASIG5V.n993 ASIG5V.n957 2.2505
R42941 ASIG5V.n998 ASIG5V.n997 2.2505
R42942 ASIG5V.n995 ASIG5V.n955 2.2505
R42943 ASIG5V.n1003 ASIG5V.n1002 2.2505
R42944 ASIG5V.n1005 ASIG5V.n953 2.2505
R42945 ASIG5V.n1010 ASIG5V.n1009 2.2505
R42946 ASIG5V.n1007 ASIG5V.n951 2.2505
R42947 ASIG5V.n1015 ASIG5V.n1014 2.2505
R42948 ASIG5V.n1017 ASIG5V.n949 2.2505
R42949 ASIG5V.n1022 ASIG5V.n1021 2.2505
R42950 ASIG5V.n1019 ASIG5V.n947 2.2505
R42951 ASIG5V.n1027 ASIG5V.n1026 2.2505
R42952 ASIG5V.n1029 ASIG5V.n945 2.2505
R42953 ASIG5V.n1034 ASIG5V.n1033 2.2505
R42954 ASIG5V.n1031 ASIG5V.n943 2.2505
R42955 ASIG5V.n1039 ASIG5V.n1038 2.2505
R42956 ASIG5V.n1041 ASIG5V.n941 2.2505
R42957 ASIG5V.n1046 ASIG5V.n1045 2.2505
R42958 ASIG5V.n1043 ASIG5V.n939 2.2505
R42959 ASIG5V.n1051 ASIG5V.n1050 2.2505
R42960 ASIG5V.n1053 ASIG5V.n937 2.2505
R42961 ASIG5V.n1058 ASIG5V.n1057 2.2505
R42962 ASIG5V.n1055 ASIG5V.n935 2.2505
R42963 ASIG5V.n1063 ASIG5V.n1062 2.2505
R42964 ASIG5V.n1065 ASIG5V.n933 2.2505
R42965 ASIG5V.n1070 ASIG5V.n1069 2.2505
R42966 ASIG5V.n1067 ASIG5V.n931 2.2505
R42967 ASIG5V.n1075 ASIG5V.n1074 2.2505
R42968 ASIG5V.n1077 ASIG5V.n929 2.2505
R42969 ASIG5V.n1082 ASIG5V.n1081 2.2505
R42970 ASIG5V.n1079 ASIG5V.n927 2.2505
R42971 ASIG5V.n1087 ASIG5V.n1086 2.2505
R42972 ASIG5V.n1089 ASIG5V.n925 2.2505
R42973 ASIG5V.n1094 ASIG5V.n1093 2.2505
R42974 ASIG5V.n1091 ASIG5V.n923 2.2505
R42975 ASIG5V.n1099 ASIG5V.n1098 2.2505
R42976 ASIG5V.n1101 ASIG5V.n921 2.2505
R42977 ASIG5V.n1106 ASIG5V.n1105 2.2505
R42978 ASIG5V.n1103 ASIG5V.n919 2.2505
R42979 ASIG5V.n1111 ASIG5V.n1110 2.2505
R42980 ASIG5V.n1113 ASIG5V.n917 2.2505
R42981 ASIG5V.n1118 ASIG5V.n1117 2.2505
R42982 ASIG5V.n1115 ASIG5V.n915 2.2505
R42983 ASIG5V.n1123 ASIG5V.n1122 2.2505
R42984 ASIG5V.n1125 ASIG5V.n913 2.2505
R42985 ASIG5V.n1130 ASIG5V.n1129 2.2505
R42986 ASIG5V.n1127 ASIG5V.n911 2.2505
R42987 ASIG5V.n1135 ASIG5V.n1134 2.2505
R42988 ASIG5V.n1137 ASIG5V.n909 2.2505
R42989 ASIG5V.n1142 ASIG5V.n1141 2.2505
R42990 ASIG5V.n1139 ASIG5V.n907 2.2505
R42991 ASIG5V.n1147 ASIG5V.n1146 2.2505
R42992 ASIG5V.n1149 ASIG5V.n905 2.2505
R42993 ASIG5V.n1154 ASIG5V.n1153 2.2505
R42994 ASIG5V.n1151 ASIG5V.n903 2.2505
R42995 ASIG5V.n1159 ASIG5V.n1158 2.2505
R42996 ASIG5V.n1161 ASIG5V.n901 2.2505
R42997 ASIG5V.n1166 ASIG5V.n1165 2.2505
R42998 ASIG5V.n1163 ASIG5V.n899 2.2505
R42999 ASIG5V.n1171 ASIG5V.n1170 2.2505
R43000 ASIG5V.n1173 ASIG5V.n897 2.2505
R43001 ASIG5V.n1178 ASIG5V.n1177 2.2505
R43002 ASIG5V.n1175 ASIG5V.n895 2.2505
R43003 ASIG5V.n1183 ASIG5V.n1182 2.2505
R43004 ASIG5V.n1185 ASIG5V.n893 2.2505
R43005 ASIG5V.n1190 ASIG5V.n1189 2.2505
R43006 ASIG5V.n1187 ASIG5V.n891 2.2505
R43007 ASIG5V.n1195 ASIG5V.n1194 2.2505
R43008 ASIG5V.n1197 ASIG5V.n889 2.2505
R43009 ASIG5V.n1202 ASIG5V.n1201 2.2505
R43010 ASIG5V.n1199 ASIG5V.n887 2.2505
R43011 ASIG5V.n1208 ASIG5V.n1207 2.2505
R43012 ASIG5V.n1210 ASIG5V.n885 2.2505
R43013 ASIG5V.n1212 ASIG5V.n884 2.2505
R43014 ASIG5V.n1215 ASIG5V.n1214 2.2505
R43015 ASIG5V.n1270 ASIG5V.n1220 2.2505
R43016 ASIG5V.n12264 ASIG5V.n12263 2.2505
R43017 ASIG5V.n12262 ASIG5V.n1273 2.2505
R43018 ASIG5V.n12261 ASIG5V.n12260 2.2505
R43019 ASIG5V.n12256 ASIG5V.n1274 2.2505
R43020 ASIG5V.n12252 ASIG5V.n12251 2.2505
R43021 ASIG5V.n12250 ASIG5V.n1275 2.2505
R43022 ASIG5V.n12249 ASIG5V.n12248 2.2505
R43023 ASIG5V.n12244 ASIG5V.n1276 2.2505
R43024 ASIG5V.n12240 ASIG5V.n12239 2.2505
R43025 ASIG5V.n12238 ASIG5V.n1277 2.2505
R43026 ASIG5V.n12237 ASIG5V.n12236 2.2505
R43027 ASIG5V.n12232 ASIG5V.n1278 2.2505
R43028 ASIG5V.n12228 ASIG5V.n12227 2.2505
R43029 ASIG5V.n12226 ASIG5V.n1279 2.2505
R43030 ASIG5V.n12225 ASIG5V.n12224 2.2505
R43031 ASIG5V.n12220 ASIG5V.n1280 2.2505
R43032 ASIG5V.n12216 ASIG5V.n12215 2.2505
R43033 ASIG5V.n12214 ASIG5V.n1281 2.2505
R43034 ASIG5V.n12213 ASIG5V.n12212 2.2505
R43035 ASIG5V.n12208 ASIG5V.n1282 2.2505
R43036 ASIG5V.n12204 ASIG5V.n12203 2.2505
R43037 ASIG5V.n12202 ASIG5V.n1283 2.2505
R43038 ASIG5V.n12201 ASIG5V.n12200 2.2505
R43039 ASIG5V.n12196 ASIG5V.n1284 2.2505
R43040 ASIG5V.n12192 ASIG5V.n12191 2.2505
R43041 ASIG5V.n12190 ASIG5V.n1285 2.2505
R43042 ASIG5V.n12189 ASIG5V.n12188 2.2505
R43043 ASIG5V.n12184 ASIG5V.n1286 2.2505
R43044 ASIG5V.n12180 ASIG5V.n12179 2.2505
R43045 ASIG5V.n12178 ASIG5V.n1287 2.2505
R43046 ASIG5V.n12177 ASIG5V.n12176 2.2505
R43047 ASIG5V.n12172 ASIG5V.n1288 2.2505
R43048 ASIG5V.n12168 ASIG5V.n12167 2.2505
R43049 ASIG5V.n12166 ASIG5V.n1289 2.2505
R43050 ASIG5V.n12165 ASIG5V.n12164 2.2505
R43051 ASIG5V.n12160 ASIG5V.n1290 2.2505
R43052 ASIG5V.n12156 ASIG5V.n12155 2.2505
R43053 ASIG5V.n12154 ASIG5V.n1291 2.2505
R43054 ASIG5V.n12153 ASIG5V.n12152 2.2505
R43055 ASIG5V.n12148 ASIG5V.n1292 2.2505
R43056 ASIG5V.n12144 ASIG5V.n12143 2.2505
R43057 ASIG5V.n12142 ASIG5V.n1293 2.2505
R43058 ASIG5V.n12141 ASIG5V.n12140 2.2505
R43059 ASIG5V.n12136 ASIG5V.n1294 2.2505
R43060 ASIG5V.n12132 ASIG5V.n12131 2.2505
R43061 ASIG5V.n12130 ASIG5V.n1295 2.2505
R43062 ASIG5V.n12129 ASIG5V.n12128 2.2505
R43063 ASIG5V.n12124 ASIG5V.n1296 2.2505
R43064 ASIG5V.n12120 ASIG5V.n12119 2.2505
R43065 ASIG5V.n12118 ASIG5V.n1297 2.2505
R43066 ASIG5V.n12117 ASIG5V.n12116 2.2505
R43067 ASIG5V.n12112 ASIG5V.n1298 2.2505
R43068 ASIG5V.n12108 ASIG5V.n12107 2.2505
R43069 ASIG5V.n12106 ASIG5V.n1299 2.2505
R43070 ASIG5V.n12105 ASIG5V.n12104 2.2505
R43071 ASIG5V.n12100 ASIG5V.n1300 2.2505
R43072 ASIG5V.n12096 ASIG5V.n12095 2.2505
R43073 ASIG5V.n12094 ASIG5V.n1301 2.2505
R43074 ASIG5V.n12093 ASIG5V.n12092 2.2505
R43075 ASIG5V.n12088 ASIG5V.n1302 2.2505
R43076 ASIG5V.n12084 ASIG5V.n12083 2.2505
R43077 ASIG5V.n12082 ASIG5V.n1303 2.2505
R43078 ASIG5V.n12081 ASIG5V.n12080 2.2505
R43079 ASIG5V.n12076 ASIG5V.n1304 2.2505
R43080 ASIG5V.n12072 ASIG5V.n12071 2.2505
R43081 ASIG5V.n12070 ASIG5V.n1305 2.2505
R43082 ASIG5V.n12069 ASIG5V.n12068 2.2505
R43083 ASIG5V.n12064 ASIG5V.n1306 2.2505
R43084 ASIG5V.n12060 ASIG5V.n12059 2.2505
R43085 ASIG5V.n12058 ASIG5V.n1307 2.2505
R43086 ASIG5V.n12057 ASIG5V.n12056 2.2505
R43087 ASIG5V.n12052 ASIG5V.n1308 2.2505
R43088 ASIG5V.n12048 ASIG5V.n12047 2.2505
R43089 ASIG5V.n12046 ASIG5V.n1309 2.2505
R43090 ASIG5V.n12045 ASIG5V.n12044 2.2505
R43091 ASIG5V.n12040 ASIG5V.n1310 2.2505
R43092 ASIG5V.n12036 ASIG5V.n12035 2.2505
R43093 ASIG5V.n12034 ASIG5V.n1311 2.2505
R43094 ASIG5V.n12033 ASIG5V.n12032 2.2505
R43095 ASIG5V.n12028 ASIG5V.n1312 2.2505
R43096 ASIG5V.n12024 ASIG5V.n12023 2.2505
R43097 ASIG5V.n12022 ASIG5V.n1315 2.2505
R43098 ASIG5V.n12021 ASIG5V.n12020 2.2505
R43099 ASIG5V.n12020 ASIG5V.n1268 2.2505
R43100 ASIG5V.n1315 ASIG5V.n1314 2.2505
R43101 ASIG5V.n12025 ASIG5V.n12024 2.2505
R43102 ASIG5V.n12028 ASIG5V.n12027 2.2505
R43103 ASIG5V.n12032 ASIG5V.n12031 2.2505
R43104 ASIG5V.n12029 ASIG5V.n1311 2.2505
R43105 ASIG5V.n12037 ASIG5V.n12036 2.2505
R43106 ASIG5V.n12040 ASIG5V.n12039 2.2505
R43107 ASIG5V.n12044 ASIG5V.n12043 2.2505
R43108 ASIG5V.n12041 ASIG5V.n1309 2.2505
R43109 ASIG5V.n12049 ASIG5V.n12048 2.2505
R43110 ASIG5V.n12052 ASIG5V.n12051 2.2505
R43111 ASIG5V.n12056 ASIG5V.n12055 2.2505
R43112 ASIG5V.n12053 ASIG5V.n1307 2.2505
R43113 ASIG5V.n12061 ASIG5V.n12060 2.2505
R43114 ASIG5V.n12064 ASIG5V.n12063 2.2505
R43115 ASIG5V.n12068 ASIG5V.n12067 2.2505
R43116 ASIG5V.n12065 ASIG5V.n1305 2.2505
R43117 ASIG5V.n12073 ASIG5V.n12072 2.2505
R43118 ASIG5V.n12076 ASIG5V.n12075 2.2505
R43119 ASIG5V.n12080 ASIG5V.n12079 2.2505
R43120 ASIG5V.n12077 ASIG5V.n1303 2.2505
R43121 ASIG5V.n12085 ASIG5V.n12084 2.2505
R43122 ASIG5V.n12088 ASIG5V.n12087 2.2505
R43123 ASIG5V.n12092 ASIG5V.n12091 2.2505
R43124 ASIG5V.n12089 ASIG5V.n1301 2.2505
R43125 ASIG5V.n12097 ASIG5V.n12096 2.2505
R43126 ASIG5V.n12100 ASIG5V.n12099 2.2505
R43127 ASIG5V.n12104 ASIG5V.n12103 2.2505
R43128 ASIG5V.n12101 ASIG5V.n1299 2.2505
R43129 ASIG5V.n12109 ASIG5V.n12108 2.2505
R43130 ASIG5V.n12112 ASIG5V.n12111 2.2505
R43131 ASIG5V.n12116 ASIG5V.n12115 2.2505
R43132 ASIG5V.n12113 ASIG5V.n1297 2.2505
R43133 ASIG5V.n12121 ASIG5V.n12120 2.2505
R43134 ASIG5V.n12124 ASIG5V.n12123 2.2505
R43135 ASIG5V.n12128 ASIG5V.n12127 2.2505
R43136 ASIG5V.n12125 ASIG5V.n1295 2.2505
R43137 ASIG5V.n12133 ASIG5V.n12132 2.2505
R43138 ASIG5V.n12136 ASIG5V.n12135 2.2505
R43139 ASIG5V.n12140 ASIG5V.n12139 2.2505
R43140 ASIG5V.n12137 ASIG5V.n1293 2.2505
R43141 ASIG5V.n12145 ASIG5V.n12144 2.2505
R43142 ASIG5V.n12148 ASIG5V.n12147 2.2505
R43143 ASIG5V.n12152 ASIG5V.n12151 2.2505
R43144 ASIG5V.n12149 ASIG5V.n1291 2.2505
R43145 ASIG5V.n12157 ASIG5V.n12156 2.2505
R43146 ASIG5V.n12160 ASIG5V.n12159 2.2505
R43147 ASIG5V.n12164 ASIG5V.n12163 2.2505
R43148 ASIG5V.n12161 ASIG5V.n1289 2.2505
R43149 ASIG5V.n12169 ASIG5V.n12168 2.2505
R43150 ASIG5V.n12172 ASIG5V.n12171 2.2505
R43151 ASIG5V.n12176 ASIG5V.n12175 2.2505
R43152 ASIG5V.n12173 ASIG5V.n1287 2.2505
R43153 ASIG5V.n12181 ASIG5V.n12180 2.2505
R43154 ASIG5V.n12184 ASIG5V.n12183 2.2505
R43155 ASIG5V.n12188 ASIG5V.n12187 2.2505
R43156 ASIG5V.n12185 ASIG5V.n1285 2.2505
R43157 ASIG5V.n12193 ASIG5V.n12192 2.2505
R43158 ASIG5V.n12196 ASIG5V.n12195 2.2505
R43159 ASIG5V.n12200 ASIG5V.n12199 2.2505
R43160 ASIG5V.n12197 ASIG5V.n1283 2.2505
R43161 ASIG5V.n12205 ASIG5V.n12204 2.2505
R43162 ASIG5V.n12208 ASIG5V.n12207 2.2505
R43163 ASIG5V.n12212 ASIG5V.n12211 2.2505
R43164 ASIG5V.n12209 ASIG5V.n1281 2.2505
R43165 ASIG5V.n12217 ASIG5V.n12216 2.2505
R43166 ASIG5V.n12220 ASIG5V.n12219 2.2505
R43167 ASIG5V.n12224 ASIG5V.n12223 2.2505
R43168 ASIG5V.n12221 ASIG5V.n1279 2.2505
R43169 ASIG5V.n12229 ASIG5V.n12228 2.2505
R43170 ASIG5V.n12232 ASIG5V.n12231 2.2505
R43171 ASIG5V.n12236 ASIG5V.n12235 2.2505
R43172 ASIG5V.n12233 ASIG5V.n1277 2.2505
R43173 ASIG5V.n12241 ASIG5V.n12240 2.2505
R43174 ASIG5V.n12244 ASIG5V.n12243 2.2505
R43175 ASIG5V.n12248 ASIG5V.n12247 2.2505
R43176 ASIG5V.n12245 ASIG5V.n1275 2.2505
R43177 ASIG5V.n12253 ASIG5V.n12252 2.2505
R43178 ASIG5V.n12256 ASIG5V.n12255 2.2505
R43179 ASIG5V.n12260 ASIG5V.n12259 2.2505
R43180 ASIG5V.n12257 ASIG5V.n1273 2.2505
R43181 ASIG5V.n12265 ASIG5V.n12264 2.2505
R43182 ASIG5V.n12267 ASIG5V.n1270 2.2505
R43183 ASIG5V.n12006 ASIG5V.n1663 2.2505
R43184 ASIG5V.n1662 ASIG5V.n1418 2.2505
R43185 ASIG5V.n1661 ASIG5V.n1660 2.2505
R43186 ASIG5V.n1658 ASIG5V.n1419 2.2505
R43187 ASIG5V.n1656 ASIG5V.n1654 2.2505
R43188 ASIG5V.n1653 ASIG5V.n1421 2.2505
R43189 ASIG5V.n1652 ASIG5V.n1651 2.2505
R43190 ASIG5V.n1649 ASIG5V.n1422 2.2505
R43191 ASIG5V.n1647 ASIG5V.n1645 2.2505
R43192 ASIG5V.n1644 ASIG5V.n1424 2.2505
R43193 ASIG5V.n1643 ASIG5V.n1642 2.2505
R43194 ASIG5V.n1640 ASIG5V.n1425 2.2505
R43195 ASIG5V.n1638 ASIG5V.n1636 2.2505
R43196 ASIG5V.n1635 ASIG5V.n1427 2.2505
R43197 ASIG5V.n1634 ASIG5V.n1633 2.2505
R43198 ASIG5V.n1631 ASIG5V.n1428 2.2505
R43199 ASIG5V.n1629 ASIG5V.n1627 2.2505
R43200 ASIG5V.n1626 ASIG5V.n1430 2.2505
R43201 ASIG5V.n1625 ASIG5V.n1624 2.2505
R43202 ASIG5V.n1622 ASIG5V.n1431 2.2505
R43203 ASIG5V.n1620 ASIG5V.n1618 2.2505
R43204 ASIG5V.n1617 ASIG5V.n1433 2.2505
R43205 ASIG5V.n1616 ASIG5V.n1615 2.2505
R43206 ASIG5V.n1613 ASIG5V.n1434 2.2505
R43207 ASIG5V.n1611 ASIG5V.n1609 2.2505
R43208 ASIG5V.n1608 ASIG5V.n1436 2.2505
R43209 ASIG5V.n1607 ASIG5V.n1606 2.2505
R43210 ASIG5V.n1604 ASIG5V.n1437 2.2505
R43211 ASIG5V.n1602 ASIG5V.n1600 2.2505
R43212 ASIG5V.n1599 ASIG5V.n1439 2.2505
R43213 ASIG5V.n1598 ASIG5V.n1597 2.2505
R43214 ASIG5V.n1595 ASIG5V.n1440 2.2505
R43215 ASIG5V.n1593 ASIG5V.n1591 2.2505
R43216 ASIG5V.n1590 ASIG5V.n1442 2.2505
R43217 ASIG5V.n1589 ASIG5V.n1588 2.2505
R43218 ASIG5V.n1586 ASIG5V.n1443 2.2505
R43219 ASIG5V.n1584 ASIG5V.n1582 2.2505
R43220 ASIG5V.n1581 ASIG5V.n1445 2.2505
R43221 ASIG5V.n1580 ASIG5V.n1579 2.2505
R43222 ASIG5V.n1577 ASIG5V.n1446 2.2505
R43223 ASIG5V.n1575 ASIG5V.n1573 2.2505
R43224 ASIG5V.n1572 ASIG5V.n1448 2.2505
R43225 ASIG5V.n1571 ASIG5V.n1570 2.2505
R43226 ASIG5V.n1568 ASIG5V.n1449 2.2505
R43227 ASIG5V.n1566 ASIG5V.n1564 2.2505
R43228 ASIG5V.n1563 ASIG5V.n1451 2.2505
R43229 ASIG5V.n1562 ASIG5V.n1561 2.2505
R43230 ASIG5V.n1559 ASIG5V.n1452 2.2505
R43231 ASIG5V.n1557 ASIG5V.n1555 2.2505
R43232 ASIG5V.n1554 ASIG5V.n1454 2.2505
R43233 ASIG5V.n1553 ASIG5V.n1552 2.2505
R43234 ASIG5V.n1550 ASIG5V.n1455 2.2505
R43235 ASIG5V.n1548 ASIG5V.n1546 2.2505
R43236 ASIG5V.n1545 ASIG5V.n1457 2.2505
R43237 ASIG5V.n1544 ASIG5V.n1543 2.2505
R43238 ASIG5V.n1541 ASIG5V.n1458 2.2505
R43239 ASIG5V.n1539 ASIG5V.n1537 2.2505
R43240 ASIG5V.n1536 ASIG5V.n1460 2.2505
R43241 ASIG5V.n1535 ASIG5V.n1534 2.2505
R43242 ASIG5V.n1532 ASIG5V.n1461 2.2505
R43243 ASIG5V.n1530 ASIG5V.n1528 2.2505
R43244 ASIG5V.n1527 ASIG5V.n1463 2.2505
R43245 ASIG5V.n1526 ASIG5V.n1525 2.2505
R43246 ASIG5V.n1523 ASIG5V.n1464 2.2505
R43247 ASIG5V.n1521 ASIG5V.n1519 2.2505
R43248 ASIG5V.n1518 ASIG5V.n1466 2.2505
R43249 ASIG5V.n1517 ASIG5V.n1516 2.2505
R43250 ASIG5V.n1514 ASIG5V.n1467 2.2505
R43251 ASIG5V.n1512 ASIG5V.n1510 2.2505
R43252 ASIG5V.n1509 ASIG5V.n1469 2.2505
R43253 ASIG5V.n1508 ASIG5V.n1507 2.2505
R43254 ASIG5V.n1505 ASIG5V.n1470 2.2505
R43255 ASIG5V.n1503 ASIG5V.n1501 2.2505
R43256 ASIG5V.n1500 ASIG5V.n1472 2.2505
R43257 ASIG5V.n1499 ASIG5V.n1498 2.2505
R43258 ASIG5V.n1496 ASIG5V.n1473 2.2505
R43259 ASIG5V.n1494 ASIG5V.n1492 2.2505
R43260 ASIG5V.n1491 ASIG5V.n1475 2.2505
R43261 ASIG5V.n1490 ASIG5V.n1489 2.2505
R43262 ASIG5V.n1487 ASIG5V.n1476 2.2505
R43263 ASIG5V.n1485 ASIG5V.n1483 2.2505
R43264 ASIG5V.n1482 ASIG5V.n1478 2.2505
R43265 ASIG5V.n1481 ASIG5V.n1480 2.2505
R43266 ASIG5V.n1479 ASIG5V.n1372 2.2505
R43267 ASIG5V.n12009 ASIG5V.n1372 2.2505
R43268 ASIG5V.n1480 ASIG5V.n1371 2.2505
R43269 ASIG5V.n1478 ASIG5V.n1477 2.2505
R43270 ASIG5V.n1485 ASIG5V.n1484 2.2505
R43271 ASIG5V.n1487 ASIG5V.n1486 2.2505
R43272 ASIG5V.n1489 ASIG5V.n1488 2.2505
R43273 ASIG5V.n1475 ASIG5V.n1474 2.2505
R43274 ASIG5V.n1494 ASIG5V.n1493 2.2505
R43275 ASIG5V.n1496 ASIG5V.n1495 2.2505
R43276 ASIG5V.n1498 ASIG5V.n1497 2.2505
R43277 ASIG5V.n1472 ASIG5V.n1471 2.2505
R43278 ASIG5V.n1503 ASIG5V.n1502 2.2505
R43279 ASIG5V.n1505 ASIG5V.n1504 2.2505
R43280 ASIG5V.n1507 ASIG5V.n1506 2.2505
R43281 ASIG5V.n1469 ASIG5V.n1468 2.2505
R43282 ASIG5V.n1512 ASIG5V.n1511 2.2505
R43283 ASIG5V.n1514 ASIG5V.n1513 2.2505
R43284 ASIG5V.n1516 ASIG5V.n1515 2.2505
R43285 ASIG5V.n1466 ASIG5V.n1465 2.2505
R43286 ASIG5V.n1521 ASIG5V.n1520 2.2505
R43287 ASIG5V.n1523 ASIG5V.n1522 2.2505
R43288 ASIG5V.n1525 ASIG5V.n1524 2.2505
R43289 ASIG5V.n1463 ASIG5V.n1462 2.2505
R43290 ASIG5V.n1530 ASIG5V.n1529 2.2505
R43291 ASIG5V.n1532 ASIG5V.n1531 2.2505
R43292 ASIG5V.n1534 ASIG5V.n1533 2.2505
R43293 ASIG5V.n1460 ASIG5V.n1459 2.2505
R43294 ASIG5V.n1539 ASIG5V.n1538 2.2505
R43295 ASIG5V.n1541 ASIG5V.n1540 2.2505
R43296 ASIG5V.n1543 ASIG5V.n1542 2.2505
R43297 ASIG5V.n1457 ASIG5V.n1456 2.2505
R43298 ASIG5V.n1548 ASIG5V.n1547 2.2505
R43299 ASIG5V.n1550 ASIG5V.n1549 2.2505
R43300 ASIG5V.n1552 ASIG5V.n1551 2.2505
R43301 ASIG5V.n1454 ASIG5V.n1453 2.2505
R43302 ASIG5V.n1557 ASIG5V.n1556 2.2505
R43303 ASIG5V.n1559 ASIG5V.n1558 2.2505
R43304 ASIG5V.n1561 ASIG5V.n1560 2.2505
R43305 ASIG5V.n1451 ASIG5V.n1450 2.2505
R43306 ASIG5V.n1566 ASIG5V.n1565 2.2505
R43307 ASIG5V.n1568 ASIG5V.n1567 2.2505
R43308 ASIG5V.n1570 ASIG5V.n1569 2.2505
R43309 ASIG5V.n1448 ASIG5V.n1447 2.2505
R43310 ASIG5V.n1575 ASIG5V.n1574 2.2505
R43311 ASIG5V.n1577 ASIG5V.n1576 2.2505
R43312 ASIG5V.n1579 ASIG5V.n1578 2.2505
R43313 ASIG5V.n1445 ASIG5V.n1444 2.2505
R43314 ASIG5V.n1584 ASIG5V.n1583 2.2505
R43315 ASIG5V.n1586 ASIG5V.n1585 2.2505
R43316 ASIG5V.n1588 ASIG5V.n1587 2.2505
R43317 ASIG5V.n1442 ASIG5V.n1441 2.2505
R43318 ASIG5V.n1593 ASIG5V.n1592 2.2505
R43319 ASIG5V.n1595 ASIG5V.n1594 2.2505
R43320 ASIG5V.n1597 ASIG5V.n1596 2.2505
R43321 ASIG5V.n1439 ASIG5V.n1438 2.2505
R43322 ASIG5V.n1602 ASIG5V.n1601 2.2505
R43323 ASIG5V.n1604 ASIG5V.n1603 2.2505
R43324 ASIG5V.n1606 ASIG5V.n1605 2.2505
R43325 ASIG5V.n1436 ASIG5V.n1435 2.2505
R43326 ASIG5V.n1611 ASIG5V.n1610 2.2505
R43327 ASIG5V.n1613 ASIG5V.n1612 2.2505
R43328 ASIG5V.n1615 ASIG5V.n1614 2.2505
R43329 ASIG5V.n1433 ASIG5V.n1432 2.2505
R43330 ASIG5V.n1620 ASIG5V.n1619 2.2505
R43331 ASIG5V.n1622 ASIG5V.n1621 2.2505
R43332 ASIG5V.n1624 ASIG5V.n1623 2.2505
R43333 ASIG5V.n1430 ASIG5V.n1429 2.2505
R43334 ASIG5V.n1629 ASIG5V.n1628 2.2505
R43335 ASIG5V.n1631 ASIG5V.n1630 2.2505
R43336 ASIG5V.n1633 ASIG5V.n1632 2.2505
R43337 ASIG5V.n1427 ASIG5V.n1426 2.2505
R43338 ASIG5V.n1638 ASIG5V.n1637 2.2505
R43339 ASIG5V.n1640 ASIG5V.n1639 2.2505
R43340 ASIG5V.n1642 ASIG5V.n1641 2.2505
R43341 ASIG5V.n1424 ASIG5V.n1423 2.2505
R43342 ASIG5V.n1647 ASIG5V.n1646 2.2505
R43343 ASIG5V.n1649 ASIG5V.n1648 2.2505
R43344 ASIG5V.n1651 ASIG5V.n1650 2.2505
R43345 ASIG5V.n1421 ASIG5V.n1420 2.2505
R43346 ASIG5V.n1656 ASIG5V.n1655 2.2505
R43347 ASIG5V.n1658 ASIG5V.n1657 2.2505
R43348 ASIG5V.n1660 ASIG5V.n1659 2.2505
R43349 ASIG5V.n1418 ASIG5V.n1417 2.2505
R43350 ASIG5V.n12007 ASIG5V.n12006 2.2505
R43351 ASIG5V.n11992 ASIG5V.n11991 2.2505
R43352 ASIG5V.n11990 ASIG5V.n1765 2.2505
R43353 ASIG5V.n11989 ASIG5V.n11988 2.2505
R43354 ASIG5V.n11986 ASIG5V.n1766 2.2505
R43355 ASIG5V.n11984 ASIG5V.n11982 2.2505
R43356 ASIG5V.n11981 ASIG5V.n1768 2.2505
R43357 ASIG5V.n11980 ASIG5V.n11979 2.2505
R43358 ASIG5V.n11977 ASIG5V.n1769 2.2505
R43359 ASIG5V.n11975 ASIG5V.n11973 2.2505
R43360 ASIG5V.n11972 ASIG5V.n1771 2.2505
R43361 ASIG5V.n11971 ASIG5V.n11970 2.2505
R43362 ASIG5V.n11968 ASIG5V.n1772 2.2505
R43363 ASIG5V.n11966 ASIG5V.n11964 2.2505
R43364 ASIG5V.n11963 ASIG5V.n1774 2.2505
R43365 ASIG5V.n11962 ASIG5V.n11961 2.2505
R43366 ASIG5V.n11959 ASIG5V.n1775 2.2505
R43367 ASIG5V.n11957 ASIG5V.n11955 2.2505
R43368 ASIG5V.n11954 ASIG5V.n1777 2.2505
R43369 ASIG5V.n11953 ASIG5V.n11952 2.2505
R43370 ASIG5V.n11950 ASIG5V.n1778 2.2505
R43371 ASIG5V.n11948 ASIG5V.n11946 2.2505
R43372 ASIG5V.n11945 ASIG5V.n1780 2.2505
R43373 ASIG5V.n11944 ASIG5V.n11943 2.2505
R43374 ASIG5V.n11941 ASIG5V.n1781 2.2505
R43375 ASIG5V.n11939 ASIG5V.n11937 2.2505
R43376 ASIG5V.n11936 ASIG5V.n1783 2.2505
R43377 ASIG5V.n11935 ASIG5V.n11934 2.2505
R43378 ASIG5V.n11932 ASIG5V.n1784 2.2505
R43379 ASIG5V.n11930 ASIG5V.n11928 2.2505
R43380 ASIG5V.n11927 ASIG5V.n1786 2.2505
R43381 ASIG5V.n11926 ASIG5V.n11925 2.2505
R43382 ASIG5V.n11923 ASIG5V.n1787 2.2505
R43383 ASIG5V.n11921 ASIG5V.n11919 2.2505
R43384 ASIG5V.n11918 ASIG5V.n1789 2.2505
R43385 ASIG5V.n11917 ASIG5V.n11916 2.2505
R43386 ASIG5V.n11914 ASIG5V.n1790 2.2505
R43387 ASIG5V.n11912 ASIG5V.n11910 2.2505
R43388 ASIG5V.n11909 ASIG5V.n1792 2.2505
R43389 ASIG5V.n11908 ASIG5V.n11907 2.2505
R43390 ASIG5V.n11905 ASIG5V.n1793 2.2505
R43391 ASIG5V.n11903 ASIG5V.n11901 2.2505
R43392 ASIG5V.n11900 ASIG5V.n1795 2.2505
R43393 ASIG5V.n11899 ASIG5V.n11898 2.2505
R43394 ASIG5V.n11896 ASIG5V.n1796 2.2505
R43395 ASIG5V.n11894 ASIG5V.n11892 2.2505
R43396 ASIG5V.n11891 ASIG5V.n1798 2.2505
R43397 ASIG5V.n11890 ASIG5V.n11889 2.2505
R43398 ASIG5V.n11887 ASIG5V.n1799 2.2505
R43399 ASIG5V.n11885 ASIG5V.n11883 2.2505
R43400 ASIG5V.n11882 ASIG5V.n1801 2.2505
R43401 ASIG5V.n11881 ASIG5V.n11880 2.2505
R43402 ASIG5V.n11878 ASIG5V.n1802 2.2505
R43403 ASIG5V.n11876 ASIG5V.n11874 2.2505
R43404 ASIG5V.n11873 ASIG5V.n1804 2.2505
R43405 ASIG5V.n11872 ASIG5V.n11871 2.2505
R43406 ASIG5V.n11869 ASIG5V.n1805 2.2505
R43407 ASIG5V.n11867 ASIG5V.n11865 2.2505
R43408 ASIG5V.n11864 ASIG5V.n1807 2.2505
R43409 ASIG5V.n11863 ASIG5V.n11862 2.2505
R43410 ASIG5V.n11860 ASIG5V.n1808 2.2505
R43411 ASIG5V.n11858 ASIG5V.n11856 2.2505
R43412 ASIG5V.n11855 ASIG5V.n1810 2.2505
R43413 ASIG5V.n11854 ASIG5V.n11853 2.2505
R43414 ASIG5V.n11851 ASIG5V.n1811 2.2505
R43415 ASIG5V.n11849 ASIG5V.n11847 2.2505
R43416 ASIG5V.n11846 ASIG5V.n1813 2.2505
R43417 ASIG5V.n11845 ASIG5V.n11844 2.2505
R43418 ASIG5V.n11842 ASIG5V.n1814 2.2505
R43419 ASIG5V.n11840 ASIG5V.n11838 2.2505
R43420 ASIG5V.n11837 ASIG5V.n1816 2.2505
R43421 ASIG5V.n11836 ASIG5V.n11835 2.2505
R43422 ASIG5V.n11833 ASIG5V.n1817 2.2505
R43423 ASIG5V.n11831 ASIG5V.n11829 2.2505
R43424 ASIG5V.n11828 ASIG5V.n1819 2.2505
R43425 ASIG5V.n11827 ASIG5V.n11826 2.2505
R43426 ASIG5V.n11824 ASIG5V.n1820 2.2505
R43427 ASIG5V.n11822 ASIG5V.n11820 2.2505
R43428 ASIG5V.n11819 ASIG5V.n1822 2.2505
R43429 ASIG5V.n11818 ASIG5V.n11817 2.2505
R43430 ASIG5V.n11815 ASIG5V.n1823 2.2505
R43431 ASIG5V.n11813 ASIG5V.n11811 2.2505
R43432 ASIG5V.n11810 ASIG5V.n1825 2.2505
R43433 ASIG5V.n11809 ASIG5V.n11808 2.2505
R43434 ASIG5V.n11807 ASIG5V.n1720 2.2505
R43435 ASIG5V.n11995 ASIG5V.n1720 2.2505
R43436 ASIG5V.n11808 ASIG5V.n1718 2.2505
R43437 ASIG5V.n1825 ASIG5V.n1824 2.2505
R43438 ASIG5V.n11813 ASIG5V.n11812 2.2505
R43439 ASIG5V.n11815 ASIG5V.n11814 2.2505
R43440 ASIG5V.n11817 ASIG5V.n11816 2.2505
R43441 ASIG5V.n1822 ASIG5V.n1821 2.2505
R43442 ASIG5V.n11822 ASIG5V.n11821 2.2505
R43443 ASIG5V.n11824 ASIG5V.n11823 2.2505
R43444 ASIG5V.n11826 ASIG5V.n11825 2.2505
R43445 ASIG5V.n1819 ASIG5V.n1818 2.2505
R43446 ASIG5V.n11831 ASIG5V.n11830 2.2505
R43447 ASIG5V.n11833 ASIG5V.n11832 2.2505
R43448 ASIG5V.n11835 ASIG5V.n11834 2.2505
R43449 ASIG5V.n1816 ASIG5V.n1815 2.2505
R43450 ASIG5V.n11840 ASIG5V.n11839 2.2505
R43451 ASIG5V.n11842 ASIG5V.n11841 2.2505
R43452 ASIG5V.n11844 ASIG5V.n11843 2.2505
R43453 ASIG5V.n1813 ASIG5V.n1812 2.2505
R43454 ASIG5V.n11849 ASIG5V.n11848 2.2505
R43455 ASIG5V.n11851 ASIG5V.n11850 2.2505
R43456 ASIG5V.n11853 ASIG5V.n11852 2.2505
R43457 ASIG5V.n1810 ASIG5V.n1809 2.2505
R43458 ASIG5V.n11858 ASIG5V.n11857 2.2505
R43459 ASIG5V.n11860 ASIG5V.n11859 2.2505
R43460 ASIG5V.n11862 ASIG5V.n11861 2.2505
R43461 ASIG5V.n1807 ASIG5V.n1806 2.2505
R43462 ASIG5V.n11867 ASIG5V.n11866 2.2505
R43463 ASIG5V.n11869 ASIG5V.n11868 2.2505
R43464 ASIG5V.n11871 ASIG5V.n11870 2.2505
R43465 ASIG5V.n1804 ASIG5V.n1803 2.2505
R43466 ASIG5V.n11876 ASIG5V.n11875 2.2505
R43467 ASIG5V.n11878 ASIG5V.n11877 2.2505
R43468 ASIG5V.n11880 ASIG5V.n11879 2.2505
R43469 ASIG5V.n1801 ASIG5V.n1800 2.2505
R43470 ASIG5V.n11885 ASIG5V.n11884 2.2505
R43471 ASIG5V.n11887 ASIG5V.n11886 2.2505
R43472 ASIG5V.n11889 ASIG5V.n11888 2.2505
R43473 ASIG5V.n1798 ASIG5V.n1797 2.2505
R43474 ASIG5V.n11894 ASIG5V.n11893 2.2505
R43475 ASIG5V.n11896 ASIG5V.n11895 2.2505
R43476 ASIG5V.n11898 ASIG5V.n11897 2.2505
R43477 ASIG5V.n1795 ASIG5V.n1794 2.2505
R43478 ASIG5V.n11903 ASIG5V.n11902 2.2505
R43479 ASIG5V.n11905 ASIG5V.n11904 2.2505
R43480 ASIG5V.n11907 ASIG5V.n11906 2.2505
R43481 ASIG5V.n1792 ASIG5V.n1791 2.2505
R43482 ASIG5V.n11912 ASIG5V.n11911 2.2505
R43483 ASIG5V.n11914 ASIG5V.n11913 2.2505
R43484 ASIG5V.n11916 ASIG5V.n11915 2.2505
R43485 ASIG5V.n1789 ASIG5V.n1788 2.2505
R43486 ASIG5V.n11921 ASIG5V.n11920 2.2505
R43487 ASIG5V.n11923 ASIG5V.n11922 2.2505
R43488 ASIG5V.n11925 ASIG5V.n11924 2.2505
R43489 ASIG5V.n1786 ASIG5V.n1785 2.2505
R43490 ASIG5V.n11930 ASIG5V.n11929 2.2505
R43491 ASIG5V.n11932 ASIG5V.n11931 2.2505
R43492 ASIG5V.n11934 ASIG5V.n11933 2.2505
R43493 ASIG5V.n1783 ASIG5V.n1782 2.2505
R43494 ASIG5V.n11939 ASIG5V.n11938 2.2505
R43495 ASIG5V.n11941 ASIG5V.n11940 2.2505
R43496 ASIG5V.n11943 ASIG5V.n11942 2.2505
R43497 ASIG5V.n1780 ASIG5V.n1779 2.2505
R43498 ASIG5V.n11948 ASIG5V.n11947 2.2505
R43499 ASIG5V.n11950 ASIG5V.n11949 2.2505
R43500 ASIG5V.n11952 ASIG5V.n11951 2.2505
R43501 ASIG5V.n1777 ASIG5V.n1776 2.2505
R43502 ASIG5V.n11957 ASIG5V.n11956 2.2505
R43503 ASIG5V.n11959 ASIG5V.n11958 2.2505
R43504 ASIG5V.n11961 ASIG5V.n11960 2.2505
R43505 ASIG5V.n1774 ASIG5V.n1773 2.2505
R43506 ASIG5V.n11966 ASIG5V.n11965 2.2505
R43507 ASIG5V.n11968 ASIG5V.n11967 2.2505
R43508 ASIG5V.n11970 ASIG5V.n11969 2.2505
R43509 ASIG5V.n1771 ASIG5V.n1770 2.2505
R43510 ASIG5V.n11975 ASIG5V.n11974 2.2505
R43511 ASIG5V.n11977 ASIG5V.n11976 2.2505
R43512 ASIG5V.n11979 ASIG5V.n11978 2.2505
R43513 ASIG5V.n1768 ASIG5V.n1767 2.2505
R43514 ASIG5V.n11984 ASIG5V.n11983 2.2505
R43515 ASIG5V.n11986 ASIG5V.n11985 2.2505
R43516 ASIG5V.n11988 ASIG5V.n11987 2.2505
R43517 ASIG5V.n1765 ASIG5V.n1764 2.2505
R43518 ASIG5V.n11993 ASIG5V.n11992 2.2505
R43519 ASIG5V.n1907 ASIG5V.n1854 2.2505
R43520 ASIG5V.n2194 ASIG5V.n2193 2.2505
R43521 ASIG5V.n2192 ASIG5V.n1908 2.2505
R43522 ASIG5V.n2191 ASIG5V.n2190 2.2505
R43523 ASIG5V.n2186 ASIG5V.n1909 2.2505
R43524 ASIG5V.n2182 ASIG5V.n2181 2.2505
R43525 ASIG5V.n2180 ASIG5V.n1910 2.2505
R43526 ASIG5V.n2179 ASIG5V.n2178 2.2505
R43527 ASIG5V.n2174 ASIG5V.n1911 2.2505
R43528 ASIG5V.n2170 ASIG5V.n2169 2.2505
R43529 ASIG5V.n2168 ASIG5V.n1912 2.2505
R43530 ASIG5V.n2167 ASIG5V.n2166 2.2505
R43531 ASIG5V.n2162 ASIG5V.n1913 2.2505
R43532 ASIG5V.n2158 ASIG5V.n2157 2.2505
R43533 ASIG5V.n2156 ASIG5V.n1914 2.2505
R43534 ASIG5V.n2155 ASIG5V.n2154 2.2505
R43535 ASIG5V.n2150 ASIG5V.n1915 2.2505
R43536 ASIG5V.n2146 ASIG5V.n2145 2.2505
R43537 ASIG5V.n2144 ASIG5V.n1916 2.2505
R43538 ASIG5V.n2143 ASIG5V.n2142 2.2505
R43539 ASIG5V.n2138 ASIG5V.n1917 2.2505
R43540 ASIG5V.n2134 ASIG5V.n2133 2.2505
R43541 ASIG5V.n2132 ASIG5V.n1918 2.2505
R43542 ASIG5V.n2131 ASIG5V.n2130 2.2505
R43543 ASIG5V.n2126 ASIG5V.n1919 2.2505
R43544 ASIG5V.n2122 ASIG5V.n2121 2.2505
R43545 ASIG5V.n2120 ASIG5V.n1920 2.2505
R43546 ASIG5V.n2119 ASIG5V.n2118 2.2505
R43547 ASIG5V.n2114 ASIG5V.n1921 2.2505
R43548 ASIG5V.n2110 ASIG5V.n2109 2.2505
R43549 ASIG5V.n2108 ASIG5V.n1922 2.2505
R43550 ASIG5V.n2107 ASIG5V.n2106 2.2505
R43551 ASIG5V.n2102 ASIG5V.n1923 2.2505
R43552 ASIG5V.n2098 ASIG5V.n2097 2.2505
R43553 ASIG5V.n2096 ASIG5V.n1924 2.2505
R43554 ASIG5V.n2095 ASIG5V.n2094 2.2505
R43555 ASIG5V.n2090 ASIG5V.n1925 2.2505
R43556 ASIG5V.n2086 ASIG5V.n2085 2.2505
R43557 ASIG5V.n2084 ASIG5V.n1926 2.2505
R43558 ASIG5V.n2083 ASIG5V.n2082 2.2505
R43559 ASIG5V.n2078 ASIG5V.n1927 2.2505
R43560 ASIG5V.n2074 ASIG5V.n2073 2.2505
R43561 ASIG5V.n2072 ASIG5V.n1928 2.2505
R43562 ASIG5V.n2071 ASIG5V.n2070 2.2505
R43563 ASIG5V.n2066 ASIG5V.n1929 2.2505
R43564 ASIG5V.n2062 ASIG5V.n2061 2.2505
R43565 ASIG5V.n2060 ASIG5V.n1930 2.2505
R43566 ASIG5V.n2059 ASIG5V.n2058 2.2505
R43567 ASIG5V.n2054 ASIG5V.n1931 2.2505
R43568 ASIG5V.n2050 ASIG5V.n2049 2.2505
R43569 ASIG5V.n2048 ASIG5V.n1932 2.2505
R43570 ASIG5V.n2047 ASIG5V.n2046 2.2505
R43571 ASIG5V.n2042 ASIG5V.n1933 2.2505
R43572 ASIG5V.n2038 ASIG5V.n2037 2.2505
R43573 ASIG5V.n2036 ASIG5V.n1934 2.2505
R43574 ASIG5V.n2035 ASIG5V.n2034 2.2505
R43575 ASIG5V.n2030 ASIG5V.n1935 2.2505
R43576 ASIG5V.n2026 ASIG5V.n2025 2.2505
R43577 ASIG5V.n2024 ASIG5V.n1936 2.2505
R43578 ASIG5V.n2023 ASIG5V.n2022 2.2505
R43579 ASIG5V.n2018 ASIG5V.n1937 2.2505
R43580 ASIG5V.n2014 ASIG5V.n2013 2.2505
R43581 ASIG5V.n2012 ASIG5V.n1938 2.2505
R43582 ASIG5V.n2011 ASIG5V.n2010 2.2505
R43583 ASIG5V.n2006 ASIG5V.n1939 2.2505
R43584 ASIG5V.n2002 ASIG5V.n2001 2.2505
R43585 ASIG5V.n2000 ASIG5V.n1940 2.2505
R43586 ASIG5V.n1999 ASIG5V.n1998 2.2505
R43587 ASIG5V.n1994 ASIG5V.n1941 2.2505
R43588 ASIG5V.n1990 ASIG5V.n1989 2.2505
R43589 ASIG5V.n1988 ASIG5V.n1942 2.2505
R43590 ASIG5V.n1987 ASIG5V.n1986 2.2505
R43591 ASIG5V.n1982 ASIG5V.n1943 2.2505
R43592 ASIG5V.n1978 ASIG5V.n1977 2.2505
R43593 ASIG5V.n1976 ASIG5V.n1944 2.2505
R43594 ASIG5V.n1975 ASIG5V.n1974 2.2505
R43595 ASIG5V.n1970 ASIG5V.n1945 2.2505
R43596 ASIG5V.n1966 ASIG5V.n1965 2.2505
R43597 ASIG5V.n1964 ASIG5V.n1946 2.2505
R43598 ASIG5V.n1963 ASIG5V.n1962 2.2505
R43599 ASIG5V.n1958 ASIG5V.n1947 2.2505
R43600 ASIG5V.n1954 ASIG5V.n1953 2.2505
R43601 ASIG5V.n1952 ASIG5V.n1951 2.2505
R43602 ASIG5V.n1948 ASIG5V.n1842 2.2505
R43603 ASIG5V.n1948 ASIG5V.n1906 2.2505
R43604 ASIG5V.n1951 ASIG5V.n1950 2.2505
R43605 ASIG5V.n1955 ASIG5V.n1954 2.2505
R43606 ASIG5V.n1958 ASIG5V.n1957 2.2505
R43607 ASIG5V.n1962 ASIG5V.n1961 2.2505
R43608 ASIG5V.n1959 ASIG5V.n1946 2.2505
R43609 ASIG5V.n1967 ASIG5V.n1966 2.2505
R43610 ASIG5V.n1970 ASIG5V.n1969 2.2505
R43611 ASIG5V.n1974 ASIG5V.n1973 2.2505
R43612 ASIG5V.n1971 ASIG5V.n1944 2.2505
R43613 ASIG5V.n1979 ASIG5V.n1978 2.2505
R43614 ASIG5V.n1982 ASIG5V.n1981 2.2505
R43615 ASIG5V.n1986 ASIG5V.n1985 2.2505
R43616 ASIG5V.n1983 ASIG5V.n1942 2.2505
R43617 ASIG5V.n1991 ASIG5V.n1990 2.2505
R43618 ASIG5V.n1994 ASIG5V.n1993 2.2505
R43619 ASIG5V.n1998 ASIG5V.n1997 2.2505
R43620 ASIG5V.n1995 ASIG5V.n1940 2.2505
R43621 ASIG5V.n2003 ASIG5V.n2002 2.2505
R43622 ASIG5V.n2006 ASIG5V.n2005 2.2505
R43623 ASIG5V.n2010 ASIG5V.n2009 2.2505
R43624 ASIG5V.n2007 ASIG5V.n1938 2.2505
R43625 ASIG5V.n2015 ASIG5V.n2014 2.2505
R43626 ASIG5V.n2018 ASIG5V.n2017 2.2505
R43627 ASIG5V.n2022 ASIG5V.n2021 2.2505
R43628 ASIG5V.n2019 ASIG5V.n1936 2.2505
R43629 ASIG5V.n2027 ASIG5V.n2026 2.2505
R43630 ASIG5V.n2030 ASIG5V.n2029 2.2505
R43631 ASIG5V.n2034 ASIG5V.n2033 2.2505
R43632 ASIG5V.n2031 ASIG5V.n1934 2.2505
R43633 ASIG5V.n2039 ASIG5V.n2038 2.2505
R43634 ASIG5V.n2042 ASIG5V.n2041 2.2505
R43635 ASIG5V.n2046 ASIG5V.n2045 2.2505
R43636 ASIG5V.n2043 ASIG5V.n1932 2.2505
R43637 ASIG5V.n2051 ASIG5V.n2050 2.2505
R43638 ASIG5V.n2054 ASIG5V.n2053 2.2505
R43639 ASIG5V.n2058 ASIG5V.n2057 2.2505
R43640 ASIG5V.n2055 ASIG5V.n1930 2.2505
R43641 ASIG5V.n2063 ASIG5V.n2062 2.2505
R43642 ASIG5V.n2066 ASIG5V.n2065 2.2505
R43643 ASIG5V.n2070 ASIG5V.n2069 2.2505
R43644 ASIG5V.n2067 ASIG5V.n1928 2.2505
R43645 ASIG5V.n2075 ASIG5V.n2074 2.2505
R43646 ASIG5V.n2078 ASIG5V.n2077 2.2505
R43647 ASIG5V.n2082 ASIG5V.n2081 2.2505
R43648 ASIG5V.n2079 ASIG5V.n1926 2.2505
R43649 ASIG5V.n2087 ASIG5V.n2086 2.2505
R43650 ASIG5V.n2090 ASIG5V.n2089 2.2505
R43651 ASIG5V.n2094 ASIG5V.n2093 2.2505
R43652 ASIG5V.n2091 ASIG5V.n1924 2.2505
R43653 ASIG5V.n2099 ASIG5V.n2098 2.2505
R43654 ASIG5V.n2102 ASIG5V.n2101 2.2505
R43655 ASIG5V.n2106 ASIG5V.n2105 2.2505
R43656 ASIG5V.n2103 ASIG5V.n1922 2.2505
R43657 ASIG5V.n2111 ASIG5V.n2110 2.2505
R43658 ASIG5V.n2114 ASIG5V.n2113 2.2505
R43659 ASIG5V.n2118 ASIG5V.n2117 2.2505
R43660 ASIG5V.n2115 ASIG5V.n1920 2.2505
R43661 ASIG5V.n2123 ASIG5V.n2122 2.2505
R43662 ASIG5V.n2126 ASIG5V.n2125 2.2505
R43663 ASIG5V.n2130 ASIG5V.n2129 2.2505
R43664 ASIG5V.n2127 ASIG5V.n1918 2.2505
R43665 ASIG5V.n2135 ASIG5V.n2134 2.2505
R43666 ASIG5V.n2138 ASIG5V.n2137 2.2505
R43667 ASIG5V.n2142 ASIG5V.n2141 2.2505
R43668 ASIG5V.n2139 ASIG5V.n1916 2.2505
R43669 ASIG5V.n2147 ASIG5V.n2146 2.2505
R43670 ASIG5V.n2150 ASIG5V.n2149 2.2505
R43671 ASIG5V.n2154 ASIG5V.n2153 2.2505
R43672 ASIG5V.n2151 ASIG5V.n1914 2.2505
R43673 ASIG5V.n2159 ASIG5V.n2158 2.2505
R43674 ASIG5V.n2162 ASIG5V.n2161 2.2505
R43675 ASIG5V.n2166 ASIG5V.n2165 2.2505
R43676 ASIG5V.n2163 ASIG5V.n1912 2.2505
R43677 ASIG5V.n2171 ASIG5V.n2170 2.2505
R43678 ASIG5V.n2174 ASIG5V.n2173 2.2505
R43679 ASIG5V.n2178 ASIG5V.n2177 2.2505
R43680 ASIG5V.n2175 ASIG5V.n1910 2.2505
R43681 ASIG5V.n2183 ASIG5V.n2182 2.2505
R43682 ASIG5V.n2186 ASIG5V.n2185 2.2505
R43683 ASIG5V.n2190 ASIG5V.n2189 2.2505
R43684 ASIG5V.n2187 ASIG5V.n1908 2.2505
R43685 ASIG5V.n2195 ASIG5V.n2194 2.2505
R43686 ASIG5V.n2197 ASIG5V.n1907 2.2505
R43687 ASIG5V.n2264 ASIG5V.n2206 2.2505
R43688 ASIG5V.n2551 ASIG5V.n2550 2.2505
R43689 ASIG5V.n2549 ASIG5V.n2265 2.2505
R43690 ASIG5V.n2548 ASIG5V.n2547 2.2505
R43691 ASIG5V.n2543 ASIG5V.n2266 2.2505
R43692 ASIG5V.n2539 ASIG5V.n2538 2.2505
R43693 ASIG5V.n2537 ASIG5V.n2267 2.2505
R43694 ASIG5V.n2536 ASIG5V.n2535 2.2505
R43695 ASIG5V.n2531 ASIG5V.n2268 2.2505
R43696 ASIG5V.n2527 ASIG5V.n2526 2.2505
R43697 ASIG5V.n2525 ASIG5V.n2269 2.2505
R43698 ASIG5V.n2524 ASIG5V.n2523 2.2505
R43699 ASIG5V.n2519 ASIG5V.n2270 2.2505
R43700 ASIG5V.n2515 ASIG5V.n2514 2.2505
R43701 ASIG5V.n2513 ASIG5V.n2271 2.2505
R43702 ASIG5V.n2512 ASIG5V.n2511 2.2505
R43703 ASIG5V.n2507 ASIG5V.n2272 2.2505
R43704 ASIG5V.n2503 ASIG5V.n2502 2.2505
R43705 ASIG5V.n2501 ASIG5V.n2273 2.2505
R43706 ASIG5V.n2500 ASIG5V.n2499 2.2505
R43707 ASIG5V.n2495 ASIG5V.n2274 2.2505
R43708 ASIG5V.n2491 ASIG5V.n2490 2.2505
R43709 ASIG5V.n2489 ASIG5V.n2275 2.2505
R43710 ASIG5V.n2488 ASIG5V.n2487 2.2505
R43711 ASIG5V.n2483 ASIG5V.n2276 2.2505
R43712 ASIG5V.n2479 ASIG5V.n2478 2.2505
R43713 ASIG5V.n2477 ASIG5V.n2277 2.2505
R43714 ASIG5V.n2476 ASIG5V.n2475 2.2505
R43715 ASIG5V.n2471 ASIG5V.n2278 2.2505
R43716 ASIG5V.n2467 ASIG5V.n2466 2.2505
R43717 ASIG5V.n2465 ASIG5V.n2279 2.2505
R43718 ASIG5V.n2464 ASIG5V.n2463 2.2505
R43719 ASIG5V.n2459 ASIG5V.n2280 2.2505
R43720 ASIG5V.n2455 ASIG5V.n2454 2.2505
R43721 ASIG5V.n2453 ASIG5V.n2281 2.2505
R43722 ASIG5V.n2452 ASIG5V.n2451 2.2505
R43723 ASIG5V.n2447 ASIG5V.n2282 2.2505
R43724 ASIG5V.n2443 ASIG5V.n2442 2.2505
R43725 ASIG5V.n2441 ASIG5V.n2283 2.2505
R43726 ASIG5V.n2440 ASIG5V.n2439 2.2505
R43727 ASIG5V.n2435 ASIG5V.n2284 2.2505
R43728 ASIG5V.n2431 ASIG5V.n2430 2.2505
R43729 ASIG5V.n2429 ASIG5V.n2285 2.2505
R43730 ASIG5V.n2428 ASIG5V.n2427 2.2505
R43731 ASIG5V.n2423 ASIG5V.n2286 2.2505
R43732 ASIG5V.n2419 ASIG5V.n2418 2.2505
R43733 ASIG5V.n2417 ASIG5V.n2287 2.2505
R43734 ASIG5V.n2416 ASIG5V.n2415 2.2505
R43735 ASIG5V.n2411 ASIG5V.n2288 2.2505
R43736 ASIG5V.n2407 ASIG5V.n2406 2.2505
R43737 ASIG5V.n2405 ASIG5V.n2289 2.2505
R43738 ASIG5V.n2404 ASIG5V.n2403 2.2505
R43739 ASIG5V.n2399 ASIG5V.n2290 2.2505
R43740 ASIG5V.n2395 ASIG5V.n2394 2.2505
R43741 ASIG5V.n2393 ASIG5V.n2291 2.2505
R43742 ASIG5V.n2392 ASIG5V.n2391 2.2505
R43743 ASIG5V.n2387 ASIG5V.n2292 2.2505
R43744 ASIG5V.n2383 ASIG5V.n2382 2.2505
R43745 ASIG5V.n2381 ASIG5V.n2293 2.2505
R43746 ASIG5V.n2380 ASIG5V.n2379 2.2505
R43747 ASIG5V.n2375 ASIG5V.n2294 2.2505
R43748 ASIG5V.n2371 ASIG5V.n2370 2.2505
R43749 ASIG5V.n2369 ASIG5V.n2295 2.2505
R43750 ASIG5V.n2368 ASIG5V.n2367 2.2505
R43751 ASIG5V.n2363 ASIG5V.n2296 2.2505
R43752 ASIG5V.n2359 ASIG5V.n2358 2.2505
R43753 ASIG5V.n2357 ASIG5V.n2297 2.2505
R43754 ASIG5V.n2356 ASIG5V.n2355 2.2505
R43755 ASIG5V.n2351 ASIG5V.n2298 2.2505
R43756 ASIG5V.n2347 ASIG5V.n2346 2.2505
R43757 ASIG5V.n2345 ASIG5V.n2299 2.2505
R43758 ASIG5V.n2344 ASIG5V.n2343 2.2505
R43759 ASIG5V.n2339 ASIG5V.n2300 2.2505
R43760 ASIG5V.n2335 ASIG5V.n2334 2.2505
R43761 ASIG5V.n2333 ASIG5V.n2301 2.2505
R43762 ASIG5V.n2332 ASIG5V.n2331 2.2505
R43763 ASIG5V.n2327 ASIG5V.n2302 2.2505
R43764 ASIG5V.n2323 ASIG5V.n2322 2.2505
R43765 ASIG5V.n2321 ASIG5V.n2303 2.2505
R43766 ASIG5V.n2320 ASIG5V.n2319 2.2505
R43767 ASIG5V.n2315 ASIG5V.n2304 2.2505
R43768 ASIG5V.n2311 ASIG5V.n2310 2.2505
R43769 ASIG5V.n2309 ASIG5V.n2308 2.2505
R43770 ASIG5V.n2305 ASIG5V.n2218 2.2505
R43771 ASIG5V.n2305 ASIG5V.n2263 2.2505
R43772 ASIG5V.n2308 ASIG5V.n2307 2.2505
R43773 ASIG5V.n2312 ASIG5V.n2311 2.2505
R43774 ASIG5V.n2315 ASIG5V.n2314 2.2505
R43775 ASIG5V.n2319 ASIG5V.n2318 2.2505
R43776 ASIG5V.n2316 ASIG5V.n2303 2.2505
R43777 ASIG5V.n2324 ASIG5V.n2323 2.2505
R43778 ASIG5V.n2327 ASIG5V.n2326 2.2505
R43779 ASIG5V.n2331 ASIG5V.n2330 2.2505
R43780 ASIG5V.n2328 ASIG5V.n2301 2.2505
R43781 ASIG5V.n2336 ASIG5V.n2335 2.2505
R43782 ASIG5V.n2339 ASIG5V.n2338 2.2505
R43783 ASIG5V.n2343 ASIG5V.n2342 2.2505
R43784 ASIG5V.n2340 ASIG5V.n2299 2.2505
R43785 ASIG5V.n2348 ASIG5V.n2347 2.2505
R43786 ASIG5V.n2351 ASIG5V.n2350 2.2505
R43787 ASIG5V.n2355 ASIG5V.n2354 2.2505
R43788 ASIG5V.n2352 ASIG5V.n2297 2.2505
R43789 ASIG5V.n2360 ASIG5V.n2359 2.2505
R43790 ASIG5V.n2363 ASIG5V.n2362 2.2505
R43791 ASIG5V.n2367 ASIG5V.n2366 2.2505
R43792 ASIG5V.n2364 ASIG5V.n2295 2.2505
R43793 ASIG5V.n2372 ASIG5V.n2371 2.2505
R43794 ASIG5V.n2375 ASIG5V.n2374 2.2505
R43795 ASIG5V.n2379 ASIG5V.n2378 2.2505
R43796 ASIG5V.n2376 ASIG5V.n2293 2.2505
R43797 ASIG5V.n2384 ASIG5V.n2383 2.2505
R43798 ASIG5V.n2387 ASIG5V.n2386 2.2505
R43799 ASIG5V.n2391 ASIG5V.n2390 2.2505
R43800 ASIG5V.n2388 ASIG5V.n2291 2.2505
R43801 ASIG5V.n2396 ASIG5V.n2395 2.2505
R43802 ASIG5V.n2399 ASIG5V.n2398 2.2505
R43803 ASIG5V.n2403 ASIG5V.n2402 2.2505
R43804 ASIG5V.n2400 ASIG5V.n2289 2.2505
R43805 ASIG5V.n2408 ASIG5V.n2407 2.2505
R43806 ASIG5V.n2411 ASIG5V.n2410 2.2505
R43807 ASIG5V.n2415 ASIG5V.n2414 2.2505
R43808 ASIG5V.n2412 ASIG5V.n2287 2.2505
R43809 ASIG5V.n2420 ASIG5V.n2419 2.2505
R43810 ASIG5V.n2423 ASIG5V.n2422 2.2505
R43811 ASIG5V.n2427 ASIG5V.n2426 2.2505
R43812 ASIG5V.n2424 ASIG5V.n2285 2.2505
R43813 ASIG5V.n2432 ASIG5V.n2431 2.2505
R43814 ASIG5V.n2435 ASIG5V.n2434 2.2505
R43815 ASIG5V.n2439 ASIG5V.n2438 2.2505
R43816 ASIG5V.n2436 ASIG5V.n2283 2.2505
R43817 ASIG5V.n2444 ASIG5V.n2443 2.2505
R43818 ASIG5V.n2447 ASIG5V.n2446 2.2505
R43819 ASIG5V.n2451 ASIG5V.n2450 2.2505
R43820 ASIG5V.n2448 ASIG5V.n2281 2.2505
R43821 ASIG5V.n2456 ASIG5V.n2455 2.2505
R43822 ASIG5V.n2459 ASIG5V.n2458 2.2505
R43823 ASIG5V.n2463 ASIG5V.n2462 2.2505
R43824 ASIG5V.n2460 ASIG5V.n2279 2.2505
R43825 ASIG5V.n2468 ASIG5V.n2467 2.2505
R43826 ASIG5V.n2471 ASIG5V.n2470 2.2505
R43827 ASIG5V.n2475 ASIG5V.n2474 2.2505
R43828 ASIG5V.n2472 ASIG5V.n2277 2.2505
R43829 ASIG5V.n2480 ASIG5V.n2479 2.2505
R43830 ASIG5V.n2483 ASIG5V.n2482 2.2505
R43831 ASIG5V.n2487 ASIG5V.n2486 2.2505
R43832 ASIG5V.n2484 ASIG5V.n2275 2.2505
R43833 ASIG5V.n2492 ASIG5V.n2491 2.2505
R43834 ASIG5V.n2495 ASIG5V.n2494 2.2505
R43835 ASIG5V.n2499 ASIG5V.n2498 2.2505
R43836 ASIG5V.n2496 ASIG5V.n2273 2.2505
R43837 ASIG5V.n2504 ASIG5V.n2503 2.2505
R43838 ASIG5V.n2507 ASIG5V.n2506 2.2505
R43839 ASIG5V.n2511 ASIG5V.n2510 2.2505
R43840 ASIG5V.n2508 ASIG5V.n2271 2.2505
R43841 ASIG5V.n2516 ASIG5V.n2515 2.2505
R43842 ASIG5V.n2519 ASIG5V.n2518 2.2505
R43843 ASIG5V.n2523 ASIG5V.n2522 2.2505
R43844 ASIG5V.n2520 ASIG5V.n2269 2.2505
R43845 ASIG5V.n2528 ASIG5V.n2527 2.2505
R43846 ASIG5V.n2531 ASIG5V.n2530 2.2505
R43847 ASIG5V.n2535 ASIG5V.n2534 2.2505
R43848 ASIG5V.n2532 ASIG5V.n2267 2.2505
R43849 ASIG5V.n2540 ASIG5V.n2539 2.2505
R43850 ASIG5V.n2543 ASIG5V.n2542 2.2505
R43851 ASIG5V.n2547 ASIG5V.n2546 2.2505
R43852 ASIG5V.n2544 ASIG5V.n2265 2.2505
R43853 ASIG5V.n2552 ASIG5V.n2551 2.2505
R43854 ASIG5V.n2554 ASIG5V.n2264 2.2505
R43855 ASIG5V.n11765 ASIG5V.n2614 2.2505
R43856 ASIG5V.n11767 ASIG5V.n11766 2.2505
R43857 ASIG5V.n2901 ASIG5V.n2617 2.2505
R43858 ASIG5V.n2900 ASIG5V.n2899 2.2505
R43859 ASIG5V.n2895 ASIG5V.n2618 2.2505
R43860 ASIG5V.n2891 ASIG5V.n2890 2.2505
R43861 ASIG5V.n2889 ASIG5V.n2619 2.2505
R43862 ASIG5V.n2888 ASIG5V.n2887 2.2505
R43863 ASIG5V.n2883 ASIG5V.n2620 2.2505
R43864 ASIG5V.n2879 ASIG5V.n2878 2.2505
R43865 ASIG5V.n2877 ASIG5V.n2621 2.2505
R43866 ASIG5V.n2876 ASIG5V.n2875 2.2505
R43867 ASIG5V.n2871 ASIG5V.n2622 2.2505
R43868 ASIG5V.n2867 ASIG5V.n2866 2.2505
R43869 ASIG5V.n2865 ASIG5V.n2623 2.2505
R43870 ASIG5V.n2864 ASIG5V.n2863 2.2505
R43871 ASIG5V.n2859 ASIG5V.n2624 2.2505
R43872 ASIG5V.n2855 ASIG5V.n2854 2.2505
R43873 ASIG5V.n2853 ASIG5V.n2625 2.2505
R43874 ASIG5V.n2852 ASIG5V.n2851 2.2505
R43875 ASIG5V.n2847 ASIG5V.n2626 2.2505
R43876 ASIG5V.n2843 ASIG5V.n2842 2.2505
R43877 ASIG5V.n2841 ASIG5V.n2627 2.2505
R43878 ASIG5V.n2840 ASIG5V.n2839 2.2505
R43879 ASIG5V.n2835 ASIG5V.n2628 2.2505
R43880 ASIG5V.n2831 ASIG5V.n2830 2.2505
R43881 ASIG5V.n2829 ASIG5V.n2629 2.2505
R43882 ASIG5V.n2828 ASIG5V.n2827 2.2505
R43883 ASIG5V.n2823 ASIG5V.n2630 2.2505
R43884 ASIG5V.n2819 ASIG5V.n2818 2.2505
R43885 ASIG5V.n2817 ASIG5V.n2631 2.2505
R43886 ASIG5V.n2816 ASIG5V.n2815 2.2505
R43887 ASIG5V.n2811 ASIG5V.n2632 2.2505
R43888 ASIG5V.n2807 ASIG5V.n2806 2.2505
R43889 ASIG5V.n2805 ASIG5V.n2633 2.2505
R43890 ASIG5V.n2804 ASIG5V.n2803 2.2505
R43891 ASIG5V.n2799 ASIG5V.n2634 2.2505
R43892 ASIG5V.n2795 ASIG5V.n2794 2.2505
R43893 ASIG5V.n2793 ASIG5V.n2635 2.2505
R43894 ASIG5V.n2792 ASIG5V.n2791 2.2505
R43895 ASIG5V.n2787 ASIG5V.n2636 2.2505
R43896 ASIG5V.n2783 ASIG5V.n2782 2.2505
R43897 ASIG5V.n2781 ASIG5V.n2637 2.2505
R43898 ASIG5V.n2780 ASIG5V.n2779 2.2505
R43899 ASIG5V.n2775 ASIG5V.n2638 2.2505
R43900 ASIG5V.n2771 ASIG5V.n2770 2.2505
R43901 ASIG5V.n2769 ASIG5V.n2639 2.2505
R43902 ASIG5V.n2768 ASIG5V.n2767 2.2505
R43903 ASIG5V.n2763 ASIG5V.n2640 2.2505
R43904 ASIG5V.n2759 ASIG5V.n2758 2.2505
R43905 ASIG5V.n2757 ASIG5V.n2641 2.2505
R43906 ASIG5V.n2756 ASIG5V.n2755 2.2505
R43907 ASIG5V.n2751 ASIG5V.n2642 2.2505
R43908 ASIG5V.n2747 ASIG5V.n2746 2.2505
R43909 ASIG5V.n2745 ASIG5V.n2643 2.2505
R43910 ASIG5V.n2744 ASIG5V.n2743 2.2505
R43911 ASIG5V.n2739 ASIG5V.n2644 2.2505
R43912 ASIG5V.n2735 ASIG5V.n2734 2.2505
R43913 ASIG5V.n2733 ASIG5V.n2645 2.2505
R43914 ASIG5V.n2732 ASIG5V.n2731 2.2505
R43915 ASIG5V.n2727 ASIG5V.n2646 2.2505
R43916 ASIG5V.n2723 ASIG5V.n2722 2.2505
R43917 ASIG5V.n2721 ASIG5V.n2647 2.2505
R43918 ASIG5V.n2720 ASIG5V.n2719 2.2505
R43919 ASIG5V.n2715 ASIG5V.n2648 2.2505
R43920 ASIG5V.n2711 ASIG5V.n2710 2.2505
R43921 ASIG5V.n2709 ASIG5V.n2649 2.2505
R43922 ASIG5V.n2708 ASIG5V.n2707 2.2505
R43923 ASIG5V.n2703 ASIG5V.n2650 2.2505
R43924 ASIG5V.n2699 ASIG5V.n2698 2.2505
R43925 ASIG5V.n2697 ASIG5V.n2651 2.2505
R43926 ASIG5V.n2696 ASIG5V.n2695 2.2505
R43927 ASIG5V.n2691 ASIG5V.n2652 2.2505
R43928 ASIG5V.n2687 ASIG5V.n2686 2.2505
R43929 ASIG5V.n2685 ASIG5V.n2653 2.2505
R43930 ASIG5V.n2684 ASIG5V.n2683 2.2505
R43931 ASIG5V.n2679 ASIG5V.n2654 2.2505
R43932 ASIG5V.n2675 ASIG5V.n2674 2.2505
R43933 ASIG5V.n2673 ASIG5V.n2655 2.2505
R43934 ASIG5V.n2672 ASIG5V.n2671 2.2505
R43935 ASIG5V.n2667 ASIG5V.n2656 2.2505
R43936 ASIG5V.n2663 ASIG5V.n2662 2.2505
R43937 ASIG5V.n2661 ASIG5V.n2660 2.2505
R43938 ASIG5V.n2657 ASIG5V.n2563 2.2505
R43939 ASIG5V.n2657 ASIG5V.n2611 2.2505
R43940 ASIG5V.n2660 ASIG5V.n2659 2.2505
R43941 ASIG5V.n2664 ASIG5V.n2663 2.2505
R43942 ASIG5V.n2667 ASIG5V.n2666 2.2505
R43943 ASIG5V.n2671 ASIG5V.n2670 2.2505
R43944 ASIG5V.n2668 ASIG5V.n2655 2.2505
R43945 ASIG5V.n2676 ASIG5V.n2675 2.2505
R43946 ASIG5V.n2679 ASIG5V.n2678 2.2505
R43947 ASIG5V.n2683 ASIG5V.n2682 2.2505
R43948 ASIG5V.n2680 ASIG5V.n2653 2.2505
R43949 ASIG5V.n2688 ASIG5V.n2687 2.2505
R43950 ASIG5V.n2691 ASIG5V.n2690 2.2505
R43951 ASIG5V.n2695 ASIG5V.n2694 2.2505
R43952 ASIG5V.n2692 ASIG5V.n2651 2.2505
R43953 ASIG5V.n2700 ASIG5V.n2699 2.2505
R43954 ASIG5V.n2703 ASIG5V.n2702 2.2505
R43955 ASIG5V.n2707 ASIG5V.n2706 2.2505
R43956 ASIG5V.n2704 ASIG5V.n2649 2.2505
R43957 ASIG5V.n2712 ASIG5V.n2711 2.2505
R43958 ASIG5V.n2715 ASIG5V.n2714 2.2505
R43959 ASIG5V.n2719 ASIG5V.n2718 2.2505
R43960 ASIG5V.n2716 ASIG5V.n2647 2.2505
R43961 ASIG5V.n2724 ASIG5V.n2723 2.2505
R43962 ASIG5V.n2727 ASIG5V.n2726 2.2505
R43963 ASIG5V.n2731 ASIG5V.n2730 2.2505
R43964 ASIG5V.n2728 ASIG5V.n2645 2.2505
R43965 ASIG5V.n2736 ASIG5V.n2735 2.2505
R43966 ASIG5V.n2739 ASIG5V.n2738 2.2505
R43967 ASIG5V.n2743 ASIG5V.n2742 2.2505
R43968 ASIG5V.n2740 ASIG5V.n2643 2.2505
R43969 ASIG5V.n2748 ASIG5V.n2747 2.2505
R43970 ASIG5V.n2751 ASIG5V.n2750 2.2505
R43971 ASIG5V.n2755 ASIG5V.n2754 2.2505
R43972 ASIG5V.n2752 ASIG5V.n2641 2.2505
R43973 ASIG5V.n2760 ASIG5V.n2759 2.2505
R43974 ASIG5V.n2763 ASIG5V.n2762 2.2505
R43975 ASIG5V.n2767 ASIG5V.n2766 2.2505
R43976 ASIG5V.n2764 ASIG5V.n2639 2.2505
R43977 ASIG5V.n2772 ASIG5V.n2771 2.2505
R43978 ASIG5V.n2775 ASIG5V.n2774 2.2505
R43979 ASIG5V.n2779 ASIG5V.n2778 2.2505
R43980 ASIG5V.n2776 ASIG5V.n2637 2.2505
R43981 ASIG5V.n2784 ASIG5V.n2783 2.2505
R43982 ASIG5V.n2787 ASIG5V.n2786 2.2505
R43983 ASIG5V.n2791 ASIG5V.n2790 2.2505
R43984 ASIG5V.n2788 ASIG5V.n2635 2.2505
R43985 ASIG5V.n2796 ASIG5V.n2795 2.2505
R43986 ASIG5V.n2799 ASIG5V.n2798 2.2505
R43987 ASIG5V.n2803 ASIG5V.n2802 2.2505
R43988 ASIG5V.n2800 ASIG5V.n2633 2.2505
R43989 ASIG5V.n2808 ASIG5V.n2807 2.2505
R43990 ASIG5V.n2811 ASIG5V.n2810 2.2505
R43991 ASIG5V.n2815 ASIG5V.n2814 2.2505
R43992 ASIG5V.n2812 ASIG5V.n2631 2.2505
R43993 ASIG5V.n2820 ASIG5V.n2819 2.2505
R43994 ASIG5V.n2823 ASIG5V.n2822 2.2505
R43995 ASIG5V.n2827 ASIG5V.n2826 2.2505
R43996 ASIG5V.n2824 ASIG5V.n2629 2.2505
R43997 ASIG5V.n2832 ASIG5V.n2831 2.2505
R43998 ASIG5V.n2835 ASIG5V.n2834 2.2505
R43999 ASIG5V.n2839 ASIG5V.n2838 2.2505
R44000 ASIG5V.n2836 ASIG5V.n2627 2.2505
R44001 ASIG5V.n2844 ASIG5V.n2843 2.2505
R44002 ASIG5V.n2847 ASIG5V.n2846 2.2505
R44003 ASIG5V.n2851 ASIG5V.n2850 2.2505
R44004 ASIG5V.n2848 ASIG5V.n2625 2.2505
R44005 ASIG5V.n2856 ASIG5V.n2855 2.2505
R44006 ASIG5V.n2859 ASIG5V.n2858 2.2505
R44007 ASIG5V.n2863 ASIG5V.n2862 2.2505
R44008 ASIG5V.n2860 ASIG5V.n2623 2.2505
R44009 ASIG5V.n2868 ASIG5V.n2867 2.2505
R44010 ASIG5V.n2871 ASIG5V.n2870 2.2505
R44011 ASIG5V.n2875 ASIG5V.n2874 2.2505
R44012 ASIG5V.n2872 ASIG5V.n2621 2.2505
R44013 ASIG5V.n2880 ASIG5V.n2879 2.2505
R44014 ASIG5V.n2883 ASIG5V.n2882 2.2505
R44015 ASIG5V.n2887 ASIG5V.n2886 2.2505
R44016 ASIG5V.n2884 ASIG5V.n2619 2.2505
R44017 ASIG5V.n2892 ASIG5V.n2891 2.2505
R44018 ASIG5V.n2895 ASIG5V.n2894 2.2505
R44019 ASIG5V.n2899 ASIG5V.n2898 2.2505
R44020 ASIG5V.n2896 ASIG5V.n2617 2.2505
R44021 ASIG5V.n11768 ASIG5V.n11767 2.2505
R44022 ASIG5V.n11770 ASIG5V.n2614 2.2505
R44023 ASIG5V.n2957 ASIG5V.n2909 2.2505
R44024 ASIG5V.n11747 ASIG5V.n11746 2.2505
R44025 ASIG5V.n11745 ASIG5V.n2959 2.2505
R44026 ASIG5V.n11744 ASIG5V.n11743 2.2505
R44027 ASIG5V.n11739 ASIG5V.n2960 2.2505
R44028 ASIG5V.n11735 ASIG5V.n11734 2.2505
R44029 ASIG5V.n11733 ASIG5V.n2961 2.2505
R44030 ASIG5V.n11732 ASIG5V.n11731 2.2505
R44031 ASIG5V.n11727 ASIG5V.n2962 2.2505
R44032 ASIG5V.n11723 ASIG5V.n11722 2.2505
R44033 ASIG5V.n11721 ASIG5V.n2963 2.2505
R44034 ASIG5V.n11720 ASIG5V.n11719 2.2505
R44035 ASIG5V.n11715 ASIG5V.n2964 2.2505
R44036 ASIG5V.n11711 ASIG5V.n11710 2.2505
R44037 ASIG5V.n11709 ASIG5V.n2965 2.2505
R44038 ASIG5V.n11708 ASIG5V.n11707 2.2505
R44039 ASIG5V.n11703 ASIG5V.n2966 2.2505
R44040 ASIG5V.n11699 ASIG5V.n11698 2.2505
R44041 ASIG5V.n11697 ASIG5V.n2967 2.2505
R44042 ASIG5V.n11696 ASIG5V.n11695 2.2505
R44043 ASIG5V.n11691 ASIG5V.n2968 2.2505
R44044 ASIG5V.n11687 ASIG5V.n11686 2.2505
R44045 ASIG5V.n11685 ASIG5V.n2969 2.2505
R44046 ASIG5V.n11684 ASIG5V.n11683 2.2505
R44047 ASIG5V.n11679 ASIG5V.n2970 2.2505
R44048 ASIG5V.n11675 ASIG5V.n11674 2.2505
R44049 ASIG5V.n11673 ASIG5V.n2971 2.2505
R44050 ASIG5V.n11672 ASIG5V.n11671 2.2505
R44051 ASIG5V.n11667 ASIG5V.n2972 2.2505
R44052 ASIG5V.n11663 ASIG5V.n11662 2.2505
R44053 ASIG5V.n11661 ASIG5V.n2973 2.2505
R44054 ASIG5V.n11660 ASIG5V.n11659 2.2505
R44055 ASIG5V.n11655 ASIG5V.n2974 2.2505
R44056 ASIG5V.n11651 ASIG5V.n11650 2.2505
R44057 ASIG5V.n11649 ASIG5V.n2975 2.2505
R44058 ASIG5V.n11648 ASIG5V.n11647 2.2505
R44059 ASIG5V.n11643 ASIG5V.n2976 2.2505
R44060 ASIG5V.n11639 ASIG5V.n11638 2.2505
R44061 ASIG5V.n11637 ASIG5V.n2977 2.2505
R44062 ASIG5V.n11636 ASIG5V.n11635 2.2505
R44063 ASIG5V.n11631 ASIG5V.n2978 2.2505
R44064 ASIG5V.n11627 ASIG5V.n11626 2.2505
R44065 ASIG5V.n11625 ASIG5V.n2979 2.2505
R44066 ASIG5V.n11624 ASIG5V.n11623 2.2505
R44067 ASIG5V.n11619 ASIG5V.n2980 2.2505
R44068 ASIG5V.n11615 ASIG5V.n11614 2.2505
R44069 ASIG5V.n11613 ASIG5V.n2981 2.2505
R44070 ASIG5V.n11612 ASIG5V.n11611 2.2505
R44071 ASIG5V.n11607 ASIG5V.n2982 2.2505
R44072 ASIG5V.n11603 ASIG5V.n11602 2.2505
R44073 ASIG5V.n11601 ASIG5V.n2983 2.2505
R44074 ASIG5V.n11600 ASIG5V.n11599 2.2505
R44075 ASIG5V.n11595 ASIG5V.n2984 2.2505
R44076 ASIG5V.n11591 ASIG5V.n11590 2.2505
R44077 ASIG5V.n11589 ASIG5V.n2985 2.2505
R44078 ASIG5V.n11588 ASIG5V.n11587 2.2505
R44079 ASIG5V.n11583 ASIG5V.n2986 2.2505
R44080 ASIG5V.n11579 ASIG5V.n11578 2.2505
R44081 ASIG5V.n11577 ASIG5V.n2987 2.2505
R44082 ASIG5V.n11576 ASIG5V.n11575 2.2505
R44083 ASIG5V.n11571 ASIG5V.n2988 2.2505
R44084 ASIG5V.n11567 ASIG5V.n11566 2.2505
R44085 ASIG5V.n11565 ASIG5V.n2989 2.2505
R44086 ASIG5V.n11564 ASIG5V.n11563 2.2505
R44087 ASIG5V.n11559 ASIG5V.n2990 2.2505
R44088 ASIG5V.n11555 ASIG5V.n11554 2.2505
R44089 ASIG5V.n11553 ASIG5V.n2991 2.2505
R44090 ASIG5V.n11552 ASIG5V.n11551 2.2505
R44091 ASIG5V.n11547 ASIG5V.n2992 2.2505
R44092 ASIG5V.n11543 ASIG5V.n11542 2.2505
R44093 ASIG5V.n11541 ASIG5V.n2993 2.2505
R44094 ASIG5V.n11540 ASIG5V.n11539 2.2505
R44095 ASIG5V.n11535 ASIG5V.n2994 2.2505
R44096 ASIG5V.n11531 ASIG5V.n11530 2.2505
R44097 ASIG5V.n11529 ASIG5V.n2995 2.2505
R44098 ASIG5V.n11528 ASIG5V.n11527 2.2505
R44099 ASIG5V.n11523 ASIG5V.n2996 2.2505
R44100 ASIG5V.n11519 ASIG5V.n11518 2.2505
R44101 ASIG5V.n11517 ASIG5V.n2997 2.2505
R44102 ASIG5V.n11516 ASIG5V.n11515 2.2505
R44103 ASIG5V.n11511 ASIG5V.n2998 2.2505
R44104 ASIG5V.n11507 ASIG5V.n11506 2.2505
R44105 ASIG5V.n11505 ASIG5V.n3001 2.2505
R44106 ASIG5V.n11504 ASIG5V.n11503 2.2505
R44107 ASIG5V.n11503 ASIG5V.n2955 2.2505
R44108 ASIG5V.n3001 ASIG5V.n3000 2.2505
R44109 ASIG5V.n11508 ASIG5V.n11507 2.2505
R44110 ASIG5V.n11511 ASIG5V.n11510 2.2505
R44111 ASIG5V.n11515 ASIG5V.n11514 2.2505
R44112 ASIG5V.n11512 ASIG5V.n2997 2.2505
R44113 ASIG5V.n11520 ASIG5V.n11519 2.2505
R44114 ASIG5V.n11523 ASIG5V.n11522 2.2505
R44115 ASIG5V.n11527 ASIG5V.n11526 2.2505
R44116 ASIG5V.n11524 ASIG5V.n2995 2.2505
R44117 ASIG5V.n11532 ASIG5V.n11531 2.2505
R44118 ASIG5V.n11535 ASIG5V.n11534 2.2505
R44119 ASIG5V.n11539 ASIG5V.n11538 2.2505
R44120 ASIG5V.n11536 ASIG5V.n2993 2.2505
R44121 ASIG5V.n11544 ASIG5V.n11543 2.2505
R44122 ASIG5V.n11547 ASIG5V.n11546 2.2505
R44123 ASIG5V.n11551 ASIG5V.n11550 2.2505
R44124 ASIG5V.n11548 ASIG5V.n2991 2.2505
R44125 ASIG5V.n11556 ASIG5V.n11555 2.2505
R44126 ASIG5V.n11559 ASIG5V.n11558 2.2505
R44127 ASIG5V.n11563 ASIG5V.n11562 2.2505
R44128 ASIG5V.n11560 ASIG5V.n2989 2.2505
R44129 ASIG5V.n11568 ASIG5V.n11567 2.2505
R44130 ASIG5V.n11571 ASIG5V.n11570 2.2505
R44131 ASIG5V.n11575 ASIG5V.n11574 2.2505
R44132 ASIG5V.n11572 ASIG5V.n2987 2.2505
R44133 ASIG5V.n11580 ASIG5V.n11579 2.2505
R44134 ASIG5V.n11583 ASIG5V.n11582 2.2505
R44135 ASIG5V.n11587 ASIG5V.n11586 2.2505
R44136 ASIG5V.n11584 ASIG5V.n2985 2.2505
R44137 ASIG5V.n11592 ASIG5V.n11591 2.2505
R44138 ASIG5V.n11595 ASIG5V.n11594 2.2505
R44139 ASIG5V.n11599 ASIG5V.n11598 2.2505
R44140 ASIG5V.n11596 ASIG5V.n2983 2.2505
R44141 ASIG5V.n11604 ASIG5V.n11603 2.2505
R44142 ASIG5V.n11607 ASIG5V.n11606 2.2505
R44143 ASIG5V.n11611 ASIG5V.n11610 2.2505
R44144 ASIG5V.n11608 ASIG5V.n2981 2.2505
R44145 ASIG5V.n11616 ASIG5V.n11615 2.2505
R44146 ASIG5V.n11619 ASIG5V.n11618 2.2505
R44147 ASIG5V.n11623 ASIG5V.n11622 2.2505
R44148 ASIG5V.n11620 ASIG5V.n2979 2.2505
R44149 ASIG5V.n11628 ASIG5V.n11627 2.2505
R44150 ASIG5V.n11631 ASIG5V.n11630 2.2505
R44151 ASIG5V.n11635 ASIG5V.n11634 2.2505
R44152 ASIG5V.n11632 ASIG5V.n2977 2.2505
R44153 ASIG5V.n11640 ASIG5V.n11639 2.2505
R44154 ASIG5V.n11643 ASIG5V.n11642 2.2505
R44155 ASIG5V.n11647 ASIG5V.n11646 2.2505
R44156 ASIG5V.n11644 ASIG5V.n2975 2.2505
R44157 ASIG5V.n11652 ASIG5V.n11651 2.2505
R44158 ASIG5V.n11655 ASIG5V.n11654 2.2505
R44159 ASIG5V.n11659 ASIG5V.n11658 2.2505
R44160 ASIG5V.n11656 ASIG5V.n2973 2.2505
R44161 ASIG5V.n11664 ASIG5V.n11663 2.2505
R44162 ASIG5V.n11667 ASIG5V.n11666 2.2505
R44163 ASIG5V.n11671 ASIG5V.n11670 2.2505
R44164 ASIG5V.n11668 ASIG5V.n2971 2.2505
R44165 ASIG5V.n11676 ASIG5V.n11675 2.2505
R44166 ASIG5V.n11679 ASIG5V.n11678 2.2505
R44167 ASIG5V.n11683 ASIG5V.n11682 2.2505
R44168 ASIG5V.n11680 ASIG5V.n2969 2.2505
R44169 ASIG5V.n11688 ASIG5V.n11687 2.2505
R44170 ASIG5V.n11691 ASIG5V.n11690 2.2505
R44171 ASIG5V.n11695 ASIG5V.n11694 2.2505
R44172 ASIG5V.n11692 ASIG5V.n2967 2.2505
R44173 ASIG5V.n11700 ASIG5V.n11699 2.2505
R44174 ASIG5V.n11703 ASIG5V.n11702 2.2505
R44175 ASIG5V.n11707 ASIG5V.n11706 2.2505
R44176 ASIG5V.n11704 ASIG5V.n2965 2.2505
R44177 ASIG5V.n11712 ASIG5V.n11711 2.2505
R44178 ASIG5V.n11715 ASIG5V.n11714 2.2505
R44179 ASIG5V.n11719 ASIG5V.n11718 2.2505
R44180 ASIG5V.n11716 ASIG5V.n2963 2.2505
R44181 ASIG5V.n11724 ASIG5V.n11723 2.2505
R44182 ASIG5V.n11727 ASIG5V.n11726 2.2505
R44183 ASIG5V.n11731 ASIG5V.n11730 2.2505
R44184 ASIG5V.n11728 ASIG5V.n2961 2.2505
R44185 ASIG5V.n11736 ASIG5V.n11735 2.2505
R44186 ASIG5V.n11739 ASIG5V.n11738 2.2505
R44187 ASIG5V.n11743 ASIG5V.n11742 2.2505
R44188 ASIG5V.n11740 ASIG5V.n2959 2.2505
R44189 ASIG5V.n11748 ASIG5V.n11747 2.2505
R44190 ASIG5V.n11750 ASIG5V.n2957 2.2505
R44191 ASIG5V.n11193 ASIG5V.n9969 2.2505
R44192 ASIG5V.n11481 ASIG5V.n11480 2.2505
R44193 ASIG5V.n11479 ASIG5V.n11194 2.2505
R44194 ASIG5V.n11478 ASIG5V.n11477 2.2505
R44195 ASIG5V.n11473 ASIG5V.n11195 2.2505
R44196 ASIG5V.n11469 ASIG5V.n11468 2.2505
R44197 ASIG5V.n11467 ASIG5V.n11196 2.2505
R44198 ASIG5V.n11466 ASIG5V.n11465 2.2505
R44199 ASIG5V.n11461 ASIG5V.n11197 2.2505
R44200 ASIG5V.n11457 ASIG5V.n11456 2.2505
R44201 ASIG5V.n11455 ASIG5V.n11198 2.2505
R44202 ASIG5V.n11454 ASIG5V.n11453 2.2505
R44203 ASIG5V.n11449 ASIG5V.n11199 2.2505
R44204 ASIG5V.n11445 ASIG5V.n11444 2.2505
R44205 ASIG5V.n11443 ASIG5V.n11200 2.2505
R44206 ASIG5V.n11442 ASIG5V.n11441 2.2505
R44207 ASIG5V.n11437 ASIG5V.n11201 2.2505
R44208 ASIG5V.n11433 ASIG5V.n11432 2.2505
R44209 ASIG5V.n11431 ASIG5V.n11202 2.2505
R44210 ASIG5V.n11430 ASIG5V.n11429 2.2505
R44211 ASIG5V.n11425 ASIG5V.n11203 2.2505
R44212 ASIG5V.n11421 ASIG5V.n11420 2.2505
R44213 ASIG5V.n11419 ASIG5V.n11204 2.2505
R44214 ASIG5V.n11418 ASIG5V.n11417 2.2505
R44215 ASIG5V.n11413 ASIG5V.n11205 2.2505
R44216 ASIG5V.n11409 ASIG5V.n11408 2.2505
R44217 ASIG5V.n11407 ASIG5V.n11206 2.2505
R44218 ASIG5V.n11406 ASIG5V.n11405 2.2505
R44219 ASIG5V.n11401 ASIG5V.n11207 2.2505
R44220 ASIG5V.n11397 ASIG5V.n11396 2.2505
R44221 ASIG5V.n11395 ASIG5V.n11208 2.2505
R44222 ASIG5V.n11394 ASIG5V.n11393 2.2505
R44223 ASIG5V.n11389 ASIG5V.n11209 2.2505
R44224 ASIG5V.n11385 ASIG5V.n11384 2.2505
R44225 ASIG5V.n11383 ASIG5V.n11210 2.2505
R44226 ASIG5V.n11382 ASIG5V.n11381 2.2505
R44227 ASIG5V.n11377 ASIG5V.n11211 2.2505
R44228 ASIG5V.n11373 ASIG5V.n11372 2.2505
R44229 ASIG5V.n11371 ASIG5V.n11212 2.2505
R44230 ASIG5V.n11370 ASIG5V.n11369 2.2505
R44231 ASIG5V.n11365 ASIG5V.n11213 2.2505
R44232 ASIG5V.n11361 ASIG5V.n11360 2.2505
R44233 ASIG5V.n11359 ASIG5V.n11214 2.2505
R44234 ASIG5V.n11358 ASIG5V.n11357 2.2505
R44235 ASIG5V.n11353 ASIG5V.n11215 2.2505
R44236 ASIG5V.n11349 ASIG5V.n11348 2.2505
R44237 ASIG5V.n11347 ASIG5V.n11216 2.2505
R44238 ASIG5V.n11346 ASIG5V.n11345 2.2505
R44239 ASIG5V.n11341 ASIG5V.n11217 2.2505
R44240 ASIG5V.n11337 ASIG5V.n11336 2.2505
R44241 ASIG5V.n11335 ASIG5V.n11218 2.2505
R44242 ASIG5V.n11334 ASIG5V.n11333 2.2505
R44243 ASIG5V.n11329 ASIG5V.n11219 2.2505
R44244 ASIG5V.n11325 ASIG5V.n11324 2.2505
R44245 ASIG5V.n11323 ASIG5V.n11220 2.2505
R44246 ASIG5V.n11322 ASIG5V.n11321 2.2505
R44247 ASIG5V.n11317 ASIG5V.n11221 2.2505
R44248 ASIG5V.n11313 ASIG5V.n11312 2.2505
R44249 ASIG5V.n11311 ASIG5V.n11222 2.2505
R44250 ASIG5V.n11310 ASIG5V.n11309 2.2505
R44251 ASIG5V.n11305 ASIG5V.n11223 2.2505
R44252 ASIG5V.n11301 ASIG5V.n11300 2.2505
R44253 ASIG5V.n11299 ASIG5V.n11224 2.2505
R44254 ASIG5V.n11298 ASIG5V.n11297 2.2505
R44255 ASIG5V.n11293 ASIG5V.n11225 2.2505
R44256 ASIG5V.n11289 ASIG5V.n11288 2.2505
R44257 ASIG5V.n11287 ASIG5V.n11226 2.2505
R44258 ASIG5V.n11286 ASIG5V.n11285 2.2505
R44259 ASIG5V.n11281 ASIG5V.n11227 2.2505
R44260 ASIG5V.n11277 ASIG5V.n11276 2.2505
R44261 ASIG5V.n11275 ASIG5V.n11228 2.2505
R44262 ASIG5V.n11274 ASIG5V.n11273 2.2505
R44263 ASIG5V.n11269 ASIG5V.n11229 2.2505
R44264 ASIG5V.n11265 ASIG5V.n11264 2.2505
R44265 ASIG5V.n11263 ASIG5V.n11230 2.2505
R44266 ASIG5V.n11262 ASIG5V.n11261 2.2505
R44267 ASIG5V.n11257 ASIG5V.n11231 2.2505
R44268 ASIG5V.n11253 ASIG5V.n11252 2.2505
R44269 ASIG5V.n11251 ASIG5V.n11232 2.2505
R44270 ASIG5V.n11250 ASIG5V.n11249 2.2505
R44271 ASIG5V.n11245 ASIG5V.n11233 2.2505
R44272 ASIG5V.n11241 ASIG5V.n11240 2.2505
R44273 ASIG5V.n11239 ASIG5V.n11236 2.2505
R44274 ASIG5V.n11238 ASIG5V.n11237 2.2505
R44275 ASIG5V.n11237 ASIG5V.n10015 2.2505
R44276 ASIG5V.n11236 ASIG5V.n11235 2.2505
R44277 ASIG5V.n11242 ASIG5V.n11241 2.2505
R44278 ASIG5V.n11245 ASIG5V.n11244 2.2505
R44279 ASIG5V.n11249 ASIG5V.n11248 2.2505
R44280 ASIG5V.n11246 ASIG5V.n11232 2.2505
R44281 ASIG5V.n11254 ASIG5V.n11253 2.2505
R44282 ASIG5V.n11257 ASIG5V.n11256 2.2505
R44283 ASIG5V.n11261 ASIG5V.n11260 2.2505
R44284 ASIG5V.n11258 ASIG5V.n11230 2.2505
R44285 ASIG5V.n11266 ASIG5V.n11265 2.2505
R44286 ASIG5V.n11269 ASIG5V.n11268 2.2505
R44287 ASIG5V.n11273 ASIG5V.n11272 2.2505
R44288 ASIG5V.n11270 ASIG5V.n11228 2.2505
R44289 ASIG5V.n11278 ASIG5V.n11277 2.2505
R44290 ASIG5V.n11281 ASIG5V.n11280 2.2505
R44291 ASIG5V.n11285 ASIG5V.n11284 2.2505
R44292 ASIG5V.n11282 ASIG5V.n11226 2.2505
R44293 ASIG5V.n11290 ASIG5V.n11289 2.2505
R44294 ASIG5V.n11293 ASIG5V.n11292 2.2505
R44295 ASIG5V.n11297 ASIG5V.n11296 2.2505
R44296 ASIG5V.n11294 ASIG5V.n11224 2.2505
R44297 ASIG5V.n11302 ASIG5V.n11301 2.2505
R44298 ASIG5V.n11305 ASIG5V.n11304 2.2505
R44299 ASIG5V.n11309 ASIG5V.n11308 2.2505
R44300 ASIG5V.n11306 ASIG5V.n11222 2.2505
R44301 ASIG5V.n11314 ASIG5V.n11313 2.2505
R44302 ASIG5V.n11317 ASIG5V.n11316 2.2505
R44303 ASIG5V.n11321 ASIG5V.n11320 2.2505
R44304 ASIG5V.n11318 ASIG5V.n11220 2.2505
R44305 ASIG5V.n11326 ASIG5V.n11325 2.2505
R44306 ASIG5V.n11329 ASIG5V.n11328 2.2505
R44307 ASIG5V.n11333 ASIG5V.n11332 2.2505
R44308 ASIG5V.n11330 ASIG5V.n11218 2.2505
R44309 ASIG5V.n11338 ASIG5V.n11337 2.2505
R44310 ASIG5V.n11341 ASIG5V.n11340 2.2505
R44311 ASIG5V.n11345 ASIG5V.n11344 2.2505
R44312 ASIG5V.n11342 ASIG5V.n11216 2.2505
R44313 ASIG5V.n11350 ASIG5V.n11349 2.2505
R44314 ASIG5V.n11353 ASIG5V.n11352 2.2505
R44315 ASIG5V.n11357 ASIG5V.n11356 2.2505
R44316 ASIG5V.n11354 ASIG5V.n11214 2.2505
R44317 ASIG5V.n11362 ASIG5V.n11361 2.2505
R44318 ASIG5V.n11365 ASIG5V.n11364 2.2505
R44319 ASIG5V.n11369 ASIG5V.n11368 2.2505
R44320 ASIG5V.n11366 ASIG5V.n11212 2.2505
R44321 ASIG5V.n11374 ASIG5V.n11373 2.2505
R44322 ASIG5V.n11377 ASIG5V.n11376 2.2505
R44323 ASIG5V.n11381 ASIG5V.n11380 2.2505
R44324 ASIG5V.n11378 ASIG5V.n11210 2.2505
R44325 ASIG5V.n11386 ASIG5V.n11385 2.2505
R44326 ASIG5V.n11389 ASIG5V.n11388 2.2505
R44327 ASIG5V.n11393 ASIG5V.n11392 2.2505
R44328 ASIG5V.n11390 ASIG5V.n11208 2.2505
R44329 ASIG5V.n11398 ASIG5V.n11397 2.2505
R44330 ASIG5V.n11401 ASIG5V.n11400 2.2505
R44331 ASIG5V.n11405 ASIG5V.n11404 2.2505
R44332 ASIG5V.n11402 ASIG5V.n11206 2.2505
R44333 ASIG5V.n11410 ASIG5V.n11409 2.2505
R44334 ASIG5V.n11413 ASIG5V.n11412 2.2505
R44335 ASIG5V.n11417 ASIG5V.n11416 2.2505
R44336 ASIG5V.n11414 ASIG5V.n11204 2.2505
R44337 ASIG5V.n11422 ASIG5V.n11421 2.2505
R44338 ASIG5V.n11425 ASIG5V.n11424 2.2505
R44339 ASIG5V.n11429 ASIG5V.n11428 2.2505
R44340 ASIG5V.n11426 ASIG5V.n11202 2.2505
R44341 ASIG5V.n11434 ASIG5V.n11433 2.2505
R44342 ASIG5V.n11437 ASIG5V.n11436 2.2505
R44343 ASIG5V.n11441 ASIG5V.n11440 2.2505
R44344 ASIG5V.n11438 ASIG5V.n11200 2.2505
R44345 ASIG5V.n11446 ASIG5V.n11445 2.2505
R44346 ASIG5V.n11449 ASIG5V.n11448 2.2505
R44347 ASIG5V.n11453 ASIG5V.n11452 2.2505
R44348 ASIG5V.n11450 ASIG5V.n11198 2.2505
R44349 ASIG5V.n11458 ASIG5V.n11457 2.2505
R44350 ASIG5V.n11461 ASIG5V.n11460 2.2505
R44351 ASIG5V.n11465 ASIG5V.n11464 2.2505
R44352 ASIG5V.n11462 ASIG5V.n11196 2.2505
R44353 ASIG5V.n11470 ASIG5V.n11469 2.2505
R44354 ASIG5V.n11473 ASIG5V.n11472 2.2505
R44355 ASIG5V.n11477 ASIG5V.n11476 2.2505
R44356 ASIG5V.n11474 ASIG5V.n11194 2.2505
R44357 ASIG5V.n11482 ASIG5V.n11481 2.2505
R44358 ASIG5V.n11484 ASIG5V.n11193 2.2505
R44359 ASIG5V.n4770 ASIG5V.n3623 2.2505
R44360 ASIG5V.n4769 ASIG5V.n4767 2.2505
R44361 ASIG5V.n4766 ASIG5V.n3717 2.2505
R44362 ASIG5V.n4765 ASIG5V.n4764 2.2505
R44363 ASIG5V.n4762 ASIG5V.n3718 2.2505
R44364 ASIG5V.n4760 ASIG5V.n4758 2.2505
R44365 ASIG5V.n4757 ASIG5V.n3720 2.2505
R44366 ASIG5V.n4756 ASIG5V.n4755 2.2505
R44367 ASIG5V.n4753 ASIG5V.n3721 2.2505
R44368 ASIG5V.n4751 ASIG5V.n4749 2.2505
R44369 ASIG5V.n4748 ASIG5V.n3723 2.2505
R44370 ASIG5V.n4747 ASIG5V.n4746 2.2505
R44371 ASIG5V.n4744 ASIG5V.n3724 2.2505
R44372 ASIG5V.n4742 ASIG5V.n4740 2.2505
R44373 ASIG5V.n4739 ASIG5V.n3726 2.2505
R44374 ASIG5V.n4738 ASIG5V.n4737 2.2505
R44375 ASIG5V.n4735 ASIG5V.n3727 2.2505
R44376 ASIG5V.n4733 ASIG5V.n4731 2.2505
R44377 ASIG5V.n4730 ASIG5V.n3729 2.2505
R44378 ASIG5V.n4729 ASIG5V.n4728 2.2505
R44379 ASIG5V.n4726 ASIG5V.n3730 2.2505
R44380 ASIG5V.n4724 ASIG5V.n4722 2.2505
R44381 ASIG5V.n4721 ASIG5V.n3732 2.2505
R44382 ASIG5V.n4720 ASIG5V.n4719 2.2505
R44383 ASIG5V.n4717 ASIG5V.n3733 2.2505
R44384 ASIG5V.n4715 ASIG5V.n4713 2.2505
R44385 ASIG5V.n4712 ASIG5V.n3735 2.2505
R44386 ASIG5V.n4711 ASIG5V.n4710 2.2505
R44387 ASIG5V.n4708 ASIG5V.n3736 2.2505
R44388 ASIG5V.n4706 ASIG5V.n4704 2.2505
R44389 ASIG5V.n4703 ASIG5V.n3738 2.2505
R44390 ASIG5V.n4702 ASIG5V.n4701 2.2505
R44391 ASIG5V.n4699 ASIG5V.n3739 2.2505
R44392 ASIG5V.n4697 ASIG5V.n4695 2.2505
R44393 ASIG5V.n4694 ASIG5V.n3741 2.2505
R44394 ASIG5V.n4693 ASIG5V.n4692 2.2505
R44395 ASIG5V.n4690 ASIG5V.n3742 2.2505
R44396 ASIG5V.n4688 ASIG5V.n4686 2.2505
R44397 ASIG5V.n4685 ASIG5V.n3744 2.2505
R44398 ASIG5V.n4684 ASIG5V.n4683 2.2505
R44399 ASIG5V.n4681 ASIG5V.n3745 2.2505
R44400 ASIG5V.n4679 ASIG5V.n4677 2.2505
R44401 ASIG5V.n4676 ASIG5V.n3747 2.2505
R44402 ASIG5V.n4675 ASIG5V.n4674 2.2505
R44403 ASIG5V.n4672 ASIG5V.n3748 2.2505
R44404 ASIG5V.n4670 ASIG5V.n4668 2.2505
R44405 ASIG5V.n4667 ASIG5V.n3750 2.2505
R44406 ASIG5V.n4666 ASIG5V.n4665 2.2505
R44407 ASIG5V.n4663 ASIG5V.n3751 2.2505
R44408 ASIG5V.n4661 ASIG5V.n4659 2.2505
R44409 ASIG5V.n4658 ASIG5V.n3753 2.2505
R44410 ASIG5V.n4657 ASIG5V.n4656 2.2505
R44411 ASIG5V.n4654 ASIG5V.n3754 2.2505
R44412 ASIG5V.n4652 ASIG5V.n4650 2.2505
R44413 ASIG5V.n4649 ASIG5V.n3756 2.2505
R44414 ASIG5V.n4648 ASIG5V.n4647 2.2505
R44415 ASIG5V.n4645 ASIG5V.n3757 2.2505
R44416 ASIG5V.n4643 ASIG5V.n4641 2.2505
R44417 ASIG5V.n4640 ASIG5V.n3759 2.2505
R44418 ASIG5V.n4639 ASIG5V.n4638 2.2505
R44419 ASIG5V.n4636 ASIG5V.n3760 2.2505
R44420 ASIG5V.n4634 ASIG5V.n4632 2.2505
R44421 ASIG5V.n4631 ASIG5V.n3762 2.2505
R44422 ASIG5V.n4630 ASIG5V.n4629 2.2505
R44423 ASIG5V.n4627 ASIG5V.n3763 2.2505
R44424 ASIG5V.n4625 ASIG5V.n4623 2.2505
R44425 ASIG5V.n4622 ASIG5V.n3765 2.2505
R44426 ASIG5V.n4621 ASIG5V.n4620 2.2505
R44427 ASIG5V.n4618 ASIG5V.n3766 2.2505
R44428 ASIG5V.n4616 ASIG5V.n4614 2.2505
R44429 ASIG5V.n4613 ASIG5V.n3768 2.2505
R44430 ASIG5V.n4612 ASIG5V.n4611 2.2505
R44431 ASIG5V.n4609 ASIG5V.n3769 2.2505
R44432 ASIG5V.n4607 ASIG5V.n4605 2.2505
R44433 ASIG5V.n4604 ASIG5V.n3771 2.2505
R44434 ASIG5V.n4603 ASIG5V.n4602 2.2505
R44435 ASIG5V.n4600 ASIG5V.n3772 2.2505
R44436 ASIG5V.n4598 ASIG5V.n4596 2.2505
R44437 ASIG5V.n4595 ASIG5V.n3774 2.2505
R44438 ASIG5V.n4594 ASIG5V.n4593 2.2505
R44439 ASIG5V.n4591 ASIG5V.n3775 2.2505
R44440 ASIG5V.n4589 ASIG5V.n4587 2.2505
R44441 ASIG5V.n4586 ASIG5V.n3776 2.2505
R44442 ASIG5V.n4585 ASIG5V.n3673 2.2505
R44443 ASIG5V.n4773 ASIG5V.n3673 2.2505
R44444 ASIG5V.n3776 ASIG5V.n3671 2.2505
R44445 ASIG5V.n4589 ASIG5V.n4588 2.2505
R44446 ASIG5V.n4591 ASIG5V.n4590 2.2505
R44447 ASIG5V.n4593 ASIG5V.n4592 2.2505
R44448 ASIG5V.n3774 ASIG5V.n3773 2.2505
R44449 ASIG5V.n4598 ASIG5V.n4597 2.2505
R44450 ASIG5V.n4600 ASIG5V.n4599 2.2505
R44451 ASIG5V.n4602 ASIG5V.n4601 2.2505
R44452 ASIG5V.n3771 ASIG5V.n3770 2.2505
R44453 ASIG5V.n4607 ASIG5V.n4606 2.2505
R44454 ASIG5V.n4609 ASIG5V.n4608 2.2505
R44455 ASIG5V.n4611 ASIG5V.n4610 2.2505
R44456 ASIG5V.n3768 ASIG5V.n3767 2.2505
R44457 ASIG5V.n4616 ASIG5V.n4615 2.2505
R44458 ASIG5V.n4618 ASIG5V.n4617 2.2505
R44459 ASIG5V.n4620 ASIG5V.n4619 2.2505
R44460 ASIG5V.n3765 ASIG5V.n3764 2.2505
R44461 ASIG5V.n4625 ASIG5V.n4624 2.2505
R44462 ASIG5V.n4627 ASIG5V.n4626 2.2505
R44463 ASIG5V.n4629 ASIG5V.n4628 2.2505
R44464 ASIG5V.n3762 ASIG5V.n3761 2.2505
R44465 ASIG5V.n4634 ASIG5V.n4633 2.2505
R44466 ASIG5V.n4636 ASIG5V.n4635 2.2505
R44467 ASIG5V.n4638 ASIG5V.n4637 2.2505
R44468 ASIG5V.n3759 ASIG5V.n3758 2.2505
R44469 ASIG5V.n4643 ASIG5V.n4642 2.2505
R44470 ASIG5V.n4645 ASIG5V.n4644 2.2505
R44471 ASIG5V.n4647 ASIG5V.n4646 2.2505
R44472 ASIG5V.n3756 ASIG5V.n3755 2.2505
R44473 ASIG5V.n4652 ASIG5V.n4651 2.2505
R44474 ASIG5V.n4654 ASIG5V.n4653 2.2505
R44475 ASIG5V.n4656 ASIG5V.n4655 2.2505
R44476 ASIG5V.n3753 ASIG5V.n3752 2.2505
R44477 ASIG5V.n4661 ASIG5V.n4660 2.2505
R44478 ASIG5V.n4663 ASIG5V.n4662 2.2505
R44479 ASIG5V.n4665 ASIG5V.n4664 2.2505
R44480 ASIG5V.n3750 ASIG5V.n3749 2.2505
R44481 ASIG5V.n4670 ASIG5V.n4669 2.2505
R44482 ASIG5V.n4672 ASIG5V.n4671 2.2505
R44483 ASIG5V.n4674 ASIG5V.n4673 2.2505
R44484 ASIG5V.n3747 ASIG5V.n3746 2.2505
R44485 ASIG5V.n4679 ASIG5V.n4678 2.2505
R44486 ASIG5V.n4681 ASIG5V.n4680 2.2505
R44487 ASIG5V.n4683 ASIG5V.n4682 2.2505
R44488 ASIG5V.n3744 ASIG5V.n3743 2.2505
R44489 ASIG5V.n4688 ASIG5V.n4687 2.2505
R44490 ASIG5V.n4690 ASIG5V.n4689 2.2505
R44491 ASIG5V.n4692 ASIG5V.n4691 2.2505
R44492 ASIG5V.n3741 ASIG5V.n3740 2.2505
R44493 ASIG5V.n4697 ASIG5V.n4696 2.2505
R44494 ASIG5V.n4699 ASIG5V.n4698 2.2505
R44495 ASIG5V.n4701 ASIG5V.n4700 2.2505
R44496 ASIG5V.n3738 ASIG5V.n3737 2.2505
R44497 ASIG5V.n4706 ASIG5V.n4705 2.2505
R44498 ASIG5V.n4708 ASIG5V.n4707 2.2505
R44499 ASIG5V.n4710 ASIG5V.n4709 2.2505
R44500 ASIG5V.n3735 ASIG5V.n3734 2.2505
R44501 ASIG5V.n4715 ASIG5V.n4714 2.2505
R44502 ASIG5V.n4717 ASIG5V.n4716 2.2505
R44503 ASIG5V.n4719 ASIG5V.n4718 2.2505
R44504 ASIG5V.n3732 ASIG5V.n3731 2.2505
R44505 ASIG5V.n4724 ASIG5V.n4723 2.2505
R44506 ASIG5V.n4726 ASIG5V.n4725 2.2505
R44507 ASIG5V.n4728 ASIG5V.n4727 2.2505
R44508 ASIG5V.n3729 ASIG5V.n3728 2.2505
R44509 ASIG5V.n4733 ASIG5V.n4732 2.2505
R44510 ASIG5V.n4735 ASIG5V.n4734 2.2505
R44511 ASIG5V.n4737 ASIG5V.n4736 2.2505
R44512 ASIG5V.n3726 ASIG5V.n3725 2.2505
R44513 ASIG5V.n4742 ASIG5V.n4741 2.2505
R44514 ASIG5V.n4744 ASIG5V.n4743 2.2505
R44515 ASIG5V.n4746 ASIG5V.n4745 2.2505
R44516 ASIG5V.n3723 ASIG5V.n3722 2.2505
R44517 ASIG5V.n4751 ASIG5V.n4750 2.2505
R44518 ASIG5V.n4753 ASIG5V.n4752 2.2505
R44519 ASIG5V.n4755 ASIG5V.n4754 2.2505
R44520 ASIG5V.n3720 ASIG5V.n3719 2.2505
R44521 ASIG5V.n4760 ASIG5V.n4759 2.2505
R44522 ASIG5V.n4762 ASIG5V.n4761 2.2505
R44523 ASIG5V.n4764 ASIG5V.n4763 2.2505
R44524 ASIG5V.n3717 ASIG5V.n3716 2.2505
R44525 ASIG5V.n4769 ASIG5V.n4768 2.2505
R44526 ASIG5V.n4771 ASIG5V.n4770 2.2505
R44527 ASIG5V.n3840 ASIG5V.n3839 2.2505
R44528 ASIG5V.n4557 ASIG5V.n4556 2.2505
R44529 ASIG5V.n4558 ASIG5V.n3787 2.2505
R44530 ASIG5V.n4561 ASIG5V.n3830 2.2505
R44531 ASIG5V.n3780 ASIG5V.n3627 2.2505
R44532 ASIG5V.n4778 ASIG5V.n4777 2.2505
R44533 ASIG5V.n3621 ASIG5V.n3620 2.2505
R44534 ASIG5V.n4786 ASIG5V.n4785 2.2505
R44535 ASIG5V.n4800 ASIG5V.n4799 2.2505
R44536 ASIG5V.n3277 ASIG5V.n3271 2.2505
R44537 ASIG5V.n4807 ASIG5V.n4806 2.2505
R44538 ASIG5V.n5066 ASIG5V.n5065 2.2505
R44539 ASIG5V.n3171 ASIG5V.n3169 2.2505
R44540 ASIG5V.n9743 ASIG5V.n9742 2.2505
R44541 ASIG5V.n9736 ASIG5V.n9735 2.2505
R44542 ASIG5V.n5117 ASIG5V.n5073 2.2505
R44543 ASIG5V.n5459 ASIG5V.n5123 2.2505
R44544 ASIG5V.n9422 ASIG5V.n5166 2.2505
R44545 ASIG5V.n9421 ASIG5V.n9420 2.2505
R44546 ASIG5V.n5510 ASIG5V.n5463 2.2505
R44547 ASIG5V.n5560 ASIG5V.n5553 2.2505
R44548 ASIG5V.n7977 ASIG5V.n5565 2.2505
R44549 ASIG5V.n9407 ASIG5V.n9406 2.2505
R44550 ASIG5V.n6254 ASIG5V.n6253 2.2505
R44551 ASIG5V.n6251 ASIG5V.n5912 2.2505
R44552 ASIG5V.n6250 ASIG5V.n5957 2.2505
R44553 ASIG5V.n6263 ASIG5V.n6261 2.2505
R44554 ASIG5V.n9384 ASIG5V.n9383 2.2505
R44555 ASIG5V.n6437 ASIG5V.n6310 2.2505
R44556 ASIG5V.n6433 ASIG5V.n6431 2.2505
R44557 ASIG5V.n9185 ASIG5V.n9184 2.2505
R44558 ASIG5V.n9178 ASIG5V.n9177 2.2505
R44559 ASIG5V.n6545 ASIG5V.n6444 2.2505
R44560 ASIG5V.n6881 ASIG5V.n6587 2.2505
R44561 ASIG5V.n6884 ASIG5V.n6632 2.2505
R44562 ASIG5V.n7239 ASIG5V.n6889 2.2505
R44563 ASIG5V.n8907 ASIG5V.n8906 2.2505
R44564 ASIG5V.n8270 ASIG5V.n8269 2.2505
R44565 ASIG5V.n8267 ASIG5V.n8171 2.2505
R44566 ASIG5V.n8266 ASIG5V.n8217 2.2505
R44567 ASIG5V.n8276 ASIG5V.n8275 2.2505
R44568 ASIG5V.n8883 ASIG5V.n8882 2.2505
R44569 ASIG5V.n12537 ASIG5V.n12536 2.2505
R44570 ASIG5V.n8582 ASIG5V.n3 2.2505
R44571 ASIG5V.n12530 ASIG5V.n12529 2.2505
R44572 ASIG5V.n512 ASIG5V.n508 2.2505
R44573 ASIG5V.n514 ASIG5V.n513 2.2505
R44574 ASIG5V.n515 ASIG5V.n173 2.2505
R44575 ASIG5V.n12313 ASIG5V.n216 2.2505
R44576 ASIG5V.n12312 ASIG5V.n12311 2.2505
R44577 ASIG5V.n528 ASIG5V.n519 2.2505
R44578 ASIG5V.n12291 ASIG5V.n571 2.2505
R44579 ASIG5V.n12290 ASIG5V.n12289 2.2505
R44580 ASIG5V.n876 ASIG5V.n864 2.2505
R44581 ASIG5V.n12278 ASIG5V.n12277 2.2505
R44582 ASIG5V.n1271 ASIG5V.n880 2.2505
R44583 ASIG5V.n12270 ASIG5V.n12269 2.2505
R44584 ASIG5V.n1326 ASIG5V.n1225 2.2505
R44585 ASIG5V.n1664 ASIG5V.n1328 2.2505
R44586 ASIG5V.n1667 ASIG5V.n1370 2.2505
R44587 ASIG5V.n1674 ASIG5V.n1672 2.2505
R44588 ASIG5V.n11999 ASIG5V.n11998 2.2505
R44589 ASIG5V.n1860 ASIG5V.n1721 2.2505
R44590 ASIG5V.n1862 ASIG5V.n1861 2.2505
R44591 ASIG5V.n2201 ASIG5V.n2200 2.2505
R44592 ASIG5V.n1850 ASIG5V.n1848 2.2505
R44593 ASIG5V.n11791 ASIG5V.n11790 2.2505
R44594 ASIG5V.n2556 ASIG5V.n1851 2.2505
R44595 ASIG5V.n11783 ASIG5V.n11782 2.2505
R44596 ASIG5V.n2213 ASIG5V.n2211 2.2505
R44597 ASIG5V.n11761 ASIG5V.n2569 2.2505
R44598 ASIG5V.n11760 ASIG5V.n2612 2.2505
R44599 ASIG5V.n11759 ASIG5V.n2907 2.2505
R44600 ASIG5V.n11753 ASIG5V.n11752 2.2505
R44601 ASIG5V.n9965 ASIG5V.n2912 2.2505
R44602 ASIG5V.n11494 ASIG5V.n11493 2.2505
R44603 ASIG5V.n11487 ASIG5V.n11486 2.2505
R44604 ASIG5V.n10016 ASIG5V.n9972 2.2505
R44605 ASIG5V.n10363 ASIG5V.n10025 2.2505
R44606 ASIG5V.n10366 ASIG5V.n10068 2.2505
R44607 ASIG5V.n10423 ASIG5V.n10371 2.2505
R44608 ASIG5V.n11174 ASIG5V.n11173 2.2505
R44609 ASIG5V.n10484 ASIG5V.n10482 2.2505
R44610 ASIG5V.n10919 ASIG5V.n10918 2.2505
R44611 ASIG5V.n10703 ASIG5V.n10485 2.2505
R44612 ASIG5V.n4309 ASIG5V.n3829 2.2505
R44613 ASIG5V.n4552 ASIG5V.n4551 2.2505
R44614 ASIG5V.n4311 ASIG5V.n4310 2.2505
R44615 ASIG5V.n4547 ASIG5V.n4546 2.2505
R44616 ASIG5V.n4545 ASIG5V.n4544 2.2505
R44617 ASIG5V.n4543 ASIG5V.n4315 2.2505
R44618 ASIG5V.n4314 ASIG5V.n4313 2.2505
R44619 ASIG5V.n4539 ASIG5V.n4538 2.2505
R44620 ASIG5V.n4537 ASIG5V.n4536 2.2505
R44621 ASIG5V.n4535 ASIG5V.n4319 2.2505
R44622 ASIG5V.n4318 ASIG5V.n4317 2.2505
R44623 ASIG5V.n4531 ASIG5V.n4530 2.2505
R44624 ASIG5V.n4529 ASIG5V.n4528 2.2505
R44625 ASIG5V.n4527 ASIG5V.n4323 2.2505
R44626 ASIG5V.n4322 ASIG5V.n4321 2.2505
R44627 ASIG5V.n4523 ASIG5V.n4522 2.2505
R44628 ASIG5V.n4521 ASIG5V.n4520 2.2505
R44629 ASIG5V.n4519 ASIG5V.n4327 2.2505
R44630 ASIG5V.n4326 ASIG5V.n4325 2.2505
R44631 ASIG5V.n4515 ASIG5V.n4514 2.2505
R44632 ASIG5V.n4513 ASIG5V.n4512 2.2505
R44633 ASIG5V.n4511 ASIG5V.n4331 2.2505
R44634 ASIG5V.n4330 ASIG5V.n4329 2.2505
R44635 ASIG5V.n4507 ASIG5V.n4506 2.2505
R44636 ASIG5V.n4505 ASIG5V.n4504 2.2505
R44637 ASIG5V.n4503 ASIG5V.n4335 2.2505
R44638 ASIG5V.n4334 ASIG5V.n4333 2.2505
R44639 ASIG5V.n4499 ASIG5V.n4498 2.2505
R44640 ASIG5V.n4497 ASIG5V.n4496 2.2505
R44641 ASIG5V.n4495 ASIG5V.n4339 2.2505
R44642 ASIG5V.n4338 ASIG5V.n4337 2.2505
R44643 ASIG5V.n4491 ASIG5V.n4490 2.2505
R44644 ASIG5V.n4489 ASIG5V.n4488 2.2505
R44645 ASIG5V.n4487 ASIG5V.n4343 2.2505
R44646 ASIG5V.n4342 ASIG5V.n4341 2.2505
R44647 ASIG5V.n4483 ASIG5V.n4482 2.2505
R44648 ASIG5V.n4481 ASIG5V.n4480 2.2505
R44649 ASIG5V.n4479 ASIG5V.n4347 2.2505
R44650 ASIG5V.n4346 ASIG5V.n4345 2.2505
R44651 ASIG5V.n4475 ASIG5V.n4474 2.2505
R44652 ASIG5V.n4473 ASIG5V.n4472 2.2505
R44653 ASIG5V.n4471 ASIG5V.n4351 2.2505
R44654 ASIG5V.n4350 ASIG5V.n4349 2.2505
R44655 ASIG5V.n4467 ASIG5V.n4466 2.2505
R44656 ASIG5V.n4465 ASIG5V.n4464 2.2505
R44657 ASIG5V.n4463 ASIG5V.n4355 2.2505
R44658 ASIG5V.n4354 ASIG5V.n4353 2.2505
R44659 ASIG5V.n4459 ASIG5V.n4458 2.2505
R44660 ASIG5V.n4457 ASIG5V.n4456 2.2505
R44661 ASIG5V.n4455 ASIG5V.n4359 2.2505
R44662 ASIG5V.n4358 ASIG5V.n4357 2.2505
R44663 ASIG5V.n4451 ASIG5V.n4450 2.2505
R44664 ASIG5V.n4449 ASIG5V.n4448 2.2505
R44665 ASIG5V.n4447 ASIG5V.n4363 2.2505
R44666 ASIG5V.n4362 ASIG5V.n4361 2.2505
R44667 ASIG5V.n4443 ASIG5V.n4442 2.2505
R44668 ASIG5V.n4441 ASIG5V.n4440 2.2505
R44669 ASIG5V.n4439 ASIG5V.n4367 2.2505
R44670 ASIG5V.n4366 ASIG5V.n4365 2.2505
R44671 ASIG5V.n4435 ASIG5V.n4434 2.2505
R44672 ASIG5V.n4433 ASIG5V.n4432 2.2505
R44673 ASIG5V.n4431 ASIG5V.n4371 2.2505
R44674 ASIG5V.n4370 ASIG5V.n4369 2.2505
R44675 ASIG5V.n4427 ASIG5V.n4426 2.2505
R44676 ASIG5V.n4425 ASIG5V.n4424 2.2505
R44677 ASIG5V.n4423 ASIG5V.n4375 2.2505
R44678 ASIG5V.n4374 ASIG5V.n4373 2.2505
R44679 ASIG5V.n4419 ASIG5V.n4418 2.2505
R44680 ASIG5V.n4417 ASIG5V.n4416 2.2505
R44681 ASIG5V.n4415 ASIG5V.n4379 2.2505
R44682 ASIG5V.n4378 ASIG5V.n4377 2.2505
R44683 ASIG5V.n4411 ASIG5V.n4410 2.2505
R44684 ASIG5V.n4409 ASIG5V.n4408 2.2505
R44685 ASIG5V.n4407 ASIG5V.n4383 2.2505
R44686 ASIG5V.n4382 ASIG5V.n4381 2.2505
R44687 ASIG5V.n4403 ASIG5V.n4402 2.2505
R44688 ASIG5V.n4401 ASIG5V.n4400 2.2505
R44689 ASIG5V.n4399 ASIG5V.n4387 2.2505
R44690 ASIG5V.n4386 ASIG5V.n4385 2.2505
R44691 ASIG5V.n4395 ASIG5V.n4394 2.2505
R44692 ASIG5V.n4393 ASIG5V.n4392 2.2505
R44693 ASIG5V.n4391 ASIG5V.n4389 2.2505
R44694 ASIG5V.n3834 ASIG5V.n3833 2.2505
R44695 ASIG5V.n4567 ASIG5V.n4566 2.2505
R44696 ASIG5V.n11181 ASIG5V.n10362 2.2505
R44697 ASIG5V.n10361 ASIG5V.n10072 2.2505
R44698 ASIG5V.n10360 ASIG5V.n10359 2.2505
R44699 ASIG5V.n10074 ASIG5V.n10073 2.2505
R44700 ASIG5V.n10179 ASIG5V.n10178 2.2505
R44701 ASIG5V.n10180 ASIG5V.n10176 2.2505
R44702 ASIG5V.n10183 ASIG5V.n10181 2.2505
R44703 ASIG5V.n10185 ASIG5V.n10174 2.2505
R44704 ASIG5V.n10188 ASIG5V.n10187 2.2505
R44705 ASIG5V.n10189 ASIG5V.n10173 2.2505
R44706 ASIG5V.n10192 ASIG5V.n10190 2.2505
R44707 ASIG5V.n10194 ASIG5V.n10171 2.2505
R44708 ASIG5V.n10197 ASIG5V.n10196 2.2505
R44709 ASIG5V.n10198 ASIG5V.n10170 2.2505
R44710 ASIG5V.n10201 ASIG5V.n10199 2.2505
R44711 ASIG5V.n10203 ASIG5V.n10168 2.2505
R44712 ASIG5V.n10206 ASIG5V.n10205 2.2505
R44713 ASIG5V.n10207 ASIG5V.n10167 2.2505
R44714 ASIG5V.n10210 ASIG5V.n10208 2.2505
R44715 ASIG5V.n10212 ASIG5V.n10165 2.2505
R44716 ASIG5V.n10215 ASIG5V.n10214 2.2505
R44717 ASIG5V.n10216 ASIG5V.n10164 2.2505
R44718 ASIG5V.n10219 ASIG5V.n10217 2.2505
R44719 ASIG5V.n10221 ASIG5V.n10162 2.2505
R44720 ASIG5V.n10224 ASIG5V.n10223 2.2505
R44721 ASIG5V.n10225 ASIG5V.n10161 2.2505
R44722 ASIG5V.n10228 ASIG5V.n10226 2.2505
R44723 ASIG5V.n10230 ASIG5V.n10159 2.2505
R44724 ASIG5V.n10233 ASIG5V.n10232 2.2505
R44725 ASIG5V.n10234 ASIG5V.n10158 2.2505
R44726 ASIG5V.n10237 ASIG5V.n10235 2.2505
R44727 ASIG5V.n10239 ASIG5V.n10156 2.2505
R44728 ASIG5V.n10242 ASIG5V.n10241 2.2505
R44729 ASIG5V.n10243 ASIG5V.n10155 2.2505
R44730 ASIG5V.n10246 ASIG5V.n10244 2.2505
R44731 ASIG5V.n10248 ASIG5V.n10153 2.2505
R44732 ASIG5V.n10251 ASIG5V.n10250 2.2505
R44733 ASIG5V.n10252 ASIG5V.n10152 2.2505
R44734 ASIG5V.n10255 ASIG5V.n10253 2.2505
R44735 ASIG5V.n10257 ASIG5V.n10150 2.2505
R44736 ASIG5V.n10260 ASIG5V.n10259 2.2505
R44737 ASIG5V.n10261 ASIG5V.n10149 2.2505
R44738 ASIG5V.n10264 ASIG5V.n10262 2.2505
R44739 ASIG5V.n10266 ASIG5V.n10147 2.2505
R44740 ASIG5V.n10269 ASIG5V.n10268 2.2505
R44741 ASIG5V.n10270 ASIG5V.n10146 2.2505
R44742 ASIG5V.n10273 ASIG5V.n10271 2.2505
R44743 ASIG5V.n10275 ASIG5V.n10144 2.2505
R44744 ASIG5V.n10278 ASIG5V.n10277 2.2505
R44745 ASIG5V.n10279 ASIG5V.n10143 2.2505
R44746 ASIG5V.n10282 ASIG5V.n10280 2.2505
R44747 ASIG5V.n10284 ASIG5V.n10141 2.2505
R44748 ASIG5V.n10287 ASIG5V.n10286 2.2505
R44749 ASIG5V.n10288 ASIG5V.n10140 2.2505
R44750 ASIG5V.n10291 ASIG5V.n10289 2.2505
R44751 ASIG5V.n10293 ASIG5V.n10138 2.2505
R44752 ASIG5V.n10296 ASIG5V.n10295 2.2505
R44753 ASIG5V.n10297 ASIG5V.n10137 2.2505
R44754 ASIG5V.n10300 ASIG5V.n10298 2.2505
R44755 ASIG5V.n10302 ASIG5V.n10135 2.2505
R44756 ASIG5V.n10305 ASIG5V.n10304 2.2505
R44757 ASIG5V.n10306 ASIG5V.n10134 2.2505
R44758 ASIG5V.n10309 ASIG5V.n10307 2.2505
R44759 ASIG5V.n10311 ASIG5V.n10132 2.2505
R44760 ASIG5V.n10314 ASIG5V.n10313 2.2505
R44761 ASIG5V.n10315 ASIG5V.n10131 2.2505
R44762 ASIG5V.n10318 ASIG5V.n10316 2.2505
R44763 ASIG5V.n10320 ASIG5V.n10129 2.2505
R44764 ASIG5V.n10323 ASIG5V.n10322 2.2505
R44765 ASIG5V.n10324 ASIG5V.n10128 2.2505
R44766 ASIG5V.n10327 ASIG5V.n10325 2.2505
R44767 ASIG5V.n10329 ASIG5V.n10126 2.2505
R44768 ASIG5V.n10332 ASIG5V.n10331 2.2505
R44769 ASIG5V.n10333 ASIG5V.n10125 2.2505
R44770 ASIG5V.n10336 ASIG5V.n10334 2.2505
R44771 ASIG5V.n10338 ASIG5V.n10123 2.2505
R44772 ASIG5V.n10341 ASIG5V.n10340 2.2505
R44773 ASIG5V.n10342 ASIG5V.n10122 2.2505
R44774 ASIG5V.n10345 ASIG5V.n10343 2.2505
R44775 ASIG5V.n10347 ASIG5V.n10120 2.2505
R44776 ASIG5V.n10350 ASIG5V.n10349 2.2505
R44777 ASIG5V.n10351 ASIG5V.n10118 2.2505
R44778 ASIG5V.n10353 ASIG5V.n10352 2.2505
R44779 ASIG5V.n10119 ASIG5V.n10116 2.2505
R44780 ASIG5V.n10116 ASIG5V.n10067 2.2505
R44781 ASIG5V.n10354 ASIG5V.n10353 2.2505
R44782 ASIG5V.n10118 ASIG5V.n10117 2.2505
R44783 ASIG5V.n10349 ASIG5V.n10348 2.2505
R44784 ASIG5V.n10347 ASIG5V.n10346 2.2505
R44785 ASIG5V.n10345 ASIG5V.n10344 2.2505
R44786 ASIG5V.n10122 ASIG5V.n10121 2.2505
R44787 ASIG5V.n10340 ASIG5V.n10339 2.2505
R44788 ASIG5V.n10338 ASIG5V.n10337 2.2505
R44789 ASIG5V.n10336 ASIG5V.n10335 2.2505
R44790 ASIG5V.n10125 ASIG5V.n10124 2.2505
R44791 ASIG5V.n10331 ASIG5V.n10330 2.2505
R44792 ASIG5V.n10329 ASIG5V.n10328 2.2505
R44793 ASIG5V.n10327 ASIG5V.n10326 2.2505
R44794 ASIG5V.n10128 ASIG5V.n10127 2.2505
R44795 ASIG5V.n10322 ASIG5V.n10321 2.2505
R44796 ASIG5V.n10320 ASIG5V.n10319 2.2505
R44797 ASIG5V.n10318 ASIG5V.n10317 2.2505
R44798 ASIG5V.n10131 ASIG5V.n10130 2.2505
R44799 ASIG5V.n10313 ASIG5V.n10312 2.2505
R44800 ASIG5V.n10311 ASIG5V.n10310 2.2505
R44801 ASIG5V.n10309 ASIG5V.n10308 2.2505
R44802 ASIG5V.n10134 ASIG5V.n10133 2.2505
R44803 ASIG5V.n10304 ASIG5V.n10303 2.2505
R44804 ASIG5V.n10302 ASIG5V.n10301 2.2505
R44805 ASIG5V.n10300 ASIG5V.n10299 2.2505
R44806 ASIG5V.n10137 ASIG5V.n10136 2.2505
R44807 ASIG5V.n10295 ASIG5V.n10294 2.2505
R44808 ASIG5V.n10293 ASIG5V.n10292 2.2505
R44809 ASIG5V.n10291 ASIG5V.n10290 2.2505
R44810 ASIG5V.n10140 ASIG5V.n10139 2.2505
R44811 ASIG5V.n10286 ASIG5V.n10285 2.2505
R44812 ASIG5V.n10284 ASIG5V.n10283 2.2505
R44813 ASIG5V.n10282 ASIG5V.n10281 2.2505
R44814 ASIG5V.n10143 ASIG5V.n10142 2.2505
R44815 ASIG5V.n10277 ASIG5V.n10276 2.2505
R44816 ASIG5V.n10275 ASIG5V.n10274 2.2505
R44817 ASIG5V.n10273 ASIG5V.n10272 2.2505
R44818 ASIG5V.n10146 ASIG5V.n10145 2.2505
R44819 ASIG5V.n10268 ASIG5V.n10267 2.2505
R44820 ASIG5V.n10266 ASIG5V.n10265 2.2505
R44821 ASIG5V.n10264 ASIG5V.n10263 2.2505
R44822 ASIG5V.n10149 ASIG5V.n10148 2.2505
R44823 ASIG5V.n10259 ASIG5V.n10258 2.2505
R44824 ASIG5V.n10257 ASIG5V.n10256 2.2505
R44825 ASIG5V.n10255 ASIG5V.n10254 2.2505
R44826 ASIG5V.n10152 ASIG5V.n10151 2.2505
R44827 ASIG5V.n10250 ASIG5V.n10249 2.2505
R44828 ASIG5V.n10248 ASIG5V.n10247 2.2505
R44829 ASIG5V.n10246 ASIG5V.n10245 2.2505
R44830 ASIG5V.n10155 ASIG5V.n10154 2.2505
R44831 ASIG5V.n10241 ASIG5V.n10240 2.2505
R44832 ASIG5V.n10239 ASIG5V.n10238 2.2505
R44833 ASIG5V.n10237 ASIG5V.n10236 2.2505
R44834 ASIG5V.n10158 ASIG5V.n10157 2.2505
R44835 ASIG5V.n10232 ASIG5V.n10231 2.2505
R44836 ASIG5V.n10230 ASIG5V.n10229 2.2505
R44837 ASIG5V.n10228 ASIG5V.n10227 2.2505
R44838 ASIG5V.n10161 ASIG5V.n10160 2.2505
R44839 ASIG5V.n10223 ASIG5V.n10222 2.2505
R44840 ASIG5V.n10221 ASIG5V.n10220 2.2505
R44841 ASIG5V.n10219 ASIG5V.n10218 2.2505
R44842 ASIG5V.n10164 ASIG5V.n10163 2.2505
R44843 ASIG5V.n10214 ASIG5V.n10213 2.2505
R44844 ASIG5V.n10212 ASIG5V.n10211 2.2505
R44845 ASIG5V.n10210 ASIG5V.n10209 2.2505
R44846 ASIG5V.n10167 ASIG5V.n10166 2.2505
R44847 ASIG5V.n10205 ASIG5V.n10204 2.2505
R44848 ASIG5V.n10203 ASIG5V.n10202 2.2505
R44849 ASIG5V.n10201 ASIG5V.n10200 2.2505
R44850 ASIG5V.n10170 ASIG5V.n10169 2.2505
R44851 ASIG5V.n10196 ASIG5V.n10195 2.2505
R44852 ASIG5V.n10194 ASIG5V.n10193 2.2505
R44853 ASIG5V.n10192 ASIG5V.n10191 2.2505
R44854 ASIG5V.n10173 ASIG5V.n10172 2.2505
R44855 ASIG5V.n10187 ASIG5V.n10186 2.2505
R44856 ASIG5V.n10185 ASIG5V.n10184 2.2505
R44857 ASIG5V.n10183 ASIG5V.n10182 2.2505
R44858 ASIG5V.n10176 ASIG5V.n10175 2.2505
R44859 ASIG5V.n10178 ASIG5V.n10177 2.2505
R44860 ASIG5V.n10075 ASIG5V.n10074 2.2505
R44861 ASIG5V.n10359 ASIG5V.n10358 2.2505
R44862 ASIG5V.n10072 ASIG5V.n10071 2.2505
R44863 ASIG5V.n11182 ASIG5V.n11181 2.2505
R44864 ASIG5V.n4250 ASIG5V.n3839 2.2505
R44865 ASIG5V.n4557 ASIG5V.n3838 2.2505
R44866 ASIG5V.n4559 ASIG5V.n4558 2.2505
R44867 ASIG5V.n4562 ASIG5V.n4561 2.2505
R44868 ASIG5V.n3627 ASIG5V.n3625 2.2505
R44869 ASIG5V.n4779 ASIG5V.n4778 2.2505
R44870 ASIG5V.n3622 ASIG5V.n3621 2.2505
R44871 ASIG5V.n4785 ASIG5V.n4784 2.2505
R44872 ASIG5V.n4801 ASIG5V.n4800 2.2505
R44873 ASIG5V.n3272 ASIG5V.n3271 2.2505
R44874 ASIG5V.n4806 ASIG5V.n4805 2.2505
R44875 ASIG5V.n5067 ASIG5V.n5066 2.2505
R44876 ASIG5V.n3173 ASIG5V.n3171 2.2505
R44877 ASIG5V.n9742 ASIG5V.n9741 2.2505
R44878 ASIG5V.n9737 ASIG5V.n9736 2.2505
R44879 ASIG5V.n5073 ASIG5V.n5072 2.2505
R44880 ASIG5V.n5460 ASIG5V.n5459 2.2505
R44881 ASIG5V.n9423 ASIG5V.n9422 2.2505
R44882 ASIG5V.n9421 ASIG5V.n5462 2.2505
R44883 ASIG5V.n5558 ASIG5V.n5463 2.2505
R44884 ASIG5V.n9412 ASIG5V.n5560 2.2505
R44885 ASIG5V.n5565 ASIG5V.n5559 2.2505
R44886 ASIG5V.n9408 ASIG5V.n9407 2.2505
R44887 ASIG5V.n6255 ASIG5V.n6254 2.2505
R44888 ASIG5V.n6251 ASIG5V.n6248 2.2505
R44889 ASIG5V.n9389 ASIG5V.n6250 2.2505
R44890 ASIG5V.n6261 ASIG5V.n6249 2.2505
R44891 ASIG5V.n9385 ASIG5V.n9384 2.2505
R44892 ASIG5V.n6438 ASIG5V.n6437 2.2505
R44893 ASIG5V.n6435 ASIG5V.n6433 2.2505
R44894 ASIG5V.n9184 ASIG5V.n9183 2.2505
R44895 ASIG5V.n9179 ASIG5V.n9178 2.2505
R44896 ASIG5V.n6444 ASIG5V.n6443 2.2505
R44897 ASIG5V.n6882 ASIG5V.n6881 2.2505
R44898 ASIG5V.n8912 ASIG5V.n6884 2.2505
R44899 ASIG5V.n6889 ASIG5V.n6883 2.2505
R44900 ASIG5V.n8908 ASIG5V.n8907 2.2505
R44901 ASIG5V.n8271 ASIG5V.n8270 2.2505
R44902 ASIG5V.n8267 ASIG5V.n8264 2.2505
R44903 ASIG5V.n8888 ASIG5V.n8266 2.2505
R44904 ASIG5V.n8275 ASIG5V.n8265 2.2505
R44905 ASIG5V.n8884 ASIG5V.n8883 2.2505
R44906 ASIG5V.n12536 ASIG5V.n12535 2.2505
R44907 ASIG5V.n5 ASIG5V.n3 2.2505
R44908 ASIG5V.n12531 ASIG5V.n12530 2.2505
R44909 ASIG5V.n512 ASIG5V.n511 2.2505
R44910 ASIG5V.n514 ASIG5V.n507 2.2505
R44911 ASIG5V.n516 ASIG5V.n515 2.2505
R44912 ASIG5V.n12314 ASIG5V.n12313 2.2505
R44913 ASIG5V.n12312 ASIG5V.n518 2.2505
R44914 ASIG5V.n861 ASIG5V.n519 2.2505
R44915 ASIG5V.n12292 ASIG5V.n12291 2.2505
R44916 ASIG5V.n12290 ASIG5V.n863 2.2505
R44917 ASIG5V.n1217 ASIG5V.n864 2.2505
R44918 ASIG5V.n12277 ASIG5V.n12276 2.2505
R44919 ASIG5V.n882 ASIG5V.n880 2.2505
R44920 ASIG5V.n12271 ASIG5V.n12270 2.2505
R44921 ASIG5V.n1225 ASIG5V.n1223 2.2505
R44922 ASIG5V.n1665 ASIG5V.n1664 2.2505
R44923 ASIG5V.n12004 ASIG5V.n1667 2.2505
R44924 ASIG5V.n1672 ASIG5V.n1666 2.2505
R44925 ASIG5V.n12000 ASIG5V.n11999 2.2505
R44926 ASIG5V.n1860 ASIG5V.n1859 2.2505
R44927 ASIG5V.n1862 ASIG5V.n1856 2.2505
R44928 ASIG5V.n2202 ASIG5V.n2201 2.2505
R44929 ASIG5V.n1852 ASIG5V.n1850 2.2505
R44930 ASIG5V.n11790 ASIG5V.n11789 2.2505
R44931 ASIG5V.n1853 ASIG5V.n1851 2.2505
R44932 ASIG5V.n11784 ASIG5V.n11783 2.2505
R44933 ASIG5V.n2211 ASIG5V.n2209 2.2505
R44934 ASIG5V.n11762 ASIG5V.n11761 2.2505
R44935 ASIG5V.n11760 ASIG5V.n2904 2.2505
R44936 ASIG5V.n11759 ASIG5V.n11758 2.2505
R44937 ASIG5V.n11754 ASIG5V.n11753 2.2505
R44938 ASIG5V.n2912 ASIG5V.n2911 2.2505
R44939 ASIG5V.n11493 ASIG5V.n11492 2.2505
R44940 ASIG5V.n11488 ASIG5V.n11487 2.2505
R44941 ASIG5V.n9972 ASIG5V.n9971 2.2505
R44942 ASIG5V.n10364 ASIG5V.n10363 2.2505
R44943 ASIG5V.n11179 ASIG5V.n10366 2.2505
R44944 ASIG5V.n10371 ASIG5V.n10365 2.2505
R44945 ASIG5V.n11175 ASIG5V.n11174 2.2505
R44946 ASIG5V.n10486 ASIG5V.n10484 2.2505
R44947 ASIG5V.n10918 ASIG5V.n10917 2.2505
R44948 ASIG5V.n10487 ASIG5V.n10485 2.2505
R44949 ASIG5V.n10463 ASIG5V.n10415 2.2505
R44950 ASIG5V.n11161 ASIG5V.n11160 2.2505
R44951 ASIG5V.n10465 ASIG5V.n10464 2.2505
R44952 ASIG5V.n11156 ASIG5V.n11155 2.2505
R44953 ASIG5V.n11154 ASIG5V.n11153 2.2505
R44954 ASIG5V.n11152 ASIG5V.n10930 2.2505
R44955 ASIG5V.n10929 ASIG5V.n10928 2.2505
R44956 ASIG5V.n11148 ASIG5V.n11147 2.2505
R44957 ASIG5V.n11146 ASIG5V.n11145 2.2505
R44958 ASIG5V.n11144 ASIG5V.n10934 2.2505
R44959 ASIG5V.n10933 ASIG5V.n10932 2.2505
R44960 ASIG5V.n11140 ASIG5V.n11139 2.2505
R44961 ASIG5V.n11138 ASIG5V.n11137 2.2505
R44962 ASIG5V.n11136 ASIG5V.n10938 2.2505
R44963 ASIG5V.n10937 ASIG5V.n10936 2.2505
R44964 ASIG5V.n11132 ASIG5V.n11131 2.2505
R44965 ASIG5V.n11130 ASIG5V.n11129 2.2505
R44966 ASIG5V.n11128 ASIG5V.n10942 2.2505
R44967 ASIG5V.n10941 ASIG5V.n10940 2.2505
R44968 ASIG5V.n11124 ASIG5V.n11123 2.2505
R44969 ASIG5V.n11122 ASIG5V.n11121 2.2505
R44970 ASIG5V.n11120 ASIG5V.n10946 2.2505
R44971 ASIG5V.n10945 ASIG5V.n10944 2.2505
R44972 ASIG5V.n11116 ASIG5V.n11115 2.2505
R44973 ASIG5V.n11114 ASIG5V.n11113 2.2505
R44974 ASIG5V.n11112 ASIG5V.n10950 2.2505
R44975 ASIG5V.n10949 ASIG5V.n10948 2.2505
R44976 ASIG5V.n11108 ASIG5V.n11107 2.2505
R44977 ASIG5V.n11106 ASIG5V.n11105 2.2505
R44978 ASIG5V.n11104 ASIG5V.n10954 2.2505
R44979 ASIG5V.n10953 ASIG5V.n10952 2.2505
R44980 ASIG5V.n11100 ASIG5V.n11099 2.2505
R44981 ASIG5V.n11098 ASIG5V.n11097 2.2505
R44982 ASIG5V.n11096 ASIG5V.n10958 2.2505
R44983 ASIG5V.n10957 ASIG5V.n10956 2.2505
R44984 ASIG5V.n11092 ASIG5V.n11091 2.2505
R44985 ASIG5V.n11090 ASIG5V.n11089 2.2505
R44986 ASIG5V.n11088 ASIG5V.n10962 2.2505
R44987 ASIG5V.n10961 ASIG5V.n10960 2.2505
R44988 ASIG5V.n11084 ASIG5V.n11083 2.2505
R44989 ASIG5V.n11082 ASIG5V.n11081 2.2505
R44990 ASIG5V.n11080 ASIG5V.n10966 2.2505
R44991 ASIG5V.n10965 ASIG5V.n10964 2.2505
R44992 ASIG5V.n11076 ASIG5V.n11075 2.2505
R44993 ASIG5V.n11074 ASIG5V.n11073 2.2505
R44994 ASIG5V.n11072 ASIG5V.n10970 2.2505
R44995 ASIG5V.n10969 ASIG5V.n10968 2.2505
R44996 ASIG5V.n11068 ASIG5V.n11067 2.2505
R44997 ASIG5V.n11066 ASIG5V.n11065 2.2505
R44998 ASIG5V.n11064 ASIG5V.n10974 2.2505
R44999 ASIG5V.n10973 ASIG5V.n10972 2.2505
R45000 ASIG5V.n11060 ASIG5V.n11059 2.2505
R45001 ASIG5V.n11058 ASIG5V.n11057 2.2505
R45002 ASIG5V.n11056 ASIG5V.n10978 2.2505
R45003 ASIG5V.n10977 ASIG5V.n10976 2.2505
R45004 ASIG5V.n11052 ASIG5V.n11051 2.2505
R45005 ASIG5V.n11050 ASIG5V.n11049 2.2505
R45006 ASIG5V.n11048 ASIG5V.n10982 2.2505
R45007 ASIG5V.n10981 ASIG5V.n10980 2.2505
R45008 ASIG5V.n11044 ASIG5V.n11043 2.2505
R45009 ASIG5V.n11042 ASIG5V.n11041 2.2505
R45010 ASIG5V.n11040 ASIG5V.n10986 2.2505
R45011 ASIG5V.n10985 ASIG5V.n10984 2.2505
R45012 ASIG5V.n11036 ASIG5V.n11035 2.2505
R45013 ASIG5V.n11034 ASIG5V.n11033 2.2505
R45014 ASIG5V.n11032 ASIG5V.n10990 2.2505
R45015 ASIG5V.n10989 ASIG5V.n10988 2.2505
R45016 ASIG5V.n11028 ASIG5V.n11027 2.2505
R45017 ASIG5V.n11026 ASIG5V.n11025 2.2505
R45018 ASIG5V.n11024 ASIG5V.n10994 2.2505
R45019 ASIG5V.n10993 ASIG5V.n10992 2.2505
R45020 ASIG5V.n11020 ASIG5V.n11019 2.2505
R45021 ASIG5V.n11018 ASIG5V.n11017 2.2505
R45022 ASIG5V.n11016 ASIG5V.n10998 2.2505
R45023 ASIG5V.n10997 ASIG5V.n10996 2.2505
R45024 ASIG5V.n11012 ASIG5V.n11011 2.2505
R45025 ASIG5V.n11010 ASIG5V.n11009 2.2505
R45026 ASIG5V.n11008 ASIG5V.n11002 2.2505
R45027 ASIG5V.n11001 ASIG5V.n11000 2.2505
R45028 ASIG5V.n11004 ASIG5V.n11003 2.2505
R45029 ASIG5V.n10422 ASIG5V.n10421 2.2505
R45030 ASIG5V.n11166 ASIG5V.n11165 2.2505
R45031 ASIG5V.n10419 ASIG5V.n10418 2.2505
R45032 ASIG5V.n11171 ASIG5V.n11170 2.2505
R45033 ASIG5V.n11170 ASIG5V.n11169 2.2505
R45034 ASIG5V.n11168 ASIG5V.n10419 2.2505
R45035 ASIG5V.n11167 ASIG5V.n11166 2.2505
R45036 ASIG5V.n10421 ASIG5V.n10420 2.2505
R45037 ASIG5V.n11005 ASIG5V.n11004 2.2505
R45038 ASIG5V.n11006 ASIG5V.n11001 2.2505
R45039 ASIG5V.n11008 ASIG5V.n11007 2.2505
R45040 ASIG5V.n11010 ASIG5V.n10999 2.2505
R45041 ASIG5V.n11013 ASIG5V.n11012 2.2505
R45042 ASIG5V.n11014 ASIG5V.n10997 2.2505
R45043 ASIG5V.n11016 ASIG5V.n11015 2.2505
R45044 ASIG5V.n11018 ASIG5V.n10995 2.2505
R45045 ASIG5V.n11021 ASIG5V.n11020 2.2505
R45046 ASIG5V.n11022 ASIG5V.n10993 2.2505
R45047 ASIG5V.n11024 ASIG5V.n11023 2.2505
R45048 ASIG5V.n11026 ASIG5V.n10991 2.2505
R45049 ASIG5V.n11029 ASIG5V.n11028 2.2505
R45050 ASIG5V.n11030 ASIG5V.n10989 2.2505
R45051 ASIG5V.n11032 ASIG5V.n11031 2.2505
R45052 ASIG5V.n11034 ASIG5V.n10987 2.2505
R45053 ASIG5V.n11037 ASIG5V.n11036 2.2505
R45054 ASIG5V.n11038 ASIG5V.n10985 2.2505
R45055 ASIG5V.n11040 ASIG5V.n11039 2.2505
R45056 ASIG5V.n11042 ASIG5V.n10983 2.2505
R45057 ASIG5V.n11045 ASIG5V.n11044 2.2505
R45058 ASIG5V.n11046 ASIG5V.n10981 2.2505
R45059 ASIG5V.n11048 ASIG5V.n11047 2.2505
R45060 ASIG5V.n11050 ASIG5V.n10979 2.2505
R45061 ASIG5V.n11053 ASIG5V.n11052 2.2505
R45062 ASIG5V.n11054 ASIG5V.n10977 2.2505
R45063 ASIG5V.n11056 ASIG5V.n11055 2.2505
R45064 ASIG5V.n11058 ASIG5V.n10975 2.2505
R45065 ASIG5V.n11061 ASIG5V.n11060 2.2505
R45066 ASIG5V.n11062 ASIG5V.n10973 2.2505
R45067 ASIG5V.n11064 ASIG5V.n11063 2.2505
R45068 ASIG5V.n11066 ASIG5V.n10971 2.2505
R45069 ASIG5V.n11069 ASIG5V.n11068 2.2505
R45070 ASIG5V.n11070 ASIG5V.n10969 2.2505
R45071 ASIG5V.n11072 ASIG5V.n11071 2.2505
R45072 ASIG5V.n11074 ASIG5V.n10967 2.2505
R45073 ASIG5V.n11077 ASIG5V.n11076 2.2505
R45074 ASIG5V.n11078 ASIG5V.n10965 2.2505
R45075 ASIG5V.n11080 ASIG5V.n11079 2.2505
R45076 ASIG5V.n11082 ASIG5V.n10963 2.2505
R45077 ASIG5V.n11085 ASIG5V.n11084 2.2505
R45078 ASIG5V.n11086 ASIG5V.n10961 2.2505
R45079 ASIG5V.n11088 ASIG5V.n11087 2.2505
R45080 ASIG5V.n11090 ASIG5V.n10959 2.2505
R45081 ASIG5V.n11093 ASIG5V.n11092 2.2505
R45082 ASIG5V.n11094 ASIG5V.n10957 2.2505
R45083 ASIG5V.n11096 ASIG5V.n11095 2.2505
R45084 ASIG5V.n11098 ASIG5V.n10955 2.2505
R45085 ASIG5V.n11101 ASIG5V.n11100 2.2505
R45086 ASIG5V.n11102 ASIG5V.n10953 2.2505
R45087 ASIG5V.n11104 ASIG5V.n11103 2.2505
R45088 ASIG5V.n11106 ASIG5V.n10951 2.2505
R45089 ASIG5V.n11109 ASIG5V.n11108 2.2505
R45090 ASIG5V.n11110 ASIG5V.n10949 2.2505
R45091 ASIG5V.n11112 ASIG5V.n11111 2.2505
R45092 ASIG5V.n11114 ASIG5V.n10947 2.2505
R45093 ASIG5V.n11117 ASIG5V.n11116 2.2505
R45094 ASIG5V.n11118 ASIG5V.n10945 2.2505
R45095 ASIG5V.n11120 ASIG5V.n11119 2.2505
R45096 ASIG5V.n11122 ASIG5V.n10943 2.2505
R45097 ASIG5V.n11125 ASIG5V.n11124 2.2505
R45098 ASIG5V.n11126 ASIG5V.n10941 2.2505
R45099 ASIG5V.n11128 ASIG5V.n11127 2.2505
R45100 ASIG5V.n11130 ASIG5V.n10939 2.2505
R45101 ASIG5V.n11133 ASIG5V.n11132 2.2505
R45102 ASIG5V.n11134 ASIG5V.n10937 2.2505
R45103 ASIG5V.n11136 ASIG5V.n11135 2.2505
R45104 ASIG5V.n11138 ASIG5V.n10935 2.2505
R45105 ASIG5V.n11141 ASIG5V.n11140 2.2505
R45106 ASIG5V.n11142 ASIG5V.n10933 2.2505
R45107 ASIG5V.n11144 ASIG5V.n11143 2.2505
R45108 ASIG5V.n11146 ASIG5V.n10931 2.2505
R45109 ASIG5V.n11149 ASIG5V.n11148 2.2505
R45110 ASIG5V.n11150 ASIG5V.n10929 2.2505
R45111 ASIG5V.n11152 ASIG5V.n11151 2.2505
R45112 ASIG5V.n11154 ASIG5V.n10927 2.2505
R45113 ASIG5V.n11157 ASIG5V.n11156 2.2505
R45114 ASIG5V.n11158 ASIG5V.n10465 2.2505
R45115 ASIG5V.n11160 ASIG5V.n11159 2.2505
R45116 ASIG5V.n10926 ASIG5V.n10463 2.2505
R45117 ASIG5V.n4250 ASIG5V.n4249 2.2505
R45118 ASIG5V.n3838 ASIG5V.n3837 2.2505
R45119 ASIG5V.n4560 ASIG5V.n4559 2.2505
R45120 ASIG5V.n4563 ASIG5V.n4562 2.2505
R45121 ASIG5V.n3625 ASIG5V.n3624 2.2505
R45122 ASIG5V.n4780 ASIG5V.n4779 2.2505
R45123 ASIG5V.n4782 ASIG5V.n3622 2.2505
R45124 ASIG5V.n4784 ASIG5V.n4783 2.2505
R45125 ASIG5V.n4802 ASIG5V.n4801 2.2505
R45126 ASIG5V.n4803 ASIG5V.n3272 2.2505
R45127 ASIG5V.n4805 ASIG5V.n4804 2.2505
R45128 ASIG5V.n5068 ASIG5V.n5067 2.2505
R45129 ASIG5V.n5069 ASIG5V.n3173 2.2505
R45130 ASIG5V.n9741 ASIG5V.n9740 2.2505
R45131 ASIG5V.n9738 ASIG5V.n9737 2.2505
R45132 ASIG5V.n5072 ASIG5V.n5071 2.2505
R45133 ASIG5V.n5460 ASIG5V.n5457 2.2505
R45134 ASIG5V.n9424 ASIG5V.n9423 2.2505
R45135 ASIG5V.n5462 ASIG5V.n5458 2.2505
R45136 ASIG5V.n5561 ASIG5V.n5558 2.2505
R45137 ASIG5V.n9412 ASIG5V.n9411 2.2505
R45138 ASIG5V.n9410 ASIG5V.n5559 2.2505
R45139 ASIG5V.n9409 ASIG5V.n9408 2.2505
R45140 ASIG5V.n6256 ASIG5V.n6255 2.2505
R45141 ASIG5V.n6257 ASIG5V.n6248 2.2505
R45142 ASIG5V.n9389 ASIG5V.n9388 2.2505
R45143 ASIG5V.n9387 ASIG5V.n6249 2.2505
R45144 ASIG5V.n9386 ASIG5V.n9385 2.2505
R45145 ASIG5V.n6439 ASIG5V.n6438 2.2505
R45146 ASIG5V.n6440 ASIG5V.n6435 2.2505
R45147 ASIG5V.n9183 ASIG5V.n9182 2.2505
R45148 ASIG5V.n9180 ASIG5V.n9179 2.2505
R45149 ASIG5V.n6443 ASIG5V.n6442 2.2505
R45150 ASIG5V.n6885 ASIG5V.n6882 2.2505
R45151 ASIG5V.n8912 ASIG5V.n8911 2.2505
R45152 ASIG5V.n8910 ASIG5V.n6883 2.2505
R45153 ASIG5V.n8909 ASIG5V.n8908 2.2505
R45154 ASIG5V.n8272 ASIG5V.n8271 2.2505
R45155 ASIG5V.n8273 ASIG5V.n8264 2.2505
R45156 ASIG5V.n8888 ASIG5V.n8887 2.2505
R45157 ASIG5V.n8886 ASIG5V.n8265 2.2505
R45158 ASIG5V.n8885 ASIG5V.n8884 2.2505
R45159 ASIG5V.n12535 ASIG5V.n12534 2.2505
R45160 ASIG5V.n12533 ASIG5V.n5 2.2505
R45161 ASIG5V.n12532 ASIG5V.n12531 2.2505
R45162 ASIG5V.n511 ASIG5V.n510 2.2505
R45163 ASIG5V.n509 ASIG5V.n507 2.2505
R45164 ASIG5V.n516 ASIG5V.n505 2.2505
R45165 ASIG5V.n12315 ASIG5V.n12314 2.2505
R45166 ASIG5V.n518 ASIG5V.n506 2.2505
R45167 ASIG5V.n861 ASIG5V.n859 2.2505
R45168 ASIG5V.n12293 ASIG5V.n12292 2.2505
R45169 ASIG5V.n863 ASIG5V.n860 2.2505
R45170 ASIG5V.n1218 ASIG5V.n1217 2.2505
R45171 ASIG5V.n12276 ASIG5V.n12275 2.2505
R45172 ASIG5V.n12274 ASIG5V.n882 2.2505
R45173 ASIG5V.n12272 ASIG5V.n12271 2.2505
R45174 ASIG5V.n1223 ASIG5V.n1221 2.2505
R45175 ASIG5V.n1668 ASIG5V.n1665 2.2505
R45176 ASIG5V.n12004 ASIG5V.n12003 2.2505
R45177 ASIG5V.n12002 ASIG5V.n1666 2.2505
R45178 ASIG5V.n12001 ASIG5V.n12000 2.2505
R45179 ASIG5V.n1859 ASIG5V.n1858 2.2505
R45180 ASIG5V.n1856 ASIG5V.n1855 2.2505
R45181 ASIG5V.n2203 ASIG5V.n2202 2.2505
R45182 ASIG5V.n2205 ASIG5V.n1852 2.2505
R45183 ASIG5V.n11789 ASIG5V.n11788 2.2505
R45184 ASIG5V.n11787 ASIG5V.n1853 2.2505
R45185 ASIG5V.n11785 ASIG5V.n11784 2.2505
R45186 ASIG5V.n2209 ASIG5V.n2207 2.2505
R45187 ASIG5V.n11763 ASIG5V.n11762 2.2505
R45188 ASIG5V.n2904 ASIG5V.n2902 2.2505
R45189 ASIG5V.n11758 ASIG5V.n11757 2.2505
R45190 ASIG5V.n11755 ASIG5V.n11754 2.2505
R45191 ASIG5V.n2911 ASIG5V.n2910 2.2505
R45192 ASIG5V.n11492 ASIG5V.n11491 2.2505
R45193 ASIG5V.n11489 ASIG5V.n11488 2.2505
R45194 ASIG5V.n9971 ASIG5V.n9970 2.2505
R45195 ASIG5V.n10367 ASIG5V.n10364 2.2505
R45196 ASIG5V.n11179 ASIG5V.n11178 2.2505
R45197 ASIG5V.n11177 ASIG5V.n10365 2.2505
R45198 ASIG5V.n11176 ASIG5V.n11175 2.2505
R45199 ASIG5V.n10488 ASIG5V.n10486 2.2505
R45200 ASIG5V.n10917 ASIG5V.n10916 2.2505
R45201 ASIG5V.n10915 ASIG5V.n10487 2.2505
R45202 ASIG5V.n4566 ASIG5V.n4565 2.2505
R45203 ASIG5V.n3836 ASIG5V.n3834 2.2505
R45204 ASIG5V.n4391 ASIG5V.n4390 2.2505
R45205 ASIG5V.n4393 ASIG5V.n4388 2.2505
R45206 ASIG5V.n4396 ASIG5V.n4395 2.2505
R45207 ASIG5V.n4397 ASIG5V.n4386 2.2505
R45208 ASIG5V.n4399 ASIG5V.n4398 2.2505
R45209 ASIG5V.n4401 ASIG5V.n4384 2.2505
R45210 ASIG5V.n4404 ASIG5V.n4403 2.2505
R45211 ASIG5V.n4405 ASIG5V.n4382 2.2505
R45212 ASIG5V.n4407 ASIG5V.n4406 2.2505
R45213 ASIG5V.n4409 ASIG5V.n4380 2.2505
R45214 ASIG5V.n4412 ASIG5V.n4411 2.2505
R45215 ASIG5V.n4413 ASIG5V.n4378 2.2505
R45216 ASIG5V.n4415 ASIG5V.n4414 2.2505
R45217 ASIG5V.n4417 ASIG5V.n4376 2.2505
R45218 ASIG5V.n4420 ASIG5V.n4419 2.2505
R45219 ASIG5V.n4421 ASIG5V.n4374 2.2505
R45220 ASIG5V.n4423 ASIG5V.n4422 2.2505
R45221 ASIG5V.n4425 ASIG5V.n4372 2.2505
R45222 ASIG5V.n4428 ASIG5V.n4427 2.2505
R45223 ASIG5V.n4429 ASIG5V.n4370 2.2505
R45224 ASIG5V.n4431 ASIG5V.n4430 2.2505
R45225 ASIG5V.n4433 ASIG5V.n4368 2.2505
R45226 ASIG5V.n4436 ASIG5V.n4435 2.2505
R45227 ASIG5V.n4437 ASIG5V.n4366 2.2505
R45228 ASIG5V.n4439 ASIG5V.n4438 2.2505
R45229 ASIG5V.n4441 ASIG5V.n4364 2.2505
R45230 ASIG5V.n4444 ASIG5V.n4443 2.2505
R45231 ASIG5V.n4445 ASIG5V.n4362 2.2505
R45232 ASIG5V.n4447 ASIG5V.n4446 2.2505
R45233 ASIG5V.n4449 ASIG5V.n4360 2.2505
R45234 ASIG5V.n4452 ASIG5V.n4451 2.2505
R45235 ASIG5V.n4453 ASIG5V.n4358 2.2505
R45236 ASIG5V.n4455 ASIG5V.n4454 2.2505
R45237 ASIG5V.n4457 ASIG5V.n4356 2.2505
R45238 ASIG5V.n4460 ASIG5V.n4459 2.2505
R45239 ASIG5V.n4461 ASIG5V.n4354 2.2505
R45240 ASIG5V.n4463 ASIG5V.n4462 2.2505
R45241 ASIG5V.n4465 ASIG5V.n4352 2.2505
R45242 ASIG5V.n4468 ASIG5V.n4467 2.2505
R45243 ASIG5V.n4469 ASIG5V.n4350 2.2505
R45244 ASIG5V.n4471 ASIG5V.n4470 2.2505
R45245 ASIG5V.n4473 ASIG5V.n4348 2.2505
R45246 ASIG5V.n4476 ASIG5V.n4475 2.2505
R45247 ASIG5V.n4477 ASIG5V.n4346 2.2505
R45248 ASIG5V.n4479 ASIG5V.n4478 2.2505
R45249 ASIG5V.n4481 ASIG5V.n4344 2.2505
R45250 ASIG5V.n4484 ASIG5V.n4483 2.2505
R45251 ASIG5V.n4485 ASIG5V.n4342 2.2505
R45252 ASIG5V.n4487 ASIG5V.n4486 2.2505
R45253 ASIG5V.n4489 ASIG5V.n4340 2.2505
R45254 ASIG5V.n4492 ASIG5V.n4491 2.2505
R45255 ASIG5V.n4493 ASIG5V.n4338 2.2505
R45256 ASIG5V.n4495 ASIG5V.n4494 2.2505
R45257 ASIG5V.n4497 ASIG5V.n4336 2.2505
R45258 ASIG5V.n4500 ASIG5V.n4499 2.2505
R45259 ASIG5V.n4501 ASIG5V.n4334 2.2505
R45260 ASIG5V.n4503 ASIG5V.n4502 2.2505
R45261 ASIG5V.n4505 ASIG5V.n4332 2.2505
R45262 ASIG5V.n4508 ASIG5V.n4507 2.2505
R45263 ASIG5V.n4509 ASIG5V.n4330 2.2505
R45264 ASIG5V.n4511 ASIG5V.n4510 2.2505
R45265 ASIG5V.n4513 ASIG5V.n4328 2.2505
R45266 ASIG5V.n4516 ASIG5V.n4515 2.2505
R45267 ASIG5V.n4517 ASIG5V.n4326 2.2505
R45268 ASIG5V.n4519 ASIG5V.n4518 2.2505
R45269 ASIG5V.n4521 ASIG5V.n4324 2.2505
R45270 ASIG5V.n4524 ASIG5V.n4523 2.2505
R45271 ASIG5V.n4525 ASIG5V.n4322 2.2505
R45272 ASIG5V.n4527 ASIG5V.n4526 2.2505
R45273 ASIG5V.n4529 ASIG5V.n4320 2.2505
R45274 ASIG5V.n4532 ASIG5V.n4531 2.2505
R45275 ASIG5V.n4533 ASIG5V.n4318 2.2505
R45276 ASIG5V.n4535 ASIG5V.n4534 2.2505
R45277 ASIG5V.n4537 ASIG5V.n4316 2.2505
R45278 ASIG5V.n4540 ASIG5V.n4539 2.2505
R45279 ASIG5V.n4541 ASIG5V.n4314 2.2505
R45280 ASIG5V.n4543 ASIG5V.n4542 2.2505
R45281 ASIG5V.n4545 ASIG5V.n4312 2.2505
R45282 ASIG5V.n4548 ASIG5V.n4547 2.2505
R45283 ASIG5V.n4549 ASIG5V.n4311 2.2505
R45284 ASIG5V.n4551 ASIG5V.n4550 2.2505
R45285 ASIG5V.n4309 ASIG5V.n3783 2.2505
R45286 ASIG5V.n10547 ASIG5V.n10494 2.24752
R45287 ASIG5V.n3907 ASIG5V.n3855 2.24752
R45288 ASIG5V.n10550 ASIG5V.n10493 2.24752
R45289 ASIG5V.n10549 ASIG5V.n10492 2.24752
R45290 ASIG5V.n10553 ASIG5V.n10493 2.24752
R45291 ASIG5V.n10552 ASIG5V.n10492 2.24752
R45292 ASIG5V.n10556 ASIG5V.n10493 2.24752
R45293 ASIG5V.n10555 ASIG5V.n10492 2.24752
R45294 ASIG5V.n10559 ASIG5V.n10493 2.24752
R45295 ASIG5V.n10558 ASIG5V.n10492 2.24752
R45296 ASIG5V.n10562 ASIG5V.n10493 2.24752
R45297 ASIG5V.n10561 ASIG5V.n10492 2.24752
R45298 ASIG5V.n10565 ASIG5V.n10493 2.24752
R45299 ASIG5V.n10564 ASIG5V.n10492 2.24752
R45300 ASIG5V.n10568 ASIG5V.n10493 2.24752
R45301 ASIG5V.n10567 ASIG5V.n10492 2.24752
R45302 ASIG5V.n10571 ASIG5V.n10493 2.24752
R45303 ASIG5V.n10570 ASIG5V.n10492 2.24752
R45304 ASIG5V.n10574 ASIG5V.n10493 2.24752
R45305 ASIG5V.n10573 ASIG5V.n10492 2.24752
R45306 ASIG5V.n10577 ASIG5V.n10493 2.24752
R45307 ASIG5V.n10576 ASIG5V.n10492 2.24752
R45308 ASIG5V.n10580 ASIG5V.n10493 2.24752
R45309 ASIG5V.n10579 ASIG5V.n10492 2.24752
R45310 ASIG5V.n10583 ASIG5V.n10493 2.24752
R45311 ASIG5V.n10582 ASIG5V.n10492 2.24752
R45312 ASIG5V.n10586 ASIG5V.n10493 2.24752
R45313 ASIG5V.n10585 ASIG5V.n10492 2.24752
R45314 ASIG5V.n10589 ASIG5V.n10493 2.24752
R45315 ASIG5V.n10588 ASIG5V.n10492 2.24752
R45316 ASIG5V.n10592 ASIG5V.n10493 2.24752
R45317 ASIG5V.n10591 ASIG5V.n10492 2.24752
R45318 ASIG5V.n10595 ASIG5V.n10493 2.24752
R45319 ASIG5V.n10594 ASIG5V.n10492 2.24752
R45320 ASIG5V.n10598 ASIG5V.n10493 2.24752
R45321 ASIG5V.n10597 ASIG5V.n10492 2.24752
R45322 ASIG5V.n10601 ASIG5V.n10493 2.24752
R45323 ASIG5V.n10600 ASIG5V.n10492 2.24752
R45324 ASIG5V.n10604 ASIG5V.n10493 2.24752
R45325 ASIG5V.n10603 ASIG5V.n10492 2.24752
R45326 ASIG5V.n10607 ASIG5V.n10493 2.24752
R45327 ASIG5V.n10606 ASIG5V.n10492 2.24752
R45328 ASIG5V.n10610 ASIG5V.n10493 2.24752
R45329 ASIG5V.n10609 ASIG5V.n10492 2.24752
R45330 ASIG5V.n10613 ASIG5V.n10493 2.24752
R45331 ASIG5V.n10612 ASIG5V.n10492 2.24752
R45332 ASIG5V.n10616 ASIG5V.n10493 2.24752
R45333 ASIG5V.n10615 ASIG5V.n10492 2.24752
R45334 ASIG5V.n10619 ASIG5V.n10493 2.24752
R45335 ASIG5V.n10618 ASIG5V.n10492 2.24752
R45336 ASIG5V.n10622 ASIG5V.n10493 2.24752
R45337 ASIG5V.n10621 ASIG5V.n10492 2.24752
R45338 ASIG5V.n10625 ASIG5V.n10493 2.24752
R45339 ASIG5V.n10624 ASIG5V.n10492 2.24752
R45340 ASIG5V.n10628 ASIG5V.n10493 2.24752
R45341 ASIG5V.n10627 ASIG5V.n10492 2.24752
R45342 ASIG5V.n10631 ASIG5V.n10493 2.24752
R45343 ASIG5V.n10630 ASIG5V.n10492 2.24752
R45344 ASIG5V.n10634 ASIG5V.n10493 2.24752
R45345 ASIG5V.n10633 ASIG5V.n10492 2.24752
R45346 ASIG5V.n10637 ASIG5V.n10493 2.24752
R45347 ASIG5V.n10636 ASIG5V.n10492 2.24752
R45348 ASIG5V.n10640 ASIG5V.n10493 2.24752
R45349 ASIG5V.n10639 ASIG5V.n10492 2.24752
R45350 ASIG5V.n10643 ASIG5V.n10493 2.24752
R45351 ASIG5V.n10642 ASIG5V.n10492 2.24752
R45352 ASIG5V.n10646 ASIG5V.n10493 2.24752
R45353 ASIG5V.n10645 ASIG5V.n10492 2.24752
R45354 ASIG5V.n10649 ASIG5V.n10493 2.24752
R45355 ASIG5V.n10648 ASIG5V.n10492 2.24752
R45356 ASIG5V.n10652 ASIG5V.n10493 2.24752
R45357 ASIG5V.n10651 ASIG5V.n10492 2.24752
R45358 ASIG5V.n10655 ASIG5V.n10493 2.24752
R45359 ASIG5V.n10654 ASIG5V.n10492 2.24752
R45360 ASIG5V.n10658 ASIG5V.n10493 2.24752
R45361 ASIG5V.n10657 ASIG5V.n10492 2.24752
R45362 ASIG5V.n10661 ASIG5V.n10493 2.24752
R45363 ASIG5V.n10660 ASIG5V.n10492 2.24752
R45364 ASIG5V.n10664 ASIG5V.n10493 2.24752
R45365 ASIG5V.n10663 ASIG5V.n10492 2.24752
R45366 ASIG5V.n10667 ASIG5V.n10493 2.24752
R45367 ASIG5V.n10666 ASIG5V.n10492 2.24752
R45368 ASIG5V.n10670 ASIG5V.n10493 2.24752
R45369 ASIG5V.n10669 ASIG5V.n10492 2.24752
R45370 ASIG5V.n10673 ASIG5V.n10493 2.24752
R45371 ASIG5V.n10672 ASIG5V.n10492 2.24752
R45372 ASIG5V.n10676 ASIG5V.n10493 2.24752
R45373 ASIG5V.n10675 ASIG5V.n10492 2.24752
R45374 ASIG5V.n10679 ASIG5V.n10493 2.24752
R45375 ASIG5V.n10678 ASIG5V.n10492 2.24752
R45376 ASIG5V.n10682 ASIG5V.n10493 2.24752
R45377 ASIG5V.n10681 ASIG5V.n10492 2.24752
R45378 ASIG5V.n10685 ASIG5V.n10493 2.24752
R45379 ASIG5V.n10684 ASIG5V.n10492 2.24752
R45380 ASIG5V.n10688 ASIG5V.n10493 2.24752
R45381 ASIG5V.n10687 ASIG5V.n10492 2.24752
R45382 ASIG5V.n10691 ASIG5V.n10493 2.24752
R45383 ASIG5V.n10690 ASIG5V.n10492 2.24752
R45384 ASIG5V.n3851 ASIG5V.n3846 2.24752
R45385 ASIG5V.n10701 ASIG5V.n10695 2.24752
R45386 ASIG5V.n4258 ASIG5V.n3851 2.24752
R45387 ASIG5V.n10702 ASIG5V.n10701 2.24752
R45388 ASIG5V.n4051 ASIG5V.n3854 2.24752
R45389 ASIG5V.n3910 ASIG5V.n3855 2.24752
R45390 ASIG5V.n4051 ASIG5V.n4050 2.24752
R45391 ASIG5V.n3912 ASIG5V.n3855 2.24752
R45392 ASIG5V.n4051 ASIG5V.n4049 2.24752
R45393 ASIG5V.n3914 ASIG5V.n3855 2.24752
R45394 ASIG5V.n4051 ASIG5V.n4048 2.24752
R45395 ASIG5V.n3916 ASIG5V.n3855 2.24752
R45396 ASIG5V.n4051 ASIG5V.n4047 2.24752
R45397 ASIG5V.n3918 ASIG5V.n3855 2.24752
R45398 ASIG5V.n4051 ASIG5V.n4046 2.24752
R45399 ASIG5V.n3920 ASIG5V.n3855 2.24752
R45400 ASIG5V.n4051 ASIG5V.n4045 2.24752
R45401 ASIG5V.n3922 ASIG5V.n3855 2.24752
R45402 ASIG5V.n4051 ASIG5V.n4044 2.24752
R45403 ASIG5V.n3924 ASIG5V.n3855 2.24752
R45404 ASIG5V.n4051 ASIG5V.n4043 2.24752
R45405 ASIG5V.n3926 ASIG5V.n3855 2.24752
R45406 ASIG5V.n4051 ASIG5V.n4042 2.24752
R45407 ASIG5V.n3928 ASIG5V.n3855 2.24752
R45408 ASIG5V.n4051 ASIG5V.n4041 2.24752
R45409 ASIG5V.n3930 ASIG5V.n3855 2.24752
R45410 ASIG5V.n4051 ASIG5V.n4040 2.24752
R45411 ASIG5V.n3932 ASIG5V.n3855 2.24752
R45412 ASIG5V.n4051 ASIG5V.n4039 2.24752
R45413 ASIG5V.n3934 ASIG5V.n3855 2.24752
R45414 ASIG5V.n4051 ASIG5V.n4038 2.24752
R45415 ASIG5V.n3936 ASIG5V.n3855 2.24752
R45416 ASIG5V.n4051 ASIG5V.n4037 2.24752
R45417 ASIG5V.n3938 ASIG5V.n3855 2.24752
R45418 ASIG5V.n4051 ASIG5V.n4036 2.24752
R45419 ASIG5V.n3940 ASIG5V.n3855 2.24752
R45420 ASIG5V.n4051 ASIG5V.n4035 2.24752
R45421 ASIG5V.n3942 ASIG5V.n3855 2.24752
R45422 ASIG5V.n4051 ASIG5V.n4034 2.24752
R45423 ASIG5V.n3944 ASIG5V.n3855 2.24752
R45424 ASIG5V.n4051 ASIG5V.n4033 2.24752
R45425 ASIG5V.n3946 ASIG5V.n3855 2.24752
R45426 ASIG5V.n4051 ASIG5V.n4032 2.24752
R45427 ASIG5V.n3948 ASIG5V.n3855 2.24752
R45428 ASIG5V.n4051 ASIG5V.n4031 2.24752
R45429 ASIG5V.n3950 ASIG5V.n3855 2.24752
R45430 ASIG5V.n4051 ASIG5V.n4030 2.24752
R45431 ASIG5V.n3952 ASIG5V.n3855 2.24752
R45432 ASIG5V.n4051 ASIG5V.n4029 2.24752
R45433 ASIG5V.n3954 ASIG5V.n3855 2.24752
R45434 ASIG5V.n4051 ASIG5V.n4028 2.24752
R45435 ASIG5V.n3956 ASIG5V.n3855 2.24752
R45436 ASIG5V.n4051 ASIG5V.n4027 2.24752
R45437 ASIG5V.n3958 ASIG5V.n3855 2.24752
R45438 ASIG5V.n4051 ASIG5V.n4026 2.24752
R45439 ASIG5V.n3960 ASIG5V.n3855 2.24752
R45440 ASIG5V.n4051 ASIG5V.n4025 2.24752
R45441 ASIG5V.n3962 ASIG5V.n3855 2.24752
R45442 ASIG5V.n4051 ASIG5V.n4024 2.24752
R45443 ASIG5V.n3964 ASIG5V.n3855 2.24752
R45444 ASIG5V.n4051 ASIG5V.n4023 2.24752
R45445 ASIG5V.n3966 ASIG5V.n3855 2.24752
R45446 ASIG5V.n4051 ASIG5V.n4022 2.24752
R45447 ASIG5V.n3968 ASIG5V.n3855 2.24752
R45448 ASIG5V.n4051 ASIG5V.n4021 2.24752
R45449 ASIG5V.n3970 ASIG5V.n3855 2.24752
R45450 ASIG5V.n4051 ASIG5V.n4020 2.24752
R45451 ASIG5V.n3972 ASIG5V.n3855 2.24752
R45452 ASIG5V.n4051 ASIG5V.n4019 2.24752
R45453 ASIG5V.n3974 ASIG5V.n3855 2.24752
R45454 ASIG5V.n4051 ASIG5V.n4018 2.24752
R45455 ASIG5V.n3976 ASIG5V.n3855 2.24752
R45456 ASIG5V.n4051 ASIG5V.n4017 2.24752
R45457 ASIG5V.n3978 ASIG5V.n3855 2.24752
R45458 ASIG5V.n4051 ASIG5V.n4016 2.24752
R45459 ASIG5V.n3980 ASIG5V.n3855 2.24752
R45460 ASIG5V.n4051 ASIG5V.n4015 2.24752
R45461 ASIG5V.n3982 ASIG5V.n3855 2.24752
R45462 ASIG5V.n4051 ASIG5V.n4014 2.24752
R45463 ASIG5V.n3984 ASIG5V.n3855 2.24752
R45464 ASIG5V.n4051 ASIG5V.n4013 2.24752
R45465 ASIG5V.n3986 ASIG5V.n3855 2.24752
R45466 ASIG5V.n4051 ASIG5V.n4012 2.24752
R45467 ASIG5V.n3988 ASIG5V.n3855 2.24752
R45468 ASIG5V.n4051 ASIG5V.n4011 2.24752
R45469 ASIG5V.n3990 ASIG5V.n3855 2.24752
R45470 ASIG5V.n4051 ASIG5V.n4010 2.24752
R45471 ASIG5V.n3992 ASIG5V.n3855 2.24752
R45472 ASIG5V.n4051 ASIG5V.n4009 2.24752
R45473 ASIG5V.n3994 ASIG5V.n3855 2.24752
R45474 ASIG5V.n4051 ASIG5V.n4008 2.24752
R45475 ASIG5V.n3996 ASIG5V.n3855 2.24752
R45476 ASIG5V.n4051 ASIG5V.n4007 2.24752
R45477 ASIG5V.n3998 ASIG5V.n3855 2.24752
R45478 ASIG5V.n4051 ASIG5V.n4006 2.24752
R45479 ASIG5V.n4000 ASIG5V.n3855 2.24752
R45480 ASIG5V.n4051 ASIG5V.n4005 2.24752
R45481 ASIG5V.n4002 ASIG5V.n3855 2.24752
R45482 ASIG5V.n4051 ASIG5V.n4004 2.24752
R45483 ASIG5V.n4052 ASIG5V.n4051 2.24752
R45484 ASIG5V.n8099 ASIG5V.n3083 2.24636
R45485 ASIG5V.n8104 ASIG5V.n8103 2.24636
R45486 ASIG5V.n8107 ASIG5V.n8106 2.24636
R45487 ASIG5V.n9886 ASIG5V.n3081 2.24636
R45488 ASIG5V.n9883 ASIG5V.n3078 2.24636
R45489 ASIG5V.n9891 ASIG5V.n9890 2.24636
R45490 ASIG5V.n8110 ASIG5V.n8109 2.24636
R45491 ASIG5V.n8116 ASIG5V.n7463 2.24636
R45492 ASIG5V.n7634 ASIG5V.n7633 2.24636
R45493 ASIG5V.n7629 ASIG5V.n7628 2.24636
R45494 ASIG5V.n7625 ASIG5V.n7624 2.24636
R45495 ASIG5V.n8092 ASIG5V.n7475 2.24636
R45496 ASIG5V.n8093 ASIG5V.n7473 2.24636
R45497 ASIG5V.n8090 ASIG5V.n7476 2.24636
R45498 ASIG5V.n9876 ASIG5V.n3087 2.24636
R45499 ASIG5V.n9877 ASIG5V.n3085 2.24636
R45500 ASIG5V.n9874 ASIG5V.n3088 2.24636
R45501 ASIG5V.n7319 ASIG5V.n7315 2.24636
R45502 ASIG5V.n8117 ASIG5V.n7321 2.24636
R45503 ASIG5V.n8121 ASIG5V.n8120 2.24636
R45504 ASIG5V.n8124 ASIG5V.n8123 2.24636
R45505 ASIG5V.n8129 ASIG5V.n7309 2.24636
R45506 ASIG5V.n7617 ASIG5V.n7616 2.24636
R45507 ASIG5V.n7612 ASIG5V.n7611 2.24636
R45508 ASIG5V.n7608 ASIG5V.n7607 2.24636
R45509 ASIG5V.n7636 ASIG5V.n7571 2.24636
R45510 ASIG5V.n7640 ASIG5V.n7639 2.24636
R45511 ASIG5V.n7643 ASIG5V.n7642 2.24636
R45512 ASIG5V.n8083 ASIG5V.n7482 2.24636
R45513 ASIG5V.n8084 ASIG5V.n7480 2.24636
R45514 ASIG5V.n8081 ASIG5V.n7483 2.24636
R45515 ASIG5V.n9867 ASIG5V.n3094 2.24636
R45516 ASIG5V.n9868 ASIG5V.n3092 2.24636
R45517 ASIG5V.n9865 ASIG5V.n3095 2.24636
R45518 ASIG5V.n7298 ASIG5V.n7294 2.24636
R45519 ASIG5V.n8130 ASIG5V.n7300 2.24636
R45520 ASIG5V.n7459 ASIG5V.n7458 2.24636
R45521 ASIG5V.n7454 ASIG5V.n7453 2.24636
R45522 ASIG5V.n8134 ASIG5V.n8133 2.24636
R45523 ASIG5V.n7456 ASIG5V.n7449 2.24636
R45524 ASIG5V.n8137 ASIG5V.n8136 2.24636
R45525 ASIG5V.n8142 ASIG5V.n7289 2.24636
R45526 ASIG5V.n7592 ASIG5V.n7579 2.24636
R45527 ASIG5V.n7585 ASIG5V.n7580 2.24636
R45528 ASIG5V.n7590 ASIG5V.n7589 2.24636
R45529 ASIG5V.n7597 ASIG5V.n7566 2.24636
R45530 ASIG5V.n7595 ASIG5V.n7576 2.24636
R45531 ASIG5V.n7599 ASIG5V.n7593 2.24636
R45532 ASIG5V.n7645 ASIG5V.n7563 2.24636
R45533 ASIG5V.n7649 ASIG5V.n7648 2.24636
R45534 ASIG5V.n7652 ASIG5V.n7651 2.24636
R45535 ASIG5V.n8074 ASIG5V.n7489 2.24636
R45536 ASIG5V.n8075 ASIG5V.n7487 2.24636
R45537 ASIG5V.n8072 ASIG5V.n7490 2.24636
R45538 ASIG5V.n9858 ASIG5V.n3101 2.24636
R45539 ASIG5V.n9859 ASIG5V.n3099 2.24636
R45540 ASIG5V.n9856 ASIG5V.n3102 2.24636
R45541 ASIG5V.n7278 ASIG5V.n7274 2.24636
R45542 ASIG5V.n8143 ASIG5V.n7280 2.24636
R45543 ASIG5V.n7365 ASIG5V.n7303 2.24636
R45544 ASIG5V.n7448 ASIG5V.n7447 2.24636
R45545 ASIG5V.n7443 ASIG5V.n7442 2.24636
R45546 ASIG5V.n7374 ASIG5V.n7373 2.24636
R45547 ASIG5V.n8147 ASIG5V.n8146 2.24636
R45548 ASIG5V.n7445 ASIG5V.n7438 2.24636
R45549 ASIG5V.n7377 ASIG5V.n7376 2.24636
R45550 ASIG5V.n8150 ASIG5V.n8149 2.24636
R45551 ASIG5V.n8155 ASIG5V.n7268 2.24636
R45552 ASIG5V.n7688 ASIG5V.n7687 2.24636
R45553 ASIG5V.n7694 ASIG5V.n7693 2.24636
R45554 ASIG5V.n7697 ASIG5V.n7696 2.24636
R45555 ASIG5V.n7677 ASIG5V.n7676 2.24636
R45556 ASIG5V.n7683 ASIG5V.n7682 2.24636
R45557 ASIG5V.n7686 ASIG5V.n7685 2.24636
R45558 ASIG5V.n7666 ASIG5V.n7665 2.24636
R45559 ASIG5V.n7672 ASIG5V.n7671 2.24636
R45560 ASIG5V.n7675 ASIG5V.n7674 2.24636
R45561 ASIG5V.n7655 ASIG5V.n7654 2.24636
R45562 ASIG5V.n7661 ASIG5V.n7660 2.24636
R45563 ASIG5V.n7664 ASIG5V.n7663 2.24636
R45564 ASIG5V.n8065 ASIG5V.n7496 2.24636
R45565 ASIG5V.n8066 ASIG5V.n7494 2.24636
R45566 ASIG5V.n8063 ASIG5V.n7497 2.24636
R45567 ASIG5V.n9849 ASIG5V.n3108 2.24636
R45568 ASIG5V.n9850 ASIG5V.n3106 2.24636
R45569 ASIG5V.n9847 ASIG5V.n3109 2.24636
R45570 ASIG5V.n7698 ASIG5V.n7542 2.24636
R45571 ASIG5V.n8156 ASIG5V.n7260 2.24636
R45572 ASIG5V.n7350 ASIG5V.n7283 2.24636
R45573 ASIG5V.n7378 ASIG5V.n7358 2.24636
R45574 ASIG5V.n7437 ASIG5V.n7436 2.24636
R45575 ASIG5V.n7432 ASIG5V.n7431 2.24636
R45576 ASIG5V.n7382 ASIG5V.n7381 2.24636
R45577 ASIG5V.n7356 ASIG5V.n7351 2.24636
R45578 ASIG5V.n7266 ASIG5V.n7261 2.24636
R45579 ASIG5V.n7434 ASIG5V.n7427 2.24636
R45580 ASIG5V.n7385 ASIG5V.n7384 2.24636
R45581 ASIG5V.n7391 ASIG5V.n7348 2.24636
R45582 ASIG5V.n8161 ASIG5V.n7257 2.24636
R45583 ASIG5V.n7704 ASIG5V.n7703 2.24636
R45584 ASIG5V.n9764 ASIG5V.n3149 2.24636
R45585 ASIG5V.n9757 ASIG5V.n3150 2.24636
R45586 ASIG5V.n9762 ASIG5V.n9761 2.24636
R45587 ASIG5V.n9776 ASIG5V.n3144 2.24636
R45588 ASIG5V.n9770 ASIG5V.n3145 2.24636
R45589 ASIG5V.n9768 ASIG5V.n9765 2.24636
R45590 ASIG5V.n9788 ASIG5V.n3139 2.24636
R45591 ASIG5V.n9782 ASIG5V.n3140 2.24636
R45592 ASIG5V.n9780 ASIG5V.n9777 2.24636
R45593 ASIG5V.n9800 ASIG5V.n3134 2.24636
R45594 ASIG5V.n9794 ASIG5V.n3135 2.24636
R45595 ASIG5V.n9792 ASIG5V.n9789 2.24636
R45596 ASIG5V.n9812 ASIG5V.n3129 2.24636
R45597 ASIG5V.n9806 ASIG5V.n3130 2.24636
R45598 ASIG5V.n9804 ASIG5V.n9801 2.24636
R45599 ASIG5V.n9824 ASIG5V.n3124 2.24636
R45600 ASIG5V.n9818 ASIG5V.n3125 2.24636
R45601 ASIG5V.n9816 ASIG5V.n9813 2.24636
R45602 ASIG5V.n9831 ASIG5V.n3122 2.24636
R45603 ASIG5V.n9832 ASIG5V.n3120 2.24636
R45604 ASIG5V.n9829 ASIG5V.n9825 2.24636
R45605 ASIG5V.n9754 ASIG5V.n3155 2.24636
R45606 ASIG5V.n7705 ASIG5V.n7534 2.24636
R45607 ASIG5V.n8162 ASIG5V.n7249 2.24636
R45608 ASIG5V.n7398 ASIG5V.n7392 2.24636
R45609 ASIG5V.n7407 ASIG5V.n7338 2.24636
R45610 ASIG5V.n7426 ASIG5V.n7425 2.24636
R45611 ASIG5V.n7421 ASIG5V.n7420 2.24636
R45612 ASIG5V.n7408 ASIG5V.n7336 2.24636
R45613 ASIG5V.n7399 ASIG5V.n7345 2.24636
R45614 ASIG5V.n7255 ASIG5V.n7250 2.24636
R45615 ASIG5V.n7709 ASIG5V.n7708 2.24636
R45616 ASIG5V.n7423 ASIG5V.n1841 2.24636
R45617 ASIG5V.n7405 ASIG5V.n7341 2.24636
R45618 ASIG5V.n7396 ASIG5V.n169 2.24636
R45619 ASIG5V.n8167 ASIG5V.n7246 2.24636
R45620 ASIG5V.n7712 ASIG5V.n7711 2.24636
R45621 ASIG5V.n9752 ASIG5V.n9751 2.24636
R45622 ASIG5V.n9944 ASIG5V.n9943 2.24636
R45623 ASIG5V.n9949 ASIG5V.n9948 2.24636
R45624 ASIG5V.n9952 ASIG5V.n9951 2.24636
R45625 ASIG5V.n9937 ASIG5V.n3014 2.24636
R45626 ASIG5V.n3020 ASIG5V.n3015 2.24636
R45627 ASIG5V.n9942 ASIG5V.n3011 2.24636
R45628 ASIG5V.n9931 ASIG5V.n3025 2.24636
R45629 ASIG5V.n3031 ASIG5V.n3026 2.24636
R45630 ASIG5V.n9936 ASIG5V.n3022 2.24636
R45631 ASIG5V.n9925 ASIG5V.n3036 2.24636
R45632 ASIG5V.n3042 ASIG5V.n3037 2.24636
R45633 ASIG5V.n9930 ASIG5V.n3033 2.24636
R45634 ASIG5V.n9919 ASIG5V.n3047 2.24636
R45635 ASIG5V.n3053 ASIG5V.n3048 2.24636
R45636 ASIG5V.n9924 ASIG5V.n3044 2.24636
R45637 ASIG5V.n9913 ASIG5V.n3058 2.24636
R45638 ASIG5V.n3064 ASIG5V.n3059 2.24636
R45639 ASIG5V.n9918 ASIG5V.n3055 2.24636
R45640 ASIG5V.n9907 ASIG5V.n3069 2.24636
R45641 ASIG5V.n3075 ASIG5V.n3070 2.24636
R45642 ASIG5V.n9912 ASIG5V.n3066 2.24636
R45643 ASIG5V.n9901 ASIG5V.n9894 2.24636
R45644 ASIG5V.n9900 ASIG5V.n9895 2.24636
R45645 ASIG5V.n9906 ASIG5V.n3077 2.24636
R45646 ASIG5V.n7995 ASIG5V.n7530 2.24636
R45647 ASIG5V.n7989 ASIG5V.n7531 2.24636
R45648 ASIG5V.n7986 ASIG5V.n7983 2.24636
R45649 ASIG5V.n8006 ASIG5V.n7525 2.24636
R45650 ASIG5V.n7998 ASIG5V.n7526 2.24636
R45651 ASIG5V.n8001 ASIG5V.n7996 2.24636
R45652 ASIG5V.n8017 ASIG5V.n7520 2.24636
R45653 ASIG5V.n8009 ASIG5V.n7521 2.24636
R45654 ASIG5V.n8012 ASIG5V.n8007 2.24636
R45655 ASIG5V.n8028 ASIG5V.n7515 2.24636
R45656 ASIG5V.n8020 ASIG5V.n7516 2.24636
R45657 ASIG5V.n8023 ASIG5V.n8018 2.24636
R45658 ASIG5V.n8039 ASIG5V.n7510 2.24636
R45659 ASIG5V.n8031 ASIG5V.n7511 2.24636
R45660 ASIG5V.n8034 ASIG5V.n8029 2.24636
R45661 ASIG5V.n8050 ASIG5V.n7505 2.24636
R45662 ASIG5V.n8042 ASIG5V.n7506 2.24636
R45663 ASIG5V.n8045 ASIG5V.n8040 2.24636
R45664 ASIG5V.n8055 ASIG5V.n7503 2.24636
R45665 ASIG5V.n8053 ASIG5V.n7501 2.24636
R45666 ASIG5V.n8057 ASIG5V.n8051 2.24636
R45667 ASIG5V.n9840 ASIG5V.n3115 2.24636
R45668 ASIG5V.n9841 ASIG5V.n3113 2.24636
R45669 ASIG5V.n9838 ASIG5V.n3116 2.24636
R45670 ASIG5V.n8105 ASIG5V.n7471 2.24552
R45671 ASIG5V.n8101 ASIG5V.n8100 2.24552
R45672 ASIG5V.n8102 ASIG5V.n7469 2.24552
R45673 ASIG5V.n8100 ASIG5V.n7468 2.24552
R45674 ASIG5V.n9889 ASIG5V.n9888 2.24552
R45675 ASIG5V.n9885 ASIG5V.n9884 2.24552
R45676 ASIG5V.n9887 ASIG5V.n3084 2.24552
R45677 ASIG5V.n9885 ASIG5V.n3082 2.24552
R45678 ASIG5V.n8108 ASIG5V.n7467 2.24552
R45679 ASIG5V.n8112 ASIG5V.n8111 2.24552
R45680 ASIG5V.n8113 ASIG5V.n7467 2.24552
R45681 ASIG5V.n7462 ASIG5V.n3056 2.24552
R45682 ASIG5V.n7632 ASIG5V.n7630 2.24552
R45683 ASIG5V.n7635 ASIG5V.n7622 2.24552
R45684 ASIG5V.n7627 ASIG5V.n7623 2.24552
R45685 ASIG5V.n7635 ASIG5V.n7621 2.24552
R45686 ASIG5V.n7479 ASIG5V.n7478 2.24552
R45687 ASIG5V.n8095 ASIG5V.n8094 2.24552
R45688 ASIG5V.n8091 ASIG5V.n7477 2.24552
R45689 ASIG5V.n8098 ASIG5V.n8097 2.24552
R45690 ASIG5V.n3091 ASIG5V.n3090 2.24552
R45691 ASIG5V.n9879 ASIG5V.n9878 2.24552
R45692 ASIG5V.n9875 ASIG5V.n3089 2.24552
R45693 ASIG5V.n9882 ASIG5V.n9881 2.24552
R45694 ASIG5V.n7314 ASIG5V.n7313 2.24552
R45695 ASIG5V.n8122 ASIG5V.n8118 2.24552
R45696 ASIG5V.n8125 ASIG5V.n7322 2.24552
R45697 ASIG5V.n7318 ASIG5V.n7316 2.24552
R45698 ASIG5V.n8119 ASIG5V.n7460 2.24552
R45699 ASIG5V.n7317 ASIG5V.n7313 2.24552
R45700 ASIG5V.n7323 ASIG5V.n3045 2.24552
R45701 ASIG5V.n8126 ASIG5V.n7308 2.24552
R45702 ASIG5V.n7610 ASIG5V.n7574 2.24552
R45703 ASIG5V.n7615 ASIG5V.n7614 2.24552
R45704 ASIG5V.n7606 ASIG5V.n7575 2.24552
R45705 ASIG5V.n7615 ASIG5V.n7605 2.24552
R45706 ASIG5V.n7641 ASIG5V.n7619 2.24552
R45707 ASIG5V.n7644 ASIG5V.n7572 2.24552
R45708 ASIG5V.n7638 ASIG5V.n7618 2.24552
R45709 ASIG5V.n7637 ASIG5V.n7573 2.24552
R45710 ASIG5V.n7486 ASIG5V.n7485 2.24552
R45711 ASIG5V.n8086 ASIG5V.n8085 2.24552
R45712 ASIG5V.n8082 ASIG5V.n7484 2.24552
R45713 ASIG5V.n8089 ASIG5V.n8088 2.24552
R45714 ASIG5V.n3098 ASIG5V.n3097 2.24552
R45715 ASIG5V.n9870 ASIG5V.n9869 2.24552
R45716 ASIG5V.n9866 ASIG5V.n3096 2.24552
R45717 ASIG5V.n9873 ASIG5V.n9872 2.24552
R45718 ASIG5V.n7293 ASIG5V.n7292 2.24552
R45719 ASIG5V.n8135 ASIG5V.n7305 2.24552
R45720 ASIG5V.n7455 ASIG5V.n7324 2.24552
R45721 ASIG5V.n7452 ASIG5V.n7307 2.24552
R45722 ASIG5V.n8138 ASIG5V.n7301 2.24552
R45723 ASIG5V.n7297 ASIG5V.n7295 2.24552
R45724 ASIG5V.n7457 ASIG5V.n7325 2.24552
R45725 ASIG5V.n8132 ASIG5V.n7304 2.24552
R45726 ASIG5V.n7296 ASIG5V.n7292 2.24552
R45727 ASIG5V.n7450 ASIG5V.n3034 2.24552
R45728 ASIG5V.n8131 ASIG5V.n7302 2.24552
R45729 ASIG5V.n8139 ASIG5V.n7288 2.24552
R45730 ASIG5V.n7588 ASIG5V.n7578 2.24552
R45731 ASIG5V.n7584 ASIG5V.n7552 2.24552
R45732 ASIG5V.n7587 ASIG5V.n7586 2.24552
R45733 ASIG5V.n7583 ASIG5V.n7552 2.24552
R45734 ASIG5V.n7601 ASIG5V.n7600 2.24552
R45735 ASIG5V.n7594 ASIG5V.n7557 2.24552
R45736 ASIG5V.n7598 ASIG5V.n7596 2.24552
R45737 ASIG5V.n7604 ASIG5V.n7603 2.24552
R45738 ASIG5V.n7650 ASIG5V.n7568 2.24552
R45739 ASIG5V.n7653 ASIG5V.n7564 2.24552
R45740 ASIG5V.n7647 ASIG5V.n7567 2.24552
R45741 ASIG5V.n7646 ASIG5V.n7565 2.24552
R45742 ASIG5V.n7493 ASIG5V.n7492 2.24552
R45743 ASIG5V.n8077 ASIG5V.n8076 2.24552
R45744 ASIG5V.n8073 ASIG5V.n7491 2.24552
R45745 ASIG5V.n8080 ASIG5V.n8079 2.24552
R45746 ASIG5V.n3105 ASIG5V.n3104 2.24552
R45747 ASIG5V.n9861 ASIG5V.n9860 2.24552
R45748 ASIG5V.n9857 ASIG5V.n3103 2.24552
R45749 ASIG5V.n9864 ASIG5V.n9863 2.24552
R45750 ASIG5V.n7273 ASIG5V.n7272 2.24552
R45751 ASIG5V.n8148 ASIG5V.n7285 2.24552
R45752 ASIG5V.n7375 ASIG5V.n7368 2.24552
R45753 ASIG5V.n7444 ASIG5V.n7327 2.24552
R45754 ASIG5V.n7441 ASIG5V.n7328 2.24552
R45755 ASIG5V.n7371 ASIG5V.n7287 2.24552
R45756 ASIG5V.n8151 ASIG5V.n7281 2.24552
R45757 ASIG5V.n7277 ASIG5V.n7275 2.24552
R45758 ASIG5V.n7446 ASIG5V.n7329 2.24552
R45759 ASIG5V.n7372 ASIG5V.n7366 2.24552
R45760 ASIG5V.n8145 ASIG5V.n7284 2.24552
R45761 ASIG5V.n7276 ASIG5V.n7272 2.24552
R45762 ASIG5V.n7439 ASIG5V.n3023 2.24552
R45763 ASIG5V.n7369 ASIG5V.n7364 2.24552
R45764 ASIG5V.n8144 ASIG5V.n7282 2.24552
R45765 ASIG5V.n8152 ASIG5V.n7267 2.24552
R45766 ASIG5V.n7695 ASIG5V.n7689 2.24552
R45767 ASIG5V.n7691 ASIG5V.n7523 2.24552
R45768 ASIG5V.n7692 ASIG5V.n7546 2.24552
R45769 ASIG5V.n7545 ASIG5V.n7523 2.24552
R45770 ASIG5V.n7684 ASIG5V.n7551 2.24552
R45771 ASIG5V.n7680 ASIG5V.n7518 2.24552
R45772 ASIG5V.n7681 ASIG5V.n7549 2.24552
R45773 ASIG5V.n7678 ASIG5V.n7548 2.24552
R45774 ASIG5V.n7673 ASIG5V.n7556 2.24552
R45775 ASIG5V.n7669 ASIG5V.n7513 2.24552
R45776 ASIG5V.n7670 ASIG5V.n7554 2.24552
R45777 ASIG5V.n7667 ASIG5V.n7553 2.24552
R45778 ASIG5V.n7662 ASIG5V.n7561 2.24552
R45779 ASIG5V.n7658 ASIG5V.n7508 2.24552
R45780 ASIG5V.n7659 ASIG5V.n7559 2.24552
R45781 ASIG5V.n7656 ASIG5V.n7558 2.24552
R45782 ASIG5V.n7500 ASIG5V.n7499 2.24552
R45783 ASIG5V.n8068 ASIG5V.n8067 2.24552
R45784 ASIG5V.n8064 ASIG5V.n7498 2.24552
R45785 ASIG5V.n8071 ASIG5V.n8070 2.24552
R45786 ASIG5V.n3112 ASIG5V.n3111 2.24552
R45787 ASIG5V.n9852 ASIG5V.n9851 2.24552
R45788 ASIG5V.n9848 ASIG5V.n3110 2.24552
R45789 ASIG5V.n9855 ASIG5V.n9854 2.24552
R45790 ASIG5V.n7699 ASIG5V.n7540 2.24552
R45791 ASIG5V.n7265 ASIG5V.n7262 2.24552
R45792 ASIG5V.n7355 ASIG5V.n7352 2.24552
R45793 ASIG5V.n7383 ASIG5V.n7362 2.24552
R45794 ASIG5V.n7433 ASIG5V.n7331 2.24552
R45795 ASIG5V.n7430 ASIG5V.n7332 2.24552
R45796 ASIG5V.n7386 ASIG5V.n7359 2.24552
R45797 ASIG5V.n7390 ASIG5V.n7389 2.24552
R45798 ASIG5V.n8160 ASIG5V.n8159 2.24552
R45799 ASIG5V.n7702 ASIG5V.n7701 2.24552
R45800 ASIG5V.n7435 ASIG5V.n7333 2.24552
R45801 ASIG5V.n7380 ASIG5V.n7361 2.24552
R45802 ASIG5V.n7354 ASIG5V.n7353 2.24552
R45803 ASIG5V.n7264 ASIG5V.n7263 2.24552
R45804 ASIG5V.n7543 ASIG5V.n7540 2.24552
R45805 ASIG5V.n7428 ASIG5V.n3012 2.24552
R45806 ASIG5V.n7379 ASIG5V.n7360 2.24552
R45807 ASIG5V.n7387 ASIG5V.n7347 2.24552
R45808 ASIG5V.n8157 ASIG5V.n7256 2.24552
R45809 ASIG5V.n7539 ASIG5V.n7258 2.24552
R45810 ASIG5V.n9760 ASIG5V.n3148 2.24552
R45811 ASIG5V.n9756 ASIG5V.n9755 2.24552
R45812 ASIG5V.n9759 ASIG5V.n9758 2.24552
R45813 ASIG5V.n9755 ASIG5V.n3154 2.24552
R45814 ASIG5V.n9769 ASIG5V.n3143 2.24552
R45815 ASIG5V.n9772 ASIG5V.n9771 2.24552
R45816 ASIG5V.n9767 ASIG5V.n9766 2.24552
R45817 ASIG5V.n9775 ASIG5V.n9774 2.24552
R45818 ASIG5V.n9781 ASIG5V.n3138 2.24552
R45819 ASIG5V.n9784 ASIG5V.n9783 2.24552
R45820 ASIG5V.n9779 ASIG5V.n9778 2.24552
R45821 ASIG5V.n9787 ASIG5V.n9786 2.24552
R45822 ASIG5V.n9793 ASIG5V.n3133 2.24552
R45823 ASIG5V.n9796 ASIG5V.n9795 2.24552
R45824 ASIG5V.n9791 ASIG5V.n9790 2.24552
R45825 ASIG5V.n9799 ASIG5V.n9798 2.24552
R45826 ASIG5V.n9805 ASIG5V.n3128 2.24552
R45827 ASIG5V.n9808 ASIG5V.n9807 2.24552
R45828 ASIG5V.n9803 ASIG5V.n9802 2.24552
R45829 ASIG5V.n9811 ASIG5V.n9810 2.24552
R45830 ASIG5V.n9817 ASIG5V.n3123 2.24552
R45831 ASIG5V.n9820 ASIG5V.n9819 2.24552
R45832 ASIG5V.n9815 ASIG5V.n9814 2.24552
R45833 ASIG5V.n9823 ASIG5V.n9822 2.24552
R45834 ASIG5V.n9828 ASIG5V.n9827 2.24552
R45835 ASIG5V.n9834 ASIG5V.n9833 2.24552
R45836 ASIG5V.n9830 ASIG5V.n9826 2.24552
R45837 ASIG5V.n9837 ASIG5V.n9836 2.24552
R45838 ASIG5V.n3159 ASIG5V.n3156 2.24552
R45839 ASIG5V.n7710 ASIG5V.n7706 2.24552
R45840 ASIG5V.n7254 ASIG5V.n7251 2.24552
R45841 ASIG5V.n7395 ASIG5V.n7394 2.24552
R45842 ASIG5V.n7344 ASIG5V.n7343 2.24552
R45843 ASIG5V.n7422 ASIG5V.n7335 2.24552
R45844 ASIG5V.n7419 ASIG5V.n7414 2.24552
R45845 ASIG5V.n7410 ASIG5V.n7409 2.24552
R45846 ASIG5V.n7401 ASIG5V.n7400 2.24552
R45847 ASIG5V.n8166 ASIG5V.n8165 2.24552
R45848 ASIG5V.n7713 ASIG5V.n7535 2.24552
R45849 ASIG5V.n9750 ASIG5V.n9749 2.24552
R45850 ASIG5V.n7424 ASIG5V.n7415 2.24552
R45851 ASIG5V.n7406 ASIG5V.n7342 2.24552
R45852 ASIG5V.n7397 ASIG5V.n7393 2.24552
R45853 ASIG5V.n7253 ASIG5V.n7252 2.24552
R45854 ASIG5V.n7707 ASIG5V.n7537 2.24552
R45855 ASIG5V.n3160 ASIG5V.n3159 2.24552
R45856 ASIG5V.n7417 ASIG5V.n3009 2.24552
R45857 ASIG5V.n7413 ASIG5V.n7412 2.24552
R45858 ASIG5V.n7404 ASIG5V.n7403 2.24552
R45859 ASIG5V.n8163 ASIG5V.n7245 2.24552
R45860 ASIG5V.n7536 ASIG5V.n7247 2.24552
R45861 ASIG5V.n7988 ASIG5V.n3162 2.24552
R45862 ASIG5V.n9950 ASIG5V.n3007 2.24552
R45863 ASIG5V.n9946 ASIG5V.n9945 2.24552
R45864 ASIG5V.n9947 ASIG5V.n3005 2.24552
R45865 ASIG5V.n9945 ASIG5V.n3003 2.24552
R45866 ASIG5V.n3019 ASIG5V.n3016 2.24552
R45867 ASIG5V.n9941 ASIG5V.n9940 2.24552
R45868 ASIG5V.n3018 ASIG5V.n3017 2.24552
R45869 ASIG5V.n9938 ASIG5V.n3010 2.24552
R45870 ASIG5V.n3030 ASIG5V.n3027 2.24552
R45871 ASIG5V.n9935 ASIG5V.n9934 2.24552
R45872 ASIG5V.n3029 ASIG5V.n3028 2.24552
R45873 ASIG5V.n9932 ASIG5V.n3021 2.24552
R45874 ASIG5V.n3041 ASIG5V.n3038 2.24552
R45875 ASIG5V.n9929 ASIG5V.n9928 2.24552
R45876 ASIG5V.n3040 ASIG5V.n3039 2.24552
R45877 ASIG5V.n9926 ASIG5V.n3032 2.24552
R45878 ASIG5V.n3052 ASIG5V.n3049 2.24552
R45879 ASIG5V.n9923 ASIG5V.n9922 2.24552
R45880 ASIG5V.n3051 ASIG5V.n3050 2.24552
R45881 ASIG5V.n9920 ASIG5V.n3043 2.24552
R45882 ASIG5V.n3063 ASIG5V.n3060 2.24552
R45883 ASIG5V.n9917 ASIG5V.n9916 2.24552
R45884 ASIG5V.n3062 ASIG5V.n3061 2.24552
R45885 ASIG5V.n9914 ASIG5V.n3054 2.24552
R45886 ASIG5V.n3074 ASIG5V.n3071 2.24552
R45887 ASIG5V.n9911 ASIG5V.n9910 2.24552
R45888 ASIG5V.n3073 ASIG5V.n3072 2.24552
R45889 ASIG5V.n9908 ASIG5V.n3065 2.24552
R45890 ASIG5V.n9899 ASIG5V.n9896 2.24552
R45891 ASIG5V.n9905 ASIG5V.n9904 2.24552
R45892 ASIG5V.n9898 ASIG5V.n9897 2.24552
R45893 ASIG5V.n9902 ASIG5V.n3076 2.24552
R45894 ASIG5V.n7987 ASIG5V.n7529 2.24552
R45895 ASIG5V.n7991 ASIG5V.n7990 2.24552
R45896 ASIG5V.n7985 ASIG5V.n7984 2.24552
R45897 ASIG5V.n7994 ASIG5V.n7993 2.24552
R45898 ASIG5V.n8002 ASIG5V.n7524 2.24552
R45899 ASIG5V.n7997 ASIG5V.n3153 2.24552
R45900 ASIG5V.n8000 ASIG5V.n7999 2.24552
R45901 ASIG5V.n8005 ASIG5V.n8004 2.24552
R45902 ASIG5V.n8013 ASIG5V.n7519 2.24552
R45903 ASIG5V.n8008 ASIG5V.n3147 2.24552
R45904 ASIG5V.n8011 ASIG5V.n8010 2.24552
R45905 ASIG5V.n8016 ASIG5V.n8015 2.24552
R45906 ASIG5V.n8024 ASIG5V.n7514 2.24552
R45907 ASIG5V.n8019 ASIG5V.n3142 2.24552
R45908 ASIG5V.n8022 ASIG5V.n8021 2.24552
R45909 ASIG5V.n8027 ASIG5V.n8026 2.24552
R45910 ASIG5V.n8035 ASIG5V.n7509 2.24552
R45911 ASIG5V.n8030 ASIG5V.n3137 2.24552
R45912 ASIG5V.n8033 ASIG5V.n8032 2.24552
R45913 ASIG5V.n8038 ASIG5V.n8037 2.24552
R45914 ASIG5V.n8046 ASIG5V.n7504 2.24552
R45915 ASIG5V.n8041 ASIG5V.n3132 2.24552
R45916 ASIG5V.n8044 ASIG5V.n8043 2.24552
R45917 ASIG5V.n8049 ASIG5V.n8048 2.24552
R45918 ASIG5V.n8059 ASIG5V.n8058 2.24552
R45919 ASIG5V.n8052 ASIG5V.n3127 2.24552
R45920 ASIG5V.n8056 ASIG5V.n8054 2.24552
R45921 ASIG5V.n8062 ASIG5V.n8061 2.24552
R45922 ASIG5V.n3119 ASIG5V.n3118 2.24552
R45923 ASIG5V.n9843 ASIG5V.n9842 2.24552
R45924 ASIG5V.n9839 ASIG5V.n3117 2.24552
R45925 ASIG5V.n9846 ASIG5V.n9845 2.24552
R45926 ASIG5V.n10356 ASIG5V.n10355 2.24164
R45927 ASIG5V.n11183 ASIG5V.n10066 2.24164
R45928 ASIG5V.n10356 ASIG5V.n10115 2.24164
R45929 ASIG5V.n11183 ASIG5V.n10065 2.24164
R45930 ASIG5V.n10356 ASIG5V.n10114 2.24164
R45931 ASIG5V.n11183 ASIG5V.n10064 2.24164
R45932 ASIG5V.n10356 ASIG5V.n10113 2.24164
R45933 ASIG5V.n11183 ASIG5V.n10063 2.24164
R45934 ASIG5V.n10356 ASIG5V.n10112 2.24164
R45935 ASIG5V.n11183 ASIG5V.n10062 2.24164
R45936 ASIG5V.n10356 ASIG5V.n10111 2.24164
R45937 ASIG5V.n11183 ASIG5V.n10061 2.24164
R45938 ASIG5V.n10356 ASIG5V.n10110 2.24164
R45939 ASIG5V.n11183 ASIG5V.n10060 2.24164
R45940 ASIG5V.n10356 ASIG5V.n10109 2.24164
R45941 ASIG5V.n11183 ASIG5V.n10059 2.24164
R45942 ASIG5V.n10356 ASIG5V.n10108 2.24164
R45943 ASIG5V.n11183 ASIG5V.n10058 2.24164
R45944 ASIG5V.n10356 ASIG5V.n10107 2.24164
R45945 ASIG5V.n11183 ASIG5V.n10057 2.24164
R45946 ASIG5V.n10356 ASIG5V.n10106 2.24164
R45947 ASIG5V.n11183 ASIG5V.n10056 2.24164
R45948 ASIG5V.n10356 ASIG5V.n10105 2.24164
R45949 ASIG5V.n11183 ASIG5V.n10055 2.24164
R45950 ASIG5V.n10356 ASIG5V.n10104 2.24164
R45951 ASIG5V.n11183 ASIG5V.n10054 2.24164
R45952 ASIG5V.n10356 ASIG5V.n10103 2.24164
R45953 ASIG5V.n11183 ASIG5V.n10053 2.24164
R45954 ASIG5V.n10356 ASIG5V.n10102 2.24164
R45955 ASIG5V.n11183 ASIG5V.n10052 2.24164
R45956 ASIG5V.n10356 ASIG5V.n10101 2.24164
R45957 ASIG5V.n11183 ASIG5V.n10051 2.24164
R45958 ASIG5V.n10356 ASIG5V.n10100 2.24164
R45959 ASIG5V.n11183 ASIG5V.n10050 2.24164
R45960 ASIG5V.n10356 ASIG5V.n10099 2.24164
R45961 ASIG5V.n11183 ASIG5V.n10049 2.24164
R45962 ASIG5V.n10356 ASIG5V.n10098 2.24164
R45963 ASIG5V.n11183 ASIG5V.n10048 2.24164
R45964 ASIG5V.n10356 ASIG5V.n10097 2.24164
R45965 ASIG5V.n11183 ASIG5V.n10047 2.24164
R45966 ASIG5V.n10356 ASIG5V.n10096 2.24164
R45967 ASIG5V.n11183 ASIG5V.n10046 2.24164
R45968 ASIG5V.n10356 ASIG5V.n10095 2.24164
R45969 ASIG5V.n11183 ASIG5V.n10045 2.24164
R45970 ASIG5V.n10356 ASIG5V.n10094 2.24164
R45971 ASIG5V.n11183 ASIG5V.n10044 2.24164
R45972 ASIG5V.n10356 ASIG5V.n10093 2.24164
R45973 ASIG5V.n11183 ASIG5V.n10043 2.24164
R45974 ASIG5V.n10356 ASIG5V.n10092 2.24164
R45975 ASIG5V.n11183 ASIG5V.n10042 2.24164
R45976 ASIG5V.n10356 ASIG5V.n10091 2.24164
R45977 ASIG5V.n11183 ASIG5V.n10041 2.24164
R45978 ASIG5V.n10356 ASIG5V.n10090 2.24164
R45979 ASIG5V.n11183 ASIG5V.n10040 2.24164
R45980 ASIG5V.n10356 ASIG5V.n10089 2.24164
R45981 ASIG5V.n11183 ASIG5V.n10039 2.24164
R45982 ASIG5V.n10356 ASIG5V.n10088 2.24164
R45983 ASIG5V.n11183 ASIG5V.n10038 2.24164
R45984 ASIG5V.n10356 ASIG5V.n10087 2.24164
R45985 ASIG5V.n11183 ASIG5V.n10037 2.24164
R45986 ASIG5V.n10356 ASIG5V.n10086 2.24164
R45987 ASIG5V.n11183 ASIG5V.n10036 2.24164
R45988 ASIG5V.n10356 ASIG5V.n10085 2.24164
R45989 ASIG5V.n11183 ASIG5V.n10035 2.24164
R45990 ASIG5V.n10356 ASIG5V.n10084 2.24164
R45991 ASIG5V.n11183 ASIG5V.n10034 2.24164
R45992 ASIG5V.n10356 ASIG5V.n10083 2.24164
R45993 ASIG5V.n11183 ASIG5V.n10033 2.24164
R45994 ASIG5V.n10356 ASIG5V.n10082 2.24164
R45995 ASIG5V.n11183 ASIG5V.n10032 2.24164
R45996 ASIG5V.n10356 ASIG5V.n10081 2.24164
R45997 ASIG5V.n11183 ASIG5V.n10031 2.24164
R45998 ASIG5V.n10356 ASIG5V.n10080 2.24164
R45999 ASIG5V.n11183 ASIG5V.n10030 2.24164
R46000 ASIG5V.n10356 ASIG5V.n10079 2.24164
R46001 ASIG5V.n11183 ASIG5V.n10029 2.24164
R46002 ASIG5V.n10356 ASIG5V.n10078 2.24164
R46003 ASIG5V.n11183 ASIG5V.n10028 2.24164
R46004 ASIG5V.n10356 ASIG5V.n10077 2.24164
R46005 ASIG5V.n11183 ASIG5V.n10027 2.24164
R46006 ASIG5V.n10357 ASIG5V.n10356 2.24164
R46007 ASIG5V.n11183 ASIG5V.n10026 2.24164
R46008 ASIG5V.n10356 ASIG5V.n10070 2.24164
R46009 ASIG5V.n11234 ASIG5V.n9966 2.24164
R46010 ASIG5V.n11485 ASIG5V.n10014 2.24164
R46011 ASIG5V.n11243 ASIG5V.n9966 2.24164
R46012 ASIG5V.n11485 ASIG5V.n10013 2.24164
R46013 ASIG5V.n11247 ASIG5V.n9966 2.24164
R46014 ASIG5V.n11485 ASIG5V.n10012 2.24164
R46015 ASIG5V.n11255 ASIG5V.n9966 2.24164
R46016 ASIG5V.n11485 ASIG5V.n10011 2.24164
R46017 ASIG5V.n11259 ASIG5V.n9966 2.24164
R46018 ASIG5V.n11485 ASIG5V.n10010 2.24164
R46019 ASIG5V.n11267 ASIG5V.n9966 2.24164
R46020 ASIG5V.n11485 ASIG5V.n10009 2.24164
R46021 ASIG5V.n11271 ASIG5V.n9966 2.24164
R46022 ASIG5V.n11485 ASIG5V.n10008 2.24164
R46023 ASIG5V.n11279 ASIG5V.n9966 2.24164
R46024 ASIG5V.n11485 ASIG5V.n10007 2.24164
R46025 ASIG5V.n11283 ASIG5V.n9966 2.24164
R46026 ASIG5V.n11485 ASIG5V.n10006 2.24164
R46027 ASIG5V.n11291 ASIG5V.n9966 2.24164
R46028 ASIG5V.n11485 ASIG5V.n10005 2.24164
R46029 ASIG5V.n11295 ASIG5V.n9966 2.24164
R46030 ASIG5V.n11485 ASIG5V.n10004 2.24164
R46031 ASIG5V.n11303 ASIG5V.n9966 2.24164
R46032 ASIG5V.n11485 ASIG5V.n10003 2.24164
R46033 ASIG5V.n11307 ASIG5V.n9966 2.24164
R46034 ASIG5V.n11485 ASIG5V.n10002 2.24164
R46035 ASIG5V.n11315 ASIG5V.n9966 2.24164
R46036 ASIG5V.n11485 ASIG5V.n10001 2.24164
R46037 ASIG5V.n11319 ASIG5V.n9966 2.24164
R46038 ASIG5V.n11485 ASIG5V.n10000 2.24164
R46039 ASIG5V.n11327 ASIG5V.n9966 2.24164
R46040 ASIG5V.n11485 ASIG5V.n9999 2.24164
R46041 ASIG5V.n11331 ASIG5V.n9966 2.24164
R46042 ASIG5V.n11485 ASIG5V.n9998 2.24164
R46043 ASIG5V.n11339 ASIG5V.n9966 2.24164
R46044 ASIG5V.n11485 ASIG5V.n9997 2.24164
R46045 ASIG5V.n11343 ASIG5V.n9966 2.24164
R46046 ASIG5V.n11485 ASIG5V.n9996 2.24164
R46047 ASIG5V.n11351 ASIG5V.n9966 2.24164
R46048 ASIG5V.n11485 ASIG5V.n9995 2.24164
R46049 ASIG5V.n11355 ASIG5V.n9966 2.24164
R46050 ASIG5V.n11485 ASIG5V.n9994 2.24164
R46051 ASIG5V.n11363 ASIG5V.n9966 2.24164
R46052 ASIG5V.n11485 ASIG5V.n9993 2.24164
R46053 ASIG5V.n11367 ASIG5V.n9966 2.24164
R46054 ASIG5V.n11485 ASIG5V.n9992 2.24164
R46055 ASIG5V.n11375 ASIG5V.n9966 2.24164
R46056 ASIG5V.n11485 ASIG5V.n9991 2.24164
R46057 ASIG5V.n11379 ASIG5V.n9966 2.24164
R46058 ASIG5V.n11485 ASIG5V.n9990 2.24164
R46059 ASIG5V.n11387 ASIG5V.n9966 2.24164
R46060 ASIG5V.n11485 ASIG5V.n9989 2.24164
R46061 ASIG5V.n11391 ASIG5V.n9966 2.24164
R46062 ASIG5V.n11485 ASIG5V.n9988 2.24164
R46063 ASIG5V.n11399 ASIG5V.n9966 2.24164
R46064 ASIG5V.n11485 ASIG5V.n9987 2.24164
R46065 ASIG5V.n11403 ASIG5V.n9966 2.24164
R46066 ASIG5V.n11485 ASIG5V.n9986 2.24164
R46067 ASIG5V.n11411 ASIG5V.n9966 2.24164
R46068 ASIG5V.n11485 ASIG5V.n9985 2.24164
R46069 ASIG5V.n11415 ASIG5V.n9966 2.24164
R46070 ASIG5V.n11485 ASIG5V.n9984 2.24164
R46071 ASIG5V.n11423 ASIG5V.n9966 2.24164
R46072 ASIG5V.n11485 ASIG5V.n9983 2.24164
R46073 ASIG5V.n11427 ASIG5V.n9966 2.24164
R46074 ASIG5V.n11485 ASIG5V.n9982 2.24164
R46075 ASIG5V.n11435 ASIG5V.n9966 2.24164
R46076 ASIG5V.n11485 ASIG5V.n9981 2.24164
R46077 ASIG5V.n11439 ASIG5V.n9966 2.24164
R46078 ASIG5V.n11485 ASIG5V.n9980 2.24164
R46079 ASIG5V.n11447 ASIG5V.n9966 2.24164
R46080 ASIG5V.n11485 ASIG5V.n9979 2.24164
R46081 ASIG5V.n11451 ASIG5V.n9966 2.24164
R46082 ASIG5V.n11485 ASIG5V.n9978 2.24164
R46083 ASIG5V.n11459 ASIG5V.n9966 2.24164
R46084 ASIG5V.n11485 ASIG5V.n9977 2.24164
R46085 ASIG5V.n11463 ASIG5V.n9966 2.24164
R46086 ASIG5V.n11485 ASIG5V.n9976 2.24164
R46087 ASIG5V.n11471 ASIG5V.n9966 2.24164
R46088 ASIG5V.n11485 ASIG5V.n9975 2.24164
R46089 ASIG5V.n11475 ASIG5V.n9966 2.24164
R46090 ASIG5V.n11485 ASIG5V.n9974 2.24164
R46091 ASIG5V.n11483 ASIG5V.n9966 2.24164
R46092 ASIG5V.n2999 ASIG5V.n2958 2.24164
R46093 ASIG5V.n11751 ASIG5V.n2954 2.24164
R46094 ASIG5V.n11509 ASIG5V.n2958 2.24164
R46095 ASIG5V.n11751 ASIG5V.n2953 2.24164
R46096 ASIG5V.n11513 ASIG5V.n2958 2.24164
R46097 ASIG5V.n11751 ASIG5V.n2952 2.24164
R46098 ASIG5V.n11521 ASIG5V.n2958 2.24164
R46099 ASIG5V.n11751 ASIG5V.n2951 2.24164
R46100 ASIG5V.n11525 ASIG5V.n2958 2.24164
R46101 ASIG5V.n11751 ASIG5V.n2950 2.24164
R46102 ASIG5V.n11533 ASIG5V.n2958 2.24164
R46103 ASIG5V.n11751 ASIG5V.n2949 2.24164
R46104 ASIG5V.n11537 ASIG5V.n2958 2.24164
R46105 ASIG5V.n11751 ASIG5V.n2948 2.24164
R46106 ASIG5V.n11545 ASIG5V.n2958 2.24164
R46107 ASIG5V.n11751 ASIG5V.n2947 2.24164
R46108 ASIG5V.n11549 ASIG5V.n2958 2.24164
R46109 ASIG5V.n11751 ASIG5V.n2946 2.24164
R46110 ASIG5V.n11557 ASIG5V.n2958 2.24164
R46111 ASIG5V.n11751 ASIG5V.n2945 2.24164
R46112 ASIG5V.n11561 ASIG5V.n2958 2.24164
R46113 ASIG5V.n11751 ASIG5V.n2944 2.24164
R46114 ASIG5V.n11569 ASIG5V.n2958 2.24164
R46115 ASIG5V.n11751 ASIG5V.n2943 2.24164
R46116 ASIG5V.n11573 ASIG5V.n2958 2.24164
R46117 ASIG5V.n11751 ASIG5V.n2942 2.24164
R46118 ASIG5V.n11581 ASIG5V.n2958 2.24164
R46119 ASIG5V.n11751 ASIG5V.n2941 2.24164
R46120 ASIG5V.n11585 ASIG5V.n2958 2.24164
R46121 ASIG5V.n11751 ASIG5V.n2940 2.24164
R46122 ASIG5V.n11593 ASIG5V.n2958 2.24164
R46123 ASIG5V.n11751 ASIG5V.n2939 2.24164
R46124 ASIG5V.n11597 ASIG5V.n2958 2.24164
R46125 ASIG5V.n11751 ASIG5V.n2938 2.24164
R46126 ASIG5V.n11605 ASIG5V.n2958 2.24164
R46127 ASIG5V.n11751 ASIG5V.n2937 2.24164
R46128 ASIG5V.n11609 ASIG5V.n2958 2.24164
R46129 ASIG5V.n11751 ASIG5V.n2936 2.24164
R46130 ASIG5V.n11617 ASIG5V.n2958 2.24164
R46131 ASIG5V.n11751 ASIG5V.n2935 2.24164
R46132 ASIG5V.n11621 ASIG5V.n2958 2.24164
R46133 ASIG5V.n11751 ASIG5V.n2934 2.24164
R46134 ASIG5V.n11629 ASIG5V.n2958 2.24164
R46135 ASIG5V.n11751 ASIG5V.n2933 2.24164
R46136 ASIG5V.n11633 ASIG5V.n2958 2.24164
R46137 ASIG5V.n11751 ASIG5V.n2932 2.24164
R46138 ASIG5V.n11641 ASIG5V.n2958 2.24164
R46139 ASIG5V.n11751 ASIG5V.n2931 2.24164
R46140 ASIG5V.n11645 ASIG5V.n2958 2.24164
R46141 ASIG5V.n11751 ASIG5V.n2930 2.24164
R46142 ASIG5V.n11653 ASIG5V.n2958 2.24164
R46143 ASIG5V.n11751 ASIG5V.n2929 2.24164
R46144 ASIG5V.n11657 ASIG5V.n2958 2.24164
R46145 ASIG5V.n11751 ASIG5V.n2928 2.24164
R46146 ASIG5V.n11665 ASIG5V.n2958 2.24164
R46147 ASIG5V.n11751 ASIG5V.n2927 2.24164
R46148 ASIG5V.n11669 ASIG5V.n2958 2.24164
R46149 ASIG5V.n11751 ASIG5V.n2926 2.24164
R46150 ASIG5V.n11677 ASIG5V.n2958 2.24164
R46151 ASIG5V.n11751 ASIG5V.n2925 2.24164
R46152 ASIG5V.n11681 ASIG5V.n2958 2.24164
R46153 ASIG5V.n11751 ASIG5V.n2924 2.24164
R46154 ASIG5V.n11689 ASIG5V.n2958 2.24164
R46155 ASIG5V.n11751 ASIG5V.n2923 2.24164
R46156 ASIG5V.n11693 ASIG5V.n2958 2.24164
R46157 ASIG5V.n11751 ASIG5V.n2922 2.24164
R46158 ASIG5V.n11701 ASIG5V.n2958 2.24164
R46159 ASIG5V.n11751 ASIG5V.n2921 2.24164
R46160 ASIG5V.n11705 ASIG5V.n2958 2.24164
R46161 ASIG5V.n11751 ASIG5V.n2920 2.24164
R46162 ASIG5V.n11713 ASIG5V.n2958 2.24164
R46163 ASIG5V.n11751 ASIG5V.n2919 2.24164
R46164 ASIG5V.n11717 ASIG5V.n2958 2.24164
R46165 ASIG5V.n11751 ASIG5V.n2918 2.24164
R46166 ASIG5V.n11725 ASIG5V.n2958 2.24164
R46167 ASIG5V.n11751 ASIG5V.n2917 2.24164
R46168 ASIG5V.n11729 ASIG5V.n2958 2.24164
R46169 ASIG5V.n11751 ASIG5V.n2916 2.24164
R46170 ASIG5V.n11737 ASIG5V.n2958 2.24164
R46171 ASIG5V.n11751 ASIG5V.n2915 2.24164
R46172 ASIG5V.n11741 ASIG5V.n2958 2.24164
R46173 ASIG5V.n11751 ASIG5V.n2914 2.24164
R46174 ASIG5V.n11749 ASIG5V.n2958 2.24164
R46175 ASIG5V.n2658 ASIG5V.n2616 2.24164
R46176 ASIG5V.n11771 ASIG5V.n2610 2.24164
R46177 ASIG5V.n2665 ASIG5V.n2616 2.24164
R46178 ASIG5V.n11771 ASIG5V.n2609 2.24164
R46179 ASIG5V.n2669 ASIG5V.n2616 2.24164
R46180 ASIG5V.n11771 ASIG5V.n2608 2.24164
R46181 ASIG5V.n2677 ASIG5V.n2616 2.24164
R46182 ASIG5V.n11771 ASIG5V.n2607 2.24164
R46183 ASIG5V.n2681 ASIG5V.n2616 2.24164
R46184 ASIG5V.n11771 ASIG5V.n2606 2.24164
R46185 ASIG5V.n2689 ASIG5V.n2616 2.24164
R46186 ASIG5V.n11771 ASIG5V.n2605 2.24164
R46187 ASIG5V.n2693 ASIG5V.n2616 2.24164
R46188 ASIG5V.n11771 ASIG5V.n2604 2.24164
R46189 ASIG5V.n2701 ASIG5V.n2616 2.24164
R46190 ASIG5V.n11771 ASIG5V.n2603 2.24164
R46191 ASIG5V.n2705 ASIG5V.n2616 2.24164
R46192 ASIG5V.n11771 ASIG5V.n2602 2.24164
R46193 ASIG5V.n2713 ASIG5V.n2616 2.24164
R46194 ASIG5V.n11771 ASIG5V.n2601 2.24164
R46195 ASIG5V.n2717 ASIG5V.n2616 2.24164
R46196 ASIG5V.n11771 ASIG5V.n2600 2.24164
R46197 ASIG5V.n2725 ASIG5V.n2616 2.24164
R46198 ASIG5V.n11771 ASIG5V.n2599 2.24164
R46199 ASIG5V.n2729 ASIG5V.n2616 2.24164
R46200 ASIG5V.n11771 ASIG5V.n2598 2.24164
R46201 ASIG5V.n2737 ASIG5V.n2616 2.24164
R46202 ASIG5V.n11771 ASIG5V.n2597 2.24164
R46203 ASIG5V.n2741 ASIG5V.n2616 2.24164
R46204 ASIG5V.n11771 ASIG5V.n2596 2.24164
R46205 ASIG5V.n2749 ASIG5V.n2616 2.24164
R46206 ASIG5V.n11771 ASIG5V.n2595 2.24164
R46207 ASIG5V.n2753 ASIG5V.n2616 2.24164
R46208 ASIG5V.n11771 ASIG5V.n2594 2.24164
R46209 ASIG5V.n2761 ASIG5V.n2616 2.24164
R46210 ASIG5V.n11771 ASIG5V.n2593 2.24164
R46211 ASIG5V.n2765 ASIG5V.n2616 2.24164
R46212 ASIG5V.n11771 ASIG5V.n2592 2.24164
R46213 ASIG5V.n2773 ASIG5V.n2616 2.24164
R46214 ASIG5V.n11771 ASIG5V.n2591 2.24164
R46215 ASIG5V.n2777 ASIG5V.n2616 2.24164
R46216 ASIG5V.n11771 ASIG5V.n2590 2.24164
R46217 ASIG5V.n2785 ASIG5V.n2616 2.24164
R46218 ASIG5V.n11771 ASIG5V.n2589 2.24164
R46219 ASIG5V.n2789 ASIG5V.n2616 2.24164
R46220 ASIG5V.n11771 ASIG5V.n2588 2.24164
R46221 ASIG5V.n2797 ASIG5V.n2616 2.24164
R46222 ASIG5V.n11771 ASIG5V.n2587 2.24164
R46223 ASIG5V.n2801 ASIG5V.n2616 2.24164
R46224 ASIG5V.n11771 ASIG5V.n2586 2.24164
R46225 ASIG5V.n2809 ASIG5V.n2616 2.24164
R46226 ASIG5V.n11771 ASIG5V.n2585 2.24164
R46227 ASIG5V.n2813 ASIG5V.n2616 2.24164
R46228 ASIG5V.n11771 ASIG5V.n2584 2.24164
R46229 ASIG5V.n2821 ASIG5V.n2616 2.24164
R46230 ASIG5V.n11771 ASIG5V.n2583 2.24164
R46231 ASIG5V.n2825 ASIG5V.n2616 2.24164
R46232 ASIG5V.n11771 ASIG5V.n2582 2.24164
R46233 ASIG5V.n2833 ASIG5V.n2616 2.24164
R46234 ASIG5V.n11771 ASIG5V.n2581 2.24164
R46235 ASIG5V.n2837 ASIG5V.n2616 2.24164
R46236 ASIG5V.n11771 ASIG5V.n2580 2.24164
R46237 ASIG5V.n2845 ASIG5V.n2616 2.24164
R46238 ASIG5V.n11771 ASIG5V.n2579 2.24164
R46239 ASIG5V.n2849 ASIG5V.n2616 2.24164
R46240 ASIG5V.n11771 ASIG5V.n2578 2.24164
R46241 ASIG5V.n2857 ASIG5V.n2616 2.24164
R46242 ASIG5V.n11771 ASIG5V.n2577 2.24164
R46243 ASIG5V.n2861 ASIG5V.n2616 2.24164
R46244 ASIG5V.n11771 ASIG5V.n2576 2.24164
R46245 ASIG5V.n2869 ASIG5V.n2616 2.24164
R46246 ASIG5V.n11771 ASIG5V.n2575 2.24164
R46247 ASIG5V.n2873 ASIG5V.n2616 2.24164
R46248 ASIG5V.n11771 ASIG5V.n2574 2.24164
R46249 ASIG5V.n2881 ASIG5V.n2616 2.24164
R46250 ASIG5V.n11771 ASIG5V.n2573 2.24164
R46251 ASIG5V.n2885 ASIG5V.n2616 2.24164
R46252 ASIG5V.n11771 ASIG5V.n2572 2.24164
R46253 ASIG5V.n2893 ASIG5V.n2616 2.24164
R46254 ASIG5V.n11771 ASIG5V.n2571 2.24164
R46255 ASIG5V.n2897 ASIG5V.n2616 2.24164
R46256 ASIG5V.n11771 ASIG5V.n2570 2.24164
R46257 ASIG5V.n11769 ASIG5V.n2616 2.24164
R46258 ASIG5V.n2306 ASIG5V.n2221 2.24164
R46259 ASIG5V.n2555 ASIG5V.n2262 2.24164
R46260 ASIG5V.n2313 ASIG5V.n2221 2.24164
R46261 ASIG5V.n2555 ASIG5V.n2261 2.24164
R46262 ASIG5V.n2317 ASIG5V.n2221 2.24164
R46263 ASIG5V.n2555 ASIG5V.n2260 2.24164
R46264 ASIG5V.n2325 ASIG5V.n2221 2.24164
R46265 ASIG5V.n2555 ASIG5V.n2259 2.24164
R46266 ASIG5V.n2329 ASIG5V.n2221 2.24164
R46267 ASIG5V.n2555 ASIG5V.n2258 2.24164
R46268 ASIG5V.n2337 ASIG5V.n2221 2.24164
R46269 ASIG5V.n2555 ASIG5V.n2257 2.24164
R46270 ASIG5V.n2341 ASIG5V.n2221 2.24164
R46271 ASIG5V.n2555 ASIG5V.n2256 2.24164
R46272 ASIG5V.n2349 ASIG5V.n2221 2.24164
R46273 ASIG5V.n2555 ASIG5V.n2255 2.24164
R46274 ASIG5V.n2353 ASIG5V.n2221 2.24164
R46275 ASIG5V.n2555 ASIG5V.n2254 2.24164
R46276 ASIG5V.n2361 ASIG5V.n2221 2.24164
R46277 ASIG5V.n2555 ASIG5V.n2253 2.24164
R46278 ASIG5V.n2365 ASIG5V.n2221 2.24164
R46279 ASIG5V.n2555 ASIG5V.n2252 2.24164
R46280 ASIG5V.n2373 ASIG5V.n2221 2.24164
R46281 ASIG5V.n2555 ASIG5V.n2251 2.24164
R46282 ASIG5V.n2377 ASIG5V.n2221 2.24164
R46283 ASIG5V.n2555 ASIG5V.n2250 2.24164
R46284 ASIG5V.n2385 ASIG5V.n2221 2.24164
R46285 ASIG5V.n2555 ASIG5V.n2249 2.24164
R46286 ASIG5V.n2389 ASIG5V.n2221 2.24164
R46287 ASIG5V.n2555 ASIG5V.n2248 2.24164
R46288 ASIG5V.n2397 ASIG5V.n2221 2.24164
R46289 ASIG5V.n2555 ASIG5V.n2247 2.24164
R46290 ASIG5V.n2401 ASIG5V.n2221 2.24164
R46291 ASIG5V.n2555 ASIG5V.n2246 2.24164
R46292 ASIG5V.n2409 ASIG5V.n2221 2.24164
R46293 ASIG5V.n2555 ASIG5V.n2245 2.24164
R46294 ASIG5V.n2413 ASIG5V.n2221 2.24164
R46295 ASIG5V.n2555 ASIG5V.n2244 2.24164
R46296 ASIG5V.n2421 ASIG5V.n2221 2.24164
R46297 ASIG5V.n2555 ASIG5V.n2243 2.24164
R46298 ASIG5V.n2425 ASIG5V.n2221 2.24164
R46299 ASIG5V.n2555 ASIG5V.n2242 2.24164
R46300 ASIG5V.n2433 ASIG5V.n2221 2.24164
R46301 ASIG5V.n2555 ASIG5V.n2241 2.24164
R46302 ASIG5V.n2437 ASIG5V.n2221 2.24164
R46303 ASIG5V.n2555 ASIG5V.n2240 2.24164
R46304 ASIG5V.n2445 ASIG5V.n2221 2.24164
R46305 ASIG5V.n2555 ASIG5V.n2239 2.24164
R46306 ASIG5V.n2449 ASIG5V.n2221 2.24164
R46307 ASIG5V.n2555 ASIG5V.n2238 2.24164
R46308 ASIG5V.n2457 ASIG5V.n2221 2.24164
R46309 ASIG5V.n2555 ASIG5V.n2237 2.24164
R46310 ASIG5V.n2461 ASIG5V.n2221 2.24164
R46311 ASIG5V.n2555 ASIG5V.n2236 2.24164
R46312 ASIG5V.n2469 ASIG5V.n2221 2.24164
R46313 ASIG5V.n2555 ASIG5V.n2235 2.24164
R46314 ASIG5V.n2473 ASIG5V.n2221 2.24164
R46315 ASIG5V.n2555 ASIG5V.n2234 2.24164
R46316 ASIG5V.n2481 ASIG5V.n2221 2.24164
R46317 ASIG5V.n2555 ASIG5V.n2233 2.24164
R46318 ASIG5V.n2485 ASIG5V.n2221 2.24164
R46319 ASIG5V.n2555 ASIG5V.n2232 2.24164
R46320 ASIG5V.n2493 ASIG5V.n2221 2.24164
R46321 ASIG5V.n2555 ASIG5V.n2231 2.24164
R46322 ASIG5V.n2497 ASIG5V.n2221 2.24164
R46323 ASIG5V.n2555 ASIG5V.n2230 2.24164
R46324 ASIG5V.n2505 ASIG5V.n2221 2.24164
R46325 ASIG5V.n2555 ASIG5V.n2229 2.24164
R46326 ASIG5V.n2509 ASIG5V.n2221 2.24164
R46327 ASIG5V.n2555 ASIG5V.n2228 2.24164
R46328 ASIG5V.n2517 ASIG5V.n2221 2.24164
R46329 ASIG5V.n2555 ASIG5V.n2227 2.24164
R46330 ASIG5V.n2521 ASIG5V.n2221 2.24164
R46331 ASIG5V.n2555 ASIG5V.n2226 2.24164
R46332 ASIG5V.n2529 ASIG5V.n2221 2.24164
R46333 ASIG5V.n2555 ASIG5V.n2225 2.24164
R46334 ASIG5V.n2533 ASIG5V.n2221 2.24164
R46335 ASIG5V.n2555 ASIG5V.n2224 2.24164
R46336 ASIG5V.n2541 ASIG5V.n2221 2.24164
R46337 ASIG5V.n2555 ASIG5V.n2223 2.24164
R46338 ASIG5V.n2545 ASIG5V.n2221 2.24164
R46339 ASIG5V.n2555 ASIG5V.n2222 2.24164
R46340 ASIG5V.n2553 ASIG5V.n2221 2.24164
R46341 ASIG5V.n1949 ASIG5V.n1864 2.24164
R46342 ASIG5V.n2198 ASIG5V.n1905 2.24164
R46343 ASIG5V.n1956 ASIG5V.n1864 2.24164
R46344 ASIG5V.n2198 ASIG5V.n1904 2.24164
R46345 ASIG5V.n1960 ASIG5V.n1864 2.24164
R46346 ASIG5V.n2198 ASIG5V.n1903 2.24164
R46347 ASIG5V.n1968 ASIG5V.n1864 2.24164
R46348 ASIG5V.n2198 ASIG5V.n1902 2.24164
R46349 ASIG5V.n1972 ASIG5V.n1864 2.24164
R46350 ASIG5V.n2198 ASIG5V.n1901 2.24164
R46351 ASIG5V.n1980 ASIG5V.n1864 2.24164
R46352 ASIG5V.n2198 ASIG5V.n1900 2.24164
R46353 ASIG5V.n1984 ASIG5V.n1864 2.24164
R46354 ASIG5V.n2198 ASIG5V.n1899 2.24164
R46355 ASIG5V.n1992 ASIG5V.n1864 2.24164
R46356 ASIG5V.n2198 ASIG5V.n1898 2.24164
R46357 ASIG5V.n1996 ASIG5V.n1864 2.24164
R46358 ASIG5V.n2198 ASIG5V.n1897 2.24164
R46359 ASIG5V.n2004 ASIG5V.n1864 2.24164
R46360 ASIG5V.n2198 ASIG5V.n1896 2.24164
R46361 ASIG5V.n2008 ASIG5V.n1864 2.24164
R46362 ASIG5V.n2198 ASIG5V.n1895 2.24164
R46363 ASIG5V.n2016 ASIG5V.n1864 2.24164
R46364 ASIG5V.n2198 ASIG5V.n1894 2.24164
R46365 ASIG5V.n2020 ASIG5V.n1864 2.24164
R46366 ASIG5V.n2198 ASIG5V.n1893 2.24164
R46367 ASIG5V.n2028 ASIG5V.n1864 2.24164
R46368 ASIG5V.n2198 ASIG5V.n1892 2.24164
R46369 ASIG5V.n2032 ASIG5V.n1864 2.24164
R46370 ASIG5V.n2198 ASIG5V.n1891 2.24164
R46371 ASIG5V.n2040 ASIG5V.n1864 2.24164
R46372 ASIG5V.n2198 ASIG5V.n1890 2.24164
R46373 ASIG5V.n2044 ASIG5V.n1864 2.24164
R46374 ASIG5V.n2198 ASIG5V.n1889 2.24164
R46375 ASIG5V.n2052 ASIG5V.n1864 2.24164
R46376 ASIG5V.n2198 ASIG5V.n1888 2.24164
R46377 ASIG5V.n2056 ASIG5V.n1864 2.24164
R46378 ASIG5V.n2198 ASIG5V.n1887 2.24164
R46379 ASIG5V.n2064 ASIG5V.n1864 2.24164
R46380 ASIG5V.n2198 ASIG5V.n1886 2.24164
R46381 ASIG5V.n2068 ASIG5V.n1864 2.24164
R46382 ASIG5V.n2198 ASIG5V.n1885 2.24164
R46383 ASIG5V.n2076 ASIG5V.n1864 2.24164
R46384 ASIG5V.n2198 ASIG5V.n1884 2.24164
R46385 ASIG5V.n2080 ASIG5V.n1864 2.24164
R46386 ASIG5V.n2198 ASIG5V.n1883 2.24164
R46387 ASIG5V.n2088 ASIG5V.n1864 2.24164
R46388 ASIG5V.n2198 ASIG5V.n1882 2.24164
R46389 ASIG5V.n2092 ASIG5V.n1864 2.24164
R46390 ASIG5V.n2198 ASIG5V.n1881 2.24164
R46391 ASIG5V.n2100 ASIG5V.n1864 2.24164
R46392 ASIG5V.n2198 ASIG5V.n1880 2.24164
R46393 ASIG5V.n2104 ASIG5V.n1864 2.24164
R46394 ASIG5V.n2198 ASIG5V.n1879 2.24164
R46395 ASIG5V.n2112 ASIG5V.n1864 2.24164
R46396 ASIG5V.n2198 ASIG5V.n1878 2.24164
R46397 ASIG5V.n2116 ASIG5V.n1864 2.24164
R46398 ASIG5V.n2198 ASIG5V.n1877 2.24164
R46399 ASIG5V.n2124 ASIG5V.n1864 2.24164
R46400 ASIG5V.n2198 ASIG5V.n1876 2.24164
R46401 ASIG5V.n2128 ASIG5V.n1864 2.24164
R46402 ASIG5V.n2198 ASIG5V.n1875 2.24164
R46403 ASIG5V.n2136 ASIG5V.n1864 2.24164
R46404 ASIG5V.n2198 ASIG5V.n1874 2.24164
R46405 ASIG5V.n2140 ASIG5V.n1864 2.24164
R46406 ASIG5V.n2198 ASIG5V.n1873 2.24164
R46407 ASIG5V.n2148 ASIG5V.n1864 2.24164
R46408 ASIG5V.n2198 ASIG5V.n1872 2.24164
R46409 ASIG5V.n2152 ASIG5V.n1864 2.24164
R46410 ASIG5V.n2198 ASIG5V.n1871 2.24164
R46411 ASIG5V.n2160 ASIG5V.n1864 2.24164
R46412 ASIG5V.n2198 ASIG5V.n1870 2.24164
R46413 ASIG5V.n2164 ASIG5V.n1864 2.24164
R46414 ASIG5V.n2198 ASIG5V.n1869 2.24164
R46415 ASIG5V.n2172 ASIG5V.n1864 2.24164
R46416 ASIG5V.n2198 ASIG5V.n1868 2.24164
R46417 ASIG5V.n2176 ASIG5V.n1864 2.24164
R46418 ASIG5V.n2198 ASIG5V.n1867 2.24164
R46419 ASIG5V.n2184 ASIG5V.n1864 2.24164
R46420 ASIG5V.n2198 ASIG5V.n1866 2.24164
R46421 ASIG5V.n2188 ASIG5V.n1864 2.24164
R46422 ASIG5V.n2198 ASIG5V.n1865 2.24164
R46423 ASIG5V.n2196 ASIG5V.n1864 2.24164
R46424 ASIG5V.n11997 ASIG5V.n11996 2.24164
R46425 ASIG5V.n11994 ASIG5V.n1762 2.24164
R46426 ASIG5V.n11997 ASIG5V.n1716 2.24164
R46427 ASIG5V.n11994 ASIG5V.n1761 2.24164
R46428 ASIG5V.n11997 ASIG5V.n1715 2.24164
R46429 ASIG5V.n11994 ASIG5V.n1760 2.24164
R46430 ASIG5V.n11997 ASIG5V.n1714 2.24164
R46431 ASIG5V.n11994 ASIG5V.n1759 2.24164
R46432 ASIG5V.n11997 ASIG5V.n1713 2.24164
R46433 ASIG5V.n11994 ASIG5V.n1758 2.24164
R46434 ASIG5V.n11997 ASIG5V.n1712 2.24164
R46435 ASIG5V.n11994 ASIG5V.n1757 2.24164
R46436 ASIG5V.n11997 ASIG5V.n1711 2.24164
R46437 ASIG5V.n11994 ASIG5V.n1756 2.24164
R46438 ASIG5V.n11997 ASIG5V.n1710 2.24164
R46439 ASIG5V.n11994 ASIG5V.n1755 2.24164
R46440 ASIG5V.n11997 ASIG5V.n1709 2.24164
R46441 ASIG5V.n11994 ASIG5V.n1754 2.24164
R46442 ASIG5V.n11997 ASIG5V.n1708 2.24164
R46443 ASIG5V.n11994 ASIG5V.n1753 2.24164
R46444 ASIG5V.n11997 ASIG5V.n1707 2.24164
R46445 ASIG5V.n11994 ASIG5V.n1752 2.24164
R46446 ASIG5V.n11997 ASIG5V.n1706 2.24164
R46447 ASIG5V.n11994 ASIG5V.n1751 2.24164
R46448 ASIG5V.n11997 ASIG5V.n1705 2.24164
R46449 ASIG5V.n11994 ASIG5V.n1750 2.24164
R46450 ASIG5V.n11997 ASIG5V.n1704 2.24164
R46451 ASIG5V.n11994 ASIG5V.n1749 2.24164
R46452 ASIG5V.n11997 ASIG5V.n1703 2.24164
R46453 ASIG5V.n11994 ASIG5V.n1748 2.24164
R46454 ASIG5V.n11997 ASIG5V.n1702 2.24164
R46455 ASIG5V.n11994 ASIG5V.n1747 2.24164
R46456 ASIG5V.n11997 ASIG5V.n1701 2.24164
R46457 ASIG5V.n11994 ASIG5V.n1746 2.24164
R46458 ASIG5V.n11997 ASIG5V.n1700 2.24164
R46459 ASIG5V.n11994 ASIG5V.n1745 2.24164
R46460 ASIG5V.n11997 ASIG5V.n1699 2.24164
R46461 ASIG5V.n11994 ASIG5V.n1744 2.24164
R46462 ASIG5V.n11997 ASIG5V.n1698 2.24164
R46463 ASIG5V.n11994 ASIG5V.n1743 2.24164
R46464 ASIG5V.n11997 ASIG5V.n1697 2.24164
R46465 ASIG5V.n11994 ASIG5V.n1742 2.24164
R46466 ASIG5V.n11997 ASIG5V.n1696 2.24164
R46467 ASIG5V.n11994 ASIG5V.n1741 2.24164
R46468 ASIG5V.n11997 ASIG5V.n1695 2.24164
R46469 ASIG5V.n11994 ASIG5V.n1740 2.24164
R46470 ASIG5V.n11997 ASIG5V.n1694 2.24164
R46471 ASIG5V.n11994 ASIG5V.n1739 2.24164
R46472 ASIG5V.n11997 ASIG5V.n1693 2.24164
R46473 ASIG5V.n11994 ASIG5V.n1738 2.24164
R46474 ASIG5V.n11997 ASIG5V.n1692 2.24164
R46475 ASIG5V.n11994 ASIG5V.n1737 2.24164
R46476 ASIG5V.n11997 ASIG5V.n1691 2.24164
R46477 ASIG5V.n11994 ASIG5V.n1736 2.24164
R46478 ASIG5V.n11997 ASIG5V.n1690 2.24164
R46479 ASIG5V.n11994 ASIG5V.n1735 2.24164
R46480 ASIG5V.n11997 ASIG5V.n1689 2.24164
R46481 ASIG5V.n11994 ASIG5V.n1734 2.24164
R46482 ASIG5V.n11997 ASIG5V.n1688 2.24164
R46483 ASIG5V.n11994 ASIG5V.n1733 2.24164
R46484 ASIG5V.n11997 ASIG5V.n1687 2.24164
R46485 ASIG5V.n11994 ASIG5V.n1732 2.24164
R46486 ASIG5V.n11997 ASIG5V.n1686 2.24164
R46487 ASIG5V.n11994 ASIG5V.n1731 2.24164
R46488 ASIG5V.n11997 ASIG5V.n1685 2.24164
R46489 ASIG5V.n11994 ASIG5V.n1730 2.24164
R46490 ASIG5V.n11997 ASIG5V.n1684 2.24164
R46491 ASIG5V.n11994 ASIG5V.n1729 2.24164
R46492 ASIG5V.n11997 ASIG5V.n1683 2.24164
R46493 ASIG5V.n11994 ASIG5V.n1728 2.24164
R46494 ASIG5V.n11997 ASIG5V.n1682 2.24164
R46495 ASIG5V.n11994 ASIG5V.n1727 2.24164
R46496 ASIG5V.n11997 ASIG5V.n1681 2.24164
R46497 ASIG5V.n11994 ASIG5V.n1726 2.24164
R46498 ASIG5V.n11997 ASIG5V.n1680 2.24164
R46499 ASIG5V.n11994 ASIG5V.n1725 2.24164
R46500 ASIG5V.n11997 ASIG5V.n1679 2.24164
R46501 ASIG5V.n11994 ASIG5V.n1724 2.24164
R46502 ASIG5V.n11997 ASIG5V.n1678 2.24164
R46503 ASIG5V.n11994 ASIG5V.n1723 2.24164
R46504 ASIG5V.n11997 ASIG5V.n1677 2.24164
R46505 ASIG5V.n11994 ASIG5V.n1722 2.24164
R46506 ASIG5V.n11997 ASIG5V.n1676 2.24164
R46507 ASIG5V.n12011 ASIG5V.n12010 2.24164
R46508 ASIG5V.n12008 ASIG5V.n1414 2.24164
R46509 ASIG5V.n12011 ASIG5V.n1369 2.24164
R46510 ASIG5V.n12008 ASIG5V.n1413 2.24164
R46511 ASIG5V.n12011 ASIG5V.n1368 2.24164
R46512 ASIG5V.n12008 ASIG5V.n1412 2.24164
R46513 ASIG5V.n12011 ASIG5V.n1367 2.24164
R46514 ASIG5V.n12008 ASIG5V.n1411 2.24164
R46515 ASIG5V.n12011 ASIG5V.n1366 2.24164
R46516 ASIG5V.n12008 ASIG5V.n1410 2.24164
R46517 ASIG5V.n12011 ASIG5V.n1365 2.24164
R46518 ASIG5V.n12008 ASIG5V.n1409 2.24164
R46519 ASIG5V.n12011 ASIG5V.n1364 2.24164
R46520 ASIG5V.n12008 ASIG5V.n1408 2.24164
R46521 ASIG5V.n12011 ASIG5V.n1363 2.24164
R46522 ASIG5V.n12008 ASIG5V.n1407 2.24164
R46523 ASIG5V.n12011 ASIG5V.n1362 2.24164
R46524 ASIG5V.n12008 ASIG5V.n1406 2.24164
R46525 ASIG5V.n12011 ASIG5V.n1361 2.24164
R46526 ASIG5V.n12008 ASIG5V.n1405 2.24164
R46527 ASIG5V.n12011 ASIG5V.n1360 2.24164
R46528 ASIG5V.n12008 ASIG5V.n1404 2.24164
R46529 ASIG5V.n12011 ASIG5V.n1359 2.24164
R46530 ASIG5V.n12008 ASIG5V.n1403 2.24164
R46531 ASIG5V.n12011 ASIG5V.n1358 2.24164
R46532 ASIG5V.n12008 ASIG5V.n1402 2.24164
R46533 ASIG5V.n12011 ASIG5V.n1357 2.24164
R46534 ASIG5V.n12008 ASIG5V.n1401 2.24164
R46535 ASIG5V.n12011 ASIG5V.n1356 2.24164
R46536 ASIG5V.n12008 ASIG5V.n1400 2.24164
R46537 ASIG5V.n12011 ASIG5V.n1355 2.24164
R46538 ASIG5V.n12008 ASIG5V.n1399 2.24164
R46539 ASIG5V.n12011 ASIG5V.n1354 2.24164
R46540 ASIG5V.n12008 ASIG5V.n1398 2.24164
R46541 ASIG5V.n12011 ASIG5V.n1353 2.24164
R46542 ASIG5V.n12008 ASIG5V.n1397 2.24164
R46543 ASIG5V.n12011 ASIG5V.n1352 2.24164
R46544 ASIG5V.n12008 ASIG5V.n1396 2.24164
R46545 ASIG5V.n12011 ASIG5V.n1351 2.24164
R46546 ASIG5V.n12008 ASIG5V.n1395 2.24164
R46547 ASIG5V.n12011 ASIG5V.n1350 2.24164
R46548 ASIG5V.n12008 ASIG5V.n1394 2.24164
R46549 ASIG5V.n12011 ASIG5V.n1349 2.24164
R46550 ASIG5V.n12008 ASIG5V.n1393 2.24164
R46551 ASIG5V.n12011 ASIG5V.n1348 2.24164
R46552 ASIG5V.n12008 ASIG5V.n1392 2.24164
R46553 ASIG5V.n12011 ASIG5V.n1347 2.24164
R46554 ASIG5V.n12008 ASIG5V.n1391 2.24164
R46555 ASIG5V.n12011 ASIG5V.n1346 2.24164
R46556 ASIG5V.n12008 ASIG5V.n1390 2.24164
R46557 ASIG5V.n12011 ASIG5V.n1345 2.24164
R46558 ASIG5V.n12008 ASIG5V.n1389 2.24164
R46559 ASIG5V.n12011 ASIG5V.n1344 2.24164
R46560 ASIG5V.n12008 ASIG5V.n1388 2.24164
R46561 ASIG5V.n12011 ASIG5V.n1343 2.24164
R46562 ASIG5V.n12008 ASIG5V.n1387 2.24164
R46563 ASIG5V.n12011 ASIG5V.n1342 2.24164
R46564 ASIG5V.n12008 ASIG5V.n1386 2.24164
R46565 ASIG5V.n12011 ASIG5V.n1341 2.24164
R46566 ASIG5V.n12008 ASIG5V.n1385 2.24164
R46567 ASIG5V.n12011 ASIG5V.n1340 2.24164
R46568 ASIG5V.n12008 ASIG5V.n1384 2.24164
R46569 ASIG5V.n12011 ASIG5V.n1339 2.24164
R46570 ASIG5V.n12008 ASIG5V.n1383 2.24164
R46571 ASIG5V.n12011 ASIG5V.n1338 2.24164
R46572 ASIG5V.n12008 ASIG5V.n1382 2.24164
R46573 ASIG5V.n12011 ASIG5V.n1337 2.24164
R46574 ASIG5V.n12008 ASIG5V.n1381 2.24164
R46575 ASIG5V.n12011 ASIG5V.n1336 2.24164
R46576 ASIG5V.n12008 ASIG5V.n1380 2.24164
R46577 ASIG5V.n12011 ASIG5V.n1335 2.24164
R46578 ASIG5V.n12008 ASIG5V.n1379 2.24164
R46579 ASIG5V.n12011 ASIG5V.n1334 2.24164
R46580 ASIG5V.n12008 ASIG5V.n1378 2.24164
R46581 ASIG5V.n12011 ASIG5V.n1333 2.24164
R46582 ASIG5V.n12008 ASIG5V.n1377 2.24164
R46583 ASIG5V.n12011 ASIG5V.n1332 2.24164
R46584 ASIG5V.n12008 ASIG5V.n1376 2.24164
R46585 ASIG5V.n12011 ASIG5V.n1331 2.24164
R46586 ASIG5V.n12008 ASIG5V.n1375 2.24164
R46587 ASIG5V.n12011 ASIG5V.n1330 2.24164
R46588 ASIG5V.n12008 ASIG5V.n1374 2.24164
R46589 ASIG5V.n12011 ASIG5V.n1329 2.24164
R46590 ASIG5V.n1313 ASIG5V.n1272 2.24164
R46591 ASIG5V.n12268 ASIG5V.n1267 2.24164
R46592 ASIG5V.n12026 ASIG5V.n1272 2.24164
R46593 ASIG5V.n12268 ASIG5V.n1266 2.24164
R46594 ASIG5V.n12030 ASIG5V.n1272 2.24164
R46595 ASIG5V.n12268 ASIG5V.n1265 2.24164
R46596 ASIG5V.n12038 ASIG5V.n1272 2.24164
R46597 ASIG5V.n12268 ASIG5V.n1264 2.24164
R46598 ASIG5V.n12042 ASIG5V.n1272 2.24164
R46599 ASIG5V.n12268 ASIG5V.n1263 2.24164
R46600 ASIG5V.n12050 ASIG5V.n1272 2.24164
R46601 ASIG5V.n12268 ASIG5V.n1262 2.24164
R46602 ASIG5V.n12054 ASIG5V.n1272 2.24164
R46603 ASIG5V.n12268 ASIG5V.n1261 2.24164
R46604 ASIG5V.n12062 ASIG5V.n1272 2.24164
R46605 ASIG5V.n12268 ASIG5V.n1260 2.24164
R46606 ASIG5V.n12066 ASIG5V.n1272 2.24164
R46607 ASIG5V.n12268 ASIG5V.n1259 2.24164
R46608 ASIG5V.n12074 ASIG5V.n1272 2.24164
R46609 ASIG5V.n12268 ASIG5V.n1258 2.24164
R46610 ASIG5V.n12078 ASIG5V.n1272 2.24164
R46611 ASIG5V.n12268 ASIG5V.n1257 2.24164
R46612 ASIG5V.n12086 ASIG5V.n1272 2.24164
R46613 ASIG5V.n12268 ASIG5V.n1256 2.24164
R46614 ASIG5V.n12090 ASIG5V.n1272 2.24164
R46615 ASIG5V.n12268 ASIG5V.n1255 2.24164
R46616 ASIG5V.n12098 ASIG5V.n1272 2.24164
R46617 ASIG5V.n12268 ASIG5V.n1254 2.24164
R46618 ASIG5V.n12102 ASIG5V.n1272 2.24164
R46619 ASIG5V.n12268 ASIG5V.n1253 2.24164
R46620 ASIG5V.n12110 ASIG5V.n1272 2.24164
R46621 ASIG5V.n12268 ASIG5V.n1252 2.24164
R46622 ASIG5V.n12114 ASIG5V.n1272 2.24164
R46623 ASIG5V.n12268 ASIG5V.n1251 2.24164
R46624 ASIG5V.n12122 ASIG5V.n1272 2.24164
R46625 ASIG5V.n12268 ASIG5V.n1250 2.24164
R46626 ASIG5V.n12126 ASIG5V.n1272 2.24164
R46627 ASIG5V.n12268 ASIG5V.n1249 2.24164
R46628 ASIG5V.n12134 ASIG5V.n1272 2.24164
R46629 ASIG5V.n12268 ASIG5V.n1248 2.24164
R46630 ASIG5V.n12138 ASIG5V.n1272 2.24164
R46631 ASIG5V.n12268 ASIG5V.n1247 2.24164
R46632 ASIG5V.n12146 ASIG5V.n1272 2.24164
R46633 ASIG5V.n12268 ASIG5V.n1246 2.24164
R46634 ASIG5V.n12150 ASIG5V.n1272 2.24164
R46635 ASIG5V.n12268 ASIG5V.n1245 2.24164
R46636 ASIG5V.n12158 ASIG5V.n1272 2.24164
R46637 ASIG5V.n12268 ASIG5V.n1244 2.24164
R46638 ASIG5V.n12162 ASIG5V.n1272 2.24164
R46639 ASIG5V.n12268 ASIG5V.n1243 2.24164
R46640 ASIG5V.n12170 ASIG5V.n1272 2.24164
R46641 ASIG5V.n12268 ASIG5V.n1242 2.24164
R46642 ASIG5V.n12174 ASIG5V.n1272 2.24164
R46643 ASIG5V.n12268 ASIG5V.n1241 2.24164
R46644 ASIG5V.n12182 ASIG5V.n1272 2.24164
R46645 ASIG5V.n12268 ASIG5V.n1240 2.24164
R46646 ASIG5V.n12186 ASIG5V.n1272 2.24164
R46647 ASIG5V.n12268 ASIG5V.n1239 2.24164
R46648 ASIG5V.n12194 ASIG5V.n1272 2.24164
R46649 ASIG5V.n12268 ASIG5V.n1238 2.24164
R46650 ASIG5V.n12198 ASIG5V.n1272 2.24164
R46651 ASIG5V.n12268 ASIG5V.n1237 2.24164
R46652 ASIG5V.n12206 ASIG5V.n1272 2.24164
R46653 ASIG5V.n12268 ASIG5V.n1236 2.24164
R46654 ASIG5V.n12210 ASIG5V.n1272 2.24164
R46655 ASIG5V.n12268 ASIG5V.n1235 2.24164
R46656 ASIG5V.n12218 ASIG5V.n1272 2.24164
R46657 ASIG5V.n12268 ASIG5V.n1234 2.24164
R46658 ASIG5V.n12222 ASIG5V.n1272 2.24164
R46659 ASIG5V.n12268 ASIG5V.n1233 2.24164
R46660 ASIG5V.n12230 ASIG5V.n1272 2.24164
R46661 ASIG5V.n12268 ASIG5V.n1232 2.24164
R46662 ASIG5V.n12234 ASIG5V.n1272 2.24164
R46663 ASIG5V.n12268 ASIG5V.n1231 2.24164
R46664 ASIG5V.n12242 ASIG5V.n1272 2.24164
R46665 ASIG5V.n12268 ASIG5V.n1230 2.24164
R46666 ASIG5V.n12246 ASIG5V.n1272 2.24164
R46667 ASIG5V.n12268 ASIG5V.n1229 2.24164
R46668 ASIG5V.n12254 ASIG5V.n1272 2.24164
R46669 ASIG5V.n12268 ASIG5V.n1228 2.24164
R46670 ASIG5V.n12258 ASIG5V.n1272 2.24164
R46671 ASIG5V.n12268 ASIG5V.n1227 2.24164
R46672 ASIG5V.n12266 ASIG5V.n1272 2.24164
R46673 ASIG5V.n968 ASIG5V.n866 2.24164
R46674 ASIG5V.n970 ASIG5V.n877 2.24164
R46675 ASIG5V.n972 ASIG5V.n866 2.24164
R46676 ASIG5V.n962 ASIG5V.n877 2.24164
R46677 ASIG5V.n980 ASIG5V.n866 2.24164
R46678 ASIG5V.n982 ASIG5V.n877 2.24164
R46679 ASIG5V.n984 ASIG5V.n866 2.24164
R46680 ASIG5V.n958 ASIG5V.n877 2.24164
R46681 ASIG5V.n992 ASIG5V.n866 2.24164
R46682 ASIG5V.n994 ASIG5V.n877 2.24164
R46683 ASIG5V.n996 ASIG5V.n866 2.24164
R46684 ASIG5V.n954 ASIG5V.n877 2.24164
R46685 ASIG5V.n1004 ASIG5V.n866 2.24164
R46686 ASIG5V.n1006 ASIG5V.n877 2.24164
R46687 ASIG5V.n1008 ASIG5V.n866 2.24164
R46688 ASIG5V.n950 ASIG5V.n877 2.24164
R46689 ASIG5V.n1016 ASIG5V.n866 2.24164
R46690 ASIG5V.n1018 ASIG5V.n877 2.24164
R46691 ASIG5V.n1020 ASIG5V.n866 2.24164
R46692 ASIG5V.n946 ASIG5V.n877 2.24164
R46693 ASIG5V.n1028 ASIG5V.n866 2.24164
R46694 ASIG5V.n1030 ASIG5V.n877 2.24164
R46695 ASIG5V.n1032 ASIG5V.n866 2.24164
R46696 ASIG5V.n942 ASIG5V.n877 2.24164
R46697 ASIG5V.n1040 ASIG5V.n866 2.24164
R46698 ASIG5V.n1042 ASIG5V.n877 2.24164
R46699 ASIG5V.n1044 ASIG5V.n866 2.24164
R46700 ASIG5V.n938 ASIG5V.n877 2.24164
R46701 ASIG5V.n1052 ASIG5V.n866 2.24164
R46702 ASIG5V.n1054 ASIG5V.n877 2.24164
R46703 ASIG5V.n1056 ASIG5V.n866 2.24164
R46704 ASIG5V.n934 ASIG5V.n877 2.24164
R46705 ASIG5V.n1064 ASIG5V.n866 2.24164
R46706 ASIG5V.n1066 ASIG5V.n877 2.24164
R46707 ASIG5V.n1068 ASIG5V.n866 2.24164
R46708 ASIG5V.n930 ASIG5V.n877 2.24164
R46709 ASIG5V.n1076 ASIG5V.n866 2.24164
R46710 ASIG5V.n1078 ASIG5V.n877 2.24164
R46711 ASIG5V.n1080 ASIG5V.n866 2.24164
R46712 ASIG5V.n926 ASIG5V.n877 2.24164
R46713 ASIG5V.n1088 ASIG5V.n866 2.24164
R46714 ASIG5V.n1090 ASIG5V.n877 2.24164
R46715 ASIG5V.n1092 ASIG5V.n866 2.24164
R46716 ASIG5V.n922 ASIG5V.n877 2.24164
R46717 ASIG5V.n1100 ASIG5V.n866 2.24164
R46718 ASIG5V.n1102 ASIG5V.n877 2.24164
R46719 ASIG5V.n1104 ASIG5V.n866 2.24164
R46720 ASIG5V.n918 ASIG5V.n877 2.24164
R46721 ASIG5V.n1112 ASIG5V.n866 2.24164
R46722 ASIG5V.n1114 ASIG5V.n877 2.24164
R46723 ASIG5V.n1116 ASIG5V.n866 2.24164
R46724 ASIG5V.n914 ASIG5V.n877 2.24164
R46725 ASIG5V.n1124 ASIG5V.n866 2.24164
R46726 ASIG5V.n1126 ASIG5V.n877 2.24164
R46727 ASIG5V.n1128 ASIG5V.n866 2.24164
R46728 ASIG5V.n910 ASIG5V.n877 2.24164
R46729 ASIG5V.n1136 ASIG5V.n866 2.24164
R46730 ASIG5V.n1138 ASIG5V.n877 2.24164
R46731 ASIG5V.n1140 ASIG5V.n866 2.24164
R46732 ASIG5V.n906 ASIG5V.n877 2.24164
R46733 ASIG5V.n1148 ASIG5V.n866 2.24164
R46734 ASIG5V.n1150 ASIG5V.n877 2.24164
R46735 ASIG5V.n1152 ASIG5V.n866 2.24164
R46736 ASIG5V.n902 ASIG5V.n877 2.24164
R46737 ASIG5V.n1160 ASIG5V.n866 2.24164
R46738 ASIG5V.n1162 ASIG5V.n877 2.24164
R46739 ASIG5V.n1164 ASIG5V.n866 2.24164
R46740 ASIG5V.n898 ASIG5V.n877 2.24164
R46741 ASIG5V.n1172 ASIG5V.n866 2.24164
R46742 ASIG5V.n1174 ASIG5V.n877 2.24164
R46743 ASIG5V.n1176 ASIG5V.n866 2.24164
R46744 ASIG5V.n894 ASIG5V.n877 2.24164
R46745 ASIG5V.n1184 ASIG5V.n866 2.24164
R46746 ASIG5V.n1186 ASIG5V.n877 2.24164
R46747 ASIG5V.n1188 ASIG5V.n866 2.24164
R46748 ASIG5V.n890 ASIG5V.n877 2.24164
R46749 ASIG5V.n1196 ASIG5V.n866 2.24164
R46750 ASIG5V.n1198 ASIG5V.n877 2.24164
R46751 ASIG5V.n1200 ASIG5V.n866 2.24164
R46752 ASIG5V.n886 ASIG5V.n877 2.24164
R46753 ASIG5V.n1209 ASIG5V.n866 2.24164
R46754 ASIG5V.n1211 ASIG5V.n877 2.24164
R46755 ASIG5V.n1213 ASIG5V.n866 2.24164
R46756 ASIG5V.n615 ASIG5V.n521 2.24164
R46757 ASIG5V.n12301 ASIG5V.n569 2.24164
R46758 ASIG5V.n622 ASIG5V.n521 2.24164
R46759 ASIG5V.n12301 ASIG5V.n568 2.24164
R46760 ASIG5V.n626 ASIG5V.n521 2.24164
R46761 ASIG5V.n12301 ASIG5V.n567 2.24164
R46762 ASIG5V.n634 ASIG5V.n521 2.24164
R46763 ASIG5V.n12301 ASIG5V.n566 2.24164
R46764 ASIG5V.n638 ASIG5V.n521 2.24164
R46765 ASIG5V.n12301 ASIG5V.n565 2.24164
R46766 ASIG5V.n646 ASIG5V.n521 2.24164
R46767 ASIG5V.n12301 ASIG5V.n564 2.24164
R46768 ASIG5V.n650 ASIG5V.n521 2.24164
R46769 ASIG5V.n12301 ASIG5V.n563 2.24164
R46770 ASIG5V.n658 ASIG5V.n521 2.24164
R46771 ASIG5V.n12301 ASIG5V.n562 2.24164
R46772 ASIG5V.n662 ASIG5V.n521 2.24164
R46773 ASIG5V.n12301 ASIG5V.n561 2.24164
R46774 ASIG5V.n670 ASIG5V.n521 2.24164
R46775 ASIG5V.n12301 ASIG5V.n560 2.24164
R46776 ASIG5V.n674 ASIG5V.n521 2.24164
R46777 ASIG5V.n12301 ASIG5V.n559 2.24164
R46778 ASIG5V.n682 ASIG5V.n521 2.24164
R46779 ASIG5V.n12301 ASIG5V.n558 2.24164
R46780 ASIG5V.n686 ASIG5V.n521 2.24164
R46781 ASIG5V.n12301 ASIG5V.n557 2.24164
R46782 ASIG5V.n694 ASIG5V.n521 2.24164
R46783 ASIG5V.n12301 ASIG5V.n556 2.24164
R46784 ASIG5V.n698 ASIG5V.n521 2.24164
R46785 ASIG5V.n12301 ASIG5V.n555 2.24164
R46786 ASIG5V.n706 ASIG5V.n521 2.24164
R46787 ASIG5V.n12301 ASIG5V.n554 2.24164
R46788 ASIG5V.n710 ASIG5V.n521 2.24164
R46789 ASIG5V.n12301 ASIG5V.n553 2.24164
R46790 ASIG5V.n718 ASIG5V.n521 2.24164
R46791 ASIG5V.n12301 ASIG5V.n552 2.24164
R46792 ASIG5V.n722 ASIG5V.n521 2.24164
R46793 ASIG5V.n12301 ASIG5V.n551 2.24164
R46794 ASIG5V.n730 ASIG5V.n521 2.24164
R46795 ASIG5V.n12301 ASIG5V.n550 2.24164
R46796 ASIG5V.n734 ASIG5V.n521 2.24164
R46797 ASIG5V.n12301 ASIG5V.n549 2.24164
R46798 ASIG5V.n742 ASIG5V.n521 2.24164
R46799 ASIG5V.n12301 ASIG5V.n548 2.24164
R46800 ASIG5V.n746 ASIG5V.n521 2.24164
R46801 ASIG5V.n12301 ASIG5V.n547 2.24164
R46802 ASIG5V.n754 ASIG5V.n521 2.24164
R46803 ASIG5V.n12301 ASIG5V.n546 2.24164
R46804 ASIG5V.n758 ASIG5V.n521 2.24164
R46805 ASIG5V.n12301 ASIG5V.n545 2.24164
R46806 ASIG5V.n766 ASIG5V.n521 2.24164
R46807 ASIG5V.n12301 ASIG5V.n544 2.24164
R46808 ASIG5V.n770 ASIG5V.n521 2.24164
R46809 ASIG5V.n12301 ASIG5V.n543 2.24164
R46810 ASIG5V.n778 ASIG5V.n521 2.24164
R46811 ASIG5V.n12301 ASIG5V.n542 2.24164
R46812 ASIG5V.n782 ASIG5V.n521 2.24164
R46813 ASIG5V.n12301 ASIG5V.n541 2.24164
R46814 ASIG5V.n790 ASIG5V.n521 2.24164
R46815 ASIG5V.n12301 ASIG5V.n540 2.24164
R46816 ASIG5V.n794 ASIG5V.n521 2.24164
R46817 ASIG5V.n12301 ASIG5V.n539 2.24164
R46818 ASIG5V.n802 ASIG5V.n521 2.24164
R46819 ASIG5V.n12301 ASIG5V.n538 2.24164
R46820 ASIG5V.n806 ASIG5V.n521 2.24164
R46821 ASIG5V.n12301 ASIG5V.n537 2.24164
R46822 ASIG5V.n814 ASIG5V.n521 2.24164
R46823 ASIG5V.n12301 ASIG5V.n536 2.24164
R46824 ASIG5V.n818 ASIG5V.n521 2.24164
R46825 ASIG5V.n12301 ASIG5V.n535 2.24164
R46826 ASIG5V.n826 ASIG5V.n521 2.24164
R46827 ASIG5V.n12301 ASIG5V.n534 2.24164
R46828 ASIG5V.n830 ASIG5V.n521 2.24164
R46829 ASIG5V.n12301 ASIG5V.n533 2.24164
R46830 ASIG5V.n838 ASIG5V.n521 2.24164
R46831 ASIG5V.n12301 ASIG5V.n532 2.24164
R46832 ASIG5V.n842 ASIG5V.n521 2.24164
R46833 ASIG5V.n12301 ASIG5V.n531 2.24164
R46834 ASIG5V.n850 ASIG5V.n521 2.24164
R46835 ASIG5V.n12301 ASIG5V.n530 2.24164
R46836 ASIG5V.n854 ASIG5V.n521 2.24164
R46837 ASIG5V.n12301 ASIG5V.n529 2.24164
R46838 ASIG5V.n12299 ASIG5V.n521 2.24164
R46839 ASIG5V.n261 ASIG5V.n219 2.24164
R46840 ASIG5V.n12323 ASIG5V.n214 2.24164
R46841 ASIG5V.n268 ASIG5V.n219 2.24164
R46842 ASIG5V.n12323 ASIG5V.n213 2.24164
R46843 ASIG5V.n272 ASIG5V.n219 2.24164
R46844 ASIG5V.n12323 ASIG5V.n212 2.24164
R46845 ASIG5V.n280 ASIG5V.n219 2.24164
R46846 ASIG5V.n12323 ASIG5V.n211 2.24164
R46847 ASIG5V.n284 ASIG5V.n219 2.24164
R46848 ASIG5V.n12323 ASIG5V.n210 2.24164
R46849 ASIG5V.n292 ASIG5V.n219 2.24164
R46850 ASIG5V.n12323 ASIG5V.n209 2.24164
R46851 ASIG5V.n296 ASIG5V.n219 2.24164
R46852 ASIG5V.n12323 ASIG5V.n208 2.24164
R46853 ASIG5V.n304 ASIG5V.n219 2.24164
R46854 ASIG5V.n12323 ASIG5V.n207 2.24164
R46855 ASIG5V.n308 ASIG5V.n219 2.24164
R46856 ASIG5V.n12323 ASIG5V.n206 2.24164
R46857 ASIG5V.n316 ASIG5V.n219 2.24164
R46858 ASIG5V.n12323 ASIG5V.n205 2.24164
R46859 ASIG5V.n320 ASIG5V.n219 2.24164
R46860 ASIG5V.n12323 ASIG5V.n204 2.24164
R46861 ASIG5V.n328 ASIG5V.n219 2.24164
R46862 ASIG5V.n12323 ASIG5V.n203 2.24164
R46863 ASIG5V.n332 ASIG5V.n219 2.24164
R46864 ASIG5V.n12323 ASIG5V.n202 2.24164
R46865 ASIG5V.n340 ASIG5V.n219 2.24164
R46866 ASIG5V.n12323 ASIG5V.n201 2.24164
R46867 ASIG5V.n344 ASIG5V.n219 2.24164
R46868 ASIG5V.n12323 ASIG5V.n200 2.24164
R46869 ASIG5V.n352 ASIG5V.n219 2.24164
R46870 ASIG5V.n12323 ASIG5V.n199 2.24164
R46871 ASIG5V.n356 ASIG5V.n219 2.24164
R46872 ASIG5V.n12323 ASIG5V.n198 2.24164
R46873 ASIG5V.n364 ASIG5V.n219 2.24164
R46874 ASIG5V.n12323 ASIG5V.n197 2.24164
R46875 ASIG5V.n368 ASIG5V.n219 2.24164
R46876 ASIG5V.n12323 ASIG5V.n196 2.24164
R46877 ASIG5V.n376 ASIG5V.n219 2.24164
R46878 ASIG5V.n12323 ASIG5V.n195 2.24164
R46879 ASIG5V.n380 ASIG5V.n219 2.24164
R46880 ASIG5V.n12323 ASIG5V.n194 2.24164
R46881 ASIG5V.n388 ASIG5V.n219 2.24164
R46882 ASIG5V.n12323 ASIG5V.n193 2.24164
R46883 ASIG5V.n392 ASIG5V.n219 2.24164
R46884 ASIG5V.n12323 ASIG5V.n192 2.24164
R46885 ASIG5V.n400 ASIG5V.n219 2.24164
R46886 ASIG5V.n12323 ASIG5V.n191 2.24164
R46887 ASIG5V.n404 ASIG5V.n219 2.24164
R46888 ASIG5V.n12323 ASIG5V.n190 2.24164
R46889 ASIG5V.n412 ASIG5V.n219 2.24164
R46890 ASIG5V.n12323 ASIG5V.n189 2.24164
R46891 ASIG5V.n416 ASIG5V.n219 2.24164
R46892 ASIG5V.n12323 ASIG5V.n188 2.24164
R46893 ASIG5V.n424 ASIG5V.n219 2.24164
R46894 ASIG5V.n12323 ASIG5V.n187 2.24164
R46895 ASIG5V.n428 ASIG5V.n219 2.24164
R46896 ASIG5V.n12323 ASIG5V.n186 2.24164
R46897 ASIG5V.n436 ASIG5V.n219 2.24164
R46898 ASIG5V.n12323 ASIG5V.n185 2.24164
R46899 ASIG5V.n440 ASIG5V.n219 2.24164
R46900 ASIG5V.n12323 ASIG5V.n184 2.24164
R46901 ASIG5V.n448 ASIG5V.n219 2.24164
R46902 ASIG5V.n12323 ASIG5V.n183 2.24164
R46903 ASIG5V.n452 ASIG5V.n219 2.24164
R46904 ASIG5V.n12323 ASIG5V.n182 2.24164
R46905 ASIG5V.n460 ASIG5V.n219 2.24164
R46906 ASIG5V.n12323 ASIG5V.n181 2.24164
R46907 ASIG5V.n464 ASIG5V.n219 2.24164
R46908 ASIG5V.n12323 ASIG5V.n180 2.24164
R46909 ASIG5V.n472 ASIG5V.n219 2.24164
R46910 ASIG5V.n12323 ASIG5V.n179 2.24164
R46911 ASIG5V.n476 ASIG5V.n219 2.24164
R46912 ASIG5V.n12323 ASIG5V.n178 2.24164
R46913 ASIG5V.n484 ASIG5V.n219 2.24164
R46914 ASIG5V.n12323 ASIG5V.n177 2.24164
R46915 ASIG5V.n488 ASIG5V.n219 2.24164
R46916 ASIG5V.n12323 ASIG5V.n176 2.24164
R46917 ASIG5V.n496 ASIG5V.n219 2.24164
R46918 ASIG5V.n12323 ASIG5V.n175 2.24164
R46919 ASIG5V.n500 ASIG5V.n219 2.24164
R46920 ASIG5V.n12323 ASIG5V.n174 2.24164
R46921 ASIG5V.n12321 ASIG5V.n219 2.24164
R46922 ASIG5V.n12528 ASIG5V.n12527 2.24164
R46923 ASIG5V.n12525 ASIG5V.n97 2.24164
R46924 ASIG5V.n12528 ASIG5V.n51 2.24164
R46925 ASIG5V.n12525 ASIG5V.n96 2.24164
R46926 ASIG5V.n12528 ASIG5V.n50 2.24164
R46927 ASIG5V.n12525 ASIG5V.n95 2.24164
R46928 ASIG5V.n12528 ASIG5V.n49 2.24164
R46929 ASIG5V.n12525 ASIG5V.n94 2.24164
R46930 ASIG5V.n12528 ASIG5V.n48 2.24164
R46931 ASIG5V.n12525 ASIG5V.n93 2.24164
R46932 ASIG5V.n12528 ASIG5V.n47 2.24164
R46933 ASIG5V.n12525 ASIG5V.n92 2.24164
R46934 ASIG5V.n12528 ASIG5V.n46 2.24164
R46935 ASIG5V.n12525 ASIG5V.n91 2.24164
R46936 ASIG5V.n12528 ASIG5V.n45 2.24164
R46937 ASIG5V.n12525 ASIG5V.n90 2.24164
R46938 ASIG5V.n12528 ASIG5V.n44 2.24164
R46939 ASIG5V.n12525 ASIG5V.n89 2.24164
R46940 ASIG5V.n12528 ASIG5V.n43 2.24164
R46941 ASIG5V.n12525 ASIG5V.n88 2.24164
R46942 ASIG5V.n12528 ASIG5V.n42 2.24164
R46943 ASIG5V.n12525 ASIG5V.n87 2.24164
R46944 ASIG5V.n12528 ASIG5V.n41 2.24164
R46945 ASIG5V.n12525 ASIG5V.n86 2.24164
R46946 ASIG5V.n12528 ASIG5V.n40 2.24164
R46947 ASIG5V.n12525 ASIG5V.n85 2.24164
R46948 ASIG5V.n12528 ASIG5V.n39 2.24164
R46949 ASIG5V.n12525 ASIG5V.n84 2.24164
R46950 ASIG5V.n12528 ASIG5V.n38 2.24164
R46951 ASIG5V.n12525 ASIG5V.n83 2.24164
R46952 ASIG5V.n12528 ASIG5V.n37 2.24164
R46953 ASIG5V.n12525 ASIG5V.n82 2.24164
R46954 ASIG5V.n12528 ASIG5V.n36 2.24164
R46955 ASIG5V.n12525 ASIG5V.n81 2.24164
R46956 ASIG5V.n12528 ASIG5V.n35 2.24164
R46957 ASIG5V.n12525 ASIG5V.n80 2.24164
R46958 ASIG5V.n12528 ASIG5V.n34 2.24164
R46959 ASIG5V.n12525 ASIG5V.n79 2.24164
R46960 ASIG5V.n12528 ASIG5V.n33 2.24164
R46961 ASIG5V.n12525 ASIG5V.n78 2.24164
R46962 ASIG5V.n12528 ASIG5V.n32 2.24164
R46963 ASIG5V.n12525 ASIG5V.n77 2.24164
R46964 ASIG5V.n12528 ASIG5V.n31 2.24164
R46965 ASIG5V.n12525 ASIG5V.n76 2.24164
R46966 ASIG5V.n12528 ASIG5V.n30 2.24164
R46967 ASIG5V.n12525 ASIG5V.n75 2.24164
R46968 ASIG5V.n12528 ASIG5V.n29 2.24164
R46969 ASIG5V.n12525 ASIG5V.n74 2.24164
R46970 ASIG5V.n12528 ASIG5V.n28 2.24164
R46971 ASIG5V.n12525 ASIG5V.n73 2.24164
R46972 ASIG5V.n12528 ASIG5V.n27 2.24164
R46973 ASIG5V.n12525 ASIG5V.n72 2.24164
R46974 ASIG5V.n12528 ASIG5V.n26 2.24164
R46975 ASIG5V.n12525 ASIG5V.n71 2.24164
R46976 ASIG5V.n12528 ASIG5V.n25 2.24164
R46977 ASIG5V.n12525 ASIG5V.n70 2.24164
R46978 ASIG5V.n12528 ASIG5V.n24 2.24164
R46979 ASIG5V.n12525 ASIG5V.n69 2.24164
R46980 ASIG5V.n12528 ASIG5V.n23 2.24164
R46981 ASIG5V.n12525 ASIG5V.n68 2.24164
R46982 ASIG5V.n12528 ASIG5V.n22 2.24164
R46983 ASIG5V.n12525 ASIG5V.n67 2.24164
R46984 ASIG5V.n12528 ASIG5V.n21 2.24164
R46985 ASIG5V.n12525 ASIG5V.n66 2.24164
R46986 ASIG5V.n12528 ASIG5V.n20 2.24164
R46987 ASIG5V.n12525 ASIG5V.n65 2.24164
R46988 ASIG5V.n12528 ASIG5V.n19 2.24164
R46989 ASIG5V.n12525 ASIG5V.n64 2.24164
R46990 ASIG5V.n12528 ASIG5V.n18 2.24164
R46991 ASIG5V.n12525 ASIG5V.n63 2.24164
R46992 ASIG5V.n12528 ASIG5V.n17 2.24164
R46993 ASIG5V.n12525 ASIG5V.n62 2.24164
R46994 ASIG5V.n12528 ASIG5V.n16 2.24164
R46995 ASIG5V.n12525 ASIG5V.n61 2.24164
R46996 ASIG5V.n12528 ASIG5V.n15 2.24164
R46997 ASIG5V.n12525 ASIG5V.n60 2.24164
R46998 ASIG5V.n12528 ASIG5V.n14 2.24164
R46999 ASIG5V.n12525 ASIG5V.n59 2.24164
R47000 ASIG5V.n12528 ASIG5V.n13 2.24164
R47001 ASIG5V.n12525 ASIG5V.n58 2.24164
R47002 ASIG5V.n12528 ASIG5V.n12 2.24164
R47003 ASIG5V.n12525 ASIG5V.n57 2.24164
R47004 ASIG5V.n12528 ASIG5V.n11 2.24164
R47005 ASIG5V.n8881 ASIG5V.n8880 2.24164
R47006 ASIG5V.n8589 ASIG5V.n1 2.24164
R47007 ASIG5V.n8881 ASIG5V.n8318 2.24164
R47008 ASIG5V.n8871 ASIG5V.n1 2.24164
R47009 ASIG5V.n8881 ASIG5V.n8317 2.24164
R47010 ASIG5V.n8866 ASIG5V.n1 2.24164
R47011 ASIG5V.n8881 ASIG5V.n8316 2.24164
R47012 ASIG5V.n8859 ASIG5V.n1 2.24164
R47013 ASIG5V.n8881 ASIG5V.n8315 2.24164
R47014 ASIG5V.n8854 ASIG5V.n1 2.24164
R47015 ASIG5V.n8881 ASIG5V.n8314 2.24164
R47016 ASIG5V.n8847 ASIG5V.n1 2.24164
R47017 ASIG5V.n8881 ASIG5V.n8313 2.24164
R47018 ASIG5V.n8842 ASIG5V.n1 2.24164
R47019 ASIG5V.n8881 ASIG5V.n8312 2.24164
R47020 ASIG5V.n8835 ASIG5V.n1 2.24164
R47021 ASIG5V.n8881 ASIG5V.n8311 2.24164
R47022 ASIG5V.n8830 ASIG5V.n1 2.24164
R47023 ASIG5V.n8881 ASIG5V.n8310 2.24164
R47024 ASIG5V.n8823 ASIG5V.n1 2.24164
R47025 ASIG5V.n8881 ASIG5V.n8309 2.24164
R47026 ASIG5V.n8818 ASIG5V.n1 2.24164
R47027 ASIG5V.n8881 ASIG5V.n8308 2.24164
R47028 ASIG5V.n8811 ASIG5V.n1 2.24164
R47029 ASIG5V.n8881 ASIG5V.n8307 2.24164
R47030 ASIG5V.n8806 ASIG5V.n1 2.24164
R47031 ASIG5V.n8881 ASIG5V.n8306 2.24164
R47032 ASIG5V.n8799 ASIG5V.n1 2.24164
R47033 ASIG5V.n8881 ASIG5V.n8305 2.24164
R47034 ASIG5V.n8794 ASIG5V.n1 2.24164
R47035 ASIG5V.n8881 ASIG5V.n8304 2.24164
R47036 ASIG5V.n8787 ASIG5V.n1 2.24164
R47037 ASIG5V.n8881 ASIG5V.n8303 2.24164
R47038 ASIG5V.n8782 ASIG5V.n1 2.24164
R47039 ASIG5V.n8881 ASIG5V.n8302 2.24164
R47040 ASIG5V.n8775 ASIG5V.n1 2.24164
R47041 ASIG5V.n8881 ASIG5V.n8301 2.24164
R47042 ASIG5V.n8770 ASIG5V.n1 2.24164
R47043 ASIG5V.n8881 ASIG5V.n8300 2.24164
R47044 ASIG5V.n8763 ASIG5V.n1 2.24164
R47045 ASIG5V.n8881 ASIG5V.n8299 2.24164
R47046 ASIG5V.n8758 ASIG5V.n1 2.24164
R47047 ASIG5V.n8881 ASIG5V.n8298 2.24164
R47048 ASIG5V.n8751 ASIG5V.n1 2.24164
R47049 ASIG5V.n8881 ASIG5V.n8297 2.24164
R47050 ASIG5V.n8746 ASIG5V.n1 2.24164
R47051 ASIG5V.n8881 ASIG5V.n8296 2.24164
R47052 ASIG5V.n8739 ASIG5V.n1 2.24164
R47053 ASIG5V.n8881 ASIG5V.n8295 2.24164
R47054 ASIG5V.n8734 ASIG5V.n1 2.24164
R47055 ASIG5V.n8881 ASIG5V.n8294 2.24164
R47056 ASIG5V.n8727 ASIG5V.n1 2.24164
R47057 ASIG5V.n8881 ASIG5V.n8293 2.24164
R47058 ASIG5V.n8722 ASIG5V.n1 2.24164
R47059 ASIG5V.n8881 ASIG5V.n8292 2.24164
R47060 ASIG5V.n8715 ASIG5V.n1 2.24164
R47061 ASIG5V.n8881 ASIG5V.n8291 2.24164
R47062 ASIG5V.n8710 ASIG5V.n1 2.24164
R47063 ASIG5V.n8881 ASIG5V.n8290 2.24164
R47064 ASIG5V.n8703 ASIG5V.n1 2.24164
R47065 ASIG5V.n8881 ASIG5V.n8289 2.24164
R47066 ASIG5V.n8698 ASIG5V.n1 2.24164
R47067 ASIG5V.n8881 ASIG5V.n8288 2.24164
R47068 ASIG5V.n8691 ASIG5V.n1 2.24164
R47069 ASIG5V.n8881 ASIG5V.n8287 2.24164
R47070 ASIG5V.n8686 ASIG5V.n1 2.24164
R47071 ASIG5V.n8881 ASIG5V.n8286 2.24164
R47072 ASIG5V.n8679 ASIG5V.n1 2.24164
R47073 ASIG5V.n8881 ASIG5V.n8285 2.24164
R47074 ASIG5V.n8674 ASIG5V.n1 2.24164
R47075 ASIG5V.n8881 ASIG5V.n8284 2.24164
R47076 ASIG5V.n8667 ASIG5V.n1 2.24164
R47077 ASIG5V.n8881 ASIG5V.n8283 2.24164
R47078 ASIG5V.n8662 ASIG5V.n1 2.24164
R47079 ASIG5V.n8881 ASIG5V.n8282 2.24164
R47080 ASIG5V.n8655 ASIG5V.n1 2.24164
R47081 ASIG5V.n8881 ASIG5V.n8281 2.24164
R47082 ASIG5V.n8650 ASIG5V.n1 2.24164
R47083 ASIG5V.n8881 ASIG5V.n8280 2.24164
R47084 ASIG5V.n8643 ASIG5V.n1 2.24164
R47085 ASIG5V.n8881 ASIG5V.n8279 2.24164
R47086 ASIG5V.n8638 ASIG5V.n1 2.24164
R47087 ASIG5V.n8881 ASIG5V.n8278 2.24164
R47088 ASIG5V.n8895 ASIG5V.n8894 2.24164
R47089 ASIG5V.n8892 ASIG5V.n8258 2.24164
R47090 ASIG5V.n8895 ASIG5V.n8212 2.24164
R47091 ASIG5V.n8892 ASIG5V.n8257 2.24164
R47092 ASIG5V.n8895 ASIG5V.n8211 2.24164
R47093 ASIG5V.n8892 ASIG5V.n8256 2.24164
R47094 ASIG5V.n8895 ASIG5V.n8210 2.24164
R47095 ASIG5V.n8892 ASIG5V.n8255 2.24164
R47096 ASIG5V.n8895 ASIG5V.n8209 2.24164
R47097 ASIG5V.n8892 ASIG5V.n8254 2.24164
R47098 ASIG5V.n8895 ASIG5V.n8208 2.24164
R47099 ASIG5V.n8892 ASIG5V.n8253 2.24164
R47100 ASIG5V.n8895 ASIG5V.n8207 2.24164
R47101 ASIG5V.n8892 ASIG5V.n8252 2.24164
R47102 ASIG5V.n8895 ASIG5V.n8206 2.24164
R47103 ASIG5V.n8892 ASIG5V.n8251 2.24164
R47104 ASIG5V.n8895 ASIG5V.n8205 2.24164
R47105 ASIG5V.n8892 ASIG5V.n8250 2.24164
R47106 ASIG5V.n8895 ASIG5V.n8204 2.24164
R47107 ASIG5V.n8892 ASIG5V.n8249 2.24164
R47108 ASIG5V.n8895 ASIG5V.n8203 2.24164
R47109 ASIG5V.n8892 ASIG5V.n8248 2.24164
R47110 ASIG5V.n8895 ASIG5V.n8202 2.24164
R47111 ASIG5V.n8892 ASIG5V.n8247 2.24164
R47112 ASIG5V.n8895 ASIG5V.n8201 2.24164
R47113 ASIG5V.n8892 ASIG5V.n8246 2.24164
R47114 ASIG5V.n8895 ASIG5V.n8200 2.24164
R47115 ASIG5V.n8892 ASIG5V.n8245 2.24164
R47116 ASIG5V.n8895 ASIG5V.n8199 2.24164
R47117 ASIG5V.n8892 ASIG5V.n8244 2.24164
R47118 ASIG5V.n8895 ASIG5V.n8198 2.24164
R47119 ASIG5V.n8892 ASIG5V.n8243 2.24164
R47120 ASIG5V.n8895 ASIG5V.n8197 2.24164
R47121 ASIG5V.n8892 ASIG5V.n8242 2.24164
R47122 ASIG5V.n8895 ASIG5V.n8196 2.24164
R47123 ASIG5V.n8892 ASIG5V.n8241 2.24164
R47124 ASIG5V.n8895 ASIG5V.n8195 2.24164
R47125 ASIG5V.n8892 ASIG5V.n8240 2.24164
R47126 ASIG5V.n8895 ASIG5V.n8194 2.24164
R47127 ASIG5V.n8892 ASIG5V.n8239 2.24164
R47128 ASIG5V.n8895 ASIG5V.n8193 2.24164
R47129 ASIG5V.n8892 ASIG5V.n8238 2.24164
R47130 ASIG5V.n8895 ASIG5V.n8192 2.24164
R47131 ASIG5V.n8892 ASIG5V.n8237 2.24164
R47132 ASIG5V.n8895 ASIG5V.n8191 2.24164
R47133 ASIG5V.n8892 ASIG5V.n8236 2.24164
R47134 ASIG5V.n8895 ASIG5V.n8190 2.24164
R47135 ASIG5V.n8892 ASIG5V.n8235 2.24164
R47136 ASIG5V.n8895 ASIG5V.n8189 2.24164
R47137 ASIG5V.n8892 ASIG5V.n8234 2.24164
R47138 ASIG5V.n8895 ASIG5V.n8188 2.24164
R47139 ASIG5V.n8892 ASIG5V.n8233 2.24164
R47140 ASIG5V.n8895 ASIG5V.n8187 2.24164
R47141 ASIG5V.n8892 ASIG5V.n8232 2.24164
R47142 ASIG5V.n8895 ASIG5V.n8186 2.24164
R47143 ASIG5V.n8892 ASIG5V.n8231 2.24164
R47144 ASIG5V.n8895 ASIG5V.n8185 2.24164
R47145 ASIG5V.n8892 ASIG5V.n8230 2.24164
R47146 ASIG5V.n8895 ASIG5V.n8184 2.24164
R47147 ASIG5V.n8892 ASIG5V.n8229 2.24164
R47148 ASIG5V.n8895 ASIG5V.n8183 2.24164
R47149 ASIG5V.n8892 ASIG5V.n8228 2.24164
R47150 ASIG5V.n8895 ASIG5V.n8182 2.24164
R47151 ASIG5V.n8892 ASIG5V.n8227 2.24164
R47152 ASIG5V.n8895 ASIG5V.n8181 2.24164
R47153 ASIG5V.n8892 ASIG5V.n8226 2.24164
R47154 ASIG5V.n8895 ASIG5V.n8180 2.24164
R47155 ASIG5V.n8892 ASIG5V.n8225 2.24164
R47156 ASIG5V.n8895 ASIG5V.n8179 2.24164
R47157 ASIG5V.n8892 ASIG5V.n8224 2.24164
R47158 ASIG5V.n8895 ASIG5V.n8178 2.24164
R47159 ASIG5V.n8892 ASIG5V.n8223 2.24164
R47160 ASIG5V.n8895 ASIG5V.n8177 2.24164
R47161 ASIG5V.n8892 ASIG5V.n8222 2.24164
R47162 ASIG5V.n8895 ASIG5V.n8176 2.24164
R47163 ASIG5V.n8892 ASIG5V.n8221 2.24164
R47164 ASIG5V.n8895 ASIG5V.n8175 2.24164
R47165 ASIG5V.n8892 ASIG5V.n8220 2.24164
R47166 ASIG5V.n8895 ASIG5V.n8174 2.24164
R47167 ASIG5V.n8892 ASIG5V.n8219 2.24164
R47168 ASIG5V.n8895 ASIG5V.n8173 2.24164
R47169 ASIG5V.n8892 ASIG5V.n8218 2.24164
R47170 ASIG5V.n8895 ASIG5V.n8172 2.24164
R47171 ASIG5V.n7228 ASIG5V.n6891 2.24164
R47172 ASIG5V.n7226 ASIG5V.n6892 2.24164
R47173 ASIG5V.n6899 ASIG5V.n6891 2.24164
R47174 ASIG5V.n6904 ASIG5V.n6892 2.24164
R47175 ASIG5V.n7218 ASIG5V.n6891 2.24164
R47176 ASIG5V.n7216 ASIG5V.n6892 2.24164
R47177 ASIG5V.n6905 ASIG5V.n6891 2.24164
R47178 ASIG5V.n6910 ASIG5V.n6892 2.24164
R47179 ASIG5V.n7208 ASIG5V.n6891 2.24164
R47180 ASIG5V.n7206 ASIG5V.n6892 2.24164
R47181 ASIG5V.n6911 ASIG5V.n6891 2.24164
R47182 ASIG5V.n6916 ASIG5V.n6892 2.24164
R47183 ASIG5V.n7198 ASIG5V.n6891 2.24164
R47184 ASIG5V.n7196 ASIG5V.n6892 2.24164
R47185 ASIG5V.n6917 ASIG5V.n6891 2.24164
R47186 ASIG5V.n6922 ASIG5V.n6892 2.24164
R47187 ASIG5V.n7188 ASIG5V.n6891 2.24164
R47188 ASIG5V.n7186 ASIG5V.n6892 2.24164
R47189 ASIG5V.n6923 ASIG5V.n6891 2.24164
R47190 ASIG5V.n6928 ASIG5V.n6892 2.24164
R47191 ASIG5V.n7178 ASIG5V.n6891 2.24164
R47192 ASIG5V.n7176 ASIG5V.n6892 2.24164
R47193 ASIG5V.n6929 ASIG5V.n6891 2.24164
R47194 ASIG5V.n6934 ASIG5V.n6892 2.24164
R47195 ASIG5V.n7168 ASIG5V.n6891 2.24164
R47196 ASIG5V.n7166 ASIG5V.n6892 2.24164
R47197 ASIG5V.n6935 ASIG5V.n6891 2.24164
R47198 ASIG5V.n6940 ASIG5V.n6892 2.24164
R47199 ASIG5V.n7158 ASIG5V.n6891 2.24164
R47200 ASIG5V.n7156 ASIG5V.n6892 2.24164
R47201 ASIG5V.n6941 ASIG5V.n6891 2.24164
R47202 ASIG5V.n6946 ASIG5V.n6892 2.24164
R47203 ASIG5V.n7148 ASIG5V.n6891 2.24164
R47204 ASIG5V.n7146 ASIG5V.n6892 2.24164
R47205 ASIG5V.n6947 ASIG5V.n6891 2.24164
R47206 ASIG5V.n6952 ASIG5V.n6892 2.24164
R47207 ASIG5V.n7138 ASIG5V.n6891 2.24164
R47208 ASIG5V.n7136 ASIG5V.n6892 2.24164
R47209 ASIG5V.n6953 ASIG5V.n6891 2.24164
R47210 ASIG5V.n6958 ASIG5V.n6892 2.24164
R47211 ASIG5V.n7128 ASIG5V.n6891 2.24164
R47212 ASIG5V.n7126 ASIG5V.n6892 2.24164
R47213 ASIG5V.n6959 ASIG5V.n6891 2.24164
R47214 ASIG5V.n6964 ASIG5V.n6892 2.24164
R47215 ASIG5V.n7118 ASIG5V.n6891 2.24164
R47216 ASIG5V.n7116 ASIG5V.n6892 2.24164
R47217 ASIG5V.n6965 ASIG5V.n6891 2.24164
R47218 ASIG5V.n6970 ASIG5V.n6892 2.24164
R47219 ASIG5V.n7108 ASIG5V.n6891 2.24164
R47220 ASIG5V.n7106 ASIG5V.n6892 2.24164
R47221 ASIG5V.n6971 ASIG5V.n6891 2.24164
R47222 ASIG5V.n6976 ASIG5V.n6892 2.24164
R47223 ASIG5V.n7098 ASIG5V.n6891 2.24164
R47224 ASIG5V.n7096 ASIG5V.n6892 2.24164
R47225 ASIG5V.n6977 ASIG5V.n6891 2.24164
R47226 ASIG5V.n6982 ASIG5V.n6892 2.24164
R47227 ASIG5V.n7088 ASIG5V.n6891 2.24164
R47228 ASIG5V.n7086 ASIG5V.n6892 2.24164
R47229 ASIG5V.n6983 ASIG5V.n6891 2.24164
R47230 ASIG5V.n6988 ASIG5V.n6892 2.24164
R47231 ASIG5V.n7078 ASIG5V.n6891 2.24164
R47232 ASIG5V.n7076 ASIG5V.n6892 2.24164
R47233 ASIG5V.n6989 ASIG5V.n6891 2.24164
R47234 ASIG5V.n6994 ASIG5V.n6892 2.24164
R47235 ASIG5V.n7068 ASIG5V.n6891 2.24164
R47236 ASIG5V.n7066 ASIG5V.n6892 2.24164
R47237 ASIG5V.n6995 ASIG5V.n6891 2.24164
R47238 ASIG5V.n7000 ASIG5V.n6892 2.24164
R47239 ASIG5V.n7058 ASIG5V.n6891 2.24164
R47240 ASIG5V.n7056 ASIG5V.n6892 2.24164
R47241 ASIG5V.n7001 ASIG5V.n6891 2.24164
R47242 ASIG5V.n7006 ASIG5V.n6892 2.24164
R47243 ASIG5V.n7048 ASIG5V.n6891 2.24164
R47244 ASIG5V.n7046 ASIG5V.n6892 2.24164
R47245 ASIG5V.n7007 ASIG5V.n6891 2.24164
R47246 ASIG5V.n7012 ASIG5V.n6892 2.24164
R47247 ASIG5V.n7038 ASIG5V.n6891 2.24164
R47248 ASIG5V.n7036 ASIG5V.n6892 2.24164
R47249 ASIG5V.n7013 ASIG5V.n6891 2.24164
R47250 ASIG5V.n7018 ASIG5V.n6892 2.24164
R47251 ASIG5V.n7028 ASIG5V.n6891 2.24164
R47252 ASIG5V.n7026 ASIG5V.n6892 2.24164
R47253 ASIG5V.n7019 ASIG5V.n6891 2.24164
R47254 ASIG5V.n8919 ASIG5V.n8918 2.24164
R47255 ASIG5V.n8916 ASIG5V.n6631 2.24164
R47256 ASIG5V.n8919 ASIG5V.n6586 2.24164
R47257 ASIG5V.n8916 ASIG5V.n6630 2.24164
R47258 ASIG5V.n8919 ASIG5V.n6585 2.24164
R47259 ASIG5V.n8916 ASIG5V.n6629 2.24164
R47260 ASIG5V.n8919 ASIG5V.n6584 2.24164
R47261 ASIG5V.n8916 ASIG5V.n6628 2.24164
R47262 ASIG5V.n8919 ASIG5V.n6583 2.24164
R47263 ASIG5V.n8916 ASIG5V.n6627 2.24164
R47264 ASIG5V.n8919 ASIG5V.n6582 2.24164
R47265 ASIG5V.n8916 ASIG5V.n6626 2.24164
R47266 ASIG5V.n8919 ASIG5V.n6581 2.24164
R47267 ASIG5V.n8916 ASIG5V.n6625 2.24164
R47268 ASIG5V.n8919 ASIG5V.n6580 2.24164
R47269 ASIG5V.n8916 ASIG5V.n6624 2.24164
R47270 ASIG5V.n8919 ASIG5V.n6579 2.24164
R47271 ASIG5V.n8916 ASIG5V.n6623 2.24164
R47272 ASIG5V.n8919 ASIG5V.n6578 2.24164
R47273 ASIG5V.n8916 ASIG5V.n6622 2.24164
R47274 ASIG5V.n8919 ASIG5V.n6577 2.24164
R47275 ASIG5V.n8916 ASIG5V.n6621 2.24164
R47276 ASIG5V.n8919 ASIG5V.n6576 2.24164
R47277 ASIG5V.n8916 ASIG5V.n6620 2.24164
R47278 ASIG5V.n8919 ASIG5V.n6575 2.24164
R47279 ASIG5V.n8916 ASIG5V.n6619 2.24164
R47280 ASIG5V.n8919 ASIG5V.n6574 2.24164
R47281 ASIG5V.n8916 ASIG5V.n6618 2.24164
R47282 ASIG5V.n8919 ASIG5V.n6573 2.24164
R47283 ASIG5V.n8916 ASIG5V.n6617 2.24164
R47284 ASIG5V.n8919 ASIG5V.n6572 2.24164
R47285 ASIG5V.n8916 ASIG5V.n6616 2.24164
R47286 ASIG5V.n8919 ASIG5V.n6571 2.24164
R47287 ASIG5V.n8916 ASIG5V.n6615 2.24164
R47288 ASIG5V.n8919 ASIG5V.n6570 2.24164
R47289 ASIG5V.n8916 ASIG5V.n6614 2.24164
R47290 ASIG5V.n8919 ASIG5V.n6569 2.24164
R47291 ASIG5V.n8916 ASIG5V.n6613 2.24164
R47292 ASIG5V.n8919 ASIG5V.n6568 2.24164
R47293 ASIG5V.n8916 ASIG5V.n6612 2.24164
R47294 ASIG5V.n8919 ASIG5V.n6567 2.24164
R47295 ASIG5V.n8916 ASIG5V.n6611 2.24164
R47296 ASIG5V.n8919 ASIG5V.n6566 2.24164
R47297 ASIG5V.n8916 ASIG5V.n6610 2.24164
R47298 ASIG5V.n8919 ASIG5V.n6565 2.24164
R47299 ASIG5V.n8916 ASIG5V.n6609 2.24164
R47300 ASIG5V.n8919 ASIG5V.n6564 2.24164
R47301 ASIG5V.n8916 ASIG5V.n6608 2.24164
R47302 ASIG5V.n8919 ASIG5V.n6563 2.24164
R47303 ASIG5V.n8916 ASIG5V.n6607 2.24164
R47304 ASIG5V.n8919 ASIG5V.n6562 2.24164
R47305 ASIG5V.n8916 ASIG5V.n6606 2.24164
R47306 ASIG5V.n8919 ASIG5V.n6561 2.24164
R47307 ASIG5V.n8916 ASIG5V.n6605 2.24164
R47308 ASIG5V.n8919 ASIG5V.n6560 2.24164
R47309 ASIG5V.n8916 ASIG5V.n6604 2.24164
R47310 ASIG5V.n8919 ASIG5V.n6559 2.24164
R47311 ASIG5V.n8916 ASIG5V.n6603 2.24164
R47312 ASIG5V.n8919 ASIG5V.n6558 2.24164
R47313 ASIG5V.n8916 ASIG5V.n6602 2.24164
R47314 ASIG5V.n8919 ASIG5V.n6557 2.24164
R47315 ASIG5V.n8916 ASIG5V.n6601 2.24164
R47316 ASIG5V.n8919 ASIG5V.n6556 2.24164
R47317 ASIG5V.n8916 ASIG5V.n6600 2.24164
R47318 ASIG5V.n8919 ASIG5V.n6555 2.24164
R47319 ASIG5V.n8916 ASIG5V.n6599 2.24164
R47320 ASIG5V.n8919 ASIG5V.n6554 2.24164
R47321 ASIG5V.n8916 ASIG5V.n6598 2.24164
R47322 ASIG5V.n8919 ASIG5V.n6553 2.24164
R47323 ASIG5V.n8916 ASIG5V.n6597 2.24164
R47324 ASIG5V.n8919 ASIG5V.n6552 2.24164
R47325 ASIG5V.n8916 ASIG5V.n6596 2.24164
R47326 ASIG5V.n8919 ASIG5V.n6551 2.24164
R47327 ASIG5V.n8916 ASIG5V.n6595 2.24164
R47328 ASIG5V.n8919 ASIG5V.n6550 2.24164
R47329 ASIG5V.n8916 ASIG5V.n6594 2.24164
R47330 ASIG5V.n8919 ASIG5V.n6549 2.24164
R47331 ASIG5V.n8916 ASIG5V.n6593 2.24164
R47332 ASIG5V.n8919 ASIG5V.n6548 2.24164
R47333 ASIG5V.n8916 ASIG5V.n6592 2.24164
R47334 ASIG5V.n8919 ASIG5V.n6547 2.24164
R47335 ASIG5V.n8916 ASIG5V.n6591 2.24164
R47336 ASIG5V.n8919 ASIG5V.n6546 2.24164
R47337 ASIG5V.n6530 ASIG5V.n6432 2.24164
R47338 ASIG5V.n9176 ASIG5V.n6486 2.24164
R47339 ASIG5V.n8934 ASIG5V.n6432 2.24164
R47340 ASIG5V.n9176 ASIG5V.n6485 2.24164
R47341 ASIG5V.n8938 ASIG5V.n6432 2.24164
R47342 ASIG5V.n9176 ASIG5V.n6484 2.24164
R47343 ASIG5V.n8946 ASIG5V.n6432 2.24164
R47344 ASIG5V.n9176 ASIG5V.n6483 2.24164
R47345 ASIG5V.n8950 ASIG5V.n6432 2.24164
R47346 ASIG5V.n9176 ASIG5V.n6482 2.24164
R47347 ASIG5V.n8958 ASIG5V.n6432 2.24164
R47348 ASIG5V.n9176 ASIG5V.n6481 2.24164
R47349 ASIG5V.n8962 ASIG5V.n6432 2.24164
R47350 ASIG5V.n9176 ASIG5V.n6480 2.24164
R47351 ASIG5V.n8970 ASIG5V.n6432 2.24164
R47352 ASIG5V.n9176 ASIG5V.n6479 2.24164
R47353 ASIG5V.n8974 ASIG5V.n6432 2.24164
R47354 ASIG5V.n9176 ASIG5V.n6478 2.24164
R47355 ASIG5V.n8982 ASIG5V.n6432 2.24164
R47356 ASIG5V.n9176 ASIG5V.n6477 2.24164
R47357 ASIG5V.n8986 ASIG5V.n6432 2.24164
R47358 ASIG5V.n9176 ASIG5V.n6476 2.24164
R47359 ASIG5V.n8994 ASIG5V.n6432 2.24164
R47360 ASIG5V.n9176 ASIG5V.n6475 2.24164
R47361 ASIG5V.n8998 ASIG5V.n6432 2.24164
R47362 ASIG5V.n9176 ASIG5V.n6474 2.24164
R47363 ASIG5V.n9006 ASIG5V.n6432 2.24164
R47364 ASIG5V.n9176 ASIG5V.n6473 2.24164
R47365 ASIG5V.n9010 ASIG5V.n6432 2.24164
R47366 ASIG5V.n9176 ASIG5V.n6472 2.24164
R47367 ASIG5V.n9018 ASIG5V.n6432 2.24164
R47368 ASIG5V.n9176 ASIG5V.n6471 2.24164
R47369 ASIG5V.n9022 ASIG5V.n6432 2.24164
R47370 ASIG5V.n9176 ASIG5V.n6470 2.24164
R47371 ASIG5V.n9030 ASIG5V.n6432 2.24164
R47372 ASIG5V.n9176 ASIG5V.n6469 2.24164
R47373 ASIG5V.n9034 ASIG5V.n6432 2.24164
R47374 ASIG5V.n9176 ASIG5V.n6468 2.24164
R47375 ASIG5V.n9042 ASIG5V.n6432 2.24164
R47376 ASIG5V.n9176 ASIG5V.n6467 2.24164
R47377 ASIG5V.n9046 ASIG5V.n6432 2.24164
R47378 ASIG5V.n9176 ASIG5V.n6466 2.24164
R47379 ASIG5V.n9054 ASIG5V.n6432 2.24164
R47380 ASIG5V.n9176 ASIG5V.n6465 2.24164
R47381 ASIG5V.n9058 ASIG5V.n6432 2.24164
R47382 ASIG5V.n9176 ASIG5V.n6464 2.24164
R47383 ASIG5V.n9066 ASIG5V.n6432 2.24164
R47384 ASIG5V.n9176 ASIG5V.n6463 2.24164
R47385 ASIG5V.n9070 ASIG5V.n6432 2.24164
R47386 ASIG5V.n9176 ASIG5V.n6462 2.24164
R47387 ASIG5V.n9078 ASIG5V.n6432 2.24164
R47388 ASIG5V.n9176 ASIG5V.n6461 2.24164
R47389 ASIG5V.n9082 ASIG5V.n6432 2.24164
R47390 ASIG5V.n9176 ASIG5V.n6460 2.24164
R47391 ASIG5V.n9090 ASIG5V.n6432 2.24164
R47392 ASIG5V.n9176 ASIG5V.n6459 2.24164
R47393 ASIG5V.n9094 ASIG5V.n6432 2.24164
R47394 ASIG5V.n9176 ASIG5V.n6458 2.24164
R47395 ASIG5V.n9102 ASIG5V.n6432 2.24164
R47396 ASIG5V.n9176 ASIG5V.n6457 2.24164
R47397 ASIG5V.n9106 ASIG5V.n6432 2.24164
R47398 ASIG5V.n9176 ASIG5V.n6456 2.24164
R47399 ASIG5V.n9114 ASIG5V.n6432 2.24164
R47400 ASIG5V.n9176 ASIG5V.n6455 2.24164
R47401 ASIG5V.n9118 ASIG5V.n6432 2.24164
R47402 ASIG5V.n9176 ASIG5V.n6454 2.24164
R47403 ASIG5V.n9126 ASIG5V.n6432 2.24164
R47404 ASIG5V.n9176 ASIG5V.n6453 2.24164
R47405 ASIG5V.n9130 ASIG5V.n6432 2.24164
R47406 ASIG5V.n9176 ASIG5V.n6452 2.24164
R47407 ASIG5V.n9138 ASIG5V.n6432 2.24164
R47408 ASIG5V.n9176 ASIG5V.n6451 2.24164
R47409 ASIG5V.n9142 ASIG5V.n6432 2.24164
R47410 ASIG5V.n9176 ASIG5V.n6450 2.24164
R47411 ASIG5V.n9150 ASIG5V.n6432 2.24164
R47412 ASIG5V.n9176 ASIG5V.n6449 2.24164
R47413 ASIG5V.n9154 ASIG5V.n6432 2.24164
R47414 ASIG5V.n9176 ASIG5V.n6448 2.24164
R47415 ASIG5V.n9162 ASIG5V.n6432 2.24164
R47416 ASIG5V.n9176 ASIG5V.n6447 2.24164
R47417 ASIG5V.n9166 ASIG5V.n6432 2.24164
R47418 ASIG5V.n9176 ASIG5V.n6446 2.24164
R47419 ASIG5V.n9174 ASIG5V.n6432 2.24164
R47420 ASIG5V.n9382 ASIG5V.n9381 2.24164
R47421 ASIG5V.n9379 ASIG5V.n6351 2.24164
R47422 ASIG5V.n9382 ASIG5V.n6305 2.24164
R47423 ASIG5V.n9379 ASIG5V.n6350 2.24164
R47424 ASIG5V.n9382 ASIG5V.n6304 2.24164
R47425 ASIG5V.n9379 ASIG5V.n6349 2.24164
R47426 ASIG5V.n9382 ASIG5V.n6303 2.24164
R47427 ASIG5V.n9379 ASIG5V.n6348 2.24164
R47428 ASIG5V.n9382 ASIG5V.n6302 2.24164
R47429 ASIG5V.n9379 ASIG5V.n6347 2.24164
R47430 ASIG5V.n9382 ASIG5V.n6301 2.24164
R47431 ASIG5V.n9379 ASIG5V.n6346 2.24164
R47432 ASIG5V.n9382 ASIG5V.n6300 2.24164
R47433 ASIG5V.n9379 ASIG5V.n6345 2.24164
R47434 ASIG5V.n9382 ASIG5V.n6299 2.24164
R47435 ASIG5V.n9379 ASIG5V.n6344 2.24164
R47436 ASIG5V.n9382 ASIG5V.n6298 2.24164
R47437 ASIG5V.n9379 ASIG5V.n6343 2.24164
R47438 ASIG5V.n9382 ASIG5V.n6297 2.24164
R47439 ASIG5V.n9379 ASIG5V.n6342 2.24164
R47440 ASIG5V.n9382 ASIG5V.n6296 2.24164
R47441 ASIG5V.n9379 ASIG5V.n6341 2.24164
R47442 ASIG5V.n9382 ASIG5V.n6295 2.24164
R47443 ASIG5V.n9379 ASIG5V.n6340 2.24164
R47444 ASIG5V.n9382 ASIG5V.n6294 2.24164
R47445 ASIG5V.n9379 ASIG5V.n6339 2.24164
R47446 ASIG5V.n9382 ASIG5V.n6293 2.24164
R47447 ASIG5V.n9379 ASIG5V.n6338 2.24164
R47448 ASIG5V.n9382 ASIG5V.n6292 2.24164
R47449 ASIG5V.n9379 ASIG5V.n6337 2.24164
R47450 ASIG5V.n9382 ASIG5V.n6291 2.24164
R47451 ASIG5V.n9379 ASIG5V.n6336 2.24164
R47452 ASIG5V.n9382 ASIG5V.n6290 2.24164
R47453 ASIG5V.n9379 ASIG5V.n6335 2.24164
R47454 ASIG5V.n9382 ASIG5V.n6289 2.24164
R47455 ASIG5V.n9379 ASIG5V.n6334 2.24164
R47456 ASIG5V.n9382 ASIG5V.n6288 2.24164
R47457 ASIG5V.n9379 ASIG5V.n6333 2.24164
R47458 ASIG5V.n9382 ASIG5V.n6287 2.24164
R47459 ASIG5V.n9379 ASIG5V.n6332 2.24164
R47460 ASIG5V.n9382 ASIG5V.n6286 2.24164
R47461 ASIG5V.n9379 ASIG5V.n6331 2.24164
R47462 ASIG5V.n9382 ASIG5V.n6285 2.24164
R47463 ASIG5V.n9379 ASIG5V.n6330 2.24164
R47464 ASIG5V.n9382 ASIG5V.n6284 2.24164
R47465 ASIG5V.n9379 ASIG5V.n6329 2.24164
R47466 ASIG5V.n9382 ASIG5V.n6283 2.24164
R47467 ASIG5V.n9379 ASIG5V.n6328 2.24164
R47468 ASIG5V.n9382 ASIG5V.n6282 2.24164
R47469 ASIG5V.n9379 ASIG5V.n6327 2.24164
R47470 ASIG5V.n9382 ASIG5V.n6281 2.24164
R47471 ASIG5V.n9379 ASIG5V.n6326 2.24164
R47472 ASIG5V.n9382 ASIG5V.n6280 2.24164
R47473 ASIG5V.n9379 ASIG5V.n6325 2.24164
R47474 ASIG5V.n9382 ASIG5V.n6279 2.24164
R47475 ASIG5V.n9379 ASIG5V.n6324 2.24164
R47476 ASIG5V.n9382 ASIG5V.n6278 2.24164
R47477 ASIG5V.n9379 ASIG5V.n6323 2.24164
R47478 ASIG5V.n9382 ASIG5V.n6277 2.24164
R47479 ASIG5V.n9379 ASIG5V.n6322 2.24164
R47480 ASIG5V.n9382 ASIG5V.n6276 2.24164
R47481 ASIG5V.n9379 ASIG5V.n6321 2.24164
R47482 ASIG5V.n9382 ASIG5V.n6275 2.24164
R47483 ASIG5V.n9379 ASIG5V.n6320 2.24164
R47484 ASIG5V.n9382 ASIG5V.n6274 2.24164
R47485 ASIG5V.n9379 ASIG5V.n6319 2.24164
R47486 ASIG5V.n9382 ASIG5V.n6273 2.24164
R47487 ASIG5V.n9379 ASIG5V.n6318 2.24164
R47488 ASIG5V.n9382 ASIG5V.n6272 2.24164
R47489 ASIG5V.n9379 ASIG5V.n6317 2.24164
R47490 ASIG5V.n9382 ASIG5V.n6271 2.24164
R47491 ASIG5V.n9379 ASIG5V.n6316 2.24164
R47492 ASIG5V.n9382 ASIG5V.n6270 2.24164
R47493 ASIG5V.n9379 ASIG5V.n6315 2.24164
R47494 ASIG5V.n9382 ASIG5V.n6269 2.24164
R47495 ASIG5V.n9379 ASIG5V.n6314 2.24164
R47496 ASIG5V.n9382 ASIG5V.n6268 2.24164
R47497 ASIG5V.n9379 ASIG5V.n6313 2.24164
R47498 ASIG5V.n9382 ASIG5V.n6267 2.24164
R47499 ASIG5V.n9379 ASIG5V.n6312 2.24164
R47500 ASIG5V.n9382 ASIG5V.n6266 2.24164
R47501 ASIG5V.n9379 ASIG5V.n6311 2.24164
R47502 ASIG5V.n9382 ASIG5V.n6265 2.24164
R47503 ASIG5V.n9396 ASIG5V.n9395 2.24164
R47504 ASIG5V.n9393 ASIG5V.n5998 2.24164
R47505 ASIG5V.n9396 ASIG5V.n5953 2.24164
R47506 ASIG5V.n9393 ASIG5V.n5997 2.24164
R47507 ASIG5V.n9396 ASIG5V.n5952 2.24164
R47508 ASIG5V.n9393 ASIG5V.n5996 2.24164
R47509 ASIG5V.n9396 ASIG5V.n5951 2.24164
R47510 ASIG5V.n9393 ASIG5V.n5995 2.24164
R47511 ASIG5V.n9396 ASIG5V.n5950 2.24164
R47512 ASIG5V.n9393 ASIG5V.n5994 2.24164
R47513 ASIG5V.n9396 ASIG5V.n5949 2.24164
R47514 ASIG5V.n9393 ASIG5V.n5993 2.24164
R47515 ASIG5V.n9396 ASIG5V.n5948 2.24164
R47516 ASIG5V.n9393 ASIG5V.n5992 2.24164
R47517 ASIG5V.n9396 ASIG5V.n5947 2.24164
R47518 ASIG5V.n9393 ASIG5V.n5991 2.24164
R47519 ASIG5V.n9396 ASIG5V.n5946 2.24164
R47520 ASIG5V.n9393 ASIG5V.n5990 2.24164
R47521 ASIG5V.n9396 ASIG5V.n5945 2.24164
R47522 ASIG5V.n9393 ASIG5V.n5989 2.24164
R47523 ASIG5V.n9396 ASIG5V.n5944 2.24164
R47524 ASIG5V.n9393 ASIG5V.n5988 2.24164
R47525 ASIG5V.n9396 ASIG5V.n5943 2.24164
R47526 ASIG5V.n9393 ASIG5V.n5987 2.24164
R47527 ASIG5V.n9396 ASIG5V.n5942 2.24164
R47528 ASIG5V.n9393 ASIG5V.n5986 2.24164
R47529 ASIG5V.n9396 ASIG5V.n5941 2.24164
R47530 ASIG5V.n9393 ASIG5V.n5985 2.24164
R47531 ASIG5V.n9396 ASIG5V.n5940 2.24164
R47532 ASIG5V.n9393 ASIG5V.n5984 2.24164
R47533 ASIG5V.n9396 ASIG5V.n5939 2.24164
R47534 ASIG5V.n9393 ASIG5V.n5983 2.24164
R47535 ASIG5V.n9396 ASIG5V.n5938 2.24164
R47536 ASIG5V.n9393 ASIG5V.n5982 2.24164
R47537 ASIG5V.n9396 ASIG5V.n5937 2.24164
R47538 ASIG5V.n9393 ASIG5V.n5981 2.24164
R47539 ASIG5V.n9396 ASIG5V.n5936 2.24164
R47540 ASIG5V.n9393 ASIG5V.n5980 2.24164
R47541 ASIG5V.n9396 ASIG5V.n5935 2.24164
R47542 ASIG5V.n9393 ASIG5V.n5979 2.24164
R47543 ASIG5V.n9396 ASIG5V.n5934 2.24164
R47544 ASIG5V.n9393 ASIG5V.n5978 2.24164
R47545 ASIG5V.n9396 ASIG5V.n5933 2.24164
R47546 ASIG5V.n9393 ASIG5V.n5977 2.24164
R47547 ASIG5V.n9396 ASIG5V.n5932 2.24164
R47548 ASIG5V.n9393 ASIG5V.n5976 2.24164
R47549 ASIG5V.n9396 ASIG5V.n5931 2.24164
R47550 ASIG5V.n9393 ASIG5V.n5975 2.24164
R47551 ASIG5V.n9396 ASIG5V.n5930 2.24164
R47552 ASIG5V.n9393 ASIG5V.n5974 2.24164
R47553 ASIG5V.n9396 ASIG5V.n5929 2.24164
R47554 ASIG5V.n9393 ASIG5V.n5973 2.24164
R47555 ASIG5V.n9396 ASIG5V.n5928 2.24164
R47556 ASIG5V.n9393 ASIG5V.n5972 2.24164
R47557 ASIG5V.n9396 ASIG5V.n5927 2.24164
R47558 ASIG5V.n9393 ASIG5V.n5971 2.24164
R47559 ASIG5V.n9396 ASIG5V.n5926 2.24164
R47560 ASIG5V.n9393 ASIG5V.n5970 2.24164
R47561 ASIG5V.n9396 ASIG5V.n5925 2.24164
R47562 ASIG5V.n9393 ASIG5V.n5969 2.24164
R47563 ASIG5V.n9396 ASIG5V.n5924 2.24164
R47564 ASIG5V.n9393 ASIG5V.n5968 2.24164
R47565 ASIG5V.n9396 ASIG5V.n5923 2.24164
R47566 ASIG5V.n9393 ASIG5V.n5967 2.24164
R47567 ASIG5V.n9396 ASIG5V.n5922 2.24164
R47568 ASIG5V.n9393 ASIG5V.n5966 2.24164
R47569 ASIG5V.n9396 ASIG5V.n5921 2.24164
R47570 ASIG5V.n9393 ASIG5V.n5965 2.24164
R47571 ASIG5V.n9396 ASIG5V.n5920 2.24164
R47572 ASIG5V.n9393 ASIG5V.n5964 2.24164
R47573 ASIG5V.n9396 ASIG5V.n5919 2.24164
R47574 ASIG5V.n9393 ASIG5V.n5963 2.24164
R47575 ASIG5V.n9396 ASIG5V.n5918 2.24164
R47576 ASIG5V.n9393 ASIG5V.n5962 2.24164
R47577 ASIG5V.n9396 ASIG5V.n5917 2.24164
R47578 ASIG5V.n9393 ASIG5V.n5961 2.24164
R47579 ASIG5V.n9396 ASIG5V.n5916 2.24164
R47580 ASIG5V.n9393 ASIG5V.n5960 2.24164
R47581 ASIG5V.n9396 ASIG5V.n5915 2.24164
R47582 ASIG5V.n9393 ASIG5V.n5959 2.24164
R47583 ASIG5V.n9396 ASIG5V.n5914 2.24164
R47584 ASIG5V.n9393 ASIG5V.n5958 2.24164
R47585 ASIG5V.n9396 ASIG5V.n5913 2.24164
R47586 ASIG5V.n5904 ASIG5V.n5567 2.24164
R47587 ASIG5V.n5902 ASIG5V.n5568 2.24164
R47588 ASIG5V.n5575 ASIG5V.n5567 2.24164
R47589 ASIG5V.n5580 ASIG5V.n5568 2.24164
R47590 ASIG5V.n5894 ASIG5V.n5567 2.24164
R47591 ASIG5V.n5892 ASIG5V.n5568 2.24164
R47592 ASIG5V.n5581 ASIG5V.n5567 2.24164
R47593 ASIG5V.n5586 ASIG5V.n5568 2.24164
R47594 ASIG5V.n5884 ASIG5V.n5567 2.24164
R47595 ASIG5V.n5882 ASIG5V.n5568 2.24164
R47596 ASIG5V.n5587 ASIG5V.n5567 2.24164
R47597 ASIG5V.n5592 ASIG5V.n5568 2.24164
R47598 ASIG5V.n5874 ASIG5V.n5567 2.24164
R47599 ASIG5V.n5872 ASIG5V.n5568 2.24164
R47600 ASIG5V.n5593 ASIG5V.n5567 2.24164
R47601 ASIG5V.n5598 ASIG5V.n5568 2.24164
R47602 ASIG5V.n5864 ASIG5V.n5567 2.24164
R47603 ASIG5V.n5862 ASIG5V.n5568 2.24164
R47604 ASIG5V.n5599 ASIG5V.n5567 2.24164
R47605 ASIG5V.n5604 ASIG5V.n5568 2.24164
R47606 ASIG5V.n5854 ASIG5V.n5567 2.24164
R47607 ASIG5V.n5852 ASIG5V.n5568 2.24164
R47608 ASIG5V.n5605 ASIG5V.n5567 2.24164
R47609 ASIG5V.n5610 ASIG5V.n5568 2.24164
R47610 ASIG5V.n5844 ASIG5V.n5567 2.24164
R47611 ASIG5V.n5842 ASIG5V.n5568 2.24164
R47612 ASIG5V.n5611 ASIG5V.n5567 2.24164
R47613 ASIG5V.n5616 ASIG5V.n5568 2.24164
R47614 ASIG5V.n5834 ASIG5V.n5567 2.24164
R47615 ASIG5V.n5832 ASIG5V.n5568 2.24164
R47616 ASIG5V.n5617 ASIG5V.n5567 2.24164
R47617 ASIG5V.n5622 ASIG5V.n5568 2.24164
R47618 ASIG5V.n5824 ASIG5V.n5567 2.24164
R47619 ASIG5V.n5822 ASIG5V.n5568 2.24164
R47620 ASIG5V.n5623 ASIG5V.n5567 2.24164
R47621 ASIG5V.n5628 ASIG5V.n5568 2.24164
R47622 ASIG5V.n5814 ASIG5V.n5567 2.24164
R47623 ASIG5V.n5812 ASIG5V.n5568 2.24164
R47624 ASIG5V.n5629 ASIG5V.n5567 2.24164
R47625 ASIG5V.n5634 ASIG5V.n5568 2.24164
R47626 ASIG5V.n5804 ASIG5V.n5567 2.24164
R47627 ASIG5V.n5802 ASIG5V.n5568 2.24164
R47628 ASIG5V.n5635 ASIG5V.n5567 2.24164
R47629 ASIG5V.n5640 ASIG5V.n5568 2.24164
R47630 ASIG5V.n5794 ASIG5V.n5567 2.24164
R47631 ASIG5V.n5792 ASIG5V.n5568 2.24164
R47632 ASIG5V.n5641 ASIG5V.n5567 2.24164
R47633 ASIG5V.n5646 ASIG5V.n5568 2.24164
R47634 ASIG5V.n5784 ASIG5V.n5567 2.24164
R47635 ASIG5V.n5782 ASIG5V.n5568 2.24164
R47636 ASIG5V.n5647 ASIG5V.n5567 2.24164
R47637 ASIG5V.n5652 ASIG5V.n5568 2.24164
R47638 ASIG5V.n5774 ASIG5V.n5567 2.24164
R47639 ASIG5V.n5772 ASIG5V.n5568 2.24164
R47640 ASIG5V.n5653 ASIG5V.n5567 2.24164
R47641 ASIG5V.n5658 ASIG5V.n5568 2.24164
R47642 ASIG5V.n5764 ASIG5V.n5567 2.24164
R47643 ASIG5V.n5762 ASIG5V.n5568 2.24164
R47644 ASIG5V.n5659 ASIG5V.n5567 2.24164
R47645 ASIG5V.n5664 ASIG5V.n5568 2.24164
R47646 ASIG5V.n5754 ASIG5V.n5567 2.24164
R47647 ASIG5V.n5752 ASIG5V.n5568 2.24164
R47648 ASIG5V.n5665 ASIG5V.n5567 2.24164
R47649 ASIG5V.n5670 ASIG5V.n5568 2.24164
R47650 ASIG5V.n5744 ASIG5V.n5567 2.24164
R47651 ASIG5V.n5742 ASIG5V.n5568 2.24164
R47652 ASIG5V.n5671 ASIG5V.n5567 2.24164
R47653 ASIG5V.n5676 ASIG5V.n5568 2.24164
R47654 ASIG5V.n5734 ASIG5V.n5567 2.24164
R47655 ASIG5V.n5732 ASIG5V.n5568 2.24164
R47656 ASIG5V.n5677 ASIG5V.n5567 2.24164
R47657 ASIG5V.n5682 ASIG5V.n5568 2.24164
R47658 ASIG5V.n5724 ASIG5V.n5567 2.24164
R47659 ASIG5V.n5722 ASIG5V.n5568 2.24164
R47660 ASIG5V.n5683 ASIG5V.n5567 2.24164
R47661 ASIG5V.n5688 ASIG5V.n5568 2.24164
R47662 ASIG5V.n5714 ASIG5V.n5567 2.24164
R47663 ASIG5V.n5712 ASIG5V.n5568 2.24164
R47664 ASIG5V.n5689 ASIG5V.n5567 2.24164
R47665 ASIG5V.n5694 ASIG5V.n5568 2.24164
R47666 ASIG5V.n5704 ASIG5V.n5567 2.24164
R47667 ASIG5V.n5702 ASIG5V.n5568 2.24164
R47668 ASIG5V.n5695 ASIG5V.n5567 2.24164
R47669 ASIG5V.n9419 ASIG5V.n9418 2.24164
R47670 ASIG5V.n9416 ASIG5V.n5552 2.24164
R47671 ASIG5V.n9419 ASIG5V.n5505 2.24164
R47672 ASIG5V.n9416 ASIG5V.n5551 2.24164
R47673 ASIG5V.n9419 ASIG5V.n5504 2.24164
R47674 ASIG5V.n9416 ASIG5V.n5550 2.24164
R47675 ASIG5V.n9419 ASIG5V.n5503 2.24164
R47676 ASIG5V.n9416 ASIG5V.n5549 2.24164
R47677 ASIG5V.n9419 ASIG5V.n5502 2.24164
R47678 ASIG5V.n9416 ASIG5V.n5548 2.24164
R47679 ASIG5V.n9419 ASIG5V.n5501 2.24164
R47680 ASIG5V.n9416 ASIG5V.n5547 2.24164
R47681 ASIG5V.n9419 ASIG5V.n5500 2.24164
R47682 ASIG5V.n9416 ASIG5V.n5546 2.24164
R47683 ASIG5V.n9419 ASIG5V.n5499 2.24164
R47684 ASIG5V.n9416 ASIG5V.n5545 2.24164
R47685 ASIG5V.n9419 ASIG5V.n5498 2.24164
R47686 ASIG5V.n9416 ASIG5V.n5544 2.24164
R47687 ASIG5V.n9419 ASIG5V.n5497 2.24164
R47688 ASIG5V.n9416 ASIG5V.n5543 2.24164
R47689 ASIG5V.n9419 ASIG5V.n5496 2.24164
R47690 ASIG5V.n9416 ASIG5V.n5542 2.24164
R47691 ASIG5V.n9419 ASIG5V.n5495 2.24164
R47692 ASIG5V.n9416 ASIG5V.n5541 2.24164
R47693 ASIG5V.n9419 ASIG5V.n5494 2.24164
R47694 ASIG5V.n9416 ASIG5V.n5540 2.24164
R47695 ASIG5V.n9419 ASIG5V.n5493 2.24164
R47696 ASIG5V.n9416 ASIG5V.n5539 2.24164
R47697 ASIG5V.n9419 ASIG5V.n5492 2.24164
R47698 ASIG5V.n9416 ASIG5V.n5538 2.24164
R47699 ASIG5V.n9419 ASIG5V.n5491 2.24164
R47700 ASIG5V.n9416 ASIG5V.n5537 2.24164
R47701 ASIG5V.n9419 ASIG5V.n5490 2.24164
R47702 ASIG5V.n9416 ASIG5V.n5536 2.24164
R47703 ASIG5V.n9419 ASIG5V.n5489 2.24164
R47704 ASIG5V.n9416 ASIG5V.n5535 2.24164
R47705 ASIG5V.n9419 ASIG5V.n5488 2.24164
R47706 ASIG5V.n9416 ASIG5V.n5534 2.24164
R47707 ASIG5V.n9419 ASIG5V.n5487 2.24164
R47708 ASIG5V.n9416 ASIG5V.n5533 2.24164
R47709 ASIG5V.n9419 ASIG5V.n5486 2.24164
R47710 ASIG5V.n9416 ASIG5V.n5532 2.24164
R47711 ASIG5V.n9419 ASIG5V.n5485 2.24164
R47712 ASIG5V.n9416 ASIG5V.n5531 2.24164
R47713 ASIG5V.n9419 ASIG5V.n5484 2.24164
R47714 ASIG5V.n9416 ASIG5V.n5530 2.24164
R47715 ASIG5V.n9419 ASIG5V.n5483 2.24164
R47716 ASIG5V.n9416 ASIG5V.n5529 2.24164
R47717 ASIG5V.n9419 ASIG5V.n5482 2.24164
R47718 ASIG5V.n9416 ASIG5V.n5528 2.24164
R47719 ASIG5V.n9419 ASIG5V.n5481 2.24164
R47720 ASIG5V.n9416 ASIG5V.n5527 2.24164
R47721 ASIG5V.n9419 ASIG5V.n5480 2.24164
R47722 ASIG5V.n9416 ASIG5V.n5526 2.24164
R47723 ASIG5V.n9419 ASIG5V.n5479 2.24164
R47724 ASIG5V.n9416 ASIG5V.n5525 2.24164
R47725 ASIG5V.n9419 ASIG5V.n5478 2.24164
R47726 ASIG5V.n9416 ASIG5V.n5524 2.24164
R47727 ASIG5V.n9419 ASIG5V.n5477 2.24164
R47728 ASIG5V.n9416 ASIG5V.n5523 2.24164
R47729 ASIG5V.n9419 ASIG5V.n5476 2.24164
R47730 ASIG5V.n9416 ASIG5V.n5522 2.24164
R47731 ASIG5V.n9419 ASIG5V.n5475 2.24164
R47732 ASIG5V.n9416 ASIG5V.n5521 2.24164
R47733 ASIG5V.n9419 ASIG5V.n5474 2.24164
R47734 ASIG5V.n9416 ASIG5V.n5520 2.24164
R47735 ASIG5V.n9419 ASIG5V.n5473 2.24164
R47736 ASIG5V.n9416 ASIG5V.n5519 2.24164
R47737 ASIG5V.n9419 ASIG5V.n5472 2.24164
R47738 ASIG5V.n9416 ASIG5V.n5518 2.24164
R47739 ASIG5V.n9419 ASIG5V.n5471 2.24164
R47740 ASIG5V.n9416 ASIG5V.n5517 2.24164
R47741 ASIG5V.n9419 ASIG5V.n5470 2.24164
R47742 ASIG5V.n9416 ASIG5V.n5516 2.24164
R47743 ASIG5V.n9419 ASIG5V.n5469 2.24164
R47744 ASIG5V.n9416 ASIG5V.n5515 2.24164
R47745 ASIG5V.n9419 ASIG5V.n5468 2.24164
R47746 ASIG5V.n9416 ASIG5V.n5514 2.24164
R47747 ASIG5V.n9419 ASIG5V.n5467 2.24164
R47748 ASIG5V.n9416 ASIG5V.n5513 2.24164
R47749 ASIG5V.n9419 ASIG5V.n5466 2.24164
R47750 ASIG5V.n9416 ASIG5V.n5512 2.24164
R47751 ASIG5V.n9419 ASIG5V.n5465 2.24164
R47752 ASIG5V.n5211 ASIG5V.n5170 2.24164
R47753 ASIG5V.n9432 ASIG5V.n5164 2.24164
R47754 ASIG5V.n5220 ASIG5V.n5170 2.24164
R47755 ASIG5V.n9432 ASIG5V.n5163 2.24164
R47756 ASIG5V.n5224 ASIG5V.n5170 2.24164
R47757 ASIG5V.n9432 ASIG5V.n5162 2.24164
R47758 ASIG5V.n5232 ASIG5V.n5170 2.24164
R47759 ASIG5V.n9432 ASIG5V.n5161 2.24164
R47760 ASIG5V.n5236 ASIG5V.n5170 2.24164
R47761 ASIG5V.n9432 ASIG5V.n5160 2.24164
R47762 ASIG5V.n5244 ASIG5V.n5170 2.24164
R47763 ASIG5V.n9432 ASIG5V.n5159 2.24164
R47764 ASIG5V.n5248 ASIG5V.n5170 2.24164
R47765 ASIG5V.n9432 ASIG5V.n5158 2.24164
R47766 ASIG5V.n5256 ASIG5V.n5170 2.24164
R47767 ASIG5V.n9432 ASIG5V.n5157 2.24164
R47768 ASIG5V.n5260 ASIG5V.n5170 2.24164
R47769 ASIG5V.n9432 ASIG5V.n5156 2.24164
R47770 ASIG5V.n5268 ASIG5V.n5170 2.24164
R47771 ASIG5V.n9432 ASIG5V.n5155 2.24164
R47772 ASIG5V.n5272 ASIG5V.n5170 2.24164
R47773 ASIG5V.n9432 ASIG5V.n5154 2.24164
R47774 ASIG5V.n5280 ASIG5V.n5170 2.24164
R47775 ASIG5V.n9432 ASIG5V.n5153 2.24164
R47776 ASIG5V.n5284 ASIG5V.n5170 2.24164
R47777 ASIG5V.n9432 ASIG5V.n5152 2.24164
R47778 ASIG5V.n5292 ASIG5V.n5170 2.24164
R47779 ASIG5V.n9432 ASIG5V.n5151 2.24164
R47780 ASIG5V.n5296 ASIG5V.n5170 2.24164
R47781 ASIG5V.n9432 ASIG5V.n5150 2.24164
R47782 ASIG5V.n5304 ASIG5V.n5170 2.24164
R47783 ASIG5V.n9432 ASIG5V.n5149 2.24164
R47784 ASIG5V.n5308 ASIG5V.n5170 2.24164
R47785 ASIG5V.n9432 ASIG5V.n5148 2.24164
R47786 ASIG5V.n5316 ASIG5V.n5170 2.24164
R47787 ASIG5V.n9432 ASIG5V.n5147 2.24164
R47788 ASIG5V.n5320 ASIG5V.n5170 2.24164
R47789 ASIG5V.n9432 ASIG5V.n5146 2.24164
R47790 ASIG5V.n5328 ASIG5V.n5170 2.24164
R47791 ASIG5V.n9432 ASIG5V.n5145 2.24164
R47792 ASIG5V.n5332 ASIG5V.n5170 2.24164
R47793 ASIG5V.n9432 ASIG5V.n5144 2.24164
R47794 ASIG5V.n5340 ASIG5V.n5170 2.24164
R47795 ASIG5V.n9432 ASIG5V.n5143 2.24164
R47796 ASIG5V.n5344 ASIG5V.n5170 2.24164
R47797 ASIG5V.n9432 ASIG5V.n5142 2.24164
R47798 ASIG5V.n5352 ASIG5V.n5170 2.24164
R47799 ASIG5V.n9432 ASIG5V.n5141 2.24164
R47800 ASIG5V.n5356 ASIG5V.n5170 2.24164
R47801 ASIG5V.n9432 ASIG5V.n5140 2.24164
R47802 ASIG5V.n5364 ASIG5V.n5170 2.24164
R47803 ASIG5V.n9432 ASIG5V.n5139 2.24164
R47804 ASIG5V.n5368 ASIG5V.n5170 2.24164
R47805 ASIG5V.n9432 ASIG5V.n5138 2.24164
R47806 ASIG5V.n5376 ASIG5V.n5170 2.24164
R47807 ASIG5V.n9432 ASIG5V.n5137 2.24164
R47808 ASIG5V.n5380 ASIG5V.n5170 2.24164
R47809 ASIG5V.n9432 ASIG5V.n5136 2.24164
R47810 ASIG5V.n5388 ASIG5V.n5170 2.24164
R47811 ASIG5V.n9432 ASIG5V.n5135 2.24164
R47812 ASIG5V.n5392 ASIG5V.n5170 2.24164
R47813 ASIG5V.n9432 ASIG5V.n5134 2.24164
R47814 ASIG5V.n5400 ASIG5V.n5170 2.24164
R47815 ASIG5V.n9432 ASIG5V.n5133 2.24164
R47816 ASIG5V.n5404 ASIG5V.n5170 2.24164
R47817 ASIG5V.n9432 ASIG5V.n5132 2.24164
R47818 ASIG5V.n5412 ASIG5V.n5170 2.24164
R47819 ASIG5V.n9432 ASIG5V.n5131 2.24164
R47820 ASIG5V.n5416 ASIG5V.n5170 2.24164
R47821 ASIG5V.n9432 ASIG5V.n5130 2.24164
R47822 ASIG5V.n5424 ASIG5V.n5170 2.24164
R47823 ASIG5V.n9432 ASIG5V.n5129 2.24164
R47824 ASIG5V.n5428 ASIG5V.n5170 2.24164
R47825 ASIG5V.n9432 ASIG5V.n5128 2.24164
R47826 ASIG5V.n5436 ASIG5V.n5170 2.24164
R47827 ASIG5V.n9432 ASIG5V.n5127 2.24164
R47828 ASIG5V.n5440 ASIG5V.n5170 2.24164
R47829 ASIG5V.n9432 ASIG5V.n5126 2.24164
R47830 ASIG5V.n5448 ASIG5V.n5170 2.24164
R47831 ASIG5V.n9432 ASIG5V.n5125 2.24164
R47832 ASIG5V.n5452 ASIG5V.n5170 2.24164
R47833 ASIG5V.n9432 ASIG5V.n5124 2.24164
R47834 ASIG5V.n9430 ASIG5V.n5170 2.24164
R47835 ASIG5V.n9483 ASIG5V.n3170 2.24164
R47836 ASIG5V.n9734 ASIG5V.n5115 2.24164
R47837 ASIG5V.n9492 ASIG5V.n3170 2.24164
R47838 ASIG5V.n9734 ASIG5V.n5114 2.24164
R47839 ASIG5V.n9496 ASIG5V.n3170 2.24164
R47840 ASIG5V.n9734 ASIG5V.n5113 2.24164
R47841 ASIG5V.n9504 ASIG5V.n3170 2.24164
R47842 ASIG5V.n9734 ASIG5V.n5112 2.24164
R47843 ASIG5V.n9508 ASIG5V.n3170 2.24164
R47844 ASIG5V.n9734 ASIG5V.n5111 2.24164
R47845 ASIG5V.n9516 ASIG5V.n3170 2.24164
R47846 ASIG5V.n9734 ASIG5V.n5110 2.24164
R47847 ASIG5V.n9520 ASIG5V.n3170 2.24164
R47848 ASIG5V.n9734 ASIG5V.n5109 2.24164
R47849 ASIG5V.n9528 ASIG5V.n3170 2.24164
R47850 ASIG5V.n9734 ASIG5V.n5108 2.24164
R47851 ASIG5V.n9532 ASIG5V.n3170 2.24164
R47852 ASIG5V.n9734 ASIG5V.n5107 2.24164
R47853 ASIG5V.n9540 ASIG5V.n3170 2.24164
R47854 ASIG5V.n9734 ASIG5V.n5106 2.24164
R47855 ASIG5V.n9544 ASIG5V.n3170 2.24164
R47856 ASIG5V.n9734 ASIG5V.n5105 2.24164
R47857 ASIG5V.n9552 ASIG5V.n3170 2.24164
R47858 ASIG5V.n9734 ASIG5V.n5104 2.24164
R47859 ASIG5V.n9556 ASIG5V.n3170 2.24164
R47860 ASIG5V.n9734 ASIG5V.n5103 2.24164
R47861 ASIG5V.n9564 ASIG5V.n3170 2.24164
R47862 ASIG5V.n9734 ASIG5V.n5102 2.24164
R47863 ASIG5V.n9568 ASIG5V.n3170 2.24164
R47864 ASIG5V.n9734 ASIG5V.n5101 2.24164
R47865 ASIG5V.n9576 ASIG5V.n3170 2.24164
R47866 ASIG5V.n9734 ASIG5V.n5100 2.24164
R47867 ASIG5V.n9580 ASIG5V.n3170 2.24164
R47868 ASIG5V.n9734 ASIG5V.n5099 2.24164
R47869 ASIG5V.n9588 ASIG5V.n3170 2.24164
R47870 ASIG5V.n9734 ASIG5V.n5098 2.24164
R47871 ASIG5V.n9592 ASIG5V.n3170 2.24164
R47872 ASIG5V.n9734 ASIG5V.n5097 2.24164
R47873 ASIG5V.n9600 ASIG5V.n3170 2.24164
R47874 ASIG5V.n9734 ASIG5V.n5096 2.24164
R47875 ASIG5V.n9604 ASIG5V.n3170 2.24164
R47876 ASIG5V.n9734 ASIG5V.n5095 2.24164
R47877 ASIG5V.n9612 ASIG5V.n3170 2.24164
R47878 ASIG5V.n9734 ASIG5V.n5094 2.24164
R47879 ASIG5V.n9616 ASIG5V.n3170 2.24164
R47880 ASIG5V.n9734 ASIG5V.n5093 2.24164
R47881 ASIG5V.n9624 ASIG5V.n3170 2.24164
R47882 ASIG5V.n9734 ASIG5V.n5092 2.24164
R47883 ASIG5V.n9628 ASIG5V.n3170 2.24164
R47884 ASIG5V.n9734 ASIG5V.n5091 2.24164
R47885 ASIG5V.n9636 ASIG5V.n3170 2.24164
R47886 ASIG5V.n9734 ASIG5V.n5090 2.24164
R47887 ASIG5V.n9640 ASIG5V.n3170 2.24164
R47888 ASIG5V.n9734 ASIG5V.n5089 2.24164
R47889 ASIG5V.n9648 ASIG5V.n3170 2.24164
R47890 ASIG5V.n9734 ASIG5V.n5088 2.24164
R47891 ASIG5V.n9652 ASIG5V.n3170 2.24164
R47892 ASIG5V.n9734 ASIG5V.n5087 2.24164
R47893 ASIG5V.n9660 ASIG5V.n3170 2.24164
R47894 ASIG5V.n9734 ASIG5V.n5086 2.24164
R47895 ASIG5V.n9664 ASIG5V.n3170 2.24164
R47896 ASIG5V.n9734 ASIG5V.n5085 2.24164
R47897 ASIG5V.n9672 ASIG5V.n3170 2.24164
R47898 ASIG5V.n9734 ASIG5V.n5084 2.24164
R47899 ASIG5V.n9676 ASIG5V.n3170 2.24164
R47900 ASIG5V.n9734 ASIG5V.n5083 2.24164
R47901 ASIG5V.n9684 ASIG5V.n3170 2.24164
R47902 ASIG5V.n9734 ASIG5V.n5082 2.24164
R47903 ASIG5V.n9688 ASIG5V.n3170 2.24164
R47904 ASIG5V.n9734 ASIG5V.n5081 2.24164
R47905 ASIG5V.n9696 ASIG5V.n3170 2.24164
R47906 ASIG5V.n9734 ASIG5V.n5080 2.24164
R47907 ASIG5V.n9700 ASIG5V.n3170 2.24164
R47908 ASIG5V.n9734 ASIG5V.n5079 2.24164
R47909 ASIG5V.n9708 ASIG5V.n3170 2.24164
R47910 ASIG5V.n9734 ASIG5V.n5078 2.24164
R47911 ASIG5V.n9712 ASIG5V.n3170 2.24164
R47912 ASIG5V.n9734 ASIG5V.n5077 2.24164
R47913 ASIG5V.n9720 ASIG5V.n3170 2.24164
R47914 ASIG5V.n9734 ASIG5V.n5076 2.24164
R47915 ASIG5V.n9724 ASIG5V.n3170 2.24164
R47916 ASIG5V.n9734 ASIG5V.n5075 2.24164
R47917 ASIG5V.n9732 ASIG5V.n3170 2.24164
R47918 ASIG5V.n3264 ASIG5V.n3223 2.24164
R47919 ASIG5V.n5064 ASIG5V.n3219 2.24164
R47920 ASIG5V.n4821 ASIG5V.n3223 2.24164
R47921 ASIG5V.n5064 ASIG5V.n3218 2.24164
R47922 ASIG5V.n4825 ASIG5V.n3223 2.24164
R47923 ASIG5V.n5064 ASIG5V.n3217 2.24164
R47924 ASIG5V.n4833 ASIG5V.n3223 2.24164
R47925 ASIG5V.n5064 ASIG5V.n3216 2.24164
R47926 ASIG5V.n4837 ASIG5V.n3223 2.24164
R47927 ASIG5V.n5064 ASIG5V.n3215 2.24164
R47928 ASIG5V.n4845 ASIG5V.n3223 2.24164
R47929 ASIG5V.n5064 ASIG5V.n3214 2.24164
R47930 ASIG5V.n4849 ASIG5V.n3223 2.24164
R47931 ASIG5V.n5064 ASIG5V.n3213 2.24164
R47932 ASIG5V.n4857 ASIG5V.n3223 2.24164
R47933 ASIG5V.n5064 ASIG5V.n3212 2.24164
R47934 ASIG5V.n4861 ASIG5V.n3223 2.24164
R47935 ASIG5V.n5064 ASIG5V.n3211 2.24164
R47936 ASIG5V.n4869 ASIG5V.n3223 2.24164
R47937 ASIG5V.n5064 ASIG5V.n3210 2.24164
R47938 ASIG5V.n4873 ASIG5V.n3223 2.24164
R47939 ASIG5V.n5064 ASIG5V.n3209 2.24164
R47940 ASIG5V.n4881 ASIG5V.n3223 2.24164
R47941 ASIG5V.n5064 ASIG5V.n3208 2.24164
R47942 ASIG5V.n4885 ASIG5V.n3223 2.24164
R47943 ASIG5V.n5064 ASIG5V.n3207 2.24164
R47944 ASIG5V.n4893 ASIG5V.n3223 2.24164
R47945 ASIG5V.n5064 ASIG5V.n3206 2.24164
R47946 ASIG5V.n4897 ASIG5V.n3223 2.24164
R47947 ASIG5V.n5064 ASIG5V.n3205 2.24164
R47948 ASIG5V.n4905 ASIG5V.n3223 2.24164
R47949 ASIG5V.n5064 ASIG5V.n3204 2.24164
R47950 ASIG5V.n4909 ASIG5V.n3223 2.24164
R47951 ASIG5V.n5064 ASIG5V.n3203 2.24164
R47952 ASIG5V.n4917 ASIG5V.n3223 2.24164
R47953 ASIG5V.n5064 ASIG5V.n3202 2.24164
R47954 ASIG5V.n4921 ASIG5V.n3223 2.24164
R47955 ASIG5V.n5064 ASIG5V.n3201 2.24164
R47956 ASIG5V.n4929 ASIG5V.n3223 2.24164
R47957 ASIG5V.n5064 ASIG5V.n3200 2.24164
R47958 ASIG5V.n4933 ASIG5V.n3223 2.24164
R47959 ASIG5V.n5064 ASIG5V.n3199 2.24164
R47960 ASIG5V.n4941 ASIG5V.n3223 2.24164
R47961 ASIG5V.n5064 ASIG5V.n3198 2.24164
R47962 ASIG5V.n4945 ASIG5V.n3223 2.24164
R47963 ASIG5V.n5064 ASIG5V.n3197 2.24164
R47964 ASIG5V.n4953 ASIG5V.n3223 2.24164
R47965 ASIG5V.n5064 ASIG5V.n3196 2.24164
R47966 ASIG5V.n4957 ASIG5V.n3223 2.24164
R47967 ASIG5V.n5064 ASIG5V.n3195 2.24164
R47968 ASIG5V.n4965 ASIG5V.n3223 2.24164
R47969 ASIG5V.n5064 ASIG5V.n3194 2.24164
R47970 ASIG5V.n4969 ASIG5V.n3223 2.24164
R47971 ASIG5V.n5064 ASIG5V.n3193 2.24164
R47972 ASIG5V.n4977 ASIG5V.n3223 2.24164
R47973 ASIG5V.n5064 ASIG5V.n3192 2.24164
R47974 ASIG5V.n4981 ASIG5V.n3223 2.24164
R47975 ASIG5V.n5064 ASIG5V.n3191 2.24164
R47976 ASIG5V.n4989 ASIG5V.n3223 2.24164
R47977 ASIG5V.n5064 ASIG5V.n3190 2.24164
R47978 ASIG5V.n4993 ASIG5V.n3223 2.24164
R47979 ASIG5V.n5064 ASIG5V.n3189 2.24164
R47980 ASIG5V.n5001 ASIG5V.n3223 2.24164
R47981 ASIG5V.n5064 ASIG5V.n3188 2.24164
R47982 ASIG5V.n5005 ASIG5V.n3223 2.24164
R47983 ASIG5V.n5064 ASIG5V.n3187 2.24164
R47984 ASIG5V.n5013 ASIG5V.n3223 2.24164
R47985 ASIG5V.n5064 ASIG5V.n3186 2.24164
R47986 ASIG5V.n5017 ASIG5V.n3223 2.24164
R47987 ASIG5V.n5064 ASIG5V.n3185 2.24164
R47988 ASIG5V.n5025 ASIG5V.n3223 2.24164
R47989 ASIG5V.n5064 ASIG5V.n3184 2.24164
R47990 ASIG5V.n5029 ASIG5V.n3223 2.24164
R47991 ASIG5V.n5064 ASIG5V.n3183 2.24164
R47992 ASIG5V.n5037 ASIG5V.n3223 2.24164
R47993 ASIG5V.n5064 ASIG5V.n3182 2.24164
R47994 ASIG5V.n5041 ASIG5V.n3223 2.24164
R47995 ASIG5V.n5064 ASIG5V.n3181 2.24164
R47996 ASIG5V.n5049 ASIG5V.n3223 2.24164
R47997 ASIG5V.n5064 ASIG5V.n3180 2.24164
R47998 ASIG5V.n5053 ASIG5V.n3223 2.24164
R47999 ASIG5V.n5064 ASIG5V.n3179 2.24164
R48000 ASIG5V.n5062 ASIG5V.n3223 2.24164
R48001 ASIG5V.n3613 ASIG5V.n3276 2.24164
R48002 ASIG5V.n3611 ASIG5V.n3278 2.24164
R48003 ASIG5V.n3284 ASIG5V.n3276 2.24164
R48004 ASIG5V.n3289 ASIG5V.n3278 2.24164
R48005 ASIG5V.n3603 ASIG5V.n3276 2.24164
R48006 ASIG5V.n3601 ASIG5V.n3278 2.24164
R48007 ASIG5V.n3290 ASIG5V.n3276 2.24164
R48008 ASIG5V.n3295 ASIG5V.n3278 2.24164
R48009 ASIG5V.n3593 ASIG5V.n3276 2.24164
R48010 ASIG5V.n3591 ASIG5V.n3278 2.24164
R48011 ASIG5V.n3296 ASIG5V.n3276 2.24164
R48012 ASIG5V.n3301 ASIG5V.n3278 2.24164
R48013 ASIG5V.n3583 ASIG5V.n3276 2.24164
R48014 ASIG5V.n3581 ASIG5V.n3278 2.24164
R48015 ASIG5V.n3302 ASIG5V.n3276 2.24164
R48016 ASIG5V.n3307 ASIG5V.n3278 2.24164
R48017 ASIG5V.n3573 ASIG5V.n3276 2.24164
R48018 ASIG5V.n3571 ASIG5V.n3278 2.24164
R48019 ASIG5V.n3308 ASIG5V.n3276 2.24164
R48020 ASIG5V.n3313 ASIG5V.n3278 2.24164
R48021 ASIG5V.n3563 ASIG5V.n3276 2.24164
R48022 ASIG5V.n3561 ASIG5V.n3278 2.24164
R48023 ASIG5V.n3314 ASIG5V.n3276 2.24164
R48024 ASIG5V.n3319 ASIG5V.n3278 2.24164
R48025 ASIG5V.n3553 ASIG5V.n3276 2.24164
R48026 ASIG5V.n3551 ASIG5V.n3278 2.24164
R48027 ASIG5V.n3320 ASIG5V.n3276 2.24164
R48028 ASIG5V.n3325 ASIG5V.n3278 2.24164
R48029 ASIG5V.n3543 ASIG5V.n3276 2.24164
R48030 ASIG5V.n3541 ASIG5V.n3278 2.24164
R48031 ASIG5V.n3326 ASIG5V.n3276 2.24164
R48032 ASIG5V.n3331 ASIG5V.n3278 2.24164
R48033 ASIG5V.n3533 ASIG5V.n3276 2.24164
R48034 ASIG5V.n3531 ASIG5V.n3278 2.24164
R48035 ASIG5V.n3332 ASIG5V.n3276 2.24164
R48036 ASIG5V.n3337 ASIG5V.n3278 2.24164
R48037 ASIG5V.n3523 ASIG5V.n3276 2.24164
R48038 ASIG5V.n3521 ASIG5V.n3278 2.24164
R48039 ASIG5V.n3338 ASIG5V.n3276 2.24164
R48040 ASIG5V.n3343 ASIG5V.n3278 2.24164
R48041 ASIG5V.n3513 ASIG5V.n3276 2.24164
R48042 ASIG5V.n3511 ASIG5V.n3278 2.24164
R48043 ASIG5V.n3344 ASIG5V.n3276 2.24164
R48044 ASIG5V.n3349 ASIG5V.n3278 2.24164
R48045 ASIG5V.n3503 ASIG5V.n3276 2.24164
R48046 ASIG5V.n3501 ASIG5V.n3278 2.24164
R48047 ASIG5V.n3350 ASIG5V.n3276 2.24164
R48048 ASIG5V.n3355 ASIG5V.n3278 2.24164
R48049 ASIG5V.n3493 ASIG5V.n3276 2.24164
R48050 ASIG5V.n3491 ASIG5V.n3278 2.24164
R48051 ASIG5V.n3356 ASIG5V.n3276 2.24164
R48052 ASIG5V.n3361 ASIG5V.n3278 2.24164
R48053 ASIG5V.n3483 ASIG5V.n3276 2.24164
R48054 ASIG5V.n3481 ASIG5V.n3278 2.24164
R48055 ASIG5V.n3362 ASIG5V.n3276 2.24164
R48056 ASIG5V.n3367 ASIG5V.n3278 2.24164
R48057 ASIG5V.n3473 ASIG5V.n3276 2.24164
R48058 ASIG5V.n3471 ASIG5V.n3278 2.24164
R48059 ASIG5V.n3368 ASIG5V.n3276 2.24164
R48060 ASIG5V.n3373 ASIG5V.n3278 2.24164
R48061 ASIG5V.n3463 ASIG5V.n3276 2.24164
R48062 ASIG5V.n3461 ASIG5V.n3278 2.24164
R48063 ASIG5V.n3374 ASIG5V.n3276 2.24164
R48064 ASIG5V.n3379 ASIG5V.n3278 2.24164
R48065 ASIG5V.n3453 ASIG5V.n3276 2.24164
R48066 ASIG5V.n3451 ASIG5V.n3278 2.24164
R48067 ASIG5V.n3380 ASIG5V.n3276 2.24164
R48068 ASIG5V.n3385 ASIG5V.n3278 2.24164
R48069 ASIG5V.n3443 ASIG5V.n3276 2.24164
R48070 ASIG5V.n3441 ASIG5V.n3278 2.24164
R48071 ASIG5V.n3386 ASIG5V.n3276 2.24164
R48072 ASIG5V.n3391 ASIG5V.n3278 2.24164
R48073 ASIG5V.n3433 ASIG5V.n3276 2.24164
R48074 ASIG5V.n3431 ASIG5V.n3278 2.24164
R48075 ASIG5V.n3392 ASIG5V.n3276 2.24164
R48076 ASIG5V.n3397 ASIG5V.n3278 2.24164
R48077 ASIG5V.n3423 ASIG5V.n3276 2.24164
R48078 ASIG5V.n3421 ASIG5V.n3278 2.24164
R48079 ASIG5V.n3398 ASIG5V.n3276 2.24164
R48080 ASIG5V.n3403 ASIG5V.n3278 2.24164
R48081 ASIG5V.n3413 ASIG5V.n3276 2.24164
R48082 ASIG5V.n3411 ASIG5V.n3278 2.24164
R48083 ASIG5V.n3404 ASIG5V.n3276 2.24164
R48084 ASIG5V.n4776 ASIG5V.n4774 2.24164
R48085 ASIG5V.n4772 ASIG5V.n3675 2.24164
R48086 ASIG5V.n4776 ASIG5V.n3670 2.24164
R48087 ASIG5V.n4772 ASIG5V.n3676 2.24164
R48088 ASIG5V.n4776 ASIG5V.n3669 2.24164
R48089 ASIG5V.n4772 ASIG5V.n3677 2.24164
R48090 ASIG5V.n4776 ASIG5V.n3668 2.24164
R48091 ASIG5V.n4772 ASIG5V.n3678 2.24164
R48092 ASIG5V.n4776 ASIG5V.n3667 2.24164
R48093 ASIG5V.n4772 ASIG5V.n3679 2.24164
R48094 ASIG5V.n4776 ASIG5V.n3666 2.24164
R48095 ASIG5V.n4772 ASIG5V.n3680 2.24164
R48096 ASIG5V.n4776 ASIG5V.n3665 2.24164
R48097 ASIG5V.n4772 ASIG5V.n3681 2.24164
R48098 ASIG5V.n4776 ASIG5V.n3664 2.24164
R48099 ASIG5V.n4772 ASIG5V.n3682 2.24164
R48100 ASIG5V.n4776 ASIG5V.n3663 2.24164
R48101 ASIG5V.n4772 ASIG5V.n3683 2.24164
R48102 ASIG5V.n4776 ASIG5V.n3662 2.24164
R48103 ASIG5V.n4772 ASIG5V.n3684 2.24164
R48104 ASIG5V.n4776 ASIG5V.n3661 2.24164
R48105 ASIG5V.n4772 ASIG5V.n3685 2.24164
R48106 ASIG5V.n4776 ASIG5V.n3660 2.24164
R48107 ASIG5V.n4772 ASIG5V.n3686 2.24164
R48108 ASIG5V.n4776 ASIG5V.n3659 2.24164
R48109 ASIG5V.n4772 ASIG5V.n3687 2.24164
R48110 ASIG5V.n4776 ASIG5V.n3658 2.24164
R48111 ASIG5V.n4772 ASIG5V.n3688 2.24164
R48112 ASIG5V.n4776 ASIG5V.n3657 2.24164
R48113 ASIG5V.n4772 ASIG5V.n3689 2.24164
R48114 ASIG5V.n4776 ASIG5V.n3656 2.24164
R48115 ASIG5V.n4772 ASIG5V.n3690 2.24164
R48116 ASIG5V.n4776 ASIG5V.n3655 2.24164
R48117 ASIG5V.n4772 ASIG5V.n3691 2.24164
R48118 ASIG5V.n4776 ASIG5V.n3654 2.24164
R48119 ASIG5V.n4772 ASIG5V.n3692 2.24164
R48120 ASIG5V.n4776 ASIG5V.n3653 2.24164
R48121 ASIG5V.n4772 ASIG5V.n3693 2.24164
R48122 ASIG5V.n4776 ASIG5V.n3652 2.24164
R48123 ASIG5V.n4772 ASIG5V.n3694 2.24164
R48124 ASIG5V.n4776 ASIG5V.n3651 2.24164
R48125 ASIG5V.n4772 ASIG5V.n3695 2.24164
R48126 ASIG5V.n4776 ASIG5V.n3650 2.24164
R48127 ASIG5V.n4772 ASIG5V.n3696 2.24164
R48128 ASIG5V.n4776 ASIG5V.n3649 2.24164
R48129 ASIG5V.n4772 ASIG5V.n3697 2.24164
R48130 ASIG5V.n4776 ASIG5V.n3648 2.24164
R48131 ASIG5V.n4772 ASIG5V.n3698 2.24164
R48132 ASIG5V.n4776 ASIG5V.n3647 2.24164
R48133 ASIG5V.n4772 ASIG5V.n3699 2.24164
R48134 ASIG5V.n4776 ASIG5V.n3646 2.24164
R48135 ASIG5V.n4772 ASIG5V.n3700 2.24164
R48136 ASIG5V.n4776 ASIG5V.n3645 2.24164
R48137 ASIG5V.n4772 ASIG5V.n3701 2.24164
R48138 ASIG5V.n4776 ASIG5V.n3644 2.24164
R48139 ASIG5V.n4772 ASIG5V.n3702 2.24164
R48140 ASIG5V.n4776 ASIG5V.n3643 2.24164
R48141 ASIG5V.n4772 ASIG5V.n3703 2.24164
R48142 ASIG5V.n4776 ASIG5V.n3642 2.24164
R48143 ASIG5V.n4772 ASIG5V.n3704 2.24164
R48144 ASIG5V.n4776 ASIG5V.n3641 2.24164
R48145 ASIG5V.n4772 ASIG5V.n3705 2.24164
R48146 ASIG5V.n4776 ASIG5V.n3640 2.24164
R48147 ASIG5V.n4772 ASIG5V.n3706 2.24164
R48148 ASIG5V.n4776 ASIG5V.n3639 2.24164
R48149 ASIG5V.n4772 ASIG5V.n3707 2.24164
R48150 ASIG5V.n4776 ASIG5V.n3638 2.24164
R48151 ASIG5V.n4772 ASIG5V.n3708 2.24164
R48152 ASIG5V.n4776 ASIG5V.n3637 2.24164
R48153 ASIG5V.n4772 ASIG5V.n3709 2.24164
R48154 ASIG5V.n4776 ASIG5V.n3636 2.24164
R48155 ASIG5V.n4772 ASIG5V.n3710 2.24164
R48156 ASIG5V.n4776 ASIG5V.n3635 2.24164
R48157 ASIG5V.n4772 ASIG5V.n3711 2.24164
R48158 ASIG5V.n4776 ASIG5V.n3634 2.24164
R48159 ASIG5V.n4772 ASIG5V.n3712 2.24164
R48160 ASIG5V.n4776 ASIG5V.n3633 2.24164
R48161 ASIG5V.n4772 ASIG5V.n3713 2.24164
R48162 ASIG5V.n4776 ASIG5V.n3632 2.24164
R48163 ASIG5V.n4772 ASIG5V.n3714 2.24164
R48164 ASIG5V.n4776 ASIG5V.n3631 2.24164
R48165 ASIG5V.n4772 ASIG5V.n3715 2.24164
R48166 ASIG5V.n4776 ASIG5V.n3630 2.24164
R48167 ASIG5V.n11163 ASIG5V.n11162 2.24164
R48168 ASIG5V.n11172 ASIG5V.n10414 2.24164
R48169 ASIG5V.n11163 ASIG5V.n10462 2.24164
R48170 ASIG5V.n11172 ASIG5V.n10413 2.24164
R48171 ASIG5V.n11163 ASIG5V.n10461 2.24164
R48172 ASIG5V.n11172 ASIG5V.n10412 2.24164
R48173 ASIG5V.n11163 ASIG5V.n10460 2.24164
R48174 ASIG5V.n11172 ASIG5V.n10411 2.24164
R48175 ASIG5V.n11163 ASIG5V.n10459 2.24164
R48176 ASIG5V.n11172 ASIG5V.n10410 2.24164
R48177 ASIG5V.n11163 ASIG5V.n10458 2.24164
R48178 ASIG5V.n11172 ASIG5V.n10409 2.24164
R48179 ASIG5V.n11163 ASIG5V.n10457 2.24164
R48180 ASIG5V.n11172 ASIG5V.n10408 2.24164
R48181 ASIG5V.n11163 ASIG5V.n10456 2.24164
R48182 ASIG5V.n11172 ASIG5V.n10407 2.24164
R48183 ASIG5V.n11163 ASIG5V.n10455 2.24164
R48184 ASIG5V.n11172 ASIG5V.n10406 2.24164
R48185 ASIG5V.n11163 ASIG5V.n10454 2.24164
R48186 ASIG5V.n11172 ASIG5V.n10405 2.24164
R48187 ASIG5V.n11163 ASIG5V.n10453 2.24164
R48188 ASIG5V.n11172 ASIG5V.n10404 2.24164
R48189 ASIG5V.n11163 ASIG5V.n10452 2.24164
R48190 ASIG5V.n11172 ASIG5V.n10403 2.24164
R48191 ASIG5V.n11163 ASIG5V.n10451 2.24164
R48192 ASIG5V.n11172 ASIG5V.n10402 2.24164
R48193 ASIG5V.n11163 ASIG5V.n10450 2.24164
R48194 ASIG5V.n11172 ASIG5V.n10401 2.24164
R48195 ASIG5V.n11163 ASIG5V.n10449 2.24164
R48196 ASIG5V.n11172 ASIG5V.n10400 2.24164
R48197 ASIG5V.n11163 ASIG5V.n10448 2.24164
R48198 ASIG5V.n11172 ASIG5V.n10399 2.24164
R48199 ASIG5V.n11163 ASIG5V.n10447 2.24164
R48200 ASIG5V.n11172 ASIG5V.n10398 2.24164
R48201 ASIG5V.n11163 ASIG5V.n10446 2.24164
R48202 ASIG5V.n11172 ASIG5V.n10397 2.24164
R48203 ASIG5V.n11163 ASIG5V.n10445 2.24164
R48204 ASIG5V.n11172 ASIG5V.n10396 2.24164
R48205 ASIG5V.n11163 ASIG5V.n10444 2.24164
R48206 ASIG5V.n11172 ASIG5V.n10395 2.24164
R48207 ASIG5V.n11163 ASIG5V.n10443 2.24164
R48208 ASIG5V.n11172 ASIG5V.n10394 2.24164
R48209 ASIG5V.n11163 ASIG5V.n10442 2.24164
R48210 ASIG5V.n11172 ASIG5V.n10393 2.24164
R48211 ASIG5V.n11163 ASIG5V.n10441 2.24164
R48212 ASIG5V.n11172 ASIG5V.n10392 2.24164
R48213 ASIG5V.n11163 ASIG5V.n10440 2.24164
R48214 ASIG5V.n11172 ASIG5V.n10391 2.24164
R48215 ASIG5V.n11163 ASIG5V.n10439 2.24164
R48216 ASIG5V.n11172 ASIG5V.n10390 2.24164
R48217 ASIG5V.n11163 ASIG5V.n10438 2.24164
R48218 ASIG5V.n11172 ASIG5V.n10389 2.24164
R48219 ASIG5V.n11163 ASIG5V.n10437 2.24164
R48220 ASIG5V.n11172 ASIG5V.n10388 2.24164
R48221 ASIG5V.n11163 ASIG5V.n10436 2.24164
R48222 ASIG5V.n11172 ASIG5V.n10387 2.24164
R48223 ASIG5V.n11163 ASIG5V.n10435 2.24164
R48224 ASIG5V.n11172 ASIG5V.n10386 2.24164
R48225 ASIG5V.n11163 ASIG5V.n10434 2.24164
R48226 ASIG5V.n11172 ASIG5V.n10385 2.24164
R48227 ASIG5V.n11163 ASIG5V.n10433 2.24164
R48228 ASIG5V.n11172 ASIG5V.n10384 2.24164
R48229 ASIG5V.n11163 ASIG5V.n10432 2.24164
R48230 ASIG5V.n11172 ASIG5V.n10383 2.24164
R48231 ASIG5V.n11163 ASIG5V.n10431 2.24164
R48232 ASIG5V.n11172 ASIG5V.n10382 2.24164
R48233 ASIG5V.n11163 ASIG5V.n10430 2.24164
R48234 ASIG5V.n11172 ASIG5V.n10381 2.24164
R48235 ASIG5V.n11163 ASIG5V.n10429 2.24164
R48236 ASIG5V.n11172 ASIG5V.n10380 2.24164
R48237 ASIG5V.n11163 ASIG5V.n10428 2.24164
R48238 ASIG5V.n11172 ASIG5V.n10379 2.24164
R48239 ASIG5V.n11163 ASIG5V.n10427 2.24164
R48240 ASIG5V.n11172 ASIG5V.n10378 2.24164
R48241 ASIG5V.n11163 ASIG5V.n10426 2.24164
R48242 ASIG5V.n11172 ASIG5V.n10377 2.24164
R48243 ASIG5V.n11163 ASIG5V.n10425 2.24164
R48244 ASIG5V.n11172 ASIG5V.n10376 2.24164
R48245 ASIG5V.n11163 ASIG5V.n10424 2.24164
R48246 ASIG5V.n11172 ASIG5V.n10375 2.24164
R48247 ASIG5V.n11164 ASIG5V.n11163 2.24164
R48248 ASIG5V.n11172 ASIG5V.n10374 2.24164
R48249 ASIG5V.n11163 ASIG5V.n10417 2.24164
R48250 ASIG5V.n4554 ASIG5V.n4553 2.24164
R48251 ASIG5V.n4568 ASIG5V.n3828 2.24164
R48252 ASIG5V.n4554 ASIG5V.n4308 2.24164
R48253 ASIG5V.n4568 ASIG5V.n3827 2.24164
R48254 ASIG5V.n4554 ASIG5V.n4307 2.24164
R48255 ASIG5V.n4568 ASIG5V.n3826 2.24164
R48256 ASIG5V.n4554 ASIG5V.n4306 2.24164
R48257 ASIG5V.n4568 ASIG5V.n3825 2.24164
R48258 ASIG5V.n4554 ASIG5V.n4305 2.24164
R48259 ASIG5V.n4568 ASIG5V.n3824 2.24164
R48260 ASIG5V.n4554 ASIG5V.n4304 2.24164
R48261 ASIG5V.n4568 ASIG5V.n3823 2.24164
R48262 ASIG5V.n4554 ASIG5V.n4303 2.24164
R48263 ASIG5V.n4568 ASIG5V.n3822 2.24164
R48264 ASIG5V.n4554 ASIG5V.n4302 2.24164
R48265 ASIG5V.n4568 ASIG5V.n3821 2.24164
R48266 ASIG5V.n4554 ASIG5V.n4301 2.24164
R48267 ASIG5V.n4568 ASIG5V.n3820 2.24164
R48268 ASIG5V.n4554 ASIG5V.n4300 2.24164
R48269 ASIG5V.n4568 ASIG5V.n3819 2.24164
R48270 ASIG5V.n4554 ASIG5V.n4299 2.24164
R48271 ASIG5V.n4568 ASIG5V.n3818 2.24164
R48272 ASIG5V.n4554 ASIG5V.n4298 2.24164
R48273 ASIG5V.n4568 ASIG5V.n3817 2.24164
R48274 ASIG5V.n4554 ASIG5V.n4297 2.24164
R48275 ASIG5V.n4568 ASIG5V.n3816 2.24164
R48276 ASIG5V.n4554 ASIG5V.n4296 2.24164
R48277 ASIG5V.n4568 ASIG5V.n3815 2.24164
R48278 ASIG5V.n4554 ASIG5V.n4295 2.24164
R48279 ASIG5V.n4568 ASIG5V.n3814 2.24164
R48280 ASIG5V.n4554 ASIG5V.n4294 2.24164
R48281 ASIG5V.n4568 ASIG5V.n3813 2.24164
R48282 ASIG5V.n4554 ASIG5V.n4293 2.24164
R48283 ASIG5V.n4568 ASIG5V.n3812 2.24164
R48284 ASIG5V.n4554 ASIG5V.n4292 2.24164
R48285 ASIG5V.n4568 ASIG5V.n3811 2.24164
R48286 ASIG5V.n4554 ASIG5V.n4291 2.24164
R48287 ASIG5V.n4568 ASIG5V.n3810 2.24164
R48288 ASIG5V.n4554 ASIG5V.n4290 2.24164
R48289 ASIG5V.n4568 ASIG5V.n3809 2.24164
R48290 ASIG5V.n4554 ASIG5V.n4289 2.24164
R48291 ASIG5V.n4568 ASIG5V.n3808 2.24164
R48292 ASIG5V.n4554 ASIG5V.n4288 2.24164
R48293 ASIG5V.n4568 ASIG5V.n3807 2.24164
R48294 ASIG5V.n4554 ASIG5V.n4287 2.24164
R48295 ASIG5V.n4568 ASIG5V.n3806 2.24164
R48296 ASIG5V.n4554 ASIG5V.n4286 2.24164
R48297 ASIG5V.n4568 ASIG5V.n3805 2.24164
R48298 ASIG5V.n4554 ASIG5V.n4285 2.24164
R48299 ASIG5V.n4568 ASIG5V.n3804 2.24164
R48300 ASIG5V.n4554 ASIG5V.n4284 2.24164
R48301 ASIG5V.n4568 ASIG5V.n3803 2.24164
R48302 ASIG5V.n4554 ASIG5V.n4283 2.24164
R48303 ASIG5V.n4568 ASIG5V.n3802 2.24164
R48304 ASIG5V.n4554 ASIG5V.n4282 2.24164
R48305 ASIG5V.n4568 ASIG5V.n3801 2.24164
R48306 ASIG5V.n4554 ASIG5V.n4281 2.24164
R48307 ASIG5V.n4568 ASIG5V.n3800 2.24164
R48308 ASIG5V.n4554 ASIG5V.n4280 2.24164
R48309 ASIG5V.n4568 ASIG5V.n3799 2.24164
R48310 ASIG5V.n4554 ASIG5V.n4279 2.24164
R48311 ASIG5V.n4568 ASIG5V.n3798 2.24164
R48312 ASIG5V.n4554 ASIG5V.n4278 2.24164
R48313 ASIG5V.n4568 ASIG5V.n3797 2.24164
R48314 ASIG5V.n4554 ASIG5V.n4277 2.24164
R48315 ASIG5V.n4568 ASIG5V.n3796 2.24164
R48316 ASIG5V.n4554 ASIG5V.n4276 2.24164
R48317 ASIG5V.n4568 ASIG5V.n3795 2.24164
R48318 ASIG5V.n4554 ASIG5V.n4275 2.24164
R48319 ASIG5V.n4568 ASIG5V.n3794 2.24164
R48320 ASIG5V.n4554 ASIG5V.n4274 2.24164
R48321 ASIG5V.n4568 ASIG5V.n3793 2.24164
R48322 ASIG5V.n4554 ASIG5V.n4273 2.24164
R48323 ASIG5V.n4568 ASIG5V.n3792 2.24164
R48324 ASIG5V.n4554 ASIG5V.n4272 2.24164
R48325 ASIG5V.n4568 ASIG5V.n3791 2.24164
R48326 ASIG5V.n4554 ASIG5V.n4271 2.24164
R48327 ASIG5V.n4568 ASIG5V.n3790 2.24164
R48328 ASIG5V.n4554 ASIG5V.n4270 2.24164
R48329 ASIG5V.n4568 ASIG5V.n3789 2.24164
R48330 ASIG5V.n4554 ASIG5V.n4269 2.24164
R48331 ASIG5V.n4568 ASIG5V.n3788 2.24164
R48332 ASIG5V.n4554 ASIG5V.n3832 2.24164
R48333 ASIG5V.n4268 ASIG5V.n4267 1.1255
R48334 ASIG5V.n4555 ASIG5V.n3786 1.1255
R48335 ASIG5V.n4570 ASIG5V.n4569 1.1255
R48336 ASIG5V.n4577 ASIG5V.n3781 1.1255
R48337 ASIG5V.n4578 ASIG5V.n3674 1.1255
R48338 ASIG5V.n4579 ASIG5V.n3629 1.1255
R48339 ASIG5V.n4775 ASIG5V.n3619 1.1255
R48340 ASIG5V.n4788 ASIG5V.n4787 1.1255
R48341 ASIG5V.n4789 ASIG5V.n3276 1.1255
R48342 ASIG5V.n4798 ASIG5V.n4797 1.1255
R48343 ASIG5V.n3270 ASIG5V.n3269 1.1255
R48344 ASIG5V.n4809 ASIG5V.n4808 1.1255
R48345 ASIG5V.n4811 ASIG5V.n3178 1.1255
R48346 ASIG5V.n3221 ASIG5V.n3167 1.1255
R48347 ASIG5V.n9745 ASIG5V.n9744 1.1255
R48348 ASIG5V.n5074 ASIG5V.n3168 1.1255
R48349 ASIG5V.n9441 ASIG5V.n9440 1.1255
R48350 ASIG5V.n5169 ASIG5V.n5118 1.1255
R48351 ASIG5V.n9434 ASIG5V.n9433 1.1255
R48352 ASIG5V.n7966 ASIG5V.n7963 1.1255
R48353 ASIG5V.n7967 ASIG5V.n5464 1.1255
R48354 ASIG5V.n7968 ASIG5V.n5506 1.1255
R48355 ASIG5V.n7974 ASIG5V.n5511 1.1255
R48356 ASIG5V.n7976 ASIG5V.n7975 1.1255
R48357 ASIG5V.n7979 ASIG5V.n7978 1.1255
R48358 ASIG5V.n9405 ASIG5V.n9404 1.1255
R48359 ASIG5V.n6252 ASIG5V.n5570 1.1255
R48360 ASIG5V.n9398 ASIG5V.n9397 1.1255
R48361 ASIG5V.n6418 ASIG5V.n5954 1.1255
R48362 ASIG5V.n6424 ASIG5V.n5999 1.1255
R48363 ASIG5V.n6425 ASIG5V.n6264 1.1255
R48364 ASIG5V.n6426 ASIG5V.n6306 1.1255
R48365 ASIG5V.n9188 ASIG5V.n6352 1.1255
R48366 ASIG5V.n9187 ASIG5V.n9186 1.1255
R48367 ASIG5V.n6445 ASIG5V.n6430 1.1255
R48368 ASIG5V.n6539 ASIG5V.n6488 1.1255
R48369 ASIG5V.n6544 ASIG5V.n6542 1.1255
R48370 ASIG5V.n8921 ASIG5V.n8920 1.1255
R48371 ASIG5V.n7236 ASIG5V.n6590 1.1255
R48372 ASIG5V.n7238 ASIG5V.n7237 1.1255
R48373 ASIG5V.n7241 ASIG5V.n7240 1.1255
R48374 ASIG5V.n8905 ASIG5V.n8904 1.1255
R48375 ASIG5V.n8268 ASIG5V.n6894 1.1255
R48376 ASIG5V.n8897 ASIG5V.n8896 1.1255
R48377 ASIG5V.n8213 ASIG5V.n8170 1.1255
R48378 ASIG5V.n8572 ASIG5V.n8259 1.1255
R48379 ASIG5V.n8573 ASIG5V.n8277 1.1255
R48380 ASIG5V.n8574 ASIG5V.n0 1.1255
R48381 ASIG5V.n8584 ASIG5V.n8583 1.1255
R48382 ASIG5V.n8581 ASIG5V.n10 1.1255
R48383 ASIG5V.n8580 ASIG5V.n52 1.1255
R48384 ASIG5V.n12334 ASIG5V.n56 1.1255
R48385 ASIG5V.n12333 ASIG5V.n98 1.1255
R48386 ASIG5V.n12332 ASIG5V.n166 1.1255
R48387 ASIG5V.n12325 ASIG5V.n12324 1.1255
R48388 ASIG5V.n520 ASIG5V.n172 1.1255
R48389 ASIG5V.n12310 ASIG5V.n12309 1.1255
R48390 ASIG5V.n12303 ASIG5V.n12302 1.1255
R48391 ASIG5V.n865 ASIG5V.n527 1.1255
R48392 ASIG5V.n12288 ASIG5V.n12287 1.1255
R48393 ASIG5V.n875 ASIG5V.n867 1.1255
R48394 ASIG5V.n12280 ASIG5V.n12279 1.1255
R48395 ASIG5V.n878 ASIG5V.n874 1.1255
R48396 ASIG5V.n1319 ASIG5V.n1226 1.1255
R48397 ASIG5V.n1321 ASIG5V.n1269 1.1255
R48398 ASIG5V.n1327 ASIG5V.n1324 1.1255
R48399 ASIG5V.n12013 ASIG5V.n12012 1.1255
R48400 ASIG5V.n1832 ASIG5V.n1373 1.1255
R48401 ASIG5V.n1833 ASIG5V.n1415 1.1255
R48402 ASIG5V.n1834 ASIG5V.n1675 1.1255
R48403 ASIG5V.n11803 ASIG5V.n1717 1.1255
R48404 ASIG5V.n11802 ASIG5V.n1763 1.1255
R48405 ASIG5V.n11801 ASIG5V.n1839 1.1255
R48406 ASIG5V.n2199 ASIG5V.n1838 1.1255
R48407 ASIG5V.n11793 ASIG5V.n11792 1.1255
R48408 ASIG5V.n1849 ASIG5V.n1847 1.1255
R48409 ASIG5V.n2558 ASIG5V.n2557 1.1255
R48410 ASIG5V.n2214 ASIG5V.n2212 1.1255
R48411 ASIG5V.n11781 ASIG5V.n11780 1.1255
R48412 ASIG5V.n2615 ASIG5V.n2215 1.1255
R48413 ASIG5V.n11773 ASIG5V.n11772 1.1255
R48414 ASIG5V.n2906 ASIG5V.n2568 1.1255
R48415 ASIG5V.n9958 ASIG5V.n9957 1.1255
R48416 ASIG5V.n9960 ASIG5V.n2913 1.1255
R48417 ASIG5V.n9963 ASIG5V.n2956 1.1255
R48418 ASIG5V.n11496 ASIG5V.n11495 1.1255
R48419 ASIG5V.n10017 ASIG5V.n9973 1.1255
R48420 ASIG5V.n11192 ASIG5V.n11191 1.1255
R48421 ASIG5V.n10076 ASIG5V.n10018 1.1255
R48422 ASIG5V.n11185 ASIG5V.n11184 1.1255
R48423 ASIG5V.n10473 ASIG5V.n10472 1.1255
R48424 ASIG5V.n10471 ASIG5V.n10470 1.1255
R48425 ASIG5V.n10479 ASIG5V.n10373 1.1255
R48426 ASIG5V.n10922 ASIG5V.n10416 1.1255
R48427 ASIG5V.n10921 ASIG5V.n10920 1.1255
R48428 ASIG5V.n10483 ASIG5V.n10481 1.1255
R48429 ASIG5V.n4267 ASIG5V.n4266 1.1255
R48430 ASIG5V.n3786 ASIG5V.n3785 1.1255
R48431 ASIG5V.n4571 ASIG5V.n4570 1.1255
R48432 ASIG5V.n4577 ASIG5V.n4576 1.1255
R48433 ASIG5V.n4578 ASIG5V.n3778 1.1255
R48434 ASIG5V.n4580 ASIG5V.n4579 1.1255
R48435 ASIG5V.n4582 ASIG5V.n3619 1.1255
R48436 ASIG5V.n4788 ASIG5V.n3618 1.1255
R48437 ASIG5V.n4790 ASIG5V.n4789 1.1255
R48438 ASIG5V.n4797 ASIG5V.n4796 1.1255
R48439 ASIG5V.n3281 ASIG5V.n3269 1.1255
R48440 ASIG5V.n4809 ASIG5V.n3268 1.1255
R48441 ASIG5V.n4813 ASIG5V.n4811 1.1255
R48442 ASIG5V.n3167 ASIG5V.n3165 1.1255
R48443 ASIG5V.n9746 ASIG5V.n9745 1.1255
R48444 ASIG5V.n3168 ASIG5V.n3166 1.1255
R48445 ASIG5V.n9440 ASIG5V.n9439 1.1255
R48446 ASIG5V.n5119 ASIG5V.n5118 1.1255
R48447 ASIG5V.n9435 ASIG5V.n9434 1.1255
R48448 ASIG5V.n7966 ASIG5V.n7965 1.1255
R48449 ASIG5V.n7967 ASIG5V.n7962 1.1255
R48450 ASIG5V.n7969 ASIG5V.n7968 1.1255
R48451 ASIG5V.n7974 ASIG5V.n7973 1.1255
R48452 ASIG5V.n7975 ASIG5V.n7715 1.1255
R48453 ASIG5V.n7980 ASIG5V.n7979 1.1255
R48454 ASIG5V.n9404 ASIG5V.n9403 1.1255
R48455 ASIG5V.n5572 ASIG5V.n5570 1.1255
R48456 ASIG5V.n9399 ASIG5V.n9398 1.1255
R48457 ASIG5V.n6419 ASIG5V.n6418 1.1255
R48458 ASIG5V.n6424 ASIG5V.n6423 1.1255
R48459 ASIG5V.n6425 ASIG5V.n6417 1.1255
R48460 ASIG5V.n6427 ASIG5V.n6426 1.1255
R48461 ASIG5V.n9189 ASIG5V.n9188 1.1255
R48462 ASIG5V.n9187 ASIG5V.n6429 1.1255
R48463 ASIG5V.n6536 ASIG5V.n6430 1.1255
R48464 ASIG5V.n8926 ASIG5V.n6539 1.1255
R48465 ASIG5V.n6542 ASIG5V.n6537 1.1255
R48466 ASIG5V.n8922 ASIG5V.n8921 1.1255
R48467 ASIG5V.n7236 ASIG5V.n7235 1.1255
R48468 ASIG5V.n7237 ASIG5V.n7233 1.1255
R48469 ASIG5V.n7242 ASIG5V.n7241 1.1255
R48470 ASIG5V.n8904 ASIG5V.n8903 1.1255
R48471 ASIG5V.n6896 ASIG5V.n6894 1.1255
R48472 ASIG5V.n8898 ASIG5V.n8897 1.1255
R48473 ASIG5V.n8170 ASIG5V.n8169 1.1255
R48474 ASIG5V.n8572 ASIG5V.n8571 1.1255
R48475 ASIG5V.n8573 ASIG5V.n8323 1.1255
R48476 ASIG5V.n8575 ASIG5V.n8574 1.1255
R48477 ASIG5V.n8585 ASIG5V.n8584 1.1255
R48478 ASIG5V.n8581 ASIG5V.n8578 1.1255
R48479 ASIG5V.n8580 ASIG5V.n8579 1.1255
R48480 ASIG5V.n12335 ASIG5V.n12334 1.1255
R48481 ASIG5V.n12333 ASIG5V.n164 1.1255
R48482 ASIG5V.n12332 ASIG5V.n12331 1.1255
R48483 ASIG5V.n12326 ASIG5V.n12325 1.1255
R48484 ASIG5V.n172 ASIG5V.n171 1.1255
R48485 ASIG5V.n12309 ASIG5V.n12308 1.1255
R48486 ASIG5V.n12304 ASIG5V.n12303 1.1255
R48487 ASIG5V.n527 ASIG5V.n526 1.1255
R48488 ASIG5V.n12287 ASIG5V.n12286 1.1255
R48489 ASIG5V.n868 ASIG5V.n867 1.1255
R48490 ASIG5V.n12281 ASIG5V.n12280 1.1255
R48491 ASIG5V.n874 ASIG5V.n872 1.1255
R48492 ASIG5V.n1319 ASIG5V.n1317 1.1255
R48493 ASIG5V.n12018 ASIG5V.n1321 1.1255
R48494 ASIG5V.n1324 ASIG5V.n1318 1.1255
R48495 ASIG5V.n12014 ASIG5V.n12013 1.1255
R48496 ASIG5V.n1832 ASIG5V.n1831 1.1255
R48497 ASIG5V.n1833 ASIG5V.n1828 1.1255
R48498 ASIG5V.n1835 ASIG5V.n1834 1.1255
R48499 ASIG5V.n11804 ASIG5V.n11803 1.1255
R48500 ASIG5V.n11802 ASIG5V.n1837 1.1255
R48501 ASIG5V.n11801 ASIG5V.n11800 1.1255
R48502 ASIG5V.n1840 ASIG5V.n1838 1.1255
R48503 ASIG5V.n11794 ASIG5V.n11793 1.1255
R48504 ASIG5V.n1847 ASIG5V.n1845 1.1255
R48505 ASIG5V.n2559 ASIG5V.n2558 1.1255
R48506 ASIG5V.n2216 ASIG5V.n2214 1.1255
R48507 ASIG5V.n11780 ASIG5V.n11779 1.1255
R48508 ASIG5V.n2217 ASIG5V.n2215 1.1255
R48509 ASIG5V.n11774 ASIG5V.n11773 1.1255
R48510 ASIG5V.n2568 ASIG5V.n2566 1.1255
R48511 ASIG5V.n9958 ASIG5V.n9955 1.1255
R48512 ASIG5V.n11501 ASIG5V.n9960 1.1255
R48513 ASIG5V.n9963 ASIG5V.n9956 1.1255
R48514 ASIG5V.n11497 ASIG5V.n11496 1.1255
R48515 ASIG5V.n10019 ASIG5V.n10017 1.1255
R48516 ASIG5V.n11191 ASIG5V.n11190 1.1255
R48517 ASIG5V.n10020 ASIG5V.n10018 1.1255
R48518 ASIG5V.n11186 ASIG5V.n11185 1.1255
R48519 ASIG5V.n10474 ASIG5V.n10473 1.1255
R48520 ASIG5V.n10477 ASIG5V.n10470 1.1255
R48521 ASIG5V.n10479 ASIG5V.n10478 1.1255
R48522 ASIG5V.n10923 ASIG5V.n10922 1.1255
R48523 ASIG5V.n10921 ASIG5V.n10469 1.1255
R48524 ASIG5V.n10707 ASIG5V.n10481 1.1255
R48525 ASIG5V.n10708 ASIG5V.n10707 1.1255
R48526 ASIG5V.n10469 ASIG5V.n10467 1.1255
R48527 ASIG5V.n10924 ASIG5V.n10923 1.1255
R48528 ASIG5V.n10478 ASIG5V.n10466 1.1255
R48529 ASIG5V.n10477 ASIG5V.n10476 1.1255
R48530 ASIG5V.n10475 ASIG5V.n10474 1.1255
R48531 ASIG5V.n11187 ASIG5V.n11186 1.1255
R48532 ASIG5V.n11188 ASIG5V.n10020 1.1255
R48533 ASIG5V.n11190 ASIG5V.n11189 1.1255
R48534 ASIG5V.n10021 ASIG5V.n10019 1.1255
R48535 ASIG5V.n11498 ASIG5V.n11497 1.1255
R48536 ASIG5V.n11499 ASIG5V.n9956 1.1255
R48537 ASIG5V.n11501 ASIG5V.n11500 1.1255
R48538 ASIG5V.n9955 ASIG5V.n9954 1.1255
R48539 ASIG5V.n2566 ASIG5V.n2564 1.1255
R48540 ASIG5V.n11775 ASIG5V.n11774 1.1255
R48541 ASIG5V.n11777 ASIG5V.n2217 1.1255
R48542 ASIG5V.n11779 ASIG5V.n11778 1.1255
R48543 ASIG5V.n2562 ASIG5V.n2216 1.1255
R48544 ASIG5V.n2560 ASIG5V.n2559 1.1255
R48545 ASIG5V.n1845 ASIG5V.n1843 1.1255
R48546 ASIG5V.n11795 ASIG5V.n11794 1.1255
R48547 ASIG5V.n11797 ASIG5V.n1840 1.1255
R48548 ASIG5V.n11800 ASIG5V.n11799 1.1255
R48549 ASIG5V.n1837 ASIG5V.n1827 1.1255
R48550 ASIG5V.n11805 ASIG5V.n11804 1.1255
R48551 ASIG5V.n1835 ASIG5V.n1826 1.1255
R48552 ASIG5V.n1829 ASIG5V.n1828 1.1255
R48553 ASIG5V.n1831 ASIG5V.n1830 1.1255
R48554 ASIG5V.n12015 ASIG5V.n12014 1.1255
R48555 ASIG5V.n12016 ASIG5V.n1318 1.1255
R48556 ASIG5V.n12018 ASIG5V.n12017 1.1255
R48557 ASIG5V.n7339 ASIG5V.n1317 1.1255
R48558 ASIG5V.n872 ASIG5V.n870 1.1255
R48559 ASIG5V.n12282 ASIG5V.n12281 1.1255
R48560 ASIG5V.n12284 ASIG5V.n868 1.1255
R48561 ASIG5V.n12286 ASIG5V.n12285 1.1255
R48562 ASIG5V.n526 ASIG5V.n525 1.1255
R48563 ASIG5V.n12305 ASIG5V.n12304 1.1255
R48564 ASIG5V.n12308 ASIG5V.n12307 1.1255
R48565 ASIG5V.n171 ASIG5V.n170 1.1255
R48566 ASIG5V.n12327 ASIG5V.n12326 1.1255
R48567 ASIG5V.n12331 ASIG5V.n12330 1.1255
R48568 ASIG5V.n164 ASIG5V.n162 1.1255
R48569 ASIG5V.n12336 ASIG5V.n12335 1.1255
R48570 ASIG5V.n8579 ASIG5V.n161 1.1255
R48571 ASIG5V.n8578 ASIG5V.n8577 1.1255
R48572 ASIG5V.n8586 ASIG5V.n8585 1.1255
R48573 ASIG5V.n8576 ASIG5V.n8575 1.1255
R48574 ASIG5V.n8323 ASIG5V.n8322 1.1255
R48575 ASIG5V.n8571 ASIG5V.n8570 1.1255
R48576 ASIG5V.n8169 ASIG5V.n8168 1.1255
R48577 ASIG5V.n8899 ASIG5V.n8898 1.1255
R48578 ASIG5V.n8900 ASIG5V.n6896 1.1255
R48579 ASIG5V.n8903 ASIG5V.n8902 1.1255
R48580 ASIG5V.n7243 ASIG5V.n7242 1.1255
R48581 ASIG5V.n7233 ASIG5V.n7232 1.1255
R48582 ASIG5V.n7235 ASIG5V.n7234 1.1255
R48583 ASIG5V.n8923 ASIG5V.n8922 1.1255
R48584 ASIG5V.n8924 ASIG5V.n6537 1.1255
R48585 ASIG5V.n8926 ASIG5V.n8925 1.1255
R48586 ASIG5V.n6536 ASIG5V.n6535 1.1255
R48587 ASIG5V.n6534 ASIG5V.n6429 1.1255
R48588 ASIG5V.n9190 ASIG5V.n9189 1.1255
R48589 ASIG5V.n6427 ASIG5V.n6415 1.1255
R48590 ASIG5V.n6421 ASIG5V.n6417 1.1255
R48591 ASIG5V.n6423 ASIG5V.n6422 1.1255
R48592 ASIG5V.n6420 ASIG5V.n6419 1.1255
R48593 ASIG5V.n9400 ASIG5V.n9399 1.1255
R48594 ASIG5V.n9401 ASIG5V.n5572 1.1255
R48595 ASIG5V.n9403 ASIG5V.n9402 1.1255
R48596 ASIG5V.n7981 ASIG5V.n7980 1.1255
R48597 ASIG5V.n7715 ASIG5V.n7714 1.1255
R48598 ASIG5V.n7973 ASIG5V.n7972 1.1255
R48599 ASIG5V.n7970 ASIG5V.n7969 1.1255
R48600 ASIG5V.n7962 ASIG5V.n7961 1.1255
R48601 ASIG5V.n7965 ASIG5V.n7964 1.1255
R48602 ASIG5V.n9436 ASIG5V.n9435 1.1255
R48603 ASIG5V.n9437 ASIG5V.n5119 1.1255
R48604 ASIG5V.n9439 ASIG5V.n9438 1.1255
R48605 ASIG5V.n3166 ASIG5V.n3164 1.1255
R48606 ASIG5V.n9747 ASIG5V.n9746 1.1255
R48607 ASIG5V.n3165 ASIG5V.n3163 1.1255
R48608 ASIG5V.n4813 ASIG5V.n4812 1.1255
R48609 ASIG5V.n4793 ASIG5V.n3268 1.1255
R48610 ASIG5V.n4794 ASIG5V.n3281 1.1255
R48611 ASIG5V.n4796 ASIG5V.n4795 1.1255
R48612 ASIG5V.n4791 ASIG5V.n4790 1.1255
R48613 ASIG5V.n3618 ASIG5V.n3617 1.1255
R48614 ASIG5V.n4583 ASIG5V.n4582 1.1255
R48615 ASIG5V.n4580 ASIG5V.n3777 1.1255
R48616 ASIG5V.n4574 ASIG5V.n3778 1.1255
R48617 ASIG5V.n4576 ASIG5V.n4575 1.1255
R48618 ASIG5V.n4572 ASIG5V.n4571 1.1255
R48619 ASIG5V.n3785 ASIG5V.n3784 1.1255
R48620 ASIG5V.n4266 ASIG5V.n4265 1.1255
R48621 ASIG5V.n10914 ASIG5V.n10913 0.902975
R48622 ASIG5V.n4248 ASIG5V.n4247 0.902975
R48623 ASIG5V.n10814 ASIG5V.n10812 0.9005
R48624 ASIG5V.n10815 ASIG5V.n10811 0.9005
R48625 ASIG5V.n10816 ASIG5V.n10810 0.9005
R48626 ASIG5V.n10817 ASIG5V.n10809 0.9005
R48627 ASIG5V.n10818 ASIG5V.n10808 0.9005
R48628 ASIG5V.n10819 ASIG5V.n10807 0.9005
R48629 ASIG5V.n10820 ASIG5V.n10806 0.9005
R48630 ASIG5V.n10821 ASIG5V.n10805 0.9005
R48631 ASIG5V.n10822 ASIG5V.n10804 0.9005
R48632 ASIG5V.n10823 ASIG5V.n10803 0.9005
R48633 ASIG5V.n10824 ASIG5V.n10802 0.9005
R48634 ASIG5V.n10825 ASIG5V.n10801 0.9005
R48635 ASIG5V.n10826 ASIG5V.n10800 0.9005
R48636 ASIG5V.n10827 ASIG5V.n10799 0.9005
R48637 ASIG5V.n10828 ASIG5V.n10798 0.9005
R48638 ASIG5V.n10829 ASIG5V.n10797 0.9005
R48639 ASIG5V.n10830 ASIG5V.n10796 0.9005
R48640 ASIG5V.n10831 ASIG5V.n10795 0.9005
R48641 ASIG5V.n10832 ASIG5V.n10794 0.9005
R48642 ASIG5V.n10833 ASIG5V.n10793 0.9005
R48643 ASIG5V.n10834 ASIG5V.n10792 0.9005
R48644 ASIG5V.n10835 ASIG5V.n10791 0.9005
R48645 ASIG5V.n10836 ASIG5V.n10790 0.9005
R48646 ASIG5V.n10837 ASIG5V.n10789 0.9005
R48647 ASIG5V.n10838 ASIG5V.n10788 0.9005
R48648 ASIG5V.n10839 ASIG5V.n10787 0.9005
R48649 ASIG5V.n10840 ASIG5V.n10786 0.9005
R48650 ASIG5V.n10841 ASIG5V.n10785 0.9005
R48651 ASIG5V.n10842 ASIG5V.n10784 0.9005
R48652 ASIG5V.n10843 ASIG5V.n10783 0.9005
R48653 ASIG5V.n10844 ASIG5V.n10782 0.9005
R48654 ASIG5V.n10845 ASIG5V.n10781 0.9005
R48655 ASIG5V.n10846 ASIG5V.n10780 0.9005
R48656 ASIG5V.n10847 ASIG5V.n10779 0.9005
R48657 ASIG5V.n10848 ASIG5V.n10778 0.9005
R48658 ASIG5V.n10849 ASIG5V.n10777 0.9005
R48659 ASIG5V.n10850 ASIG5V.n10776 0.9005
R48660 ASIG5V.n10851 ASIG5V.n10775 0.9005
R48661 ASIG5V.n10852 ASIG5V.n10774 0.9005
R48662 ASIG5V.n10853 ASIG5V.n10773 0.9005
R48663 ASIG5V.n10854 ASIG5V.n10772 0.9005
R48664 ASIG5V.n10855 ASIG5V.n10771 0.9005
R48665 ASIG5V.n10856 ASIG5V.n10770 0.9005
R48666 ASIG5V.n10857 ASIG5V.n10769 0.9005
R48667 ASIG5V.n10858 ASIG5V.n10768 0.9005
R48668 ASIG5V.n10859 ASIG5V.n10767 0.9005
R48669 ASIG5V.n10860 ASIG5V.n10766 0.9005
R48670 ASIG5V.n10861 ASIG5V.n10765 0.9005
R48671 ASIG5V.n10862 ASIG5V.n10764 0.9005
R48672 ASIG5V.n10863 ASIG5V.n10763 0.9005
R48673 ASIG5V.n10864 ASIG5V.n10762 0.9005
R48674 ASIG5V.n10865 ASIG5V.n10761 0.9005
R48675 ASIG5V.n10866 ASIG5V.n10760 0.9005
R48676 ASIG5V.n10867 ASIG5V.n10759 0.9005
R48677 ASIG5V.n10868 ASIG5V.n10758 0.9005
R48678 ASIG5V.n10869 ASIG5V.n10757 0.9005
R48679 ASIG5V.n10870 ASIG5V.n10756 0.9005
R48680 ASIG5V.n10871 ASIG5V.n10755 0.9005
R48681 ASIG5V.n10872 ASIG5V.n10754 0.9005
R48682 ASIG5V.n10873 ASIG5V.n10753 0.9005
R48683 ASIG5V.n10874 ASIG5V.n10752 0.9005
R48684 ASIG5V.n10875 ASIG5V.n10751 0.9005
R48685 ASIG5V.n10876 ASIG5V.n10750 0.9005
R48686 ASIG5V.n10877 ASIG5V.n10749 0.9005
R48687 ASIG5V.n10878 ASIG5V.n10748 0.9005
R48688 ASIG5V.n10879 ASIG5V.n10747 0.9005
R48689 ASIG5V.n10880 ASIG5V.n10746 0.9005
R48690 ASIG5V.n10881 ASIG5V.n10745 0.9005
R48691 ASIG5V.n10882 ASIG5V.n10744 0.9005
R48692 ASIG5V.n10883 ASIG5V.n10743 0.9005
R48693 ASIG5V.n10884 ASIG5V.n10742 0.9005
R48694 ASIG5V.n10885 ASIG5V.n10741 0.9005
R48695 ASIG5V.n10886 ASIG5V.n10740 0.9005
R48696 ASIG5V.n10887 ASIG5V.n10739 0.9005
R48697 ASIG5V.n10888 ASIG5V.n10738 0.9005
R48698 ASIG5V.n10889 ASIG5V.n10737 0.9005
R48699 ASIG5V.n10890 ASIG5V.n10736 0.9005
R48700 ASIG5V.n10891 ASIG5V.n10735 0.9005
R48701 ASIG5V.n10892 ASIG5V.n10734 0.9005
R48702 ASIG5V.n10893 ASIG5V.n10733 0.9005
R48703 ASIG5V.n10894 ASIG5V.n10732 0.9005
R48704 ASIG5V.n10895 ASIG5V.n10731 0.9005
R48705 ASIG5V.n10896 ASIG5V.n10730 0.9005
R48706 ASIG5V.n10897 ASIG5V.n10729 0.9005
R48707 ASIG5V.n10898 ASIG5V.n10728 0.9005
R48708 ASIG5V.n10899 ASIG5V.n10727 0.9005
R48709 ASIG5V.n10900 ASIG5V.n10726 0.9005
R48710 ASIG5V.n10901 ASIG5V.n10725 0.9005
R48711 ASIG5V.n10902 ASIG5V.n10724 0.9005
R48712 ASIG5V.n10903 ASIG5V.n10723 0.9005
R48713 ASIG5V.n10904 ASIG5V.n10722 0.9005
R48714 ASIG5V.n10905 ASIG5V.n10721 0.9005
R48715 ASIG5V.n10906 ASIG5V.n10720 0.9005
R48716 ASIG5V.n10907 ASIG5V.n10719 0.9005
R48717 ASIG5V.n10908 ASIG5V.n10718 0.9005
R48718 ASIG5V.n10909 ASIG5V.n10717 0.9005
R48719 ASIG5V.n10716 ASIG5V.n10692 0.9005
R48720 ASIG5V.n10813 ASIG5V.n10489 0.9005
R48721 ASIG5V.n10813 ASIG5V.n10548 0.9005
R48722 ASIG5V.n10814 ASIG5V.n10545 0.9005
R48723 ASIG5V.n10815 ASIG5V.n10551 0.9005
R48724 ASIG5V.n10816 ASIG5V.n10544 0.9005
R48725 ASIG5V.n10817 ASIG5V.n10554 0.9005
R48726 ASIG5V.n10818 ASIG5V.n10543 0.9005
R48727 ASIG5V.n10819 ASIG5V.n10557 0.9005
R48728 ASIG5V.n10820 ASIG5V.n10542 0.9005
R48729 ASIG5V.n10821 ASIG5V.n10560 0.9005
R48730 ASIG5V.n10822 ASIG5V.n10541 0.9005
R48731 ASIG5V.n10823 ASIG5V.n10563 0.9005
R48732 ASIG5V.n10824 ASIG5V.n10540 0.9005
R48733 ASIG5V.n10825 ASIG5V.n10566 0.9005
R48734 ASIG5V.n10826 ASIG5V.n10539 0.9005
R48735 ASIG5V.n10827 ASIG5V.n10569 0.9005
R48736 ASIG5V.n10828 ASIG5V.n10538 0.9005
R48737 ASIG5V.n10829 ASIG5V.n10572 0.9005
R48738 ASIG5V.n10830 ASIG5V.n10537 0.9005
R48739 ASIG5V.n10831 ASIG5V.n10575 0.9005
R48740 ASIG5V.n10832 ASIG5V.n10536 0.9005
R48741 ASIG5V.n10833 ASIG5V.n10578 0.9005
R48742 ASIG5V.n10834 ASIG5V.n10535 0.9005
R48743 ASIG5V.n10835 ASIG5V.n10581 0.9005
R48744 ASIG5V.n10836 ASIG5V.n10534 0.9005
R48745 ASIG5V.n10837 ASIG5V.n10584 0.9005
R48746 ASIG5V.n10838 ASIG5V.n10533 0.9005
R48747 ASIG5V.n10839 ASIG5V.n10587 0.9005
R48748 ASIG5V.n10840 ASIG5V.n10532 0.9005
R48749 ASIG5V.n10841 ASIG5V.n10590 0.9005
R48750 ASIG5V.n10842 ASIG5V.n10531 0.9005
R48751 ASIG5V.n10843 ASIG5V.n10593 0.9005
R48752 ASIG5V.n10844 ASIG5V.n10530 0.9005
R48753 ASIG5V.n10845 ASIG5V.n10596 0.9005
R48754 ASIG5V.n10846 ASIG5V.n10529 0.9005
R48755 ASIG5V.n10847 ASIG5V.n10599 0.9005
R48756 ASIG5V.n10848 ASIG5V.n10528 0.9005
R48757 ASIG5V.n10849 ASIG5V.n10602 0.9005
R48758 ASIG5V.n10850 ASIG5V.n10527 0.9005
R48759 ASIG5V.n10851 ASIG5V.n10605 0.9005
R48760 ASIG5V.n10852 ASIG5V.n10526 0.9005
R48761 ASIG5V.n10853 ASIG5V.n10608 0.9005
R48762 ASIG5V.n10854 ASIG5V.n10525 0.9005
R48763 ASIG5V.n10855 ASIG5V.n10611 0.9005
R48764 ASIG5V.n10856 ASIG5V.n10524 0.9005
R48765 ASIG5V.n10857 ASIG5V.n10614 0.9005
R48766 ASIG5V.n10858 ASIG5V.n10523 0.9005
R48767 ASIG5V.n10859 ASIG5V.n10617 0.9005
R48768 ASIG5V.n10860 ASIG5V.n10522 0.9005
R48769 ASIG5V.n10861 ASIG5V.n10620 0.9005
R48770 ASIG5V.n10862 ASIG5V.n10521 0.9005
R48771 ASIG5V.n10863 ASIG5V.n10623 0.9005
R48772 ASIG5V.n10864 ASIG5V.n10520 0.9005
R48773 ASIG5V.n10865 ASIG5V.n10626 0.9005
R48774 ASIG5V.n10866 ASIG5V.n10519 0.9005
R48775 ASIG5V.n10867 ASIG5V.n10629 0.9005
R48776 ASIG5V.n10868 ASIG5V.n10518 0.9005
R48777 ASIG5V.n10869 ASIG5V.n10632 0.9005
R48778 ASIG5V.n10870 ASIG5V.n10517 0.9005
R48779 ASIG5V.n10871 ASIG5V.n10635 0.9005
R48780 ASIG5V.n10872 ASIG5V.n10516 0.9005
R48781 ASIG5V.n10873 ASIG5V.n10638 0.9005
R48782 ASIG5V.n10874 ASIG5V.n10515 0.9005
R48783 ASIG5V.n10875 ASIG5V.n10641 0.9005
R48784 ASIG5V.n10876 ASIG5V.n10514 0.9005
R48785 ASIG5V.n10877 ASIG5V.n10644 0.9005
R48786 ASIG5V.n10878 ASIG5V.n10513 0.9005
R48787 ASIG5V.n10879 ASIG5V.n10647 0.9005
R48788 ASIG5V.n10880 ASIG5V.n10512 0.9005
R48789 ASIG5V.n10881 ASIG5V.n10650 0.9005
R48790 ASIG5V.n10882 ASIG5V.n10511 0.9005
R48791 ASIG5V.n10883 ASIG5V.n10653 0.9005
R48792 ASIG5V.n10884 ASIG5V.n10510 0.9005
R48793 ASIG5V.n10885 ASIG5V.n10656 0.9005
R48794 ASIG5V.n10886 ASIG5V.n10509 0.9005
R48795 ASIG5V.n10887 ASIG5V.n10659 0.9005
R48796 ASIG5V.n10888 ASIG5V.n10508 0.9005
R48797 ASIG5V.n10889 ASIG5V.n10662 0.9005
R48798 ASIG5V.n10890 ASIG5V.n10507 0.9005
R48799 ASIG5V.n10891 ASIG5V.n10665 0.9005
R48800 ASIG5V.n10892 ASIG5V.n10506 0.9005
R48801 ASIG5V.n10893 ASIG5V.n10668 0.9005
R48802 ASIG5V.n10894 ASIG5V.n10505 0.9005
R48803 ASIG5V.n10895 ASIG5V.n10671 0.9005
R48804 ASIG5V.n10896 ASIG5V.n10504 0.9005
R48805 ASIG5V.n10897 ASIG5V.n10674 0.9005
R48806 ASIG5V.n10898 ASIG5V.n10503 0.9005
R48807 ASIG5V.n10899 ASIG5V.n10677 0.9005
R48808 ASIG5V.n10900 ASIG5V.n10502 0.9005
R48809 ASIG5V.n10901 ASIG5V.n10680 0.9005
R48810 ASIG5V.n10902 ASIG5V.n10501 0.9005
R48811 ASIG5V.n10903 ASIG5V.n10683 0.9005
R48812 ASIG5V.n10904 ASIG5V.n10500 0.9005
R48813 ASIG5V.n10905 ASIG5V.n10686 0.9005
R48814 ASIG5V.n10906 ASIG5V.n10499 0.9005
R48815 ASIG5V.n10907 ASIG5V.n10689 0.9005
R48816 ASIG5V.n10908 ASIG5V.n10498 0.9005
R48817 ASIG5V.n10910 ASIG5V.n10909 0.9005
R48818 ASIG5V.n10692 ASIG5V.n10497 0.9005
R48819 ASIG5V.n10913 ASIG5V.n10912 0.9005
R48820 ASIG5V.n4101 ASIG5V.n3856 0.9005
R48821 ASIG5V.n4103 ASIG5V.n4102 0.9005
R48822 ASIG5V.n4104 ASIG5V.n4100 0.9005
R48823 ASIG5V.n4106 ASIG5V.n4105 0.9005
R48824 ASIG5V.n4107 ASIG5V.n4099 0.9005
R48825 ASIG5V.n4109 ASIG5V.n4108 0.9005
R48826 ASIG5V.n4110 ASIG5V.n4098 0.9005
R48827 ASIG5V.n4112 ASIG5V.n4111 0.9005
R48828 ASIG5V.n4113 ASIG5V.n4097 0.9005
R48829 ASIG5V.n4115 ASIG5V.n4114 0.9005
R48830 ASIG5V.n4116 ASIG5V.n4096 0.9005
R48831 ASIG5V.n4118 ASIG5V.n4117 0.9005
R48832 ASIG5V.n4119 ASIG5V.n4095 0.9005
R48833 ASIG5V.n4121 ASIG5V.n4120 0.9005
R48834 ASIG5V.n4122 ASIG5V.n4094 0.9005
R48835 ASIG5V.n4124 ASIG5V.n4123 0.9005
R48836 ASIG5V.n4125 ASIG5V.n4093 0.9005
R48837 ASIG5V.n4127 ASIG5V.n4126 0.9005
R48838 ASIG5V.n4128 ASIG5V.n4092 0.9005
R48839 ASIG5V.n4130 ASIG5V.n4129 0.9005
R48840 ASIG5V.n4131 ASIG5V.n4091 0.9005
R48841 ASIG5V.n4133 ASIG5V.n4132 0.9005
R48842 ASIG5V.n4134 ASIG5V.n4090 0.9005
R48843 ASIG5V.n4136 ASIG5V.n4135 0.9005
R48844 ASIG5V.n4137 ASIG5V.n4089 0.9005
R48845 ASIG5V.n4139 ASIG5V.n4138 0.9005
R48846 ASIG5V.n4140 ASIG5V.n4088 0.9005
R48847 ASIG5V.n4142 ASIG5V.n4141 0.9005
R48848 ASIG5V.n4143 ASIG5V.n4087 0.9005
R48849 ASIG5V.n4145 ASIG5V.n4144 0.9005
R48850 ASIG5V.n4146 ASIG5V.n4086 0.9005
R48851 ASIG5V.n4148 ASIG5V.n4147 0.9005
R48852 ASIG5V.n4149 ASIG5V.n4085 0.9005
R48853 ASIG5V.n4151 ASIG5V.n4150 0.9005
R48854 ASIG5V.n4152 ASIG5V.n4084 0.9005
R48855 ASIG5V.n4154 ASIG5V.n4153 0.9005
R48856 ASIG5V.n4155 ASIG5V.n4083 0.9005
R48857 ASIG5V.n4157 ASIG5V.n4156 0.9005
R48858 ASIG5V.n4158 ASIG5V.n4082 0.9005
R48859 ASIG5V.n4160 ASIG5V.n4159 0.9005
R48860 ASIG5V.n4161 ASIG5V.n4081 0.9005
R48861 ASIG5V.n4163 ASIG5V.n4162 0.9005
R48862 ASIG5V.n4164 ASIG5V.n4080 0.9005
R48863 ASIG5V.n4166 ASIG5V.n4165 0.9005
R48864 ASIG5V.n4167 ASIG5V.n4079 0.9005
R48865 ASIG5V.n4169 ASIG5V.n4168 0.9005
R48866 ASIG5V.n4170 ASIG5V.n4078 0.9005
R48867 ASIG5V.n4172 ASIG5V.n4171 0.9005
R48868 ASIG5V.n4173 ASIG5V.n4077 0.9005
R48869 ASIG5V.n4175 ASIG5V.n4174 0.9005
R48870 ASIG5V.n4176 ASIG5V.n4076 0.9005
R48871 ASIG5V.n4178 ASIG5V.n4177 0.9005
R48872 ASIG5V.n4179 ASIG5V.n4075 0.9005
R48873 ASIG5V.n4181 ASIG5V.n4180 0.9005
R48874 ASIG5V.n4182 ASIG5V.n4074 0.9005
R48875 ASIG5V.n4184 ASIG5V.n4183 0.9005
R48876 ASIG5V.n4185 ASIG5V.n4073 0.9005
R48877 ASIG5V.n4187 ASIG5V.n4186 0.9005
R48878 ASIG5V.n4188 ASIG5V.n4072 0.9005
R48879 ASIG5V.n4190 ASIG5V.n4189 0.9005
R48880 ASIG5V.n4191 ASIG5V.n4071 0.9005
R48881 ASIG5V.n4193 ASIG5V.n4192 0.9005
R48882 ASIG5V.n4194 ASIG5V.n4070 0.9005
R48883 ASIG5V.n4196 ASIG5V.n4195 0.9005
R48884 ASIG5V.n4197 ASIG5V.n4069 0.9005
R48885 ASIG5V.n4199 ASIG5V.n4198 0.9005
R48886 ASIG5V.n4200 ASIG5V.n4068 0.9005
R48887 ASIG5V.n4202 ASIG5V.n4201 0.9005
R48888 ASIG5V.n4203 ASIG5V.n4067 0.9005
R48889 ASIG5V.n4205 ASIG5V.n4204 0.9005
R48890 ASIG5V.n4206 ASIG5V.n4066 0.9005
R48891 ASIG5V.n4208 ASIG5V.n4207 0.9005
R48892 ASIG5V.n4209 ASIG5V.n4065 0.9005
R48893 ASIG5V.n4211 ASIG5V.n4210 0.9005
R48894 ASIG5V.n4212 ASIG5V.n4064 0.9005
R48895 ASIG5V.n4214 ASIG5V.n4213 0.9005
R48896 ASIG5V.n4215 ASIG5V.n4063 0.9005
R48897 ASIG5V.n4217 ASIG5V.n4216 0.9005
R48898 ASIG5V.n4218 ASIG5V.n4062 0.9005
R48899 ASIG5V.n4220 ASIG5V.n4219 0.9005
R48900 ASIG5V.n4221 ASIG5V.n4061 0.9005
R48901 ASIG5V.n4223 ASIG5V.n4222 0.9005
R48902 ASIG5V.n4224 ASIG5V.n4060 0.9005
R48903 ASIG5V.n4226 ASIG5V.n4225 0.9005
R48904 ASIG5V.n4227 ASIG5V.n4059 0.9005
R48905 ASIG5V.n4229 ASIG5V.n4228 0.9005
R48906 ASIG5V.n4230 ASIG5V.n4058 0.9005
R48907 ASIG5V.n4232 ASIG5V.n4231 0.9005
R48908 ASIG5V.n4233 ASIG5V.n4057 0.9005
R48909 ASIG5V.n4235 ASIG5V.n4234 0.9005
R48910 ASIG5V.n4236 ASIG5V.n4056 0.9005
R48911 ASIG5V.n4238 ASIG5V.n4237 0.9005
R48912 ASIG5V.n4239 ASIG5V.n4055 0.9005
R48913 ASIG5V.n4241 ASIG5V.n4240 0.9005
R48914 ASIG5V.n4242 ASIG5V.n4054 0.9005
R48915 ASIG5V.n4244 ASIG5V.n4243 0.9005
R48916 ASIG5V.n4245 ASIG5V.n4053 0.9005
R48917 ASIG5V.n4252 ASIG5V.n4246 0.9005
R48918 ASIG5V.n4247 ASIG5V.n3909 0.9005
R48919 ASIG5V.n4053 ASIG5V.n3908 0.9005
R48920 ASIG5V.n4256 ASIG5V.n3856 0.9005
R48921 ASIG5V.n4103 ASIG5V.n3906 0.9005
R48922 ASIG5V.n4104 ASIG5V.n3911 0.9005
R48923 ASIG5V.n4105 ASIG5V.n3905 0.9005
R48924 ASIG5V.n4099 ASIG5V.n3913 0.9005
R48925 ASIG5V.n4109 ASIG5V.n3904 0.9005
R48926 ASIG5V.n4110 ASIG5V.n3915 0.9005
R48927 ASIG5V.n4111 ASIG5V.n3903 0.9005
R48928 ASIG5V.n4097 ASIG5V.n3917 0.9005
R48929 ASIG5V.n4115 ASIG5V.n3902 0.9005
R48930 ASIG5V.n4116 ASIG5V.n3919 0.9005
R48931 ASIG5V.n4117 ASIG5V.n3901 0.9005
R48932 ASIG5V.n4095 ASIG5V.n3921 0.9005
R48933 ASIG5V.n4121 ASIG5V.n3900 0.9005
R48934 ASIG5V.n4122 ASIG5V.n3923 0.9005
R48935 ASIG5V.n4123 ASIG5V.n3899 0.9005
R48936 ASIG5V.n4093 ASIG5V.n3925 0.9005
R48937 ASIG5V.n4127 ASIG5V.n3898 0.9005
R48938 ASIG5V.n4128 ASIG5V.n3927 0.9005
R48939 ASIG5V.n4129 ASIG5V.n3897 0.9005
R48940 ASIG5V.n4091 ASIG5V.n3929 0.9005
R48941 ASIG5V.n4133 ASIG5V.n3896 0.9005
R48942 ASIG5V.n4134 ASIG5V.n3931 0.9005
R48943 ASIG5V.n4135 ASIG5V.n3895 0.9005
R48944 ASIG5V.n4089 ASIG5V.n3933 0.9005
R48945 ASIG5V.n4139 ASIG5V.n3894 0.9005
R48946 ASIG5V.n4140 ASIG5V.n3935 0.9005
R48947 ASIG5V.n4141 ASIG5V.n3893 0.9005
R48948 ASIG5V.n4087 ASIG5V.n3937 0.9005
R48949 ASIG5V.n4145 ASIG5V.n3892 0.9005
R48950 ASIG5V.n4146 ASIG5V.n3939 0.9005
R48951 ASIG5V.n4147 ASIG5V.n3891 0.9005
R48952 ASIG5V.n4085 ASIG5V.n3941 0.9005
R48953 ASIG5V.n4151 ASIG5V.n3890 0.9005
R48954 ASIG5V.n4152 ASIG5V.n3943 0.9005
R48955 ASIG5V.n4153 ASIG5V.n3889 0.9005
R48956 ASIG5V.n4083 ASIG5V.n3945 0.9005
R48957 ASIG5V.n4157 ASIG5V.n3888 0.9005
R48958 ASIG5V.n4158 ASIG5V.n3947 0.9005
R48959 ASIG5V.n4159 ASIG5V.n3887 0.9005
R48960 ASIG5V.n4081 ASIG5V.n3949 0.9005
R48961 ASIG5V.n4163 ASIG5V.n3886 0.9005
R48962 ASIG5V.n4164 ASIG5V.n3951 0.9005
R48963 ASIG5V.n4165 ASIG5V.n3885 0.9005
R48964 ASIG5V.n4079 ASIG5V.n3953 0.9005
R48965 ASIG5V.n4169 ASIG5V.n3884 0.9005
R48966 ASIG5V.n4170 ASIG5V.n3955 0.9005
R48967 ASIG5V.n4171 ASIG5V.n3883 0.9005
R48968 ASIG5V.n4077 ASIG5V.n3957 0.9005
R48969 ASIG5V.n4175 ASIG5V.n3882 0.9005
R48970 ASIG5V.n4176 ASIG5V.n3959 0.9005
R48971 ASIG5V.n4177 ASIG5V.n3881 0.9005
R48972 ASIG5V.n4075 ASIG5V.n3961 0.9005
R48973 ASIG5V.n4181 ASIG5V.n3880 0.9005
R48974 ASIG5V.n4182 ASIG5V.n3963 0.9005
R48975 ASIG5V.n4183 ASIG5V.n3879 0.9005
R48976 ASIG5V.n4073 ASIG5V.n3965 0.9005
R48977 ASIG5V.n4187 ASIG5V.n3878 0.9005
R48978 ASIG5V.n4188 ASIG5V.n3967 0.9005
R48979 ASIG5V.n4189 ASIG5V.n3877 0.9005
R48980 ASIG5V.n4071 ASIG5V.n3969 0.9005
R48981 ASIG5V.n4193 ASIG5V.n3876 0.9005
R48982 ASIG5V.n4194 ASIG5V.n3971 0.9005
R48983 ASIG5V.n4195 ASIG5V.n3875 0.9005
R48984 ASIG5V.n4069 ASIG5V.n3973 0.9005
R48985 ASIG5V.n4199 ASIG5V.n3874 0.9005
R48986 ASIG5V.n4200 ASIG5V.n3975 0.9005
R48987 ASIG5V.n4201 ASIG5V.n3873 0.9005
R48988 ASIG5V.n4067 ASIG5V.n3977 0.9005
R48989 ASIG5V.n4205 ASIG5V.n3872 0.9005
R48990 ASIG5V.n4206 ASIG5V.n3979 0.9005
R48991 ASIG5V.n4207 ASIG5V.n3871 0.9005
R48992 ASIG5V.n4065 ASIG5V.n3981 0.9005
R48993 ASIG5V.n4211 ASIG5V.n3870 0.9005
R48994 ASIG5V.n4212 ASIG5V.n3983 0.9005
R48995 ASIG5V.n4213 ASIG5V.n3869 0.9005
R48996 ASIG5V.n4063 ASIG5V.n3985 0.9005
R48997 ASIG5V.n4217 ASIG5V.n3868 0.9005
R48998 ASIG5V.n4218 ASIG5V.n3987 0.9005
R48999 ASIG5V.n4219 ASIG5V.n3867 0.9005
R49000 ASIG5V.n4061 ASIG5V.n3989 0.9005
R49001 ASIG5V.n4223 ASIG5V.n3866 0.9005
R49002 ASIG5V.n4224 ASIG5V.n3991 0.9005
R49003 ASIG5V.n4225 ASIG5V.n3865 0.9005
R49004 ASIG5V.n4059 ASIG5V.n3993 0.9005
R49005 ASIG5V.n4229 ASIG5V.n3864 0.9005
R49006 ASIG5V.n4230 ASIG5V.n3995 0.9005
R49007 ASIG5V.n4231 ASIG5V.n3863 0.9005
R49008 ASIG5V.n4057 ASIG5V.n3997 0.9005
R49009 ASIG5V.n4235 ASIG5V.n3862 0.9005
R49010 ASIG5V.n4236 ASIG5V.n3999 0.9005
R49011 ASIG5V.n4237 ASIG5V.n3861 0.9005
R49012 ASIG5V.n4055 ASIG5V.n4001 0.9005
R49013 ASIG5V.n4241 ASIG5V.n3860 0.9005
R49014 ASIG5V.n4242 ASIG5V.n4003 0.9005
R49015 ASIG5V.n4243 ASIG5V.n3859 0.9005
R49016 ASIG5V.n4254 ASIG5V.n4252 0.9005
R49017 ASIG5V.n10711 ASIG5V.n10710 0.757975
R49018 ASIG5V.n4259 ASIG5V.n3843 0.757975
R49019 ASIG5V.n10694 ASIG5V.n10693 0.7505
R49020 ASIG5V.n10715 ASIG5V.n10714 0.7505
R49021 ASIG5V.n10714 ASIG5V.n10713 0.7505
R49022 ASIG5V.n10700 ASIG5V.n10694 0.7505
R49023 ASIG5V.n10705 ASIG5V.n10698 0.7505
R49024 ASIG5V.n4263 ASIG5V.n4262 0.7505
R49025 ASIG5V.n3845 ASIG5V.n3844 0.7505
R49026 ASIG5V.n4257 ASIG5V.n3845 0.7505
R49027 ASIG5V.n4262 ASIG5V.n4261 0.7505
R49028 ASIG5V.n3853 ASIG5V.n3852 0.7505
R49029 ASIG5V.n8124 ASIG5V.n7459 0.478669
R49030 ASIG5V.n8130 ASIG5V.n8129 0.478669
R49031 ASIG5V.n7607 ASIG5V.n7294 0.478669
R49032 ASIG5V.n7593 ASIG5V.n7592 0.478669
R49033 ASIG5V.n7677 ASIG5V.n7675 0.478669
R49034 ASIG5V.n9789 ASIG5V.n9788 0.478669
R49035 ASIG5V.n9925 ASIG5V.n9924 0.478669
R49036 ASIG5V.n8029 ASIG5V.n8028 0.478669
R49037 ASIG5V.n10710 ASIG5V.n10709 0.383312
R49038 ASIG5V.n4264 ASIG5V.n3843 0.383312
R49039 ASIG5V.n11798 ASIG5V.n1841 0.296012
R49040 ASIG5V.n7341 ASIG5V.n7340 0.296012
R49041 ASIG5V.n12328 ASIG5V.n169 0.296012
R49042 ASIG5V.n8901 ASIG5V.n8167 0.296012
R49043 ASIG5V.n7712 ASIG5V.n6416 0.296012
R49044 ASIG5V.n9752 ASIG5V.n9748 0.296012
R49045 ASIG5V.n9953 ASIG5V.n9952 0.296012
R49046 ASIG5V.n7983 ASIG5V.n7982 0.296012
R49047 ASIG5V.n9891 ASIG5V.n3083 0.161366
R49048 ASIG5V.n8109 ASIG5V.n8107 0.161366
R49049 ASIG5V.n8117 ASIG5V.n8116 0.161366
R49050 ASIG5V.n7449 ASIG5V.n7448 0.161366
R49051 ASIG5V.n7438 ASIG5V.n7437 0.161366
R49052 ASIG5V.n7427 ASIG5V.n7426 0.161366
R49053 ASIG5V.n7475 ASIG5V.n3088 0.161366
R49054 ASIG5V.n7633 ASIG5V.n7476 0.161366
R49055 ASIG5V.n7624 ASIG5V.n7315 0.161366
R49056 ASIG5V.n8137 ASIG5V.n7303 0.161366
R49057 ASIG5V.n7378 ASIG5V.n7377 0.161366
R49058 ASIG5V.n7385 ASIG5V.n7338 0.161366
R49059 ASIG5V.n7482 ASIG5V.n3095 0.161366
R49060 ASIG5V.n7636 ASIG5V.n7483 0.161366
R49061 ASIG5V.n7643 ASIG5V.n7617 0.161366
R49062 ASIG5V.n8143 ASIG5V.n8142 0.161366
R49063 ASIG5V.n8150 ASIG5V.n7283 0.161366
R49064 ASIG5V.n7392 ASIG5V.n7391 0.161366
R49065 ASIG5V.n7489 ASIG5V.n3102 0.161366
R49066 ASIG5V.n7645 ASIG5V.n7490 0.161366
R49067 ASIG5V.n7652 ASIG5V.n7566 0.161366
R49068 ASIG5V.n7590 ASIG5V.n7274 0.161366
R49069 ASIG5V.n8156 ASIG5V.n8155 0.161366
R49070 ASIG5V.n8162 ASIG5V.n8161 0.161366
R49071 ASIG5V.n7496 ASIG5V.n3109 0.161366
R49072 ASIG5V.n7655 ASIG5V.n7497 0.161366
R49073 ASIG5V.n7666 ASIG5V.n7664 0.161366
R49074 ASIG5V.n7688 ASIG5V.n7686 0.161366
R49075 ASIG5V.n7698 ASIG5V.n7697 0.161366
R49076 ASIG5V.n7705 ASIG5V.n7704 0.161366
R49077 ASIG5V.n9825 ASIG5V.n9824 0.161366
R49078 ASIG5V.n9813 ASIG5V.n9812 0.161366
R49079 ASIG5V.n9801 ASIG5V.n9800 0.161366
R49080 ASIG5V.n9777 ASIG5V.n9776 0.161366
R49081 ASIG5V.n9765 ASIG5V.n9764 0.161366
R49082 ASIG5V.n9762 ASIG5V.n9754 0.161366
R49083 ASIG5V.n9907 ASIG5V.n9906 0.161366
R49084 ASIG5V.n9913 ASIG5V.n9912 0.161366
R49085 ASIG5V.n9919 ASIG5V.n9918 0.161366
R49086 ASIG5V.n9931 ASIG5V.n9930 0.161366
R49087 ASIG5V.n9937 ASIG5V.n9936 0.161366
R49088 ASIG5V.n9943 ASIG5V.n9942 0.161366
R49089 ASIG5V.n7503 ASIG5V.n3116 0.161366
R49090 ASIG5V.n8051 ASIG5V.n8050 0.161366
R49091 ASIG5V.n8040 ASIG5V.n8039 0.161366
R49092 ASIG5V.n8018 ASIG5V.n8017 0.161366
R49093 ASIG5V.n8007 ASIG5V.n8006 0.161366
R49094 ASIG5V.n7996 ASIG5V.n7995 0.161366
R49095 ASIG5V.n9843 ASIG5V.n9837 0.1151
R49096 ASIG5V.n9852 ASIG5V.n9846 0.1151
R49097 ASIG5V.n9861 ASIG5V.n9855 0.1151
R49098 ASIG5V.n9879 ASIG5V.n9873 0.1151
R49099 ASIG5V.n9885 ASIG5V.n9882 0.1151
R49100 ASIG5V.n9905 ASIG5V.n9892 0.1151
R49101 ASIG5V.n9823 ASIG5V.n3127 0.1151
R49102 ASIG5V.n8068 ASIG5V.n8062 0.1151
R49103 ASIG5V.n8077 ASIG5V.n8071 0.1151
R49104 ASIG5V.n8095 ASIG5V.n8089 0.1151
R49105 ASIG5V.n8100 ASIG5V.n8098 0.1151
R49106 ASIG5V.n9911 ASIG5V.n3067 0.1151
R49107 ASIG5V.n9811 ASIG5V.n3132 0.1151
R49108 ASIG5V.n8049 ASIG5V.n7508 0.1151
R49109 ASIG5V.n7656 ASIG5V.n7653 0.1151
R49110 ASIG5V.n7637 ASIG5V.n7635 0.1151
R49111 ASIG5V.n8115 ASIG5V.n7464 0.1151
R49112 ASIG5V.n9917 ASIG5V.n3056 0.1151
R49113 ASIG5V.n9799 ASIG5V.n3137 0.1151
R49114 ASIG5V.n8038 ASIG5V.n7513 0.1151
R49115 ASIG5V.n7667 ASIG5V.n7557 0.1151
R49116 ASIG5V.n8128 ASIG5V.n7310 0.1151
R49117 ASIG5V.n8126 ASIG5V.n8125 0.1151
R49118 ASIG5V.n9923 ASIG5V.n3045 0.1151
R49119 ASIG5V.n9787 ASIG5V.n3142 0.1151
R49120 ASIG5V.n8027 ASIG5V.n7518 0.1151
R49121 ASIG5V.n7678 ASIG5V.n7552 0.1151
R49122 ASIG5V.n8139 ASIG5V.n8138 0.1151
R49123 ASIG5V.n8131 ASIG5V.n7307 0.1151
R49124 ASIG5V.n9929 ASIG5V.n3034 0.1151
R49125 ASIG5V.n9775 ASIG5V.n3147 0.1151
R49126 ASIG5V.n8016 ASIG5V.n7523 0.1151
R49127 ASIG5V.n8154 ASIG5V.n7269 0.1151
R49128 ASIG5V.n8144 ASIG5V.n7287 0.1151
R49129 ASIG5V.n7369 ASIG5V.n7328 0.1151
R49130 ASIG5V.n9935 ASIG5V.n3023 0.1151
R49131 ASIG5V.n9763 ASIG5V.n3153 0.1151
R49132 ASIG5V.n8005 ASIG5V.n7528 0.1151
R49133 ASIG5V.n8160 ASIG5V.n7258 0.1151
R49134 ASIG5V.n7387 ASIG5V.n7386 0.1151
R49135 ASIG5V.n7379 ASIG5V.n7332 0.1151
R49136 ASIG5V.n9941 ASIG5V.n3012 0.1151
R49137 ASIG5V.n7991 ASIG5V.n7988 0.1151
R49138 ASIG5V.n7994 ASIG5V.n7713 0.1151
R49139 ASIG5V.n8166 ASIG5V.n7247 0.1151
R49140 ASIG5V.n7410 ASIG5V.n7404 0.1151
R49141 ASIG5V.n7414 ASIG5V.n7413 0.1151
R49142 ASIG5V.n9945 ASIG5V.n3009 0.1151
R49143 ASIG5V ASIG5V.n9864 0.0881
R49144 ASIG5V.n9870 ASIG5V 0.0881
R49145 ASIG5V ASIG5V.n8080 0.0881
R49146 ASIG5V.n8086 ASIG5V 0.0881
R49147 ASIG5V.n7646 ASIG5V 0.0881
R49148 ASIG5V ASIG5V.n7644 0.0881
R49149 ASIG5V ASIG5V.n7604 0.0881
R49150 ASIG5V.n7615 ASIG5V 0.0881
R49151 ASIG5V.n7591 ASIG5V 0.0881
R49152 ASIG5V.n8141 ASIG5V 0.0881
R49153 ASIG5V.n8152 ASIG5V 0.0881
R49154 ASIG5V ASIG5V.n8151 0.0881
R49155 ASIG5V.n8157 ASIG5V 0.0881
R49156 ASIG5V.n7390 ASIG5V 0.0881
R49157 ASIG5V.n8163 ASIG5V 0.0881
R49158 ASIG5V.n7401 ASIG5V 0.0881
R49159 ASIG5V.n10352 ASIG5V.n10119 0.0380882
R49160 ASIG5V.n10352 ASIG5V.n10351 0.0380882
R49161 ASIG5V.n10351 ASIG5V.n10350 0.0380882
R49162 ASIG5V.n10350 ASIG5V.n10120 0.0380882
R49163 ASIG5V.n10343 ASIG5V.n10120 0.0380882
R49164 ASIG5V.n10343 ASIG5V.n10342 0.0380882
R49165 ASIG5V.n10342 ASIG5V.n10341 0.0380882
R49166 ASIG5V.n10341 ASIG5V.n10123 0.0380882
R49167 ASIG5V.n10334 ASIG5V.n10123 0.0380882
R49168 ASIG5V.n10334 ASIG5V.n10333 0.0380882
R49169 ASIG5V.n10333 ASIG5V.n10332 0.0380882
R49170 ASIG5V.n10332 ASIG5V.n10126 0.0380882
R49171 ASIG5V.n10325 ASIG5V.n10126 0.0380882
R49172 ASIG5V.n10325 ASIG5V.n10324 0.0380882
R49173 ASIG5V.n10324 ASIG5V.n10323 0.0380882
R49174 ASIG5V.n10323 ASIG5V.n10129 0.0380882
R49175 ASIG5V.n10316 ASIG5V.n10129 0.0380882
R49176 ASIG5V.n10316 ASIG5V.n10315 0.0380882
R49177 ASIG5V.n10315 ASIG5V.n10314 0.0380882
R49178 ASIG5V.n10314 ASIG5V.n10132 0.0380882
R49179 ASIG5V.n10307 ASIG5V.n10132 0.0380882
R49180 ASIG5V.n10307 ASIG5V.n10306 0.0380882
R49181 ASIG5V.n10306 ASIG5V.n10305 0.0380882
R49182 ASIG5V.n10305 ASIG5V.n10135 0.0380882
R49183 ASIG5V.n10298 ASIG5V.n10135 0.0380882
R49184 ASIG5V.n10298 ASIG5V.n10297 0.0380882
R49185 ASIG5V.n10297 ASIG5V.n10296 0.0380882
R49186 ASIG5V.n10296 ASIG5V.n10138 0.0380882
R49187 ASIG5V.n10289 ASIG5V.n10138 0.0380882
R49188 ASIG5V.n10289 ASIG5V.n10288 0.0380882
R49189 ASIG5V.n10288 ASIG5V.n10287 0.0380882
R49190 ASIG5V.n10287 ASIG5V.n10141 0.0380882
R49191 ASIG5V.n10280 ASIG5V.n10141 0.0380882
R49192 ASIG5V.n10280 ASIG5V.n10279 0.0380882
R49193 ASIG5V.n10279 ASIG5V.n10278 0.0380882
R49194 ASIG5V.n10278 ASIG5V.n10144 0.0380882
R49195 ASIG5V.n10271 ASIG5V.n10144 0.0380882
R49196 ASIG5V.n10271 ASIG5V.n10270 0.0380882
R49197 ASIG5V.n10270 ASIG5V.n10269 0.0380882
R49198 ASIG5V.n10269 ASIG5V.n10147 0.0380882
R49199 ASIG5V.n10262 ASIG5V.n10147 0.0380882
R49200 ASIG5V.n10262 ASIG5V.n10261 0.0380882
R49201 ASIG5V.n10261 ASIG5V.n10260 0.0380882
R49202 ASIG5V.n10260 ASIG5V.n10150 0.0380882
R49203 ASIG5V.n10253 ASIG5V.n10150 0.0380882
R49204 ASIG5V.n10253 ASIG5V.n10252 0.0380882
R49205 ASIG5V.n10252 ASIG5V.n10251 0.0380882
R49206 ASIG5V.n10251 ASIG5V.n10153 0.0380882
R49207 ASIG5V.n10244 ASIG5V.n10153 0.0380882
R49208 ASIG5V.n10244 ASIG5V.n10243 0.0380882
R49209 ASIG5V.n10243 ASIG5V.n10242 0.0380882
R49210 ASIG5V.n10242 ASIG5V.n10156 0.0380882
R49211 ASIG5V.n10235 ASIG5V.n10156 0.0380882
R49212 ASIG5V.n10235 ASIG5V.n10234 0.0380882
R49213 ASIG5V.n10234 ASIG5V.n10233 0.0380882
R49214 ASIG5V.n10233 ASIG5V.n10159 0.0380882
R49215 ASIG5V.n10226 ASIG5V.n10159 0.0380882
R49216 ASIG5V.n10226 ASIG5V.n10225 0.0380882
R49217 ASIG5V.n10225 ASIG5V.n10224 0.0380882
R49218 ASIG5V.n10224 ASIG5V.n10162 0.0380882
R49219 ASIG5V.n10217 ASIG5V.n10162 0.0380882
R49220 ASIG5V.n10217 ASIG5V.n10216 0.0380882
R49221 ASIG5V.n10216 ASIG5V.n10215 0.0380882
R49222 ASIG5V.n10215 ASIG5V.n10165 0.0380882
R49223 ASIG5V.n10208 ASIG5V.n10165 0.0380882
R49224 ASIG5V.n10208 ASIG5V.n10207 0.0380882
R49225 ASIG5V.n10207 ASIG5V.n10206 0.0380882
R49226 ASIG5V.n10206 ASIG5V.n10168 0.0380882
R49227 ASIG5V.n10199 ASIG5V.n10168 0.0380882
R49228 ASIG5V.n10199 ASIG5V.n10198 0.0380882
R49229 ASIG5V.n10198 ASIG5V.n10197 0.0380882
R49230 ASIG5V.n10197 ASIG5V.n10171 0.0380882
R49231 ASIG5V.n10190 ASIG5V.n10171 0.0380882
R49232 ASIG5V.n10190 ASIG5V.n10189 0.0380882
R49233 ASIG5V.n10189 ASIG5V.n10188 0.0380882
R49234 ASIG5V.n10188 ASIG5V.n10174 0.0380882
R49235 ASIG5V.n10181 ASIG5V.n10174 0.0380882
R49236 ASIG5V.n10181 ASIG5V.n10180 0.0380882
R49237 ASIG5V.n10180 ASIG5V.n10179 0.0380882
R49238 ASIG5V.n10179 ASIG5V.n10073 0.0380882
R49239 ASIG5V.n10360 ASIG5V.n10073 0.0380882
R49240 ASIG5V.n10361 ASIG5V.n10360 0.0380882
R49241 ASIG5V.n10362 ASIG5V.n10361 0.0380882
R49242 ASIG5V.n3616 ASIG5V.n3282 0.0380882
R49243 ASIG5V.n3608 ASIG5V.n3282 0.0380882
R49244 ASIG5V.n3608 ASIG5V.n3607 0.0380882
R49245 ASIG5V.n3607 ASIG5V.n3606 0.0380882
R49246 ASIG5V.n3606 ASIG5V.n3286 0.0380882
R49247 ASIG5V.n3598 ASIG5V.n3286 0.0380882
R49248 ASIG5V.n3598 ASIG5V.n3597 0.0380882
R49249 ASIG5V.n3597 ASIG5V.n3596 0.0380882
R49250 ASIG5V.n3596 ASIG5V.n3292 0.0380882
R49251 ASIG5V.n3588 ASIG5V.n3292 0.0380882
R49252 ASIG5V.n3588 ASIG5V.n3587 0.0380882
R49253 ASIG5V.n3587 ASIG5V.n3586 0.0380882
R49254 ASIG5V.n3586 ASIG5V.n3298 0.0380882
R49255 ASIG5V.n3578 ASIG5V.n3298 0.0380882
R49256 ASIG5V.n3578 ASIG5V.n3577 0.0380882
R49257 ASIG5V.n3577 ASIG5V.n3576 0.0380882
R49258 ASIG5V.n3576 ASIG5V.n3304 0.0380882
R49259 ASIG5V.n3568 ASIG5V.n3304 0.0380882
R49260 ASIG5V.n3568 ASIG5V.n3567 0.0380882
R49261 ASIG5V.n3567 ASIG5V.n3566 0.0380882
R49262 ASIG5V.n3566 ASIG5V.n3310 0.0380882
R49263 ASIG5V.n3558 ASIG5V.n3310 0.0380882
R49264 ASIG5V.n3558 ASIG5V.n3557 0.0380882
R49265 ASIG5V.n3557 ASIG5V.n3556 0.0380882
R49266 ASIG5V.n3556 ASIG5V.n3316 0.0380882
R49267 ASIG5V.n3548 ASIG5V.n3316 0.0380882
R49268 ASIG5V.n3548 ASIG5V.n3547 0.0380882
R49269 ASIG5V.n3547 ASIG5V.n3546 0.0380882
R49270 ASIG5V.n3546 ASIG5V.n3322 0.0380882
R49271 ASIG5V.n3538 ASIG5V.n3322 0.0380882
R49272 ASIG5V.n3538 ASIG5V.n3537 0.0380882
R49273 ASIG5V.n3537 ASIG5V.n3536 0.0380882
R49274 ASIG5V.n3536 ASIG5V.n3328 0.0380882
R49275 ASIG5V.n3528 ASIG5V.n3328 0.0380882
R49276 ASIG5V.n3528 ASIG5V.n3527 0.0380882
R49277 ASIG5V.n3527 ASIG5V.n3526 0.0380882
R49278 ASIG5V.n3526 ASIG5V.n3334 0.0380882
R49279 ASIG5V.n3518 ASIG5V.n3334 0.0380882
R49280 ASIG5V.n3518 ASIG5V.n3517 0.0380882
R49281 ASIG5V.n3517 ASIG5V.n3516 0.0380882
R49282 ASIG5V.n3516 ASIG5V.n3340 0.0380882
R49283 ASIG5V.n3508 ASIG5V.n3340 0.0380882
R49284 ASIG5V.n3508 ASIG5V.n3507 0.0380882
R49285 ASIG5V.n3507 ASIG5V.n3506 0.0380882
R49286 ASIG5V.n3506 ASIG5V.n3346 0.0380882
R49287 ASIG5V.n3498 ASIG5V.n3346 0.0380882
R49288 ASIG5V.n3498 ASIG5V.n3497 0.0380882
R49289 ASIG5V.n3497 ASIG5V.n3496 0.0380882
R49290 ASIG5V.n3496 ASIG5V.n3352 0.0380882
R49291 ASIG5V.n3488 ASIG5V.n3352 0.0380882
R49292 ASIG5V.n3488 ASIG5V.n3487 0.0380882
R49293 ASIG5V.n3487 ASIG5V.n3486 0.0380882
R49294 ASIG5V.n3486 ASIG5V.n3358 0.0380882
R49295 ASIG5V.n3478 ASIG5V.n3358 0.0380882
R49296 ASIG5V.n3478 ASIG5V.n3477 0.0380882
R49297 ASIG5V.n3477 ASIG5V.n3476 0.0380882
R49298 ASIG5V.n3476 ASIG5V.n3364 0.0380882
R49299 ASIG5V.n3468 ASIG5V.n3364 0.0380882
R49300 ASIG5V.n3468 ASIG5V.n3467 0.0380882
R49301 ASIG5V.n3467 ASIG5V.n3466 0.0380882
R49302 ASIG5V.n3466 ASIG5V.n3370 0.0380882
R49303 ASIG5V.n3458 ASIG5V.n3370 0.0380882
R49304 ASIG5V.n3458 ASIG5V.n3457 0.0380882
R49305 ASIG5V.n3457 ASIG5V.n3456 0.0380882
R49306 ASIG5V.n3456 ASIG5V.n3376 0.0380882
R49307 ASIG5V.n3448 ASIG5V.n3376 0.0380882
R49308 ASIG5V.n3448 ASIG5V.n3447 0.0380882
R49309 ASIG5V.n3447 ASIG5V.n3446 0.0380882
R49310 ASIG5V.n3446 ASIG5V.n3382 0.0380882
R49311 ASIG5V.n3438 ASIG5V.n3382 0.0380882
R49312 ASIG5V.n3438 ASIG5V.n3437 0.0380882
R49313 ASIG5V.n3437 ASIG5V.n3436 0.0380882
R49314 ASIG5V.n3436 ASIG5V.n3388 0.0380882
R49315 ASIG5V.n3428 ASIG5V.n3388 0.0380882
R49316 ASIG5V.n3428 ASIG5V.n3427 0.0380882
R49317 ASIG5V.n3427 ASIG5V.n3426 0.0380882
R49318 ASIG5V.n3426 ASIG5V.n3394 0.0380882
R49319 ASIG5V.n3418 ASIG5V.n3394 0.0380882
R49320 ASIG5V.n3418 ASIG5V.n3417 0.0380882
R49321 ASIG5V.n3417 ASIG5V.n3416 0.0380882
R49322 ASIG5V.n3416 ASIG5V.n3400 0.0380882
R49323 ASIG5V.n3408 ASIG5V.n3400 0.0380882
R49324 ASIG5V.n3408 ASIG5V.n3407 0.0380882
R49325 ASIG5V.n3615 ASIG5V.n3283 0.0380882
R49326 ASIG5V.n3609 ASIG5V.n3283 0.0380882
R49327 ASIG5V.n3609 ASIG5V.n3285 0.0380882
R49328 ASIG5V.n3605 ASIG5V.n3285 0.0380882
R49329 ASIG5V.n3605 ASIG5V.n3287 0.0380882
R49330 ASIG5V.n3599 ASIG5V.n3287 0.0380882
R49331 ASIG5V.n3599 ASIG5V.n3291 0.0380882
R49332 ASIG5V.n3595 ASIG5V.n3291 0.0380882
R49333 ASIG5V.n3595 ASIG5V.n3293 0.0380882
R49334 ASIG5V.n3589 ASIG5V.n3293 0.0380882
R49335 ASIG5V.n3589 ASIG5V.n3297 0.0380882
R49336 ASIG5V.n3585 ASIG5V.n3297 0.0380882
R49337 ASIG5V.n3585 ASIG5V.n3299 0.0380882
R49338 ASIG5V.n3579 ASIG5V.n3299 0.0380882
R49339 ASIG5V.n3579 ASIG5V.n3303 0.0380882
R49340 ASIG5V.n3575 ASIG5V.n3303 0.0380882
R49341 ASIG5V.n3575 ASIG5V.n3305 0.0380882
R49342 ASIG5V.n3569 ASIG5V.n3305 0.0380882
R49343 ASIG5V.n3569 ASIG5V.n3309 0.0380882
R49344 ASIG5V.n3565 ASIG5V.n3309 0.0380882
R49345 ASIG5V.n3565 ASIG5V.n3311 0.0380882
R49346 ASIG5V.n3559 ASIG5V.n3311 0.0380882
R49347 ASIG5V.n3559 ASIG5V.n3315 0.0380882
R49348 ASIG5V.n3555 ASIG5V.n3315 0.0380882
R49349 ASIG5V.n3555 ASIG5V.n3317 0.0380882
R49350 ASIG5V.n3549 ASIG5V.n3317 0.0380882
R49351 ASIG5V.n3549 ASIG5V.n3321 0.0380882
R49352 ASIG5V.n3545 ASIG5V.n3321 0.0380882
R49353 ASIG5V.n3545 ASIG5V.n3323 0.0380882
R49354 ASIG5V.n3539 ASIG5V.n3323 0.0380882
R49355 ASIG5V.n3539 ASIG5V.n3327 0.0380882
R49356 ASIG5V.n3535 ASIG5V.n3327 0.0380882
R49357 ASIG5V.n3535 ASIG5V.n3329 0.0380882
R49358 ASIG5V.n3529 ASIG5V.n3329 0.0380882
R49359 ASIG5V.n3529 ASIG5V.n3333 0.0380882
R49360 ASIG5V.n3525 ASIG5V.n3333 0.0380882
R49361 ASIG5V.n3525 ASIG5V.n3335 0.0380882
R49362 ASIG5V.n3519 ASIG5V.n3335 0.0380882
R49363 ASIG5V.n3519 ASIG5V.n3339 0.0380882
R49364 ASIG5V.n3515 ASIG5V.n3339 0.0380882
R49365 ASIG5V.n3515 ASIG5V.n3341 0.0380882
R49366 ASIG5V.n3509 ASIG5V.n3341 0.0380882
R49367 ASIG5V.n3509 ASIG5V.n3345 0.0380882
R49368 ASIG5V.n3505 ASIG5V.n3345 0.0380882
R49369 ASIG5V.n3505 ASIG5V.n3347 0.0380882
R49370 ASIG5V.n3499 ASIG5V.n3347 0.0380882
R49371 ASIG5V.n3499 ASIG5V.n3351 0.0380882
R49372 ASIG5V.n3495 ASIG5V.n3351 0.0380882
R49373 ASIG5V.n3495 ASIG5V.n3353 0.0380882
R49374 ASIG5V.n3489 ASIG5V.n3353 0.0380882
R49375 ASIG5V.n3489 ASIG5V.n3357 0.0380882
R49376 ASIG5V.n3485 ASIG5V.n3357 0.0380882
R49377 ASIG5V.n3485 ASIG5V.n3359 0.0380882
R49378 ASIG5V.n3479 ASIG5V.n3359 0.0380882
R49379 ASIG5V.n3479 ASIG5V.n3363 0.0380882
R49380 ASIG5V.n3475 ASIG5V.n3363 0.0380882
R49381 ASIG5V.n3475 ASIG5V.n3365 0.0380882
R49382 ASIG5V.n3469 ASIG5V.n3365 0.0380882
R49383 ASIG5V.n3469 ASIG5V.n3369 0.0380882
R49384 ASIG5V.n3465 ASIG5V.n3369 0.0380882
R49385 ASIG5V.n3465 ASIG5V.n3371 0.0380882
R49386 ASIG5V.n3459 ASIG5V.n3371 0.0380882
R49387 ASIG5V.n3459 ASIG5V.n3375 0.0380882
R49388 ASIG5V.n3455 ASIG5V.n3375 0.0380882
R49389 ASIG5V.n3455 ASIG5V.n3377 0.0380882
R49390 ASIG5V.n3449 ASIG5V.n3377 0.0380882
R49391 ASIG5V.n3449 ASIG5V.n3381 0.0380882
R49392 ASIG5V.n3445 ASIG5V.n3381 0.0380882
R49393 ASIG5V.n3445 ASIG5V.n3383 0.0380882
R49394 ASIG5V.n3439 ASIG5V.n3383 0.0380882
R49395 ASIG5V.n3439 ASIG5V.n3387 0.0380882
R49396 ASIG5V.n3435 ASIG5V.n3387 0.0380882
R49397 ASIG5V.n3435 ASIG5V.n3389 0.0380882
R49398 ASIG5V.n3429 ASIG5V.n3389 0.0380882
R49399 ASIG5V.n3429 ASIG5V.n3393 0.0380882
R49400 ASIG5V.n3425 ASIG5V.n3393 0.0380882
R49401 ASIG5V.n3425 ASIG5V.n3395 0.0380882
R49402 ASIG5V.n3419 ASIG5V.n3395 0.0380882
R49403 ASIG5V.n3419 ASIG5V.n3399 0.0380882
R49404 ASIG5V.n3415 ASIG5V.n3399 0.0380882
R49405 ASIG5V.n3415 ASIG5V.n3401 0.0380882
R49406 ASIG5V.n3409 ASIG5V.n3401 0.0380882
R49407 ASIG5V.n3409 ASIG5V.n3406 0.0380882
R49408 ASIG5V.n4817 ASIG5V.n4816 0.0380882
R49409 ASIG5V.n4818 ASIG5V.n4817 0.0380882
R49410 ASIG5V.n4818 ASIG5V.n3263 0.0380882
R49411 ASIG5V.n4828 ASIG5V.n3263 0.0380882
R49412 ASIG5V.n4829 ASIG5V.n4828 0.0380882
R49413 ASIG5V.n4830 ASIG5V.n4829 0.0380882
R49414 ASIG5V.n4830 ASIG5V.n3261 0.0380882
R49415 ASIG5V.n4840 ASIG5V.n3261 0.0380882
R49416 ASIG5V.n4841 ASIG5V.n4840 0.0380882
R49417 ASIG5V.n4842 ASIG5V.n4841 0.0380882
R49418 ASIG5V.n4842 ASIG5V.n3259 0.0380882
R49419 ASIG5V.n4852 ASIG5V.n3259 0.0380882
R49420 ASIG5V.n4853 ASIG5V.n4852 0.0380882
R49421 ASIG5V.n4854 ASIG5V.n4853 0.0380882
R49422 ASIG5V.n4854 ASIG5V.n3257 0.0380882
R49423 ASIG5V.n4864 ASIG5V.n3257 0.0380882
R49424 ASIG5V.n4865 ASIG5V.n4864 0.0380882
R49425 ASIG5V.n4866 ASIG5V.n4865 0.0380882
R49426 ASIG5V.n4866 ASIG5V.n3255 0.0380882
R49427 ASIG5V.n4876 ASIG5V.n3255 0.0380882
R49428 ASIG5V.n4877 ASIG5V.n4876 0.0380882
R49429 ASIG5V.n4878 ASIG5V.n4877 0.0380882
R49430 ASIG5V.n4878 ASIG5V.n3253 0.0380882
R49431 ASIG5V.n4888 ASIG5V.n3253 0.0380882
R49432 ASIG5V.n4889 ASIG5V.n4888 0.0380882
R49433 ASIG5V.n4890 ASIG5V.n4889 0.0380882
R49434 ASIG5V.n4890 ASIG5V.n3251 0.0380882
R49435 ASIG5V.n4900 ASIG5V.n3251 0.0380882
R49436 ASIG5V.n4901 ASIG5V.n4900 0.0380882
R49437 ASIG5V.n4902 ASIG5V.n4901 0.0380882
R49438 ASIG5V.n4902 ASIG5V.n3249 0.0380882
R49439 ASIG5V.n4912 ASIG5V.n3249 0.0380882
R49440 ASIG5V.n4913 ASIG5V.n4912 0.0380882
R49441 ASIG5V.n4914 ASIG5V.n4913 0.0380882
R49442 ASIG5V.n4914 ASIG5V.n3247 0.0380882
R49443 ASIG5V.n4924 ASIG5V.n3247 0.0380882
R49444 ASIG5V.n4925 ASIG5V.n4924 0.0380882
R49445 ASIG5V.n4926 ASIG5V.n4925 0.0380882
R49446 ASIG5V.n4926 ASIG5V.n3245 0.0380882
R49447 ASIG5V.n4936 ASIG5V.n3245 0.0380882
R49448 ASIG5V.n4937 ASIG5V.n4936 0.0380882
R49449 ASIG5V.n4938 ASIG5V.n4937 0.0380882
R49450 ASIG5V.n4938 ASIG5V.n3243 0.0380882
R49451 ASIG5V.n4948 ASIG5V.n3243 0.0380882
R49452 ASIG5V.n4949 ASIG5V.n4948 0.0380882
R49453 ASIG5V.n4950 ASIG5V.n4949 0.0380882
R49454 ASIG5V.n4950 ASIG5V.n3241 0.0380882
R49455 ASIG5V.n4960 ASIG5V.n3241 0.0380882
R49456 ASIG5V.n4961 ASIG5V.n4960 0.0380882
R49457 ASIG5V.n4962 ASIG5V.n4961 0.0380882
R49458 ASIG5V.n4962 ASIG5V.n3239 0.0380882
R49459 ASIG5V.n4972 ASIG5V.n3239 0.0380882
R49460 ASIG5V.n4973 ASIG5V.n4972 0.0380882
R49461 ASIG5V.n4974 ASIG5V.n4973 0.0380882
R49462 ASIG5V.n4974 ASIG5V.n3237 0.0380882
R49463 ASIG5V.n4984 ASIG5V.n3237 0.0380882
R49464 ASIG5V.n4985 ASIG5V.n4984 0.0380882
R49465 ASIG5V.n4986 ASIG5V.n4985 0.0380882
R49466 ASIG5V.n4986 ASIG5V.n3235 0.0380882
R49467 ASIG5V.n4996 ASIG5V.n3235 0.0380882
R49468 ASIG5V.n4997 ASIG5V.n4996 0.0380882
R49469 ASIG5V.n4998 ASIG5V.n4997 0.0380882
R49470 ASIG5V.n4998 ASIG5V.n3233 0.0380882
R49471 ASIG5V.n5008 ASIG5V.n3233 0.0380882
R49472 ASIG5V.n5009 ASIG5V.n5008 0.0380882
R49473 ASIG5V.n5010 ASIG5V.n5009 0.0380882
R49474 ASIG5V.n5010 ASIG5V.n3231 0.0380882
R49475 ASIG5V.n5020 ASIG5V.n3231 0.0380882
R49476 ASIG5V.n5021 ASIG5V.n5020 0.0380882
R49477 ASIG5V.n5022 ASIG5V.n5021 0.0380882
R49478 ASIG5V.n5022 ASIG5V.n3229 0.0380882
R49479 ASIG5V.n5032 ASIG5V.n3229 0.0380882
R49480 ASIG5V.n5033 ASIG5V.n5032 0.0380882
R49481 ASIG5V.n5034 ASIG5V.n5033 0.0380882
R49482 ASIG5V.n5034 ASIG5V.n3227 0.0380882
R49483 ASIG5V.n5044 ASIG5V.n3227 0.0380882
R49484 ASIG5V.n5045 ASIG5V.n5044 0.0380882
R49485 ASIG5V.n5046 ASIG5V.n5045 0.0380882
R49486 ASIG5V.n5046 ASIG5V.n3225 0.0380882
R49487 ASIG5V.n5056 ASIG5V.n3225 0.0380882
R49488 ASIG5V.n5057 ASIG5V.n5056 0.0380882
R49489 ASIG5V.n5059 ASIG5V.n5057 0.0380882
R49490 ASIG5V.n5059 ASIG5V.n5058 0.0380882
R49491 ASIG5V.n4815 ASIG5V.n3266 0.0380882
R49492 ASIG5V.n4819 ASIG5V.n3266 0.0380882
R49493 ASIG5V.n4823 ASIG5V.n4819 0.0380882
R49494 ASIG5V.n4827 ASIG5V.n4823 0.0380882
R49495 ASIG5V.n4827 ASIG5V.n3262 0.0380882
R49496 ASIG5V.n4831 ASIG5V.n3262 0.0380882
R49497 ASIG5V.n4835 ASIG5V.n4831 0.0380882
R49498 ASIG5V.n4839 ASIG5V.n4835 0.0380882
R49499 ASIG5V.n4839 ASIG5V.n3260 0.0380882
R49500 ASIG5V.n4843 ASIG5V.n3260 0.0380882
R49501 ASIG5V.n4847 ASIG5V.n4843 0.0380882
R49502 ASIG5V.n4851 ASIG5V.n4847 0.0380882
R49503 ASIG5V.n4851 ASIG5V.n3258 0.0380882
R49504 ASIG5V.n4855 ASIG5V.n3258 0.0380882
R49505 ASIG5V.n4859 ASIG5V.n4855 0.0380882
R49506 ASIG5V.n4863 ASIG5V.n4859 0.0380882
R49507 ASIG5V.n4863 ASIG5V.n3256 0.0380882
R49508 ASIG5V.n4867 ASIG5V.n3256 0.0380882
R49509 ASIG5V.n4871 ASIG5V.n4867 0.0380882
R49510 ASIG5V.n4875 ASIG5V.n4871 0.0380882
R49511 ASIG5V.n4875 ASIG5V.n3254 0.0380882
R49512 ASIG5V.n4879 ASIG5V.n3254 0.0380882
R49513 ASIG5V.n4883 ASIG5V.n4879 0.0380882
R49514 ASIG5V.n4887 ASIG5V.n4883 0.0380882
R49515 ASIG5V.n4887 ASIG5V.n3252 0.0380882
R49516 ASIG5V.n4891 ASIG5V.n3252 0.0380882
R49517 ASIG5V.n4895 ASIG5V.n4891 0.0380882
R49518 ASIG5V.n4899 ASIG5V.n4895 0.0380882
R49519 ASIG5V.n4899 ASIG5V.n3250 0.0380882
R49520 ASIG5V.n4903 ASIG5V.n3250 0.0380882
R49521 ASIG5V.n4907 ASIG5V.n4903 0.0380882
R49522 ASIG5V.n4911 ASIG5V.n4907 0.0380882
R49523 ASIG5V.n4911 ASIG5V.n3248 0.0380882
R49524 ASIG5V.n4915 ASIG5V.n3248 0.0380882
R49525 ASIG5V.n4919 ASIG5V.n4915 0.0380882
R49526 ASIG5V.n4923 ASIG5V.n4919 0.0380882
R49527 ASIG5V.n4923 ASIG5V.n3246 0.0380882
R49528 ASIG5V.n4927 ASIG5V.n3246 0.0380882
R49529 ASIG5V.n4931 ASIG5V.n4927 0.0380882
R49530 ASIG5V.n4935 ASIG5V.n4931 0.0380882
R49531 ASIG5V.n4935 ASIG5V.n3244 0.0380882
R49532 ASIG5V.n4939 ASIG5V.n3244 0.0380882
R49533 ASIG5V.n4943 ASIG5V.n4939 0.0380882
R49534 ASIG5V.n4947 ASIG5V.n4943 0.0380882
R49535 ASIG5V.n4947 ASIG5V.n3242 0.0380882
R49536 ASIG5V.n4951 ASIG5V.n3242 0.0380882
R49537 ASIG5V.n4955 ASIG5V.n4951 0.0380882
R49538 ASIG5V.n4959 ASIG5V.n4955 0.0380882
R49539 ASIG5V.n4959 ASIG5V.n3240 0.0380882
R49540 ASIG5V.n4963 ASIG5V.n3240 0.0380882
R49541 ASIG5V.n4967 ASIG5V.n4963 0.0380882
R49542 ASIG5V.n4971 ASIG5V.n4967 0.0380882
R49543 ASIG5V.n4971 ASIG5V.n3238 0.0380882
R49544 ASIG5V.n4975 ASIG5V.n3238 0.0380882
R49545 ASIG5V.n4979 ASIG5V.n4975 0.0380882
R49546 ASIG5V.n4983 ASIG5V.n4979 0.0380882
R49547 ASIG5V.n4983 ASIG5V.n3236 0.0380882
R49548 ASIG5V.n4987 ASIG5V.n3236 0.0380882
R49549 ASIG5V.n4991 ASIG5V.n4987 0.0380882
R49550 ASIG5V.n4995 ASIG5V.n4991 0.0380882
R49551 ASIG5V.n4995 ASIG5V.n3234 0.0380882
R49552 ASIG5V.n4999 ASIG5V.n3234 0.0380882
R49553 ASIG5V.n5003 ASIG5V.n4999 0.0380882
R49554 ASIG5V.n5007 ASIG5V.n5003 0.0380882
R49555 ASIG5V.n5007 ASIG5V.n3232 0.0380882
R49556 ASIG5V.n5011 ASIG5V.n3232 0.0380882
R49557 ASIG5V.n5015 ASIG5V.n5011 0.0380882
R49558 ASIG5V.n5019 ASIG5V.n5015 0.0380882
R49559 ASIG5V.n5019 ASIG5V.n3230 0.0380882
R49560 ASIG5V.n5023 ASIG5V.n3230 0.0380882
R49561 ASIG5V.n5027 ASIG5V.n5023 0.0380882
R49562 ASIG5V.n5031 ASIG5V.n5027 0.0380882
R49563 ASIG5V.n5031 ASIG5V.n3228 0.0380882
R49564 ASIG5V.n5035 ASIG5V.n3228 0.0380882
R49565 ASIG5V.n5039 ASIG5V.n5035 0.0380882
R49566 ASIG5V.n5043 ASIG5V.n5039 0.0380882
R49567 ASIG5V.n5043 ASIG5V.n3226 0.0380882
R49568 ASIG5V.n5047 ASIG5V.n3226 0.0380882
R49569 ASIG5V.n5051 ASIG5V.n5047 0.0380882
R49570 ASIG5V.n5055 ASIG5V.n5051 0.0380882
R49571 ASIG5V.n5055 ASIG5V.n3224 0.0380882
R49572 ASIG5V.n5060 ASIG5V.n3224 0.0380882
R49573 ASIG5V.n5060 ASIG5V.n3222 0.0380882
R49574 ASIG5V.n9488 ASIG5V.n9487 0.0380882
R49575 ASIG5V.n9489 ASIG5V.n9488 0.0380882
R49576 ASIG5V.n9489 ASIG5V.n9482 0.0380882
R49577 ASIG5V.n9499 ASIG5V.n9482 0.0380882
R49578 ASIG5V.n9500 ASIG5V.n9499 0.0380882
R49579 ASIG5V.n9501 ASIG5V.n9500 0.0380882
R49580 ASIG5V.n9501 ASIG5V.n9480 0.0380882
R49581 ASIG5V.n9511 ASIG5V.n9480 0.0380882
R49582 ASIG5V.n9512 ASIG5V.n9511 0.0380882
R49583 ASIG5V.n9513 ASIG5V.n9512 0.0380882
R49584 ASIG5V.n9513 ASIG5V.n9478 0.0380882
R49585 ASIG5V.n9523 ASIG5V.n9478 0.0380882
R49586 ASIG5V.n9524 ASIG5V.n9523 0.0380882
R49587 ASIG5V.n9525 ASIG5V.n9524 0.0380882
R49588 ASIG5V.n9525 ASIG5V.n9476 0.0380882
R49589 ASIG5V.n9535 ASIG5V.n9476 0.0380882
R49590 ASIG5V.n9536 ASIG5V.n9535 0.0380882
R49591 ASIG5V.n9537 ASIG5V.n9536 0.0380882
R49592 ASIG5V.n9537 ASIG5V.n9474 0.0380882
R49593 ASIG5V.n9547 ASIG5V.n9474 0.0380882
R49594 ASIG5V.n9548 ASIG5V.n9547 0.0380882
R49595 ASIG5V.n9549 ASIG5V.n9548 0.0380882
R49596 ASIG5V.n9549 ASIG5V.n9472 0.0380882
R49597 ASIG5V.n9559 ASIG5V.n9472 0.0380882
R49598 ASIG5V.n9560 ASIG5V.n9559 0.0380882
R49599 ASIG5V.n9561 ASIG5V.n9560 0.0380882
R49600 ASIG5V.n9561 ASIG5V.n9470 0.0380882
R49601 ASIG5V.n9571 ASIG5V.n9470 0.0380882
R49602 ASIG5V.n9572 ASIG5V.n9571 0.0380882
R49603 ASIG5V.n9573 ASIG5V.n9572 0.0380882
R49604 ASIG5V.n9573 ASIG5V.n9468 0.0380882
R49605 ASIG5V.n9583 ASIG5V.n9468 0.0380882
R49606 ASIG5V.n9584 ASIG5V.n9583 0.0380882
R49607 ASIG5V.n9585 ASIG5V.n9584 0.0380882
R49608 ASIG5V.n9585 ASIG5V.n9466 0.0380882
R49609 ASIG5V.n9595 ASIG5V.n9466 0.0380882
R49610 ASIG5V.n9596 ASIG5V.n9595 0.0380882
R49611 ASIG5V.n9597 ASIG5V.n9596 0.0380882
R49612 ASIG5V.n9597 ASIG5V.n9464 0.0380882
R49613 ASIG5V.n9607 ASIG5V.n9464 0.0380882
R49614 ASIG5V.n9608 ASIG5V.n9607 0.0380882
R49615 ASIG5V.n9609 ASIG5V.n9608 0.0380882
R49616 ASIG5V.n9609 ASIG5V.n9462 0.0380882
R49617 ASIG5V.n9619 ASIG5V.n9462 0.0380882
R49618 ASIG5V.n9620 ASIG5V.n9619 0.0380882
R49619 ASIG5V.n9621 ASIG5V.n9620 0.0380882
R49620 ASIG5V.n9621 ASIG5V.n9460 0.0380882
R49621 ASIG5V.n9631 ASIG5V.n9460 0.0380882
R49622 ASIG5V.n9632 ASIG5V.n9631 0.0380882
R49623 ASIG5V.n9633 ASIG5V.n9632 0.0380882
R49624 ASIG5V.n9633 ASIG5V.n9458 0.0380882
R49625 ASIG5V.n9643 ASIG5V.n9458 0.0380882
R49626 ASIG5V.n9644 ASIG5V.n9643 0.0380882
R49627 ASIG5V.n9645 ASIG5V.n9644 0.0380882
R49628 ASIG5V.n9645 ASIG5V.n9456 0.0380882
R49629 ASIG5V.n9655 ASIG5V.n9456 0.0380882
R49630 ASIG5V.n9656 ASIG5V.n9655 0.0380882
R49631 ASIG5V.n9657 ASIG5V.n9656 0.0380882
R49632 ASIG5V.n9657 ASIG5V.n9454 0.0380882
R49633 ASIG5V.n9667 ASIG5V.n9454 0.0380882
R49634 ASIG5V.n9668 ASIG5V.n9667 0.0380882
R49635 ASIG5V.n9669 ASIG5V.n9668 0.0380882
R49636 ASIG5V.n9669 ASIG5V.n9452 0.0380882
R49637 ASIG5V.n9679 ASIG5V.n9452 0.0380882
R49638 ASIG5V.n9680 ASIG5V.n9679 0.0380882
R49639 ASIG5V.n9681 ASIG5V.n9680 0.0380882
R49640 ASIG5V.n9681 ASIG5V.n9450 0.0380882
R49641 ASIG5V.n9691 ASIG5V.n9450 0.0380882
R49642 ASIG5V.n9692 ASIG5V.n9691 0.0380882
R49643 ASIG5V.n9693 ASIG5V.n9692 0.0380882
R49644 ASIG5V.n9693 ASIG5V.n9448 0.0380882
R49645 ASIG5V.n9703 ASIG5V.n9448 0.0380882
R49646 ASIG5V.n9704 ASIG5V.n9703 0.0380882
R49647 ASIG5V.n9705 ASIG5V.n9704 0.0380882
R49648 ASIG5V.n9705 ASIG5V.n9446 0.0380882
R49649 ASIG5V.n9715 ASIG5V.n9446 0.0380882
R49650 ASIG5V.n9716 ASIG5V.n9715 0.0380882
R49651 ASIG5V.n9717 ASIG5V.n9716 0.0380882
R49652 ASIG5V.n9717 ASIG5V.n9444 0.0380882
R49653 ASIG5V.n9727 ASIG5V.n9444 0.0380882
R49654 ASIG5V.n9728 ASIG5V.n9727 0.0380882
R49655 ASIG5V.n9729 ASIG5V.n9728 0.0380882
R49656 ASIG5V.n9729 ASIG5V.n5070 0.0380882
R49657 ASIG5V.n9486 ASIG5V.n9485 0.0380882
R49658 ASIG5V.n9490 ASIG5V.n9485 0.0380882
R49659 ASIG5V.n9494 ASIG5V.n9490 0.0380882
R49660 ASIG5V.n9498 ASIG5V.n9494 0.0380882
R49661 ASIG5V.n9498 ASIG5V.n9481 0.0380882
R49662 ASIG5V.n9502 ASIG5V.n9481 0.0380882
R49663 ASIG5V.n9506 ASIG5V.n9502 0.0380882
R49664 ASIG5V.n9510 ASIG5V.n9506 0.0380882
R49665 ASIG5V.n9510 ASIG5V.n9479 0.0380882
R49666 ASIG5V.n9514 ASIG5V.n9479 0.0380882
R49667 ASIG5V.n9518 ASIG5V.n9514 0.0380882
R49668 ASIG5V.n9522 ASIG5V.n9518 0.0380882
R49669 ASIG5V.n9522 ASIG5V.n9477 0.0380882
R49670 ASIG5V.n9526 ASIG5V.n9477 0.0380882
R49671 ASIG5V.n9530 ASIG5V.n9526 0.0380882
R49672 ASIG5V.n9534 ASIG5V.n9530 0.0380882
R49673 ASIG5V.n9534 ASIG5V.n9475 0.0380882
R49674 ASIG5V.n9538 ASIG5V.n9475 0.0380882
R49675 ASIG5V.n9542 ASIG5V.n9538 0.0380882
R49676 ASIG5V.n9546 ASIG5V.n9542 0.0380882
R49677 ASIG5V.n9546 ASIG5V.n9473 0.0380882
R49678 ASIG5V.n9550 ASIG5V.n9473 0.0380882
R49679 ASIG5V.n9554 ASIG5V.n9550 0.0380882
R49680 ASIG5V.n9558 ASIG5V.n9554 0.0380882
R49681 ASIG5V.n9558 ASIG5V.n9471 0.0380882
R49682 ASIG5V.n9562 ASIG5V.n9471 0.0380882
R49683 ASIG5V.n9566 ASIG5V.n9562 0.0380882
R49684 ASIG5V.n9570 ASIG5V.n9566 0.0380882
R49685 ASIG5V.n9570 ASIG5V.n9469 0.0380882
R49686 ASIG5V.n9574 ASIG5V.n9469 0.0380882
R49687 ASIG5V.n9578 ASIG5V.n9574 0.0380882
R49688 ASIG5V.n9582 ASIG5V.n9578 0.0380882
R49689 ASIG5V.n9582 ASIG5V.n9467 0.0380882
R49690 ASIG5V.n9586 ASIG5V.n9467 0.0380882
R49691 ASIG5V.n9590 ASIG5V.n9586 0.0380882
R49692 ASIG5V.n9594 ASIG5V.n9590 0.0380882
R49693 ASIG5V.n9594 ASIG5V.n9465 0.0380882
R49694 ASIG5V.n9598 ASIG5V.n9465 0.0380882
R49695 ASIG5V.n9602 ASIG5V.n9598 0.0380882
R49696 ASIG5V.n9606 ASIG5V.n9602 0.0380882
R49697 ASIG5V.n9606 ASIG5V.n9463 0.0380882
R49698 ASIG5V.n9610 ASIG5V.n9463 0.0380882
R49699 ASIG5V.n9614 ASIG5V.n9610 0.0380882
R49700 ASIG5V.n9618 ASIG5V.n9614 0.0380882
R49701 ASIG5V.n9618 ASIG5V.n9461 0.0380882
R49702 ASIG5V.n9622 ASIG5V.n9461 0.0380882
R49703 ASIG5V.n9626 ASIG5V.n9622 0.0380882
R49704 ASIG5V.n9630 ASIG5V.n9626 0.0380882
R49705 ASIG5V.n9630 ASIG5V.n9459 0.0380882
R49706 ASIG5V.n9634 ASIG5V.n9459 0.0380882
R49707 ASIG5V.n9638 ASIG5V.n9634 0.0380882
R49708 ASIG5V.n9642 ASIG5V.n9638 0.0380882
R49709 ASIG5V.n9642 ASIG5V.n9457 0.0380882
R49710 ASIG5V.n9646 ASIG5V.n9457 0.0380882
R49711 ASIG5V.n9650 ASIG5V.n9646 0.0380882
R49712 ASIG5V.n9654 ASIG5V.n9650 0.0380882
R49713 ASIG5V.n9654 ASIG5V.n9455 0.0380882
R49714 ASIG5V.n9658 ASIG5V.n9455 0.0380882
R49715 ASIG5V.n9662 ASIG5V.n9658 0.0380882
R49716 ASIG5V.n9666 ASIG5V.n9662 0.0380882
R49717 ASIG5V.n9666 ASIG5V.n9453 0.0380882
R49718 ASIG5V.n9670 ASIG5V.n9453 0.0380882
R49719 ASIG5V.n9674 ASIG5V.n9670 0.0380882
R49720 ASIG5V.n9678 ASIG5V.n9674 0.0380882
R49721 ASIG5V.n9678 ASIG5V.n9451 0.0380882
R49722 ASIG5V.n9682 ASIG5V.n9451 0.0380882
R49723 ASIG5V.n9686 ASIG5V.n9682 0.0380882
R49724 ASIG5V.n9690 ASIG5V.n9686 0.0380882
R49725 ASIG5V.n9690 ASIG5V.n9449 0.0380882
R49726 ASIG5V.n9694 ASIG5V.n9449 0.0380882
R49727 ASIG5V.n9698 ASIG5V.n9694 0.0380882
R49728 ASIG5V.n9702 ASIG5V.n9698 0.0380882
R49729 ASIG5V.n9702 ASIG5V.n9447 0.0380882
R49730 ASIG5V.n9706 ASIG5V.n9447 0.0380882
R49731 ASIG5V.n9710 ASIG5V.n9706 0.0380882
R49732 ASIG5V.n9714 ASIG5V.n9710 0.0380882
R49733 ASIG5V.n9714 ASIG5V.n9445 0.0380882
R49734 ASIG5V.n9718 ASIG5V.n9445 0.0380882
R49735 ASIG5V.n9722 ASIG5V.n9718 0.0380882
R49736 ASIG5V.n9726 ASIG5V.n9722 0.0380882
R49737 ASIG5V.n9726 ASIG5V.n9443 0.0380882
R49738 ASIG5V.n9730 ASIG5V.n9443 0.0380882
R49739 ASIG5V.n9730 ASIG5V.n9442 0.0380882
R49740 ASIG5V.n5216 ASIG5V.n5215 0.0380882
R49741 ASIG5V.n5217 ASIG5V.n5216 0.0380882
R49742 ASIG5V.n5217 ASIG5V.n5210 0.0380882
R49743 ASIG5V.n5227 ASIG5V.n5210 0.0380882
R49744 ASIG5V.n5228 ASIG5V.n5227 0.0380882
R49745 ASIG5V.n5229 ASIG5V.n5228 0.0380882
R49746 ASIG5V.n5229 ASIG5V.n5208 0.0380882
R49747 ASIG5V.n5239 ASIG5V.n5208 0.0380882
R49748 ASIG5V.n5240 ASIG5V.n5239 0.0380882
R49749 ASIG5V.n5241 ASIG5V.n5240 0.0380882
R49750 ASIG5V.n5241 ASIG5V.n5206 0.0380882
R49751 ASIG5V.n5251 ASIG5V.n5206 0.0380882
R49752 ASIG5V.n5252 ASIG5V.n5251 0.0380882
R49753 ASIG5V.n5253 ASIG5V.n5252 0.0380882
R49754 ASIG5V.n5253 ASIG5V.n5204 0.0380882
R49755 ASIG5V.n5263 ASIG5V.n5204 0.0380882
R49756 ASIG5V.n5264 ASIG5V.n5263 0.0380882
R49757 ASIG5V.n5265 ASIG5V.n5264 0.0380882
R49758 ASIG5V.n5265 ASIG5V.n5202 0.0380882
R49759 ASIG5V.n5275 ASIG5V.n5202 0.0380882
R49760 ASIG5V.n5276 ASIG5V.n5275 0.0380882
R49761 ASIG5V.n5277 ASIG5V.n5276 0.0380882
R49762 ASIG5V.n5277 ASIG5V.n5200 0.0380882
R49763 ASIG5V.n5287 ASIG5V.n5200 0.0380882
R49764 ASIG5V.n5288 ASIG5V.n5287 0.0380882
R49765 ASIG5V.n5289 ASIG5V.n5288 0.0380882
R49766 ASIG5V.n5289 ASIG5V.n5198 0.0380882
R49767 ASIG5V.n5299 ASIG5V.n5198 0.0380882
R49768 ASIG5V.n5300 ASIG5V.n5299 0.0380882
R49769 ASIG5V.n5301 ASIG5V.n5300 0.0380882
R49770 ASIG5V.n5301 ASIG5V.n5196 0.0380882
R49771 ASIG5V.n5311 ASIG5V.n5196 0.0380882
R49772 ASIG5V.n5312 ASIG5V.n5311 0.0380882
R49773 ASIG5V.n5313 ASIG5V.n5312 0.0380882
R49774 ASIG5V.n5313 ASIG5V.n5194 0.0380882
R49775 ASIG5V.n5323 ASIG5V.n5194 0.0380882
R49776 ASIG5V.n5324 ASIG5V.n5323 0.0380882
R49777 ASIG5V.n5325 ASIG5V.n5324 0.0380882
R49778 ASIG5V.n5325 ASIG5V.n5192 0.0380882
R49779 ASIG5V.n5335 ASIG5V.n5192 0.0380882
R49780 ASIG5V.n5336 ASIG5V.n5335 0.0380882
R49781 ASIG5V.n5337 ASIG5V.n5336 0.0380882
R49782 ASIG5V.n5337 ASIG5V.n5190 0.0380882
R49783 ASIG5V.n5347 ASIG5V.n5190 0.0380882
R49784 ASIG5V.n5348 ASIG5V.n5347 0.0380882
R49785 ASIG5V.n5349 ASIG5V.n5348 0.0380882
R49786 ASIG5V.n5349 ASIG5V.n5188 0.0380882
R49787 ASIG5V.n5359 ASIG5V.n5188 0.0380882
R49788 ASIG5V.n5360 ASIG5V.n5359 0.0380882
R49789 ASIG5V.n5361 ASIG5V.n5360 0.0380882
R49790 ASIG5V.n5361 ASIG5V.n5186 0.0380882
R49791 ASIG5V.n5371 ASIG5V.n5186 0.0380882
R49792 ASIG5V.n5372 ASIG5V.n5371 0.0380882
R49793 ASIG5V.n5373 ASIG5V.n5372 0.0380882
R49794 ASIG5V.n5373 ASIG5V.n5184 0.0380882
R49795 ASIG5V.n5383 ASIG5V.n5184 0.0380882
R49796 ASIG5V.n5384 ASIG5V.n5383 0.0380882
R49797 ASIG5V.n5385 ASIG5V.n5384 0.0380882
R49798 ASIG5V.n5385 ASIG5V.n5182 0.0380882
R49799 ASIG5V.n5395 ASIG5V.n5182 0.0380882
R49800 ASIG5V.n5396 ASIG5V.n5395 0.0380882
R49801 ASIG5V.n5397 ASIG5V.n5396 0.0380882
R49802 ASIG5V.n5397 ASIG5V.n5180 0.0380882
R49803 ASIG5V.n5407 ASIG5V.n5180 0.0380882
R49804 ASIG5V.n5408 ASIG5V.n5407 0.0380882
R49805 ASIG5V.n5409 ASIG5V.n5408 0.0380882
R49806 ASIG5V.n5409 ASIG5V.n5178 0.0380882
R49807 ASIG5V.n5419 ASIG5V.n5178 0.0380882
R49808 ASIG5V.n5420 ASIG5V.n5419 0.0380882
R49809 ASIG5V.n5421 ASIG5V.n5420 0.0380882
R49810 ASIG5V.n5421 ASIG5V.n5176 0.0380882
R49811 ASIG5V.n5431 ASIG5V.n5176 0.0380882
R49812 ASIG5V.n5432 ASIG5V.n5431 0.0380882
R49813 ASIG5V.n5433 ASIG5V.n5432 0.0380882
R49814 ASIG5V.n5433 ASIG5V.n5174 0.0380882
R49815 ASIG5V.n5443 ASIG5V.n5174 0.0380882
R49816 ASIG5V.n5444 ASIG5V.n5443 0.0380882
R49817 ASIG5V.n5445 ASIG5V.n5444 0.0380882
R49818 ASIG5V.n5445 ASIG5V.n5172 0.0380882
R49819 ASIG5V.n5455 ASIG5V.n5172 0.0380882
R49820 ASIG5V.n5456 ASIG5V.n5455 0.0380882
R49821 ASIG5V.n9427 ASIG5V.n5456 0.0380882
R49822 ASIG5V.n9427 ASIG5V.n9426 0.0380882
R49823 ASIG5V.n5214 ASIG5V.n5213 0.0380882
R49824 ASIG5V.n5218 ASIG5V.n5213 0.0380882
R49825 ASIG5V.n5222 ASIG5V.n5218 0.0380882
R49826 ASIG5V.n5226 ASIG5V.n5222 0.0380882
R49827 ASIG5V.n5226 ASIG5V.n5209 0.0380882
R49828 ASIG5V.n5230 ASIG5V.n5209 0.0380882
R49829 ASIG5V.n5234 ASIG5V.n5230 0.0380882
R49830 ASIG5V.n5238 ASIG5V.n5234 0.0380882
R49831 ASIG5V.n5238 ASIG5V.n5207 0.0380882
R49832 ASIG5V.n5242 ASIG5V.n5207 0.0380882
R49833 ASIG5V.n5246 ASIG5V.n5242 0.0380882
R49834 ASIG5V.n5250 ASIG5V.n5246 0.0380882
R49835 ASIG5V.n5250 ASIG5V.n5205 0.0380882
R49836 ASIG5V.n5254 ASIG5V.n5205 0.0380882
R49837 ASIG5V.n5258 ASIG5V.n5254 0.0380882
R49838 ASIG5V.n5262 ASIG5V.n5258 0.0380882
R49839 ASIG5V.n5262 ASIG5V.n5203 0.0380882
R49840 ASIG5V.n5266 ASIG5V.n5203 0.0380882
R49841 ASIG5V.n5270 ASIG5V.n5266 0.0380882
R49842 ASIG5V.n5274 ASIG5V.n5270 0.0380882
R49843 ASIG5V.n5274 ASIG5V.n5201 0.0380882
R49844 ASIG5V.n5278 ASIG5V.n5201 0.0380882
R49845 ASIG5V.n5282 ASIG5V.n5278 0.0380882
R49846 ASIG5V.n5286 ASIG5V.n5282 0.0380882
R49847 ASIG5V.n5286 ASIG5V.n5199 0.0380882
R49848 ASIG5V.n5290 ASIG5V.n5199 0.0380882
R49849 ASIG5V.n5294 ASIG5V.n5290 0.0380882
R49850 ASIG5V.n5298 ASIG5V.n5294 0.0380882
R49851 ASIG5V.n5298 ASIG5V.n5197 0.0380882
R49852 ASIG5V.n5302 ASIG5V.n5197 0.0380882
R49853 ASIG5V.n5306 ASIG5V.n5302 0.0380882
R49854 ASIG5V.n5310 ASIG5V.n5306 0.0380882
R49855 ASIG5V.n5310 ASIG5V.n5195 0.0380882
R49856 ASIG5V.n5314 ASIG5V.n5195 0.0380882
R49857 ASIG5V.n5318 ASIG5V.n5314 0.0380882
R49858 ASIG5V.n5322 ASIG5V.n5318 0.0380882
R49859 ASIG5V.n5322 ASIG5V.n5193 0.0380882
R49860 ASIG5V.n5326 ASIG5V.n5193 0.0380882
R49861 ASIG5V.n5330 ASIG5V.n5326 0.0380882
R49862 ASIG5V.n5334 ASIG5V.n5330 0.0380882
R49863 ASIG5V.n5334 ASIG5V.n5191 0.0380882
R49864 ASIG5V.n5338 ASIG5V.n5191 0.0380882
R49865 ASIG5V.n5342 ASIG5V.n5338 0.0380882
R49866 ASIG5V.n5346 ASIG5V.n5342 0.0380882
R49867 ASIG5V.n5346 ASIG5V.n5189 0.0380882
R49868 ASIG5V.n5350 ASIG5V.n5189 0.0380882
R49869 ASIG5V.n5354 ASIG5V.n5350 0.0380882
R49870 ASIG5V.n5358 ASIG5V.n5354 0.0380882
R49871 ASIG5V.n5358 ASIG5V.n5187 0.0380882
R49872 ASIG5V.n5362 ASIG5V.n5187 0.0380882
R49873 ASIG5V.n5366 ASIG5V.n5362 0.0380882
R49874 ASIG5V.n5370 ASIG5V.n5366 0.0380882
R49875 ASIG5V.n5370 ASIG5V.n5185 0.0380882
R49876 ASIG5V.n5374 ASIG5V.n5185 0.0380882
R49877 ASIG5V.n5378 ASIG5V.n5374 0.0380882
R49878 ASIG5V.n5382 ASIG5V.n5378 0.0380882
R49879 ASIG5V.n5382 ASIG5V.n5183 0.0380882
R49880 ASIG5V.n5386 ASIG5V.n5183 0.0380882
R49881 ASIG5V.n5390 ASIG5V.n5386 0.0380882
R49882 ASIG5V.n5394 ASIG5V.n5390 0.0380882
R49883 ASIG5V.n5394 ASIG5V.n5181 0.0380882
R49884 ASIG5V.n5398 ASIG5V.n5181 0.0380882
R49885 ASIG5V.n5402 ASIG5V.n5398 0.0380882
R49886 ASIG5V.n5406 ASIG5V.n5402 0.0380882
R49887 ASIG5V.n5406 ASIG5V.n5179 0.0380882
R49888 ASIG5V.n5410 ASIG5V.n5179 0.0380882
R49889 ASIG5V.n5414 ASIG5V.n5410 0.0380882
R49890 ASIG5V.n5418 ASIG5V.n5414 0.0380882
R49891 ASIG5V.n5418 ASIG5V.n5177 0.0380882
R49892 ASIG5V.n5422 ASIG5V.n5177 0.0380882
R49893 ASIG5V.n5426 ASIG5V.n5422 0.0380882
R49894 ASIG5V.n5430 ASIG5V.n5426 0.0380882
R49895 ASIG5V.n5430 ASIG5V.n5175 0.0380882
R49896 ASIG5V.n5434 ASIG5V.n5175 0.0380882
R49897 ASIG5V.n5438 ASIG5V.n5434 0.0380882
R49898 ASIG5V.n5442 ASIG5V.n5438 0.0380882
R49899 ASIG5V.n5442 ASIG5V.n5173 0.0380882
R49900 ASIG5V.n5446 ASIG5V.n5173 0.0380882
R49901 ASIG5V.n5450 ASIG5V.n5446 0.0380882
R49902 ASIG5V.n5454 ASIG5V.n5450 0.0380882
R49903 ASIG5V.n5454 ASIG5V.n5171 0.0380882
R49904 ASIG5V.n9428 ASIG5V.n5171 0.0380882
R49905 ASIG5V.n9428 ASIG5V.n5168 0.0380882
R49906 ASIG5V.n7960 ASIG5V.n7959 0.0380882
R49907 ASIG5V.n7959 ASIG5V.n7717 0.0380882
R49908 ASIG5V.n7953 ASIG5V.n7717 0.0380882
R49909 ASIG5V.n7953 ASIG5V.n7952 0.0380882
R49910 ASIG5V.n7952 ASIG5V.n7951 0.0380882
R49911 ASIG5V.n7951 ASIG5V.n7720 0.0380882
R49912 ASIG5V.n7944 ASIG5V.n7720 0.0380882
R49913 ASIG5V.n7944 ASIG5V.n7943 0.0380882
R49914 ASIG5V.n7943 ASIG5V.n7942 0.0380882
R49915 ASIG5V.n7942 ASIG5V.n7723 0.0380882
R49916 ASIG5V.n7935 ASIG5V.n7723 0.0380882
R49917 ASIG5V.n7935 ASIG5V.n7934 0.0380882
R49918 ASIG5V.n7934 ASIG5V.n7933 0.0380882
R49919 ASIG5V.n7933 ASIG5V.n7726 0.0380882
R49920 ASIG5V.n7926 ASIG5V.n7726 0.0380882
R49921 ASIG5V.n7926 ASIG5V.n7925 0.0380882
R49922 ASIG5V.n7925 ASIG5V.n7924 0.0380882
R49923 ASIG5V.n7924 ASIG5V.n7729 0.0380882
R49924 ASIG5V.n7917 ASIG5V.n7729 0.0380882
R49925 ASIG5V.n7917 ASIG5V.n7916 0.0380882
R49926 ASIG5V.n7916 ASIG5V.n7915 0.0380882
R49927 ASIG5V.n7915 ASIG5V.n7732 0.0380882
R49928 ASIG5V.n7908 ASIG5V.n7732 0.0380882
R49929 ASIG5V.n7908 ASIG5V.n7907 0.0380882
R49930 ASIG5V.n7907 ASIG5V.n7906 0.0380882
R49931 ASIG5V.n7906 ASIG5V.n7735 0.0380882
R49932 ASIG5V.n7899 ASIG5V.n7735 0.0380882
R49933 ASIG5V.n7899 ASIG5V.n7898 0.0380882
R49934 ASIG5V.n7898 ASIG5V.n7897 0.0380882
R49935 ASIG5V.n7897 ASIG5V.n7738 0.0380882
R49936 ASIG5V.n7890 ASIG5V.n7738 0.0380882
R49937 ASIG5V.n7890 ASIG5V.n7889 0.0380882
R49938 ASIG5V.n7889 ASIG5V.n7888 0.0380882
R49939 ASIG5V.n7888 ASIG5V.n7741 0.0380882
R49940 ASIG5V.n7881 ASIG5V.n7741 0.0380882
R49941 ASIG5V.n7881 ASIG5V.n7880 0.0380882
R49942 ASIG5V.n7880 ASIG5V.n7879 0.0380882
R49943 ASIG5V.n7879 ASIG5V.n7744 0.0380882
R49944 ASIG5V.n7872 ASIG5V.n7744 0.0380882
R49945 ASIG5V.n7872 ASIG5V.n7871 0.0380882
R49946 ASIG5V.n7871 ASIG5V.n7870 0.0380882
R49947 ASIG5V.n7870 ASIG5V.n7747 0.0380882
R49948 ASIG5V.n7863 ASIG5V.n7747 0.0380882
R49949 ASIG5V.n7863 ASIG5V.n7862 0.0380882
R49950 ASIG5V.n7862 ASIG5V.n7861 0.0380882
R49951 ASIG5V.n7861 ASIG5V.n7750 0.0380882
R49952 ASIG5V.n7854 ASIG5V.n7750 0.0380882
R49953 ASIG5V.n7854 ASIG5V.n7853 0.0380882
R49954 ASIG5V.n7853 ASIG5V.n7852 0.0380882
R49955 ASIG5V.n7852 ASIG5V.n7753 0.0380882
R49956 ASIG5V.n7845 ASIG5V.n7753 0.0380882
R49957 ASIG5V.n7845 ASIG5V.n7844 0.0380882
R49958 ASIG5V.n7844 ASIG5V.n7843 0.0380882
R49959 ASIG5V.n7843 ASIG5V.n7756 0.0380882
R49960 ASIG5V.n7836 ASIG5V.n7756 0.0380882
R49961 ASIG5V.n7836 ASIG5V.n7835 0.0380882
R49962 ASIG5V.n7835 ASIG5V.n7834 0.0380882
R49963 ASIG5V.n7834 ASIG5V.n7759 0.0380882
R49964 ASIG5V.n7827 ASIG5V.n7759 0.0380882
R49965 ASIG5V.n7827 ASIG5V.n7826 0.0380882
R49966 ASIG5V.n7826 ASIG5V.n7825 0.0380882
R49967 ASIG5V.n7825 ASIG5V.n7762 0.0380882
R49968 ASIG5V.n7818 ASIG5V.n7762 0.0380882
R49969 ASIG5V.n7818 ASIG5V.n7817 0.0380882
R49970 ASIG5V.n7817 ASIG5V.n7816 0.0380882
R49971 ASIG5V.n7816 ASIG5V.n7765 0.0380882
R49972 ASIG5V.n7809 ASIG5V.n7765 0.0380882
R49973 ASIG5V.n7809 ASIG5V.n7808 0.0380882
R49974 ASIG5V.n7808 ASIG5V.n7807 0.0380882
R49975 ASIG5V.n7807 ASIG5V.n7768 0.0380882
R49976 ASIG5V.n7800 ASIG5V.n7768 0.0380882
R49977 ASIG5V.n7800 ASIG5V.n7799 0.0380882
R49978 ASIG5V.n7799 ASIG5V.n7798 0.0380882
R49979 ASIG5V.n7798 ASIG5V.n7771 0.0380882
R49980 ASIG5V.n7791 ASIG5V.n7771 0.0380882
R49981 ASIG5V.n7791 ASIG5V.n7790 0.0380882
R49982 ASIG5V.n7790 ASIG5V.n7789 0.0380882
R49983 ASIG5V.n7789 ASIG5V.n7774 0.0380882
R49984 ASIG5V.n7782 ASIG5V.n7774 0.0380882
R49985 ASIG5V.n7782 ASIG5V.n7781 0.0380882
R49986 ASIG5V.n7781 ASIG5V.n7780 0.0380882
R49987 ASIG5V.n7780 ASIG5V.n7777 0.0380882
R49988 ASIG5V.n7777 ASIG5V.n5557 0.0380882
R49989 ASIG5V.n7958 ASIG5V.n5509 0.0380882
R49990 ASIG5V.n7958 ASIG5V.n7957 0.0380882
R49991 ASIG5V.n7957 ASIG5V.n7955 0.0380882
R49992 ASIG5V.n7955 ASIG5V.n7719 0.0380882
R49993 ASIG5V.n7950 ASIG5V.n7719 0.0380882
R49994 ASIG5V.n7950 ASIG5V.n7948 0.0380882
R49995 ASIG5V.n7948 ASIG5V.n7946 0.0380882
R49996 ASIG5V.n7946 ASIG5V.n7722 0.0380882
R49997 ASIG5V.n7941 ASIG5V.n7722 0.0380882
R49998 ASIG5V.n7941 ASIG5V.n7939 0.0380882
R49999 ASIG5V.n7939 ASIG5V.n7937 0.0380882
R50000 ASIG5V.n7937 ASIG5V.n7725 0.0380882
R50001 ASIG5V.n7932 ASIG5V.n7725 0.0380882
R50002 ASIG5V.n7932 ASIG5V.n7930 0.0380882
R50003 ASIG5V.n7930 ASIG5V.n7928 0.0380882
R50004 ASIG5V.n7928 ASIG5V.n7728 0.0380882
R50005 ASIG5V.n7923 ASIG5V.n7728 0.0380882
R50006 ASIG5V.n7923 ASIG5V.n7921 0.0380882
R50007 ASIG5V.n7921 ASIG5V.n7919 0.0380882
R50008 ASIG5V.n7919 ASIG5V.n7731 0.0380882
R50009 ASIG5V.n7914 ASIG5V.n7731 0.0380882
R50010 ASIG5V.n7914 ASIG5V.n7912 0.0380882
R50011 ASIG5V.n7912 ASIG5V.n7910 0.0380882
R50012 ASIG5V.n7910 ASIG5V.n7734 0.0380882
R50013 ASIG5V.n7905 ASIG5V.n7734 0.0380882
R50014 ASIG5V.n7905 ASIG5V.n7903 0.0380882
R50015 ASIG5V.n7903 ASIG5V.n7901 0.0380882
R50016 ASIG5V.n7901 ASIG5V.n7737 0.0380882
R50017 ASIG5V.n7896 ASIG5V.n7737 0.0380882
R50018 ASIG5V.n7896 ASIG5V.n7894 0.0380882
R50019 ASIG5V.n7894 ASIG5V.n7892 0.0380882
R50020 ASIG5V.n7892 ASIG5V.n7740 0.0380882
R50021 ASIG5V.n7887 ASIG5V.n7740 0.0380882
R50022 ASIG5V.n7887 ASIG5V.n7885 0.0380882
R50023 ASIG5V.n7885 ASIG5V.n7883 0.0380882
R50024 ASIG5V.n7883 ASIG5V.n7743 0.0380882
R50025 ASIG5V.n7878 ASIG5V.n7743 0.0380882
R50026 ASIG5V.n7878 ASIG5V.n7876 0.0380882
R50027 ASIG5V.n7876 ASIG5V.n7874 0.0380882
R50028 ASIG5V.n7874 ASIG5V.n7746 0.0380882
R50029 ASIG5V.n7869 ASIG5V.n7746 0.0380882
R50030 ASIG5V.n7869 ASIG5V.n7867 0.0380882
R50031 ASIG5V.n7867 ASIG5V.n7865 0.0380882
R50032 ASIG5V.n7865 ASIG5V.n7749 0.0380882
R50033 ASIG5V.n7860 ASIG5V.n7749 0.0380882
R50034 ASIG5V.n7860 ASIG5V.n7858 0.0380882
R50035 ASIG5V.n7858 ASIG5V.n7856 0.0380882
R50036 ASIG5V.n7856 ASIG5V.n7752 0.0380882
R50037 ASIG5V.n7851 ASIG5V.n7752 0.0380882
R50038 ASIG5V.n7851 ASIG5V.n7849 0.0380882
R50039 ASIG5V.n7849 ASIG5V.n7847 0.0380882
R50040 ASIG5V.n7847 ASIG5V.n7755 0.0380882
R50041 ASIG5V.n7842 ASIG5V.n7755 0.0380882
R50042 ASIG5V.n7842 ASIG5V.n7840 0.0380882
R50043 ASIG5V.n7840 ASIG5V.n7838 0.0380882
R50044 ASIG5V.n7838 ASIG5V.n7758 0.0380882
R50045 ASIG5V.n7833 ASIG5V.n7758 0.0380882
R50046 ASIG5V.n7833 ASIG5V.n7831 0.0380882
R50047 ASIG5V.n7831 ASIG5V.n7829 0.0380882
R50048 ASIG5V.n7829 ASIG5V.n7761 0.0380882
R50049 ASIG5V.n7824 ASIG5V.n7761 0.0380882
R50050 ASIG5V.n7824 ASIG5V.n7822 0.0380882
R50051 ASIG5V.n7822 ASIG5V.n7820 0.0380882
R50052 ASIG5V.n7820 ASIG5V.n7764 0.0380882
R50053 ASIG5V.n7815 ASIG5V.n7764 0.0380882
R50054 ASIG5V.n7815 ASIG5V.n7813 0.0380882
R50055 ASIG5V.n7813 ASIG5V.n7811 0.0380882
R50056 ASIG5V.n7811 ASIG5V.n7767 0.0380882
R50057 ASIG5V.n7806 ASIG5V.n7767 0.0380882
R50058 ASIG5V.n7806 ASIG5V.n7804 0.0380882
R50059 ASIG5V.n7804 ASIG5V.n7802 0.0380882
R50060 ASIG5V.n7802 ASIG5V.n7770 0.0380882
R50061 ASIG5V.n7797 ASIG5V.n7770 0.0380882
R50062 ASIG5V.n7797 ASIG5V.n7795 0.0380882
R50063 ASIG5V.n7795 ASIG5V.n7793 0.0380882
R50064 ASIG5V.n7793 ASIG5V.n7773 0.0380882
R50065 ASIG5V.n7788 ASIG5V.n7773 0.0380882
R50066 ASIG5V.n7788 ASIG5V.n7786 0.0380882
R50067 ASIG5V.n7786 ASIG5V.n7784 0.0380882
R50068 ASIG5V.n7784 ASIG5V.n7776 0.0380882
R50069 ASIG5V.n7779 ASIG5V.n7776 0.0380882
R50070 ASIG5V.n7779 ASIG5V.n5556 0.0380882
R50071 ASIG5V.n9414 ASIG5V.n5556 0.0380882
R50072 ASIG5V.n5907 ASIG5V.n5573 0.0380882
R50073 ASIG5V.n5899 ASIG5V.n5573 0.0380882
R50074 ASIG5V.n5899 ASIG5V.n5898 0.0380882
R50075 ASIG5V.n5898 ASIG5V.n5897 0.0380882
R50076 ASIG5V.n5897 ASIG5V.n5577 0.0380882
R50077 ASIG5V.n5889 ASIG5V.n5577 0.0380882
R50078 ASIG5V.n5889 ASIG5V.n5888 0.0380882
R50079 ASIG5V.n5888 ASIG5V.n5887 0.0380882
R50080 ASIG5V.n5887 ASIG5V.n5583 0.0380882
R50081 ASIG5V.n5879 ASIG5V.n5583 0.0380882
R50082 ASIG5V.n5879 ASIG5V.n5878 0.0380882
R50083 ASIG5V.n5878 ASIG5V.n5877 0.0380882
R50084 ASIG5V.n5877 ASIG5V.n5589 0.0380882
R50085 ASIG5V.n5869 ASIG5V.n5589 0.0380882
R50086 ASIG5V.n5869 ASIG5V.n5868 0.0380882
R50087 ASIG5V.n5868 ASIG5V.n5867 0.0380882
R50088 ASIG5V.n5867 ASIG5V.n5595 0.0380882
R50089 ASIG5V.n5859 ASIG5V.n5595 0.0380882
R50090 ASIG5V.n5859 ASIG5V.n5858 0.0380882
R50091 ASIG5V.n5858 ASIG5V.n5857 0.0380882
R50092 ASIG5V.n5857 ASIG5V.n5601 0.0380882
R50093 ASIG5V.n5849 ASIG5V.n5601 0.0380882
R50094 ASIG5V.n5849 ASIG5V.n5848 0.0380882
R50095 ASIG5V.n5848 ASIG5V.n5847 0.0380882
R50096 ASIG5V.n5847 ASIG5V.n5607 0.0380882
R50097 ASIG5V.n5839 ASIG5V.n5607 0.0380882
R50098 ASIG5V.n5839 ASIG5V.n5838 0.0380882
R50099 ASIG5V.n5838 ASIG5V.n5837 0.0380882
R50100 ASIG5V.n5837 ASIG5V.n5613 0.0380882
R50101 ASIG5V.n5829 ASIG5V.n5613 0.0380882
R50102 ASIG5V.n5829 ASIG5V.n5828 0.0380882
R50103 ASIG5V.n5828 ASIG5V.n5827 0.0380882
R50104 ASIG5V.n5827 ASIG5V.n5619 0.0380882
R50105 ASIG5V.n5819 ASIG5V.n5619 0.0380882
R50106 ASIG5V.n5819 ASIG5V.n5818 0.0380882
R50107 ASIG5V.n5818 ASIG5V.n5817 0.0380882
R50108 ASIG5V.n5817 ASIG5V.n5625 0.0380882
R50109 ASIG5V.n5809 ASIG5V.n5625 0.0380882
R50110 ASIG5V.n5809 ASIG5V.n5808 0.0380882
R50111 ASIG5V.n5808 ASIG5V.n5807 0.0380882
R50112 ASIG5V.n5807 ASIG5V.n5631 0.0380882
R50113 ASIG5V.n5799 ASIG5V.n5631 0.0380882
R50114 ASIG5V.n5799 ASIG5V.n5798 0.0380882
R50115 ASIG5V.n5798 ASIG5V.n5797 0.0380882
R50116 ASIG5V.n5797 ASIG5V.n5637 0.0380882
R50117 ASIG5V.n5789 ASIG5V.n5637 0.0380882
R50118 ASIG5V.n5789 ASIG5V.n5788 0.0380882
R50119 ASIG5V.n5788 ASIG5V.n5787 0.0380882
R50120 ASIG5V.n5787 ASIG5V.n5643 0.0380882
R50121 ASIG5V.n5779 ASIG5V.n5643 0.0380882
R50122 ASIG5V.n5779 ASIG5V.n5778 0.0380882
R50123 ASIG5V.n5778 ASIG5V.n5777 0.0380882
R50124 ASIG5V.n5777 ASIG5V.n5649 0.0380882
R50125 ASIG5V.n5769 ASIG5V.n5649 0.0380882
R50126 ASIG5V.n5769 ASIG5V.n5768 0.0380882
R50127 ASIG5V.n5768 ASIG5V.n5767 0.0380882
R50128 ASIG5V.n5767 ASIG5V.n5655 0.0380882
R50129 ASIG5V.n5759 ASIG5V.n5655 0.0380882
R50130 ASIG5V.n5759 ASIG5V.n5758 0.0380882
R50131 ASIG5V.n5758 ASIG5V.n5757 0.0380882
R50132 ASIG5V.n5757 ASIG5V.n5661 0.0380882
R50133 ASIG5V.n5749 ASIG5V.n5661 0.0380882
R50134 ASIG5V.n5749 ASIG5V.n5748 0.0380882
R50135 ASIG5V.n5748 ASIG5V.n5747 0.0380882
R50136 ASIG5V.n5747 ASIG5V.n5667 0.0380882
R50137 ASIG5V.n5739 ASIG5V.n5667 0.0380882
R50138 ASIG5V.n5739 ASIG5V.n5738 0.0380882
R50139 ASIG5V.n5738 ASIG5V.n5737 0.0380882
R50140 ASIG5V.n5737 ASIG5V.n5673 0.0380882
R50141 ASIG5V.n5729 ASIG5V.n5673 0.0380882
R50142 ASIG5V.n5729 ASIG5V.n5728 0.0380882
R50143 ASIG5V.n5728 ASIG5V.n5727 0.0380882
R50144 ASIG5V.n5727 ASIG5V.n5679 0.0380882
R50145 ASIG5V.n5719 ASIG5V.n5679 0.0380882
R50146 ASIG5V.n5719 ASIG5V.n5718 0.0380882
R50147 ASIG5V.n5718 ASIG5V.n5717 0.0380882
R50148 ASIG5V.n5717 ASIG5V.n5685 0.0380882
R50149 ASIG5V.n5709 ASIG5V.n5685 0.0380882
R50150 ASIG5V.n5709 ASIG5V.n5708 0.0380882
R50151 ASIG5V.n5708 ASIG5V.n5707 0.0380882
R50152 ASIG5V.n5707 ASIG5V.n5691 0.0380882
R50153 ASIG5V.n5699 ASIG5V.n5691 0.0380882
R50154 ASIG5V.n5699 ASIG5V.n5698 0.0380882
R50155 ASIG5V.n5906 ASIG5V.n5574 0.0380882
R50156 ASIG5V.n5900 ASIG5V.n5574 0.0380882
R50157 ASIG5V.n5900 ASIG5V.n5576 0.0380882
R50158 ASIG5V.n5896 ASIG5V.n5576 0.0380882
R50159 ASIG5V.n5896 ASIG5V.n5578 0.0380882
R50160 ASIG5V.n5890 ASIG5V.n5578 0.0380882
R50161 ASIG5V.n5890 ASIG5V.n5582 0.0380882
R50162 ASIG5V.n5886 ASIG5V.n5582 0.0380882
R50163 ASIG5V.n5886 ASIG5V.n5584 0.0380882
R50164 ASIG5V.n5880 ASIG5V.n5584 0.0380882
R50165 ASIG5V.n5880 ASIG5V.n5588 0.0380882
R50166 ASIG5V.n5876 ASIG5V.n5588 0.0380882
R50167 ASIG5V.n5876 ASIG5V.n5590 0.0380882
R50168 ASIG5V.n5870 ASIG5V.n5590 0.0380882
R50169 ASIG5V.n5870 ASIG5V.n5594 0.0380882
R50170 ASIG5V.n5866 ASIG5V.n5594 0.0380882
R50171 ASIG5V.n5866 ASIG5V.n5596 0.0380882
R50172 ASIG5V.n5860 ASIG5V.n5596 0.0380882
R50173 ASIG5V.n5860 ASIG5V.n5600 0.0380882
R50174 ASIG5V.n5856 ASIG5V.n5600 0.0380882
R50175 ASIG5V.n5856 ASIG5V.n5602 0.0380882
R50176 ASIG5V.n5850 ASIG5V.n5602 0.0380882
R50177 ASIG5V.n5850 ASIG5V.n5606 0.0380882
R50178 ASIG5V.n5846 ASIG5V.n5606 0.0380882
R50179 ASIG5V.n5846 ASIG5V.n5608 0.0380882
R50180 ASIG5V.n5840 ASIG5V.n5608 0.0380882
R50181 ASIG5V.n5840 ASIG5V.n5612 0.0380882
R50182 ASIG5V.n5836 ASIG5V.n5612 0.0380882
R50183 ASIG5V.n5836 ASIG5V.n5614 0.0380882
R50184 ASIG5V.n5830 ASIG5V.n5614 0.0380882
R50185 ASIG5V.n5830 ASIG5V.n5618 0.0380882
R50186 ASIG5V.n5826 ASIG5V.n5618 0.0380882
R50187 ASIG5V.n5826 ASIG5V.n5620 0.0380882
R50188 ASIG5V.n5820 ASIG5V.n5620 0.0380882
R50189 ASIG5V.n5820 ASIG5V.n5624 0.0380882
R50190 ASIG5V.n5816 ASIG5V.n5624 0.0380882
R50191 ASIG5V.n5816 ASIG5V.n5626 0.0380882
R50192 ASIG5V.n5810 ASIG5V.n5626 0.0380882
R50193 ASIG5V.n5810 ASIG5V.n5630 0.0380882
R50194 ASIG5V.n5806 ASIG5V.n5630 0.0380882
R50195 ASIG5V.n5806 ASIG5V.n5632 0.0380882
R50196 ASIG5V.n5800 ASIG5V.n5632 0.0380882
R50197 ASIG5V.n5800 ASIG5V.n5636 0.0380882
R50198 ASIG5V.n5796 ASIG5V.n5636 0.0380882
R50199 ASIG5V.n5796 ASIG5V.n5638 0.0380882
R50200 ASIG5V.n5790 ASIG5V.n5638 0.0380882
R50201 ASIG5V.n5790 ASIG5V.n5642 0.0380882
R50202 ASIG5V.n5786 ASIG5V.n5642 0.0380882
R50203 ASIG5V.n5786 ASIG5V.n5644 0.0380882
R50204 ASIG5V.n5780 ASIG5V.n5644 0.0380882
R50205 ASIG5V.n5780 ASIG5V.n5648 0.0380882
R50206 ASIG5V.n5776 ASIG5V.n5648 0.0380882
R50207 ASIG5V.n5776 ASIG5V.n5650 0.0380882
R50208 ASIG5V.n5770 ASIG5V.n5650 0.0380882
R50209 ASIG5V.n5770 ASIG5V.n5654 0.0380882
R50210 ASIG5V.n5766 ASIG5V.n5654 0.0380882
R50211 ASIG5V.n5766 ASIG5V.n5656 0.0380882
R50212 ASIG5V.n5760 ASIG5V.n5656 0.0380882
R50213 ASIG5V.n5760 ASIG5V.n5660 0.0380882
R50214 ASIG5V.n5756 ASIG5V.n5660 0.0380882
R50215 ASIG5V.n5756 ASIG5V.n5662 0.0380882
R50216 ASIG5V.n5750 ASIG5V.n5662 0.0380882
R50217 ASIG5V.n5750 ASIG5V.n5666 0.0380882
R50218 ASIG5V.n5746 ASIG5V.n5666 0.0380882
R50219 ASIG5V.n5746 ASIG5V.n5668 0.0380882
R50220 ASIG5V.n5740 ASIG5V.n5668 0.0380882
R50221 ASIG5V.n5740 ASIG5V.n5672 0.0380882
R50222 ASIG5V.n5736 ASIG5V.n5672 0.0380882
R50223 ASIG5V.n5736 ASIG5V.n5674 0.0380882
R50224 ASIG5V.n5730 ASIG5V.n5674 0.0380882
R50225 ASIG5V.n5730 ASIG5V.n5678 0.0380882
R50226 ASIG5V.n5726 ASIG5V.n5678 0.0380882
R50227 ASIG5V.n5726 ASIG5V.n5680 0.0380882
R50228 ASIG5V.n5720 ASIG5V.n5680 0.0380882
R50229 ASIG5V.n5720 ASIG5V.n5684 0.0380882
R50230 ASIG5V.n5716 ASIG5V.n5684 0.0380882
R50231 ASIG5V.n5716 ASIG5V.n5686 0.0380882
R50232 ASIG5V.n5710 ASIG5V.n5686 0.0380882
R50233 ASIG5V.n5710 ASIG5V.n5690 0.0380882
R50234 ASIG5V.n5706 ASIG5V.n5690 0.0380882
R50235 ASIG5V.n5706 ASIG5V.n5692 0.0380882
R50236 ASIG5V.n5700 ASIG5V.n5692 0.0380882
R50237 ASIG5V.n5700 ASIG5V.n5697 0.0380882
R50238 ASIG5V.n6065 ASIG5V.n6063 0.0380882
R50239 ASIG5V.n6066 ASIG5V.n6065 0.0380882
R50240 ASIG5V.n6067 ASIG5V.n6066 0.0380882
R50241 ASIG5V.n6067 ASIG5V.n6060 0.0380882
R50242 ASIG5V.n6074 ASIG5V.n6060 0.0380882
R50243 ASIG5V.n6075 ASIG5V.n6074 0.0380882
R50244 ASIG5V.n6076 ASIG5V.n6075 0.0380882
R50245 ASIG5V.n6076 ASIG5V.n6057 0.0380882
R50246 ASIG5V.n6083 ASIG5V.n6057 0.0380882
R50247 ASIG5V.n6084 ASIG5V.n6083 0.0380882
R50248 ASIG5V.n6085 ASIG5V.n6084 0.0380882
R50249 ASIG5V.n6085 ASIG5V.n6054 0.0380882
R50250 ASIG5V.n6092 ASIG5V.n6054 0.0380882
R50251 ASIG5V.n6093 ASIG5V.n6092 0.0380882
R50252 ASIG5V.n6094 ASIG5V.n6093 0.0380882
R50253 ASIG5V.n6094 ASIG5V.n6051 0.0380882
R50254 ASIG5V.n6101 ASIG5V.n6051 0.0380882
R50255 ASIG5V.n6102 ASIG5V.n6101 0.0380882
R50256 ASIG5V.n6103 ASIG5V.n6102 0.0380882
R50257 ASIG5V.n6103 ASIG5V.n6048 0.0380882
R50258 ASIG5V.n6110 ASIG5V.n6048 0.0380882
R50259 ASIG5V.n6111 ASIG5V.n6110 0.0380882
R50260 ASIG5V.n6112 ASIG5V.n6111 0.0380882
R50261 ASIG5V.n6112 ASIG5V.n6045 0.0380882
R50262 ASIG5V.n6119 ASIG5V.n6045 0.0380882
R50263 ASIG5V.n6120 ASIG5V.n6119 0.0380882
R50264 ASIG5V.n6121 ASIG5V.n6120 0.0380882
R50265 ASIG5V.n6121 ASIG5V.n6042 0.0380882
R50266 ASIG5V.n6128 ASIG5V.n6042 0.0380882
R50267 ASIG5V.n6129 ASIG5V.n6128 0.0380882
R50268 ASIG5V.n6130 ASIG5V.n6129 0.0380882
R50269 ASIG5V.n6130 ASIG5V.n6039 0.0380882
R50270 ASIG5V.n6137 ASIG5V.n6039 0.0380882
R50271 ASIG5V.n6138 ASIG5V.n6137 0.0380882
R50272 ASIG5V.n6139 ASIG5V.n6138 0.0380882
R50273 ASIG5V.n6139 ASIG5V.n6036 0.0380882
R50274 ASIG5V.n6146 ASIG5V.n6036 0.0380882
R50275 ASIG5V.n6147 ASIG5V.n6146 0.0380882
R50276 ASIG5V.n6148 ASIG5V.n6147 0.0380882
R50277 ASIG5V.n6148 ASIG5V.n6033 0.0380882
R50278 ASIG5V.n6155 ASIG5V.n6033 0.0380882
R50279 ASIG5V.n6156 ASIG5V.n6155 0.0380882
R50280 ASIG5V.n6157 ASIG5V.n6156 0.0380882
R50281 ASIG5V.n6157 ASIG5V.n6030 0.0380882
R50282 ASIG5V.n6164 ASIG5V.n6030 0.0380882
R50283 ASIG5V.n6165 ASIG5V.n6164 0.0380882
R50284 ASIG5V.n6166 ASIG5V.n6165 0.0380882
R50285 ASIG5V.n6166 ASIG5V.n6027 0.0380882
R50286 ASIG5V.n6173 ASIG5V.n6027 0.0380882
R50287 ASIG5V.n6174 ASIG5V.n6173 0.0380882
R50288 ASIG5V.n6175 ASIG5V.n6174 0.0380882
R50289 ASIG5V.n6175 ASIG5V.n6024 0.0380882
R50290 ASIG5V.n6182 ASIG5V.n6024 0.0380882
R50291 ASIG5V.n6183 ASIG5V.n6182 0.0380882
R50292 ASIG5V.n6184 ASIG5V.n6183 0.0380882
R50293 ASIG5V.n6184 ASIG5V.n6021 0.0380882
R50294 ASIG5V.n6191 ASIG5V.n6021 0.0380882
R50295 ASIG5V.n6192 ASIG5V.n6191 0.0380882
R50296 ASIG5V.n6193 ASIG5V.n6192 0.0380882
R50297 ASIG5V.n6193 ASIG5V.n6018 0.0380882
R50298 ASIG5V.n6200 ASIG5V.n6018 0.0380882
R50299 ASIG5V.n6201 ASIG5V.n6200 0.0380882
R50300 ASIG5V.n6202 ASIG5V.n6201 0.0380882
R50301 ASIG5V.n6202 ASIG5V.n6015 0.0380882
R50302 ASIG5V.n6209 ASIG5V.n6015 0.0380882
R50303 ASIG5V.n6210 ASIG5V.n6209 0.0380882
R50304 ASIG5V.n6211 ASIG5V.n6210 0.0380882
R50305 ASIG5V.n6211 ASIG5V.n6012 0.0380882
R50306 ASIG5V.n6218 ASIG5V.n6012 0.0380882
R50307 ASIG5V.n6219 ASIG5V.n6218 0.0380882
R50308 ASIG5V.n6220 ASIG5V.n6219 0.0380882
R50309 ASIG5V.n6220 ASIG5V.n6009 0.0380882
R50310 ASIG5V.n6227 ASIG5V.n6009 0.0380882
R50311 ASIG5V.n6228 ASIG5V.n6227 0.0380882
R50312 ASIG5V.n6229 ASIG5V.n6228 0.0380882
R50313 ASIG5V.n6229 ASIG5V.n6006 0.0380882
R50314 ASIG5V.n6236 ASIG5V.n6006 0.0380882
R50315 ASIG5V.n6237 ASIG5V.n6236 0.0380882
R50316 ASIG5V.n6238 ASIG5V.n6237 0.0380882
R50317 ASIG5V.n6238 ASIG5V.n6003 0.0380882
R50318 ASIG5V.n6245 ASIG5V.n6003 0.0380882
R50319 ASIG5V.n6246 ASIG5V.n6245 0.0380882
R50320 ASIG5V.n6247 ASIG5V.n6246 0.0380882
R50321 ASIG5V.n6064 ASIG5V.n5956 0.0380882
R50322 ASIG5V.n6064 ASIG5V.n6062 0.0380882
R50323 ASIG5V.n6069 ASIG5V.n6062 0.0380882
R50324 ASIG5V.n6071 ASIG5V.n6069 0.0380882
R50325 ASIG5V.n6073 ASIG5V.n6071 0.0380882
R50326 ASIG5V.n6073 ASIG5V.n6059 0.0380882
R50327 ASIG5V.n6078 ASIG5V.n6059 0.0380882
R50328 ASIG5V.n6080 ASIG5V.n6078 0.0380882
R50329 ASIG5V.n6082 ASIG5V.n6080 0.0380882
R50330 ASIG5V.n6082 ASIG5V.n6056 0.0380882
R50331 ASIG5V.n6087 ASIG5V.n6056 0.0380882
R50332 ASIG5V.n6089 ASIG5V.n6087 0.0380882
R50333 ASIG5V.n6091 ASIG5V.n6089 0.0380882
R50334 ASIG5V.n6091 ASIG5V.n6053 0.0380882
R50335 ASIG5V.n6096 ASIG5V.n6053 0.0380882
R50336 ASIG5V.n6098 ASIG5V.n6096 0.0380882
R50337 ASIG5V.n6100 ASIG5V.n6098 0.0380882
R50338 ASIG5V.n6100 ASIG5V.n6050 0.0380882
R50339 ASIG5V.n6105 ASIG5V.n6050 0.0380882
R50340 ASIG5V.n6107 ASIG5V.n6105 0.0380882
R50341 ASIG5V.n6109 ASIG5V.n6107 0.0380882
R50342 ASIG5V.n6109 ASIG5V.n6047 0.0380882
R50343 ASIG5V.n6114 ASIG5V.n6047 0.0380882
R50344 ASIG5V.n6116 ASIG5V.n6114 0.0380882
R50345 ASIG5V.n6118 ASIG5V.n6116 0.0380882
R50346 ASIG5V.n6118 ASIG5V.n6044 0.0380882
R50347 ASIG5V.n6123 ASIG5V.n6044 0.0380882
R50348 ASIG5V.n6125 ASIG5V.n6123 0.0380882
R50349 ASIG5V.n6127 ASIG5V.n6125 0.0380882
R50350 ASIG5V.n6127 ASIG5V.n6041 0.0380882
R50351 ASIG5V.n6132 ASIG5V.n6041 0.0380882
R50352 ASIG5V.n6134 ASIG5V.n6132 0.0380882
R50353 ASIG5V.n6136 ASIG5V.n6134 0.0380882
R50354 ASIG5V.n6136 ASIG5V.n6038 0.0380882
R50355 ASIG5V.n6141 ASIG5V.n6038 0.0380882
R50356 ASIG5V.n6143 ASIG5V.n6141 0.0380882
R50357 ASIG5V.n6145 ASIG5V.n6143 0.0380882
R50358 ASIG5V.n6145 ASIG5V.n6035 0.0380882
R50359 ASIG5V.n6150 ASIG5V.n6035 0.0380882
R50360 ASIG5V.n6152 ASIG5V.n6150 0.0380882
R50361 ASIG5V.n6154 ASIG5V.n6152 0.0380882
R50362 ASIG5V.n6154 ASIG5V.n6032 0.0380882
R50363 ASIG5V.n6159 ASIG5V.n6032 0.0380882
R50364 ASIG5V.n6161 ASIG5V.n6159 0.0380882
R50365 ASIG5V.n6163 ASIG5V.n6161 0.0380882
R50366 ASIG5V.n6163 ASIG5V.n6029 0.0380882
R50367 ASIG5V.n6168 ASIG5V.n6029 0.0380882
R50368 ASIG5V.n6170 ASIG5V.n6168 0.0380882
R50369 ASIG5V.n6172 ASIG5V.n6170 0.0380882
R50370 ASIG5V.n6172 ASIG5V.n6026 0.0380882
R50371 ASIG5V.n6177 ASIG5V.n6026 0.0380882
R50372 ASIG5V.n6179 ASIG5V.n6177 0.0380882
R50373 ASIG5V.n6181 ASIG5V.n6179 0.0380882
R50374 ASIG5V.n6181 ASIG5V.n6023 0.0380882
R50375 ASIG5V.n6186 ASIG5V.n6023 0.0380882
R50376 ASIG5V.n6188 ASIG5V.n6186 0.0380882
R50377 ASIG5V.n6190 ASIG5V.n6188 0.0380882
R50378 ASIG5V.n6190 ASIG5V.n6020 0.0380882
R50379 ASIG5V.n6195 ASIG5V.n6020 0.0380882
R50380 ASIG5V.n6197 ASIG5V.n6195 0.0380882
R50381 ASIG5V.n6199 ASIG5V.n6197 0.0380882
R50382 ASIG5V.n6199 ASIG5V.n6017 0.0380882
R50383 ASIG5V.n6204 ASIG5V.n6017 0.0380882
R50384 ASIG5V.n6206 ASIG5V.n6204 0.0380882
R50385 ASIG5V.n6208 ASIG5V.n6206 0.0380882
R50386 ASIG5V.n6208 ASIG5V.n6014 0.0380882
R50387 ASIG5V.n6213 ASIG5V.n6014 0.0380882
R50388 ASIG5V.n6215 ASIG5V.n6213 0.0380882
R50389 ASIG5V.n6217 ASIG5V.n6215 0.0380882
R50390 ASIG5V.n6217 ASIG5V.n6011 0.0380882
R50391 ASIG5V.n6222 ASIG5V.n6011 0.0380882
R50392 ASIG5V.n6224 ASIG5V.n6222 0.0380882
R50393 ASIG5V.n6226 ASIG5V.n6224 0.0380882
R50394 ASIG5V.n6226 ASIG5V.n6008 0.0380882
R50395 ASIG5V.n6231 ASIG5V.n6008 0.0380882
R50396 ASIG5V.n6233 ASIG5V.n6231 0.0380882
R50397 ASIG5V.n6235 ASIG5V.n6233 0.0380882
R50398 ASIG5V.n6235 ASIG5V.n6005 0.0380882
R50399 ASIG5V.n6240 ASIG5V.n6005 0.0380882
R50400 ASIG5V.n6242 ASIG5V.n6240 0.0380882
R50401 ASIG5V.n6244 ASIG5V.n6242 0.0380882
R50402 ASIG5V.n6244 ASIG5V.n6002 0.0380882
R50403 ASIG5V.n9391 ASIG5V.n6002 0.0380882
R50404 ASIG5V.n9194 ASIG5V.n9192 0.0380882
R50405 ASIG5V.n9195 ASIG5V.n9194 0.0380882
R50406 ASIG5V.n9196 ASIG5V.n9195 0.0380882
R50407 ASIG5V.n9196 ASIG5V.n6412 0.0380882
R50408 ASIG5V.n9203 ASIG5V.n6412 0.0380882
R50409 ASIG5V.n9204 ASIG5V.n9203 0.0380882
R50410 ASIG5V.n9205 ASIG5V.n9204 0.0380882
R50411 ASIG5V.n9205 ASIG5V.n6409 0.0380882
R50412 ASIG5V.n9212 ASIG5V.n6409 0.0380882
R50413 ASIG5V.n9213 ASIG5V.n9212 0.0380882
R50414 ASIG5V.n9214 ASIG5V.n9213 0.0380882
R50415 ASIG5V.n9214 ASIG5V.n6406 0.0380882
R50416 ASIG5V.n9221 ASIG5V.n6406 0.0380882
R50417 ASIG5V.n9222 ASIG5V.n9221 0.0380882
R50418 ASIG5V.n9223 ASIG5V.n9222 0.0380882
R50419 ASIG5V.n9223 ASIG5V.n6403 0.0380882
R50420 ASIG5V.n9230 ASIG5V.n6403 0.0380882
R50421 ASIG5V.n9231 ASIG5V.n9230 0.0380882
R50422 ASIG5V.n9232 ASIG5V.n9231 0.0380882
R50423 ASIG5V.n9232 ASIG5V.n6400 0.0380882
R50424 ASIG5V.n9239 ASIG5V.n6400 0.0380882
R50425 ASIG5V.n9240 ASIG5V.n9239 0.0380882
R50426 ASIG5V.n9241 ASIG5V.n9240 0.0380882
R50427 ASIG5V.n9241 ASIG5V.n6397 0.0380882
R50428 ASIG5V.n9248 ASIG5V.n6397 0.0380882
R50429 ASIG5V.n9249 ASIG5V.n9248 0.0380882
R50430 ASIG5V.n9250 ASIG5V.n9249 0.0380882
R50431 ASIG5V.n9250 ASIG5V.n6394 0.0380882
R50432 ASIG5V.n9257 ASIG5V.n6394 0.0380882
R50433 ASIG5V.n9258 ASIG5V.n9257 0.0380882
R50434 ASIG5V.n9259 ASIG5V.n9258 0.0380882
R50435 ASIG5V.n9259 ASIG5V.n6391 0.0380882
R50436 ASIG5V.n9266 ASIG5V.n6391 0.0380882
R50437 ASIG5V.n9267 ASIG5V.n9266 0.0380882
R50438 ASIG5V.n9268 ASIG5V.n9267 0.0380882
R50439 ASIG5V.n9268 ASIG5V.n6388 0.0380882
R50440 ASIG5V.n9275 ASIG5V.n6388 0.0380882
R50441 ASIG5V.n9276 ASIG5V.n9275 0.0380882
R50442 ASIG5V.n9277 ASIG5V.n9276 0.0380882
R50443 ASIG5V.n9277 ASIG5V.n6385 0.0380882
R50444 ASIG5V.n9284 ASIG5V.n6385 0.0380882
R50445 ASIG5V.n9285 ASIG5V.n9284 0.0380882
R50446 ASIG5V.n9286 ASIG5V.n9285 0.0380882
R50447 ASIG5V.n9286 ASIG5V.n6382 0.0380882
R50448 ASIG5V.n9293 ASIG5V.n6382 0.0380882
R50449 ASIG5V.n9294 ASIG5V.n9293 0.0380882
R50450 ASIG5V.n9295 ASIG5V.n9294 0.0380882
R50451 ASIG5V.n9295 ASIG5V.n6379 0.0380882
R50452 ASIG5V.n9302 ASIG5V.n6379 0.0380882
R50453 ASIG5V.n9303 ASIG5V.n9302 0.0380882
R50454 ASIG5V.n9304 ASIG5V.n9303 0.0380882
R50455 ASIG5V.n9304 ASIG5V.n6376 0.0380882
R50456 ASIG5V.n9311 ASIG5V.n6376 0.0380882
R50457 ASIG5V.n9312 ASIG5V.n9311 0.0380882
R50458 ASIG5V.n9313 ASIG5V.n9312 0.0380882
R50459 ASIG5V.n9313 ASIG5V.n6373 0.0380882
R50460 ASIG5V.n9320 ASIG5V.n6373 0.0380882
R50461 ASIG5V.n9321 ASIG5V.n9320 0.0380882
R50462 ASIG5V.n9322 ASIG5V.n9321 0.0380882
R50463 ASIG5V.n9322 ASIG5V.n6370 0.0380882
R50464 ASIG5V.n9329 ASIG5V.n6370 0.0380882
R50465 ASIG5V.n9330 ASIG5V.n9329 0.0380882
R50466 ASIG5V.n9331 ASIG5V.n9330 0.0380882
R50467 ASIG5V.n9331 ASIG5V.n6367 0.0380882
R50468 ASIG5V.n9338 ASIG5V.n6367 0.0380882
R50469 ASIG5V.n9339 ASIG5V.n9338 0.0380882
R50470 ASIG5V.n9340 ASIG5V.n9339 0.0380882
R50471 ASIG5V.n9340 ASIG5V.n6364 0.0380882
R50472 ASIG5V.n9347 ASIG5V.n6364 0.0380882
R50473 ASIG5V.n9348 ASIG5V.n9347 0.0380882
R50474 ASIG5V.n9349 ASIG5V.n9348 0.0380882
R50475 ASIG5V.n9349 ASIG5V.n6361 0.0380882
R50476 ASIG5V.n9356 ASIG5V.n6361 0.0380882
R50477 ASIG5V.n9357 ASIG5V.n9356 0.0380882
R50478 ASIG5V.n9358 ASIG5V.n9357 0.0380882
R50479 ASIG5V.n9358 ASIG5V.n6358 0.0380882
R50480 ASIG5V.n9365 ASIG5V.n6358 0.0380882
R50481 ASIG5V.n9366 ASIG5V.n9365 0.0380882
R50482 ASIG5V.n9367 ASIG5V.n9366 0.0380882
R50483 ASIG5V.n9367 ASIG5V.n6355 0.0380882
R50484 ASIG5V.n9374 ASIG5V.n6355 0.0380882
R50485 ASIG5V.n9375 ASIG5V.n9374 0.0380882
R50486 ASIG5V.n9376 ASIG5V.n9375 0.0380882
R50487 ASIG5V.n9193 ASIG5V.n6309 0.0380882
R50488 ASIG5V.n9193 ASIG5V.n6414 0.0380882
R50489 ASIG5V.n9198 ASIG5V.n6414 0.0380882
R50490 ASIG5V.n9200 ASIG5V.n9198 0.0380882
R50491 ASIG5V.n9202 ASIG5V.n9200 0.0380882
R50492 ASIG5V.n9202 ASIG5V.n6411 0.0380882
R50493 ASIG5V.n9207 ASIG5V.n6411 0.0380882
R50494 ASIG5V.n9209 ASIG5V.n9207 0.0380882
R50495 ASIG5V.n9211 ASIG5V.n9209 0.0380882
R50496 ASIG5V.n9211 ASIG5V.n6408 0.0380882
R50497 ASIG5V.n9216 ASIG5V.n6408 0.0380882
R50498 ASIG5V.n9218 ASIG5V.n9216 0.0380882
R50499 ASIG5V.n9220 ASIG5V.n9218 0.0380882
R50500 ASIG5V.n9220 ASIG5V.n6405 0.0380882
R50501 ASIG5V.n9225 ASIG5V.n6405 0.0380882
R50502 ASIG5V.n9227 ASIG5V.n9225 0.0380882
R50503 ASIG5V.n9229 ASIG5V.n9227 0.0380882
R50504 ASIG5V.n9229 ASIG5V.n6402 0.0380882
R50505 ASIG5V.n9234 ASIG5V.n6402 0.0380882
R50506 ASIG5V.n9236 ASIG5V.n9234 0.0380882
R50507 ASIG5V.n9238 ASIG5V.n9236 0.0380882
R50508 ASIG5V.n9238 ASIG5V.n6399 0.0380882
R50509 ASIG5V.n9243 ASIG5V.n6399 0.0380882
R50510 ASIG5V.n9245 ASIG5V.n9243 0.0380882
R50511 ASIG5V.n9247 ASIG5V.n9245 0.0380882
R50512 ASIG5V.n9247 ASIG5V.n6396 0.0380882
R50513 ASIG5V.n9252 ASIG5V.n6396 0.0380882
R50514 ASIG5V.n9254 ASIG5V.n9252 0.0380882
R50515 ASIG5V.n9256 ASIG5V.n9254 0.0380882
R50516 ASIG5V.n9256 ASIG5V.n6393 0.0380882
R50517 ASIG5V.n9261 ASIG5V.n6393 0.0380882
R50518 ASIG5V.n9263 ASIG5V.n9261 0.0380882
R50519 ASIG5V.n9265 ASIG5V.n9263 0.0380882
R50520 ASIG5V.n9265 ASIG5V.n6390 0.0380882
R50521 ASIG5V.n9270 ASIG5V.n6390 0.0380882
R50522 ASIG5V.n9272 ASIG5V.n9270 0.0380882
R50523 ASIG5V.n9274 ASIG5V.n9272 0.0380882
R50524 ASIG5V.n9274 ASIG5V.n6387 0.0380882
R50525 ASIG5V.n9279 ASIG5V.n6387 0.0380882
R50526 ASIG5V.n9281 ASIG5V.n9279 0.0380882
R50527 ASIG5V.n9283 ASIG5V.n9281 0.0380882
R50528 ASIG5V.n9283 ASIG5V.n6384 0.0380882
R50529 ASIG5V.n9288 ASIG5V.n6384 0.0380882
R50530 ASIG5V.n9290 ASIG5V.n9288 0.0380882
R50531 ASIG5V.n9292 ASIG5V.n9290 0.0380882
R50532 ASIG5V.n9292 ASIG5V.n6381 0.0380882
R50533 ASIG5V.n9297 ASIG5V.n6381 0.0380882
R50534 ASIG5V.n9299 ASIG5V.n9297 0.0380882
R50535 ASIG5V.n9301 ASIG5V.n9299 0.0380882
R50536 ASIG5V.n9301 ASIG5V.n6378 0.0380882
R50537 ASIG5V.n9306 ASIG5V.n6378 0.0380882
R50538 ASIG5V.n9308 ASIG5V.n9306 0.0380882
R50539 ASIG5V.n9310 ASIG5V.n9308 0.0380882
R50540 ASIG5V.n9310 ASIG5V.n6375 0.0380882
R50541 ASIG5V.n9315 ASIG5V.n6375 0.0380882
R50542 ASIG5V.n9317 ASIG5V.n9315 0.0380882
R50543 ASIG5V.n9319 ASIG5V.n9317 0.0380882
R50544 ASIG5V.n9319 ASIG5V.n6372 0.0380882
R50545 ASIG5V.n9324 ASIG5V.n6372 0.0380882
R50546 ASIG5V.n9326 ASIG5V.n9324 0.0380882
R50547 ASIG5V.n9328 ASIG5V.n9326 0.0380882
R50548 ASIG5V.n9328 ASIG5V.n6369 0.0380882
R50549 ASIG5V.n9333 ASIG5V.n6369 0.0380882
R50550 ASIG5V.n9335 ASIG5V.n9333 0.0380882
R50551 ASIG5V.n9337 ASIG5V.n9335 0.0380882
R50552 ASIG5V.n9337 ASIG5V.n6366 0.0380882
R50553 ASIG5V.n9342 ASIG5V.n6366 0.0380882
R50554 ASIG5V.n9344 ASIG5V.n9342 0.0380882
R50555 ASIG5V.n9346 ASIG5V.n9344 0.0380882
R50556 ASIG5V.n9346 ASIG5V.n6363 0.0380882
R50557 ASIG5V.n9351 ASIG5V.n6363 0.0380882
R50558 ASIG5V.n9353 ASIG5V.n9351 0.0380882
R50559 ASIG5V.n9355 ASIG5V.n9353 0.0380882
R50560 ASIG5V.n9355 ASIG5V.n6360 0.0380882
R50561 ASIG5V.n9360 ASIG5V.n6360 0.0380882
R50562 ASIG5V.n9362 ASIG5V.n9360 0.0380882
R50563 ASIG5V.n9364 ASIG5V.n9362 0.0380882
R50564 ASIG5V.n9364 ASIG5V.n6357 0.0380882
R50565 ASIG5V.n9369 ASIG5V.n6357 0.0380882
R50566 ASIG5V.n9371 ASIG5V.n9369 0.0380882
R50567 ASIG5V.n9373 ASIG5V.n9371 0.0380882
R50568 ASIG5V.n9373 ASIG5V.n6354 0.0380882
R50569 ASIG5V.n9377 ASIG5V.n6354 0.0380882
R50570 ASIG5V.n8930 ASIG5V.n8929 0.0380882
R50571 ASIG5V.n8931 ASIG5V.n8930 0.0380882
R50572 ASIG5V.n8931 ASIG5V.n6529 0.0380882
R50573 ASIG5V.n8941 ASIG5V.n6529 0.0380882
R50574 ASIG5V.n8942 ASIG5V.n8941 0.0380882
R50575 ASIG5V.n8943 ASIG5V.n8942 0.0380882
R50576 ASIG5V.n8943 ASIG5V.n6527 0.0380882
R50577 ASIG5V.n8953 ASIG5V.n6527 0.0380882
R50578 ASIG5V.n8954 ASIG5V.n8953 0.0380882
R50579 ASIG5V.n8955 ASIG5V.n8954 0.0380882
R50580 ASIG5V.n8955 ASIG5V.n6525 0.0380882
R50581 ASIG5V.n8965 ASIG5V.n6525 0.0380882
R50582 ASIG5V.n8966 ASIG5V.n8965 0.0380882
R50583 ASIG5V.n8967 ASIG5V.n8966 0.0380882
R50584 ASIG5V.n8967 ASIG5V.n6523 0.0380882
R50585 ASIG5V.n8977 ASIG5V.n6523 0.0380882
R50586 ASIG5V.n8978 ASIG5V.n8977 0.0380882
R50587 ASIG5V.n8979 ASIG5V.n8978 0.0380882
R50588 ASIG5V.n8979 ASIG5V.n6521 0.0380882
R50589 ASIG5V.n8989 ASIG5V.n6521 0.0380882
R50590 ASIG5V.n8990 ASIG5V.n8989 0.0380882
R50591 ASIG5V.n8991 ASIG5V.n8990 0.0380882
R50592 ASIG5V.n8991 ASIG5V.n6519 0.0380882
R50593 ASIG5V.n9001 ASIG5V.n6519 0.0380882
R50594 ASIG5V.n9002 ASIG5V.n9001 0.0380882
R50595 ASIG5V.n9003 ASIG5V.n9002 0.0380882
R50596 ASIG5V.n9003 ASIG5V.n6517 0.0380882
R50597 ASIG5V.n9013 ASIG5V.n6517 0.0380882
R50598 ASIG5V.n9014 ASIG5V.n9013 0.0380882
R50599 ASIG5V.n9015 ASIG5V.n9014 0.0380882
R50600 ASIG5V.n9015 ASIG5V.n6515 0.0380882
R50601 ASIG5V.n9025 ASIG5V.n6515 0.0380882
R50602 ASIG5V.n9026 ASIG5V.n9025 0.0380882
R50603 ASIG5V.n9027 ASIG5V.n9026 0.0380882
R50604 ASIG5V.n9027 ASIG5V.n6513 0.0380882
R50605 ASIG5V.n9037 ASIG5V.n6513 0.0380882
R50606 ASIG5V.n9038 ASIG5V.n9037 0.0380882
R50607 ASIG5V.n9039 ASIG5V.n9038 0.0380882
R50608 ASIG5V.n9039 ASIG5V.n6511 0.0380882
R50609 ASIG5V.n9049 ASIG5V.n6511 0.0380882
R50610 ASIG5V.n9050 ASIG5V.n9049 0.0380882
R50611 ASIG5V.n9051 ASIG5V.n9050 0.0380882
R50612 ASIG5V.n9051 ASIG5V.n6509 0.0380882
R50613 ASIG5V.n9061 ASIG5V.n6509 0.0380882
R50614 ASIG5V.n9062 ASIG5V.n9061 0.0380882
R50615 ASIG5V.n9063 ASIG5V.n9062 0.0380882
R50616 ASIG5V.n9063 ASIG5V.n6507 0.0380882
R50617 ASIG5V.n9073 ASIG5V.n6507 0.0380882
R50618 ASIG5V.n9074 ASIG5V.n9073 0.0380882
R50619 ASIG5V.n9075 ASIG5V.n9074 0.0380882
R50620 ASIG5V.n9075 ASIG5V.n6505 0.0380882
R50621 ASIG5V.n9085 ASIG5V.n6505 0.0380882
R50622 ASIG5V.n9086 ASIG5V.n9085 0.0380882
R50623 ASIG5V.n9087 ASIG5V.n9086 0.0380882
R50624 ASIG5V.n9087 ASIG5V.n6503 0.0380882
R50625 ASIG5V.n9097 ASIG5V.n6503 0.0380882
R50626 ASIG5V.n9098 ASIG5V.n9097 0.0380882
R50627 ASIG5V.n9099 ASIG5V.n9098 0.0380882
R50628 ASIG5V.n9099 ASIG5V.n6501 0.0380882
R50629 ASIG5V.n9109 ASIG5V.n6501 0.0380882
R50630 ASIG5V.n9110 ASIG5V.n9109 0.0380882
R50631 ASIG5V.n9111 ASIG5V.n9110 0.0380882
R50632 ASIG5V.n9111 ASIG5V.n6499 0.0380882
R50633 ASIG5V.n9121 ASIG5V.n6499 0.0380882
R50634 ASIG5V.n9122 ASIG5V.n9121 0.0380882
R50635 ASIG5V.n9123 ASIG5V.n9122 0.0380882
R50636 ASIG5V.n9123 ASIG5V.n6497 0.0380882
R50637 ASIG5V.n9133 ASIG5V.n6497 0.0380882
R50638 ASIG5V.n9134 ASIG5V.n9133 0.0380882
R50639 ASIG5V.n9135 ASIG5V.n9134 0.0380882
R50640 ASIG5V.n9135 ASIG5V.n6495 0.0380882
R50641 ASIG5V.n9145 ASIG5V.n6495 0.0380882
R50642 ASIG5V.n9146 ASIG5V.n9145 0.0380882
R50643 ASIG5V.n9147 ASIG5V.n9146 0.0380882
R50644 ASIG5V.n9147 ASIG5V.n6493 0.0380882
R50645 ASIG5V.n9157 ASIG5V.n6493 0.0380882
R50646 ASIG5V.n9158 ASIG5V.n9157 0.0380882
R50647 ASIG5V.n9159 ASIG5V.n9158 0.0380882
R50648 ASIG5V.n9159 ASIG5V.n6491 0.0380882
R50649 ASIG5V.n9169 ASIG5V.n6491 0.0380882
R50650 ASIG5V.n9170 ASIG5V.n9169 0.0380882
R50651 ASIG5V.n9171 ASIG5V.n9170 0.0380882
R50652 ASIG5V.n9171 ASIG5V.n6441 0.0380882
R50653 ASIG5V.n8928 ASIG5V.n6532 0.0380882
R50654 ASIG5V.n8932 ASIG5V.n6532 0.0380882
R50655 ASIG5V.n8936 ASIG5V.n8932 0.0380882
R50656 ASIG5V.n8940 ASIG5V.n8936 0.0380882
R50657 ASIG5V.n8940 ASIG5V.n6528 0.0380882
R50658 ASIG5V.n8944 ASIG5V.n6528 0.0380882
R50659 ASIG5V.n8948 ASIG5V.n8944 0.0380882
R50660 ASIG5V.n8952 ASIG5V.n8948 0.0380882
R50661 ASIG5V.n8952 ASIG5V.n6526 0.0380882
R50662 ASIG5V.n8956 ASIG5V.n6526 0.0380882
R50663 ASIG5V.n8960 ASIG5V.n8956 0.0380882
R50664 ASIG5V.n8964 ASIG5V.n8960 0.0380882
R50665 ASIG5V.n8964 ASIG5V.n6524 0.0380882
R50666 ASIG5V.n8968 ASIG5V.n6524 0.0380882
R50667 ASIG5V.n8972 ASIG5V.n8968 0.0380882
R50668 ASIG5V.n8976 ASIG5V.n8972 0.0380882
R50669 ASIG5V.n8976 ASIG5V.n6522 0.0380882
R50670 ASIG5V.n8980 ASIG5V.n6522 0.0380882
R50671 ASIG5V.n8984 ASIG5V.n8980 0.0380882
R50672 ASIG5V.n8988 ASIG5V.n8984 0.0380882
R50673 ASIG5V.n8988 ASIG5V.n6520 0.0380882
R50674 ASIG5V.n8992 ASIG5V.n6520 0.0380882
R50675 ASIG5V.n8996 ASIG5V.n8992 0.0380882
R50676 ASIG5V.n9000 ASIG5V.n8996 0.0380882
R50677 ASIG5V.n9000 ASIG5V.n6518 0.0380882
R50678 ASIG5V.n9004 ASIG5V.n6518 0.0380882
R50679 ASIG5V.n9008 ASIG5V.n9004 0.0380882
R50680 ASIG5V.n9012 ASIG5V.n9008 0.0380882
R50681 ASIG5V.n9012 ASIG5V.n6516 0.0380882
R50682 ASIG5V.n9016 ASIG5V.n6516 0.0380882
R50683 ASIG5V.n9020 ASIG5V.n9016 0.0380882
R50684 ASIG5V.n9024 ASIG5V.n9020 0.0380882
R50685 ASIG5V.n9024 ASIG5V.n6514 0.0380882
R50686 ASIG5V.n9028 ASIG5V.n6514 0.0380882
R50687 ASIG5V.n9032 ASIG5V.n9028 0.0380882
R50688 ASIG5V.n9036 ASIG5V.n9032 0.0380882
R50689 ASIG5V.n9036 ASIG5V.n6512 0.0380882
R50690 ASIG5V.n9040 ASIG5V.n6512 0.0380882
R50691 ASIG5V.n9044 ASIG5V.n9040 0.0380882
R50692 ASIG5V.n9048 ASIG5V.n9044 0.0380882
R50693 ASIG5V.n9048 ASIG5V.n6510 0.0380882
R50694 ASIG5V.n9052 ASIG5V.n6510 0.0380882
R50695 ASIG5V.n9056 ASIG5V.n9052 0.0380882
R50696 ASIG5V.n9060 ASIG5V.n9056 0.0380882
R50697 ASIG5V.n9060 ASIG5V.n6508 0.0380882
R50698 ASIG5V.n9064 ASIG5V.n6508 0.0380882
R50699 ASIG5V.n9068 ASIG5V.n9064 0.0380882
R50700 ASIG5V.n9072 ASIG5V.n9068 0.0380882
R50701 ASIG5V.n9072 ASIG5V.n6506 0.0380882
R50702 ASIG5V.n9076 ASIG5V.n6506 0.0380882
R50703 ASIG5V.n9080 ASIG5V.n9076 0.0380882
R50704 ASIG5V.n9084 ASIG5V.n9080 0.0380882
R50705 ASIG5V.n9084 ASIG5V.n6504 0.0380882
R50706 ASIG5V.n9088 ASIG5V.n6504 0.0380882
R50707 ASIG5V.n9092 ASIG5V.n9088 0.0380882
R50708 ASIG5V.n9096 ASIG5V.n9092 0.0380882
R50709 ASIG5V.n9096 ASIG5V.n6502 0.0380882
R50710 ASIG5V.n9100 ASIG5V.n6502 0.0380882
R50711 ASIG5V.n9104 ASIG5V.n9100 0.0380882
R50712 ASIG5V.n9108 ASIG5V.n9104 0.0380882
R50713 ASIG5V.n9108 ASIG5V.n6500 0.0380882
R50714 ASIG5V.n9112 ASIG5V.n6500 0.0380882
R50715 ASIG5V.n9116 ASIG5V.n9112 0.0380882
R50716 ASIG5V.n9120 ASIG5V.n9116 0.0380882
R50717 ASIG5V.n9120 ASIG5V.n6498 0.0380882
R50718 ASIG5V.n9124 ASIG5V.n6498 0.0380882
R50719 ASIG5V.n9128 ASIG5V.n9124 0.0380882
R50720 ASIG5V.n9132 ASIG5V.n9128 0.0380882
R50721 ASIG5V.n9132 ASIG5V.n6496 0.0380882
R50722 ASIG5V.n9136 ASIG5V.n6496 0.0380882
R50723 ASIG5V.n9140 ASIG5V.n9136 0.0380882
R50724 ASIG5V.n9144 ASIG5V.n9140 0.0380882
R50725 ASIG5V.n9144 ASIG5V.n6494 0.0380882
R50726 ASIG5V.n9148 ASIG5V.n6494 0.0380882
R50727 ASIG5V.n9152 ASIG5V.n9148 0.0380882
R50728 ASIG5V.n9156 ASIG5V.n9152 0.0380882
R50729 ASIG5V.n9156 ASIG5V.n6492 0.0380882
R50730 ASIG5V.n9160 ASIG5V.n6492 0.0380882
R50731 ASIG5V.n9164 ASIG5V.n9160 0.0380882
R50732 ASIG5V.n9168 ASIG5V.n9164 0.0380882
R50733 ASIG5V.n9168 ASIG5V.n6490 0.0380882
R50734 ASIG5V.n9172 ASIG5V.n6490 0.0380882
R50735 ASIG5V.n9172 ASIG5V.n6489 0.0380882
R50736 ASIG5V.n6698 ASIG5V.n6696 0.0380882
R50737 ASIG5V.n6699 ASIG5V.n6698 0.0380882
R50738 ASIG5V.n6700 ASIG5V.n6699 0.0380882
R50739 ASIG5V.n6700 ASIG5V.n6693 0.0380882
R50740 ASIG5V.n6707 ASIG5V.n6693 0.0380882
R50741 ASIG5V.n6708 ASIG5V.n6707 0.0380882
R50742 ASIG5V.n6709 ASIG5V.n6708 0.0380882
R50743 ASIG5V.n6709 ASIG5V.n6690 0.0380882
R50744 ASIG5V.n6716 ASIG5V.n6690 0.0380882
R50745 ASIG5V.n6717 ASIG5V.n6716 0.0380882
R50746 ASIG5V.n6718 ASIG5V.n6717 0.0380882
R50747 ASIG5V.n6718 ASIG5V.n6687 0.0380882
R50748 ASIG5V.n6725 ASIG5V.n6687 0.0380882
R50749 ASIG5V.n6726 ASIG5V.n6725 0.0380882
R50750 ASIG5V.n6727 ASIG5V.n6726 0.0380882
R50751 ASIG5V.n6727 ASIG5V.n6684 0.0380882
R50752 ASIG5V.n6734 ASIG5V.n6684 0.0380882
R50753 ASIG5V.n6735 ASIG5V.n6734 0.0380882
R50754 ASIG5V.n6736 ASIG5V.n6735 0.0380882
R50755 ASIG5V.n6736 ASIG5V.n6681 0.0380882
R50756 ASIG5V.n6743 ASIG5V.n6681 0.0380882
R50757 ASIG5V.n6744 ASIG5V.n6743 0.0380882
R50758 ASIG5V.n6745 ASIG5V.n6744 0.0380882
R50759 ASIG5V.n6745 ASIG5V.n6678 0.0380882
R50760 ASIG5V.n6752 ASIG5V.n6678 0.0380882
R50761 ASIG5V.n6753 ASIG5V.n6752 0.0380882
R50762 ASIG5V.n6754 ASIG5V.n6753 0.0380882
R50763 ASIG5V.n6754 ASIG5V.n6675 0.0380882
R50764 ASIG5V.n6761 ASIG5V.n6675 0.0380882
R50765 ASIG5V.n6762 ASIG5V.n6761 0.0380882
R50766 ASIG5V.n6763 ASIG5V.n6762 0.0380882
R50767 ASIG5V.n6763 ASIG5V.n6672 0.0380882
R50768 ASIG5V.n6770 ASIG5V.n6672 0.0380882
R50769 ASIG5V.n6771 ASIG5V.n6770 0.0380882
R50770 ASIG5V.n6772 ASIG5V.n6771 0.0380882
R50771 ASIG5V.n6772 ASIG5V.n6669 0.0380882
R50772 ASIG5V.n6779 ASIG5V.n6669 0.0380882
R50773 ASIG5V.n6780 ASIG5V.n6779 0.0380882
R50774 ASIG5V.n6781 ASIG5V.n6780 0.0380882
R50775 ASIG5V.n6781 ASIG5V.n6666 0.0380882
R50776 ASIG5V.n6788 ASIG5V.n6666 0.0380882
R50777 ASIG5V.n6789 ASIG5V.n6788 0.0380882
R50778 ASIG5V.n6790 ASIG5V.n6789 0.0380882
R50779 ASIG5V.n6790 ASIG5V.n6663 0.0380882
R50780 ASIG5V.n6797 ASIG5V.n6663 0.0380882
R50781 ASIG5V.n6798 ASIG5V.n6797 0.0380882
R50782 ASIG5V.n6799 ASIG5V.n6798 0.0380882
R50783 ASIG5V.n6799 ASIG5V.n6660 0.0380882
R50784 ASIG5V.n6806 ASIG5V.n6660 0.0380882
R50785 ASIG5V.n6807 ASIG5V.n6806 0.0380882
R50786 ASIG5V.n6808 ASIG5V.n6807 0.0380882
R50787 ASIG5V.n6808 ASIG5V.n6657 0.0380882
R50788 ASIG5V.n6815 ASIG5V.n6657 0.0380882
R50789 ASIG5V.n6816 ASIG5V.n6815 0.0380882
R50790 ASIG5V.n6817 ASIG5V.n6816 0.0380882
R50791 ASIG5V.n6817 ASIG5V.n6654 0.0380882
R50792 ASIG5V.n6824 ASIG5V.n6654 0.0380882
R50793 ASIG5V.n6825 ASIG5V.n6824 0.0380882
R50794 ASIG5V.n6826 ASIG5V.n6825 0.0380882
R50795 ASIG5V.n6826 ASIG5V.n6651 0.0380882
R50796 ASIG5V.n6833 ASIG5V.n6651 0.0380882
R50797 ASIG5V.n6834 ASIG5V.n6833 0.0380882
R50798 ASIG5V.n6835 ASIG5V.n6834 0.0380882
R50799 ASIG5V.n6835 ASIG5V.n6648 0.0380882
R50800 ASIG5V.n6842 ASIG5V.n6648 0.0380882
R50801 ASIG5V.n6843 ASIG5V.n6842 0.0380882
R50802 ASIG5V.n6844 ASIG5V.n6843 0.0380882
R50803 ASIG5V.n6844 ASIG5V.n6645 0.0380882
R50804 ASIG5V.n6851 ASIG5V.n6645 0.0380882
R50805 ASIG5V.n6852 ASIG5V.n6851 0.0380882
R50806 ASIG5V.n6853 ASIG5V.n6852 0.0380882
R50807 ASIG5V.n6853 ASIG5V.n6642 0.0380882
R50808 ASIG5V.n6860 ASIG5V.n6642 0.0380882
R50809 ASIG5V.n6861 ASIG5V.n6860 0.0380882
R50810 ASIG5V.n6862 ASIG5V.n6861 0.0380882
R50811 ASIG5V.n6862 ASIG5V.n6639 0.0380882
R50812 ASIG5V.n6869 ASIG5V.n6639 0.0380882
R50813 ASIG5V.n6870 ASIG5V.n6869 0.0380882
R50814 ASIG5V.n6871 ASIG5V.n6870 0.0380882
R50815 ASIG5V.n6871 ASIG5V.n6636 0.0380882
R50816 ASIG5V.n6878 ASIG5V.n6636 0.0380882
R50817 ASIG5V.n6879 ASIG5V.n6878 0.0380882
R50818 ASIG5V.n6880 ASIG5V.n6879 0.0380882
R50819 ASIG5V.n6697 ASIG5V.n6589 0.0380882
R50820 ASIG5V.n6697 ASIG5V.n6695 0.0380882
R50821 ASIG5V.n6702 ASIG5V.n6695 0.0380882
R50822 ASIG5V.n6704 ASIG5V.n6702 0.0380882
R50823 ASIG5V.n6706 ASIG5V.n6704 0.0380882
R50824 ASIG5V.n6706 ASIG5V.n6692 0.0380882
R50825 ASIG5V.n6711 ASIG5V.n6692 0.0380882
R50826 ASIG5V.n6713 ASIG5V.n6711 0.0380882
R50827 ASIG5V.n6715 ASIG5V.n6713 0.0380882
R50828 ASIG5V.n6715 ASIG5V.n6689 0.0380882
R50829 ASIG5V.n6720 ASIG5V.n6689 0.0380882
R50830 ASIG5V.n6722 ASIG5V.n6720 0.0380882
R50831 ASIG5V.n6724 ASIG5V.n6722 0.0380882
R50832 ASIG5V.n6724 ASIG5V.n6686 0.0380882
R50833 ASIG5V.n6729 ASIG5V.n6686 0.0380882
R50834 ASIG5V.n6731 ASIG5V.n6729 0.0380882
R50835 ASIG5V.n6733 ASIG5V.n6731 0.0380882
R50836 ASIG5V.n6733 ASIG5V.n6683 0.0380882
R50837 ASIG5V.n6738 ASIG5V.n6683 0.0380882
R50838 ASIG5V.n6740 ASIG5V.n6738 0.0380882
R50839 ASIG5V.n6742 ASIG5V.n6740 0.0380882
R50840 ASIG5V.n6742 ASIG5V.n6680 0.0380882
R50841 ASIG5V.n6747 ASIG5V.n6680 0.0380882
R50842 ASIG5V.n6749 ASIG5V.n6747 0.0380882
R50843 ASIG5V.n6751 ASIG5V.n6749 0.0380882
R50844 ASIG5V.n6751 ASIG5V.n6677 0.0380882
R50845 ASIG5V.n6756 ASIG5V.n6677 0.0380882
R50846 ASIG5V.n6758 ASIG5V.n6756 0.0380882
R50847 ASIG5V.n6760 ASIG5V.n6758 0.0380882
R50848 ASIG5V.n6760 ASIG5V.n6674 0.0380882
R50849 ASIG5V.n6765 ASIG5V.n6674 0.0380882
R50850 ASIG5V.n6767 ASIG5V.n6765 0.0380882
R50851 ASIG5V.n6769 ASIG5V.n6767 0.0380882
R50852 ASIG5V.n6769 ASIG5V.n6671 0.0380882
R50853 ASIG5V.n6774 ASIG5V.n6671 0.0380882
R50854 ASIG5V.n6776 ASIG5V.n6774 0.0380882
R50855 ASIG5V.n6778 ASIG5V.n6776 0.0380882
R50856 ASIG5V.n6778 ASIG5V.n6668 0.0380882
R50857 ASIG5V.n6783 ASIG5V.n6668 0.0380882
R50858 ASIG5V.n6785 ASIG5V.n6783 0.0380882
R50859 ASIG5V.n6787 ASIG5V.n6785 0.0380882
R50860 ASIG5V.n6787 ASIG5V.n6665 0.0380882
R50861 ASIG5V.n6792 ASIG5V.n6665 0.0380882
R50862 ASIG5V.n6794 ASIG5V.n6792 0.0380882
R50863 ASIG5V.n6796 ASIG5V.n6794 0.0380882
R50864 ASIG5V.n6796 ASIG5V.n6662 0.0380882
R50865 ASIG5V.n6801 ASIG5V.n6662 0.0380882
R50866 ASIG5V.n6803 ASIG5V.n6801 0.0380882
R50867 ASIG5V.n6805 ASIG5V.n6803 0.0380882
R50868 ASIG5V.n6805 ASIG5V.n6659 0.0380882
R50869 ASIG5V.n6810 ASIG5V.n6659 0.0380882
R50870 ASIG5V.n6812 ASIG5V.n6810 0.0380882
R50871 ASIG5V.n6814 ASIG5V.n6812 0.0380882
R50872 ASIG5V.n6814 ASIG5V.n6656 0.0380882
R50873 ASIG5V.n6819 ASIG5V.n6656 0.0380882
R50874 ASIG5V.n6821 ASIG5V.n6819 0.0380882
R50875 ASIG5V.n6823 ASIG5V.n6821 0.0380882
R50876 ASIG5V.n6823 ASIG5V.n6653 0.0380882
R50877 ASIG5V.n6828 ASIG5V.n6653 0.0380882
R50878 ASIG5V.n6830 ASIG5V.n6828 0.0380882
R50879 ASIG5V.n6832 ASIG5V.n6830 0.0380882
R50880 ASIG5V.n6832 ASIG5V.n6650 0.0380882
R50881 ASIG5V.n6837 ASIG5V.n6650 0.0380882
R50882 ASIG5V.n6839 ASIG5V.n6837 0.0380882
R50883 ASIG5V.n6841 ASIG5V.n6839 0.0380882
R50884 ASIG5V.n6841 ASIG5V.n6647 0.0380882
R50885 ASIG5V.n6846 ASIG5V.n6647 0.0380882
R50886 ASIG5V.n6848 ASIG5V.n6846 0.0380882
R50887 ASIG5V.n6850 ASIG5V.n6848 0.0380882
R50888 ASIG5V.n6850 ASIG5V.n6644 0.0380882
R50889 ASIG5V.n6855 ASIG5V.n6644 0.0380882
R50890 ASIG5V.n6857 ASIG5V.n6855 0.0380882
R50891 ASIG5V.n6859 ASIG5V.n6857 0.0380882
R50892 ASIG5V.n6859 ASIG5V.n6641 0.0380882
R50893 ASIG5V.n6864 ASIG5V.n6641 0.0380882
R50894 ASIG5V.n6866 ASIG5V.n6864 0.0380882
R50895 ASIG5V.n6868 ASIG5V.n6866 0.0380882
R50896 ASIG5V.n6868 ASIG5V.n6638 0.0380882
R50897 ASIG5V.n6873 ASIG5V.n6638 0.0380882
R50898 ASIG5V.n6875 ASIG5V.n6873 0.0380882
R50899 ASIG5V.n6877 ASIG5V.n6875 0.0380882
R50900 ASIG5V.n6877 ASIG5V.n6635 0.0380882
R50901 ASIG5V.n8914 ASIG5V.n6635 0.0380882
R50902 ASIG5V.n7231 ASIG5V.n6897 0.0380882
R50903 ASIG5V.n7223 ASIG5V.n6897 0.0380882
R50904 ASIG5V.n7223 ASIG5V.n7222 0.0380882
R50905 ASIG5V.n7222 ASIG5V.n7221 0.0380882
R50906 ASIG5V.n7221 ASIG5V.n6901 0.0380882
R50907 ASIG5V.n7213 ASIG5V.n6901 0.0380882
R50908 ASIG5V.n7213 ASIG5V.n7212 0.0380882
R50909 ASIG5V.n7212 ASIG5V.n7211 0.0380882
R50910 ASIG5V.n7211 ASIG5V.n6907 0.0380882
R50911 ASIG5V.n7203 ASIG5V.n6907 0.0380882
R50912 ASIG5V.n7203 ASIG5V.n7202 0.0380882
R50913 ASIG5V.n7202 ASIG5V.n7201 0.0380882
R50914 ASIG5V.n7201 ASIG5V.n6913 0.0380882
R50915 ASIG5V.n7193 ASIG5V.n6913 0.0380882
R50916 ASIG5V.n7193 ASIG5V.n7192 0.0380882
R50917 ASIG5V.n7192 ASIG5V.n7191 0.0380882
R50918 ASIG5V.n7191 ASIG5V.n6919 0.0380882
R50919 ASIG5V.n7183 ASIG5V.n6919 0.0380882
R50920 ASIG5V.n7183 ASIG5V.n7182 0.0380882
R50921 ASIG5V.n7182 ASIG5V.n7181 0.0380882
R50922 ASIG5V.n7181 ASIG5V.n6925 0.0380882
R50923 ASIG5V.n7173 ASIG5V.n6925 0.0380882
R50924 ASIG5V.n7173 ASIG5V.n7172 0.0380882
R50925 ASIG5V.n7172 ASIG5V.n7171 0.0380882
R50926 ASIG5V.n7171 ASIG5V.n6931 0.0380882
R50927 ASIG5V.n7163 ASIG5V.n6931 0.0380882
R50928 ASIG5V.n7163 ASIG5V.n7162 0.0380882
R50929 ASIG5V.n7162 ASIG5V.n7161 0.0380882
R50930 ASIG5V.n7161 ASIG5V.n6937 0.0380882
R50931 ASIG5V.n7153 ASIG5V.n6937 0.0380882
R50932 ASIG5V.n7153 ASIG5V.n7152 0.0380882
R50933 ASIG5V.n7152 ASIG5V.n7151 0.0380882
R50934 ASIG5V.n7151 ASIG5V.n6943 0.0380882
R50935 ASIG5V.n7143 ASIG5V.n6943 0.0380882
R50936 ASIG5V.n7143 ASIG5V.n7142 0.0380882
R50937 ASIG5V.n7142 ASIG5V.n7141 0.0380882
R50938 ASIG5V.n7141 ASIG5V.n6949 0.0380882
R50939 ASIG5V.n7133 ASIG5V.n6949 0.0380882
R50940 ASIG5V.n7133 ASIG5V.n7132 0.0380882
R50941 ASIG5V.n7132 ASIG5V.n7131 0.0380882
R50942 ASIG5V.n7131 ASIG5V.n6955 0.0380882
R50943 ASIG5V.n7123 ASIG5V.n6955 0.0380882
R50944 ASIG5V.n7123 ASIG5V.n7122 0.0380882
R50945 ASIG5V.n7122 ASIG5V.n7121 0.0380882
R50946 ASIG5V.n7121 ASIG5V.n6961 0.0380882
R50947 ASIG5V.n7113 ASIG5V.n6961 0.0380882
R50948 ASIG5V.n7113 ASIG5V.n7112 0.0380882
R50949 ASIG5V.n7112 ASIG5V.n7111 0.0380882
R50950 ASIG5V.n7111 ASIG5V.n6967 0.0380882
R50951 ASIG5V.n7103 ASIG5V.n6967 0.0380882
R50952 ASIG5V.n7103 ASIG5V.n7102 0.0380882
R50953 ASIG5V.n7102 ASIG5V.n7101 0.0380882
R50954 ASIG5V.n7101 ASIG5V.n6973 0.0380882
R50955 ASIG5V.n7093 ASIG5V.n6973 0.0380882
R50956 ASIG5V.n7093 ASIG5V.n7092 0.0380882
R50957 ASIG5V.n7092 ASIG5V.n7091 0.0380882
R50958 ASIG5V.n7091 ASIG5V.n6979 0.0380882
R50959 ASIG5V.n7083 ASIG5V.n6979 0.0380882
R50960 ASIG5V.n7083 ASIG5V.n7082 0.0380882
R50961 ASIG5V.n7082 ASIG5V.n7081 0.0380882
R50962 ASIG5V.n7081 ASIG5V.n6985 0.0380882
R50963 ASIG5V.n7073 ASIG5V.n6985 0.0380882
R50964 ASIG5V.n7073 ASIG5V.n7072 0.0380882
R50965 ASIG5V.n7072 ASIG5V.n7071 0.0380882
R50966 ASIG5V.n7071 ASIG5V.n6991 0.0380882
R50967 ASIG5V.n7063 ASIG5V.n6991 0.0380882
R50968 ASIG5V.n7063 ASIG5V.n7062 0.0380882
R50969 ASIG5V.n7062 ASIG5V.n7061 0.0380882
R50970 ASIG5V.n7061 ASIG5V.n6997 0.0380882
R50971 ASIG5V.n7053 ASIG5V.n6997 0.0380882
R50972 ASIG5V.n7053 ASIG5V.n7052 0.0380882
R50973 ASIG5V.n7052 ASIG5V.n7051 0.0380882
R50974 ASIG5V.n7051 ASIG5V.n7003 0.0380882
R50975 ASIG5V.n7043 ASIG5V.n7003 0.0380882
R50976 ASIG5V.n7043 ASIG5V.n7042 0.0380882
R50977 ASIG5V.n7042 ASIG5V.n7041 0.0380882
R50978 ASIG5V.n7041 ASIG5V.n7009 0.0380882
R50979 ASIG5V.n7033 ASIG5V.n7009 0.0380882
R50980 ASIG5V.n7033 ASIG5V.n7032 0.0380882
R50981 ASIG5V.n7032 ASIG5V.n7031 0.0380882
R50982 ASIG5V.n7031 ASIG5V.n7015 0.0380882
R50983 ASIG5V.n7023 ASIG5V.n7015 0.0380882
R50984 ASIG5V.n7023 ASIG5V.n7022 0.0380882
R50985 ASIG5V.n7230 ASIG5V.n6898 0.0380882
R50986 ASIG5V.n7224 ASIG5V.n6898 0.0380882
R50987 ASIG5V.n7224 ASIG5V.n6900 0.0380882
R50988 ASIG5V.n7220 ASIG5V.n6900 0.0380882
R50989 ASIG5V.n7220 ASIG5V.n6902 0.0380882
R50990 ASIG5V.n7214 ASIG5V.n6902 0.0380882
R50991 ASIG5V.n7214 ASIG5V.n6906 0.0380882
R50992 ASIG5V.n7210 ASIG5V.n6906 0.0380882
R50993 ASIG5V.n7210 ASIG5V.n6908 0.0380882
R50994 ASIG5V.n7204 ASIG5V.n6908 0.0380882
R50995 ASIG5V.n7204 ASIG5V.n6912 0.0380882
R50996 ASIG5V.n7200 ASIG5V.n6912 0.0380882
R50997 ASIG5V.n7200 ASIG5V.n6914 0.0380882
R50998 ASIG5V.n7194 ASIG5V.n6914 0.0380882
R50999 ASIG5V.n7194 ASIG5V.n6918 0.0380882
R51000 ASIG5V.n7190 ASIG5V.n6918 0.0380882
R51001 ASIG5V.n7190 ASIG5V.n6920 0.0380882
R51002 ASIG5V.n7184 ASIG5V.n6920 0.0380882
R51003 ASIG5V.n7184 ASIG5V.n6924 0.0380882
R51004 ASIG5V.n7180 ASIG5V.n6924 0.0380882
R51005 ASIG5V.n7180 ASIG5V.n6926 0.0380882
R51006 ASIG5V.n7174 ASIG5V.n6926 0.0380882
R51007 ASIG5V.n7174 ASIG5V.n6930 0.0380882
R51008 ASIG5V.n7170 ASIG5V.n6930 0.0380882
R51009 ASIG5V.n7170 ASIG5V.n6932 0.0380882
R51010 ASIG5V.n7164 ASIG5V.n6932 0.0380882
R51011 ASIG5V.n7164 ASIG5V.n6936 0.0380882
R51012 ASIG5V.n7160 ASIG5V.n6936 0.0380882
R51013 ASIG5V.n7160 ASIG5V.n6938 0.0380882
R51014 ASIG5V.n7154 ASIG5V.n6938 0.0380882
R51015 ASIG5V.n7154 ASIG5V.n6942 0.0380882
R51016 ASIG5V.n7150 ASIG5V.n6942 0.0380882
R51017 ASIG5V.n7150 ASIG5V.n6944 0.0380882
R51018 ASIG5V.n7144 ASIG5V.n6944 0.0380882
R51019 ASIG5V.n7144 ASIG5V.n6948 0.0380882
R51020 ASIG5V.n7140 ASIG5V.n6948 0.0380882
R51021 ASIG5V.n7140 ASIG5V.n6950 0.0380882
R51022 ASIG5V.n7134 ASIG5V.n6950 0.0380882
R51023 ASIG5V.n7134 ASIG5V.n6954 0.0380882
R51024 ASIG5V.n7130 ASIG5V.n6954 0.0380882
R51025 ASIG5V.n7130 ASIG5V.n6956 0.0380882
R51026 ASIG5V.n7124 ASIG5V.n6956 0.0380882
R51027 ASIG5V.n7124 ASIG5V.n6960 0.0380882
R51028 ASIG5V.n7120 ASIG5V.n6960 0.0380882
R51029 ASIG5V.n7120 ASIG5V.n6962 0.0380882
R51030 ASIG5V.n7114 ASIG5V.n6962 0.0380882
R51031 ASIG5V.n7114 ASIG5V.n6966 0.0380882
R51032 ASIG5V.n7110 ASIG5V.n6966 0.0380882
R51033 ASIG5V.n7110 ASIG5V.n6968 0.0380882
R51034 ASIG5V.n7104 ASIG5V.n6968 0.0380882
R51035 ASIG5V.n7104 ASIG5V.n6972 0.0380882
R51036 ASIG5V.n7100 ASIG5V.n6972 0.0380882
R51037 ASIG5V.n7100 ASIG5V.n6974 0.0380882
R51038 ASIG5V.n7094 ASIG5V.n6974 0.0380882
R51039 ASIG5V.n7094 ASIG5V.n6978 0.0380882
R51040 ASIG5V.n7090 ASIG5V.n6978 0.0380882
R51041 ASIG5V.n7090 ASIG5V.n6980 0.0380882
R51042 ASIG5V.n7084 ASIG5V.n6980 0.0380882
R51043 ASIG5V.n7084 ASIG5V.n6984 0.0380882
R51044 ASIG5V.n7080 ASIG5V.n6984 0.0380882
R51045 ASIG5V.n7080 ASIG5V.n6986 0.0380882
R51046 ASIG5V.n7074 ASIG5V.n6986 0.0380882
R51047 ASIG5V.n7074 ASIG5V.n6990 0.0380882
R51048 ASIG5V.n7070 ASIG5V.n6990 0.0380882
R51049 ASIG5V.n7070 ASIG5V.n6992 0.0380882
R51050 ASIG5V.n7064 ASIG5V.n6992 0.0380882
R51051 ASIG5V.n7064 ASIG5V.n6996 0.0380882
R51052 ASIG5V.n7060 ASIG5V.n6996 0.0380882
R51053 ASIG5V.n7060 ASIG5V.n6998 0.0380882
R51054 ASIG5V.n7054 ASIG5V.n6998 0.0380882
R51055 ASIG5V.n7054 ASIG5V.n7002 0.0380882
R51056 ASIG5V.n7050 ASIG5V.n7002 0.0380882
R51057 ASIG5V.n7050 ASIG5V.n7004 0.0380882
R51058 ASIG5V.n7044 ASIG5V.n7004 0.0380882
R51059 ASIG5V.n7044 ASIG5V.n7008 0.0380882
R51060 ASIG5V.n7040 ASIG5V.n7008 0.0380882
R51061 ASIG5V.n7040 ASIG5V.n7010 0.0380882
R51062 ASIG5V.n7034 ASIG5V.n7010 0.0380882
R51063 ASIG5V.n7034 ASIG5V.n7014 0.0380882
R51064 ASIG5V.n7030 ASIG5V.n7014 0.0380882
R51065 ASIG5V.n7030 ASIG5V.n7016 0.0380882
R51066 ASIG5V.n7024 ASIG5V.n7016 0.0380882
R51067 ASIG5V.n7024 ASIG5V.n7021 0.0380882
R51068 ASIG5V.n8568 ASIG5V.n8567 0.0380882
R51069 ASIG5V.n8567 ASIG5V.n8325 0.0380882
R51070 ASIG5V.n8561 ASIG5V.n8325 0.0380882
R51071 ASIG5V.n8561 ASIG5V.n8560 0.0380882
R51072 ASIG5V.n8560 ASIG5V.n8559 0.0380882
R51073 ASIG5V.n8559 ASIG5V.n8328 0.0380882
R51074 ASIG5V.n8552 ASIG5V.n8328 0.0380882
R51075 ASIG5V.n8552 ASIG5V.n8551 0.0380882
R51076 ASIG5V.n8551 ASIG5V.n8550 0.0380882
R51077 ASIG5V.n8550 ASIG5V.n8331 0.0380882
R51078 ASIG5V.n8543 ASIG5V.n8331 0.0380882
R51079 ASIG5V.n8543 ASIG5V.n8542 0.0380882
R51080 ASIG5V.n8542 ASIG5V.n8541 0.0380882
R51081 ASIG5V.n8541 ASIG5V.n8334 0.0380882
R51082 ASIG5V.n8534 ASIG5V.n8334 0.0380882
R51083 ASIG5V.n8534 ASIG5V.n8533 0.0380882
R51084 ASIG5V.n8533 ASIG5V.n8532 0.0380882
R51085 ASIG5V.n8532 ASIG5V.n8337 0.0380882
R51086 ASIG5V.n8525 ASIG5V.n8337 0.0380882
R51087 ASIG5V.n8525 ASIG5V.n8524 0.0380882
R51088 ASIG5V.n8524 ASIG5V.n8523 0.0380882
R51089 ASIG5V.n8523 ASIG5V.n8340 0.0380882
R51090 ASIG5V.n8516 ASIG5V.n8340 0.0380882
R51091 ASIG5V.n8516 ASIG5V.n8515 0.0380882
R51092 ASIG5V.n8515 ASIG5V.n8514 0.0380882
R51093 ASIG5V.n8514 ASIG5V.n8343 0.0380882
R51094 ASIG5V.n8507 ASIG5V.n8343 0.0380882
R51095 ASIG5V.n8507 ASIG5V.n8506 0.0380882
R51096 ASIG5V.n8506 ASIG5V.n8505 0.0380882
R51097 ASIG5V.n8505 ASIG5V.n8346 0.0380882
R51098 ASIG5V.n8498 ASIG5V.n8346 0.0380882
R51099 ASIG5V.n8498 ASIG5V.n8497 0.0380882
R51100 ASIG5V.n8497 ASIG5V.n8496 0.0380882
R51101 ASIG5V.n8496 ASIG5V.n8349 0.0380882
R51102 ASIG5V.n8489 ASIG5V.n8349 0.0380882
R51103 ASIG5V.n8489 ASIG5V.n8488 0.0380882
R51104 ASIG5V.n8488 ASIG5V.n8487 0.0380882
R51105 ASIG5V.n8487 ASIG5V.n8352 0.0380882
R51106 ASIG5V.n8480 ASIG5V.n8352 0.0380882
R51107 ASIG5V.n8480 ASIG5V.n8479 0.0380882
R51108 ASIG5V.n8479 ASIG5V.n8478 0.0380882
R51109 ASIG5V.n8478 ASIG5V.n8355 0.0380882
R51110 ASIG5V.n8471 ASIG5V.n8355 0.0380882
R51111 ASIG5V.n8471 ASIG5V.n8470 0.0380882
R51112 ASIG5V.n8470 ASIG5V.n8469 0.0380882
R51113 ASIG5V.n8469 ASIG5V.n8358 0.0380882
R51114 ASIG5V.n8462 ASIG5V.n8358 0.0380882
R51115 ASIG5V.n8462 ASIG5V.n8461 0.0380882
R51116 ASIG5V.n8461 ASIG5V.n8460 0.0380882
R51117 ASIG5V.n8460 ASIG5V.n8361 0.0380882
R51118 ASIG5V.n8453 ASIG5V.n8361 0.0380882
R51119 ASIG5V.n8453 ASIG5V.n8452 0.0380882
R51120 ASIG5V.n8452 ASIG5V.n8451 0.0380882
R51121 ASIG5V.n8451 ASIG5V.n8364 0.0380882
R51122 ASIG5V.n8444 ASIG5V.n8364 0.0380882
R51123 ASIG5V.n8444 ASIG5V.n8443 0.0380882
R51124 ASIG5V.n8443 ASIG5V.n8442 0.0380882
R51125 ASIG5V.n8442 ASIG5V.n8367 0.0380882
R51126 ASIG5V.n8435 ASIG5V.n8367 0.0380882
R51127 ASIG5V.n8435 ASIG5V.n8434 0.0380882
R51128 ASIG5V.n8434 ASIG5V.n8433 0.0380882
R51129 ASIG5V.n8433 ASIG5V.n8370 0.0380882
R51130 ASIG5V.n8426 ASIG5V.n8370 0.0380882
R51131 ASIG5V.n8426 ASIG5V.n8425 0.0380882
R51132 ASIG5V.n8425 ASIG5V.n8424 0.0380882
R51133 ASIG5V.n8424 ASIG5V.n8373 0.0380882
R51134 ASIG5V.n8417 ASIG5V.n8373 0.0380882
R51135 ASIG5V.n8417 ASIG5V.n8416 0.0380882
R51136 ASIG5V.n8416 ASIG5V.n8415 0.0380882
R51137 ASIG5V.n8415 ASIG5V.n8376 0.0380882
R51138 ASIG5V.n8408 ASIG5V.n8376 0.0380882
R51139 ASIG5V.n8408 ASIG5V.n8407 0.0380882
R51140 ASIG5V.n8407 ASIG5V.n8406 0.0380882
R51141 ASIG5V.n8406 ASIG5V.n8379 0.0380882
R51142 ASIG5V.n8399 ASIG5V.n8379 0.0380882
R51143 ASIG5V.n8399 ASIG5V.n8398 0.0380882
R51144 ASIG5V.n8398 ASIG5V.n8397 0.0380882
R51145 ASIG5V.n8397 ASIG5V.n8382 0.0380882
R51146 ASIG5V.n8390 ASIG5V.n8382 0.0380882
R51147 ASIG5V.n8390 ASIG5V.n8389 0.0380882
R51148 ASIG5V.n8389 ASIG5V.n8388 0.0380882
R51149 ASIG5V.n8388 ASIG5V.n8385 0.0380882
R51150 ASIG5V.n8385 ASIG5V.n8263 0.0380882
R51151 ASIG5V.n8566 ASIG5V.n8216 0.0380882
R51152 ASIG5V.n8566 ASIG5V.n8565 0.0380882
R51153 ASIG5V.n8565 ASIG5V.n8563 0.0380882
R51154 ASIG5V.n8563 ASIG5V.n8327 0.0380882
R51155 ASIG5V.n8558 ASIG5V.n8327 0.0380882
R51156 ASIG5V.n8558 ASIG5V.n8556 0.0380882
R51157 ASIG5V.n8556 ASIG5V.n8554 0.0380882
R51158 ASIG5V.n8554 ASIG5V.n8330 0.0380882
R51159 ASIG5V.n8549 ASIG5V.n8330 0.0380882
R51160 ASIG5V.n8549 ASIG5V.n8547 0.0380882
R51161 ASIG5V.n8547 ASIG5V.n8545 0.0380882
R51162 ASIG5V.n8545 ASIG5V.n8333 0.0380882
R51163 ASIG5V.n8540 ASIG5V.n8333 0.0380882
R51164 ASIG5V.n8540 ASIG5V.n8538 0.0380882
R51165 ASIG5V.n8538 ASIG5V.n8536 0.0380882
R51166 ASIG5V.n8536 ASIG5V.n8336 0.0380882
R51167 ASIG5V.n8531 ASIG5V.n8336 0.0380882
R51168 ASIG5V.n8531 ASIG5V.n8529 0.0380882
R51169 ASIG5V.n8529 ASIG5V.n8527 0.0380882
R51170 ASIG5V.n8527 ASIG5V.n8339 0.0380882
R51171 ASIG5V.n8522 ASIG5V.n8339 0.0380882
R51172 ASIG5V.n8522 ASIG5V.n8520 0.0380882
R51173 ASIG5V.n8520 ASIG5V.n8518 0.0380882
R51174 ASIG5V.n8518 ASIG5V.n8342 0.0380882
R51175 ASIG5V.n8513 ASIG5V.n8342 0.0380882
R51176 ASIG5V.n8513 ASIG5V.n8511 0.0380882
R51177 ASIG5V.n8511 ASIG5V.n8509 0.0380882
R51178 ASIG5V.n8509 ASIG5V.n8345 0.0380882
R51179 ASIG5V.n8504 ASIG5V.n8345 0.0380882
R51180 ASIG5V.n8504 ASIG5V.n8502 0.0380882
R51181 ASIG5V.n8502 ASIG5V.n8500 0.0380882
R51182 ASIG5V.n8500 ASIG5V.n8348 0.0380882
R51183 ASIG5V.n8495 ASIG5V.n8348 0.0380882
R51184 ASIG5V.n8495 ASIG5V.n8493 0.0380882
R51185 ASIG5V.n8493 ASIG5V.n8491 0.0380882
R51186 ASIG5V.n8491 ASIG5V.n8351 0.0380882
R51187 ASIG5V.n8486 ASIG5V.n8351 0.0380882
R51188 ASIG5V.n8486 ASIG5V.n8484 0.0380882
R51189 ASIG5V.n8484 ASIG5V.n8482 0.0380882
R51190 ASIG5V.n8482 ASIG5V.n8354 0.0380882
R51191 ASIG5V.n8477 ASIG5V.n8354 0.0380882
R51192 ASIG5V.n8477 ASIG5V.n8475 0.0380882
R51193 ASIG5V.n8475 ASIG5V.n8473 0.0380882
R51194 ASIG5V.n8473 ASIG5V.n8357 0.0380882
R51195 ASIG5V.n8468 ASIG5V.n8357 0.0380882
R51196 ASIG5V.n8468 ASIG5V.n8466 0.0380882
R51197 ASIG5V.n8466 ASIG5V.n8464 0.0380882
R51198 ASIG5V.n8464 ASIG5V.n8360 0.0380882
R51199 ASIG5V.n8459 ASIG5V.n8360 0.0380882
R51200 ASIG5V.n8459 ASIG5V.n8457 0.0380882
R51201 ASIG5V.n8457 ASIG5V.n8455 0.0380882
R51202 ASIG5V.n8455 ASIG5V.n8363 0.0380882
R51203 ASIG5V.n8450 ASIG5V.n8363 0.0380882
R51204 ASIG5V.n8450 ASIG5V.n8448 0.0380882
R51205 ASIG5V.n8448 ASIG5V.n8446 0.0380882
R51206 ASIG5V.n8446 ASIG5V.n8366 0.0380882
R51207 ASIG5V.n8441 ASIG5V.n8366 0.0380882
R51208 ASIG5V.n8441 ASIG5V.n8439 0.0380882
R51209 ASIG5V.n8439 ASIG5V.n8437 0.0380882
R51210 ASIG5V.n8437 ASIG5V.n8369 0.0380882
R51211 ASIG5V.n8432 ASIG5V.n8369 0.0380882
R51212 ASIG5V.n8432 ASIG5V.n8430 0.0380882
R51213 ASIG5V.n8430 ASIG5V.n8428 0.0380882
R51214 ASIG5V.n8428 ASIG5V.n8372 0.0380882
R51215 ASIG5V.n8423 ASIG5V.n8372 0.0380882
R51216 ASIG5V.n8423 ASIG5V.n8421 0.0380882
R51217 ASIG5V.n8421 ASIG5V.n8419 0.0380882
R51218 ASIG5V.n8419 ASIG5V.n8375 0.0380882
R51219 ASIG5V.n8414 ASIG5V.n8375 0.0380882
R51220 ASIG5V.n8414 ASIG5V.n8412 0.0380882
R51221 ASIG5V.n8412 ASIG5V.n8410 0.0380882
R51222 ASIG5V.n8410 ASIG5V.n8378 0.0380882
R51223 ASIG5V.n8405 ASIG5V.n8378 0.0380882
R51224 ASIG5V.n8405 ASIG5V.n8403 0.0380882
R51225 ASIG5V.n8403 ASIG5V.n8401 0.0380882
R51226 ASIG5V.n8401 ASIG5V.n8381 0.0380882
R51227 ASIG5V.n8396 ASIG5V.n8381 0.0380882
R51228 ASIG5V.n8396 ASIG5V.n8394 0.0380882
R51229 ASIG5V.n8394 ASIG5V.n8392 0.0380882
R51230 ASIG5V.n8392 ASIG5V.n8384 0.0380882
R51231 ASIG5V.n8387 ASIG5V.n8384 0.0380882
R51232 ASIG5V.n8387 ASIG5V.n8262 0.0380882
R51233 ASIG5V.n8890 ASIG5V.n8262 0.0380882
R51234 ASIG5V.n8876 ASIG5V.n8588 0.0380882
R51235 ASIG5V.n8876 ASIG5V.n8875 0.0380882
R51236 ASIG5V.n8875 ASIG5V.n8874 0.0380882
R51237 ASIG5V.n8874 ASIG5V.n8592 0.0380882
R51238 ASIG5V.n8864 ASIG5V.n8592 0.0380882
R51239 ASIG5V.n8864 ASIG5V.n8863 0.0380882
R51240 ASIG5V.n8863 ASIG5V.n8862 0.0380882
R51241 ASIG5V.n8862 ASIG5V.n8594 0.0380882
R51242 ASIG5V.n8852 ASIG5V.n8594 0.0380882
R51243 ASIG5V.n8852 ASIG5V.n8851 0.0380882
R51244 ASIG5V.n8851 ASIG5V.n8850 0.0380882
R51245 ASIG5V.n8850 ASIG5V.n8596 0.0380882
R51246 ASIG5V.n8840 ASIG5V.n8596 0.0380882
R51247 ASIG5V.n8840 ASIG5V.n8839 0.0380882
R51248 ASIG5V.n8839 ASIG5V.n8838 0.0380882
R51249 ASIG5V.n8838 ASIG5V.n8598 0.0380882
R51250 ASIG5V.n8828 ASIG5V.n8598 0.0380882
R51251 ASIG5V.n8828 ASIG5V.n8827 0.0380882
R51252 ASIG5V.n8827 ASIG5V.n8826 0.0380882
R51253 ASIG5V.n8826 ASIG5V.n8600 0.0380882
R51254 ASIG5V.n8816 ASIG5V.n8600 0.0380882
R51255 ASIG5V.n8816 ASIG5V.n8815 0.0380882
R51256 ASIG5V.n8815 ASIG5V.n8814 0.0380882
R51257 ASIG5V.n8814 ASIG5V.n8602 0.0380882
R51258 ASIG5V.n8804 ASIG5V.n8602 0.0380882
R51259 ASIG5V.n8804 ASIG5V.n8803 0.0380882
R51260 ASIG5V.n8803 ASIG5V.n8802 0.0380882
R51261 ASIG5V.n8802 ASIG5V.n8604 0.0380882
R51262 ASIG5V.n8792 ASIG5V.n8604 0.0380882
R51263 ASIG5V.n8792 ASIG5V.n8791 0.0380882
R51264 ASIG5V.n8791 ASIG5V.n8790 0.0380882
R51265 ASIG5V.n8790 ASIG5V.n8606 0.0380882
R51266 ASIG5V.n8780 ASIG5V.n8606 0.0380882
R51267 ASIG5V.n8780 ASIG5V.n8779 0.0380882
R51268 ASIG5V.n8779 ASIG5V.n8778 0.0380882
R51269 ASIG5V.n8778 ASIG5V.n8608 0.0380882
R51270 ASIG5V.n8768 ASIG5V.n8608 0.0380882
R51271 ASIG5V.n8768 ASIG5V.n8767 0.0380882
R51272 ASIG5V.n8767 ASIG5V.n8766 0.0380882
R51273 ASIG5V.n8766 ASIG5V.n8610 0.0380882
R51274 ASIG5V.n8756 ASIG5V.n8610 0.0380882
R51275 ASIG5V.n8756 ASIG5V.n8755 0.0380882
R51276 ASIG5V.n8755 ASIG5V.n8754 0.0380882
R51277 ASIG5V.n8754 ASIG5V.n8612 0.0380882
R51278 ASIG5V.n8744 ASIG5V.n8612 0.0380882
R51279 ASIG5V.n8744 ASIG5V.n8743 0.0380882
R51280 ASIG5V.n8743 ASIG5V.n8742 0.0380882
R51281 ASIG5V.n8742 ASIG5V.n8614 0.0380882
R51282 ASIG5V.n8732 ASIG5V.n8614 0.0380882
R51283 ASIG5V.n8732 ASIG5V.n8731 0.0380882
R51284 ASIG5V.n8731 ASIG5V.n8730 0.0380882
R51285 ASIG5V.n8730 ASIG5V.n8616 0.0380882
R51286 ASIG5V.n8720 ASIG5V.n8616 0.0380882
R51287 ASIG5V.n8720 ASIG5V.n8719 0.0380882
R51288 ASIG5V.n8719 ASIG5V.n8718 0.0380882
R51289 ASIG5V.n8718 ASIG5V.n8618 0.0380882
R51290 ASIG5V.n8708 ASIG5V.n8618 0.0380882
R51291 ASIG5V.n8708 ASIG5V.n8707 0.0380882
R51292 ASIG5V.n8707 ASIG5V.n8706 0.0380882
R51293 ASIG5V.n8706 ASIG5V.n8620 0.0380882
R51294 ASIG5V.n8696 ASIG5V.n8620 0.0380882
R51295 ASIG5V.n8696 ASIG5V.n8695 0.0380882
R51296 ASIG5V.n8695 ASIG5V.n8694 0.0380882
R51297 ASIG5V.n8694 ASIG5V.n8622 0.0380882
R51298 ASIG5V.n8684 ASIG5V.n8622 0.0380882
R51299 ASIG5V.n8684 ASIG5V.n8683 0.0380882
R51300 ASIG5V.n8683 ASIG5V.n8682 0.0380882
R51301 ASIG5V.n8682 ASIG5V.n8624 0.0380882
R51302 ASIG5V.n8672 ASIG5V.n8624 0.0380882
R51303 ASIG5V.n8672 ASIG5V.n8671 0.0380882
R51304 ASIG5V.n8671 ASIG5V.n8670 0.0380882
R51305 ASIG5V.n8670 ASIG5V.n8626 0.0380882
R51306 ASIG5V.n8660 ASIG5V.n8626 0.0380882
R51307 ASIG5V.n8660 ASIG5V.n8659 0.0380882
R51308 ASIG5V.n8659 ASIG5V.n8658 0.0380882
R51309 ASIG5V.n8658 ASIG5V.n8628 0.0380882
R51310 ASIG5V.n8648 ASIG5V.n8628 0.0380882
R51311 ASIG5V.n8648 ASIG5V.n8647 0.0380882
R51312 ASIG5V.n8647 ASIG5V.n8646 0.0380882
R51313 ASIG5V.n8646 ASIG5V.n8630 0.0380882
R51314 ASIG5V.n8636 ASIG5V.n8630 0.0380882
R51315 ASIG5V.n8636 ASIG5V.n8635 0.0380882
R51316 ASIG5V.n8635 ASIG5V.n8634 0.0380882
R51317 ASIG5V.n8878 ASIG5V.n8877 0.0380882
R51318 ASIG5V.n8877 ASIG5V.n8591 0.0380882
R51319 ASIG5V.n8873 ASIG5V.n8591 0.0380882
R51320 ASIG5V.n8873 ASIG5V.n8869 0.0380882
R51321 ASIG5V.n8869 ASIG5V.n8868 0.0380882
R51322 ASIG5V.n8868 ASIG5V.n8593 0.0380882
R51323 ASIG5V.n8861 ASIG5V.n8593 0.0380882
R51324 ASIG5V.n8861 ASIG5V.n8857 0.0380882
R51325 ASIG5V.n8857 ASIG5V.n8856 0.0380882
R51326 ASIG5V.n8856 ASIG5V.n8595 0.0380882
R51327 ASIG5V.n8849 ASIG5V.n8595 0.0380882
R51328 ASIG5V.n8849 ASIG5V.n8845 0.0380882
R51329 ASIG5V.n8845 ASIG5V.n8844 0.0380882
R51330 ASIG5V.n8844 ASIG5V.n8597 0.0380882
R51331 ASIG5V.n8837 ASIG5V.n8597 0.0380882
R51332 ASIG5V.n8837 ASIG5V.n8833 0.0380882
R51333 ASIG5V.n8833 ASIG5V.n8832 0.0380882
R51334 ASIG5V.n8832 ASIG5V.n8599 0.0380882
R51335 ASIG5V.n8825 ASIG5V.n8599 0.0380882
R51336 ASIG5V.n8825 ASIG5V.n8821 0.0380882
R51337 ASIG5V.n8821 ASIG5V.n8820 0.0380882
R51338 ASIG5V.n8820 ASIG5V.n8601 0.0380882
R51339 ASIG5V.n8813 ASIG5V.n8601 0.0380882
R51340 ASIG5V.n8813 ASIG5V.n8809 0.0380882
R51341 ASIG5V.n8809 ASIG5V.n8808 0.0380882
R51342 ASIG5V.n8808 ASIG5V.n8603 0.0380882
R51343 ASIG5V.n8801 ASIG5V.n8603 0.0380882
R51344 ASIG5V.n8801 ASIG5V.n8797 0.0380882
R51345 ASIG5V.n8797 ASIG5V.n8796 0.0380882
R51346 ASIG5V.n8796 ASIG5V.n8605 0.0380882
R51347 ASIG5V.n8789 ASIG5V.n8605 0.0380882
R51348 ASIG5V.n8789 ASIG5V.n8785 0.0380882
R51349 ASIG5V.n8785 ASIG5V.n8784 0.0380882
R51350 ASIG5V.n8784 ASIG5V.n8607 0.0380882
R51351 ASIG5V.n8777 ASIG5V.n8607 0.0380882
R51352 ASIG5V.n8777 ASIG5V.n8773 0.0380882
R51353 ASIG5V.n8773 ASIG5V.n8772 0.0380882
R51354 ASIG5V.n8772 ASIG5V.n8609 0.0380882
R51355 ASIG5V.n8765 ASIG5V.n8609 0.0380882
R51356 ASIG5V.n8765 ASIG5V.n8761 0.0380882
R51357 ASIG5V.n8761 ASIG5V.n8760 0.0380882
R51358 ASIG5V.n8760 ASIG5V.n8611 0.0380882
R51359 ASIG5V.n8753 ASIG5V.n8611 0.0380882
R51360 ASIG5V.n8753 ASIG5V.n8749 0.0380882
R51361 ASIG5V.n8749 ASIG5V.n8748 0.0380882
R51362 ASIG5V.n8748 ASIG5V.n8613 0.0380882
R51363 ASIG5V.n8741 ASIG5V.n8613 0.0380882
R51364 ASIG5V.n8741 ASIG5V.n8737 0.0380882
R51365 ASIG5V.n8737 ASIG5V.n8736 0.0380882
R51366 ASIG5V.n8736 ASIG5V.n8615 0.0380882
R51367 ASIG5V.n8729 ASIG5V.n8615 0.0380882
R51368 ASIG5V.n8729 ASIG5V.n8725 0.0380882
R51369 ASIG5V.n8725 ASIG5V.n8724 0.0380882
R51370 ASIG5V.n8724 ASIG5V.n8617 0.0380882
R51371 ASIG5V.n8717 ASIG5V.n8617 0.0380882
R51372 ASIG5V.n8717 ASIG5V.n8713 0.0380882
R51373 ASIG5V.n8713 ASIG5V.n8712 0.0380882
R51374 ASIG5V.n8712 ASIG5V.n8619 0.0380882
R51375 ASIG5V.n8705 ASIG5V.n8619 0.0380882
R51376 ASIG5V.n8705 ASIG5V.n8701 0.0380882
R51377 ASIG5V.n8701 ASIG5V.n8700 0.0380882
R51378 ASIG5V.n8700 ASIG5V.n8621 0.0380882
R51379 ASIG5V.n8693 ASIG5V.n8621 0.0380882
R51380 ASIG5V.n8693 ASIG5V.n8689 0.0380882
R51381 ASIG5V.n8689 ASIG5V.n8688 0.0380882
R51382 ASIG5V.n8688 ASIG5V.n8623 0.0380882
R51383 ASIG5V.n8681 ASIG5V.n8623 0.0380882
R51384 ASIG5V.n8681 ASIG5V.n8677 0.0380882
R51385 ASIG5V.n8677 ASIG5V.n8676 0.0380882
R51386 ASIG5V.n8676 ASIG5V.n8625 0.0380882
R51387 ASIG5V.n8669 ASIG5V.n8625 0.0380882
R51388 ASIG5V.n8669 ASIG5V.n8665 0.0380882
R51389 ASIG5V.n8665 ASIG5V.n8664 0.0380882
R51390 ASIG5V.n8664 ASIG5V.n8627 0.0380882
R51391 ASIG5V.n8657 ASIG5V.n8627 0.0380882
R51392 ASIG5V.n8657 ASIG5V.n8653 0.0380882
R51393 ASIG5V.n8653 ASIG5V.n8652 0.0380882
R51394 ASIG5V.n8652 ASIG5V.n8629 0.0380882
R51395 ASIG5V.n8645 ASIG5V.n8629 0.0380882
R51396 ASIG5V.n8645 ASIG5V.n8641 0.0380882
R51397 ASIG5V.n8641 ASIG5V.n8640 0.0380882
R51398 ASIG5V.n8640 ASIG5V.n8631 0.0380882
R51399 ASIG5V.n8633 ASIG5V.n8631 0.0380882
R51400 ASIG5V.n12340 ASIG5V.n12338 0.0380882
R51401 ASIG5V.n12341 ASIG5V.n12340 0.0380882
R51402 ASIG5V.n12342 ASIG5V.n12341 0.0380882
R51403 ASIG5V.n12342 ASIG5V.n158 0.0380882
R51404 ASIG5V.n12349 ASIG5V.n158 0.0380882
R51405 ASIG5V.n12350 ASIG5V.n12349 0.0380882
R51406 ASIG5V.n12351 ASIG5V.n12350 0.0380882
R51407 ASIG5V.n12351 ASIG5V.n155 0.0380882
R51408 ASIG5V.n12358 ASIG5V.n155 0.0380882
R51409 ASIG5V.n12359 ASIG5V.n12358 0.0380882
R51410 ASIG5V.n12360 ASIG5V.n12359 0.0380882
R51411 ASIG5V.n12360 ASIG5V.n152 0.0380882
R51412 ASIG5V.n12367 ASIG5V.n152 0.0380882
R51413 ASIG5V.n12368 ASIG5V.n12367 0.0380882
R51414 ASIG5V.n12369 ASIG5V.n12368 0.0380882
R51415 ASIG5V.n12369 ASIG5V.n149 0.0380882
R51416 ASIG5V.n12376 ASIG5V.n149 0.0380882
R51417 ASIG5V.n12377 ASIG5V.n12376 0.0380882
R51418 ASIG5V.n12378 ASIG5V.n12377 0.0380882
R51419 ASIG5V.n12378 ASIG5V.n146 0.0380882
R51420 ASIG5V.n12385 ASIG5V.n146 0.0380882
R51421 ASIG5V.n12386 ASIG5V.n12385 0.0380882
R51422 ASIG5V.n12387 ASIG5V.n12386 0.0380882
R51423 ASIG5V.n12387 ASIG5V.n143 0.0380882
R51424 ASIG5V.n12394 ASIG5V.n143 0.0380882
R51425 ASIG5V.n12395 ASIG5V.n12394 0.0380882
R51426 ASIG5V.n12396 ASIG5V.n12395 0.0380882
R51427 ASIG5V.n12396 ASIG5V.n140 0.0380882
R51428 ASIG5V.n12403 ASIG5V.n140 0.0380882
R51429 ASIG5V.n12404 ASIG5V.n12403 0.0380882
R51430 ASIG5V.n12405 ASIG5V.n12404 0.0380882
R51431 ASIG5V.n12405 ASIG5V.n137 0.0380882
R51432 ASIG5V.n12412 ASIG5V.n137 0.0380882
R51433 ASIG5V.n12413 ASIG5V.n12412 0.0380882
R51434 ASIG5V.n12414 ASIG5V.n12413 0.0380882
R51435 ASIG5V.n12414 ASIG5V.n134 0.0380882
R51436 ASIG5V.n12421 ASIG5V.n134 0.0380882
R51437 ASIG5V.n12422 ASIG5V.n12421 0.0380882
R51438 ASIG5V.n12423 ASIG5V.n12422 0.0380882
R51439 ASIG5V.n12423 ASIG5V.n131 0.0380882
R51440 ASIG5V.n12430 ASIG5V.n131 0.0380882
R51441 ASIG5V.n12431 ASIG5V.n12430 0.0380882
R51442 ASIG5V.n12432 ASIG5V.n12431 0.0380882
R51443 ASIG5V.n12432 ASIG5V.n128 0.0380882
R51444 ASIG5V.n12439 ASIG5V.n128 0.0380882
R51445 ASIG5V.n12440 ASIG5V.n12439 0.0380882
R51446 ASIG5V.n12441 ASIG5V.n12440 0.0380882
R51447 ASIG5V.n12441 ASIG5V.n125 0.0380882
R51448 ASIG5V.n12448 ASIG5V.n125 0.0380882
R51449 ASIG5V.n12449 ASIG5V.n12448 0.0380882
R51450 ASIG5V.n12450 ASIG5V.n12449 0.0380882
R51451 ASIG5V.n12450 ASIG5V.n122 0.0380882
R51452 ASIG5V.n12457 ASIG5V.n122 0.0380882
R51453 ASIG5V.n12458 ASIG5V.n12457 0.0380882
R51454 ASIG5V.n12459 ASIG5V.n12458 0.0380882
R51455 ASIG5V.n12459 ASIG5V.n119 0.0380882
R51456 ASIG5V.n12466 ASIG5V.n119 0.0380882
R51457 ASIG5V.n12467 ASIG5V.n12466 0.0380882
R51458 ASIG5V.n12468 ASIG5V.n12467 0.0380882
R51459 ASIG5V.n12468 ASIG5V.n116 0.0380882
R51460 ASIG5V.n12475 ASIG5V.n116 0.0380882
R51461 ASIG5V.n12476 ASIG5V.n12475 0.0380882
R51462 ASIG5V.n12477 ASIG5V.n12476 0.0380882
R51463 ASIG5V.n12477 ASIG5V.n113 0.0380882
R51464 ASIG5V.n12484 ASIG5V.n113 0.0380882
R51465 ASIG5V.n12485 ASIG5V.n12484 0.0380882
R51466 ASIG5V.n12486 ASIG5V.n12485 0.0380882
R51467 ASIG5V.n12486 ASIG5V.n110 0.0380882
R51468 ASIG5V.n12493 ASIG5V.n110 0.0380882
R51469 ASIG5V.n12494 ASIG5V.n12493 0.0380882
R51470 ASIG5V.n12495 ASIG5V.n12494 0.0380882
R51471 ASIG5V.n12495 ASIG5V.n107 0.0380882
R51472 ASIG5V.n12502 ASIG5V.n107 0.0380882
R51473 ASIG5V.n12503 ASIG5V.n12502 0.0380882
R51474 ASIG5V.n12504 ASIG5V.n12503 0.0380882
R51475 ASIG5V.n12504 ASIG5V.n104 0.0380882
R51476 ASIG5V.n12511 ASIG5V.n104 0.0380882
R51477 ASIG5V.n12512 ASIG5V.n12511 0.0380882
R51478 ASIG5V.n12513 ASIG5V.n12512 0.0380882
R51479 ASIG5V.n12513 ASIG5V.n101 0.0380882
R51480 ASIG5V.n12520 ASIG5V.n101 0.0380882
R51481 ASIG5V.n12521 ASIG5V.n12520 0.0380882
R51482 ASIG5V.n12522 ASIG5V.n12521 0.0380882
R51483 ASIG5V.n12339 ASIG5V.n55 0.0380882
R51484 ASIG5V.n12339 ASIG5V.n160 0.0380882
R51485 ASIG5V.n12344 ASIG5V.n160 0.0380882
R51486 ASIG5V.n12346 ASIG5V.n12344 0.0380882
R51487 ASIG5V.n12348 ASIG5V.n12346 0.0380882
R51488 ASIG5V.n12348 ASIG5V.n157 0.0380882
R51489 ASIG5V.n12353 ASIG5V.n157 0.0380882
R51490 ASIG5V.n12355 ASIG5V.n12353 0.0380882
R51491 ASIG5V.n12357 ASIG5V.n12355 0.0380882
R51492 ASIG5V.n12357 ASIG5V.n154 0.0380882
R51493 ASIG5V.n12362 ASIG5V.n154 0.0380882
R51494 ASIG5V.n12364 ASIG5V.n12362 0.0380882
R51495 ASIG5V.n12366 ASIG5V.n12364 0.0380882
R51496 ASIG5V.n12366 ASIG5V.n151 0.0380882
R51497 ASIG5V.n12371 ASIG5V.n151 0.0380882
R51498 ASIG5V.n12373 ASIG5V.n12371 0.0380882
R51499 ASIG5V.n12375 ASIG5V.n12373 0.0380882
R51500 ASIG5V.n12375 ASIG5V.n148 0.0380882
R51501 ASIG5V.n12380 ASIG5V.n148 0.0380882
R51502 ASIG5V.n12382 ASIG5V.n12380 0.0380882
R51503 ASIG5V.n12384 ASIG5V.n12382 0.0380882
R51504 ASIG5V.n12384 ASIG5V.n145 0.0380882
R51505 ASIG5V.n12389 ASIG5V.n145 0.0380882
R51506 ASIG5V.n12391 ASIG5V.n12389 0.0380882
R51507 ASIG5V.n12393 ASIG5V.n12391 0.0380882
R51508 ASIG5V.n12393 ASIG5V.n142 0.0380882
R51509 ASIG5V.n12398 ASIG5V.n142 0.0380882
R51510 ASIG5V.n12400 ASIG5V.n12398 0.0380882
R51511 ASIG5V.n12402 ASIG5V.n12400 0.0380882
R51512 ASIG5V.n12402 ASIG5V.n139 0.0380882
R51513 ASIG5V.n12407 ASIG5V.n139 0.0380882
R51514 ASIG5V.n12409 ASIG5V.n12407 0.0380882
R51515 ASIG5V.n12411 ASIG5V.n12409 0.0380882
R51516 ASIG5V.n12411 ASIG5V.n136 0.0380882
R51517 ASIG5V.n12416 ASIG5V.n136 0.0380882
R51518 ASIG5V.n12418 ASIG5V.n12416 0.0380882
R51519 ASIG5V.n12420 ASIG5V.n12418 0.0380882
R51520 ASIG5V.n12420 ASIG5V.n133 0.0380882
R51521 ASIG5V.n12425 ASIG5V.n133 0.0380882
R51522 ASIG5V.n12427 ASIG5V.n12425 0.0380882
R51523 ASIG5V.n12429 ASIG5V.n12427 0.0380882
R51524 ASIG5V.n12429 ASIG5V.n130 0.0380882
R51525 ASIG5V.n12434 ASIG5V.n130 0.0380882
R51526 ASIG5V.n12436 ASIG5V.n12434 0.0380882
R51527 ASIG5V.n12438 ASIG5V.n12436 0.0380882
R51528 ASIG5V.n12438 ASIG5V.n127 0.0380882
R51529 ASIG5V.n12443 ASIG5V.n127 0.0380882
R51530 ASIG5V.n12445 ASIG5V.n12443 0.0380882
R51531 ASIG5V.n12447 ASIG5V.n12445 0.0380882
R51532 ASIG5V.n12447 ASIG5V.n124 0.0380882
R51533 ASIG5V.n12452 ASIG5V.n124 0.0380882
R51534 ASIG5V.n12454 ASIG5V.n12452 0.0380882
R51535 ASIG5V.n12456 ASIG5V.n12454 0.0380882
R51536 ASIG5V.n12456 ASIG5V.n121 0.0380882
R51537 ASIG5V.n12461 ASIG5V.n121 0.0380882
R51538 ASIG5V.n12463 ASIG5V.n12461 0.0380882
R51539 ASIG5V.n12465 ASIG5V.n12463 0.0380882
R51540 ASIG5V.n12465 ASIG5V.n118 0.0380882
R51541 ASIG5V.n12470 ASIG5V.n118 0.0380882
R51542 ASIG5V.n12472 ASIG5V.n12470 0.0380882
R51543 ASIG5V.n12474 ASIG5V.n12472 0.0380882
R51544 ASIG5V.n12474 ASIG5V.n115 0.0380882
R51545 ASIG5V.n12479 ASIG5V.n115 0.0380882
R51546 ASIG5V.n12481 ASIG5V.n12479 0.0380882
R51547 ASIG5V.n12483 ASIG5V.n12481 0.0380882
R51548 ASIG5V.n12483 ASIG5V.n112 0.0380882
R51549 ASIG5V.n12488 ASIG5V.n112 0.0380882
R51550 ASIG5V.n12490 ASIG5V.n12488 0.0380882
R51551 ASIG5V.n12492 ASIG5V.n12490 0.0380882
R51552 ASIG5V.n12492 ASIG5V.n109 0.0380882
R51553 ASIG5V.n12497 ASIG5V.n109 0.0380882
R51554 ASIG5V.n12499 ASIG5V.n12497 0.0380882
R51555 ASIG5V.n12501 ASIG5V.n12499 0.0380882
R51556 ASIG5V.n12501 ASIG5V.n106 0.0380882
R51557 ASIG5V.n12506 ASIG5V.n106 0.0380882
R51558 ASIG5V.n12508 ASIG5V.n12506 0.0380882
R51559 ASIG5V.n12510 ASIG5V.n12508 0.0380882
R51560 ASIG5V.n12510 ASIG5V.n103 0.0380882
R51561 ASIG5V.n12515 ASIG5V.n103 0.0380882
R51562 ASIG5V.n12517 ASIG5V.n12515 0.0380882
R51563 ASIG5V.n12519 ASIG5V.n12517 0.0380882
R51564 ASIG5V.n12519 ASIG5V.n100 0.0380882
R51565 ASIG5V.n12523 ASIG5V.n100 0.0380882
R51566 ASIG5V.n264 ASIG5V.n168 0.0380882
R51567 ASIG5V.n265 ASIG5V.n264 0.0380882
R51568 ASIG5V.n265 ASIG5V.n259 0.0380882
R51569 ASIG5V.n275 ASIG5V.n259 0.0380882
R51570 ASIG5V.n276 ASIG5V.n275 0.0380882
R51571 ASIG5V.n277 ASIG5V.n276 0.0380882
R51572 ASIG5V.n277 ASIG5V.n257 0.0380882
R51573 ASIG5V.n287 ASIG5V.n257 0.0380882
R51574 ASIG5V.n288 ASIG5V.n287 0.0380882
R51575 ASIG5V.n289 ASIG5V.n288 0.0380882
R51576 ASIG5V.n289 ASIG5V.n255 0.0380882
R51577 ASIG5V.n299 ASIG5V.n255 0.0380882
R51578 ASIG5V.n300 ASIG5V.n299 0.0380882
R51579 ASIG5V.n301 ASIG5V.n300 0.0380882
R51580 ASIG5V.n301 ASIG5V.n253 0.0380882
R51581 ASIG5V.n311 ASIG5V.n253 0.0380882
R51582 ASIG5V.n312 ASIG5V.n311 0.0380882
R51583 ASIG5V.n313 ASIG5V.n312 0.0380882
R51584 ASIG5V.n313 ASIG5V.n251 0.0380882
R51585 ASIG5V.n323 ASIG5V.n251 0.0380882
R51586 ASIG5V.n324 ASIG5V.n323 0.0380882
R51587 ASIG5V.n325 ASIG5V.n324 0.0380882
R51588 ASIG5V.n325 ASIG5V.n249 0.0380882
R51589 ASIG5V.n335 ASIG5V.n249 0.0380882
R51590 ASIG5V.n336 ASIG5V.n335 0.0380882
R51591 ASIG5V.n337 ASIG5V.n336 0.0380882
R51592 ASIG5V.n337 ASIG5V.n247 0.0380882
R51593 ASIG5V.n347 ASIG5V.n247 0.0380882
R51594 ASIG5V.n348 ASIG5V.n347 0.0380882
R51595 ASIG5V.n349 ASIG5V.n348 0.0380882
R51596 ASIG5V.n349 ASIG5V.n245 0.0380882
R51597 ASIG5V.n359 ASIG5V.n245 0.0380882
R51598 ASIG5V.n360 ASIG5V.n359 0.0380882
R51599 ASIG5V.n361 ASIG5V.n360 0.0380882
R51600 ASIG5V.n361 ASIG5V.n243 0.0380882
R51601 ASIG5V.n371 ASIG5V.n243 0.0380882
R51602 ASIG5V.n372 ASIG5V.n371 0.0380882
R51603 ASIG5V.n373 ASIG5V.n372 0.0380882
R51604 ASIG5V.n373 ASIG5V.n241 0.0380882
R51605 ASIG5V.n383 ASIG5V.n241 0.0380882
R51606 ASIG5V.n384 ASIG5V.n383 0.0380882
R51607 ASIG5V.n385 ASIG5V.n384 0.0380882
R51608 ASIG5V.n385 ASIG5V.n239 0.0380882
R51609 ASIG5V.n395 ASIG5V.n239 0.0380882
R51610 ASIG5V.n396 ASIG5V.n395 0.0380882
R51611 ASIG5V.n397 ASIG5V.n396 0.0380882
R51612 ASIG5V.n397 ASIG5V.n237 0.0380882
R51613 ASIG5V.n407 ASIG5V.n237 0.0380882
R51614 ASIG5V.n408 ASIG5V.n407 0.0380882
R51615 ASIG5V.n409 ASIG5V.n408 0.0380882
R51616 ASIG5V.n409 ASIG5V.n235 0.0380882
R51617 ASIG5V.n419 ASIG5V.n235 0.0380882
R51618 ASIG5V.n420 ASIG5V.n419 0.0380882
R51619 ASIG5V.n421 ASIG5V.n420 0.0380882
R51620 ASIG5V.n421 ASIG5V.n233 0.0380882
R51621 ASIG5V.n431 ASIG5V.n233 0.0380882
R51622 ASIG5V.n432 ASIG5V.n431 0.0380882
R51623 ASIG5V.n433 ASIG5V.n432 0.0380882
R51624 ASIG5V.n433 ASIG5V.n231 0.0380882
R51625 ASIG5V.n443 ASIG5V.n231 0.0380882
R51626 ASIG5V.n444 ASIG5V.n443 0.0380882
R51627 ASIG5V.n445 ASIG5V.n444 0.0380882
R51628 ASIG5V.n445 ASIG5V.n229 0.0380882
R51629 ASIG5V.n455 ASIG5V.n229 0.0380882
R51630 ASIG5V.n456 ASIG5V.n455 0.0380882
R51631 ASIG5V.n457 ASIG5V.n456 0.0380882
R51632 ASIG5V.n457 ASIG5V.n227 0.0380882
R51633 ASIG5V.n467 ASIG5V.n227 0.0380882
R51634 ASIG5V.n468 ASIG5V.n467 0.0380882
R51635 ASIG5V.n469 ASIG5V.n468 0.0380882
R51636 ASIG5V.n469 ASIG5V.n225 0.0380882
R51637 ASIG5V.n479 ASIG5V.n225 0.0380882
R51638 ASIG5V.n480 ASIG5V.n479 0.0380882
R51639 ASIG5V.n481 ASIG5V.n480 0.0380882
R51640 ASIG5V.n481 ASIG5V.n223 0.0380882
R51641 ASIG5V.n491 ASIG5V.n223 0.0380882
R51642 ASIG5V.n492 ASIG5V.n491 0.0380882
R51643 ASIG5V.n493 ASIG5V.n492 0.0380882
R51644 ASIG5V.n493 ASIG5V.n221 0.0380882
R51645 ASIG5V.n503 ASIG5V.n221 0.0380882
R51646 ASIG5V.n504 ASIG5V.n503 0.0380882
R51647 ASIG5V.n12318 ASIG5V.n504 0.0380882
R51648 ASIG5V.n12318 ASIG5V.n12317 0.0380882
R51649 ASIG5V.n263 ASIG5V.n260 0.0380882
R51650 ASIG5V.n266 ASIG5V.n263 0.0380882
R51651 ASIG5V.n270 ASIG5V.n266 0.0380882
R51652 ASIG5V.n274 ASIG5V.n270 0.0380882
R51653 ASIG5V.n274 ASIG5V.n258 0.0380882
R51654 ASIG5V.n278 ASIG5V.n258 0.0380882
R51655 ASIG5V.n282 ASIG5V.n278 0.0380882
R51656 ASIG5V.n286 ASIG5V.n282 0.0380882
R51657 ASIG5V.n286 ASIG5V.n256 0.0380882
R51658 ASIG5V.n290 ASIG5V.n256 0.0380882
R51659 ASIG5V.n294 ASIG5V.n290 0.0380882
R51660 ASIG5V.n298 ASIG5V.n294 0.0380882
R51661 ASIG5V.n298 ASIG5V.n254 0.0380882
R51662 ASIG5V.n302 ASIG5V.n254 0.0380882
R51663 ASIG5V.n306 ASIG5V.n302 0.0380882
R51664 ASIG5V.n310 ASIG5V.n306 0.0380882
R51665 ASIG5V.n310 ASIG5V.n252 0.0380882
R51666 ASIG5V.n314 ASIG5V.n252 0.0380882
R51667 ASIG5V.n318 ASIG5V.n314 0.0380882
R51668 ASIG5V.n322 ASIG5V.n318 0.0380882
R51669 ASIG5V.n322 ASIG5V.n250 0.0380882
R51670 ASIG5V.n326 ASIG5V.n250 0.0380882
R51671 ASIG5V.n330 ASIG5V.n326 0.0380882
R51672 ASIG5V.n334 ASIG5V.n330 0.0380882
R51673 ASIG5V.n334 ASIG5V.n248 0.0380882
R51674 ASIG5V.n338 ASIG5V.n248 0.0380882
R51675 ASIG5V.n342 ASIG5V.n338 0.0380882
R51676 ASIG5V.n346 ASIG5V.n342 0.0380882
R51677 ASIG5V.n346 ASIG5V.n246 0.0380882
R51678 ASIG5V.n350 ASIG5V.n246 0.0380882
R51679 ASIG5V.n354 ASIG5V.n350 0.0380882
R51680 ASIG5V.n358 ASIG5V.n354 0.0380882
R51681 ASIG5V.n358 ASIG5V.n244 0.0380882
R51682 ASIG5V.n362 ASIG5V.n244 0.0380882
R51683 ASIG5V.n366 ASIG5V.n362 0.0380882
R51684 ASIG5V.n370 ASIG5V.n366 0.0380882
R51685 ASIG5V.n370 ASIG5V.n242 0.0380882
R51686 ASIG5V.n374 ASIG5V.n242 0.0380882
R51687 ASIG5V.n378 ASIG5V.n374 0.0380882
R51688 ASIG5V.n382 ASIG5V.n378 0.0380882
R51689 ASIG5V.n382 ASIG5V.n240 0.0380882
R51690 ASIG5V.n386 ASIG5V.n240 0.0380882
R51691 ASIG5V.n390 ASIG5V.n386 0.0380882
R51692 ASIG5V.n394 ASIG5V.n390 0.0380882
R51693 ASIG5V.n394 ASIG5V.n238 0.0380882
R51694 ASIG5V.n398 ASIG5V.n238 0.0380882
R51695 ASIG5V.n402 ASIG5V.n398 0.0380882
R51696 ASIG5V.n406 ASIG5V.n402 0.0380882
R51697 ASIG5V.n406 ASIG5V.n236 0.0380882
R51698 ASIG5V.n410 ASIG5V.n236 0.0380882
R51699 ASIG5V.n414 ASIG5V.n410 0.0380882
R51700 ASIG5V.n418 ASIG5V.n414 0.0380882
R51701 ASIG5V.n418 ASIG5V.n234 0.0380882
R51702 ASIG5V.n422 ASIG5V.n234 0.0380882
R51703 ASIG5V.n426 ASIG5V.n422 0.0380882
R51704 ASIG5V.n430 ASIG5V.n426 0.0380882
R51705 ASIG5V.n430 ASIG5V.n232 0.0380882
R51706 ASIG5V.n434 ASIG5V.n232 0.0380882
R51707 ASIG5V.n438 ASIG5V.n434 0.0380882
R51708 ASIG5V.n442 ASIG5V.n438 0.0380882
R51709 ASIG5V.n442 ASIG5V.n230 0.0380882
R51710 ASIG5V.n446 ASIG5V.n230 0.0380882
R51711 ASIG5V.n450 ASIG5V.n446 0.0380882
R51712 ASIG5V.n454 ASIG5V.n450 0.0380882
R51713 ASIG5V.n454 ASIG5V.n228 0.0380882
R51714 ASIG5V.n458 ASIG5V.n228 0.0380882
R51715 ASIG5V.n462 ASIG5V.n458 0.0380882
R51716 ASIG5V.n466 ASIG5V.n462 0.0380882
R51717 ASIG5V.n466 ASIG5V.n226 0.0380882
R51718 ASIG5V.n470 ASIG5V.n226 0.0380882
R51719 ASIG5V.n474 ASIG5V.n470 0.0380882
R51720 ASIG5V.n478 ASIG5V.n474 0.0380882
R51721 ASIG5V.n478 ASIG5V.n224 0.0380882
R51722 ASIG5V.n482 ASIG5V.n224 0.0380882
R51723 ASIG5V.n486 ASIG5V.n482 0.0380882
R51724 ASIG5V.n490 ASIG5V.n486 0.0380882
R51725 ASIG5V.n490 ASIG5V.n222 0.0380882
R51726 ASIG5V.n494 ASIG5V.n222 0.0380882
R51727 ASIG5V.n498 ASIG5V.n494 0.0380882
R51728 ASIG5V.n502 ASIG5V.n498 0.0380882
R51729 ASIG5V.n502 ASIG5V.n220 0.0380882
R51730 ASIG5V.n12319 ASIG5V.n220 0.0380882
R51731 ASIG5V.n12319 ASIG5V.n218 0.0380882
R51732 ASIG5V.n618 ASIG5V.n524 0.0380882
R51733 ASIG5V.n619 ASIG5V.n618 0.0380882
R51734 ASIG5V.n619 ASIG5V.n613 0.0380882
R51735 ASIG5V.n629 ASIG5V.n613 0.0380882
R51736 ASIG5V.n630 ASIG5V.n629 0.0380882
R51737 ASIG5V.n631 ASIG5V.n630 0.0380882
R51738 ASIG5V.n631 ASIG5V.n611 0.0380882
R51739 ASIG5V.n641 ASIG5V.n611 0.0380882
R51740 ASIG5V.n642 ASIG5V.n641 0.0380882
R51741 ASIG5V.n643 ASIG5V.n642 0.0380882
R51742 ASIG5V.n643 ASIG5V.n609 0.0380882
R51743 ASIG5V.n653 ASIG5V.n609 0.0380882
R51744 ASIG5V.n654 ASIG5V.n653 0.0380882
R51745 ASIG5V.n655 ASIG5V.n654 0.0380882
R51746 ASIG5V.n655 ASIG5V.n607 0.0380882
R51747 ASIG5V.n665 ASIG5V.n607 0.0380882
R51748 ASIG5V.n666 ASIG5V.n665 0.0380882
R51749 ASIG5V.n667 ASIG5V.n666 0.0380882
R51750 ASIG5V.n667 ASIG5V.n605 0.0380882
R51751 ASIG5V.n677 ASIG5V.n605 0.0380882
R51752 ASIG5V.n678 ASIG5V.n677 0.0380882
R51753 ASIG5V.n679 ASIG5V.n678 0.0380882
R51754 ASIG5V.n679 ASIG5V.n603 0.0380882
R51755 ASIG5V.n689 ASIG5V.n603 0.0380882
R51756 ASIG5V.n690 ASIG5V.n689 0.0380882
R51757 ASIG5V.n691 ASIG5V.n690 0.0380882
R51758 ASIG5V.n691 ASIG5V.n601 0.0380882
R51759 ASIG5V.n701 ASIG5V.n601 0.0380882
R51760 ASIG5V.n702 ASIG5V.n701 0.0380882
R51761 ASIG5V.n703 ASIG5V.n702 0.0380882
R51762 ASIG5V.n703 ASIG5V.n599 0.0380882
R51763 ASIG5V.n713 ASIG5V.n599 0.0380882
R51764 ASIG5V.n714 ASIG5V.n713 0.0380882
R51765 ASIG5V.n715 ASIG5V.n714 0.0380882
R51766 ASIG5V.n715 ASIG5V.n597 0.0380882
R51767 ASIG5V.n725 ASIG5V.n597 0.0380882
R51768 ASIG5V.n726 ASIG5V.n725 0.0380882
R51769 ASIG5V.n727 ASIG5V.n726 0.0380882
R51770 ASIG5V.n727 ASIG5V.n595 0.0380882
R51771 ASIG5V.n737 ASIG5V.n595 0.0380882
R51772 ASIG5V.n738 ASIG5V.n737 0.0380882
R51773 ASIG5V.n739 ASIG5V.n738 0.0380882
R51774 ASIG5V.n739 ASIG5V.n593 0.0380882
R51775 ASIG5V.n749 ASIG5V.n593 0.0380882
R51776 ASIG5V.n750 ASIG5V.n749 0.0380882
R51777 ASIG5V.n751 ASIG5V.n750 0.0380882
R51778 ASIG5V.n751 ASIG5V.n591 0.0380882
R51779 ASIG5V.n761 ASIG5V.n591 0.0380882
R51780 ASIG5V.n762 ASIG5V.n761 0.0380882
R51781 ASIG5V.n763 ASIG5V.n762 0.0380882
R51782 ASIG5V.n763 ASIG5V.n589 0.0380882
R51783 ASIG5V.n773 ASIG5V.n589 0.0380882
R51784 ASIG5V.n774 ASIG5V.n773 0.0380882
R51785 ASIG5V.n775 ASIG5V.n774 0.0380882
R51786 ASIG5V.n775 ASIG5V.n587 0.0380882
R51787 ASIG5V.n785 ASIG5V.n587 0.0380882
R51788 ASIG5V.n786 ASIG5V.n785 0.0380882
R51789 ASIG5V.n787 ASIG5V.n786 0.0380882
R51790 ASIG5V.n787 ASIG5V.n585 0.0380882
R51791 ASIG5V.n797 ASIG5V.n585 0.0380882
R51792 ASIG5V.n798 ASIG5V.n797 0.0380882
R51793 ASIG5V.n799 ASIG5V.n798 0.0380882
R51794 ASIG5V.n799 ASIG5V.n583 0.0380882
R51795 ASIG5V.n809 ASIG5V.n583 0.0380882
R51796 ASIG5V.n810 ASIG5V.n809 0.0380882
R51797 ASIG5V.n811 ASIG5V.n810 0.0380882
R51798 ASIG5V.n811 ASIG5V.n581 0.0380882
R51799 ASIG5V.n821 ASIG5V.n581 0.0380882
R51800 ASIG5V.n822 ASIG5V.n821 0.0380882
R51801 ASIG5V.n823 ASIG5V.n822 0.0380882
R51802 ASIG5V.n823 ASIG5V.n579 0.0380882
R51803 ASIG5V.n833 ASIG5V.n579 0.0380882
R51804 ASIG5V.n834 ASIG5V.n833 0.0380882
R51805 ASIG5V.n835 ASIG5V.n834 0.0380882
R51806 ASIG5V.n835 ASIG5V.n577 0.0380882
R51807 ASIG5V.n845 ASIG5V.n577 0.0380882
R51808 ASIG5V.n846 ASIG5V.n845 0.0380882
R51809 ASIG5V.n847 ASIG5V.n846 0.0380882
R51810 ASIG5V.n847 ASIG5V.n575 0.0380882
R51811 ASIG5V.n857 ASIG5V.n575 0.0380882
R51812 ASIG5V.n858 ASIG5V.n857 0.0380882
R51813 ASIG5V.n12296 ASIG5V.n858 0.0380882
R51814 ASIG5V.n12296 ASIG5V.n12295 0.0380882
R51815 ASIG5V.n617 ASIG5V.n614 0.0380882
R51816 ASIG5V.n620 ASIG5V.n617 0.0380882
R51817 ASIG5V.n624 ASIG5V.n620 0.0380882
R51818 ASIG5V.n628 ASIG5V.n624 0.0380882
R51819 ASIG5V.n628 ASIG5V.n612 0.0380882
R51820 ASIG5V.n632 ASIG5V.n612 0.0380882
R51821 ASIG5V.n636 ASIG5V.n632 0.0380882
R51822 ASIG5V.n640 ASIG5V.n636 0.0380882
R51823 ASIG5V.n640 ASIG5V.n610 0.0380882
R51824 ASIG5V.n644 ASIG5V.n610 0.0380882
R51825 ASIG5V.n648 ASIG5V.n644 0.0380882
R51826 ASIG5V.n652 ASIG5V.n648 0.0380882
R51827 ASIG5V.n652 ASIG5V.n608 0.0380882
R51828 ASIG5V.n656 ASIG5V.n608 0.0380882
R51829 ASIG5V.n660 ASIG5V.n656 0.0380882
R51830 ASIG5V.n664 ASIG5V.n660 0.0380882
R51831 ASIG5V.n664 ASIG5V.n606 0.0380882
R51832 ASIG5V.n668 ASIG5V.n606 0.0380882
R51833 ASIG5V.n672 ASIG5V.n668 0.0380882
R51834 ASIG5V.n676 ASIG5V.n672 0.0380882
R51835 ASIG5V.n676 ASIG5V.n604 0.0380882
R51836 ASIG5V.n680 ASIG5V.n604 0.0380882
R51837 ASIG5V.n684 ASIG5V.n680 0.0380882
R51838 ASIG5V.n688 ASIG5V.n684 0.0380882
R51839 ASIG5V.n688 ASIG5V.n602 0.0380882
R51840 ASIG5V.n692 ASIG5V.n602 0.0380882
R51841 ASIG5V.n696 ASIG5V.n692 0.0380882
R51842 ASIG5V.n700 ASIG5V.n696 0.0380882
R51843 ASIG5V.n700 ASIG5V.n600 0.0380882
R51844 ASIG5V.n704 ASIG5V.n600 0.0380882
R51845 ASIG5V.n708 ASIG5V.n704 0.0380882
R51846 ASIG5V.n712 ASIG5V.n708 0.0380882
R51847 ASIG5V.n712 ASIG5V.n598 0.0380882
R51848 ASIG5V.n716 ASIG5V.n598 0.0380882
R51849 ASIG5V.n720 ASIG5V.n716 0.0380882
R51850 ASIG5V.n724 ASIG5V.n720 0.0380882
R51851 ASIG5V.n724 ASIG5V.n596 0.0380882
R51852 ASIG5V.n728 ASIG5V.n596 0.0380882
R51853 ASIG5V.n732 ASIG5V.n728 0.0380882
R51854 ASIG5V.n736 ASIG5V.n732 0.0380882
R51855 ASIG5V.n736 ASIG5V.n594 0.0380882
R51856 ASIG5V.n740 ASIG5V.n594 0.0380882
R51857 ASIG5V.n744 ASIG5V.n740 0.0380882
R51858 ASIG5V.n748 ASIG5V.n744 0.0380882
R51859 ASIG5V.n748 ASIG5V.n592 0.0380882
R51860 ASIG5V.n752 ASIG5V.n592 0.0380882
R51861 ASIG5V.n756 ASIG5V.n752 0.0380882
R51862 ASIG5V.n760 ASIG5V.n756 0.0380882
R51863 ASIG5V.n760 ASIG5V.n590 0.0380882
R51864 ASIG5V.n764 ASIG5V.n590 0.0380882
R51865 ASIG5V.n768 ASIG5V.n764 0.0380882
R51866 ASIG5V.n772 ASIG5V.n768 0.0380882
R51867 ASIG5V.n772 ASIG5V.n588 0.0380882
R51868 ASIG5V.n776 ASIG5V.n588 0.0380882
R51869 ASIG5V.n780 ASIG5V.n776 0.0380882
R51870 ASIG5V.n784 ASIG5V.n780 0.0380882
R51871 ASIG5V.n784 ASIG5V.n586 0.0380882
R51872 ASIG5V.n788 ASIG5V.n586 0.0380882
R51873 ASIG5V.n792 ASIG5V.n788 0.0380882
R51874 ASIG5V.n796 ASIG5V.n792 0.0380882
R51875 ASIG5V.n796 ASIG5V.n584 0.0380882
R51876 ASIG5V.n800 ASIG5V.n584 0.0380882
R51877 ASIG5V.n804 ASIG5V.n800 0.0380882
R51878 ASIG5V.n808 ASIG5V.n804 0.0380882
R51879 ASIG5V.n808 ASIG5V.n582 0.0380882
R51880 ASIG5V.n812 ASIG5V.n582 0.0380882
R51881 ASIG5V.n816 ASIG5V.n812 0.0380882
R51882 ASIG5V.n820 ASIG5V.n816 0.0380882
R51883 ASIG5V.n820 ASIG5V.n580 0.0380882
R51884 ASIG5V.n824 ASIG5V.n580 0.0380882
R51885 ASIG5V.n828 ASIG5V.n824 0.0380882
R51886 ASIG5V.n832 ASIG5V.n828 0.0380882
R51887 ASIG5V.n832 ASIG5V.n578 0.0380882
R51888 ASIG5V.n836 ASIG5V.n578 0.0380882
R51889 ASIG5V.n840 ASIG5V.n836 0.0380882
R51890 ASIG5V.n844 ASIG5V.n840 0.0380882
R51891 ASIG5V.n844 ASIG5V.n576 0.0380882
R51892 ASIG5V.n848 ASIG5V.n576 0.0380882
R51893 ASIG5V.n852 ASIG5V.n848 0.0380882
R51894 ASIG5V.n856 ASIG5V.n852 0.0380882
R51895 ASIG5V.n856 ASIG5V.n574 0.0380882
R51896 ASIG5V.n12297 ASIG5V.n574 0.0380882
R51897 ASIG5V.n12297 ASIG5V.n573 0.0380882
R51898 ASIG5V.n964 ASIG5V.n869 0.0380882
R51899 ASIG5V.n975 ASIG5V.n964 0.0380882
R51900 ASIG5V.n976 ASIG5V.n975 0.0380882
R51901 ASIG5V.n977 ASIG5V.n976 0.0380882
R51902 ASIG5V.n977 ASIG5V.n960 0.0380882
R51903 ASIG5V.n987 ASIG5V.n960 0.0380882
R51904 ASIG5V.n988 ASIG5V.n987 0.0380882
R51905 ASIG5V.n989 ASIG5V.n988 0.0380882
R51906 ASIG5V.n989 ASIG5V.n956 0.0380882
R51907 ASIG5V.n999 ASIG5V.n956 0.0380882
R51908 ASIG5V.n1000 ASIG5V.n999 0.0380882
R51909 ASIG5V.n1001 ASIG5V.n1000 0.0380882
R51910 ASIG5V.n1001 ASIG5V.n952 0.0380882
R51911 ASIG5V.n1011 ASIG5V.n952 0.0380882
R51912 ASIG5V.n1012 ASIG5V.n1011 0.0380882
R51913 ASIG5V.n1013 ASIG5V.n1012 0.0380882
R51914 ASIG5V.n1013 ASIG5V.n948 0.0380882
R51915 ASIG5V.n1023 ASIG5V.n948 0.0380882
R51916 ASIG5V.n1024 ASIG5V.n1023 0.0380882
R51917 ASIG5V.n1025 ASIG5V.n1024 0.0380882
R51918 ASIG5V.n1025 ASIG5V.n944 0.0380882
R51919 ASIG5V.n1035 ASIG5V.n944 0.0380882
R51920 ASIG5V.n1036 ASIG5V.n1035 0.0380882
R51921 ASIG5V.n1037 ASIG5V.n1036 0.0380882
R51922 ASIG5V.n1037 ASIG5V.n940 0.0380882
R51923 ASIG5V.n1047 ASIG5V.n940 0.0380882
R51924 ASIG5V.n1048 ASIG5V.n1047 0.0380882
R51925 ASIG5V.n1049 ASIG5V.n1048 0.0380882
R51926 ASIG5V.n1049 ASIG5V.n936 0.0380882
R51927 ASIG5V.n1059 ASIG5V.n936 0.0380882
R51928 ASIG5V.n1060 ASIG5V.n1059 0.0380882
R51929 ASIG5V.n1061 ASIG5V.n1060 0.0380882
R51930 ASIG5V.n1061 ASIG5V.n932 0.0380882
R51931 ASIG5V.n1071 ASIG5V.n932 0.0380882
R51932 ASIG5V.n1072 ASIG5V.n1071 0.0380882
R51933 ASIG5V.n1073 ASIG5V.n1072 0.0380882
R51934 ASIG5V.n1073 ASIG5V.n928 0.0380882
R51935 ASIG5V.n1083 ASIG5V.n928 0.0380882
R51936 ASIG5V.n1084 ASIG5V.n1083 0.0380882
R51937 ASIG5V.n1085 ASIG5V.n1084 0.0380882
R51938 ASIG5V.n1085 ASIG5V.n924 0.0380882
R51939 ASIG5V.n1095 ASIG5V.n924 0.0380882
R51940 ASIG5V.n1096 ASIG5V.n1095 0.0380882
R51941 ASIG5V.n1097 ASIG5V.n1096 0.0380882
R51942 ASIG5V.n1097 ASIG5V.n920 0.0380882
R51943 ASIG5V.n1107 ASIG5V.n920 0.0380882
R51944 ASIG5V.n1108 ASIG5V.n1107 0.0380882
R51945 ASIG5V.n1109 ASIG5V.n1108 0.0380882
R51946 ASIG5V.n1109 ASIG5V.n916 0.0380882
R51947 ASIG5V.n1119 ASIG5V.n916 0.0380882
R51948 ASIG5V.n1120 ASIG5V.n1119 0.0380882
R51949 ASIG5V.n1121 ASIG5V.n1120 0.0380882
R51950 ASIG5V.n1121 ASIG5V.n912 0.0380882
R51951 ASIG5V.n1131 ASIG5V.n912 0.0380882
R51952 ASIG5V.n1132 ASIG5V.n1131 0.0380882
R51953 ASIG5V.n1133 ASIG5V.n1132 0.0380882
R51954 ASIG5V.n1133 ASIG5V.n908 0.0380882
R51955 ASIG5V.n1143 ASIG5V.n908 0.0380882
R51956 ASIG5V.n1144 ASIG5V.n1143 0.0380882
R51957 ASIG5V.n1145 ASIG5V.n1144 0.0380882
R51958 ASIG5V.n1145 ASIG5V.n904 0.0380882
R51959 ASIG5V.n1155 ASIG5V.n904 0.0380882
R51960 ASIG5V.n1156 ASIG5V.n1155 0.0380882
R51961 ASIG5V.n1157 ASIG5V.n1156 0.0380882
R51962 ASIG5V.n1157 ASIG5V.n900 0.0380882
R51963 ASIG5V.n1167 ASIG5V.n900 0.0380882
R51964 ASIG5V.n1168 ASIG5V.n1167 0.0380882
R51965 ASIG5V.n1169 ASIG5V.n1168 0.0380882
R51966 ASIG5V.n1169 ASIG5V.n896 0.0380882
R51967 ASIG5V.n1179 ASIG5V.n896 0.0380882
R51968 ASIG5V.n1180 ASIG5V.n1179 0.0380882
R51969 ASIG5V.n1181 ASIG5V.n1180 0.0380882
R51970 ASIG5V.n1181 ASIG5V.n892 0.0380882
R51971 ASIG5V.n1191 ASIG5V.n892 0.0380882
R51972 ASIG5V.n1192 ASIG5V.n1191 0.0380882
R51973 ASIG5V.n1193 ASIG5V.n1192 0.0380882
R51974 ASIG5V.n1193 ASIG5V.n888 0.0380882
R51975 ASIG5V.n1203 ASIG5V.n888 0.0380882
R51976 ASIG5V.n1204 ASIG5V.n1203 0.0380882
R51977 ASIG5V.n1206 ASIG5V.n1204 0.0380882
R51978 ASIG5V.n1206 ASIG5V.n1205 0.0380882
R51979 ASIG5V.n1205 ASIG5V.n883 0.0380882
R51980 ASIG5V.n1216 ASIG5V.n883 0.0380882
R51981 ASIG5V.n966 ASIG5V.n965 0.0380882
R51982 ASIG5V.n974 ASIG5V.n965 0.0380882
R51983 ASIG5V.n974 ASIG5V.n963 0.0380882
R51984 ASIG5V.n978 ASIG5V.n963 0.0380882
R51985 ASIG5V.n978 ASIG5V.n961 0.0380882
R51986 ASIG5V.n986 ASIG5V.n961 0.0380882
R51987 ASIG5V.n986 ASIG5V.n959 0.0380882
R51988 ASIG5V.n990 ASIG5V.n959 0.0380882
R51989 ASIG5V.n990 ASIG5V.n957 0.0380882
R51990 ASIG5V.n998 ASIG5V.n957 0.0380882
R51991 ASIG5V.n998 ASIG5V.n955 0.0380882
R51992 ASIG5V.n1002 ASIG5V.n955 0.0380882
R51993 ASIG5V.n1002 ASIG5V.n953 0.0380882
R51994 ASIG5V.n1010 ASIG5V.n953 0.0380882
R51995 ASIG5V.n1010 ASIG5V.n951 0.0380882
R51996 ASIG5V.n1014 ASIG5V.n951 0.0380882
R51997 ASIG5V.n1014 ASIG5V.n949 0.0380882
R51998 ASIG5V.n1022 ASIG5V.n949 0.0380882
R51999 ASIG5V.n1022 ASIG5V.n947 0.0380882
R52000 ASIG5V.n1026 ASIG5V.n947 0.0380882
R52001 ASIG5V.n1026 ASIG5V.n945 0.0380882
R52002 ASIG5V.n1034 ASIG5V.n945 0.0380882
R52003 ASIG5V.n1034 ASIG5V.n943 0.0380882
R52004 ASIG5V.n1038 ASIG5V.n943 0.0380882
R52005 ASIG5V.n1038 ASIG5V.n941 0.0380882
R52006 ASIG5V.n1046 ASIG5V.n941 0.0380882
R52007 ASIG5V.n1046 ASIG5V.n939 0.0380882
R52008 ASIG5V.n1050 ASIG5V.n939 0.0380882
R52009 ASIG5V.n1050 ASIG5V.n937 0.0380882
R52010 ASIG5V.n1058 ASIG5V.n937 0.0380882
R52011 ASIG5V.n1058 ASIG5V.n935 0.0380882
R52012 ASIG5V.n1062 ASIG5V.n935 0.0380882
R52013 ASIG5V.n1062 ASIG5V.n933 0.0380882
R52014 ASIG5V.n1070 ASIG5V.n933 0.0380882
R52015 ASIG5V.n1070 ASIG5V.n931 0.0380882
R52016 ASIG5V.n1074 ASIG5V.n931 0.0380882
R52017 ASIG5V.n1074 ASIG5V.n929 0.0380882
R52018 ASIG5V.n1082 ASIG5V.n929 0.0380882
R52019 ASIG5V.n1082 ASIG5V.n927 0.0380882
R52020 ASIG5V.n1086 ASIG5V.n927 0.0380882
R52021 ASIG5V.n1086 ASIG5V.n925 0.0380882
R52022 ASIG5V.n1094 ASIG5V.n925 0.0380882
R52023 ASIG5V.n1094 ASIG5V.n923 0.0380882
R52024 ASIG5V.n1098 ASIG5V.n923 0.0380882
R52025 ASIG5V.n1098 ASIG5V.n921 0.0380882
R52026 ASIG5V.n1106 ASIG5V.n921 0.0380882
R52027 ASIG5V.n1106 ASIG5V.n919 0.0380882
R52028 ASIG5V.n1110 ASIG5V.n919 0.0380882
R52029 ASIG5V.n1110 ASIG5V.n917 0.0380882
R52030 ASIG5V.n1118 ASIG5V.n917 0.0380882
R52031 ASIG5V.n1118 ASIG5V.n915 0.0380882
R52032 ASIG5V.n1122 ASIG5V.n915 0.0380882
R52033 ASIG5V.n1122 ASIG5V.n913 0.0380882
R52034 ASIG5V.n1130 ASIG5V.n913 0.0380882
R52035 ASIG5V.n1130 ASIG5V.n911 0.0380882
R52036 ASIG5V.n1134 ASIG5V.n911 0.0380882
R52037 ASIG5V.n1134 ASIG5V.n909 0.0380882
R52038 ASIG5V.n1142 ASIG5V.n909 0.0380882
R52039 ASIG5V.n1142 ASIG5V.n907 0.0380882
R52040 ASIG5V.n1146 ASIG5V.n907 0.0380882
R52041 ASIG5V.n1146 ASIG5V.n905 0.0380882
R52042 ASIG5V.n1154 ASIG5V.n905 0.0380882
R52043 ASIG5V.n1154 ASIG5V.n903 0.0380882
R52044 ASIG5V.n1158 ASIG5V.n903 0.0380882
R52045 ASIG5V.n1158 ASIG5V.n901 0.0380882
R52046 ASIG5V.n1166 ASIG5V.n901 0.0380882
R52047 ASIG5V.n1166 ASIG5V.n899 0.0380882
R52048 ASIG5V.n1170 ASIG5V.n899 0.0380882
R52049 ASIG5V.n1170 ASIG5V.n897 0.0380882
R52050 ASIG5V.n1178 ASIG5V.n897 0.0380882
R52051 ASIG5V.n1178 ASIG5V.n895 0.0380882
R52052 ASIG5V.n1182 ASIG5V.n895 0.0380882
R52053 ASIG5V.n1182 ASIG5V.n893 0.0380882
R52054 ASIG5V.n1190 ASIG5V.n893 0.0380882
R52055 ASIG5V.n1190 ASIG5V.n891 0.0380882
R52056 ASIG5V.n1194 ASIG5V.n891 0.0380882
R52057 ASIG5V.n1194 ASIG5V.n889 0.0380882
R52058 ASIG5V.n1202 ASIG5V.n889 0.0380882
R52059 ASIG5V.n1202 ASIG5V.n887 0.0380882
R52060 ASIG5V.n1207 ASIG5V.n887 0.0380882
R52061 ASIG5V.n1207 ASIG5V.n885 0.0380882
R52062 ASIG5V.n885 ASIG5V.n884 0.0380882
R52063 ASIG5V.n1215 ASIG5V.n884 0.0380882
R52064 ASIG5V.n12022 ASIG5V.n12021 0.0380882
R52065 ASIG5V.n12023 ASIG5V.n12022 0.0380882
R52066 ASIG5V.n12023 ASIG5V.n1312 0.0380882
R52067 ASIG5V.n12033 ASIG5V.n1312 0.0380882
R52068 ASIG5V.n12034 ASIG5V.n12033 0.0380882
R52069 ASIG5V.n12035 ASIG5V.n12034 0.0380882
R52070 ASIG5V.n12035 ASIG5V.n1310 0.0380882
R52071 ASIG5V.n12045 ASIG5V.n1310 0.0380882
R52072 ASIG5V.n12046 ASIG5V.n12045 0.0380882
R52073 ASIG5V.n12047 ASIG5V.n12046 0.0380882
R52074 ASIG5V.n12047 ASIG5V.n1308 0.0380882
R52075 ASIG5V.n12057 ASIG5V.n1308 0.0380882
R52076 ASIG5V.n12058 ASIG5V.n12057 0.0380882
R52077 ASIG5V.n12059 ASIG5V.n12058 0.0380882
R52078 ASIG5V.n12059 ASIG5V.n1306 0.0380882
R52079 ASIG5V.n12069 ASIG5V.n1306 0.0380882
R52080 ASIG5V.n12070 ASIG5V.n12069 0.0380882
R52081 ASIG5V.n12071 ASIG5V.n12070 0.0380882
R52082 ASIG5V.n12071 ASIG5V.n1304 0.0380882
R52083 ASIG5V.n12081 ASIG5V.n1304 0.0380882
R52084 ASIG5V.n12082 ASIG5V.n12081 0.0380882
R52085 ASIG5V.n12083 ASIG5V.n12082 0.0380882
R52086 ASIG5V.n12083 ASIG5V.n1302 0.0380882
R52087 ASIG5V.n12093 ASIG5V.n1302 0.0380882
R52088 ASIG5V.n12094 ASIG5V.n12093 0.0380882
R52089 ASIG5V.n12095 ASIG5V.n12094 0.0380882
R52090 ASIG5V.n12095 ASIG5V.n1300 0.0380882
R52091 ASIG5V.n12105 ASIG5V.n1300 0.0380882
R52092 ASIG5V.n12106 ASIG5V.n12105 0.0380882
R52093 ASIG5V.n12107 ASIG5V.n12106 0.0380882
R52094 ASIG5V.n12107 ASIG5V.n1298 0.0380882
R52095 ASIG5V.n12117 ASIG5V.n1298 0.0380882
R52096 ASIG5V.n12118 ASIG5V.n12117 0.0380882
R52097 ASIG5V.n12119 ASIG5V.n12118 0.0380882
R52098 ASIG5V.n12119 ASIG5V.n1296 0.0380882
R52099 ASIG5V.n12129 ASIG5V.n1296 0.0380882
R52100 ASIG5V.n12130 ASIG5V.n12129 0.0380882
R52101 ASIG5V.n12131 ASIG5V.n12130 0.0380882
R52102 ASIG5V.n12131 ASIG5V.n1294 0.0380882
R52103 ASIG5V.n12141 ASIG5V.n1294 0.0380882
R52104 ASIG5V.n12142 ASIG5V.n12141 0.0380882
R52105 ASIG5V.n12143 ASIG5V.n12142 0.0380882
R52106 ASIG5V.n12143 ASIG5V.n1292 0.0380882
R52107 ASIG5V.n12153 ASIG5V.n1292 0.0380882
R52108 ASIG5V.n12154 ASIG5V.n12153 0.0380882
R52109 ASIG5V.n12155 ASIG5V.n12154 0.0380882
R52110 ASIG5V.n12155 ASIG5V.n1290 0.0380882
R52111 ASIG5V.n12165 ASIG5V.n1290 0.0380882
R52112 ASIG5V.n12166 ASIG5V.n12165 0.0380882
R52113 ASIG5V.n12167 ASIG5V.n12166 0.0380882
R52114 ASIG5V.n12167 ASIG5V.n1288 0.0380882
R52115 ASIG5V.n12177 ASIG5V.n1288 0.0380882
R52116 ASIG5V.n12178 ASIG5V.n12177 0.0380882
R52117 ASIG5V.n12179 ASIG5V.n12178 0.0380882
R52118 ASIG5V.n12179 ASIG5V.n1286 0.0380882
R52119 ASIG5V.n12189 ASIG5V.n1286 0.0380882
R52120 ASIG5V.n12190 ASIG5V.n12189 0.0380882
R52121 ASIG5V.n12191 ASIG5V.n12190 0.0380882
R52122 ASIG5V.n12191 ASIG5V.n1284 0.0380882
R52123 ASIG5V.n12201 ASIG5V.n1284 0.0380882
R52124 ASIG5V.n12202 ASIG5V.n12201 0.0380882
R52125 ASIG5V.n12203 ASIG5V.n12202 0.0380882
R52126 ASIG5V.n12203 ASIG5V.n1282 0.0380882
R52127 ASIG5V.n12213 ASIG5V.n1282 0.0380882
R52128 ASIG5V.n12214 ASIG5V.n12213 0.0380882
R52129 ASIG5V.n12215 ASIG5V.n12214 0.0380882
R52130 ASIG5V.n12215 ASIG5V.n1280 0.0380882
R52131 ASIG5V.n12225 ASIG5V.n1280 0.0380882
R52132 ASIG5V.n12226 ASIG5V.n12225 0.0380882
R52133 ASIG5V.n12227 ASIG5V.n12226 0.0380882
R52134 ASIG5V.n12227 ASIG5V.n1278 0.0380882
R52135 ASIG5V.n12237 ASIG5V.n1278 0.0380882
R52136 ASIG5V.n12238 ASIG5V.n12237 0.0380882
R52137 ASIG5V.n12239 ASIG5V.n12238 0.0380882
R52138 ASIG5V.n12239 ASIG5V.n1276 0.0380882
R52139 ASIG5V.n12249 ASIG5V.n1276 0.0380882
R52140 ASIG5V.n12250 ASIG5V.n12249 0.0380882
R52141 ASIG5V.n12251 ASIG5V.n12250 0.0380882
R52142 ASIG5V.n12251 ASIG5V.n1274 0.0380882
R52143 ASIG5V.n12261 ASIG5V.n1274 0.0380882
R52144 ASIG5V.n12262 ASIG5V.n12261 0.0380882
R52145 ASIG5V.n12263 ASIG5V.n12262 0.0380882
R52146 ASIG5V.n12263 ASIG5V.n1220 0.0380882
R52147 ASIG5V.n12020 ASIG5V.n1315 0.0380882
R52148 ASIG5V.n12024 ASIG5V.n1315 0.0380882
R52149 ASIG5V.n12028 ASIG5V.n12024 0.0380882
R52150 ASIG5V.n12032 ASIG5V.n12028 0.0380882
R52151 ASIG5V.n12032 ASIG5V.n1311 0.0380882
R52152 ASIG5V.n12036 ASIG5V.n1311 0.0380882
R52153 ASIG5V.n12040 ASIG5V.n12036 0.0380882
R52154 ASIG5V.n12044 ASIG5V.n12040 0.0380882
R52155 ASIG5V.n12044 ASIG5V.n1309 0.0380882
R52156 ASIG5V.n12048 ASIG5V.n1309 0.0380882
R52157 ASIG5V.n12052 ASIG5V.n12048 0.0380882
R52158 ASIG5V.n12056 ASIG5V.n12052 0.0380882
R52159 ASIG5V.n12056 ASIG5V.n1307 0.0380882
R52160 ASIG5V.n12060 ASIG5V.n1307 0.0380882
R52161 ASIG5V.n12064 ASIG5V.n12060 0.0380882
R52162 ASIG5V.n12068 ASIG5V.n12064 0.0380882
R52163 ASIG5V.n12068 ASIG5V.n1305 0.0380882
R52164 ASIG5V.n12072 ASIG5V.n1305 0.0380882
R52165 ASIG5V.n12076 ASIG5V.n12072 0.0380882
R52166 ASIG5V.n12080 ASIG5V.n12076 0.0380882
R52167 ASIG5V.n12080 ASIG5V.n1303 0.0380882
R52168 ASIG5V.n12084 ASIG5V.n1303 0.0380882
R52169 ASIG5V.n12088 ASIG5V.n12084 0.0380882
R52170 ASIG5V.n12092 ASIG5V.n12088 0.0380882
R52171 ASIG5V.n12092 ASIG5V.n1301 0.0380882
R52172 ASIG5V.n12096 ASIG5V.n1301 0.0380882
R52173 ASIG5V.n12100 ASIG5V.n12096 0.0380882
R52174 ASIG5V.n12104 ASIG5V.n12100 0.0380882
R52175 ASIG5V.n12104 ASIG5V.n1299 0.0380882
R52176 ASIG5V.n12108 ASIG5V.n1299 0.0380882
R52177 ASIG5V.n12112 ASIG5V.n12108 0.0380882
R52178 ASIG5V.n12116 ASIG5V.n12112 0.0380882
R52179 ASIG5V.n12116 ASIG5V.n1297 0.0380882
R52180 ASIG5V.n12120 ASIG5V.n1297 0.0380882
R52181 ASIG5V.n12124 ASIG5V.n12120 0.0380882
R52182 ASIG5V.n12128 ASIG5V.n12124 0.0380882
R52183 ASIG5V.n12128 ASIG5V.n1295 0.0380882
R52184 ASIG5V.n12132 ASIG5V.n1295 0.0380882
R52185 ASIG5V.n12136 ASIG5V.n12132 0.0380882
R52186 ASIG5V.n12140 ASIG5V.n12136 0.0380882
R52187 ASIG5V.n12140 ASIG5V.n1293 0.0380882
R52188 ASIG5V.n12144 ASIG5V.n1293 0.0380882
R52189 ASIG5V.n12148 ASIG5V.n12144 0.0380882
R52190 ASIG5V.n12152 ASIG5V.n12148 0.0380882
R52191 ASIG5V.n12152 ASIG5V.n1291 0.0380882
R52192 ASIG5V.n12156 ASIG5V.n1291 0.0380882
R52193 ASIG5V.n12160 ASIG5V.n12156 0.0380882
R52194 ASIG5V.n12164 ASIG5V.n12160 0.0380882
R52195 ASIG5V.n12164 ASIG5V.n1289 0.0380882
R52196 ASIG5V.n12168 ASIG5V.n1289 0.0380882
R52197 ASIG5V.n12172 ASIG5V.n12168 0.0380882
R52198 ASIG5V.n12176 ASIG5V.n12172 0.0380882
R52199 ASIG5V.n12176 ASIG5V.n1287 0.0380882
R52200 ASIG5V.n12180 ASIG5V.n1287 0.0380882
R52201 ASIG5V.n12184 ASIG5V.n12180 0.0380882
R52202 ASIG5V.n12188 ASIG5V.n12184 0.0380882
R52203 ASIG5V.n12188 ASIG5V.n1285 0.0380882
R52204 ASIG5V.n12192 ASIG5V.n1285 0.0380882
R52205 ASIG5V.n12196 ASIG5V.n12192 0.0380882
R52206 ASIG5V.n12200 ASIG5V.n12196 0.0380882
R52207 ASIG5V.n12200 ASIG5V.n1283 0.0380882
R52208 ASIG5V.n12204 ASIG5V.n1283 0.0380882
R52209 ASIG5V.n12208 ASIG5V.n12204 0.0380882
R52210 ASIG5V.n12212 ASIG5V.n12208 0.0380882
R52211 ASIG5V.n12212 ASIG5V.n1281 0.0380882
R52212 ASIG5V.n12216 ASIG5V.n1281 0.0380882
R52213 ASIG5V.n12220 ASIG5V.n12216 0.0380882
R52214 ASIG5V.n12224 ASIG5V.n12220 0.0380882
R52215 ASIG5V.n12224 ASIG5V.n1279 0.0380882
R52216 ASIG5V.n12228 ASIG5V.n1279 0.0380882
R52217 ASIG5V.n12232 ASIG5V.n12228 0.0380882
R52218 ASIG5V.n12236 ASIG5V.n12232 0.0380882
R52219 ASIG5V.n12236 ASIG5V.n1277 0.0380882
R52220 ASIG5V.n12240 ASIG5V.n1277 0.0380882
R52221 ASIG5V.n12244 ASIG5V.n12240 0.0380882
R52222 ASIG5V.n12248 ASIG5V.n12244 0.0380882
R52223 ASIG5V.n12248 ASIG5V.n1275 0.0380882
R52224 ASIG5V.n12252 ASIG5V.n1275 0.0380882
R52225 ASIG5V.n12256 ASIG5V.n12252 0.0380882
R52226 ASIG5V.n12260 ASIG5V.n12256 0.0380882
R52227 ASIG5V.n12260 ASIG5V.n1273 0.0380882
R52228 ASIG5V.n12264 ASIG5V.n1273 0.0380882
R52229 ASIG5V.n12264 ASIG5V.n1270 0.0380882
R52230 ASIG5V.n1481 ASIG5V.n1479 0.0380882
R52231 ASIG5V.n1482 ASIG5V.n1481 0.0380882
R52232 ASIG5V.n1483 ASIG5V.n1482 0.0380882
R52233 ASIG5V.n1483 ASIG5V.n1476 0.0380882
R52234 ASIG5V.n1490 ASIG5V.n1476 0.0380882
R52235 ASIG5V.n1491 ASIG5V.n1490 0.0380882
R52236 ASIG5V.n1492 ASIG5V.n1491 0.0380882
R52237 ASIG5V.n1492 ASIG5V.n1473 0.0380882
R52238 ASIG5V.n1499 ASIG5V.n1473 0.0380882
R52239 ASIG5V.n1500 ASIG5V.n1499 0.0380882
R52240 ASIG5V.n1501 ASIG5V.n1500 0.0380882
R52241 ASIG5V.n1501 ASIG5V.n1470 0.0380882
R52242 ASIG5V.n1508 ASIG5V.n1470 0.0380882
R52243 ASIG5V.n1509 ASIG5V.n1508 0.0380882
R52244 ASIG5V.n1510 ASIG5V.n1509 0.0380882
R52245 ASIG5V.n1510 ASIG5V.n1467 0.0380882
R52246 ASIG5V.n1517 ASIG5V.n1467 0.0380882
R52247 ASIG5V.n1518 ASIG5V.n1517 0.0380882
R52248 ASIG5V.n1519 ASIG5V.n1518 0.0380882
R52249 ASIG5V.n1519 ASIG5V.n1464 0.0380882
R52250 ASIG5V.n1526 ASIG5V.n1464 0.0380882
R52251 ASIG5V.n1527 ASIG5V.n1526 0.0380882
R52252 ASIG5V.n1528 ASIG5V.n1527 0.0380882
R52253 ASIG5V.n1528 ASIG5V.n1461 0.0380882
R52254 ASIG5V.n1535 ASIG5V.n1461 0.0380882
R52255 ASIG5V.n1536 ASIG5V.n1535 0.0380882
R52256 ASIG5V.n1537 ASIG5V.n1536 0.0380882
R52257 ASIG5V.n1537 ASIG5V.n1458 0.0380882
R52258 ASIG5V.n1544 ASIG5V.n1458 0.0380882
R52259 ASIG5V.n1545 ASIG5V.n1544 0.0380882
R52260 ASIG5V.n1546 ASIG5V.n1545 0.0380882
R52261 ASIG5V.n1546 ASIG5V.n1455 0.0380882
R52262 ASIG5V.n1553 ASIG5V.n1455 0.0380882
R52263 ASIG5V.n1554 ASIG5V.n1553 0.0380882
R52264 ASIG5V.n1555 ASIG5V.n1554 0.0380882
R52265 ASIG5V.n1555 ASIG5V.n1452 0.0380882
R52266 ASIG5V.n1562 ASIG5V.n1452 0.0380882
R52267 ASIG5V.n1563 ASIG5V.n1562 0.0380882
R52268 ASIG5V.n1564 ASIG5V.n1563 0.0380882
R52269 ASIG5V.n1564 ASIG5V.n1449 0.0380882
R52270 ASIG5V.n1571 ASIG5V.n1449 0.0380882
R52271 ASIG5V.n1572 ASIG5V.n1571 0.0380882
R52272 ASIG5V.n1573 ASIG5V.n1572 0.0380882
R52273 ASIG5V.n1573 ASIG5V.n1446 0.0380882
R52274 ASIG5V.n1580 ASIG5V.n1446 0.0380882
R52275 ASIG5V.n1581 ASIG5V.n1580 0.0380882
R52276 ASIG5V.n1582 ASIG5V.n1581 0.0380882
R52277 ASIG5V.n1582 ASIG5V.n1443 0.0380882
R52278 ASIG5V.n1589 ASIG5V.n1443 0.0380882
R52279 ASIG5V.n1590 ASIG5V.n1589 0.0380882
R52280 ASIG5V.n1591 ASIG5V.n1590 0.0380882
R52281 ASIG5V.n1591 ASIG5V.n1440 0.0380882
R52282 ASIG5V.n1598 ASIG5V.n1440 0.0380882
R52283 ASIG5V.n1599 ASIG5V.n1598 0.0380882
R52284 ASIG5V.n1600 ASIG5V.n1599 0.0380882
R52285 ASIG5V.n1600 ASIG5V.n1437 0.0380882
R52286 ASIG5V.n1607 ASIG5V.n1437 0.0380882
R52287 ASIG5V.n1608 ASIG5V.n1607 0.0380882
R52288 ASIG5V.n1609 ASIG5V.n1608 0.0380882
R52289 ASIG5V.n1609 ASIG5V.n1434 0.0380882
R52290 ASIG5V.n1616 ASIG5V.n1434 0.0380882
R52291 ASIG5V.n1617 ASIG5V.n1616 0.0380882
R52292 ASIG5V.n1618 ASIG5V.n1617 0.0380882
R52293 ASIG5V.n1618 ASIG5V.n1431 0.0380882
R52294 ASIG5V.n1625 ASIG5V.n1431 0.0380882
R52295 ASIG5V.n1626 ASIG5V.n1625 0.0380882
R52296 ASIG5V.n1627 ASIG5V.n1626 0.0380882
R52297 ASIG5V.n1627 ASIG5V.n1428 0.0380882
R52298 ASIG5V.n1634 ASIG5V.n1428 0.0380882
R52299 ASIG5V.n1635 ASIG5V.n1634 0.0380882
R52300 ASIG5V.n1636 ASIG5V.n1635 0.0380882
R52301 ASIG5V.n1636 ASIG5V.n1425 0.0380882
R52302 ASIG5V.n1643 ASIG5V.n1425 0.0380882
R52303 ASIG5V.n1644 ASIG5V.n1643 0.0380882
R52304 ASIG5V.n1645 ASIG5V.n1644 0.0380882
R52305 ASIG5V.n1645 ASIG5V.n1422 0.0380882
R52306 ASIG5V.n1652 ASIG5V.n1422 0.0380882
R52307 ASIG5V.n1653 ASIG5V.n1652 0.0380882
R52308 ASIG5V.n1654 ASIG5V.n1653 0.0380882
R52309 ASIG5V.n1654 ASIG5V.n1419 0.0380882
R52310 ASIG5V.n1661 ASIG5V.n1419 0.0380882
R52311 ASIG5V.n1662 ASIG5V.n1661 0.0380882
R52312 ASIG5V.n1663 ASIG5V.n1662 0.0380882
R52313 ASIG5V.n1480 ASIG5V.n1372 0.0380882
R52314 ASIG5V.n1480 ASIG5V.n1478 0.0380882
R52315 ASIG5V.n1485 ASIG5V.n1478 0.0380882
R52316 ASIG5V.n1487 ASIG5V.n1485 0.0380882
R52317 ASIG5V.n1489 ASIG5V.n1487 0.0380882
R52318 ASIG5V.n1489 ASIG5V.n1475 0.0380882
R52319 ASIG5V.n1494 ASIG5V.n1475 0.0380882
R52320 ASIG5V.n1496 ASIG5V.n1494 0.0380882
R52321 ASIG5V.n1498 ASIG5V.n1496 0.0380882
R52322 ASIG5V.n1498 ASIG5V.n1472 0.0380882
R52323 ASIG5V.n1503 ASIG5V.n1472 0.0380882
R52324 ASIG5V.n1505 ASIG5V.n1503 0.0380882
R52325 ASIG5V.n1507 ASIG5V.n1505 0.0380882
R52326 ASIG5V.n1507 ASIG5V.n1469 0.0380882
R52327 ASIG5V.n1512 ASIG5V.n1469 0.0380882
R52328 ASIG5V.n1514 ASIG5V.n1512 0.0380882
R52329 ASIG5V.n1516 ASIG5V.n1514 0.0380882
R52330 ASIG5V.n1516 ASIG5V.n1466 0.0380882
R52331 ASIG5V.n1521 ASIG5V.n1466 0.0380882
R52332 ASIG5V.n1523 ASIG5V.n1521 0.0380882
R52333 ASIG5V.n1525 ASIG5V.n1523 0.0380882
R52334 ASIG5V.n1525 ASIG5V.n1463 0.0380882
R52335 ASIG5V.n1530 ASIG5V.n1463 0.0380882
R52336 ASIG5V.n1532 ASIG5V.n1530 0.0380882
R52337 ASIG5V.n1534 ASIG5V.n1532 0.0380882
R52338 ASIG5V.n1534 ASIG5V.n1460 0.0380882
R52339 ASIG5V.n1539 ASIG5V.n1460 0.0380882
R52340 ASIG5V.n1541 ASIG5V.n1539 0.0380882
R52341 ASIG5V.n1543 ASIG5V.n1541 0.0380882
R52342 ASIG5V.n1543 ASIG5V.n1457 0.0380882
R52343 ASIG5V.n1548 ASIG5V.n1457 0.0380882
R52344 ASIG5V.n1550 ASIG5V.n1548 0.0380882
R52345 ASIG5V.n1552 ASIG5V.n1550 0.0380882
R52346 ASIG5V.n1552 ASIG5V.n1454 0.0380882
R52347 ASIG5V.n1557 ASIG5V.n1454 0.0380882
R52348 ASIG5V.n1559 ASIG5V.n1557 0.0380882
R52349 ASIG5V.n1561 ASIG5V.n1559 0.0380882
R52350 ASIG5V.n1561 ASIG5V.n1451 0.0380882
R52351 ASIG5V.n1566 ASIG5V.n1451 0.0380882
R52352 ASIG5V.n1568 ASIG5V.n1566 0.0380882
R52353 ASIG5V.n1570 ASIG5V.n1568 0.0380882
R52354 ASIG5V.n1570 ASIG5V.n1448 0.0380882
R52355 ASIG5V.n1575 ASIG5V.n1448 0.0380882
R52356 ASIG5V.n1577 ASIG5V.n1575 0.0380882
R52357 ASIG5V.n1579 ASIG5V.n1577 0.0380882
R52358 ASIG5V.n1579 ASIG5V.n1445 0.0380882
R52359 ASIG5V.n1584 ASIG5V.n1445 0.0380882
R52360 ASIG5V.n1586 ASIG5V.n1584 0.0380882
R52361 ASIG5V.n1588 ASIG5V.n1586 0.0380882
R52362 ASIG5V.n1588 ASIG5V.n1442 0.0380882
R52363 ASIG5V.n1593 ASIG5V.n1442 0.0380882
R52364 ASIG5V.n1595 ASIG5V.n1593 0.0380882
R52365 ASIG5V.n1597 ASIG5V.n1595 0.0380882
R52366 ASIG5V.n1597 ASIG5V.n1439 0.0380882
R52367 ASIG5V.n1602 ASIG5V.n1439 0.0380882
R52368 ASIG5V.n1604 ASIG5V.n1602 0.0380882
R52369 ASIG5V.n1606 ASIG5V.n1604 0.0380882
R52370 ASIG5V.n1606 ASIG5V.n1436 0.0380882
R52371 ASIG5V.n1611 ASIG5V.n1436 0.0380882
R52372 ASIG5V.n1613 ASIG5V.n1611 0.0380882
R52373 ASIG5V.n1615 ASIG5V.n1613 0.0380882
R52374 ASIG5V.n1615 ASIG5V.n1433 0.0380882
R52375 ASIG5V.n1620 ASIG5V.n1433 0.0380882
R52376 ASIG5V.n1622 ASIG5V.n1620 0.0380882
R52377 ASIG5V.n1624 ASIG5V.n1622 0.0380882
R52378 ASIG5V.n1624 ASIG5V.n1430 0.0380882
R52379 ASIG5V.n1629 ASIG5V.n1430 0.0380882
R52380 ASIG5V.n1631 ASIG5V.n1629 0.0380882
R52381 ASIG5V.n1633 ASIG5V.n1631 0.0380882
R52382 ASIG5V.n1633 ASIG5V.n1427 0.0380882
R52383 ASIG5V.n1638 ASIG5V.n1427 0.0380882
R52384 ASIG5V.n1640 ASIG5V.n1638 0.0380882
R52385 ASIG5V.n1642 ASIG5V.n1640 0.0380882
R52386 ASIG5V.n1642 ASIG5V.n1424 0.0380882
R52387 ASIG5V.n1647 ASIG5V.n1424 0.0380882
R52388 ASIG5V.n1649 ASIG5V.n1647 0.0380882
R52389 ASIG5V.n1651 ASIG5V.n1649 0.0380882
R52390 ASIG5V.n1651 ASIG5V.n1421 0.0380882
R52391 ASIG5V.n1656 ASIG5V.n1421 0.0380882
R52392 ASIG5V.n1658 ASIG5V.n1656 0.0380882
R52393 ASIG5V.n1660 ASIG5V.n1658 0.0380882
R52394 ASIG5V.n1660 ASIG5V.n1418 0.0380882
R52395 ASIG5V.n12006 ASIG5V.n1418 0.0380882
R52396 ASIG5V.n11809 ASIG5V.n11807 0.0380882
R52397 ASIG5V.n11810 ASIG5V.n11809 0.0380882
R52398 ASIG5V.n11811 ASIG5V.n11810 0.0380882
R52399 ASIG5V.n11811 ASIG5V.n1823 0.0380882
R52400 ASIG5V.n11818 ASIG5V.n1823 0.0380882
R52401 ASIG5V.n11819 ASIG5V.n11818 0.0380882
R52402 ASIG5V.n11820 ASIG5V.n11819 0.0380882
R52403 ASIG5V.n11820 ASIG5V.n1820 0.0380882
R52404 ASIG5V.n11827 ASIG5V.n1820 0.0380882
R52405 ASIG5V.n11828 ASIG5V.n11827 0.0380882
R52406 ASIG5V.n11829 ASIG5V.n11828 0.0380882
R52407 ASIG5V.n11829 ASIG5V.n1817 0.0380882
R52408 ASIG5V.n11836 ASIG5V.n1817 0.0380882
R52409 ASIG5V.n11837 ASIG5V.n11836 0.0380882
R52410 ASIG5V.n11838 ASIG5V.n11837 0.0380882
R52411 ASIG5V.n11838 ASIG5V.n1814 0.0380882
R52412 ASIG5V.n11845 ASIG5V.n1814 0.0380882
R52413 ASIG5V.n11846 ASIG5V.n11845 0.0380882
R52414 ASIG5V.n11847 ASIG5V.n11846 0.0380882
R52415 ASIG5V.n11847 ASIG5V.n1811 0.0380882
R52416 ASIG5V.n11854 ASIG5V.n1811 0.0380882
R52417 ASIG5V.n11855 ASIG5V.n11854 0.0380882
R52418 ASIG5V.n11856 ASIG5V.n11855 0.0380882
R52419 ASIG5V.n11856 ASIG5V.n1808 0.0380882
R52420 ASIG5V.n11863 ASIG5V.n1808 0.0380882
R52421 ASIG5V.n11864 ASIG5V.n11863 0.0380882
R52422 ASIG5V.n11865 ASIG5V.n11864 0.0380882
R52423 ASIG5V.n11865 ASIG5V.n1805 0.0380882
R52424 ASIG5V.n11872 ASIG5V.n1805 0.0380882
R52425 ASIG5V.n11873 ASIG5V.n11872 0.0380882
R52426 ASIG5V.n11874 ASIG5V.n11873 0.0380882
R52427 ASIG5V.n11874 ASIG5V.n1802 0.0380882
R52428 ASIG5V.n11881 ASIG5V.n1802 0.0380882
R52429 ASIG5V.n11882 ASIG5V.n11881 0.0380882
R52430 ASIG5V.n11883 ASIG5V.n11882 0.0380882
R52431 ASIG5V.n11883 ASIG5V.n1799 0.0380882
R52432 ASIG5V.n11890 ASIG5V.n1799 0.0380882
R52433 ASIG5V.n11891 ASIG5V.n11890 0.0380882
R52434 ASIG5V.n11892 ASIG5V.n11891 0.0380882
R52435 ASIG5V.n11892 ASIG5V.n1796 0.0380882
R52436 ASIG5V.n11899 ASIG5V.n1796 0.0380882
R52437 ASIG5V.n11900 ASIG5V.n11899 0.0380882
R52438 ASIG5V.n11901 ASIG5V.n11900 0.0380882
R52439 ASIG5V.n11901 ASIG5V.n1793 0.0380882
R52440 ASIG5V.n11908 ASIG5V.n1793 0.0380882
R52441 ASIG5V.n11909 ASIG5V.n11908 0.0380882
R52442 ASIG5V.n11910 ASIG5V.n11909 0.0380882
R52443 ASIG5V.n11910 ASIG5V.n1790 0.0380882
R52444 ASIG5V.n11917 ASIG5V.n1790 0.0380882
R52445 ASIG5V.n11918 ASIG5V.n11917 0.0380882
R52446 ASIG5V.n11919 ASIG5V.n11918 0.0380882
R52447 ASIG5V.n11919 ASIG5V.n1787 0.0380882
R52448 ASIG5V.n11926 ASIG5V.n1787 0.0380882
R52449 ASIG5V.n11927 ASIG5V.n11926 0.0380882
R52450 ASIG5V.n11928 ASIG5V.n11927 0.0380882
R52451 ASIG5V.n11928 ASIG5V.n1784 0.0380882
R52452 ASIG5V.n11935 ASIG5V.n1784 0.0380882
R52453 ASIG5V.n11936 ASIG5V.n11935 0.0380882
R52454 ASIG5V.n11937 ASIG5V.n11936 0.0380882
R52455 ASIG5V.n11937 ASIG5V.n1781 0.0380882
R52456 ASIG5V.n11944 ASIG5V.n1781 0.0380882
R52457 ASIG5V.n11945 ASIG5V.n11944 0.0380882
R52458 ASIG5V.n11946 ASIG5V.n11945 0.0380882
R52459 ASIG5V.n11946 ASIG5V.n1778 0.0380882
R52460 ASIG5V.n11953 ASIG5V.n1778 0.0380882
R52461 ASIG5V.n11954 ASIG5V.n11953 0.0380882
R52462 ASIG5V.n11955 ASIG5V.n11954 0.0380882
R52463 ASIG5V.n11955 ASIG5V.n1775 0.0380882
R52464 ASIG5V.n11962 ASIG5V.n1775 0.0380882
R52465 ASIG5V.n11963 ASIG5V.n11962 0.0380882
R52466 ASIG5V.n11964 ASIG5V.n11963 0.0380882
R52467 ASIG5V.n11964 ASIG5V.n1772 0.0380882
R52468 ASIG5V.n11971 ASIG5V.n1772 0.0380882
R52469 ASIG5V.n11972 ASIG5V.n11971 0.0380882
R52470 ASIG5V.n11973 ASIG5V.n11972 0.0380882
R52471 ASIG5V.n11973 ASIG5V.n1769 0.0380882
R52472 ASIG5V.n11980 ASIG5V.n1769 0.0380882
R52473 ASIG5V.n11981 ASIG5V.n11980 0.0380882
R52474 ASIG5V.n11982 ASIG5V.n11981 0.0380882
R52475 ASIG5V.n11982 ASIG5V.n1766 0.0380882
R52476 ASIG5V.n11989 ASIG5V.n1766 0.0380882
R52477 ASIG5V.n11990 ASIG5V.n11989 0.0380882
R52478 ASIG5V.n11991 ASIG5V.n11990 0.0380882
R52479 ASIG5V.n11808 ASIG5V.n1720 0.0380882
R52480 ASIG5V.n11808 ASIG5V.n1825 0.0380882
R52481 ASIG5V.n11813 ASIG5V.n1825 0.0380882
R52482 ASIG5V.n11815 ASIG5V.n11813 0.0380882
R52483 ASIG5V.n11817 ASIG5V.n11815 0.0380882
R52484 ASIG5V.n11817 ASIG5V.n1822 0.0380882
R52485 ASIG5V.n11822 ASIG5V.n1822 0.0380882
R52486 ASIG5V.n11824 ASIG5V.n11822 0.0380882
R52487 ASIG5V.n11826 ASIG5V.n11824 0.0380882
R52488 ASIG5V.n11826 ASIG5V.n1819 0.0380882
R52489 ASIG5V.n11831 ASIG5V.n1819 0.0380882
R52490 ASIG5V.n11833 ASIG5V.n11831 0.0380882
R52491 ASIG5V.n11835 ASIG5V.n11833 0.0380882
R52492 ASIG5V.n11835 ASIG5V.n1816 0.0380882
R52493 ASIG5V.n11840 ASIG5V.n1816 0.0380882
R52494 ASIG5V.n11842 ASIG5V.n11840 0.0380882
R52495 ASIG5V.n11844 ASIG5V.n11842 0.0380882
R52496 ASIG5V.n11844 ASIG5V.n1813 0.0380882
R52497 ASIG5V.n11849 ASIG5V.n1813 0.0380882
R52498 ASIG5V.n11851 ASIG5V.n11849 0.0380882
R52499 ASIG5V.n11853 ASIG5V.n11851 0.0380882
R52500 ASIG5V.n11853 ASIG5V.n1810 0.0380882
R52501 ASIG5V.n11858 ASIG5V.n1810 0.0380882
R52502 ASIG5V.n11860 ASIG5V.n11858 0.0380882
R52503 ASIG5V.n11862 ASIG5V.n11860 0.0380882
R52504 ASIG5V.n11862 ASIG5V.n1807 0.0380882
R52505 ASIG5V.n11867 ASIG5V.n1807 0.0380882
R52506 ASIG5V.n11869 ASIG5V.n11867 0.0380882
R52507 ASIG5V.n11871 ASIG5V.n11869 0.0380882
R52508 ASIG5V.n11871 ASIG5V.n1804 0.0380882
R52509 ASIG5V.n11876 ASIG5V.n1804 0.0380882
R52510 ASIG5V.n11878 ASIG5V.n11876 0.0380882
R52511 ASIG5V.n11880 ASIG5V.n11878 0.0380882
R52512 ASIG5V.n11880 ASIG5V.n1801 0.0380882
R52513 ASIG5V.n11885 ASIG5V.n1801 0.0380882
R52514 ASIG5V.n11887 ASIG5V.n11885 0.0380882
R52515 ASIG5V.n11889 ASIG5V.n11887 0.0380882
R52516 ASIG5V.n11889 ASIG5V.n1798 0.0380882
R52517 ASIG5V.n11894 ASIG5V.n1798 0.0380882
R52518 ASIG5V.n11896 ASIG5V.n11894 0.0380882
R52519 ASIG5V.n11898 ASIG5V.n11896 0.0380882
R52520 ASIG5V.n11898 ASIG5V.n1795 0.0380882
R52521 ASIG5V.n11903 ASIG5V.n1795 0.0380882
R52522 ASIG5V.n11905 ASIG5V.n11903 0.0380882
R52523 ASIG5V.n11907 ASIG5V.n11905 0.0380882
R52524 ASIG5V.n11907 ASIG5V.n1792 0.0380882
R52525 ASIG5V.n11912 ASIG5V.n1792 0.0380882
R52526 ASIG5V.n11914 ASIG5V.n11912 0.0380882
R52527 ASIG5V.n11916 ASIG5V.n11914 0.0380882
R52528 ASIG5V.n11916 ASIG5V.n1789 0.0380882
R52529 ASIG5V.n11921 ASIG5V.n1789 0.0380882
R52530 ASIG5V.n11923 ASIG5V.n11921 0.0380882
R52531 ASIG5V.n11925 ASIG5V.n11923 0.0380882
R52532 ASIG5V.n11925 ASIG5V.n1786 0.0380882
R52533 ASIG5V.n11930 ASIG5V.n1786 0.0380882
R52534 ASIG5V.n11932 ASIG5V.n11930 0.0380882
R52535 ASIG5V.n11934 ASIG5V.n11932 0.0380882
R52536 ASIG5V.n11934 ASIG5V.n1783 0.0380882
R52537 ASIG5V.n11939 ASIG5V.n1783 0.0380882
R52538 ASIG5V.n11941 ASIG5V.n11939 0.0380882
R52539 ASIG5V.n11943 ASIG5V.n11941 0.0380882
R52540 ASIG5V.n11943 ASIG5V.n1780 0.0380882
R52541 ASIG5V.n11948 ASIG5V.n1780 0.0380882
R52542 ASIG5V.n11950 ASIG5V.n11948 0.0380882
R52543 ASIG5V.n11952 ASIG5V.n11950 0.0380882
R52544 ASIG5V.n11952 ASIG5V.n1777 0.0380882
R52545 ASIG5V.n11957 ASIG5V.n1777 0.0380882
R52546 ASIG5V.n11959 ASIG5V.n11957 0.0380882
R52547 ASIG5V.n11961 ASIG5V.n11959 0.0380882
R52548 ASIG5V.n11961 ASIG5V.n1774 0.0380882
R52549 ASIG5V.n11966 ASIG5V.n1774 0.0380882
R52550 ASIG5V.n11968 ASIG5V.n11966 0.0380882
R52551 ASIG5V.n11970 ASIG5V.n11968 0.0380882
R52552 ASIG5V.n11970 ASIG5V.n1771 0.0380882
R52553 ASIG5V.n11975 ASIG5V.n1771 0.0380882
R52554 ASIG5V.n11977 ASIG5V.n11975 0.0380882
R52555 ASIG5V.n11979 ASIG5V.n11977 0.0380882
R52556 ASIG5V.n11979 ASIG5V.n1768 0.0380882
R52557 ASIG5V.n11984 ASIG5V.n1768 0.0380882
R52558 ASIG5V.n11986 ASIG5V.n11984 0.0380882
R52559 ASIG5V.n11988 ASIG5V.n11986 0.0380882
R52560 ASIG5V.n11988 ASIG5V.n1765 0.0380882
R52561 ASIG5V.n11992 ASIG5V.n1765 0.0380882
R52562 ASIG5V.n1952 ASIG5V.n1842 0.0380882
R52563 ASIG5V.n1953 ASIG5V.n1952 0.0380882
R52564 ASIG5V.n1953 ASIG5V.n1947 0.0380882
R52565 ASIG5V.n1963 ASIG5V.n1947 0.0380882
R52566 ASIG5V.n1964 ASIG5V.n1963 0.0380882
R52567 ASIG5V.n1965 ASIG5V.n1964 0.0380882
R52568 ASIG5V.n1965 ASIG5V.n1945 0.0380882
R52569 ASIG5V.n1975 ASIG5V.n1945 0.0380882
R52570 ASIG5V.n1976 ASIG5V.n1975 0.0380882
R52571 ASIG5V.n1977 ASIG5V.n1976 0.0380882
R52572 ASIG5V.n1977 ASIG5V.n1943 0.0380882
R52573 ASIG5V.n1987 ASIG5V.n1943 0.0380882
R52574 ASIG5V.n1988 ASIG5V.n1987 0.0380882
R52575 ASIG5V.n1989 ASIG5V.n1988 0.0380882
R52576 ASIG5V.n1989 ASIG5V.n1941 0.0380882
R52577 ASIG5V.n1999 ASIG5V.n1941 0.0380882
R52578 ASIG5V.n2000 ASIG5V.n1999 0.0380882
R52579 ASIG5V.n2001 ASIG5V.n2000 0.0380882
R52580 ASIG5V.n2001 ASIG5V.n1939 0.0380882
R52581 ASIG5V.n2011 ASIG5V.n1939 0.0380882
R52582 ASIG5V.n2012 ASIG5V.n2011 0.0380882
R52583 ASIG5V.n2013 ASIG5V.n2012 0.0380882
R52584 ASIG5V.n2013 ASIG5V.n1937 0.0380882
R52585 ASIG5V.n2023 ASIG5V.n1937 0.0380882
R52586 ASIG5V.n2024 ASIG5V.n2023 0.0380882
R52587 ASIG5V.n2025 ASIG5V.n2024 0.0380882
R52588 ASIG5V.n2025 ASIG5V.n1935 0.0380882
R52589 ASIG5V.n2035 ASIG5V.n1935 0.0380882
R52590 ASIG5V.n2036 ASIG5V.n2035 0.0380882
R52591 ASIG5V.n2037 ASIG5V.n2036 0.0380882
R52592 ASIG5V.n2037 ASIG5V.n1933 0.0380882
R52593 ASIG5V.n2047 ASIG5V.n1933 0.0380882
R52594 ASIG5V.n2048 ASIG5V.n2047 0.0380882
R52595 ASIG5V.n2049 ASIG5V.n2048 0.0380882
R52596 ASIG5V.n2049 ASIG5V.n1931 0.0380882
R52597 ASIG5V.n2059 ASIG5V.n1931 0.0380882
R52598 ASIG5V.n2060 ASIG5V.n2059 0.0380882
R52599 ASIG5V.n2061 ASIG5V.n2060 0.0380882
R52600 ASIG5V.n2061 ASIG5V.n1929 0.0380882
R52601 ASIG5V.n2071 ASIG5V.n1929 0.0380882
R52602 ASIG5V.n2072 ASIG5V.n2071 0.0380882
R52603 ASIG5V.n2073 ASIG5V.n2072 0.0380882
R52604 ASIG5V.n2073 ASIG5V.n1927 0.0380882
R52605 ASIG5V.n2083 ASIG5V.n1927 0.0380882
R52606 ASIG5V.n2084 ASIG5V.n2083 0.0380882
R52607 ASIG5V.n2085 ASIG5V.n2084 0.0380882
R52608 ASIG5V.n2085 ASIG5V.n1925 0.0380882
R52609 ASIG5V.n2095 ASIG5V.n1925 0.0380882
R52610 ASIG5V.n2096 ASIG5V.n2095 0.0380882
R52611 ASIG5V.n2097 ASIG5V.n2096 0.0380882
R52612 ASIG5V.n2097 ASIG5V.n1923 0.0380882
R52613 ASIG5V.n2107 ASIG5V.n1923 0.0380882
R52614 ASIG5V.n2108 ASIG5V.n2107 0.0380882
R52615 ASIG5V.n2109 ASIG5V.n2108 0.0380882
R52616 ASIG5V.n2109 ASIG5V.n1921 0.0380882
R52617 ASIG5V.n2119 ASIG5V.n1921 0.0380882
R52618 ASIG5V.n2120 ASIG5V.n2119 0.0380882
R52619 ASIG5V.n2121 ASIG5V.n2120 0.0380882
R52620 ASIG5V.n2121 ASIG5V.n1919 0.0380882
R52621 ASIG5V.n2131 ASIG5V.n1919 0.0380882
R52622 ASIG5V.n2132 ASIG5V.n2131 0.0380882
R52623 ASIG5V.n2133 ASIG5V.n2132 0.0380882
R52624 ASIG5V.n2133 ASIG5V.n1917 0.0380882
R52625 ASIG5V.n2143 ASIG5V.n1917 0.0380882
R52626 ASIG5V.n2144 ASIG5V.n2143 0.0380882
R52627 ASIG5V.n2145 ASIG5V.n2144 0.0380882
R52628 ASIG5V.n2145 ASIG5V.n1915 0.0380882
R52629 ASIG5V.n2155 ASIG5V.n1915 0.0380882
R52630 ASIG5V.n2156 ASIG5V.n2155 0.0380882
R52631 ASIG5V.n2157 ASIG5V.n2156 0.0380882
R52632 ASIG5V.n2157 ASIG5V.n1913 0.0380882
R52633 ASIG5V.n2167 ASIG5V.n1913 0.0380882
R52634 ASIG5V.n2168 ASIG5V.n2167 0.0380882
R52635 ASIG5V.n2169 ASIG5V.n2168 0.0380882
R52636 ASIG5V.n2169 ASIG5V.n1911 0.0380882
R52637 ASIG5V.n2179 ASIG5V.n1911 0.0380882
R52638 ASIG5V.n2180 ASIG5V.n2179 0.0380882
R52639 ASIG5V.n2181 ASIG5V.n2180 0.0380882
R52640 ASIG5V.n2181 ASIG5V.n1909 0.0380882
R52641 ASIG5V.n2191 ASIG5V.n1909 0.0380882
R52642 ASIG5V.n2192 ASIG5V.n2191 0.0380882
R52643 ASIG5V.n2193 ASIG5V.n2192 0.0380882
R52644 ASIG5V.n2193 ASIG5V.n1854 0.0380882
R52645 ASIG5V.n1951 ASIG5V.n1948 0.0380882
R52646 ASIG5V.n1954 ASIG5V.n1951 0.0380882
R52647 ASIG5V.n1958 ASIG5V.n1954 0.0380882
R52648 ASIG5V.n1962 ASIG5V.n1958 0.0380882
R52649 ASIG5V.n1962 ASIG5V.n1946 0.0380882
R52650 ASIG5V.n1966 ASIG5V.n1946 0.0380882
R52651 ASIG5V.n1970 ASIG5V.n1966 0.0380882
R52652 ASIG5V.n1974 ASIG5V.n1970 0.0380882
R52653 ASIG5V.n1974 ASIG5V.n1944 0.0380882
R52654 ASIG5V.n1978 ASIG5V.n1944 0.0380882
R52655 ASIG5V.n1982 ASIG5V.n1978 0.0380882
R52656 ASIG5V.n1986 ASIG5V.n1982 0.0380882
R52657 ASIG5V.n1986 ASIG5V.n1942 0.0380882
R52658 ASIG5V.n1990 ASIG5V.n1942 0.0380882
R52659 ASIG5V.n1994 ASIG5V.n1990 0.0380882
R52660 ASIG5V.n1998 ASIG5V.n1994 0.0380882
R52661 ASIG5V.n1998 ASIG5V.n1940 0.0380882
R52662 ASIG5V.n2002 ASIG5V.n1940 0.0380882
R52663 ASIG5V.n2006 ASIG5V.n2002 0.0380882
R52664 ASIG5V.n2010 ASIG5V.n2006 0.0380882
R52665 ASIG5V.n2010 ASIG5V.n1938 0.0380882
R52666 ASIG5V.n2014 ASIG5V.n1938 0.0380882
R52667 ASIG5V.n2018 ASIG5V.n2014 0.0380882
R52668 ASIG5V.n2022 ASIG5V.n2018 0.0380882
R52669 ASIG5V.n2022 ASIG5V.n1936 0.0380882
R52670 ASIG5V.n2026 ASIG5V.n1936 0.0380882
R52671 ASIG5V.n2030 ASIG5V.n2026 0.0380882
R52672 ASIG5V.n2034 ASIG5V.n2030 0.0380882
R52673 ASIG5V.n2034 ASIG5V.n1934 0.0380882
R52674 ASIG5V.n2038 ASIG5V.n1934 0.0380882
R52675 ASIG5V.n2042 ASIG5V.n2038 0.0380882
R52676 ASIG5V.n2046 ASIG5V.n2042 0.0380882
R52677 ASIG5V.n2046 ASIG5V.n1932 0.0380882
R52678 ASIG5V.n2050 ASIG5V.n1932 0.0380882
R52679 ASIG5V.n2054 ASIG5V.n2050 0.0380882
R52680 ASIG5V.n2058 ASIG5V.n2054 0.0380882
R52681 ASIG5V.n2058 ASIG5V.n1930 0.0380882
R52682 ASIG5V.n2062 ASIG5V.n1930 0.0380882
R52683 ASIG5V.n2066 ASIG5V.n2062 0.0380882
R52684 ASIG5V.n2070 ASIG5V.n2066 0.0380882
R52685 ASIG5V.n2070 ASIG5V.n1928 0.0380882
R52686 ASIG5V.n2074 ASIG5V.n1928 0.0380882
R52687 ASIG5V.n2078 ASIG5V.n2074 0.0380882
R52688 ASIG5V.n2082 ASIG5V.n2078 0.0380882
R52689 ASIG5V.n2082 ASIG5V.n1926 0.0380882
R52690 ASIG5V.n2086 ASIG5V.n1926 0.0380882
R52691 ASIG5V.n2090 ASIG5V.n2086 0.0380882
R52692 ASIG5V.n2094 ASIG5V.n2090 0.0380882
R52693 ASIG5V.n2094 ASIG5V.n1924 0.0380882
R52694 ASIG5V.n2098 ASIG5V.n1924 0.0380882
R52695 ASIG5V.n2102 ASIG5V.n2098 0.0380882
R52696 ASIG5V.n2106 ASIG5V.n2102 0.0380882
R52697 ASIG5V.n2106 ASIG5V.n1922 0.0380882
R52698 ASIG5V.n2110 ASIG5V.n1922 0.0380882
R52699 ASIG5V.n2114 ASIG5V.n2110 0.0380882
R52700 ASIG5V.n2118 ASIG5V.n2114 0.0380882
R52701 ASIG5V.n2118 ASIG5V.n1920 0.0380882
R52702 ASIG5V.n2122 ASIG5V.n1920 0.0380882
R52703 ASIG5V.n2126 ASIG5V.n2122 0.0380882
R52704 ASIG5V.n2130 ASIG5V.n2126 0.0380882
R52705 ASIG5V.n2130 ASIG5V.n1918 0.0380882
R52706 ASIG5V.n2134 ASIG5V.n1918 0.0380882
R52707 ASIG5V.n2138 ASIG5V.n2134 0.0380882
R52708 ASIG5V.n2142 ASIG5V.n2138 0.0380882
R52709 ASIG5V.n2142 ASIG5V.n1916 0.0380882
R52710 ASIG5V.n2146 ASIG5V.n1916 0.0380882
R52711 ASIG5V.n2150 ASIG5V.n2146 0.0380882
R52712 ASIG5V.n2154 ASIG5V.n2150 0.0380882
R52713 ASIG5V.n2154 ASIG5V.n1914 0.0380882
R52714 ASIG5V.n2158 ASIG5V.n1914 0.0380882
R52715 ASIG5V.n2162 ASIG5V.n2158 0.0380882
R52716 ASIG5V.n2166 ASIG5V.n2162 0.0380882
R52717 ASIG5V.n2166 ASIG5V.n1912 0.0380882
R52718 ASIG5V.n2170 ASIG5V.n1912 0.0380882
R52719 ASIG5V.n2174 ASIG5V.n2170 0.0380882
R52720 ASIG5V.n2178 ASIG5V.n2174 0.0380882
R52721 ASIG5V.n2178 ASIG5V.n1910 0.0380882
R52722 ASIG5V.n2182 ASIG5V.n1910 0.0380882
R52723 ASIG5V.n2186 ASIG5V.n2182 0.0380882
R52724 ASIG5V.n2190 ASIG5V.n2186 0.0380882
R52725 ASIG5V.n2190 ASIG5V.n1908 0.0380882
R52726 ASIG5V.n2194 ASIG5V.n1908 0.0380882
R52727 ASIG5V.n2194 ASIG5V.n1907 0.0380882
R52728 ASIG5V.n2309 ASIG5V.n2218 0.0380882
R52729 ASIG5V.n2310 ASIG5V.n2309 0.0380882
R52730 ASIG5V.n2310 ASIG5V.n2304 0.0380882
R52731 ASIG5V.n2320 ASIG5V.n2304 0.0380882
R52732 ASIG5V.n2321 ASIG5V.n2320 0.0380882
R52733 ASIG5V.n2322 ASIG5V.n2321 0.0380882
R52734 ASIG5V.n2322 ASIG5V.n2302 0.0380882
R52735 ASIG5V.n2332 ASIG5V.n2302 0.0380882
R52736 ASIG5V.n2333 ASIG5V.n2332 0.0380882
R52737 ASIG5V.n2334 ASIG5V.n2333 0.0380882
R52738 ASIG5V.n2334 ASIG5V.n2300 0.0380882
R52739 ASIG5V.n2344 ASIG5V.n2300 0.0380882
R52740 ASIG5V.n2345 ASIG5V.n2344 0.0380882
R52741 ASIG5V.n2346 ASIG5V.n2345 0.0380882
R52742 ASIG5V.n2346 ASIG5V.n2298 0.0380882
R52743 ASIG5V.n2356 ASIG5V.n2298 0.0380882
R52744 ASIG5V.n2357 ASIG5V.n2356 0.0380882
R52745 ASIG5V.n2358 ASIG5V.n2357 0.0380882
R52746 ASIG5V.n2358 ASIG5V.n2296 0.0380882
R52747 ASIG5V.n2368 ASIG5V.n2296 0.0380882
R52748 ASIG5V.n2369 ASIG5V.n2368 0.0380882
R52749 ASIG5V.n2370 ASIG5V.n2369 0.0380882
R52750 ASIG5V.n2370 ASIG5V.n2294 0.0380882
R52751 ASIG5V.n2380 ASIG5V.n2294 0.0380882
R52752 ASIG5V.n2381 ASIG5V.n2380 0.0380882
R52753 ASIG5V.n2382 ASIG5V.n2381 0.0380882
R52754 ASIG5V.n2382 ASIG5V.n2292 0.0380882
R52755 ASIG5V.n2392 ASIG5V.n2292 0.0380882
R52756 ASIG5V.n2393 ASIG5V.n2392 0.0380882
R52757 ASIG5V.n2394 ASIG5V.n2393 0.0380882
R52758 ASIG5V.n2394 ASIG5V.n2290 0.0380882
R52759 ASIG5V.n2404 ASIG5V.n2290 0.0380882
R52760 ASIG5V.n2405 ASIG5V.n2404 0.0380882
R52761 ASIG5V.n2406 ASIG5V.n2405 0.0380882
R52762 ASIG5V.n2406 ASIG5V.n2288 0.0380882
R52763 ASIG5V.n2416 ASIG5V.n2288 0.0380882
R52764 ASIG5V.n2417 ASIG5V.n2416 0.0380882
R52765 ASIG5V.n2418 ASIG5V.n2417 0.0380882
R52766 ASIG5V.n2418 ASIG5V.n2286 0.0380882
R52767 ASIG5V.n2428 ASIG5V.n2286 0.0380882
R52768 ASIG5V.n2429 ASIG5V.n2428 0.0380882
R52769 ASIG5V.n2430 ASIG5V.n2429 0.0380882
R52770 ASIG5V.n2430 ASIG5V.n2284 0.0380882
R52771 ASIG5V.n2440 ASIG5V.n2284 0.0380882
R52772 ASIG5V.n2441 ASIG5V.n2440 0.0380882
R52773 ASIG5V.n2442 ASIG5V.n2441 0.0380882
R52774 ASIG5V.n2442 ASIG5V.n2282 0.0380882
R52775 ASIG5V.n2452 ASIG5V.n2282 0.0380882
R52776 ASIG5V.n2453 ASIG5V.n2452 0.0380882
R52777 ASIG5V.n2454 ASIG5V.n2453 0.0380882
R52778 ASIG5V.n2454 ASIG5V.n2280 0.0380882
R52779 ASIG5V.n2464 ASIG5V.n2280 0.0380882
R52780 ASIG5V.n2465 ASIG5V.n2464 0.0380882
R52781 ASIG5V.n2466 ASIG5V.n2465 0.0380882
R52782 ASIG5V.n2466 ASIG5V.n2278 0.0380882
R52783 ASIG5V.n2476 ASIG5V.n2278 0.0380882
R52784 ASIG5V.n2477 ASIG5V.n2476 0.0380882
R52785 ASIG5V.n2478 ASIG5V.n2477 0.0380882
R52786 ASIG5V.n2478 ASIG5V.n2276 0.0380882
R52787 ASIG5V.n2488 ASIG5V.n2276 0.0380882
R52788 ASIG5V.n2489 ASIG5V.n2488 0.0380882
R52789 ASIG5V.n2490 ASIG5V.n2489 0.0380882
R52790 ASIG5V.n2490 ASIG5V.n2274 0.0380882
R52791 ASIG5V.n2500 ASIG5V.n2274 0.0380882
R52792 ASIG5V.n2501 ASIG5V.n2500 0.0380882
R52793 ASIG5V.n2502 ASIG5V.n2501 0.0380882
R52794 ASIG5V.n2502 ASIG5V.n2272 0.0380882
R52795 ASIG5V.n2512 ASIG5V.n2272 0.0380882
R52796 ASIG5V.n2513 ASIG5V.n2512 0.0380882
R52797 ASIG5V.n2514 ASIG5V.n2513 0.0380882
R52798 ASIG5V.n2514 ASIG5V.n2270 0.0380882
R52799 ASIG5V.n2524 ASIG5V.n2270 0.0380882
R52800 ASIG5V.n2525 ASIG5V.n2524 0.0380882
R52801 ASIG5V.n2526 ASIG5V.n2525 0.0380882
R52802 ASIG5V.n2526 ASIG5V.n2268 0.0380882
R52803 ASIG5V.n2536 ASIG5V.n2268 0.0380882
R52804 ASIG5V.n2537 ASIG5V.n2536 0.0380882
R52805 ASIG5V.n2538 ASIG5V.n2537 0.0380882
R52806 ASIG5V.n2538 ASIG5V.n2266 0.0380882
R52807 ASIG5V.n2548 ASIG5V.n2266 0.0380882
R52808 ASIG5V.n2549 ASIG5V.n2548 0.0380882
R52809 ASIG5V.n2550 ASIG5V.n2549 0.0380882
R52810 ASIG5V.n2550 ASIG5V.n2206 0.0380882
R52811 ASIG5V.n2308 ASIG5V.n2305 0.0380882
R52812 ASIG5V.n2311 ASIG5V.n2308 0.0380882
R52813 ASIG5V.n2315 ASIG5V.n2311 0.0380882
R52814 ASIG5V.n2319 ASIG5V.n2315 0.0380882
R52815 ASIG5V.n2319 ASIG5V.n2303 0.0380882
R52816 ASIG5V.n2323 ASIG5V.n2303 0.0380882
R52817 ASIG5V.n2327 ASIG5V.n2323 0.0380882
R52818 ASIG5V.n2331 ASIG5V.n2327 0.0380882
R52819 ASIG5V.n2331 ASIG5V.n2301 0.0380882
R52820 ASIG5V.n2335 ASIG5V.n2301 0.0380882
R52821 ASIG5V.n2339 ASIG5V.n2335 0.0380882
R52822 ASIG5V.n2343 ASIG5V.n2339 0.0380882
R52823 ASIG5V.n2343 ASIG5V.n2299 0.0380882
R52824 ASIG5V.n2347 ASIG5V.n2299 0.0380882
R52825 ASIG5V.n2351 ASIG5V.n2347 0.0380882
R52826 ASIG5V.n2355 ASIG5V.n2351 0.0380882
R52827 ASIG5V.n2355 ASIG5V.n2297 0.0380882
R52828 ASIG5V.n2359 ASIG5V.n2297 0.0380882
R52829 ASIG5V.n2363 ASIG5V.n2359 0.0380882
R52830 ASIG5V.n2367 ASIG5V.n2363 0.0380882
R52831 ASIG5V.n2367 ASIG5V.n2295 0.0380882
R52832 ASIG5V.n2371 ASIG5V.n2295 0.0380882
R52833 ASIG5V.n2375 ASIG5V.n2371 0.0380882
R52834 ASIG5V.n2379 ASIG5V.n2375 0.0380882
R52835 ASIG5V.n2379 ASIG5V.n2293 0.0380882
R52836 ASIG5V.n2383 ASIG5V.n2293 0.0380882
R52837 ASIG5V.n2387 ASIG5V.n2383 0.0380882
R52838 ASIG5V.n2391 ASIG5V.n2387 0.0380882
R52839 ASIG5V.n2391 ASIG5V.n2291 0.0380882
R52840 ASIG5V.n2395 ASIG5V.n2291 0.0380882
R52841 ASIG5V.n2399 ASIG5V.n2395 0.0380882
R52842 ASIG5V.n2403 ASIG5V.n2399 0.0380882
R52843 ASIG5V.n2403 ASIG5V.n2289 0.0380882
R52844 ASIG5V.n2407 ASIG5V.n2289 0.0380882
R52845 ASIG5V.n2411 ASIG5V.n2407 0.0380882
R52846 ASIG5V.n2415 ASIG5V.n2411 0.0380882
R52847 ASIG5V.n2415 ASIG5V.n2287 0.0380882
R52848 ASIG5V.n2419 ASIG5V.n2287 0.0380882
R52849 ASIG5V.n2423 ASIG5V.n2419 0.0380882
R52850 ASIG5V.n2427 ASIG5V.n2423 0.0380882
R52851 ASIG5V.n2427 ASIG5V.n2285 0.0380882
R52852 ASIG5V.n2431 ASIG5V.n2285 0.0380882
R52853 ASIG5V.n2435 ASIG5V.n2431 0.0380882
R52854 ASIG5V.n2439 ASIG5V.n2435 0.0380882
R52855 ASIG5V.n2439 ASIG5V.n2283 0.0380882
R52856 ASIG5V.n2443 ASIG5V.n2283 0.0380882
R52857 ASIG5V.n2447 ASIG5V.n2443 0.0380882
R52858 ASIG5V.n2451 ASIG5V.n2447 0.0380882
R52859 ASIG5V.n2451 ASIG5V.n2281 0.0380882
R52860 ASIG5V.n2455 ASIG5V.n2281 0.0380882
R52861 ASIG5V.n2459 ASIG5V.n2455 0.0380882
R52862 ASIG5V.n2463 ASIG5V.n2459 0.0380882
R52863 ASIG5V.n2463 ASIG5V.n2279 0.0380882
R52864 ASIG5V.n2467 ASIG5V.n2279 0.0380882
R52865 ASIG5V.n2471 ASIG5V.n2467 0.0380882
R52866 ASIG5V.n2475 ASIG5V.n2471 0.0380882
R52867 ASIG5V.n2475 ASIG5V.n2277 0.0380882
R52868 ASIG5V.n2479 ASIG5V.n2277 0.0380882
R52869 ASIG5V.n2483 ASIG5V.n2479 0.0380882
R52870 ASIG5V.n2487 ASIG5V.n2483 0.0380882
R52871 ASIG5V.n2487 ASIG5V.n2275 0.0380882
R52872 ASIG5V.n2491 ASIG5V.n2275 0.0380882
R52873 ASIG5V.n2495 ASIG5V.n2491 0.0380882
R52874 ASIG5V.n2499 ASIG5V.n2495 0.0380882
R52875 ASIG5V.n2499 ASIG5V.n2273 0.0380882
R52876 ASIG5V.n2503 ASIG5V.n2273 0.0380882
R52877 ASIG5V.n2507 ASIG5V.n2503 0.0380882
R52878 ASIG5V.n2511 ASIG5V.n2507 0.0380882
R52879 ASIG5V.n2511 ASIG5V.n2271 0.0380882
R52880 ASIG5V.n2515 ASIG5V.n2271 0.0380882
R52881 ASIG5V.n2519 ASIG5V.n2515 0.0380882
R52882 ASIG5V.n2523 ASIG5V.n2519 0.0380882
R52883 ASIG5V.n2523 ASIG5V.n2269 0.0380882
R52884 ASIG5V.n2527 ASIG5V.n2269 0.0380882
R52885 ASIG5V.n2531 ASIG5V.n2527 0.0380882
R52886 ASIG5V.n2535 ASIG5V.n2531 0.0380882
R52887 ASIG5V.n2535 ASIG5V.n2267 0.0380882
R52888 ASIG5V.n2539 ASIG5V.n2267 0.0380882
R52889 ASIG5V.n2543 ASIG5V.n2539 0.0380882
R52890 ASIG5V.n2547 ASIG5V.n2543 0.0380882
R52891 ASIG5V.n2547 ASIG5V.n2265 0.0380882
R52892 ASIG5V.n2551 ASIG5V.n2265 0.0380882
R52893 ASIG5V.n2551 ASIG5V.n2264 0.0380882
R52894 ASIG5V.n2661 ASIG5V.n2563 0.0380882
R52895 ASIG5V.n2662 ASIG5V.n2661 0.0380882
R52896 ASIG5V.n2662 ASIG5V.n2656 0.0380882
R52897 ASIG5V.n2672 ASIG5V.n2656 0.0380882
R52898 ASIG5V.n2673 ASIG5V.n2672 0.0380882
R52899 ASIG5V.n2674 ASIG5V.n2673 0.0380882
R52900 ASIG5V.n2674 ASIG5V.n2654 0.0380882
R52901 ASIG5V.n2684 ASIG5V.n2654 0.0380882
R52902 ASIG5V.n2685 ASIG5V.n2684 0.0380882
R52903 ASIG5V.n2686 ASIG5V.n2685 0.0380882
R52904 ASIG5V.n2686 ASIG5V.n2652 0.0380882
R52905 ASIG5V.n2696 ASIG5V.n2652 0.0380882
R52906 ASIG5V.n2697 ASIG5V.n2696 0.0380882
R52907 ASIG5V.n2698 ASIG5V.n2697 0.0380882
R52908 ASIG5V.n2698 ASIG5V.n2650 0.0380882
R52909 ASIG5V.n2708 ASIG5V.n2650 0.0380882
R52910 ASIG5V.n2709 ASIG5V.n2708 0.0380882
R52911 ASIG5V.n2710 ASIG5V.n2709 0.0380882
R52912 ASIG5V.n2710 ASIG5V.n2648 0.0380882
R52913 ASIG5V.n2720 ASIG5V.n2648 0.0380882
R52914 ASIG5V.n2721 ASIG5V.n2720 0.0380882
R52915 ASIG5V.n2722 ASIG5V.n2721 0.0380882
R52916 ASIG5V.n2722 ASIG5V.n2646 0.0380882
R52917 ASIG5V.n2732 ASIG5V.n2646 0.0380882
R52918 ASIG5V.n2733 ASIG5V.n2732 0.0380882
R52919 ASIG5V.n2734 ASIG5V.n2733 0.0380882
R52920 ASIG5V.n2734 ASIG5V.n2644 0.0380882
R52921 ASIG5V.n2744 ASIG5V.n2644 0.0380882
R52922 ASIG5V.n2745 ASIG5V.n2744 0.0380882
R52923 ASIG5V.n2746 ASIG5V.n2745 0.0380882
R52924 ASIG5V.n2746 ASIG5V.n2642 0.0380882
R52925 ASIG5V.n2756 ASIG5V.n2642 0.0380882
R52926 ASIG5V.n2757 ASIG5V.n2756 0.0380882
R52927 ASIG5V.n2758 ASIG5V.n2757 0.0380882
R52928 ASIG5V.n2758 ASIG5V.n2640 0.0380882
R52929 ASIG5V.n2768 ASIG5V.n2640 0.0380882
R52930 ASIG5V.n2769 ASIG5V.n2768 0.0380882
R52931 ASIG5V.n2770 ASIG5V.n2769 0.0380882
R52932 ASIG5V.n2770 ASIG5V.n2638 0.0380882
R52933 ASIG5V.n2780 ASIG5V.n2638 0.0380882
R52934 ASIG5V.n2781 ASIG5V.n2780 0.0380882
R52935 ASIG5V.n2782 ASIG5V.n2781 0.0380882
R52936 ASIG5V.n2782 ASIG5V.n2636 0.0380882
R52937 ASIG5V.n2792 ASIG5V.n2636 0.0380882
R52938 ASIG5V.n2793 ASIG5V.n2792 0.0380882
R52939 ASIG5V.n2794 ASIG5V.n2793 0.0380882
R52940 ASIG5V.n2794 ASIG5V.n2634 0.0380882
R52941 ASIG5V.n2804 ASIG5V.n2634 0.0380882
R52942 ASIG5V.n2805 ASIG5V.n2804 0.0380882
R52943 ASIG5V.n2806 ASIG5V.n2805 0.0380882
R52944 ASIG5V.n2806 ASIG5V.n2632 0.0380882
R52945 ASIG5V.n2816 ASIG5V.n2632 0.0380882
R52946 ASIG5V.n2817 ASIG5V.n2816 0.0380882
R52947 ASIG5V.n2818 ASIG5V.n2817 0.0380882
R52948 ASIG5V.n2818 ASIG5V.n2630 0.0380882
R52949 ASIG5V.n2828 ASIG5V.n2630 0.0380882
R52950 ASIG5V.n2829 ASIG5V.n2828 0.0380882
R52951 ASIG5V.n2830 ASIG5V.n2829 0.0380882
R52952 ASIG5V.n2830 ASIG5V.n2628 0.0380882
R52953 ASIG5V.n2840 ASIG5V.n2628 0.0380882
R52954 ASIG5V.n2841 ASIG5V.n2840 0.0380882
R52955 ASIG5V.n2842 ASIG5V.n2841 0.0380882
R52956 ASIG5V.n2842 ASIG5V.n2626 0.0380882
R52957 ASIG5V.n2852 ASIG5V.n2626 0.0380882
R52958 ASIG5V.n2853 ASIG5V.n2852 0.0380882
R52959 ASIG5V.n2854 ASIG5V.n2853 0.0380882
R52960 ASIG5V.n2854 ASIG5V.n2624 0.0380882
R52961 ASIG5V.n2864 ASIG5V.n2624 0.0380882
R52962 ASIG5V.n2865 ASIG5V.n2864 0.0380882
R52963 ASIG5V.n2866 ASIG5V.n2865 0.0380882
R52964 ASIG5V.n2866 ASIG5V.n2622 0.0380882
R52965 ASIG5V.n2876 ASIG5V.n2622 0.0380882
R52966 ASIG5V.n2877 ASIG5V.n2876 0.0380882
R52967 ASIG5V.n2878 ASIG5V.n2877 0.0380882
R52968 ASIG5V.n2878 ASIG5V.n2620 0.0380882
R52969 ASIG5V.n2888 ASIG5V.n2620 0.0380882
R52970 ASIG5V.n2889 ASIG5V.n2888 0.0380882
R52971 ASIG5V.n2890 ASIG5V.n2889 0.0380882
R52972 ASIG5V.n2890 ASIG5V.n2618 0.0380882
R52973 ASIG5V.n2900 ASIG5V.n2618 0.0380882
R52974 ASIG5V.n2901 ASIG5V.n2900 0.0380882
R52975 ASIG5V.n11766 ASIG5V.n2901 0.0380882
R52976 ASIG5V.n11766 ASIG5V.n11765 0.0380882
R52977 ASIG5V.n2660 ASIG5V.n2657 0.0380882
R52978 ASIG5V.n2663 ASIG5V.n2660 0.0380882
R52979 ASIG5V.n2667 ASIG5V.n2663 0.0380882
R52980 ASIG5V.n2671 ASIG5V.n2667 0.0380882
R52981 ASIG5V.n2671 ASIG5V.n2655 0.0380882
R52982 ASIG5V.n2675 ASIG5V.n2655 0.0380882
R52983 ASIG5V.n2679 ASIG5V.n2675 0.0380882
R52984 ASIG5V.n2683 ASIG5V.n2679 0.0380882
R52985 ASIG5V.n2683 ASIG5V.n2653 0.0380882
R52986 ASIG5V.n2687 ASIG5V.n2653 0.0380882
R52987 ASIG5V.n2691 ASIG5V.n2687 0.0380882
R52988 ASIG5V.n2695 ASIG5V.n2691 0.0380882
R52989 ASIG5V.n2695 ASIG5V.n2651 0.0380882
R52990 ASIG5V.n2699 ASIG5V.n2651 0.0380882
R52991 ASIG5V.n2703 ASIG5V.n2699 0.0380882
R52992 ASIG5V.n2707 ASIG5V.n2703 0.0380882
R52993 ASIG5V.n2707 ASIG5V.n2649 0.0380882
R52994 ASIG5V.n2711 ASIG5V.n2649 0.0380882
R52995 ASIG5V.n2715 ASIG5V.n2711 0.0380882
R52996 ASIG5V.n2719 ASIG5V.n2715 0.0380882
R52997 ASIG5V.n2719 ASIG5V.n2647 0.0380882
R52998 ASIG5V.n2723 ASIG5V.n2647 0.0380882
R52999 ASIG5V.n2727 ASIG5V.n2723 0.0380882
R53000 ASIG5V.n2731 ASIG5V.n2727 0.0380882
R53001 ASIG5V.n2731 ASIG5V.n2645 0.0380882
R53002 ASIG5V.n2735 ASIG5V.n2645 0.0380882
R53003 ASIG5V.n2739 ASIG5V.n2735 0.0380882
R53004 ASIG5V.n2743 ASIG5V.n2739 0.0380882
R53005 ASIG5V.n2743 ASIG5V.n2643 0.0380882
R53006 ASIG5V.n2747 ASIG5V.n2643 0.0380882
R53007 ASIG5V.n2751 ASIG5V.n2747 0.0380882
R53008 ASIG5V.n2755 ASIG5V.n2751 0.0380882
R53009 ASIG5V.n2755 ASIG5V.n2641 0.0380882
R53010 ASIG5V.n2759 ASIG5V.n2641 0.0380882
R53011 ASIG5V.n2763 ASIG5V.n2759 0.0380882
R53012 ASIG5V.n2767 ASIG5V.n2763 0.0380882
R53013 ASIG5V.n2767 ASIG5V.n2639 0.0380882
R53014 ASIG5V.n2771 ASIG5V.n2639 0.0380882
R53015 ASIG5V.n2775 ASIG5V.n2771 0.0380882
R53016 ASIG5V.n2779 ASIG5V.n2775 0.0380882
R53017 ASIG5V.n2779 ASIG5V.n2637 0.0380882
R53018 ASIG5V.n2783 ASIG5V.n2637 0.0380882
R53019 ASIG5V.n2787 ASIG5V.n2783 0.0380882
R53020 ASIG5V.n2791 ASIG5V.n2787 0.0380882
R53021 ASIG5V.n2791 ASIG5V.n2635 0.0380882
R53022 ASIG5V.n2795 ASIG5V.n2635 0.0380882
R53023 ASIG5V.n2799 ASIG5V.n2795 0.0380882
R53024 ASIG5V.n2803 ASIG5V.n2799 0.0380882
R53025 ASIG5V.n2803 ASIG5V.n2633 0.0380882
R53026 ASIG5V.n2807 ASIG5V.n2633 0.0380882
R53027 ASIG5V.n2811 ASIG5V.n2807 0.0380882
R53028 ASIG5V.n2815 ASIG5V.n2811 0.0380882
R53029 ASIG5V.n2815 ASIG5V.n2631 0.0380882
R53030 ASIG5V.n2819 ASIG5V.n2631 0.0380882
R53031 ASIG5V.n2823 ASIG5V.n2819 0.0380882
R53032 ASIG5V.n2827 ASIG5V.n2823 0.0380882
R53033 ASIG5V.n2827 ASIG5V.n2629 0.0380882
R53034 ASIG5V.n2831 ASIG5V.n2629 0.0380882
R53035 ASIG5V.n2835 ASIG5V.n2831 0.0380882
R53036 ASIG5V.n2839 ASIG5V.n2835 0.0380882
R53037 ASIG5V.n2839 ASIG5V.n2627 0.0380882
R53038 ASIG5V.n2843 ASIG5V.n2627 0.0380882
R53039 ASIG5V.n2847 ASIG5V.n2843 0.0380882
R53040 ASIG5V.n2851 ASIG5V.n2847 0.0380882
R53041 ASIG5V.n2851 ASIG5V.n2625 0.0380882
R53042 ASIG5V.n2855 ASIG5V.n2625 0.0380882
R53043 ASIG5V.n2859 ASIG5V.n2855 0.0380882
R53044 ASIG5V.n2863 ASIG5V.n2859 0.0380882
R53045 ASIG5V.n2863 ASIG5V.n2623 0.0380882
R53046 ASIG5V.n2867 ASIG5V.n2623 0.0380882
R53047 ASIG5V.n2871 ASIG5V.n2867 0.0380882
R53048 ASIG5V.n2875 ASIG5V.n2871 0.0380882
R53049 ASIG5V.n2875 ASIG5V.n2621 0.0380882
R53050 ASIG5V.n2879 ASIG5V.n2621 0.0380882
R53051 ASIG5V.n2883 ASIG5V.n2879 0.0380882
R53052 ASIG5V.n2887 ASIG5V.n2883 0.0380882
R53053 ASIG5V.n2887 ASIG5V.n2619 0.0380882
R53054 ASIG5V.n2891 ASIG5V.n2619 0.0380882
R53055 ASIG5V.n2895 ASIG5V.n2891 0.0380882
R53056 ASIG5V.n2899 ASIG5V.n2895 0.0380882
R53057 ASIG5V.n2899 ASIG5V.n2617 0.0380882
R53058 ASIG5V.n11767 ASIG5V.n2617 0.0380882
R53059 ASIG5V.n11767 ASIG5V.n2614 0.0380882
R53060 ASIG5V.n11505 ASIG5V.n11504 0.0380882
R53061 ASIG5V.n11506 ASIG5V.n11505 0.0380882
R53062 ASIG5V.n11506 ASIG5V.n2998 0.0380882
R53063 ASIG5V.n11516 ASIG5V.n2998 0.0380882
R53064 ASIG5V.n11517 ASIG5V.n11516 0.0380882
R53065 ASIG5V.n11518 ASIG5V.n11517 0.0380882
R53066 ASIG5V.n11518 ASIG5V.n2996 0.0380882
R53067 ASIG5V.n11528 ASIG5V.n2996 0.0380882
R53068 ASIG5V.n11529 ASIG5V.n11528 0.0380882
R53069 ASIG5V.n11530 ASIG5V.n11529 0.0380882
R53070 ASIG5V.n11530 ASIG5V.n2994 0.0380882
R53071 ASIG5V.n11540 ASIG5V.n2994 0.0380882
R53072 ASIG5V.n11541 ASIG5V.n11540 0.0380882
R53073 ASIG5V.n11542 ASIG5V.n11541 0.0380882
R53074 ASIG5V.n11542 ASIG5V.n2992 0.0380882
R53075 ASIG5V.n11552 ASIG5V.n2992 0.0380882
R53076 ASIG5V.n11553 ASIG5V.n11552 0.0380882
R53077 ASIG5V.n11554 ASIG5V.n11553 0.0380882
R53078 ASIG5V.n11554 ASIG5V.n2990 0.0380882
R53079 ASIG5V.n11564 ASIG5V.n2990 0.0380882
R53080 ASIG5V.n11565 ASIG5V.n11564 0.0380882
R53081 ASIG5V.n11566 ASIG5V.n11565 0.0380882
R53082 ASIG5V.n11566 ASIG5V.n2988 0.0380882
R53083 ASIG5V.n11576 ASIG5V.n2988 0.0380882
R53084 ASIG5V.n11577 ASIG5V.n11576 0.0380882
R53085 ASIG5V.n11578 ASIG5V.n11577 0.0380882
R53086 ASIG5V.n11578 ASIG5V.n2986 0.0380882
R53087 ASIG5V.n11588 ASIG5V.n2986 0.0380882
R53088 ASIG5V.n11589 ASIG5V.n11588 0.0380882
R53089 ASIG5V.n11590 ASIG5V.n11589 0.0380882
R53090 ASIG5V.n11590 ASIG5V.n2984 0.0380882
R53091 ASIG5V.n11600 ASIG5V.n2984 0.0380882
R53092 ASIG5V.n11601 ASIG5V.n11600 0.0380882
R53093 ASIG5V.n11602 ASIG5V.n11601 0.0380882
R53094 ASIG5V.n11602 ASIG5V.n2982 0.0380882
R53095 ASIG5V.n11612 ASIG5V.n2982 0.0380882
R53096 ASIG5V.n11613 ASIG5V.n11612 0.0380882
R53097 ASIG5V.n11614 ASIG5V.n11613 0.0380882
R53098 ASIG5V.n11614 ASIG5V.n2980 0.0380882
R53099 ASIG5V.n11624 ASIG5V.n2980 0.0380882
R53100 ASIG5V.n11625 ASIG5V.n11624 0.0380882
R53101 ASIG5V.n11626 ASIG5V.n11625 0.0380882
R53102 ASIG5V.n11626 ASIG5V.n2978 0.0380882
R53103 ASIG5V.n11636 ASIG5V.n2978 0.0380882
R53104 ASIG5V.n11637 ASIG5V.n11636 0.0380882
R53105 ASIG5V.n11638 ASIG5V.n11637 0.0380882
R53106 ASIG5V.n11638 ASIG5V.n2976 0.0380882
R53107 ASIG5V.n11648 ASIG5V.n2976 0.0380882
R53108 ASIG5V.n11649 ASIG5V.n11648 0.0380882
R53109 ASIG5V.n11650 ASIG5V.n11649 0.0380882
R53110 ASIG5V.n11650 ASIG5V.n2974 0.0380882
R53111 ASIG5V.n11660 ASIG5V.n2974 0.0380882
R53112 ASIG5V.n11661 ASIG5V.n11660 0.0380882
R53113 ASIG5V.n11662 ASIG5V.n11661 0.0380882
R53114 ASIG5V.n11662 ASIG5V.n2972 0.0380882
R53115 ASIG5V.n11672 ASIG5V.n2972 0.0380882
R53116 ASIG5V.n11673 ASIG5V.n11672 0.0380882
R53117 ASIG5V.n11674 ASIG5V.n11673 0.0380882
R53118 ASIG5V.n11674 ASIG5V.n2970 0.0380882
R53119 ASIG5V.n11684 ASIG5V.n2970 0.0380882
R53120 ASIG5V.n11685 ASIG5V.n11684 0.0380882
R53121 ASIG5V.n11686 ASIG5V.n11685 0.0380882
R53122 ASIG5V.n11686 ASIG5V.n2968 0.0380882
R53123 ASIG5V.n11696 ASIG5V.n2968 0.0380882
R53124 ASIG5V.n11697 ASIG5V.n11696 0.0380882
R53125 ASIG5V.n11698 ASIG5V.n11697 0.0380882
R53126 ASIG5V.n11698 ASIG5V.n2966 0.0380882
R53127 ASIG5V.n11708 ASIG5V.n2966 0.0380882
R53128 ASIG5V.n11709 ASIG5V.n11708 0.0380882
R53129 ASIG5V.n11710 ASIG5V.n11709 0.0380882
R53130 ASIG5V.n11710 ASIG5V.n2964 0.0380882
R53131 ASIG5V.n11720 ASIG5V.n2964 0.0380882
R53132 ASIG5V.n11721 ASIG5V.n11720 0.0380882
R53133 ASIG5V.n11722 ASIG5V.n11721 0.0380882
R53134 ASIG5V.n11722 ASIG5V.n2962 0.0380882
R53135 ASIG5V.n11732 ASIG5V.n2962 0.0380882
R53136 ASIG5V.n11733 ASIG5V.n11732 0.0380882
R53137 ASIG5V.n11734 ASIG5V.n11733 0.0380882
R53138 ASIG5V.n11734 ASIG5V.n2960 0.0380882
R53139 ASIG5V.n11744 ASIG5V.n2960 0.0380882
R53140 ASIG5V.n11745 ASIG5V.n11744 0.0380882
R53141 ASIG5V.n11746 ASIG5V.n11745 0.0380882
R53142 ASIG5V.n11746 ASIG5V.n2909 0.0380882
R53143 ASIG5V.n11503 ASIG5V.n3001 0.0380882
R53144 ASIG5V.n11507 ASIG5V.n3001 0.0380882
R53145 ASIG5V.n11511 ASIG5V.n11507 0.0380882
R53146 ASIG5V.n11515 ASIG5V.n11511 0.0380882
R53147 ASIG5V.n11515 ASIG5V.n2997 0.0380882
R53148 ASIG5V.n11519 ASIG5V.n2997 0.0380882
R53149 ASIG5V.n11523 ASIG5V.n11519 0.0380882
R53150 ASIG5V.n11527 ASIG5V.n11523 0.0380882
R53151 ASIG5V.n11527 ASIG5V.n2995 0.0380882
R53152 ASIG5V.n11531 ASIG5V.n2995 0.0380882
R53153 ASIG5V.n11535 ASIG5V.n11531 0.0380882
R53154 ASIG5V.n11539 ASIG5V.n11535 0.0380882
R53155 ASIG5V.n11539 ASIG5V.n2993 0.0380882
R53156 ASIG5V.n11543 ASIG5V.n2993 0.0380882
R53157 ASIG5V.n11547 ASIG5V.n11543 0.0380882
R53158 ASIG5V.n11551 ASIG5V.n11547 0.0380882
R53159 ASIG5V.n11551 ASIG5V.n2991 0.0380882
R53160 ASIG5V.n11555 ASIG5V.n2991 0.0380882
R53161 ASIG5V.n11559 ASIG5V.n11555 0.0380882
R53162 ASIG5V.n11563 ASIG5V.n11559 0.0380882
R53163 ASIG5V.n11563 ASIG5V.n2989 0.0380882
R53164 ASIG5V.n11567 ASIG5V.n2989 0.0380882
R53165 ASIG5V.n11571 ASIG5V.n11567 0.0380882
R53166 ASIG5V.n11575 ASIG5V.n11571 0.0380882
R53167 ASIG5V.n11575 ASIG5V.n2987 0.0380882
R53168 ASIG5V.n11579 ASIG5V.n2987 0.0380882
R53169 ASIG5V.n11583 ASIG5V.n11579 0.0380882
R53170 ASIG5V.n11587 ASIG5V.n11583 0.0380882
R53171 ASIG5V.n11587 ASIG5V.n2985 0.0380882
R53172 ASIG5V.n11591 ASIG5V.n2985 0.0380882
R53173 ASIG5V.n11595 ASIG5V.n11591 0.0380882
R53174 ASIG5V.n11599 ASIG5V.n11595 0.0380882
R53175 ASIG5V.n11599 ASIG5V.n2983 0.0380882
R53176 ASIG5V.n11603 ASIG5V.n2983 0.0380882
R53177 ASIG5V.n11607 ASIG5V.n11603 0.0380882
R53178 ASIG5V.n11611 ASIG5V.n11607 0.0380882
R53179 ASIG5V.n11611 ASIG5V.n2981 0.0380882
R53180 ASIG5V.n11615 ASIG5V.n2981 0.0380882
R53181 ASIG5V.n11619 ASIG5V.n11615 0.0380882
R53182 ASIG5V.n11623 ASIG5V.n11619 0.0380882
R53183 ASIG5V.n11623 ASIG5V.n2979 0.0380882
R53184 ASIG5V.n11627 ASIG5V.n2979 0.0380882
R53185 ASIG5V.n11631 ASIG5V.n11627 0.0380882
R53186 ASIG5V.n11635 ASIG5V.n11631 0.0380882
R53187 ASIG5V.n11635 ASIG5V.n2977 0.0380882
R53188 ASIG5V.n11639 ASIG5V.n2977 0.0380882
R53189 ASIG5V.n11643 ASIG5V.n11639 0.0380882
R53190 ASIG5V.n11647 ASIG5V.n11643 0.0380882
R53191 ASIG5V.n11647 ASIG5V.n2975 0.0380882
R53192 ASIG5V.n11651 ASIG5V.n2975 0.0380882
R53193 ASIG5V.n11655 ASIG5V.n11651 0.0380882
R53194 ASIG5V.n11659 ASIG5V.n11655 0.0380882
R53195 ASIG5V.n11659 ASIG5V.n2973 0.0380882
R53196 ASIG5V.n11663 ASIG5V.n2973 0.0380882
R53197 ASIG5V.n11667 ASIG5V.n11663 0.0380882
R53198 ASIG5V.n11671 ASIG5V.n11667 0.0380882
R53199 ASIG5V.n11671 ASIG5V.n2971 0.0380882
R53200 ASIG5V.n11675 ASIG5V.n2971 0.0380882
R53201 ASIG5V.n11679 ASIG5V.n11675 0.0380882
R53202 ASIG5V.n11683 ASIG5V.n11679 0.0380882
R53203 ASIG5V.n11683 ASIG5V.n2969 0.0380882
R53204 ASIG5V.n11687 ASIG5V.n2969 0.0380882
R53205 ASIG5V.n11691 ASIG5V.n11687 0.0380882
R53206 ASIG5V.n11695 ASIG5V.n11691 0.0380882
R53207 ASIG5V.n11695 ASIG5V.n2967 0.0380882
R53208 ASIG5V.n11699 ASIG5V.n2967 0.0380882
R53209 ASIG5V.n11703 ASIG5V.n11699 0.0380882
R53210 ASIG5V.n11707 ASIG5V.n11703 0.0380882
R53211 ASIG5V.n11707 ASIG5V.n2965 0.0380882
R53212 ASIG5V.n11711 ASIG5V.n2965 0.0380882
R53213 ASIG5V.n11715 ASIG5V.n11711 0.0380882
R53214 ASIG5V.n11719 ASIG5V.n11715 0.0380882
R53215 ASIG5V.n11719 ASIG5V.n2963 0.0380882
R53216 ASIG5V.n11723 ASIG5V.n2963 0.0380882
R53217 ASIG5V.n11727 ASIG5V.n11723 0.0380882
R53218 ASIG5V.n11731 ASIG5V.n11727 0.0380882
R53219 ASIG5V.n11731 ASIG5V.n2961 0.0380882
R53220 ASIG5V.n11735 ASIG5V.n2961 0.0380882
R53221 ASIG5V.n11739 ASIG5V.n11735 0.0380882
R53222 ASIG5V.n11743 ASIG5V.n11739 0.0380882
R53223 ASIG5V.n11743 ASIG5V.n2959 0.0380882
R53224 ASIG5V.n11747 ASIG5V.n2959 0.0380882
R53225 ASIG5V.n11747 ASIG5V.n2957 0.0380882
R53226 ASIG5V.n11239 ASIG5V.n11238 0.0380882
R53227 ASIG5V.n11240 ASIG5V.n11239 0.0380882
R53228 ASIG5V.n11240 ASIG5V.n11233 0.0380882
R53229 ASIG5V.n11250 ASIG5V.n11233 0.0380882
R53230 ASIG5V.n11251 ASIG5V.n11250 0.0380882
R53231 ASIG5V.n11252 ASIG5V.n11251 0.0380882
R53232 ASIG5V.n11252 ASIG5V.n11231 0.0380882
R53233 ASIG5V.n11262 ASIG5V.n11231 0.0380882
R53234 ASIG5V.n11263 ASIG5V.n11262 0.0380882
R53235 ASIG5V.n11264 ASIG5V.n11263 0.0380882
R53236 ASIG5V.n11264 ASIG5V.n11229 0.0380882
R53237 ASIG5V.n11274 ASIG5V.n11229 0.0380882
R53238 ASIG5V.n11275 ASIG5V.n11274 0.0380882
R53239 ASIG5V.n11276 ASIG5V.n11275 0.0380882
R53240 ASIG5V.n11276 ASIG5V.n11227 0.0380882
R53241 ASIG5V.n11286 ASIG5V.n11227 0.0380882
R53242 ASIG5V.n11287 ASIG5V.n11286 0.0380882
R53243 ASIG5V.n11288 ASIG5V.n11287 0.0380882
R53244 ASIG5V.n11288 ASIG5V.n11225 0.0380882
R53245 ASIG5V.n11298 ASIG5V.n11225 0.0380882
R53246 ASIG5V.n11299 ASIG5V.n11298 0.0380882
R53247 ASIG5V.n11300 ASIG5V.n11299 0.0380882
R53248 ASIG5V.n11300 ASIG5V.n11223 0.0380882
R53249 ASIG5V.n11310 ASIG5V.n11223 0.0380882
R53250 ASIG5V.n11311 ASIG5V.n11310 0.0380882
R53251 ASIG5V.n11312 ASIG5V.n11311 0.0380882
R53252 ASIG5V.n11312 ASIG5V.n11221 0.0380882
R53253 ASIG5V.n11322 ASIG5V.n11221 0.0380882
R53254 ASIG5V.n11323 ASIG5V.n11322 0.0380882
R53255 ASIG5V.n11324 ASIG5V.n11323 0.0380882
R53256 ASIG5V.n11324 ASIG5V.n11219 0.0380882
R53257 ASIG5V.n11334 ASIG5V.n11219 0.0380882
R53258 ASIG5V.n11335 ASIG5V.n11334 0.0380882
R53259 ASIG5V.n11336 ASIG5V.n11335 0.0380882
R53260 ASIG5V.n11336 ASIG5V.n11217 0.0380882
R53261 ASIG5V.n11346 ASIG5V.n11217 0.0380882
R53262 ASIG5V.n11347 ASIG5V.n11346 0.0380882
R53263 ASIG5V.n11348 ASIG5V.n11347 0.0380882
R53264 ASIG5V.n11348 ASIG5V.n11215 0.0380882
R53265 ASIG5V.n11358 ASIG5V.n11215 0.0380882
R53266 ASIG5V.n11359 ASIG5V.n11358 0.0380882
R53267 ASIG5V.n11360 ASIG5V.n11359 0.0380882
R53268 ASIG5V.n11360 ASIG5V.n11213 0.0380882
R53269 ASIG5V.n11370 ASIG5V.n11213 0.0380882
R53270 ASIG5V.n11371 ASIG5V.n11370 0.0380882
R53271 ASIG5V.n11372 ASIG5V.n11371 0.0380882
R53272 ASIG5V.n11372 ASIG5V.n11211 0.0380882
R53273 ASIG5V.n11382 ASIG5V.n11211 0.0380882
R53274 ASIG5V.n11383 ASIG5V.n11382 0.0380882
R53275 ASIG5V.n11384 ASIG5V.n11383 0.0380882
R53276 ASIG5V.n11384 ASIG5V.n11209 0.0380882
R53277 ASIG5V.n11394 ASIG5V.n11209 0.0380882
R53278 ASIG5V.n11395 ASIG5V.n11394 0.0380882
R53279 ASIG5V.n11396 ASIG5V.n11395 0.0380882
R53280 ASIG5V.n11396 ASIG5V.n11207 0.0380882
R53281 ASIG5V.n11406 ASIG5V.n11207 0.0380882
R53282 ASIG5V.n11407 ASIG5V.n11406 0.0380882
R53283 ASIG5V.n11408 ASIG5V.n11407 0.0380882
R53284 ASIG5V.n11408 ASIG5V.n11205 0.0380882
R53285 ASIG5V.n11418 ASIG5V.n11205 0.0380882
R53286 ASIG5V.n11419 ASIG5V.n11418 0.0380882
R53287 ASIG5V.n11420 ASIG5V.n11419 0.0380882
R53288 ASIG5V.n11420 ASIG5V.n11203 0.0380882
R53289 ASIG5V.n11430 ASIG5V.n11203 0.0380882
R53290 ASIG5V.n11431 ASIG5V.n11430 0.0380882
R53291 ASIG5V.n11432 ASIG5V.n11431 0.0380882
R53292 ASIG5V.n11432 ASIG5V.n11201 0.0380882
R53293 ASIG5V.n11442 ASIG5V.n11201 0.0380882
R53294 ASIG5V.n11443 ASIG5V.n11442 0.0380882
R53295 ASIG5V.n11444 ASIG5V.n11443 0.0380882
R53296 ASIG5V.n11444 ASIG5V.n11199 0.0380882
R53297 ASIG5V.n11454 ASIG5V.n11199 0.0380882
R53298 ASIG5V.n11455 ASIG5V.n11454 0.0380882
R53299 ASIG5V.n11456 ASIG5V.n11455 0.0380882
R53300 ASIG5V.n11456 ASIG5V.n11197 0.0380882
R53301 ASIG5V.n11466 ASIG5V.n11197 0.0380882
R53302 ASIG5V.n11467 ASIG5V.n11466 0.0380882
R53303 ASIG5V.n11468 ASIG5V.n11467 0.0380882
R53304 ASIG5V.n11468 ASIG5V.n11195 0.0380882
R53305 ASIG5V.n11478 ASIG5V.n11195 0.0380882
R53306 ASIG5V.n11479 ASIG5V.n11478 0.0380882
R53307 ASIG5V.n11480 ASIG5V.n11479 0.0380882
R53308 ASIG5V.n11480 ASIG5V.n9969 0.0380882
R53309 ASIG5V.n11237 ASIG5V.n11236 0.0380882
R53310 ASIG5V.n11241 ASIG5V.n11236 0.0380882
R53311 ASIG5V.n11245 ASIG5V.n11241 0.0380882
R53312 ASIG5V.n11249 ASIG5V.n11245 0.0380882
R53313 ASIG5V.n11249 ASIG5V.n11232 0.0380882
R53314 ASIG5V.n11253 ASIG5V.n11232 0.0380882
R53315 ASIG5V.n11257 ASIG5V.n11253 0.0380882
R53316 ASIG5V.n11261 ASIG5V.n11257 0.0380882
R53317 ASIG5V.n11261 ASIG5V.n11230 0.0380882
R53318 ASIG5V.n11265 ASIG5V.n11230 0.0380882
R53319 ASIG5V.n11269 ASIG5V.n11265 0.0380882
R53320 ASIG5V.n11273 ASIG5V.n11269 0.0380882
R53321 ASIG5V.n11273 ASIG5V.n11228 0.0380882
R53322 ASIG5V.n11277 ASIG5V.n11228 0.0380882
R53323 ASIG5V.n11281 ASIG5V.n11277 0.0380882
R53324 ASIG5V.n11285 ASIG5V.n11281 0.0380882
R53325 ASIG5V.n11285 ASIG5V.n11226 0.0380882
R53326 ASIG5V.n11289 ASIG5V.n11226 0.0380882
R53327 ASIG5V.n11293 ASIG5V.n11289 0.0380882
R53328 ASIG5V.n11297 ASIG5V.n11293 0.0380882
R53329 ASIG5V.n11297 ASIG5V.n11224 0.0380882
R53330 ASIG5V.n11301 ASIG5V.n11224 0.0380882
R53331 ASIG5V.n11305 ASIG5V.n11301 0.0380882
R53332 ASIG5V.n11309 ASIG5V.n11305 0.0380882
R53333 ASIG5V.n11309 ASIG5V.n11222 0.0380882
R53334 ASIG5V.n11313 ASIG5V.n11222 0.0380882
R53335 ASIG5V.n11317 ASIG5V.n11313 0.0380882
R53336 ASIG5V.n11321 ASIG5V.n11317 0.0380882
R53337 ASIG5V.n11321 ASIG5V.n11220 0.0380882
R53338 ASIG5V.n11325 ASIG5V.n11220 0.0380882
R53339 ASIG5V.n11329 ASIG5V.n11325 0.0380882
R53340 ASIG5V.n11333 ASIG5V.n11329 0.0380882
R53341 ASIG5V.n11333 ASIG5V.n11218 0.0380882
R53342 ASIG5V.n11337 ASIG5V.n11218 0.0380882
R53343 ASIG5V.n11341 ASIG5V.n11337 0.0380882
R53344 ASIG5V.n11345 ASIG5V.n11341 0.0380882
R53345 ASIG5V.n11345 ASIG5V.n11216 0.0380882
R53346 ASIG5V.n11349 ASIG5V.n11216 0.0380882
R53347 ASIG5V.n11353 ASIG5V.n11349 0.0380882
R53348 ASIG5V.n11357 ASIG5V.n11353 0.0380882
R53349 ASIG5V.n11357 ASIG5V.n11214 0.0380882
R53350 ASIG5V.n11361 ASIG5V.n11214 0.0380882
R53351 ASIG5V.n11365 ASIG5V.n11361 0.0380882
R53352 ASIG5V.n11369 ASIG5V.n11365 0.0380882
R53353 ASIG5V.n11369 ASIG5V.n11212 0.0380882
R53354 ASIG5V.n11373 ASIG5V.n11212 0.0380882
R53355 ASIG5V.n11377 ASIG5V.n11373 0.0380882
R53356 ASIG5V.n11381 ASIG5V.n11377 0.0380882
R53357 ASIG5V.n11381 ASIG5V.n11210 0.0380882
R53358 ASIG5V.n11385 ASIG5V.n11210 0.0380882
R53359 ASIG5V.n11389 ASIG5V.n11385 0.0380882
R53360 ASIG5V.n11393 ASIG5V.n11389 0.0380882
R53361 ASIG5V.n11393 ASIG5V.n11208 0.0380882
R53362 ASIG5V.n11397 ASIG5V.n11208 0.0380882
R53363 ASIG5V.n11401 ASIG5V.n11397 0.0380882
R53364 ASIG5V.n11405 ASIG5V.n11401 0.0380882
R53365 ASIG5V.n11405 ASIG5V.n11206 0.0380882
R53366 ASIG5V.n11409 ASIG5V.n11206 0.0380882
R53367 ASIG5V.n11413 ASIG5V.n11409 0.0380882
R53368 ASIG5V.n11417 ASIG5V.n11413 0.0380882
R53369 ASIG5V.n11417 ASIG5V.n11204 0.0380882
R53370 ASIG5V.n11421 ASIG5V.n11204 0.0380882
R53371 ASIG5V.n11425 ASIG5V.n11421 0.0380882
R53372 ASIG5V.n11429 ASIG5V.n11425 0.0380882
R53373 ASIG5V.n11429 ASIG5V.n11202 0.0380882
R53374 ASIG5V.n11433 ASIG5V.n11202 0.0380882
R53375 ASIG5V.n11437 ASIG5V.n11433 0.0380882
R53376 ASIG5V.n11441 ASIG5V.n11437 0.0380882
R53377 ASIG5V.n11441 ASIG5V.n11200 0.0380882
R53378 ASIG5V.n11445 ASIG5V.n11200 0.0380882
R53379 ASIG5V.n11449 ASIG5V.n11445 0.0380882
R53380 ASIG5V.n11453 ASIG5V.n11449 0.0380882
R53381 ASIG5V.n11453 ASIG5V.n11198 0.0380882
R53382 ASIG5V.n11457 ASIG5V.n11198 0.0380882
R53383 ASIG5V.n11461 ASIG5V.n11457 0.0380882
R53384 ASIG5V.n11465 ASIG5V.n11461 0.0380882
R53385 ASIG5V.n11465 ASIG5V.n11196 0.0380882
R53386 ASIG5V.n11469 ASIG5V.n11196 0.0380882
R53387 ASIG5V.n11473 ASIG5V.n11469 0.0380882
R53388 ASIG5V.n11477 ASIG5V.n11473 0.0380882
R53389 ASIG5V.n11477 ASIG5V.n11194 0.0380882
R53390 ASIG5V.n11481 ASIG5V.n11194 0.0380882
R53391 ASIG5V.n11481 ASIG5V.n11193 0.0380882
R53392 ASIG5V.n4586 ASIG5V.n4585 0.0380882
R53393 ASIG5V.n4587 ASIG5V.n4586 0.0380882
R53394 ASIG5V.n4587 ASIG5V.n3775 0.0380882
R53395 ASIG5V.n4594 ASIG5V.n3775 0.0380882
R53396 ASIG5V.n4595 ASIG5V.n4594 0.0380882
R53397 ASIG5V.n4596 ASIG5V.n4595 0.0380882
R53398 ASIG5V.n4596 ASIG5V.n3772 0.0380882
R53399 ASIG5V.n4603 ASIG5V.n3772 0.0380882
R53400 ASIG5V.n4604 ASIG5V.n4603 0.0380882
R53401 ASIG5V.n4605 ASIG5V.n4604 0.0380882
R53402 ASIG5V.n4605 ASIG5V.n3769 0.0380882
R53403 ASIG5V.n4612 ASIG5V.n3769 0.0380882
R53404 ASIG5V.n4613 ASIG5V.n4612 0.0380882
R53405 ASIG5V.n4614 ASIG5V.n4613 0.0380882
R53406 ASIG5V.n4614 ASIG5V.n3766 0.0380882
R53407 ASIG5V.n4621 ASIG5V.n3766 0.0380882
R53408 ASIG5V.n4622 ASIG5V.n4621 0.0380882
R53409 ASIG5V.n4623 ASIG5V.n4622 0.0380882
R53410 ASIG5V.n4623 ASIG5V.n3763 0.0380882
R53411 ASIG5V.n4630 ASIG5V.n3763 0.0380882
R53412 ASIG5V.n4631 ASIG5V.n4630 0.0380882
R53413 ASIG5V.n4632 ASIG5V.n4631 0.0380882
R53414 ASIG5V.n4632 ASIG5V.n3760 0.0380882
R53415 ASIG5V.n4639 ASIG5V.n3760 0.0380882
R53416 ASIG5V.n4640 ASIG5V.n4639 0.0380882
R53417 ASIG5V.n4641 ASIG5V.n4640 0.0380882
R53418 ASIG5V.n4641 ASIG5V.n3757 0.0380882
R53419 ASIG5V.n4648 ASIG5V.n3757 0.0380882
R53420 ASIG5V.n4649 ASIG5V.n4648 0.0380882
R53421 ASIG5V.n4650 ASIG5V.n4649 0.0380882
R53422 ASIG5V.n4650 ASIG5V.n3754 0.0380882
R53423 ASIG5V.n4657 ASIG5V.n3754 0.0380882
R53424 ASIG5V.n4658 ASIG5V.n4657 0.0380882
R53425 ASIG5V.n4659 ASIG5V.n4658 0.0380882
R53426 ASIG5V.n4659 ASIG5V.n3751 0.0380882
R53427 ASIG5V.n4666 ASIG5V.n3751 0.0380882
R53428 ASIG5V.n4667 ASIG5V.n4666 0.0380882
R53429 ASIG5V.n4668 ASIG5V.n4667 0.0380882
R53430 ASIG5V.n4668 ASIG5V.n3748 0.0380882
R53431 ASIG5V.n4675 ASIG5V.n3748 0.0380882
R53432 ASIG5V.n4676 ASIG5V.n4675 0.0380882
R53433 ASIG5V.n4677 ASIG5V.n4676 0.0380882
R53434 ASIG5V.n4677 ASIG5V.n3745 0.0380882
R53435 ASIG5V.n4684 ASIG5V.n3745 0.0380882
R53436 ASIG5V.n4685 ASIG5V.n4684 0.0380882
R53437 ASIG5V.n4686 ASIG5V.n4685 0.0380882
R53438 ASIG5V.n4686 ASIG5V.n3742 0.0380882
R53439 ASIG5V.n4693 ASIG5V.n3742 0.0380882
R53440 ASIG5V.n4694 ASIG5V.n4693 0.0380882
R53441 ASIG5V.n4695 ASIG5V.n4694 0.0380882
R53442 ASIG5V.n4695 ASIG5V.n3739 0.0380882
R53443 ASIG5V.n4702 ASIG5V.n3739 0.0380882
R53444 ASIG5V.n4703 ASIG5V.n4702 0.0380882
R53445 ASIG5V.n4704 ASIG5V.n4703 0.0380882
R53446 ASIG5V.n4704 ASIG5V.n3736 0.0380882
R53447 ASIG5V.n4711 ASIG5V.n3736 0.0380882
R53448 ASIG5V.n4712 ASIG5V.n4711 0.0380882
R53449 ASIG5V.n4713 ASIG5V.n4712 0.0380882
R53450 ASIG5V.n4713 ASIG5V.n3733 0.0380882
R53451 ASIG5V.n4720 ASIG5V.n3733 0.0380882
R53452 ASIG5V.n4721 ASIG5V.n4720 0.0380882
R53453 ASIG5V.n4722 ASIG5V.n4721 0.0380882
R53454 ASIG5V.n4722 ASIG5V.n3730 0.0380882
R53455 ASIG5V.n4729 ASIG5V.n3730 0.0380882
R53456 ASIG5V.n4730 ASIG5V.n4729 0.0380882
R53457 ASIG5V.n4731 ASIG5V.n4730 0.0380882
R53458 ASIG5V.n4731 ASIG5V.n3727 0.0380882
R53459 ASIG5V.n4738 ASIG5V.n3727 0.0380882
R53460 ASIG5V.n4739 ASIG5V.n4738 0.0380882
R53461 ASIG5V.n4740 ASIG5V.n4739 0.0380882
R53462 ASIG5V.n4740 ASIG5V.n3724 0.0380882
R53463 ASIG5V.n4747 ASIG5V.n3724 0.0380882
R53464 ASIG5V.n4748 ASIG5V.n4747 0.0380882
R53465 ASIG5V.n4749 ASIG5V.n4748 0.0380882
R53466 ASIG5V.n4749 ASIG5V.n3721 0.0380882
R53467 ASIG5V.n4756 ASIG5V.n3721 0.0380882
R53468 ASIG5V.n4757 ASIG5V.n4756 0.0380882
R53469 ASIG5V.n4758 ASIG5V.n4757 0.0380882
R53470 ASIG5V.n4758 ASIG5V.n3718 0.0380882
R53471 ASIG5V.n4765 ASIG5V.n3718 0.0380882
R53472 ASIG5V.n4766 ASIG5V.n4765 0.0380882
R53473 ASIG5V.n4767 ASIG5V.n4766 0.0380882
R53474 ASIG5V.n4767 ASIG5V.n3623 0.0380882
R53475 ASIG5V.n3776 ASIG5V.n3673 0.0380882
R53476 ASIG5V.n4589 ASIG5V.n3776 0.0380882
R53477 ASIG5V.n4591 ASIG5V.n4589 0.0380882
R53478 ASIG5V.n4593 ASIG5V.n4591 0.0380882
R53479 ASIG5V.n4593 ASIG5V.n3774 0.0380882
R53480 ASIG5V.n4598 ASIG5V.n3774 0.0380882
R53481 ASIG5V.n4600 ASIG5V.n4598 0.0380882
R53482 ASIG5V.n4602 ASIG5V.n4600 0.0380882
R53483 ASIG5V.n4602 ASIG5V.n3771 0.0380882
R53484 ASIG5V.n4607 ASIG5V.n3771 0.0380882
R53485 ASIG5V.n4609 ASIG5V.n4607 0.0380882
R53486 ASIG5V.n4611 ASIG5V.n4609 0.0380882
R53487 ASIG5V.n4611 ASIG5V.n3768 0.0380882
R53488 ASIG5V.n4616 ASIG5V.n3768 0.0380882
R53489 ASIG5V.n4618 ASIG5V.n4616 0.0380882
R53490 ASIG5V.n4620 ASIG5V.n4618 0.0380882
R53491 ASIG5V.n4620 ASIG5V.n3765 0.0380882
R53492 ASIG5V.n4625 ASIG5V.n3765 0.0380882
R53493 ASIG5V.n4627 ASIG5V.n4625 0.0380882
R53494 ASIG5V.n4629 ASIG5V.n4627 0.0380882
R53495 ASIG5V.n4629 ASIG5V.n3762 0.0380882
R53496 ASIG5V.n4634 ASIG5V.n3762 0.0380882
R53497 ASIG5V.n4636 ASIG5V.n4634 0.0380882
R53498 ASIG5V.n4638 ASIG5V.n4636 0.0380882
R53499 ASIG5V.n4638 ASIG5V.n3759 0.0380882
R53500 ASIG5V.n4643 ASIG5V.n3759 0.0380882
R53501 ASIG5V.n4645 ASIG5V.n4643 0.0380882
R53502 ASIG5V.n4647 ASIG5V.n4645 0.0380882
R53503 ASIG5V.n4647 ASIG5V.n3756 0.0380882
R53504 ASIG5V.n4652 ASIG5V.n3756 0.0380882
R53505 ASIG5V.n4654 ASIG5V.n4652 0.0380882
R53506 ASIG5V.n4656 ASIG5V.n4654 0.0380882
R53507 ASIG5V.n4656 ASIG5V.n3753 0.0380882
R53508 ASIG5V.n4661 ASIG5V.n3753 0.0380882
R53509 ASIG5V.n4663 ASIG5V.n4661 0.0380882
R53510 ASIG5V.n4665 ASIG5V.n4663 0.0380882
R53511 ASIG5V.n4665 ASIG5V.n3750 0.0380882
R53512 ASIG5V.n4670 ASIG5V.n3750 0.0380882
R53513 ASIG5V.n4672 ASIG5V.n4670 0.0380882
R53514 ASIG5V.n4674 ASIG5V.n4672 0.0380882
R53515 ASIG5V.n4674 ASIG5V.n3747 0.0380882
R53516 ASIG5V.n4679 ASIG5V.n3747 0.0380882
R53517 ASIG5V.n4681 ASIG5V.n4679 0.0380882
R53518 ASIG5V.n4683 ASIG5V.n4681 0.0380882
R53519 ASIG5V.n4683 ASIG5V.n3744 0.0380882
R53520 ASIG5V.n4688 ASIG5V.n3744 0.0380882
R53521 ASIG5V.n4690 ASIG5V.n4688 0.0380882
R53522 ASIG5V.n4692 ASIG5V.n4690 0.0380882
R53523 ASIG5V.n4692 ASIG5V.n3741 0.0380882
R53524 ASIG5V.n4697 ASIG5V.n3741 0.0380882
R53525 ASIG5V.n4699 ASIG5V.n4697 0.0380882
R53526 ASIG5V.n4701 ASIG5V.n4699 0.0380882
R53527 ASIG5V.n4701 ASIG5V.n3738 0.0380882
R53528 ASIG5V.n4706 ASIG5V.n3738 0.0380882
R53529 ASIG5V.n4708 ASIG5V.n4706 0.0380882
R53530 ASIG5V.n4710 ASIG5V.n4708 0.0380882
R53531 ASIG5V.n4710 ASIG5V.n3735 0.0380882
R53532 ASIG5V.n4715 ASIG5V.n3735 0.0380882
R53533 ASIG5V.n4717 ASIG5V.n4715 0.0380882
R53534 ASIG5V.n4719 ASIG5V.n4717 0.0380882
R53535 ASIG5V.n4719 ASIG5V.n3732 0.0380882
R53536 ASIG5V.n4724 ASIG5V.n3732 0.0380882
R53537 ASIG5V.n4726 ASIG5V.n4724 0.0380882
R53538 ASIG5V.n4728 ASIG5V.n4726 0.0380882
R53539 ASIG5V.n4728 ASIG5V.n3729 0.0380882
R53540 ASIG5V.n4733 ASIG5V.n3729 0.0380882
R53541 ASIG5V.n4735 ASIG5V.n4733 0.0380882
R53542 ASIG5V.n4737 ASIG5V.n4735 0.0380882
R53543 ASIG5V.n4737 ASIG5V.n3726 0.0380882
R53544 ASIG5V.n4742 ASIG5V.n3726 0.0380882
R53545 ASIG5V.n4744 ASIG5V.n4742 0.0380882
R53546 ASIG5V.n4746 ASIG5V.n4744 0.0380882
R53547 ASIG5V.n4746 ASIG5V.n3723 0.0380882
R53548 ASIG5V.n4751 ASIG5V.n3723 0.0380882
R53549 ASIG5V.n4753 ASIG5V.n4751 0.0380882
R53550 ASIG5V.n4755 ASIG5V.n4753 0.0380882
R53551 ASIG5V.n4755 ASIG5V.n3720 0.0380882
R53552 ASIG5V.n4760 ASIG5V.n3720 0.0380882
R53553 ASIG5V.n4762 ASIG5V.n4760 0.0380882
R53554 ASIG5V.n4764 ASIG5V.n4762 0.0380882
R53555 ASIG5V.n4764 ASIG5V.n3717 0.0380882
R53556 ASIG5V.n4769 ASIG5V.n3717 0.0380882
R53557 ASIG5V.n4770 ASIG5V.n4769 0.0380882
R53558 ASIG5V.n4551 ASIG5V.n4309 0.0380882
R53559 ASIG5V.n4551 ASIG5V.n4311 0.0380882
R53560 ASIG5V.n4547 ASIG5V.n4311 0.0380882
R53561 ASIG5V.n4547 ASIG5V.n4545 0.0380882
R53562 ASIG5V.n4545 ASIG5V.n4543 0.0380882
R53563 ASIG5V.n4543 ASIG5V.n4314 0.0380882
R53564 ASIG5V.n4539 ASIG5V.n4314 0.0380882
R53565 ASIG5V.n4539 ASIG5V.n4537 0.0380882
R53566 ASIG5V.n4537 ASIG5V.n4535 0.0380882
R53567 ASIG5V.n4535 ASIG5V.n4318 0.0380882
R53568 ASIG5V.n4531 ASIG5V.n4318 0.0380882
R53569 ASIG5V.n4531 ASIG5V.n4529 0.0380882
R53570 ASIG5V.n4529 ASIG5V.n4527 0.0380882
R53571 ASIG5V.n4527 ASIG5V.n4322 0.0380882
R53572 ASIG5V.n4523 ASIG5V.n4322 0.0380882
R53573 ASIG5V.n4523 ASIG5V.n4521 0.0380882
R53574 ASIG5V.n4521 ASIG5V.n4519 0.0380882
R53575 ASIG5V.n4519 ASIG5V.n4326 0.0380882
R53576 ASIG5V.n4515 ASIG5V.n4326 0.0380882
R53577 ASIG5V.n4515 ASIG5V.n4513 0.0380882
R53578 ASIG5V.n4513 ASIG5V.n4511 0.0380882
R53579 ASIG5V.n4511 ASIG5V.n4330 0.0380882
R53580 ASIG5V.n4507 ASIG5V.n4330 0.0380882
R53581 ASIG5V.n4507 ASIG5V.n4505 0.0380882
R53582 ASIG5V.n4505 ASIG5V.n4503 0.0380882
R53583 ASIG5V.n4503 ASIG5V.n4334 0.0380882
R53584 ASIG5V.n4499 ASIG5V.n4334 0.0380882
R53585 ASIG5V.n4499 ASIG5V.n4497 0.0380882
R53586 ASIG5V.n4497 ASIG5V.n4495 0.0380882
R53587 ASIG5V.n4495 ASIG5V.n4338 0.0380882
R53588 ASIG5V.n4491 ASIG5V.n4338 0.0380882
R53589 ASIG5V.n4491 ASIG5V.n4489 0.0380882
R53590 ASIG5V.n4489 ASIG5V.n4487 0.0380882
R53591 ASIG5V.n4487 ASIG5V.n4342 0.0380882
R53592 ASIG5V.n4483 ASIG5V.n4342 0.0380882
R53593 ASIG5V.n4483 ASIG5V.n4481 0.0380882
R53594 ASIG5V.n4481 ASIG5V.n4479 0.0380882
R53595 ASIG5V.n4479 ASIG5V.n4346 0.0380882
R53596 ASIG5V.n4475 ASIG5V.n4346 0.0380882
R53597 ASIG5V.n4475 ASIG5V.n4473 0.0380882
R53598 ASIG5V.n4473 ASIG5V.n4471 0.0380882
R53599 ASIG5V.n4471 ASIG5V.n4350 0.0380882
R53600 ASIG5V.n4467 ASIG5V.n4350 0.0380882
R53601 ASIG5V.n4467 ASIG5V.n4465 0.0380882
R53602 ASIG5V.n4465 ASIG5V.n4463 0.0380882
R53603 ASIG5V.n4463 ASIG5V.n4354 0.0380882
R53604 ASIG5V.n4459 ASIG5V.n4354 0.0380882
R53605 ASIG5V.n4459 ASIG5V.n4457 0.0380882
R53606 ASIG5V.n4457 ASIG5V.n4455 0.0380882
R53607 ASIG5V.n4455 ASIG5V.n4358 0.0380882
R53608 ASIG5V.n4451 ASIG5V.n4358 0.0380882
R53609 ASIG5V.n4451 ASIG5V.n4449 0.0380882
R53610 ASIG5V.n4449 ASIG5V.n4447 0.0380882
R53611 ASIG5V.n4447 ASIG5V.n4362 0.0380882
R53612 ASIG5V.n4443 ASIG5V.n4362 0.0380882
R53613 ASIG5V.n4443 ASIG5V.n4441 0.0380882
R53614 ASIG5V.n4441 ASIG5V.n4439 0.0380882
R53615 ASIG5V.n4439 ASIG5V.n4366 0.0380882
R53616 ASIG5V.n4435 ASIG5V.n4366 0.0380882
R53617 ASIG5V.n4435 ASIG5V.n4433 0.0380882
R53618 ASIG5V.n4433 ASIG5V.n4431 0.0380882
R53619 ASIG5V.n4431 ASIG5V.n4370 0.0380882
R53620 ASIG5V.n4427 ASIG5V.n4370 0.0380882
R53621 ASIG5V.n4427 ASIG5V.n4425 0.0380882
R53622 ASIG5V.n4425 ASIG5V.n4423 0.0380882
R53623 ASIG5V.n4423 ASIG5V.n4374 0.0380882
R53624 ASIG5V.n4419 ASIG5V.n4374 0.0380882
R53625 ASIG5V.n4419 ASIG5V.n4417 0.0380882
R53626 ASIG5V.n4417 ASIG5V.n4415 0.0380882
R53627 ASIG5V.n4415 ASIG5V.n4378 0.0380882
R53628 ASIG5V.n4411 ASIG5V.n4378 0.0380882
R53629 ASIG5V.n4411 ASIG5V.n4409 0.0380882
R53630 ASIG5V.n4409 ASIG5V.n4407 0.0380882
R53631 ASIG5V.n4407 ASIG5V.n4382 0.0380882
R53632 ASIG5V.n4403 ASIG5V.n4382 0.0380882
R53633 ASIG5V.n4403 ASIG5V.n4401 0.0380882
R53634 ASIG5V.n4401 ASIG5V.n4399 0.0380882
R53635 ASIG5V.n4399 ASIG5V.n4386 0.0380882
R53636 ASIG5V.n4395 ASIG5V.n4386 0.0380882
R53637 ASIG5V.n4395 ASIG5V.n4393 0.0380882
R53638 ASIG5V.n4393 ASIG5V.n4391 0.0380882
R53639 ASIG5V.n4391 ASIG5V.n3834 0.0380882
R53640 ASIG5V.n4566 ASIG5V.n3834 0.0380882
R53641 ASIG5V.n10353 ASIG5V.n10116 0.0380882
R53642 ASIG5V.n10353 ASIG5V.n10118 0.0380882
R53643 ASIG5V.n10349 ASIG5V.n10118 0.0380882
R53644 ASIG5V.n10349 ASIG5V.n10347 0.0380882
R53645 ASIG5V.n10347 ASIG5V.n10345 0.0380882
R53646 ASIG5V.n10345 ASIG5V.n10122 0.0380882
R53647 ASIG5V.n10340 ASIG5V.n10122 0.0380882
R53648 ASIG5V.n10340 ASIG5V.n10338 0.0380882
R53649 ASIG5V.n10338 ASIG5V.n10336 0.0380882
R53650 ASIG5V.n10336 ASIG5V.n10125 0.0380882
R53651 ASIG5V.n10331 ASIG5V.n10125 0.0380882
R53652 ASIG5V.n10331 ASIG5V.n10329 0.0380882
R53653 ASIG5V.n10329 ASIG5V.n10327 0.0380882
R53654 ASIG5V.n10327 ASIG5V.n10128 0.0380882
R53655 ASIG5V.n10322 ASIG5V.n10128 0.0380882
R53656 ASIG5V.n10322 ASIG5V.n10320 0.0380882
R53657 ASIG5V.n10320 ASIG5V.n10318 0.0380882
R53658 ASIG5V.n10318 ASIG5V.n10131 0.0380882
R53659 ASIG5V.n10313 ASIG5V.n10131 0.0380882
R53660 ASIG5V.n10313 ASIG5V.n10311 0.0380882
R53661 ASIG5V.n10311 ASIG5V.n10309 0.0380882
R53662 ASIG5V.n10309 ASIG5V.n10134 0.0380882
R53663 ASIG5V.n10304 ASIG5V.n10134 0.0380882
R53664 ASIG5V.n10304 ASIG5V.n10302 0.0380882
R53665 ASIG5V.n10302 ASIG5V.n10300 0.0380882
R53666 ASIG5V.n10300 ASIG5V.n10137 0.0380882
R53667 ASIG5V.n10295 ASIG5V.n10137 0.0380882
R53668 ASIG5V.n10295 ASIG5V.n10293 0.0380882
R53669 ASIG5V.n10293 ASIG5V.n10291 0.0380882
R53670 ASIG5V.n10291 ASIG5V.n10140 0.0380882
R53671 ASIG5V.n10286 ASIG5V.n10140 0.0380882
R53672 ASIG5V.n10286 ASIG5V.n10284 0.0380882
R53673 ASIG5V.n10284 ASIG5V.n10282 0.0380882
R53674 ASIG5V.n10282 ASIG5V.n10143 0.0380882
R53675 ASIG5V.n10277 ASIG5V.n10143 0.0380882
R53676 ASIG5V.n10277 ASIG5V.n10275 0.0380882
R53677 ASIG5V.n10275 ASIG5V.n10273 0.0380882
R53678 ASIG5V.n10273 ASIG5V.n10146 0.0380882
R53679 ASIG5V.n10268 ASIG5V.n10146 0.0380882
R53680 ASIG5V.n10268 ASIG5V.n10266 0.0380882
R53681 ASIG5V.n10266 ASIG5V.n10264 0.0380882
R53682 ASIG5V.n10264 ASIG5V.n10149 0.0380882
R53683 ASIG5V.n10259 ASIG5V.n10149 0.0380882
R53684 ASIG5V.n10259 ASIG5V.n10257 0.0380882
R53685 ASIG5V.n10257 ASIG5V.n10255 0.0380882
R53686 ASIG5V.n10255 ASIG5V.n10152 0.0380882
R53687 ASIG5V.n10250 ASIG5V.n10152 0.0380882
R53688 ASIG5V.n10250 ASIG5V.n10248 0.0380882
R53689 ASIG5V.n10248 ASIG5V.n10246 0.0380882
R53690 ASIG5V.n10246 ASIG5V.n10155 0.0380882
R53691 ASIG5V.n10241 ASIG5V.n10155 0.0380882
R53692 ASIG5V.n10241 ASIG5V.n10239 0.0380882
R53693 ASIG5V.n10239 ASIG5V.n10237 0.0380882
R53694 ASIG5V.n10237 ASIG5V.n10158 0.0380882
R53695 ASIG5V.n10232 ASIG5V.n10158 0.0380882
R53696 ASIG5V.n10232 ASIG5V.n10230 0.0380882
R53697 ASIG5V.n10230 ASIG5V.n10228 0.0380882
R53698 ASIG5V.n10228 ASIG5V.n10161 0.0380882
R53699 ASIG5V.n10223 ASIG5V.n10161 0.0380882
R53700 ASIG5V.n10223 ASIG5V.n10221 0.0380882
R53701 ASIG5V.n10221 ASIG5V.n10219 0.0380882
R53702 ASIG5V.n10219 ASIG5V.n10164 0.0380882
R53703 ASIG5V.n10214 ASIG5V.n10164 0.0380882
R53704 ASIG5V.n10214 ASIG5V.n10212 0.0380882
R53705 ASIG5V.n10212 ASIG5V.n10210 0.0380882
R53706 ASIG5V.n10210 ASIG5V.n10167 0.0380882
R53707 ASIG5V.n10205 ASIG5V.n10167 0.0380882
R53708 ASIG5V.n10205 ASIG5V.n10203 0.0380882
R53709 ASIG5V.n10203 ASIG5V.n10201 0.0380882
R53710 ASIG5V.n10201 ASIG5V.n10170 0.0380882
R53711 ASIG5V.n10196 ASIG5V.n10170 0.0380882
R53712 ASIG5V.n10196 ASIG5V.n10194 0.0380882
R53713 ASIG5V.n10194 ASIG5V.n10192 0.0380882
R53714 ASIG5V.n10192 ASIG5V.n10173 0.0380882
R53715 ASIG5V.n10187 ASIG5V.n10173 0.0380882
R53716 ASIG5V.n10187 ASIG5V.n10185 0.0380882
R53717 ASIG5V.n10185 ASIG5V.n10183 0.0380882
R53718 ASIG5V.n10183 ASIG5V.n10176 0.0380882
R53719 ASIG5V.n10178 ASIG5V.n10176 0.0380882
R53720 ASIG5V.n10178 ASIG5V.n10074 0.0380882
R53721 ASIG5V.n10359 ASIG5V.n10074 0.0380882
R53722 ASIG5V.n10359 ASIG5V.n10072 0.0380882
R53723 ASIG5V.n11181 ASIG5V.n10072 0.0380882
R53724 ASIG5V.n11160 ASIG5V.n10463 0.0380882
R53725 ASIG5V.n11160 ASIG5V.n10465 0.0380882
R53726 ASIG5V.n11156 ASIG5V.n10465 0.0380882
R53727 ASIG5V.n11156 ASIG5V.n11154 0.0380882
R53728 ASIG5V.n11154 ASIG5V.n11152 0.0380882
R53729 ASIG5V.n11152 ASIG5V.n10929 0.0380882
R53730 ASIG5V.n11148 ASIG5V.n10929 0.0380882
R53731 ASIG5V.n11148 ASIG5V.n11146 0.0380882
R53732 ASIG5V.n11146 ASIG5V.n11144 0.0380882
R53733 ASIG5V.n11144 ASIG5V.n10933 0.0380882
R53734 ASIG5V.n11140 ASIG5V.n10933 0.0380882
R53735 ASIG5V.n11140 ASIG5V.n11138 0.0380882
R53736 ASIG5V.n11138 ASIG5V.n11136 0.0380882
R53737 ASIG5V.n11136 ASIG5V.n10937 0.0380882
R53738 ASIG5V.n11132 ASIG5V.n10937 0.0380882
R53739 ASIG5V.n11132 ASIG5V.n11130 0.0380882
R53740 ASIG5V.n11130 ASIG5V.n11128 0.0380882
R53741 ASIG5V.n11128 ASIG5V.n10941 0.0380882
R53742 ASIG5V.n11124 ASIG5V.n10941 0.0380882
R53743 ASIG5V.n11124 ASIG5V.n11122 0.0380882
R53744 ASIG5V.n11122 ASIG5V.n11120 0.0380882
R53745 ASIG5V.n11120 ASIG5V.n10945 0.0380882
R53746 ASIG5V.n11116 ASIG5V.n10945 0.0380882
R53747 ASIG5V.n11116 ASIG5V.n11114 0.0380882
R53748 ASIG5V.n11114 ASIG5V.n11112 0.0380882
R53749 ASIG5V.n11112 ASIG5V.n10949 0.0380882
R53750 ASIG5V.n11108 ASIG5V.n10949 0.0380882
R53751 ASIG5V.n11108 ASIG5V.n11106 0.0380882
R53752 ASIG5V.n11106 ASIG5V.n11104 0.0380882
R53753 ASIG5V.n11104 ASIG5V.n10953 0.0380882
R53754 ASIG5V.n11100 ASIG5V.n10953 0.0380882
R53755 ASIG5V.n11100 ASIG5V.n11098 0.0380882
R53756 ASIG5V.n11098 ASIG5V.n11096 0.0380882
R53757 ASIG5V.n11096 ASIG5V.n10957 0.0380882
R53758 ASIG5V.n11092 ASIG5V.n10957 0.0380882
R53759 ASIG5V.n11092 ASIG5V.n11090 0.0380882
R53760 ASIG5V.n11090 ASIG5V.n11088 0.0380882
R53761 ASIG5V.n11088 ASIG5V.n10961 0.0380882
R53762 ASIG5V.n11084 ASIG5V.n10961 0.0380882
R53763 ASIG5V.n11084 ASIG5V.n11082 0.0380882
R53764 ASIG5V.n11082 ASIG5V.n11080 0.0380882
R53765 ASIG5V.n11080 ASIG5V.n10965 0.0380882
R53766 ASIG5V.n11076 ASIG5V.n10965 0.0380882
R53767 ASIG5V.n11076 ASIG5V.n11074 0.0380882
R53768 ASIG5V.n11074 ASIG5V.n11072 0.0380882
R53769 ASIG5V.n11072 ASIG5V.n10969 0.0380882
R53770 ASIG5V.n11068 ASIG5V.n10969 0.0380882
R53771 ASIG5V.n11068 ASIG5V.n11066 0.0380882
R53772 ASIG5V.n11066 ASIG5V.n11064 0.0380882
R53773 ASIG5V.n11064 ASIG5V.n10973 0.0380882
R53774 ASIG5V.n11060 ASIG5V.n10973 0.0380882
R53775 ASIG5V.n11060 ASIG5V.n11058 0.0380882
R53776 ASIG5V.n11058 ASIG5V.n11056 0.0380882
R53777 ASIG5V.n11056 ASIG5V.n10977 0.0380882
R53778 ASIG5V.n11052 ASIG5V.n10977 0.0380882
R53779 ASIG5V.n11052 ASIG5V.n11050 0.0380882
R53780 ASIG5V.n11050 ASIG5V.n11048 0.0380882
R53781 ASIG5V.n11048 ASIG5V.n10981 0.0380882
R53782 ASIG5V.n11044 ASIG5V.n10981 0.0380882
R53783 ASIG5V.n11044 ASIG5V.n11042 0.0380882
R53784 ASIG5V.n11042 ASIG5V.n11040 0.0380882
R53785 ASIG5V.n11040 ASIG5V.n10985 0.0380882
R53786 ASIG5V.n11036 ASIG5V.n10985 0.0380882
R53787 ASIG5V.n11036 ASIG5V.n11034 0.0380882
R53788 ASIG5V.n11034 ASIG5V.n11032 0.0380882
R53789 ASIG5V.n11032 ASIG5V.n10989 0.0380882
R53790 ASIG5V.n11028 ASIG5V.n10989 0.0380882
R53791 ASIG5V.n11028 ASIG5V.n11026 0.0380882
R53792 ASIG5V.n11026 ASIG5V.n11024 0.0380882
R53793 ASIG5V.n11024 ASIG5V.n10993 0.0380882
R53794 ASIG5V.n11020 ASIG5V.n10993 0.0380882
R53795 ASIG5V.n11020 ASIG5V.n11018 0.0380882
R53796 ASIG5V.n11018 ASIG5V.n11016 0.0380882
R53797 ASIG5V.n11016 ASIG5V.n10997 0.0380882
R53798 ASIG5V.n11012 ASIG5V.n10997 0.0380882
R53799 ASIG5V.n11012 ASIG5V.n11010 0.0380882
R53800 ASIG5V.n11010 ASIG5V.n11008 0.0380882
R53801 ASIG5V.n11008 ASIG5V.n11001 0.0380882
R53802 ASIG5V.n11004 ASIG5V.n11001 0.0380882
R53803 ASIG5V.n11004 ASIG5V.n10421 0.0380882
R53804 ASIG5V.n11166 ASIG5V.n10421 0.0380882
R53805 ASIG5V.n11166 ASIG5V.n10419 0.0380882
R53806 ASIG5V.n11170 ASIG5V.n10419 0.0380882
R53807 ASIG5V.n11159 ASIG5V.n10926 0.0380882
R53808 ASIG5V.n11159 ASIG5V.n11158 0.0380882
R53809 ASIG5V.n11158 ASIG5V.n11157 0.0380882
R53810 ASIG5V.n11157 ASIG5V.n10927 0.0380882
R53811 ASIG5V.n11151 ASIG5V.n10927 0.0380882
R53812 ASIG5V.n11151 ASIG5V.n11150 0.0380882
R53813 ASIG5V.n11150 ASIG5V.n11149 0.0380882
R53814 ASIG5V.n11149 ASIG5V.n10931 0.0380882
R53815 ASIG5V.n11143 ASIG5V.n10931 0.0380882
R53816 ASIG5V.n11143 ASIG5V.n11142 0.0380882
R53817 ASIG5V.n11142 ASIG5V.n11141 0.0380882
R53818 ASIG5V.n11141 ASIG5V.n10935 0.0380882
R53819 ASIG5V.n11135 ASIG5V.n10935 0.0380882
R53820 ASIG5V.n11135 ASIG5V.n11134 0.0380882
R53821 ASIG5V.n11134 ASIG5V.n11133 0.0380882
R53822 ASIG5V.n11133 ASIG5V.n10939 0.0380882
R53823 ASIG5V.n11127 ASIG5V.n10939 0.0380882
R53824 ASIG5V.n11127 ASIG5V.n11126 0.0380882
R53825 ASIG5V.n11126 ASIG5V.n11125 0.0380882
R53826 ASIG5V.n11125 ASIG5V.n10943 0.0380882
R53827 ASIG5V.n11119 ASIG5V.n10943 0.0380882
R53828 ASIG5V.n11119 ASIG5V.n11118 0.0380882
R53829 ASIG5V.n11118 ASIG5V.n11117 0.0380882
R53830 ASIG5V.n11117 ASIG5V.n10947 0.0380882
R53831 ASIG5V.n11111 ASIG5V.n10947 0.0380882
R53832 ASIG5V.n11111 ASIG5V.n11110 0.0380882
R53833 ASIG5V.n11110 ASIG5V.n11109 0.0380882
R53834 ASIG5V.n11109 ASIG5V.n10951 0.0380882
R53835 ASIG5V.n11103 ASIG5V.n10951 0.0380882
R53836 ASIG5V.n11103 ASIG5V.n11102 0.0380882
R53837 ASIG5V.n11102 ASIG5V.n11101 0.0380882
R53838 ASIG5V.n11101 ASIG5V.n10955 0.0380882
R53839 ASIG5V.n11095 ASIG5V.n10955 0.0380882
R53840 ASIG5V.n11095 ASIG5V.n11094 0.0380882
R53841 ASIG5V.n11094 ASIG5V.n11093 0.0380882
R53842 ASIG5V.n11093 ASIG5V.n10959 0.0380882
R53843 ASIG5V.n11087 ASIG5V.n10959 0.0380882
R53844 ASIG5V.n11087 ASIG5V.n11086 0.0380882
R53845 ASIG5V.n11086 ASIG5V.n11085 0.0380882
R53846 ASIG5V.n11085 ASIG5V.n10963 0.0380882
R53847 ASIG5V.n11079 ASIG5V.n10963 0.0380882
R53848 ASIG5V.n11079 ASIG5V.n11078 0.0380882
R53849 ASIG5V.n11078 ASIG5V.n11077 0.0380882
R53850 ASIG5V.n11077 ASIG5V.n10967 0.0380882
R53851 ASIG5V.n11071 ASIG5V.n10967 0.0380882
R53852 ASIG5V.n11071 ASIG5V.n11070 0.0380882
R53853 ASIG5V.n11070 ASIG5V.n11069 0.0380882
R53854 ASIG5V.n11069 ASIG5V.n10971 0.0380882
R53855 ASIG5V.n11063 ASIG5V.n10971 0.0380882
R53856 ASIG5V.n11063 ASIG5V.n11062 0.0380882
R53857 ASIG5V.n11062 ASIG5V.n11061 0.0380882
R53858 ASIG5V.n11061 ASIG5V.n10975 0.0380882
R53859 ASIG5V.n11055 ASIG5V.n10975 0.0380882
R53860 ASIG5V.n11055 ASIG5V.n11054 0.0380882
R53861 ASIG5V.n11054 ASIG5V.n11053 0.0380882
R53862 ASIG5V.n11053 ASIG5V.n10979 0.0380882
R53863 ASIG5V.n11047 ASIG5V.n10979 0.0380882
R53864 ASIG5V.n11047 ASIG5V.n11046 0.0380882
R53865 ASIG5V.n11046 ASIG5V.n11045 0.0380882
R53866 ASIG5V.n11045 ASIG5V.n10983 0.0380882
R53867 ASIG5V.n11039 ASIG5V.n10983 0.0380882
R53868 ASIG5V.n11039 ASIG5V.n11038 0.0380882
R53869 ASIG5V.n11038 ASIG5V.n11037 0.0380882
R53870 ASIG5V.n11037 ASIG5V.n10987 0.0380882
R53871 ASIG5V.n11031 ASIG5V.n10987 0.0380882
R53872 ASIG5V.n11031 ASIG5V.n11030 0.0380882
R53873 ASIG5V.n11030 ASIG5V.n11029 0.0380882
R53874 ASIG5V.n11029 ASIG5V.n10991 0.0380882
R53875 ASIG5V.n11023 ASIG5V.n10991 0.0380882
R53876 ASIG5V.n11023 ASIG5V.n11022 0.0380882
R53877 ASIG5V.n11022 ASIG5V.n11021 0.0380882
R53878 ASIG5V.n11021 ASIG5V.n10995 0.0380882
R53879 ASIG5V.n11015 ASIG5V.n10995 0.0380882
R53880 ASIG5V.n11015 ASIG5V.n11014 0.0380882
R53881 ASIG5V.n11014 ASIG5V.n11013 0.0380882
R53882 ASIG5V.n11013 ASIG5V.n10999 0.0380882
R53883 ASIG5V.n11007 ASIG5V.n10999 0.0380882
R53884 ASIG5V.n11007 ASIG5V.n11006 0.0380882
R53885 ASIG5V.n11006 ASIG5V.n11005 0.0380882
R53886 ASIG5V.n11005 ASIG5V.n10420 0.0380882
R53887 ASIG5V.n11167 ASIG5V.n10420 0.0380882
R53888 ASIG5V.n11168 ASIG5V.n11167 0.0380882
R53889 ASIG5V.n11169 ASIG5V.n11168 0.0380882
R53890 ASIG5V.n4550 ASIG5V.n3783 0.0380882
R53891 ASIG5V.n4550 ASIG5V.n4549 0.0380882
R53892 ASIG5V.n4549 ASIG5V.n4548 0.0380882
R53893 ASIG5V.n4548 ASIG5V.n4312 0.0380882
R53894 ASIG5V.n4542 ASIG5V.n4312 0.0380882
R53895 ASIG5V.n4542 ASIG5V.n4541 0.0380882
R53896 ASIG5V.n4541 ASIG5V.n4540 0.0380882
R53897 ASIG5V.n4540 ASIG5V.n4316 0.0380882
R53898 ASIG5V.n4534 ASIG5V.n4316 0.0380882
R53899 ASIG5V.n4534 ASIG5V.n4533 0.0380882
R53900 ASIG5V.n4533 ASIG5V.n4532 0.0380882
R53901 ASIG5V.n4532 ASIG5V.n4320 0.0380882
R53902 ASIG5V.n4526 ASIG5V.n4320 0.0380882
R53903 ASIG5V.n4526 ASIG5V.n4525 0.0380882
R53904 ASIG5V.n4525 ASIG5V.n4524 0.0380882
R53905 ASIG5V.n4524 ASIG5V.n4324 0.0380882
R53906 ASIG5V.n4518 ASIG5V.n4324 0.0380882
R53907 ASIG5V.n4518 ASIG5V.n4517 0.0380882
R53908 ASIG5V.n4517 ASIG5V.n4516 0.0380882
R53909 ASIG5V.n4516 ASIG5V.n4328 0.0380882
R53910 ASIG5V.n4510 ASIG5V.n4328 0.0380882
R53911 ASIG5V.n4510 ASIG5V.n4509 0.0380882
R53912 ASIG5V.n4509 ASIG5V.n4508 0.0380882
R53913 ASIG5V.n4508 ASIG5V.n4332 0.0380882
R53914 ASIG5V.n4502 ASIG5V.n4332 0.0380882
R53915 ASIG5V.n4502 ASIG5V.n4501 0.0380882
R53916 ASIG5V.n4501 ASIG5V.n4500 0.0380882
R53917 ASIG5V.n4500 ASIG5V.n4336 0.0380882
R53918 ASIG5V.n4494 ASIG5V.n4336 0.0380882
R53919 ASIG5V.n4494 ASIG5V.n4493 0.0380882
R53920 ASIG5V.n4493 ASIG5V.n4492 0.0380882
R53921 ASIG5V.n4492 ASIG5V.n4340 0.0380882
R53922 ASIG5V.n4486 ASIG5V.n4340 0.0380882
R53923 ASIG5V.n4486 ASIG5V.n4485 0.0380882
R53924 ASIG5V.n4485 ASIG5V.n4484 0.0380882
R53925 ASIG5V.n4484 ASIG5V.n4344 0.0380882
R53926 ASIG5V.n4478 ASIG5V.n4344 0.0380882
R53927 ASIG5V.n4478 ASIG5V.n4477 0.0380882
R53928 ASIG5V.n4477 ASIG5V.n4476 0.0380882
R53929 ASIG5V.n4476 ASIG5V.n4348 0.0380882
R53930 ASIG5V.n4470 ASIG5V.n4348 0.0380882
R53931 ASIG5V.n4470 ASIG5V.n4469 0.0380882
R53932 ASIG5V.n4469 ASIG5V.n4468 0.0380882
R53933 ASIG5V.n4468 ASIG5V.n4352 0.0380882
R53934 ASIG5V.n4462 ASIG5V.n4352 0.0380882
R53935 ASIG5V.n4462 ASIG5V.n4461 0.0380882
R53936 ASIG5V.n4461 ASIG5V.n4460 0.0380882
R53937 ASIG5V.n4460 ASIG5V.n4356 0.0380882
R53938 ASIG5V.n4454 ASIG5V.n4356 0.0380882
R53939 ASIG5V.n4454 ASIG5V.n4453 0.0380882
R53940 ASIG5V.n4453 ASIG5V.n4452 0.0380882
R53941 ASIG5V.n4452 ASIG5V.n4360 0.0380882
R53942 ASIG5V.n4446 ASIG5V.n4360 0.0380882
R53943 ASIG5V.n4446 ASIG5V.n4445 0.0380882
R53944 ASIG5V.n4445 ASIG5V.n4444 0.0380882
R53945 ASIG5V.n4444 ASIG5V.n4364 0.0380882
R53946 ASIG5V.n4438 ASIG5V.n4364 0.0380882
R53947 ASIG5V.n4438 ASIG5V.n4437 0.0380882
R53948 ASIG5V.n4437 ASIG5V.n4436 0.0380882
R53949 ASIG5V.n4436 ASIG5V.n4368 0.0380882
R53950 ASIG5V.n4430 ASIG5V.n4368 0.0380882
R53951 ASIG5V.n4430 ASIG5V.n4429 0.0380882
R53952 ASIG5V.n4429 ASIG5V.n4428 0.0380882
R53953 ASIG5V.n4428 ASIG5V.n4372 0.0380882
R53954 ASIG5V.n4422 ASIG5V.n4372 0.0380882
R53955 ASIG5V.n4422 ASIG5V.n4421 0.0380882
R53956 ASIG5V.n4421 ASIG5V.n4420 0.0380882
R53957 ASIG5V.n4420 ASIG5V.n4376 0.0380882
R53958 ASIG5V.n4414 ASIG5V.n4376 0.0380882
R53959 ASIG5V.n4414 ASIG5V.n4413 0.0380882
R53960 ASIG5V.n4413 ASIG5V.n4412 0.0380882
R53961 ASIG5V.n4412 ASIG5V.n4380 0.0380882
R53962 ASIG5V.n4406 ASIG5V.n4380 0.0380882
R53963 ASIG5V.n4406 ASIG5V.n4405 0.0380882
R53964 ASIG5V.n4405 ASIG5V.n4404 0.0380882
R53965 ASIG5V.n4404 ASIG5V.n4384 0.0380882
R53966 ASIG5V.n4398 ASIG5V.n4384 0.0380882
R53967 ASIG5V.n4398 ASIG5V.n4397 0.0380882
R53968 ASIG5V.n4397 ASIG5V.n4396 0.0380882
R53969 ASIG5V.n4396 ASIG5V.n4388 0.0380882
R53970 ASIG5V.n4390 ASIG5V.n4388 0.0380882
R53971 ASIG5V.n4390 ASIG5V.n3836 0.0380882
R53972 ASIG5V.n4565 ASIG5V.n3836 0.0380882
R53973 ASIG5V.n4249 ASIG5V.n3837 0.03245
R53974 ASIG5V.n4560 ASIG5V.n3837 0.03245
R53975 ASIG5V.n4563 ASIG5V.n3624 0.03245
R53976 ASIG5V.n4780 ASIG5V.n3624 0.03245
R53977 ASIG5V.n4783 ASIG5V.n4782 0.03245
R53978 ASIG5V.n4803 ASIG5V.n4802 0.03245
R53979 ASIG5V.n4804 ASIG5V.n4803 0.03245
R53980 ASIG5V.n5069 ASIG5V.n5068 0.03245
R53981 ASIG5V.n9740 ASIG5V.n5069 0.03245
R53982 ASIG5V.n9738 ASIG5V.n5071 0.03245
R53983 ASIG5V.n5457 ASIG5V.n5071 0.03245
R53984 ASIG5V.n9424 ASIG5V.n5458 0.03245
R53985 ASIG5V.n5561 ASIG5V.n5458 0.03245
R53986 ASIG5V.n9411 ASIG5V.n9410 0.03245
R53987 ASIG5V.n9410 ASIG5V.n9409 0.03245
R53988 ASIG5V.n6257 ASIG5V.n6256 0.03245
R53989 ASIG5V.n9388 ASIG5V.n9387 0.03245
R53990 ASIG5V.n9387 ASIG5V.n9386 0.03245
R53991 ASIG5V.n6440 ASIG5V.n6439 0.03245
R53992 ASIG5V.n9182 ASIG5V.n6440 0.03245
R53993 ASIG5V.n9180 ASIG5V.n6442 0.03245
R53994 ASIG5V.n6885 ASIG5V.n6442 0.03245
R53995 ASIG5V.n8911 ASIG5V.n8910 0.03245
R53996 ASIG5V.n8910 ASIG5V.n8909 0.03245
R53997 ASIG5V.n8273 ASIG5V.n8272 0.03245
R53998 ASIG5V.n8887 ASIG5V.n8886 0.03245
R53999 ASIG5V.n8886 ASIG5V.n8885 0.03245
R54000 ASIG5V.n12534 ASIG5V.n12533 0.03245
R54001 ASIG5V.n12533 ASIG5V.n12532 0.03245
R54002 ASIG5V.n510 ASIG5V.n509 0.03245
R54003 ASIG5V.n509 ASIG5V.n505 0.03245
R54004 ASIG5V.n12315 ASIG5V.n506 0.03245
R54005 ASIG5V.n859 ASIG5V.n506 0.03245
R54006 ASIG5V.n12293 ASIG5V.n860 0.03245
R54007 ASIG5V.n1218 ASIG5V.n860 0.03245
R54008 ASIG5V.n12275 ASIG5V.n12274 0.03245
R54009 ASIG5V.n12272 ASIG5V.n1221 0.03245
R54010 ASIG5V.n1668 ASIG5V.n1221 0.03245
R54011 ASIG5V.n12003 ASIG5V.n12002 0.03245
R54012 ASIG5V.n12002 ASIG5V.n12001 0.03245
R54013 ASIG5V.n1858 ASIG5V.n1855 0.03245
R54014 ASIG5V.n2203 ASIG5V.n1855 0.03245
R54015 ASIG5V.n11788 ASIG5V.n2205 0.03245
R54016 ASIG5V.n11788 ASIG5V.n11787 0.03245
R54017 ASIG5V.n11785 ASIG5V.n2207 0.03245
R54018 ASIG5V.n11763 ASIG5V.n2902 0.03245
R54019 ASIG5V.n11757 ASIG5V.n2902 0.03245
R54020 ASIG5V.n11755 ASIG5V.n2910 0.03245
R54021 ASIG5V.n11491 ASIG5V.n2910 0.03245
R54022 ASIG5V.n11489 ASIG5V.n9970 0.03245
R54023 ASIG5V.n10367 ASIG5V.n9970 0.03245
R54024 ASIG5V.n11178 ASIG5V.n11177 0.03245
R54025 ASIG5V.n11177 ASIG5V.n11176 0.03245
R54026 ASIG5V.n10916 ASIG5V.n10488 0.03245
R54027 ASIG5V.n10916 ASIG5V.n10915 0.03245
R54028 ASIG5V.n4783 ASIG5V.n3273 0.031775
R54029 ASIG5V.n10119 ASIG5V.n10022 0.0317353
R54030 ASIG5V.n4792 ASIG5V.n3616 0.0317353
R54031 ASIG5V.n4816 ASIG5V.n3267 0.0317353
R54032 ASIG5V.n9487 ASIG5V.n3164 0.0317353
R54033 ASIG5V.n5215 ASIG5V.n5120 0.0317353
R54034 ASIG5V.n7971 ASIG5V.n7960 0.0317353
R54035 ASIG5V.n5908 ASIG5V.n5907 0.0317353
R54036 ASIG5V.n6063 ASIG5V.n5909 0.0317353
R54037 ASIG5V.n9192 ASIG5V.n9191 0.0317353
R54038 ASIG5V.n8929 ASIG5V.n6533 0.0317353
R54039 ASIG5V.n6696 ASIG5V.n6540 0.0317353
R54040 ASIG5V.n7244 ASIG5V.n7231 0.0317353
R54041 ASIG5V.n8569 ASIG5V.n8568 0.0317353
R54042 ASIG5V.n8588 ASIG5V.n8587 0.0317353
R54043 ASIG5V.n12338 ASIG5V.n12337 0.0317353
R54044 ASIG5V.n12329 ASIG5V.n168 0.0317353
R54045 ASIG5V.n12306 ASIG5V.n524 0.0317353
R54046 ASIG5V.n12283 ASIG5V.n869 0.0317353
R54047 ASIG5V.n12021 ASIG5V.n1316 0.0317353
R54048 ASIG5V.n1479 ASIG5V.n1322 0.0317353
R54049 ASIG5V.n11807 ASIG5V.n11806 0.0317353
R54050 ASIG5V.n11796 ASIG5V.n1842 0.0317353
R54051 ASIG5V.n2561 ASIG5V.n2218 0.0317353
R54052 ASIG5V.n11776 ASIG5V.n2563 0.0317353
R54053 ASIG5V.n11504 ASIG5V.n3002 0.0317353
R54054 ASIG5V.n11238 ASIG5V.n9961 0.0317353
R54055 ASIG5V.n4585 ASIG5V.n4584 0.0317353
R54056 ASIG5V.n10926 ASIG5V.n10925 0.0317353
R54057 ASIG5V.n4573 ASIG5V.n3783 0.0317353
R54058 ASIG5V.n8274 ASIG5V.n8273 0.031325
R54059 ASIG5V.n12275 ASIG5V.n1219 0.030875
R54060 ASIG5V.n11764 ASIG5V.n2207 0.030875
R54061 ASIG5V.n6256 ASIG5V.n5563 0.030425
R54062 ASIG5V.n6258 ASIG5V.n6257 0.028625
R54063 ASIG5V.n4557 ASIG5V.n3839 0.0284039
R54064 ASIG5V.n4558 ASIG5V.n4557 0.0284039
R54065 ASIG5V.n4561 ASIG5V.n3627 0.0284039
R54066 ASIG5V.n4778 ASIG5V.n3627 0.0284039
R54067 ASIG5V.n4785 ASIG5V.n3621 0.0284039
R54068 ASIG5V.n4800 ASIG5V.n3271 0.0284039
R54069 ASIG5V.n4806 ASIG5V.n3271 0.0284039
R54070 ASIG5V.n5066 ASIG5V.n3171 0.0284039
R54071 ASIG5V.n9742 ASIG5V.n3171 0.0284039
R54072 ASIG5V.n9736 ASIG5V.n5073 0.0284039
R54073 ASIG5V.n5459 ASIG5V.n5073 0.0284039
R54074 ASIG5V.n9422 ASIG5V.n9421 0.0284039
R54075 ASIG5V.n9421 ASIG5V.n5463 0.0284039
R54076 ASIG5V.n5565 ASIG5V.n5560 0.0284039
R54077 ASIG5V.n9407 ASIG5V.n5565 0.0284039
R54078 ASIG5V.n6254 ASIG5V.n6251 0.0284039
R54079 ASIG5V.n6261 ASIG5V.n6250 0.0284039
R54080 ASIG5V.n9384 ASIG5V.n6261 0.0284039
R54081 ASIG5V.n6437 ASIG5V.n6433 0.0284039
R54082 ASIG5V.n9184 ASIG5V.n6433 0.0284039
R54083 ASIG5V.n9178 ASIG5V.n6444 0.0284039
R54084 ASIG5V.n6881 ASIG5V.n6444 0.0284039
R54085 ASIG5V.n6889 ASIG5V.n6884 0.0284039
R54086 ASIG5V.n8907 ASIG5V.n6889 0.0284039
R54087 ASIG5V.n8270 ASIG5V.n8267 0.0284039
R54088 ASIG5V.n8275 ASIG5V.n8266 0.0284039
R54089 ASIG5V.n8883 ASIG5V.n8275 0.0284039
R54090 ASIG5V.n12536 ASIG5V.n3 0.0284039
R54091 ASIG5V.n12530 ASIG5V.n3 0.0284039
R54092 ASIG5V.n514 ASIG5V.n512 0.0284039
R54093 ASIG5V.n515 ASIG5V.n514 0.0284039
R54094 ASIG5V.n12313 ASIG5V.n12312 0.0284039
R54095 ASIG5V.n12312 ASIG5V.n519 0.0284039
R54096 ASIG5V.n12291 ASIG5V.n12290 0.0284039
R54097 ASIG5V.n12290 ASIG5V.n864 0.0284039
R54098 ASIG5V.n12277 ASIG5V.n880 0.0284039
R54099 ASIG5V.n12270 ASIG5V.n1225 0.0284039
R54100 ASIG5V.n1664 ASIG5V.n1225 0.0284039
R54101 ASIG5V.n1672 ASIG5V.n1667 0.0284039
R54102 ASIG5V.n11999 ASIG5V.n1672 0.0284039
R54103 ASIG5V.n1862 ASIG5V.n1860 0.0284039
R54104 ASIG5V.n2201 ASIG5V.n1862 0.0284039
R54105 ASIG5V.n11790 ASIG5V.n1850 0.0284039
R54106 ASIG5V.n11790 ASIG5V.n1851 0.0284039
R54107 ASIG5V.n11783 ASIG5V.n2211 0.0284039
R54108 ASIG5V.n11761 ASIG5V.n11760 0.0284039
R54109 ASIG5V.n11760 ASIG5V.n11759 0.0284039
R54110 ASIG5V.n11753 ASIG5V.n2912 0.0284039
R54111 ASIG5V.n11493 ASIG5V.n2912 0.0284039
R54112 ASIG5V.n11487 ASIG5V.n9972 0.0284039
R54113 ASIG5V.n10363 ASIG5V.n9972 0.0284039
R54114 ASIG5V.n10371 ASIG5V.n10366 0.0284039
R54115 ASIG5V.n11174 ASIG5V.n10371 0.0284039
R54116 ASIG5V.n10918 ASIG5V.n10484 0.0284039
R54117 ASIG5V.n10918 ASIG5V.n10485 0.0284039
R54118 ASIG5V.n4250 ASIG5V.n3838 0.0284039
R54119 ASIG5V.n4559 ASIG5V.n3838 0.0284039
R54120 ASIG5V.n4562 ASIG5V.n3625 0.0284039
R54121 ASIG5V.n4779 ASIG5V.n3625 0.0284039
R54122 ASIG5V.n4784 ASIG5V.n3622 0.0284039
R54123 ASIG5V.n4801 ASIG5V.n3272 0.0284039
R54124 ASIG5V.n4805 ASIG5V.n3272 0.0284039
R54125 ASIG5V.n5067 ASIG5V.n3173 0.0284039
R54126 ASIG5V.n9741 ASIG5V.n3173 0.0284039
R54127 ASIG5V.n9737 ASIG5V.n5072 0.0284039
R54128 ASIG5V.n5460 ASIG5V.n5072 0.0284039
R54129 ASIG5V.n9423 ASIG5V.n5462 0.0284039
R54130 ASIG5V.n5558 ASIG5V.n5462 0.0284039
R54131 ASIG5V.n9412 ASIG5V.n5559 0.0284039
R54132 ASIG5V.n9408 ASIG5V.n5559 0.0284039
R54133 ASIG5V.n6255 ASIG5V.n6248 0.0284039
R54134 ASIG5V.n9389 ASIG5V.n6249 0.0284039
R54135 ASIG5V.n9385 ASIG5V.n6249 0.0284039
R54136 ASIG5V.n6438 ASIG5V.n6435 0.0284039
R54137 ASIG5V.n9183 ASIG5V.n6435 0.0284039
R54138 ASIG5V.n9179 ASIG5V.n6443 0.0284039
R54139 ASIG5V.n6882 ASIG5V.n6443 0.0284039
R54140 ASIG5V.n8912 ASIG5V.n6883 0.0284039
R54141 ASIG5V.n8908 ASIG5V.n6883 0.0284039
R54142 ASIG5V.n8271 ASIG5V.n8264 0.0284039
R54143 ASIG5V.n8888 ASIG5V.n8265 0.0284039
R54144 ASIG5V.n8884 ASIG5V.n8265 0.0284039
R54145 ASIG5V.n12535 ASIG5V.n5 0.0284039
R54146 ASIG5V.n12531 ASIG5V.n5 0.0284039
R54147 ASIG5V.n511 ASIG5V.n507 0.0284039
R54148 ASIG5V.n516 ASIG5V.n507 0.0284039
R54149 ASIG5V.n12314 ASIG5V.n518 0.0284039
R54150 ASIG5V.n861 ASIG5V.n518 0.0284039
R54151 ASIG5V.n12292 ASIG5V.n863 0.0284039
R54152 ASIG5V.n1217 ASIG5V.n863 0.0284039
R54153 ASIG5V.n12276 ASIG5V.n882 0.0284039
R54154 ASIG5V.n12271 ASIG5V.n1223 0.0284039
R54155 ASIG5V.n1665 ASIG5V.n1223 0.0284039
R54156 ASIG5V.n12004 ASIG5V.n1666 0.0284039
R54157 ASIG5V.n12000 ASIG5V.n1666 0.0284039
R54158 ASIG5V.n1859 ASIG5V.n1856 0.0284039
R54159 ASIG5V.n2202 ASIG5V.n1856 0.0284039
R54160 ASIG5V.n11789 ASIG5V.n1852 0.0284039
R54161 ASIG5V.n11789 ASIG5V.n1853 0.0284039
R54162 ASIG5V.n11784 ASIG5V.n2209 0.0284039
R54163 ASIG5V.n11762 ASIG5V.n2904 0.0284039
R54164 ASIG5V.n11758 ASIG5V.n2904 0.0284039
R54165 ASIG5V.n11754 ASIG5V.n2911 0.0284039
R54166 ASIG5V.n11492 ASIG5V.n2911 0.0284039
R54167 ASIG5V.n11488 ASIG5V.n9971 0.0284039
R54168 ASIG5V.n10364 ASIG5V.n9971 0.0284039
R54169 ASIG5V.n11179 ASIG5V.n10365 0.0284039
R54170 ASIG5V.n11175 ASIG5V.n10365 0.0284039
R54171 ASIG5V.n10917 ASIG5V.n10486 0.0284039
R54172 ASIG5V.n10917 ASIG5V.n10487 0.0284039
R54173 ASIG5V.n12274 ASIG5V.n12273 0.028175
R54174 ASIG5V.n11786 ASIG5V.n11785 0.028175
R54175 ASIG5V.n4785 ASIG5V.n3275 0.0278144
R54176 ASIG5V.n4784 ASIG5V.n3274 0.0278144
R54177 ASIG5V.n8272 ASIG5V.n6887 0.027725
R54178 ASIG5V.n8267 ASIG5V.n8260 0.0274214
R54179 ASIG5V.n8889 ASIG5V.n8264 0.0274214
R54180 ASIG5V.n4782 ASIG5V.n4781 0.027275
R54181 ASIG5V.n12277 ASIG5V.n879 0.0270284
R54182 ASIG5V.n2613 ASIG5V.n2211 0.0270284
R54183 ASIG5V.n12276 ASIG5V.n881 0.0270284
R54184 ASIG5V.n2903 ASIG5V.n2209 0.0270284
R54185 ASIG5V.n6254 ASIG5V.n5566 0.0266354
R54186 ASIG5V.n6255 ASIG5V.n5564 0.0266354
R54187 ASIG5V.n4804 ASIG5V.n3175 0.025925
R54188 ASIG5V.n10368 ASIG5V.n10362 0.0259118
R54189 ASIG5V.n3407 ASIG5V.n3273 0.0259118
R54190 ASIG5V.n5058 ASIG5V.n3175 0.0259118
R54191 ASIG5V.n9739 ASIG5V.n5070 0.0259118
R54192 ASIG5V.n9426 ASIG5V.n9425 0.0259118
R54193 ASIG5V.n5562 ASIG5V.n5557 0.0259118
R54194 ASIG5V.n5698 ASIG5V.n5563 0.0259118
R54195 ASIG5V.n6258 ASIG5V.n6247 0.0259118
R54196 ASIG5V.n9376 ASIG5V.n6259 0.0259118
R54197 ASIG5V.n9181 ASIG5V.n6441 0.0259118
R54198 ASIG5V.n6886 ASIG5V.n6880 0.0259118
R54199 ASIG5V.n7022 ASIG5V.n6887 0.0259118
R54200 ASIG5V.n8274 ASIG5V.n8263 0.0259118
R54201 ASIG5V.n8634 ASIG5V.n6 0.0259118
R54202 ASIG5V.n12522 ASIG5V.n7 0.0259118
R54203 ASIG5V.n12317 ASIG5V.n12316 0.0259118
R54204 ASIG5V.n12295 ASIG5V.n12294 0.0259118
R54205 ASIG5V.n1219 ASIG5V.n1216 0.0259118
R54206 ASIG5V.n12273 ASIG5V.n1220 0.0259118
R54207 ASIG5V.n1669 ASIG5V.n1663 0.0259118
R54208 ASIG5V.n11991 ASIG5V.n1670 0.0259118
R54209 ASIG5V.n2204 ASIG5V.n1854 0.0259118
R54210 ASIG5V.n11786 ASIG5V.n2206 0.0259118
R54211 ASIG5V.n11765 ASIG5V.n11764 0.0259118
R54212 ASIG5V.n11756 ASIG5V.n2909 0.0259118
R54213 ASIG5V.n11490 ASIG5V.n9969 0.0259118
R54214 ASIG5V.n4781 ASIG5V.n3623 0.0259118
R54215 ASIG5V.n11169 ASIG5V.n10369 0.0259118
R54216 ASIG5V.n4565 ASIG5V.n4564 0.0259118
R54217 ASIG5V.n8885 ASIG5V.n6 0.025475
R54218 ASIG5V.n10488 ASIG5V.n10369 0.025475
R54219 ASIG5V.n10716 ASIG5V.n10715 0.0251375
R54220 ASIG5V.n10714 ASIG5V.n10692 0.0251375
R54221 ASIG5V.n10713 ASIG5V.n10497 0.0251375
R54222 ASIG5V.n4101 ASIG5V.n3844 0.0251375
R54223 ASIG5V.n3856 ASIG5V.n3845 0.0251375
R54224 ASIG5V.n4257 ASIG5V.n4256 0.0251375
R54225 ASIG5V.n6251 ASIG5V.n6000 0.0250633
R54226 ASIG5V.n9390 ASIG5V.n6248 0.0250633
R54227 ASIG5V.n12294 ASIG5V.n12293 0.025025
R54228 ASIG5V.n11757 ASIG5V.n11756 0.025025
R54229 ASIG5V.n1224 ASIG5V.n880 0.0246703
R54230 ASIG5V.n11783 ASIG5V.n2210 0.0246703
R54231 ASIG5V.n1222 ASIG5V.n882 0.0246703
R54232 ASIG5V.n11784 ASIG5V.n2208 0.0246703
R54233 ASIG5V.n9411 ASIG5V.n5562 0.024575
R54234 ASIG5V.n8270 ASIG5V.n6890 0.0242773
R54235 ASIG5V.n8271 ASIG5V.n6888 0.0242773
R54236 ASIG5V.n3628 ASIG5V.n3621 0.0238843
R54237 ASIG5V.n3626 ASIG5V.n3622 0.0238843
R54238 ASIG5V.n9386 ASIG5V.n6259 0.022775
R54239 ASIG5V.n4806 ASIG5V.n3177 0.0227052
R54240 ASIG5V.n4805 ASIG5V.n3176 0.0227052
R54241 ASIG5V.n1669 ASIG5V.n1668 0.022325
R54242 ASIG5V.n2205 ASIG5V.n2204 0.022325
R54243 ASIG5V.n8883 ASIG5V.n2 0.0223122
R54244 ASIG5V.n10484 ASIG5V.n10372 0.0223122
R54245 ASIG5V.n8884 ASIG5V.n4 0.0223122
R54246 ASIG5V.n10486 ASIG5V.n10370 0.0223122
R54247 ASIG5V.n12291 ASIG5V.n572 0.0219192
R54248 ASIG5V.n11759 ASIG5V.n2905 0.0219192
R54249 ASIG5V.n12292 ASIG5V.n862 0.0219192
R54250 ASIG5V.n11758 ASIG5V.n2908 0.0219192
R54251 ASIG5V.n8911 ASIG5V.n6886 0.021875
R54252 ASIG5V.n5560 ASIG5V.n5554 0.0215262
R54253 ASIG5V.n9413 ASIG5V.n9412 0.0215262
R54254 ASIG5V.n4564 ASIG5V.n4563 0.021425
R54255 ASIG5V.n9740 ASIG5V.n9739 0.020075
R54256 ASIG5V.n9384 ASIG5V.n6262 0.0199541
R54257 ASIG5V.n9385 ASIG5V.n6260 0.0199541
R54258 ASIG5V.n3613 ASIG5V.n3612 0.019716
R54259 ASIG5V.n3611 ASIG5V.n3610 0.019716
R54260 ASIG5V.n3610 ASIG5V.n3284 0.019716
R54261 ASIG5V.n3604 ASIG5V.n3289 0.019716
R54262 ASIG5V.n3604 ASIG5V.n3603 0.019716
R54263 ASIG5V.n3601 ASIG5V.n3600 0.019716
R54264 ASIG5V.n3600 ASIG5V.n3290 0.019716
R54265 ASIG5V.n3594 ASIG5V.n3295 0.019716
R54266 ASIG5V.n3594 ASIG5V.n3593 0.019716
R54267 ASIG5V.n3591 ASIG5V.n3590 0.019716
R54268 ASIG5V.n3590 ASIG5V.n3296 0.019716
R54269 ASIG5V.n3584 ASIG5V.n3301 0.019716
R54270 ASIG5V.n3584 ASIG5V.n3583 0.019716
R54271 ASIG5V.n3581 ASIG5V.n3580 0.019716
R54272 ASIG5V.n3580 ASIG5V.n3302 0.019716
R54273 ASIG5V.n3574 ASIG5V.n3307 0.019716
R54274 ASIG5V.n3574 ASIG5V.n3573 0.019716
R54275 ASIG5V.n3571 ASIG5V.n3570 0.019716
R54276 ASIG5V.n3570 ASIG5V.n3308 0.019716
R54277 ASIG5V.n3564 ASIG5V.n3313 0.019716
R54278 ASIG5V.n3564 ASIG5V.n3563 0.019716
R54279 ASIG5V.n3561 ASIG5V.n3560 0.019716
R54280 ASIG5V.n3560 ASIG5V.n3314 0.019716
R54281 ASIG5V.n3554 ASIG5V.n3319 0.019716
R54282 ASIG5V.n3554 ASIG5V.n3553 0.019716
R54283 ASIG5V.n3551 ASIG5V.n3550 0.019716
R54284 ASIG5V.n3550 ASIG5V.n3320 0.019716
R54285 ASIG5V.n3544 ASIG5V.n3325 0.019716
R54286 ASIG5V.n3544 ASIG5V.n3543 0.019716
R54287 ASIG5V.n3541 ASIG5V.n3540 0.019716
R54288 ASIG5V.n3540 ASIG5V.n3326 0.019716
R54289 ASIG5V.n3534 ASIG5V.n3331 0.019716
R54290 ASIG5V.n3534 ASIG5V.n3533 0.019716
R54291 ASIG5V.n3531 ASIG5V.n3530 0.019716
R54292 ASIG5V.n3530 ASIG5V.n3332 0.019716
R54293 ASIG5V.n3524 ASIG5V.n3337 0.019716
R54294 ASIG5V.n3524 ASIG5V.n3523 0.019716
R54295 ASIG5V.n3521 ASIG5V.n3520 0.019716
R54296 ASIG5V.n3520 ASIG5V.n3338 0.019716
R54297 ASIG5V.n3514 ASIG5V.n3343 0.019716
R54298 ASIG5V.n3514 ASIG5V.n3513 0.019716
R54299 ASIG5V.n3511 ASIG5V.n3510 0.019716
R54300 ASIG5V.n3510 ASIG5V.n3344 0.019716
R54301 ASIG5V.n3504 ASIG5V.n3349 0.019716
R54302 ASIG5V.n3504 ASIG5V.n3503 0.019716
R54303 ASIG5V.n3501 ASIG5V.n3500 0.019716
R54304 ASIG5V.n3500 ASIG5V.n3350 0.019716
R54305 ASIG5V.n3494 ASIG5V.n3355 0.019716
R54306 ASIG5V.n3494 ASIG5V.n3493 0.019716
R54307 ASIG5V.n3491 ASIG5V.n3490 0.019716
R54308 ASIG5V.n3490 ASIG5V.n3356 0.019716
R54309 ASIG5V.n3484 ASIG5V.n3361 0.019716
R54310 ASIG5V.n3484 ASIG5V.n3483 0.019716
R54311 ASIG5V.n3481 ASIG5V.n3480 0.019716
R54312 ASIG5V.n3480 ASIG5V.n3362 0.019716
R54313 ASIG5V.n3474 ASIG5V.n3367 0.019716
R54314 ASIG5V.n3474 ASIG5V.n3473 0.019716
R54315 ASIG5V.n3471 ASIG5V.n3470 0.019716
R54316 ASIG5V.n3470 ASIG5V.n3368 0.019716
R54317 ASIG5V.n3464 ASIG5V.n3373 0.019716
R54318 ASIG5V.n3464 ASIG5V.n3463 0.019716
R54319 ASIG5V.n3461 ASIG5V.n3460 0.019716
R54320 ASIG5V.n3460 ASIG5V.n3374 0.019716
R54321 ASIG5V.n3454 ASIG5V.n3379 0.019716
R54322 ASIG5V.n3454 ASIG5V.n3453 0.019716
R54323 ASIG5V.n3451 ASIG5V.n3450 0.019716
R54324 ASIG5V.n3450 ASIG5V.n3380 0.019716
R54325 ASIG5V.n3444 ASIG5V.n3385 0.019716
R54326 ASIG5V.n3444 ASIG5V.n3443 0.019716
R54327 ASIG5V.n3441 ASIG5V.n3440 0.019716
R54328 ASIG5V.n3440 ASIG5V.n3386 0.019716
R54329 ASIG5V.n3434 ASIG5V.n3391 0.019716
R54330 ASIG5V.n3434 ASIG5V.n3433 0.019716
R54331 ASIG5V.n3431 ASIG5V.n3430 0.019716
R54332 ASIG5V.n3430 ASIG5V.n3392 0.019716
R54333 ASIG5V.n3424 ASIG5V.n3397 0.019716
R54334 ASIG5V.n3424 ASIG5V.n3423 0.019716
R54335 ASIG5V.n3421 ASIG5V.n3420 0.019716
R54336 ASIG5V.n3420 ASIG5V.n3398 0.019716
R54337 ASIG5V.n3414 ASIG5V.n3403 0.019716
R54338 ASIG5V.n3414 ASIG5V.n3413 0.019716
R54339 ASIG5V.n3411 ASIG5V.n3410 0.019716
R54340 ASIG5V.n3410 ASIG5V.n3404 0.019716
R54341 ASIG5V.n3265 ASIG5V.n3264 0.019716
R54342 ASIG5V.n4820 ASIG5V.n3219 0.019716
R54343 ASIG5V.n4821 ASIG5V.n4820 0.019716
R54344 ASIG5V.n4826 ASIG5V.n3218 0.019716
R54345 ASIG5V.n4826 ASIG5V.n4825 0.019716
R54346 ASIG5V.n4832 ASIG5V.n3217 0.019716
R54347 ASIG5V.n4833 ASIG5V.n4832 0.019716
R54348 ASIG5V.n4838 ASIG5V.n3216 0.019716
R54349 ASIG5V.n4838 ASIG5V.n4837 0.019716
R54350 ASIG5V.n4844 ASIG5V.n3215 0.019716
R54351 ASIG5V.n4845 ASIG5V.n4844 0.019716
R54352 ASIG5V.n4850 ASIG5V.n3214 0.019716
R54353 ASIG5V.n4850 ASIG5V.n4849 0.019716
R54354 ASIG5V.n4856 ASIG5V.n3213 0.019716
R54355 ASIG5V.n4857 ASIG5V.n4856 0.019716
R54356 ASIG5V.n4862 ASIG5V.n3212 0.019716
R54357 ASIG5V.n4862 ASIG5V.n4861 0.019716
R54358 ASIG5V.n4868 ASIG5V.n3211 0.019716
R54359 ASIG5V.n4869 ASIG5V.n4868 0.019716
R54360 ASIG5V.n4874 ASIG5V.n3210 0.019716
R54361 ASIG5V.n4874 ASIG5V.n4873 0.019716
R54362 ASIG5V.n4880 ASIG5V.n3209 0.019716
R54363 ASIG5V.n4881 ASIG5V.n4880 0.019716
R54364 ASIG5V.n4886 ASIG5V.n3208 0.019716
R54365 ASIG5V.n4886 ASIG5V.n4885 0.019716
R54366 ASIG5V.n4892 ASIG5V.n3207 0.019716
R54367 ASIG5V.n4893 ASIG5V.n4892 0.019716
R54368 ASIG5V.n4898 ASIG5V.n3206 0.019716
R54369 ASIG5V.n4898 ASIG5V.n4897 0.019716
R54370 ASIG5V.n4904 ASIG5V.n3205 0.019716
R54371 ASIG5V.n4905 ASIG5V.n4904 0.019716
R54372 ASIG5V.n4910 ASIG5V.n3204 0.019716
R54373 ASIG5V.n4910 ASIG5V.n4909 0.019716
R54374 ASIG5V.n4916 ASIG5V.n3203 0.019716
R54375 ASIG5V.n4917 ASIG5V.n4916 0.019716
R54376 ASIG5V.n4922 ASIG5V.n3202 0.019716
R54377 ASIG5V.n4922 ASIG5V.n4921 0.019716
R54378 ASIG5V.n4928 ASIG5V.n3201 0.019716
R54379 ASIG5V.n4929 ASIG5V.n4928 0.019716
R54380 ASIG5V.n4934 ASIG5V.n3200 0.019716
R54381 ASIG5V.n4934 ASIG5V.n4933 0.019716
R54382 ASIG5V.n4940 ASIG5V.n3199 0.019716
R54383 ASIG5V.n4941 ASIG5V.n4940 0.019716
R54384 ASIG5V.n4946 ASIG5V.n3198 0.019716
R54385 ASIG5V.n4946 ASIG5V.n4945 0.019716
R54386 ASIG5V.n4952 ASIG5V.n3197 0.019716
R54387 ASIG5V.n4953 ASIG5V.n4952 0.019716
R54388 ASIG5V.n4958 ASIG5V.n3196 0.019716
R54389 ASIG5V.n4958 ASIG5V.n4957 0.019716
R54390 ASIG5V.n4964 ASIG5V.n3195 0.019716
R54391 ASIG5V.n4965 ASIG5V.n4964 0.019716
R54392 ASIG5V.n4970 ASIG5V.n3194 0.019716
R54393 ASIG5V.n4970 ASIG5V.n4969 0.019716
R54394 ASIG5V.n4976 ASIG5V.n3193 0.019716
R54395 ASIG5V.n4977 ASIG5V.n4976 0.019716
R54396 ASIG5V.n4982 ASIG5V.n3192 0.019716
R54397 ASIG5V.n4982 ASIG5V.n4981 0.019716
R54398 ASIG5V.n4988 ASIG5V.n3191 0.019716
R54399 ASIG5V.n4989 ASIG5V.n4988 0.019716
R54400 ASIG5V.n4994 ASIG5V.n3190 0.019716
R54401 ASIG5V.n4994 ASIG5V.n4993 0.019716
R54402 ASIG5V.n5000 ASIG5V.n3189 0.019716
R54403 ASIG5V.n5001 ASIG5V.n5000 0.019716
R54404 ASIG5V.n5006 ASIG5V.n3188 0.019716
R54405 ASIG5V.n5006 ASIG5V.n5005 0.019716
R54406 ASIG5V.n5012 ASIG5V.n3187 0.019716
R54407 ASIG5V.n5013 ASIG5V.n5012 0.019716
R54408 ASIG5V.n5018 ASIG5V.n3186 0.019716
R54409 ASIG5V.n5018 ASIG5V.n5017 0.019716
R54410 ASIG5V.n5024 ASIG5V.n3185 0.019716
R54411 ASIG5V.n5025 ASIG5V.n5024 0.019716
R54412 ASIG5V.n5030 ASIG5V.n3184 0.019716
R54413 ASIG5V.n5030 ASIG5V.n5029 0.019716
R54414 ASIG5V.n5036 ASIG5V.n3183 0.019716
R54415 ASIG5V.n5037 ASIG5V.n5036 0.019716
R54416 ASIG5V.n5042 ASIG5V.n3182 0.019716
R54417 ASIG5V.n5042 ASIG5V.n5041 0.019716
R54418 ASIG5V.n5048 ASIG5V.n3181 0.019716
R54419 ASIG5V.n5049 ASIG5V.n5048 0.019716
R54420 ASIG5V.n5054 ASIG5V.n3180 0.019716
R54421 ASIG5V.n5054 ASIG5V.n5053 0.019716
R54422 ASIG5V.n5061 ASIG5V.n3179 0.019716
R54423 ASIG5V.n5062 ASIG5V.n5061 0.019716
R54424 ASIG5V.n9484 ASIG5V.n9483 0.019716
R54425 ASIG5V.n9491 ASIG5V.n5115 0.019716
R54426 ASIG5V.n9492 ASIG5V.n9491 0.019716
R54427 ASIG5V.n9497 ASIG5V.n5114 0.019716
R54428 ASIG5V.n9497 ASIG5V.n9496 0.019716
R54429 ASIG5V.n9503 ASIG5V.n5113 0.019716
R54430 ASIG5V.n9504 ASIG5V.n9503 0.019716
R54431 ASIG5V.n9509 ASIG5V.n5112 0.019716
R54432 ASIG5V.n9509 ASIG5V.n9508 0.019716
R54433 ASIG5V.n9515 ASIG5V.n5111 0.019716
R54434 ASIG5V.n9516 ASIG5V.n9515 0.019716
R54435 ASIG5V.n9521 ASIG5V.n5110 0.019716
R54436 ASIG5V.n9521 ASIG5V.n9520 0.019716
R54437 ASIG5V.n9527 ASIG5V.n5109 0.019716
R54438 ASIG5V.n9528 ASIG5V.n9527 0.019716
R54439 ASIG5V.n9533 ASIG5V.n5108 0.019716
R54440 ASIG5V.n9533 ASIG5V.n9532 0.019716
R54441 ASIG5V.n9539 ASIG5V.n5107 0.019716
R54442 ASIG5V.n9540 ASIG5V.n9539 0.019716
R54443 ASIG5V.n9545 ASIG5V.n5106 0.019716
R54444 ASIG5V.n9545 ASIG5V.n9544 0.019716
R54445 ASIG5V.n9551 ASIG5V.n5105 0.019716
R54446 ASIG5V.n9552 ASIG5V.n9551 0.019716
R54447 ASIG5V.n9557 ASIG5V.n5104 0.019716
R54448 ASIG5V.n9557 ASIG5V.n9556 0.019716
R54449 ASIG5V.n9563 ASIG5V.n5103 0.019716
R54450 ASIG5V.n9564 ASIG5V.n9563 0.019716
R54451 ASIG5V.n9569 ASIG5V.n5102 0.019716
R54452 ASIG5V.n9569 ASIG5V.n9568 0.019716
R54453 ASIG5V.n9575 ASIG5V.n5101 0.019716
R54454 ASIG5V.n9576 ASIG5V.n9575 0.019716
R54455 ASIG5V.n9581 ASIG5V.n5100 0.019716
R54456 ASIG5V.n9581 ASIG5V.n9580 0.019716
R54457 ASIG5V.n9587 ASIG5V.n5099 0.019716
R54458 ASIG5V.n9588 ASIG5V.n9587 0.019716
R54459 ASIG5V.n9593 ASIG5V.n5098 0.019716
R54460 ASIG5V.n9593 ASIG5V.n9592 0.019716
R54461 ASIG5V.n9599 ASIG5V.n5097 0.019716
R54462 ASIG5V.n9600 ASIG5V.n9599 0.019716
R54463 ASIG5V.n9605 ASIG5V.n5096 0.019716
R54464 ASIG5V.n9605 ASIG5V.n9604 0.019716
R54465 ASIG5V.n9611 ASIG5V.n5095 0.019716
R54466 ASIG5V.n9612 ASIG5V.n9611 0.019716
R54467 ASIG5V.n9617 ASIG5V.n5094 0.019716
R54468 ASIG5V.n9617 ASIG5V.n9616 0.019716
R54469 ASIG5V.n9623 ASIG5V.n5093 0.019716
R54470 ASIG5V.n9624 ASIG5V.n9623 0.019716
R54471 ASIG5V.n9629 ASIG5V.n5092 0.019716
R54472 ASIG5V.n9629 ASIG5V.n9628 0.019716
R54473 ASIG5V.n9635 ASIG5V.n5091 0.019716
R54474 ASIG5V.n9636 ASIG5V.n9635 0.019716
R54475 ASIG5V.n9641 ASIG5V.n5090 0.019716
R54476 ASIG5V.n9641 ASIG5V.n9640 0.019716
R54477 ASIG5V.n9647 ASIG5V.n5089 0.019716
R54478 ASIG5V.n9648 ASIG5V.n9647 0.019716
R54479 ASIG5V.n9653 ASIG5V.n5088 0.019716
R54480 ASIG5V.n9653 ASIG5V.n9652 0.019716
R54481 ASIG5V.n9659 ASIG5V.n5087 0.019716
R54482 ASIG5V.n9660 ASIG5V.n9659 0.019716
R54483 ASIG5V.n9665 ASIG5V.n5086 0.019716
R54484 ASIG5V.n9665 ASIG5V.n9664 0.019716
R54485 ASIG5V.n9671 ASIG5V.n5085 0.019716
R54486 ASIG5V.n9672 ASIG5V.n9671 0.019716
R54487 ASIG5V.n9677 ASIG5V.n5084 0.019716
R54488 ASIG5V.n9677 ASIG5V.n9676 0.019716
R54489 ASIG5V.n9683 ASIG5V.n5083 0.019716
R54490 ASIG5V.n9684 ASIG5V.n9683 0.019716
R54491 ASIG5V.n9689 ASIG5V.n5082 0.019716
R54492 ASIG5V.n9689 ASIG5V.n9688 0.019716
R54493 ASIG5V.n9695 ASIG5V.n5081 0.019716
R54494 ASIG5V.n9696 ASIG5V.n9695 0.019716
R54495 ASIG5V.n9701 ASIG5V.n5080 0.019716
R54496 ASIG5V.n9701 ASIG5V.n9700 0.019716
R54497 ASIG5V.n9707 ASIG5V.n5079 0.019716
R54498 ASIG5V.n9708 ASIG5V.n9707 0.019716
R54499 ASIG5V.n9713 ASIG5V.n5078 0.019716
R54500 ASIG5V.n9713 ASIG5V.n9712 0.019716
R54501 ASIG5V.n9719 ASIG5V.n5077 0.019716
R54502 ASIG5V.n9720 ASIG5V.n9719 0.019716
R54503 ASIG5V.n9725 ASIG5V.n5076 0.019716
R54504 ASIG5V.n9725 ASIG5V.n9724 0.019716
R54505 ASIG5V.n9731 ASIG5V.n5075 0.019716
R54506 ASIG5V.n9732 ASIG5V.n9731 0.019716
R54507 ASIG5V.n5212 ASIG5V.n5211 0.019716
R54508 ASIG5V.n5219 ASIG5V.n5164 0.019716
R54509 ASIG5V.n5220 ASIG5V.n5219 0.019716
R54510 ASIG5V.n5225 ASIG5V.n5163 0.019716
R54511 ASIG5V.n5225 ASIG5V.n5224 0.019716
R54512 ASIG5V.n5231 ASIG5V.n5162 0.019716
R54513 ASIG5V.n5232 ASIG5V.n5231 0.019716
R54514 ASIG5V.n5237 ASIG5V.n5161 0.019716
R54515 ASIG5V.n5237 ASIG5V.n5236 0.019716
R54516 ASIG5V.n5243 ASIG5V.n5160 0.019716
R54517 ASIG5V.n5244 ASIG5V.n5243 0.019716
R54518 ASIG5V.n5249 ASIG5V.n5159 0.019716
R54519 ASIG5V.n5249 ASIG5V.n5248 0.019716
R54520 ASIG5V.n5255 ASIG5V.n5158 0.019716
R54521 ASIG5V.n5256 ASIG5V.n5255 0.019716
R54522 ASIG5V.n5261 ASIG5V.n5157 0.019716
R54523 ASIG5V.n5261 ASIG5V.n5260 0.019716
R54524 ASIG5V.n5267 ASIG5V.n5156 0.019716
R54525 ASIG5V.n5268 ASIG5V.n5267 0.019716
R54526 ASIG5V.n5273 ASIG5V.n5155 0.019716
R54527 ASIG5V.n5273 ASIG5V.n5272 0.019716
R54528 ASIG5V.n5279 ASIG5V.n5154 0.019716
R54529 ASIG5V.n5280 ASIG5V.n5279 0.019716
R54530 ASIG5V.n5285 ASIG5V.n5153 0.019716
R54531 ASIG5V.n5285 ASIG5V.n5284 0.019716
R54532 ASIG5V.n5291 ASIG5V.n5152 0.019716
R54533 ASIG5V.n5292 ASIG5V.n5291 0.019716
R54534 ASIG5V.n5297 ASIG5V.n5151 0.019716
R54535 ASIG5V.n5297 ASIG5V.n5296 0.019716
R54536 ASIG5V.n5303 ASIG5V.n5150 0.019716
R54537 ASIG5V.n5304 ASIG5V.n5303 0.019716
R54538 ASIG5V.n5309 ASIG5V.n5149 0.019716
R54539 ASIG5V.n5309 ASIG5V.n5308 0.019716
R54540 ASIG5V.n5315 ASIG5V.n5148 0.019716
R54541 ASIG5V.n5316 ASIG5V.n5315 0.019716
R54542 ASIG5V.n5321 ASIG5V.n5147 0.019716
R54543 ASIG5V.n5321 ASIG5V.n5320 0.019716
R54544 ASIG5V.n5327 ASIG5V.n5146 0.019716
R54545 ASIG5V.n5328 ASIG5V.n5327 0.019716
R54546 ASIG5V.n5333 ASIG5V.n5145 0.019716
R54547 ASIG5V.n5333 ASIG5V.n5332 0.019716
R54548 ASIG5V.n5339 ASIG5V.n5144 0.019716
R54549 ASIG5V.n5340 ASIG5V.n5339 0.019716
R54550 ASIG5V.n5345 ASIG5V.n5143 0.019716
R54551 ASIG5V.n5345 ASIG5V.n5344 0.019716
R54552 ASIG5V.n5351 ASIG5V.n5142 0.019716
R54553 ASIG5V.n5352 ASIG5V.n5351 0.019716
R54554 ASIG5V.n5357 ASIG5V.n5141 0.019716
R54555 ASIG5V.n5357 ASIG5V.n5356 0.019716
R54556 ASIG5V.n5363 ASIG5V.n5140 0.019716
R54557 ASIG5V.n5364 ASIG5V.n5363 0.019716
R54558 ASIG5V.n5369 ASIG5V.n5139 0.019716
R54559 ASIG5V.n5369 ASIG5V.n5368 0.019716
R54560 ASIG5V.n5375 ASIG5V.n5138 0.019716
R54561 ASIG5V.n5376 ASIG5V.n5375 0.019716
R54562 ASIG5V.n5381 ASIG5V.n5137 0.019716
R54563 ASIG5V.n5381 ASIG5V.n5380 0.019716
R54564 ASIG5V.n5387 ASIG5V.n5136 0.019716
R54565 ASIG5V.n5388 ASIG5V.n5387 0.019716
R54566 ASIG5V.n5393 ASIG5V.n5135 0.019716
R54567 ASIG5V.n5393 ASIG5V.n5392 0.019716
R54568 ASIG5V.n5399 ASIG5V.n5134 0.019716
R54569 ASIG5V.n5400 ASIG5V.n5399 0.019716
R54570 ASIG5V.n5405 ASIG5V.n5133 0.019716
R54571 ASIG5V.n5405 ASIG5V.n5404 0.019716
R54572 ASIG5V.n5411 ASIG5V.n5132 0.019716
R54573 ASIG5V.n5412 ASIG5V.n5411 0.019716
R54574 ASIG5V.n5417 ASIG5V.n5131 0.019716
R54575 ASIG5V.n5417 ASIG5V.n5416 0.019716
R54576 ASIG5V.n5423 ASIG5V.n5130 0.019716
R54577 ASIG5V.n5424 ASIG5V.n5423 0.019716
R54578 ASIG5V.n5429 ASIG5V.n5129 0.019716
R54579 ASIG5V.n5429 ASIG5V.n5428 0.019716
R54580 ASIG5V.n5435 ASIG5V.n5128 0.019716
R54581 ASIG5V.n5436 ASIG5V.n5435 0.019716
R54582 ASIG5V.n5441 ASIG5V.n5127 0.019716
R54583 ASIG5V.n5441 ASIG5V.n5440 0.019716
R54584 ASIG5V.n5447 ASIG5V.n5126 0.019716
R54585 ASIG5V.n5448 ASIG5V.n5447 0.019716
R54586 ASIG5V.n5453 ASIG5V.n5125 0.019716
R54587 ASIG5V.n5453 ASIG5V.n5452 0.019716
R54588 ASIG5V.n9429 ASIG5V.n5124 0.019716
R54589 ASIG5V.n9430 ASIG5V.n9429 0.019716
R54590 ASIG5V.n9418 ASIG5V.n5507 0.019716
R54591 ASIG5V.n7956 ASIG5V.n5552 0.019716
R54592 ASIG5V.n7956 ASIG5V.n5505 0.019716
R54593 ASIG5V.n7718 ASIG5V.n5551 0.019716
R54594 ASIG5V.n7718 ASIG5V.n5504 0.019716
R54595 ASIG5V.n7947 ASIG5V.n5550 0.019716
R54596 ASIG5V.n7947 ASIG5V.n5503 0.019716
R54597 ASIG5V.n7721 ASIG5V.n5549 0.019716
R54598 ASIG5V.n7721 ASIG5V.n5502 0.019716
R54599 ASIG5V.n7938 ASIG5V.n5548 0.019716
R54600 ASIG5V.n7938 ASIG5V.n5501 0.019716
R54601 ASIG5V.n7724 ASIG5V.n5547 0.019716
R54602 ASIG5V.n7724 ASIG5V.n5500 0.019716
R54603 ASIG5V.n7929 ASIG5V.n5546 0.019716
R54604 ASIG5V.n7929 ASIG5V.n5499 0.019716
R54605 ASIG5V.n7727 ASIG5V.n5545 0.019716
R54606 ASIG5V.n7727 ASIG5V.n5498 0.019716
R54607 ASIG5V.n7920 ASIG5V.n5544 0.019716
R54608 ASIG5V.n7920 ASIG5V.n5497 0.019716
R54609 ASIG5V.n7730 ASIG5V.n5543 0.019716
R54610 ASIG5V.n7730 ASIG5V.n5496 0.019716
R54611 ASIG5V.n7911 ASIG5V.n5542 0.019716
R54612 ASIG5V.n7911 ASIG5V.n5495 0.019716
R54613 ASIG5V.n7733 ASIG5V.n5541 0.019716
R54614 ASIG5V.n7733 ASIG5V.n5494 0.019716
R54615 ASIG5V.n7902 ASIG5V.n5540 0.019716
R54616 ASIG5V.n7902 ASIG5V.n5493 0.019716
R54617 ASIG5V.n7736 ASIG5V.n5539 0.019716
R54618 ASIG5V.n7736 ASIG5V.n5492 0.019716
R54619 ASIG5V.n7893 ASIG5V.n5538 0.019716
R54620 ASIG5V.n7893 ASIG5V.n5491 0.019716
R54621 ASIG5V.n7739 ASIG5V.n5537 0.019716
R54622 ASIG5V.n7739 ASIG5V.n5490 0.019716
R54623 ASIG5V.n7884 ASIG5V.n5536 0.019716
R54624 ASIG5V.n7884 ASIG5V.n5489 0.019716
R54625 ASIG5V.n7742 ASIG5V.n5535 0.019716
R54626 ASIG5V.n7742 ASIG5V.n5488 0.019716
R54627 ASIG5V.n7875 ASIG5V.n5534 0.019716
R54628 ASIG5V.n7875 ASIG5V.n5487 0.019716
R54629 ASIG5V.n7745 ASIG5V.n5533 0.019716
R54630 ASIG5V.n7745 ASIG5V.n5486 0.019716
R54631 ASIG5V.n7866 ASIG5V.n5532 0.019716
R54632 ASIG5V.n7866 ASIG5V.n5485 0.019716
R54633 ASIG5V.n7748 ASIG5V.n5531 0.019716
R54634 ASIG5V.n7748 ASIG5V.n5484 0.019716
R54635 ASIG5V.n7857 ASIG5V.n5530 0.019716
R54636 ASIG5V.n7857 ASIG5V.n5483 0.019716
R54637 ASIG5V.n7751 ASIG5V.n5529 0.019716
R54638 ASIG5V.n7751 ASIG5V.n5482 0.019716
R54639 ASIG5V.n7848 ASIG5V.n5528 0.019716
R54640 ASIG5V.n7848 ASIG5V.n5481 0.019716
R54641 ASIG5V.n7754 ASIG5V.n5527 0.019716
R54642 ASIG5V.n7754 ASIG5V.n5480 0.019716
R54643 ASIG5V.n7839 ASIG5V.n5526 0.019716
R54644 ASIG5V.n7839 ASIG5V.n5479 0.019716
R54645 ASIG5V.n7757 ASIG5V.n5525 0.019716
R54646 ASIG5V.n7757 ASIG5V.n5478 0.019716
R54647 ASIG5V.n7830 ASIG5V.n5524 0.019716
R54648 ASIG5V.n7830 ASIG5V.n5477 0.019716
R54649 ASIG5V.n7760 ASIG5V.n5523 0.019716
R54650 ASIG5V.n7760 ASIG5V.n5476 0.019716
R54651 ASIG5V.n7821 ASIG5V.n5522 0.019716
R54652 ASIG5V.n7821 ASIG5V.n5475 0.019716
R54653 ASIG5V.n7763 ASIG5V.n5521 0.019716
R54654 ASIG5V.n7763 ASIG5V.n5474 0.019716
R54655 ASIG5V.n7812 ASIG5V.n5520 0.019716
R54656 ASIG5V.n7812 ASIG5V.n5473 0.019716
R54657 ASIG5V.n7766 ASIG5V.n5519 0.019716
R54658 ASIG5V.n7766 ASIG5V.n5472 0.019716
R54659 ASIG5V.n7803 ASIG5V.n5518 0.019716
R54660 ASIG5V.n7803 ASIG5V.n5471 0.019716
R54661 ASIG5V.n7769 ASIG5V.n5517 0.019716
R54662 ASIG5V.n7769 ASIG5V.n5470 0.019716
R54663 ASIG5V.n7794 ASIG5V.n5516 0.019716
R54664 ASIG5V.n7794 ASIG5V.n5469 0.019716
R54665 ASIG5V.n7772 ASIG5V.n5515 0.019716
R54666 ASIG5V.n7772 ASIG5V.n5468 0.019716
R54667 ASIG5V.n7785 ASIG5V.n5514 0.019716
R54668 ASIG5V.n7785 ASIG5V.n5467 0.019716
R54669 ASIG5V.n7775 ASIG5V.n5513 0.019716
R54670 ASIG5V.n7775 ASIG5V.n5466 0.019716
R54671 ASIG5V.n5555 ASIG5V.n5512 0.019716
R54672 ASIG5V.n5555 ASIG5V.n5465 0.019716
R54673 ASIG5V.n5904 ASIG5V.n5903 0.019716
R54674 ASIG5V.n5902 ASIG5V.n5901 0.019716
R54675 ASIG5V.n5901 ASIG5V.n5575 0.019716
R54676 ASIG5V.n5895 ASIG5V.n5580 0.019716
R54677 ASIG5V.n5895 ASIG5V.n5894 0.019716
R54678 ASIG5V.n5892 ASIG5V.n5891 0.019716
R54679 ASIG5V.n5891 ASIG5V.n5581 0.019716
R54680 ASIG5V.n5885 ASIG5V.n5586 0.019716
R54681 ASIG5V.n5885 ASIG5V.n5884 0.019716
R54682 ASIG5V.n5882 ASIG5V.n5881 0.019716
R54683 ASIG5V.n5881 ASIG5V.n5587 0.019716
R54684 ASIG5V.n5875 ASIG5V.n5592 0.019716
R54685 ASIG5V.n5875 ASIG5V.n5874 0.019716
R54686 ASIG5V.n5872 ASIG5V.n5871 0.019716
R54687 ASIG5V.n5871 ASIG5V.n5593 0.019716
R54688 ASIG5V.n5865 ASIG5V.n5598 0.019716
R54689 ASIG5V.n5865 ASIG5V.n5864 0.019716
R54690 ASIG5V.n5862 ASIG5V.n5861 0.019716
R54691 ASIG5V.n5861 ASIG5V.n5599 0.019716
R54692 ASIG5V.n5855 ASIG5V.n5604 0.019716
R54693 ASIG5V.n5855 ASIG5V.n5854 0.019716
R54694 ASIG5V.n5852 ASIG5V.n5851 0.019716
R54695 ASIG5V.n5851 ASIG5V.n5605 0.019716
R54696 ASIG5V.n5845 ASIG5V.n5610 0.019716
R54697 ASIG5V.n5845 ASIG5V.n5844 0.019716
R54698 ASIG5V.n5842 ASIG5V.n5841 0.019716
R54699 ASIG5V.n5841 ASIG5V.n5611 0.019716
R54700 ASIG5V.n5835 ASIG5V.n5616 0.019716
R54701 ASIG5V.n5835 ASIG5V.n5834 0.019716
R54702 ASIG5V.n5832 ASIG5V.n5831 0.019716
R54703 ASIG5V.n5831 ASIG5V.n5617 0.019716
R54704 ASIG5V.n5825 ASIG5V.n5622 0.019716
R54705 ASIG5V.n5825 ASIG5V.n5824 0.019716
R54706 ASIG5V.n5822 ASIG5V.n5821 0.019716
R54707 ASIG5V.n5821 ASIG5V.n5623 0.019716
R54708 ASIG5V.n5815 ASIG5V.n5628 0.019716
R54709 ASIG5V.n5815 ASIG5V.n5814 0.019716
R54710 ASIG5V.n5812 ASIG5V.n5811 0.019716
R54711 ASIG5V.n5811 ASIG5V.n5629 0.019716
R54712 ASIG5V.n5805 ASIG5V.n5634 0.019716
R54713 ASIG5V.n5805 ASIG5V.n5804 0.019716
R54714 ASIG5V.n5802 ASIG5V.n5801 0.019716
R54715 ASIG5V.n5801 ASIG5V.n5635 0.019716
R54716 ASIG5V.n5795 ASIG5V.n5640 0.019716
R54717 ASIG5V.n5795 ASIG5V.n5794 0.019716
R54718 ASIG5V.n5792 ASIG5V.n5791 0.019716
R54719 ASIG5V.n5791 ASIG5V.n5641 0.019716
R54720 ASIG5V.n5785 ASIG5V.n5646 0.019716
R54721 ASIG5V.n5785 ASIG5V.n5784 0.019716
R54722 ASIG5V.n5782 ASIG5V.n5781 0.019716
R54723 ASIG5V.n5781 ASIG5V.n5647 0.019716
R54724 ASIG5V.n5775 ASIG5V.n5652 0.019716
R54725 ASIG5V.n5775 ASIG5V.n5774 0.019716
R54726 ASIG5V.n5772 ASIG5V.n5771 0.019716
R54727 ASIG5V.n5771 ASIG5V.n5653 0.019716
R54728 ASIG5V.n5765 ASIG5V.n5658 0.019716
R54729 ASIG5V.n5765 ASIG5V.n5764 0.019716
R54730 ASIG5V.n5762 ASIG5V.n5761 0.019716
R54731 ASIG5V.n5761 ASIG5V.n5659 0.019716
R54732 ASIG5V.n5755 ASIG5V.n5664 0.019716
R54733 ASIG5V.n5755 ASIG5V.n5754 0.019716
R54734 ASIG5V.n5752 ASIG5V.n5751 0.019716
R54735 ASIG5V.n5751 ASIG5V.n5665 0.019716
R54736 ASIG5V.n5745 ASIG5V.n5670 0.019716
R54737 ASIG5V.n5745 ASIG5V.n5744 0.019716
R54738 ASIG5V.n5742 ASIG5V.n5741 0.019716
R54739 ASIG5V.n5741 ASIG5V.n5671 0.019716
R54740 ASIG5V.n5735 ASIG5V.n5676 0.019716
R54741 ASIG5V.n5735 ASIG5V.n5734 0.019716
R54742 ASIG5V.n5732 ASIG5V.n5731 0.019716
R54743 ASIG5V.n5731 ASIG5V.n5677 0.019716
R54744 ASIG5V.n5725 ASIG5V.n5682 0.019716
R54745 ASIG5V.n5725 ASIG5V.n5724 0.019716
R54746 ASIG5V.n5722 ASIG5V.n5721 0.019716
R54747 ASIG5V.n5721 ASIG5V.n5683 0.019716
R54748 ASIG5V.n5715 ASIG5V.n5688 0.019716
R54749 ASIG5V.n5715 ASIG5V.n5714 0.019716
R54750 ASIG5V.n5712 ASIG5V.n5711 0.019716
R54751 ASIG5V.n5711 ASIG5V.n5689 0.019716
R54752 ASIG5V.n5705 ASIG5V.n5694 0.019716
R54753 ASIG5V.n5705 ASIG5V.n5704 0.019716
R54754 ASIG5V.n5702 ASIG5V.n5701 0.019716
R54755 ASIG5V.n5701 ASIG5V.n5695 0.019716
R54756 ASIG5V.n9395 ASIG5V.n5955 0.019716
R54757 ASIG5V.n6061 ASIG5V.n5998 0.019716
R54758 ASIG5V.n6061 ASIG5V.n5953 0.019716
R54759 ASIG5V.n6070 ASIG5V.n5997 0.019716
R54760 ASIG5V.n6070 ASIG5V.n5952 0.019716
R54761 ASIG5V.n6058 ASIG5V.n5996 0.019716
R54762 ASIG5V.n6058 ASIG5V.n5951 0.019716
R54763 ASIG5V.n6079 ASIG5V.n5995 0.019716
R54764 ASIG5V.n6079 ASIG5V.n5950 0.019716
R54765 ASIG5V.n6055 ASIG5V.n5994 0.019716
R54766 ASIG5V.n6055 ASIG5V.n5949 0.019716
R54767 ASIG5V.n6088 ASIG5V.n5993 0.019716
R54768 ASIG5V.n6088 ASIG5V.n5948 0.019716
R54769 ASIG5V.n6052 ASIG5V.n5992 0.019716
R54770 ASIG5V.n6052 ASIG5V.n5947 0.019716
R54771 ASIG5V.n6097 ASIG5V.n5991 0.019716
R54772 ASIG5V.n6097 ASIG5V.n5946 0.019716
R54773 ASIG5V.n6049 ASIG5V.n5990 0.019716
R54774 ASIG5V.n6049 ASIG5V.n5945 0.019716
R54775 ASIG5V.n6106 ASIG5V.n5989 0.019716
R54776 ASIG5V.n6106 ASIG5V.n5944 0.019716
R54777 ASIG5V.n6046 ASIG5V.n5988 0.019716
R54778 ASIG5V.n6046 ASIG5V.n5943 0.019716
R54779 ASIG5V.n6115 ASIG5V.n5987 0.019716
R54780 ASIG5V.n6115 ASIG5V.n5942 0.019716
R54781 ASIG5V.n6043 ASIG5V.n5986 0.019716
R54782 ASIG5V.n6043 ASIG5V.n5941 0.019716
R54783 ASIG5V.n6124 ASIG5V.n5985 0.019716
R54784 ASIG5V.n6124 ASIG5V.n5940 0.019716
R54785 ASIG5V.n6040 ASIG5V.n5984 0.019716
R54786 ASIG5V.n6040 ASIG5V.n5939 0.019716
R54787 ASIG5V.n6133 ASIG5V.n5983 0.019716
R54788 ASIG5V.n6133 ASIG5V.n5938 0.019716
R54789 ASIG5V.n6037 ASIG5V.n5982 0.019716
R54790 ASIG5V.n6037 ASIG5V.n5937 0.019716
R54791 ASIG5V.n6142 ASIG5V.n5981 0.019716
R54792 ASIG5V.n6142 ASIG5V.n5936 0.019716
R54793 ASIG5V.n6034 ASIG5V.n5980 0.019716
R54794 ASIG5V.n6034 ASIG5V.n5935 0.019716
R54795 ASIG5V.n6151 ASIG5V.n5979 0.019716
R54796 ASIG5V.n6151 ASIG5V.n5934 0.019716
R54797 ASIG5V.n6031 ASIG5V.n5978 0.019716
R54798 ASIG5V.n6031 ASIG5V.n5933 0.019716
R54799 ASIG5V.n6160 ASIG5V.n5977 0.019716
R54800 ASIG5V.n6160 ASIG5V.n5932 0.019716
R54801 ASIG5V.n6028 ASIG5V.n5976 0.019716
R54802 ASIG5V.n6028 ASIG5V.n5931 0.019716
R54803 ASIG5V.n6169 ASIG5V.n5975 0.019716
R54804 ASIG5V.n6169 ASIG5V.n5930 0.019716
R54805 ASIG5V.n6025 ASIG5V.n5974 0.019716
R54806 ASIG5V.n6025 ASIG5V.n5929 0.019716
R54807 ASIG5V.n6178 ASIG5V.n5973 0.019716
R54808 ASIG5V.n6178 ASIG5V.n5928 0.019716
R54809 ASIG5V.n6022 ASIG5V.n5972 0.019716
R54810 ASIG5V.n6022 ASIG5V.n5927 0.019716
R54811 ASIG5V.n6187 ASIG5V.n5971 0.019716
R54812 ASIG5V.n6187 ASIG5V.n5926 0.019716
R54813 ASIG5V.n6019 ASIG5V.n5970 0.019716
R54814 ASIG5V.n6019 ASIG5V.n5925 0.019716
R54815 ASIG5V.n6196 ASIG5V.n5969 0.019716
R54816 ASIG5V.n6196 ASIG5V.n5924 0.019716
R54817 ASIG5V.n6016 ASIG5V.n5968 0.019716
R54818 ASIG5V.n6016 ASIG5V.n5923 0.019716
R54819 ASIG5V.n6205 ASIG5V.n5967 0.019716
R54820 ASIG5V.n6205 ASIG5V.n5922 0.019716
R54821 ASIG5V.n6013 ASIG5V.n5966 0.019716
R54822 ASIG5V.n6013 ASIG5V.n5921 0.019716
R54823 ASIG5V.n6214 ASIG5V.n5965 0.019716
R54824 ASIG5V.n6214 ASIG5V.n5920 0.019716
R54825 ASIG5V.n6010 ASIG5V.n5964 0.019716
R54826 ASIG5V.n6010 ASIG5V.n5919 0.019716
R54827 ASIG5V.n6223 ASIG5V.n5963 0.019716
R54828 ASIG5V.n6223 ASIG5V.n5918 0.019716
R54829 ASIG5V.n6007 ASIG5V.n5962 0.019716
R54830 ASIG5V.n6007 ASIG5V.n5917 0.019716
R54831 ASIG5V.n6232 ASIG5V.n5961 0.019716
R54832 ASIG5V.n6232 ASIG5V.n5916 0.019716
R54833 ASIG5V.n6004 ASIG5V.n5960 0.019716
R54834 ASIG5V.n6004 ASIG5V.n5915 0.019716
R54835 ASIG5V.n6241 ASIG5V.n5959 0.019716
R54836 ASIG5V.n6241 ASIG5V.n5914 0.019716
R54837 ASIG5V.n6001 ASIG5V.n5958 0.019716
R54838 ASIG5V.n6001 ASIG5V.n5913 0.019716
R54839 ASIG5V.n9381 ASIG5V.n6307 0.019716
R54840 ASIG5V.n6413 ASIG5V.n6351 0.019716
R54841 ASIG5V.n6413 ASIG5V.n6305 0.019716
R54842 ASIG5V.n9199 ASIG5V.n6350 0.019716
R54843 ASIG5V.n9199 ASIG5V.n6304 0.019716
R54844 ASIG5V.n6410 ASIG5V.n6349 0.019716
R54845 ASIG5V.n6410 ASIG5V.n6303 0.019716
R54846 ASIG5V.n9208 ASIG5V.n6348 0.019716
R54847 ASIG5V.n9208 ASIG5V.n6302 0.019716
R54848 ASIG5V.n6407 ASIG5V.n6347 0.019716
R54849 ASIG5V.n6407 ASIG5V.n6301 0.019716
R54850 ASIG5V.n9217 ASIG5V.n6346 0.019716
R54851 ASIG5V.n9217 ASIG5V.n6300 0.019716
R54852 ASIG5V.n6404 ASIG5V.n6345 0.019716
R54853 ASIG5V.n6404 ASIG5V.n6299 0.019716
R54854 ASIG5V.n9226 ASIG5V.n6344 0.019716
R54855 ASIG5V.n9226 ASIG5V.n6298 0.019716
R54856 ASIG5V.n6401 ASIG5V.n6343 0.019716
R54857 ASIG5V.n6401 ASIG5V.n6297 0.019716
R54858 ASIG5V.n9235 ASIG5V.n6342 0.019716
R54859 ASIG5V.n9235 ASIG5V.n6296 0.019716
R54860 ASIG5V.n6398 ASIG5V.n6341 0.019716
R54861 ASIG5V.n6398 ASIG5V.n6295 0.019716
R54862 ASIG5V.n9244 ASIG5V.n6340 0.019716
R54863 ASIG5V.n9244 ASIG5V.n6294 0.019716
R54864 ASIG5V.n6395 ASIG5V.n6339 0.019716
R54865 ASIG5V.n6395 ASIG5V.n6293 0.019716
R54866 ASIG5V.n9253 ASIG5V.n6338 0.019716
R54867 ASIG5V.n9253 ASIG5V.n6292 0.019716
R54868 ASIG5V.n6392 ASIG5V.n6337 0.019716
R54869 ASIG5V.n6392 ASIG5V.n6291 0.019716
R54870 ASIG5V.n9262 ASIG5V.n6336 0.019716
R54871 ASIG5V.n9262 ASIG5V.n6290 0.019716
R54872 ASIG5V.n6389 ASIG5V.n6335 0.019716
R54873 ASIG5V.n6389 ASIG5V.n6289 0.019716
R54874 ASIG5V.n9271 ASIG5V.n6334 0.019716
R54875 ASIG5V.n9271 ASIG5V.n6288 0.019716
R54876 ASIG5V.n6386 ASIG5V.n6333 0.019716
R54877 ASIG5V.n6386 ASIG5V.n6287 0.019716
R54878 ASIG5V.n9280 ASIG5V.n6332 0.019716
R54879 ASIG5V.n9280 ASIG5V.n6286 0.019716
R54880 ASIG5V.n6383 ASIG5V.n6331 0.019716
R54881 ASIG5V.n6383 ASIG5V.n6285 0.019716
R54882 ASIG5V.n9289 ASIG5V.n6330 0.019716
R54883 ASIG5V.n9289 ASIG5V.n6284 0.019716
R54884 ASIG5V.n6380 ASIG5V.n6329 0.019716
R54885 ASIG5V.n6380 ASIG5V.n6283 0.019716
R54886 ASIG5V.n9298 ASIG5V.n6328 0.019716
R54887 ASIG5V.n9298 ASIG5V.n6282 0.019716
R54888 ASIG5V.n6377 ASIG5V.n6327 0.019716
R54889 ASIG5V.n6377 ASIG5V.n6281 0.019716
R54890 ASIG5V.n9307 ASIG5V.n6326 0.019716
R54891 ASIG5V.n9307 ASIG5V.n6280 0.019716
R54892 ASIG5V.n6374 ASIG5V.n6325 0.019716
R54893 ASIG5V.n6374 ASIG5V.n6279 0.019716
R54894 ASIG5V.n9316 ASIG5V.n6324 0.019716
R54895 ASIG5V.n9316 ASIG5V.n6278 0.019716
R54896 ASIG5V.n6371 ASIG5V.n6323 0.019716
R54897 ASIG5V.n6371 ASIG5V.n6277 0.019716
R54898 ASIG5V.n9325 ASIG5V.n6322 0.019716
R54899 ASIG5V.n9325 ASIG5V.n6276 0.019716
R54900 ASIG5V.n6368 ASIG5V.n6321 0.019716
R54901 ASIG5V.n6368 ASIG5V.n6275 0.019716
R54902 ASIG5V.n9334 ASIG5V.n6320 0.019716
R54903 ASIG5V.n9334 ASIG5V.n6274 0.019716
R54904 ASIG5V.n6365 ASIG5V.n6319 0.019716
R54905 ASIG5V.n6365 ASIG5V.n6273 0.019716
R54906 ASIG5V.n9343 ASIG5V.n6318 0.019716
R54907 ASIG5V.n9343 ASIG5V.n6272 0.019716
R54908 ASIG5V.n6362 ASIG5V.n6317 0.019716
R54909 ASIG5V.n6362 ASIG5V.n6271 0.019716
R54910 ASIG5V.n9352 ASIG5V.n6316 0.019716
R54911 ASIG5V.n9352 ASIG5V.n6270 0.019716
R54912 ASIG5V.n6359 ASIG5V.n6315 0.019716
R54913 ASIG5V.n6359 ASIG5V.n6269 0.019716
R54914 ASIG5V.n9361 ASIG5V.n6314 0.019716
R54915 ASIG5V.n9361 ASIG5V.n6268 0.019716
R54916 ASIG5V.n6356 ASIG5V.n6313 0.019716
R54917 ASIG5V.n6356 ASIG5V.n6267 0.019716
R54918 ASIG5V.n9370 ASIG5V.n6312 0.019716
R54919 ASIG5V.n9370 ASIG5V.n6266 0.019716
R54920 ASIG5V.n6353 ASIG5V.n6311 0.019716
R54921 ASIG5V.n6353 ASIG5V.n6265 0.019716
R54922 ASIG5V.n6531 ASIG5V.n6530 0.019716
R54923 ASIG5V.n8933 ASIG5V.n6486 0.019716
R54924 ASIG5V.n8934 ASIG5V.n8933 0.019716
R54925 ASIG5V.n8939 ASIG5V.n6485 0.019716
R54926 ASIG5V.n8939 ASIG5V.n8938 0.019716
R54927 ASIG5V.n8945 ASIG5V.n6484 0.019716
R54928 ASIG5V.n8946 ASIG5V.n8945 0.019716
R54929 ASIG5V.n8951 ASIG5V.n6483 0.019716
R54930 ASIG5V.n8951 ASIG5V.n8950 0.019716
R54931 ASIG5V.n8957 ASIG5V.n6482 0.019716
R54932 ASIG5V.n8958 ASIG5V.n8957 0.019716
R54933 ASIG5V.n8963 ASIG5V.n6481 0.019716
R54934 ASIG5V.n8963 ASIG5V.n8962 0.019716
R54935 ASIG5V.n8969 ASIG5V.n6480 0.019716
R54936 ASIG5V.n8970 ASIG5V.n8969 0.019716
R54937 ASIG5V.n8975 ASIG5V.n6479 0.019716
R54938 ASIG5V.n8975 ASIG5V.n8974 0.019716
R54939 ASIG5V.n8981 ASIG5V.n6478 0.019716
R54940 ASIG5V.n8982 ASIG5V.n8981 0.019716
R54941 ASIG5V.n8987 ASIG5V.n6477 0.019716
R54942 ASIG5V.n8987 ASIG5V.n8986 0.019716
R54943 ASIG5V.n8993 ASIG5V.n6476 0.019716
R54944 ASIG5V.n8994 ASIG5V.n8993 0.019716
R54945 ASIG5V.n8999 ASIG5V.n6475 0.019716
R54946 ASIG5V.n8999 ASIG5V.n8998 0.019716
R54947 ASIG5V.n9005 ASIG5V.n6474 0.019716
R54948 ASIG5V.n9006 ASIG5V.n9005 0.019716
R54949 ASIG5V.n9011 ASIG5V.n6473 0.019716
R54950 ASIG5V.n9011 ASIG5V.n9010 0.019716
R54951 ASIG5V.n9017 ASIG5V.n6472 0.019716
R54952 ASIG5V.n9018 ASIG5V.n9017 0.019716
R54953 ASIG5V.n9023 ASIG5V.n6471 0.019716
R54954 ASIG5V.n9023 ASIG5V.n9022 0.019716
R54955 ASIG5V.n9029 ASIG5V.n6470 0.019716
R54956 ASIG5V.n9030 ASIG5V.n9029 0.019716
R54957 ASIG5V.n9035 ASIG5V.n6469 0.019716
R54958 ASIG5V.n9035 ASIG5V.n9034 0.019716
R54959 ASIG5V.n9041 ASIG5V.n6468 0.019716
R54960 ASIG5V.n9042 ASIG5V.n9041 0.019716
R54961 ASIG5V.n9047 ASIG5V.n6467 0.019716
R54962 ASIG5V.n9047 ASIG5V.n9046 0.019716
R54963 ASIG5V.n9053 ASIG5V.n6466 0.019716
R54964 ASIG5V.n9054 ASIG5V.n9053 0.019716
R54965 ASIG5V.n9059 ASIG5V.n6465 0.019716
R54966 ASIG5V.n9059 ASIG5V.n9058 0.019716
R54967 ASIG5V.n9065 ASIG5V.n6464 0.019716
R54968 ASIG5V.n9066 ASIG5V.n9065 0.019716
R54969 ASIG5V.n9071 ASIG5V.n6463 0.019716
R54970 ASIG5V.n9071 ASIG5V.n9070 0.019716
R54971 ASIG5V.n9077 ASIG5V.n6462 0.019716
R54972 ASIG5V.n9078 ASIG5V.n9077 0.019716
R54973 ASIG5V.n9083 ASIG5V.n6461 0.019716
R54974 ASIG5V.n9083 ASIG5V.n9082 0.019716
R54975 ASIG5V.n9089 ASIG5V.n6460 0.019716
R54976 ASIG5V.n9090 ASIG5V.n9089 0.019716
R54977 ASIG5V.n9095 ASIG5V.n6459 0.019716
R54978 ASIG5V.n9095 ASIG5V.n9094 0.019716
R54979 ASIG5V.n9101 ASIG5V.n6458 0.019716
R54980 ASIG5V.n9102 ASIG5V.n9101 0.019716
R54981 ASIG5V.n9107 ASIG5V.n6457 0.019716
R54982 ASIG5V.n9107 ASIG5V.n9106 0.019716
R54983 ASIG5V.n9113 ASIG5V.n6456 0.019716
R54984 ASIG5V.n9114 ASIG5V.n9113 0.019716
R54985 ASIG5V.n9119 ASIG5V.n6455 0.019716
R54986 ASIG5V.n9119 ASIG5V.n9118 0.019716
R54987 ASIG5V.n9125 ASIG5V.n6454 0.019716
R54988 ASIG5V.n9126 ASIG5V.n9125 0.019716
R54989 ASIG5V.n9131 ASIG5V.n6453 0.019716
R54990 ASIG5V.n9131 ASIG5V.n9130 0.019716
R54991 ASIG5V.n9137 ASIG5V.n6452 0.019716
R54992 ASIG5V.n9138 ASIG5V.n9137 0.019716
R54993 ASIG5V.n9143 ASIG5V.n6451 0.019716
R54994 ASIG5V.n9143 ASIG5V.n9142 0.019716
R54995 ASIG5V.n9149 ASIG5V.n6450 0.019716
R54996 ASIG5V.n9150 ASIG5V.n9149 0.019716
R54997 ASIG5V.n9155 ASIG5V.n6449 0.019716
R54998 ASIG5V.n9155 ASIG5V.n9154 0.019716
R54999 ASIG5V.n9161 ASIG5V.n6448 0.019716
R55000 ASIG5V.n9162 ASIG5V.n9161 0.019716
R55001 ASIG5V.n9167 ASIG5V.n6447 0.019716
R55002 ASIG5V.n9167 ASIG5V.n9166 0.019716
R55003 ASIG5V.n9173 ASIG5V.n6446 0.019716
R55004 ASIG5V.n9174 ASIG5V.n9173 0.019716
R55005 ASIG5V.n8918 ASIG5V.n6588 0.019716
R55006 ASIG5V.n6694 ASIG5V.n6631 0.019716
R55007 ASIG5V.n6694 ASIG5V.n6586 0.019716
R55008 ASIG5V.n6703 ASIG5V.n6630 0.019716
R55009 ASIG5V.n6703 ASIG5V.n6585 0.019716
R55010 ASIG5V.n6691 ASIG5V.n6629 0.019716
R55011 ASIG5V.n6691 ASIG5V.n6584 0.019716
R55012 ASIG5V.n6712 ASIG5V.n6628 0.019716
R55013 ASIG5V.n6712 ASIG5V.n6583 0.019716
R55014 ASIG5V.n6688 ASIG5V.n6627 0.019716
R55015 ASIG5V.n6688 ASIG5V.n6582 0.019716
R55016 ASIG5V.n6721 ASIG5V.n6626 0.019716
R55017 ASIG5V.n6721 ASIG5V.n6581 0.019716
R55018 ASIG5V.n6685 ASIG5V.n6625 0.019716
R55019 ASIG5V.n6685 ASIG5V.n6580 0.019716
R55020 ASIG5V.n6730 ASIG5V.n6624 0.019716
R55021 ASIG5V.n6730 ASIG5V.n6579 0.019716
R55022 ASIG5V.n6682 ASIG5V.n6623 0.019716
R55023 ASIG5V.n6682 ASIG5V.n6578 0.019716
R55024 ASIG5V.n6739 ASIG5V.n6622 0.019716
R55025 ASIG5V.n6739 ASIG5V.n6577 0.019716
R55026 ASIG5V.n6679 ASIG5V.n6621 0.019716
R55027 ASIG5V.n6679 ASIG5V.n6576 0.019716
R55028 ASIG5V.n6748 ASIG5V.n6620 0.019716
R55029 ASIG5V.n6748 ASIG5V.n6575 0.019716
R55030 ASIG5V.n6676 ASIG5V.n6619 0.019716
R55031 ASIG5V.n6676 ASIG5V.n6574 0.019716
R55032 ASIG5V.n6757 ASIG5V.n6618 0.019716
R55033 ASIG5V.n6757 ASIG5V.n6573 0.019716
R55034 ASIG5V.n6673 ASIG5V.n6617 0.019716
R55035 ASIG5V.n6673 ASIG5V.n6572 0.019716
R55036 ASIG5V.n6766 ASIG5V.n6616 0.019716
R55037 ASIG5V.n6766 ASIG5V.n6571 0.019716
R55038 ASIG5V.n6670 ASIG5V.n6615 0.019716
R55039 ASIG5V.n6670 ASIG5V.n6570 0.019716
R55040 ASIG5V.n6775 ASIG5V.n6614 0.019716
R55041 ASIG5V.n6775 ASIG5V.n6569 0.019716
R55042 ASIG5V.n6667 ASIG5V.n6613 0.019716
R55043 ASIG5V.n6667 ASIG5V.n6568 0.019716
R55044 ASIG5V.n6784 ASIG5V.n6612 0.019716
R55045 ASIG5V.n6784 ASIG5V.n6567 0.019716
R55046 ASIG5V.n6664 ASIG5V.n6611 0.019716
R55047 ASIG5V.n6664 ASIG5V.n6566 0.019716
R55048 ASIG5V.n6793 ASIG5V.n6610 0.019716
R55049 ASIG5V.n6793 ASIG5V.n6565 0.019716
R55050 ASIG5V.n6661 ASIG5V.n6609 0.019716
R55051 ASIG5V.n6661 ASIG5V.n6564 0.019716
R55052 ASIG5V.n6802 ASIG5V.n6608 0.019716
R55053 ASIG5V.n6802 ASIG5V.n6563 0.019716
R55054 ASIG5V.n6658 ASIG5V.n6607 0.019716
R55055 ASIG5V.n6658 ASIG5V.n6562 0.019716
R55056 ASIG5V.n6811 ASIG5V.n6606 0.019716
R55057 ASIG5V.n6811 ASIG5V.n6561 0.019716
R55058 ASIG5V.n6655 ASIG5V.n6605 0.019716
R55059 ASIG5V.n6655 ASIG5V.n6560 0.019716
R55060 ASIG5V.n6820 ASIG5V.n6604 0.019716
R55061 ASIG5V.n6820 ASIG5V.n6559 0.019716
R55062 ASIG5V.n6652 ASIG5V.n6603 0.019716
R55063 ASIG5V.n6652 ASIG5V.n6558 0.019716
R55064 ASIG5V.n6829 ASIG5V.n6602 0.019716
R55065 ASIG5V.n6829 ASIG5V.n6557 0.019716
R55066 ASIG5V.n6649 ASIG5V.n6601 0.019716
R55067 ASIG5V.n6649 ASIG5V.n6556 0.019716
R55068 ASIG5V.n6838 ASIG5V.n6600 0.019716
R55069 ASIG5V.n6838 ASIG5V.n6555 0.019716
R55070 ASIG5V.n6646 ASIG5V.n6599 0.019716
R55071 ASIG5V.n6646 ASIG5V.n6554 0.019716
R55072 ASIG5V.n6847 ASIG5V.n6598 0.019716
R55073 ASIG5V.n6847 ASIG5V.n6553 0.019716
R55074 ASIG5V.n6643 ASIG5V.n6597 0.019716
R55075 ASIG5V.n6643 ASIG5V.n6552 0.019716
R55076 ASIG5V.n6856 ASIG5V.n6596 0.019716
R55077 ASIG5V.n6856 ASIG5V.n6551 0.019716
R55078 ASIG5V.n6640 ASIG5V.n6595 0.019716
R55079 ASIG5V.n6640 ASIG5V.n6550 0.019716
R55080 ASIG5V.n6865 ASIG5V.n6594 0.019716
R55081 ASIG5V.n6865 ASIG5V.n6549 0.019716
R55082 ASIG5V.n6637 ASIG5V.n6593 0.019716
R55083 ASIG5V.n6637 ASIG5V.n6548 0.019716
R55084 ASIG5V.n6874 ASIG5V.n6592 0.019716
R55085 ASIG5V.n6874 ASIG5V.n6547 0.019716
R55086 ASIG5V.n6634 ASIG5V.n6591 0.019716
R55087 ASIG5V.n6634 ASIG5V.n6546 0.019716
R55088 ASIG5V.n7228 ASIG5V.n7227 0.019716
R55089 ASIG5V.n7226 ASIG5V.n7225 0.019716
R55090 ASIG5V.n7225 ASIG5V.n6899 0.019716
R55091 ASIG5V.n7219 ASIG5V.n6904 0.019716
R55092 ASIG5V.n7219 ASIG5V.n7218 0.019716
R55093 ASIG5V.n7216 ASIG5V.n7215 0.019716
R55094 ASIG5V.n7215 ASIG5V.n6905 0.019716
R55095 ASIG5V.n7209 ASIG5V.n6910 0.019716
R55096 ASIG5V.n7209 ASIG5V.n7208 0.019716
R55097 ASIG5V.n7206 ASIG5V.n7205 0.019716
R55098 ASIG5V.n7205 ASIG5V.n6911 0.019716
R55099 ASIG5V.n7199 ASIG5V.n6916 0.019716
R55100 ASIG5V.n7199 ASIG5V.n7198 0.019716
R55101 ASIG5V.n7196 ASIG5V.n7195 0.019716
R55102 ASIG5V.n7195 ASIG5V.n6917 0.019716
R55103 ASIG5V.n7189 ASIG5V.n6922 0.019716
R55104 ASIG5V.n7189 ASIG5V.n7188 0.019716
R55105 ASIG5V.n7186 ASIG5V.n7185 0.019716
R55106 ASIG5V.n7185 ASIG5V.n6923 0.019716
R55107 ASIG5V.n7179 ASIG5V.n6928 0.019716
R55108 ASIG5V.n7179 ASIG5V.n7178 0.019716
R55109 ASIG5V.n7176 ASIG5V.n7175 0.019716
R55110 ASIG5V.n7175 ASIG5V.n6929 0.019716
R55111 ASIG5V.n7169 ASIG5V.n6934 0.019716
R55112 ASIG5V.n7169 ASIG5V.n7168 0.019716
R55113 ASIG5V.n7166 ASIG5V.n7165 0.019716
R55114 ASIG5V.n7165 ASIG5V.n6935 0.019716
R55115 ASIG5V.n7159 ASIG5V.n6940 0.019716
R55116 ASIG5V.n7159 ASIG5V.n7158 0.019716
R55117 ASIG5V.n7156 ASIG5V.n7155 0.019716
R55118 ASIG5V.n7155 ASIG5V.n6941 0.019716
R55119 ASIG5V.n7149 ASIG5V.n6946 0.019716
R55120 ASIG5V.n7149 ASIG5V.n7148 0.019716
R55121 ASIG5V.n7146 ASIG5V.n7145 0.019716
R55122 ASIG5V.n7145 ASIG5V.n6947 0.019716
R55123 ASIG5V.n7139 ASIG5V.n6952 0.019716
R55124 ASIG5V.n7139 ASIG5V.n7138 0.019716
R55125 ASIG5V.n7136 ASIG5V.n7135 0.019716
R55126 ASIG5V.n7135 ASIG5V.n6953 0.019716
R55127 ASIG5V.n7129 ASIG5V.n6958 0.019716
R55128 ASIG5V.n7129 ASIG5V.n7128 0.019716
R55129 ASIG5V.n7126 ASIG5V.n7125 0.019716
R55130 ASIG5V.n7125 ASIG5V.n6959 0.019716
R55131 ASIG5V.n7119 ASIG5V.n6964 0.019716
R55132 ASIG5V.n7119 ASIG5V.n7118 0.019716
R55133 ASIG5V.n7116 ASIG5V.n7115 0.019716
R55134 ASIG5V.n7115 ASIG5V.n6965 0.019716
R55135 ASIG5V.n7109 ASIG5V.n6970 0.019716
R55136 ASIG5V.n7109 ASIG5V.n7108 0.019716
R55137 ASIG5V.n7106 ASIG5V.n7105 0.019716
R55138 ASIG5V.n7105 ASIG5V.n6971 0.019716
R55139 ASIG5V.n7099 ASIG5V.n6976 0.019716
R55140 ASIG5V.n7099 ASIG5V.n7098 0.019716
R55141 ASIG5V.n7096 ASIG5V.n7095 0.019716
R55142 ASIG5V.n7095 ASIG5V.n6977 0.019716
R55143 ASIG5V.n7089 ASIG5V.n6982 0.019716
R55144 ASIG5V.n7089 ASIG5V.n7088 0.019716
R55145 ASIG5V.n7086 ASIG5V.n7085 0.019716
R55146 ASIG5V.n7085 ASIG5V.n6983 0.019716
R55147 ASIG5V.n7079 ASIG5V.n6988 0.019716
R55148 ASIG5V.n7079 ASIG5V.n7078 0.019716
R55149 ASIG5V.n7076 ASIG5V.n7075 0.019716
R55150 ASIG5V.n7075 ASIG5V.n6989 0.019716
R55151 ASIG5V.n7069 ASIG5V.n6994 0.019716
R55152 ASIG5V.n7069 ASIG5V.n7068 0.019716
R55153 ASIG5V.n7066 ASIG5V.n7065 0.019716
R55154 ASIG5V.n7065 ASIG5V.n6995 0.019716
R55155 ASIG5V.n7059 ASIG5V.n7000 0.019716
R55156 ASIG5V.n7059 ASIG5V.n7058 0.019716
R55157 ASIG5V.n7056 ASIG5V.n7055 0.019716
R55158 ASIG5V.n7055 ASIG5V.n7001 0.019716
R55159 ASIG5V.n7049 ASIG5V.n7006 0.019716
R55160 ASIG5V.n7049 ASIG5V.n7048 0.019716
R55161 ASIG5V.n7046 ASIG5V.n7045 0.019716
R55162 ASIG5V.n7045 ASIG5V.n7007 0.019716
R55163 ASIG5V.n7039 ASIG5V.n7012 0.019716
R55164 ASIG5V.n7039 ASIG5V.n7038 0.019716
R55165 ASIG5V.n7036 ASIG5V.n7035 0.019716
R55166 ASIG5V.n7035 ASIG5V.n7013 0.019716
R55167 ASIG5V.n7029 ASIG5V.n7018 0.019716
R55168 ASIG5V.n7029 ASIG5V.n7028 0.019716
R55169 ASIG5V.n7026 ASIG5V.n7025 0.019716
R55170 ASIG5V.n7025 ASIG5V.n7019 0.019716
R55171 ASIG5V.n8894 ASIG5V.n8214 0.019716
R55172 ASIG5V.n8564 ASIG5V.n8258 0.019716
R55173 ASIG5V.n8564 ASIG5V.n8212 0.019716
R55174 ASIG5V.n8326 ASIG5V.n8257 0.019716
R55175 ASIG5V.n8326 ASIG5V.n8211 0.019716
R55176 ASIG5V.n8555 ASIG5V.n8256 0.019716
R55177 ASIG5V.n8555 ASIG5V.n8210 0.019716
R55178 ASIG5V.n8329 ASIG5V.n8255 0.019716
R55179 ASIG5V.n8329 ASIG5V.n8209 0.019716
R55180 ASIG5V.n8546 ASIG5V.n8254 0.019716
R55181 ASIG5V.n8546 ASIG5V.n8208 0.019716
R55182 ASIG5V.n8332 ASIG5V.n8253 0.019716
R55183 ASIG5V.n8332 ASIG5V.n8207 0.019716
R55184 ASIG5V.n8537 ASIG5V.n8252 0.019716
R55185 ASIG5V.n8537 ASIG5V.n8206 0.019716
R55186 ASIG5V.n8335 ASIG5V.n8251 0.019716
R55187 ASIG5V.n8335 ASIG5V.n8205 0.019716
R55188 ASIG5V.n8528 ASIG5V.n8250 0.019716
R55189 ASIG5V.n8528 ASIG5V.n8204 0.019716
R55190 ASIG5V.n8338 ASIG5V.n8249 0.019716
R55191 ASIG5V.n8338 ASIG5V.n8203 0.019716
R55192 ASIG5V.n8519 ASIG5V.n8248 0.019716
R55193 ASIG5V.n8519 ASIG5V.n8202 0.019716
R55194 ASIG5V.n8341 ASIG5V.n8247 0.019716
R55195 ASIG5V.n8341 ASIG5V.n8201 0.019716
R55196 ASIG5V.n8510 ASIG5V.n8246 0.019716
R55197 ASIG5V.n8510 ASIG5V.n8200 0.019716
R55198 ASIG5V.n8344 ASIG5V.n8245 0.019716
R55199 ASIG5V.n8344 ASIG5V.n8199 0.019716
R55200 ASIG5V.n8501 ASIG5V.n8244 0.019716
R55201 ASIG5V.n8501 ASIG5V.n8198 0.019716
R55202 ASIG5V.n8347 ASIG5V.n8243 0.019716
R55203 ASIG5V.n8347 ASIG5V.n8197 0.019716
R55204 ASIG5V.n8492 ASIG5V.n8242 0.019716
R55205 ASIG5V.n8492 ASIG5V.n8196 0.019716
R55206 ASIG5V.n8350 ASIG5V.n8241 0.019716
R55207 ASIG5V.n8350 ASIG5V.n8195 0.019716
R55208 ASIG5V.n8483 ASIG5V.n8240 0.019716
R55209 ASIG5V.n8483 ASIG5V.n8194 0.019716
R55210 ASIG5V.n8353 ASIG5V.n8239 0.019716
R55211 ASIG5V.n8353 ASIG5V.n8193 0.019716
R55212 ASIG5V.n8474 ASIG5V.n8238 0.019716
R55213 ASIG5V.n8474 ASIG5V.n8192 0.019716
R55214 ASIG5V.n8356 ASIG5V.n8237 0.019716
R55215 ASIG5V.n8356 ASIG5V.n8191 0.019716
R55216 ASIG5V.n8465 ASIG5V.n8236 0.019716
R55217 ASIG5V.n8465 ASIG5V.n8190 0.019716
R55218 ASIG5V.n8359 ASIG5V.n8235 0.019716
R55219 ASIG5V.n8359 ASIG5V.n8189 0.019716
R55220 ASIG5V.n8456 ASIG5V.n8234 0.019716
R55221 ASIG5V.n8456 ASIG5V.n8188 0.019716
R55222 ASIG5V.n8362 ASIG5V.n8233 0.019716
R55223 ASIG5V.n8362 ASIG5V.n8187 0.019716
R55224 ASIG5V.n8447 ASIG5V.n8232 0.019716
R55225 ASIG5V.n8447 ASIG5V.n8186 0.019716
R55226 ASIG5V.n8365 ASIG5V.n8231 0.019716
R55227 ASIG5V.n8365 ASIG5V.n8185 0.019716
R55228 ASIG5V.n8438 ASIG5V.n8230 0.019716
R55229 ASIG5V.n8438 ASIG5V.n8184 0.019716
R55230 ASIG5V.n8368 ASIG5V.n8229 0.019716
R55231 ASIG5V.n8368 ASIG5V.n8183 0.019716
R55232 ASIG5V.n8429 ASIG5V.n8228 0.019716
R55233 ASIG5V.n8429 ASIG5V.n8182 0.019716
R55234 ASIG5V.n8371 ASIG5V.n8227 0.019716
R55235 ASIG5V.n8371 ASIG5V.n8181 0.019716
R55236 ASIG5V.n8420 ASIG5V.n8226 0.019716
R55237 ASIG5V.n8420 ASIG5V.n8180 0.019716
R55238 ASIG5V.n8374 ASIG5V.n8225 0.019716
R55239 ASIG5V.n8374 ASIG5V.n8179 0.019716
R55240 ASIG5V.n8411 ASIG5V.n8224 0.019716
R55241 ASIG5V.n8411 ASIG5V.n8178 0.019716
R55242 ASIG5V.n8377 ASIG5V.n8223 0.019716
R55243 ASIG5V.n8377 ASIG5V.n8177 0.019716
R55244 ASIG5V.n8402 ASIG5V.n8222 0.019716
R55245 ASIG5V.n8402 ASIG5V.n8176 0.019716
R55246 ASIG5V.n8380 ASIG5V.n8221 0.019716
R55247 ASIG5V.n8380 ASIG5V.n8175 0.019716
R55248 ASIG5V.n8393 ASIG5V.n8220 0.019716
R55249 ASIG5V.n8393 ASIG5V.n8174 0.019716
R55250 ASIG5V.n8383 ASIG5V.n8219 0.019716
R55251 ASIG5V.n8383 ASIG5V.n8173 0.019716
R55252 ASIG5V.n8261 ASIG5V.n8218 0.019716
R55253 ASIG5V.n8261 ASIG5V.n8172 0.019716
R55254 ASIG5V.n8880 ASIG5V.n8319 0.019716
R55255 ASIG5V.n8590 ASIG5V.n8589 0.019716
R55256 ASIG5V.n8590 ASIG5V.n8318 0.019716
R55257 ASIG5V.n8871 ASIG5V.n8870 0.019716
R55258 ASIG5V.n8870 ASIG5V.n8317 0.019716
R55259 ASIG5V.n8866 ASIG5V.n8865 0.019716
R55260 ASIG5V.n8865 ASIG5V.n8316 0.019716
R55261 ASIG5V.n8859 ASIG5V.n8858 0.019716
R55262 ASIG5V.n8858 ASIG5V.n8315 0.019716
R55263 ASIG5V.n8854 ASIG5V.n8853 0.019716
R55264 ASIG5V.n8853 ASIG5V.n8314 0.019716
R55265 ASIG5V.n8847 ASIG5V.n8846 0.019716
R55266 ASIG5V.n8846 ASIG5V.n8313 0.019716
R55267 ASIG5V.n8842 ASIG5V.n8841 0.019716
R55268 ASIG5V.n8841 ASIG5V.n8312 0.019716
R55269 ASIG5V.n8835 ASIG5V.n8834 0.019716
R55270 ASIG5V.n8834 ASIG5V.n8311 0.019716
R55271 ASIG5V.n8830 ASIG5V.n8829 0.019716
R55272 ASIG5V.n8829 ASIG5V.n8310 0.019716
R55273 ASIG5V.n8823 ASIG5V.n8822 0.019716
R55274 ASIG5V.n8822 ASIG5V.n8309 0.019716
R55275 ASIG5V.n8818 ASIG5V.n8817 0.019716
R55276 ASIG5V.n8817 ASIG5V.n8308 0.019716
R55277 ASIG5V.n8811 ASIG5V.n8810 0.019716
R55278 ASIG5V.n8810 ASIG5V.n8307 0.019716
R55279 ASIG5V.n8806 ASIG5V.n8805 0.019716
R55280 ASIG5V.n8805 ASIG5V.n8306 0.019716
R55281 ASIG5V.n8799 ASIG5V.n8798 0.019716
R55282 ASIG5V.n8798 ASIG5V.n8305 0.019716
R55283 ASIG5V.n8794 ASIG5V.n8793 0.019716
R55284 ASIG5V.n8793 ASIG5V.n8304 0.019716
R55285 ASIG5V.n8787 ASIG5V.n8786 0.019716
R55286 ASIG5V.n8786 ASIG5V.n8303 0.019716
R55287 ASIG5V.n8782 ASIG5V.n8781 0.019716
R55288 ASIG5V.n8781 ASIG5V.n8302 0.019716
R55289 ASIG5V.n8775 ASIG5V.n8774 0.019716
R55290 ASIG5V.n8774 ASIG5V.n8301 0.019716
R55291 ASIG5V.n8770 ASIG5V.n8769 0.019716
R55292 ASIG5V.n8769 ASIG5V.n8300 0.019716
R55293 ASIG5V.n8763 ASIG5V.n8762 0.019716
R55294 ASIG5V.n8762 ASIG5V.n8299 0.019716
R55295 ASIG5V.n8758 ASIG5V.n8757 0.019716
R55296 ASIG5V.n8757 ASIG5V.n8298 0.019716
R55297 ASIG5V.n8751 ASIG5V.n8750 0.019716
R55298 ASIG5V.n8750 ASIG5V.n8297 0.019716
R55299 ASIG5V.n8746 ASIG5V.n8745 0.019716
R55300 ASIG5V.n8745 ASIG5V.n8296 0.019716
R55301 ASIG5V.n8739 ASIG5V.n8738 0.019716
R55302 ASIG5V.n8738 ASIG5V.n8295 0.019716
R55303 ASIG5V.n8734 ASIG5V.n8733 0.019716
R55304 ASIG5V.n8733 ASIG5V.n8294 0.019716
R55305 ASIG5V.n8727 ASIG5V.n8726 0.019716
R55306 ASIG5V.n8726 ASIG5V.n8293 0.019716
R55307 ASIG5V.n8722 ASIG5V.n8721 0.019716
R55308 ASIG5V.n8721 ASIG5V.n8292 0.019716
R55309 ASIG5V.n8715 ASIG5V.n8714 0.019716
R55310 ASIG5V.n8714 ASIG5V.n8291 0.019716
R55311 ASIG5V.n8710 ASIG5V.n8709 0.019716
R55312 ASIG5V.n8709 ASIG5V.n8290 0.019716
R55313 ASIG5V.n8703 ASIG5V.n8702 0.019716
R55314 ASIG5V.n8702 ASIG5V.n8289 0.019716
R55315 ASIG5V.n8698 ASIG5V.n8697 0.019716
R55316 ASIG5V.n8697 ASIG5V.n8288 0.019716
R55317 ASIG5V.n8691 ASIG5V.n8690 0.019716
R55318 ASIG5V.n8690 ASIG5V.n8287 0.019716
R55319 ASIG5V.n8686 ASIG5V.n8685 0.019716
R55320 ASIG5V.n8685 ASIG5V.n8286 0.019716
R55321 ASIG5V.n8679 ASIG5V.n8678 0.019716
R55322 ASIG5V.n8678 ASIG5V.n8285 0.019716
R55323 ASIG5V.n8674 ASIG5V.n8673 0.019716
R55324 ASIG5V.n8673 ASIG5V.n8284 0.019716
R55325 ASIG5V.n8667 ASIG5V.n8666 0.019716
R55326 ASIG5V.n8666 ASIG5V.n8283 0.019716
R55327 ASIG5V.n8662 ASIG5V.n8661 0.019716
R55328 ASIG5V.n8661 ASIG5V.n8282 0.019716
R55329 ASIG5V.n8655 ASIG5V.n8654 0.019716
R55330 ASIG5V.n8654 ASIG5V.n8281 0.019716
R55331 ASIG5V.n8650 ASIG5V.n8649 0.019716
R55332 ASIG5V.n8649 ASIG5V.n8280 0.019716
R55333 ASIG5V.n8643 ASIG5V.n8642 0.019716
R55334 ASIG5V.n8642 ASIG5V.n8279 0.019716
R55335 ASIG5V.n8638 ASIG5V.n8637 0.019716
R55336 ASIG5V.n8637 ASIG5V.n8278 0.019716
R55337 ASIG5V.n12527 ASIG5V.n53 0.019716
R55338 ASIG5V.n159 ASIG5V.n97 0.019716
R55339 ASIG5V.n159 ASIG5V.n51 0.019716
R55340 ASIG5V.n12345 ASIG5V.n96 0.019716
R55341 ASIG5V.n12345 ASIG5V.n50 0.019716
R55342 ASIG5V.n156 ASIG5V.n95 0.019716
R55343 ASIG5V.n156 ASIG5V.n49 0.019716
R55344 ASIG5V.n12354 ASIG5V.n94 0.019716
R55345 ASIG5V.n12354 ASIG5V.n48 0.019716
R55346 ASIG5V.n153 ASIG5V.n93 0.019716
R55347 ASIG5V.n153 ASIG5V.n47 0.019716
R55348 ASIG5V.n12363 ASIG5V.n92 0.019716
R55349 ASIG5V.n12363 ASIG5V.n46 0.019716
R55350 ASIG5V.n150 ASIG5V.n91 0.019716
R55351 ASIG5V.n150 ASIG5V.n45 0.019716
R55352 ASIG5V.n12372 ASIG5V.n90 0.019716
R55353 ASIG5V.n12372 ASIG5V.n44 0.019716
R55354 ASIG5V.n147 ASIG5V.n89 0.019716
R55355 ASIG5V.n147 ASIG5V.n43 0.019716
R55356 ASIG5V.n12381 ASIG5V.n88 0.019716
R55357 ASIG5V.n12381 ASIG5V.n42 0.019716
R55358 ASIG5V.n144 ASIG5V.n87 0.019716
R55359 ASIG5V.n144 ASIG5V.n41 0.019716
R55360 ASIG5V.n12390 ASIG5V.n86 0.019716
R55361 ASIG5V.n12390 ASIG5V.n40 0.019716
R55362 ASIG5V.n141 ASIG5V.n85 0.019716
R55363 ASIG5V.n141 ASIG5V.n39 0.019716
R55364 ASIG5V.n12399 ASIG5V.n84 0.019716
R55365 ASIG5V.n12399 ASIG5V.n38 0.019716
R55366 ASIG5V.n138 ASIG5V.n83 0.019716
R55367 ASIG5V.n138 ASIG5V.n37 0.019716
R55368 ASIG5V.n12408 ASIG5V.n82 0.019716
R55369 ASIG5V.n12408 ASIG5V.n36 0.019716
R55370 ASIG5V.n135 ASIG5V.n81 0.019716
R55371 ASIG5V.n135 ASIG5V.n35 0.019716
R55372 ASIG5V.n12417 ASIG5V.n80 0.019716
R55373 ASIG5V.n12417 ASIG5V.n34 0.019716
R55374 ASIG5V.n132 ASIG5V.n79 0.019716
R55375 ASIG5V.n132 ASIG5V.n33 0.019716
R55376 ASIG5V.n12426 ASIG5V.n78 0.019716
R55377 ASIG5V.n12426 ASIG5V.n32 0.019716
R55378 ASIG5V.n129 ASIG5V.n77 0.019716
R55379 ASIG5V.n129 ASIG5V.n31 0.019716
R55380 ASIG5V.n12435 ASIG5V.n76 0.019716
R55381 ASIG5V.n12435 ASIG5V.n30 0.019716
R55382 ASIG5V.n126 ASIG5V.n75 0.019716
R55383 ASIG5V.n126 ASIG5V.n29 0.019716
R55384 ASIG5V.n12444 ASIG5V.n74 0.019716
R55385 ASIG5V.n12444 ASIG5V.n28 0.019716
R55386 ASIG5V.n123 ASIG5V.n73 0.019716
R55387 ASIG5V.n123 ASIG5V.n27 0.019716
R55388 ASIG5V.n12453 ASIG5V.n72 0.019716
R55389 ASIG5V.n12453 ASIG5V.n26 0.019716
R55390 ASIG5V.n120 ASIG5V.n71 0.019716
R55391 ASIG5V.n120 ASIG5V.n25 0.019716
R55392 ASIG5V.n12462 ASIG5V.n70 0.019716
R55393 ASIG5V.n12462 ASIG5V.n24 0.019716
R55394 ASIG5V.n117 ASIG5V.n69 0.019716
R55395 ASIG5V.n117 ASIG5V.n23 0.019716
R55396 ASIG5V.n12471 ASIG5V.n68 0.019716
R55397 ASIG5V.n12471 ASIG5V.n22 0.019716
R55398 ASIG5V.n114 ASIG5V.n67 0.019716
R55399 ASIG5V.n114 ASIG5V.n21 0.019716
R55400 ASIG5V.n12480 ASIG5V.n66 0.019716
R55401 ASIG5V.n12480 ASIG5V.n20 0.019716
R55402 ASIG5V.n111 ASIG5V.n65 0.019716
R55403 ASIG5V.n111 ASIG5V.n19 0.019716
R55404 ASIG5V.n12489 ASIG5V.n64 0.019716
R55405 ASIG5V.n12489 ASIG5V.n18 0.019716
R55406 ASIG5V.n108 ASIG5V.n63 0.019716
R55407 ASIG5V.n108 ASIG5V.n17 0.019716
R55408 ASIG5V.n12498 ASIG5V.n62 0.019716
R55409 ASIG5V.n12498 ASIG5V.n16 0.019716
R55410 ASIG5V.n105 ASIG5V.n61 0.019716
R55411 ASIG5V.n105 ASIG5V.n15 0.019716
R55412 ASIG5V.n12507 ASIG5V.n60 0.019716
R55413 ASIG5V.n12507 ASIG5V.n14 0.019716
R55414 ASIG5V.n102 ASIG5V.n59 0.019716
R55415 ASIG5V.n102 ASIG5V.n13 0.019716
R55416 ASIG5V.n12516 ASIG5V.n58 0.019716
R55417 ASIG5V.n12516 ASIG5V.n12 0.019716
R55418 ASIG5V.n99 ASIG5V.n57 0.019716
R55419 ASIG5V.n99 ASIG5V.n11 0.019716
R55420 ASIG5V.n262 ASIG5V.n261 0.019716
R55421 ASIG5V.n267 ASIG5V.n214 0.019716
R55422 ASIG5V.n268 ASIG5V.n267 0.019716
R55423 ASIG5V.n273 ASIG5V.n213 0.019716
R55424 ASIG5V.n273 ASIG5V.n272 0.019716
R55425 ASIG5V.n279 ASIG5V.n212 0.019716
R55426 ASIG5V.n280 ASIG5V.n279 0.019716
R55427 ASIG5V.n285 ASIG5V.n211 0.019716
R55428 ASIG5V.n285 ASIG5V.n284 0.019716
R55429 ASIG5V.n291 ASIG5V.n210 0.019716
R55430 ASIG5V.n292 ASIG5V.n291 0.019716
R55431 ASIG5V.n297 ASIG5V.n209 0.019716
R55432 ASIG5V.n297 ASIG5V.n296 0.019716
R55433 ASIG5V.n303 ASIG5V.n208 0.019716
R55434 ASIG5V.n304 ASIG5V.n303 0.019716
R55435 ASIG5V.n309 ASIG5V.n207 0.019716
R55436 ASIG5V.n309 ASIG5V.n308 0.019716
R55437 ASIG5V.n315 ASIG5V.n206 0.019716
R55438 ASIG5V.n316 ASIG5V.n315 0.019716
R55439 ASIG5V.n321 ASIG5V.n205 0.019716
R55440 ASIG5V.n321 ASIG5V.n320 0.019716
R55441 ASIG5V.n327 ASIG5V.n204 0.019716
R55442 ASIG5V.n328 ASIG5V.n327 0.019716
R55443 ASIG5V.n333 ASIG5V.n203 0.019716
R55444 ASIG5V.n333 ASIG5V.n332 0.019716
R55445 ASIG5V.n339 ASIG5V.n202 0.019716
R55446 ASIG5V.n340 ASIG5V.n339 0.019716
R55447 ASIG5V.n345 ASIG5V.n201 0.019716
R55448 ASIG5V.n345 ASIG5V.n344 0.019716
R55449 ASIG5V.n351 ASIG5V.n200 0.019716
R55450 ASIG5V.n352 ASIG5V.n351 0.019716
R55451 ASIG5V.n357 ASIG5V.n199 0.019716
R55452 ASIG5V.n357 ASIG5V.n356 0.019716
R55453 ASIG5V.n363 ASIG5V.n198 0.019716
R55454 ASIG5V.n364 ASIG5V.n363 0.019716
R55455 ASIG5V.n369 ASIG5V.n197 0.019716
R55456 ASIG5V.n369 ASIG5V.n368 0.019716
R55457 ASIG5V.n375 ASIG5V.n196 0.019716
R55458 ASIG5V.n376 ASIG5V.n375 0.019716
R55459 ASIG5V.n381 ASIG5V.n195 0.019716
R55460 ASIG5V.n381 ASIG5V.n380 0.019716
R55461 ASIG5V.n387 ASIG5V.n194 0.019716
R55462 ASIG5V.n388 ASIG5V.n387 0.019716
R55463 ASIG5V.n393 ASIG5V.n193 0.019716
R55464 ASIG5V.n393 ASIG5V.n392 0.019716
R55465 ASIG5V.n399 ASIG5V.n192 0.019716
R55466 ASIG5V.n400 ASIG5V.n399 0.019716
R55467 ASIG5V.n405 ASIG5V.n191 0.019716
R55468 ASIG5V.n405 ASIG5V.n404 0.019716
R55469 ASIG5V.n411 ASIG5V.n190 0.019716
R55470 ASIG5V.n412 ASIG5V.n411 0.019716
R55471 ASIG5V.n417 ASIG5V.n189 0.019716
R55472 ASIG5V.n417 ASIG5V.n416 0.019716
R55473 ASIG5V.n423 ASIG5V.n188 0.019716
R55474 ASIG5V.n424 ASIG5V.n423 0.019716
R55475 ASIG5V.n429 ASIG5V.n187 0.019716
R55476 ASIG5V.n429 ASIG5V.n428 0.019716
R55477 ASIG5V.n435 ASIG5V.n186 0.019716
R55478 ASIG5V.n436 ASIG5V.n435 0.019716
R55479 ASIG5V.n441 ASIG5V.n185 0.019716
R55480 ASIG5V.n441 ASIG5V.n440 0.019716
R55481 ASIG5V.n447 ASIG5V.n184 0.019716
R55482 ASIG5V.n448 ASIG5V.n447 0.019716
R55483 ASIG5V.n453 ASIG5V.n183 0.019716
R55484 ASIG5V.n453 ASIG5V.n452 0.019716
R55485 ASIG5V.n459 ASIG5V.n182 0.019716
R55486 ASIG5V.n460 ASIG5V.n459 0.019716
R55487 ASIG5V.n465 ASIG5V.n181 0.019716
R55488 ASIG5V.n465 ASIG5V.n464 0.019716
R55489 ASIG5V.n471 ASIG5V.n180 0.019716
R55490 ASIG5V.n472 ASIG5V.n471 0.019716
R55491 ASIG5V.n477 ASIG5V.n179 0.019716
R55492 ASIG5V.n477 ASIG5V.n476 0.019716
R55493 ASIG5V.n483 ASIG5V.n178 0.019716
R55494 ASIG5V.n484 ASIG5V.n483 0.019716
R55495 ASIG5V.n489 ASIG5V.n177 0.019716
R55496 ASIG5V.n489 ASIG5V.n488 0.019716
R55497 ASIG5V.n495 ASIG5V.n176 0.019716
R55498 ASIG5V.n496 ASIG5V.n495 0.019716
R55499 ASIG5V.n501 ASIG5V.n175 0.019716
R55500 ASIG5V.n501 ASIG5V.n500 0.019716
R55501 ASIG5V.n12320 ASIG5V.n174 0.019716
R55502 ASIG5V.n12321 ASIG5V.n12320 0.019716
R55503 ASIG5V.n616 ASIG5V.n615 0.019716
R55504 ASIG5V.n621 ASIG5V.n569 0.019716
R55505 ASIG5V.n622 ASIG5V.n621 0.019716
R55506 ASIG5V.n627 ASIG5V.n568 0.019716
R55507 ASIG5V.n627 ASIG5V.n626 0.019716
R55508 ASIG5V.n633 ASIG5V.n567 0.019716
R55509 ASIG5V.n634 ASIG5V.n633 0.019716
R55510 ASIG5V.n639 ASIG5V.n566 0.019716
R55511 ASIG5V.n639 ASIG5V.n638 0.019716
R55512 ASIG5V.n645 ASIG5V.n565 0.019716
R55513 ASIG5V.n646 ASIG5V.n645 0.019716
R55514 ASIG5V.n651 ASIG5V.n564 0.019716
R55515 ASIG5V.n651 ASIG5V.n650 0.019716
R55516 ASIG5V.n657 ASIG5V.n563 0.019716
R55517 ASIG5V.n658 ASIG5V.n657 0.019716
R55518 ASIG5V.n663 ASIG5V.n562 0.019716
R55519 ASIG5V.n663 ASIG5V.n662 0.019716
R55520 ASIG5V.n669 ASIG5V.n561 0.019716
R55521 ASIG5V.n670 ASIG5V.n669 0.019716
R55522 ASIG5V.n675 ASIG5V.n560 0.019716
R55523 ASIG5V.n675 ASIG5V.n674 0.019716
R55524 ASIG5V.n681 ASIG5V.n559 0.019716
R55525 ASIG5V.n682 ASIG5V.n681 0.019716
R55526 ASIG5V.n687 ASIG5V.n558 0.019716
R55527 ASIG5V.n687 ASIG5V.n686 0.019716
R55528 ASIG5V.n693 ASIG5V.n557 0.019716
R55529 ASIG5V.n694 ASIG5V.n693 0.019716
R55530 ASIG5V.n699 ASIG5V.n556 0.019716
R55531 ASIG5V.n699 ASIG5V.n698 0.019716
R55532 ASIG5V.n705 ASIG5V.n555 0.019716
R55533 ASIG5V.n706 ASIG5V.n705 0.019716
R55534 ASIG5V.n711 ASIG5V.n554 0.019716
R55535 ASIG5V.n711 ASIG5V.n710 0.019716
R55536 ASIG5V.n717 ASIG5V.n553 0.019716
R55537 ASIG5V.n718 ASIG5V.n717 0.019716
R55538 ASIG5V.n723 ASIG5V.n552 0.019716
R55539 ASIG5V.n723 ASIG5V.n722 0.019716
R55540 ASIG5V.n729 ASIG5V.n551 0.019716
R55541 ASIG5V.n730 ASIG5V.n729 0.019716
R55542 ASIG5V.n735 ASIG5V.n550 0.019716
R55543 ASIG5V.n735 ASIG5V.n734 0.019716
R55544 ASIG5V.n741 ASIG5V.n549 0.019716
R55545 ASIG5V.n742 ASIG5V.n741 0.019716
R55546 ASIG5V.n747 ASIG5V.n548 0.019716
R55547 ASIG5V.n747 ASIG5V.n746 0.019716
R55548 ASIG5V.n753 ASIG5V.n547 0.019716
R55549 ASIG5V.n754 ASIG5V.n753 0.019716
R55550 ASIG5V.n759 ASIG5V.n546 0.019716
R55551 ASIG5V.n759 ASIG5V.n758 0.019716
R55552 ASIG5V.n765 ASIG5V.n545 0.019716
R55553 ASIG5V.n766 ASIG5V.n765 0.019716
R55554 ASIG5V.n771 ASIG5V.n544 0.019716
R55555 ASIG5V.n771 ASIG5V.n770 0.019716
R55556 ASIG5V.n777 ASIG5V.n543 0.019716
R55557 ASIG5V.n778 ASIG5V.n777 0.019716
R55558 ASIG5V.n783 ASIG5V.n542 0.019716
R55559 ASIG5V.n783 ASIG5V.n782 0.019716
R55560 ASIG5V.n789 ASIG5V.n541 0.019716
R55561 ASIG5V.n790 ASIG5V.n789 0.019716
R55562 ASIG5V.n795 ASIG5V.n540 0.019716
R55563 ASIG5V.n795 ASIG5V.n794 0.019716
R55564 ASIG5V.n801 ASIG5V.n539 0.019716
R55565 ASIG5V.n802 ASIG5V.n801 0.019716
R55566 ASIG5V.n807 ASIG5V.n538 0.019716
R55567 ASIG5V.n807 ASIG5V.n806 0.019716
R55568 ASIG5V.n813 ASIG5V.n537 0.019716
R55569 ASIG5V.n814 ASIG5V.n813 0.019716
R55570 ASIG5V.n819 ASIG5V.n536 0.019716
R55571 ASIG5V.n819 ASIG5V.n818 0.019716
R55572 ASIG5V.n825 ASIG5V.n535 0.019716
R55573 ASIG5V.n826 ASIG5V.n825 0.019716
R55574 ASIG5V.n831 ASIG5V.n534 0.019716
R55575 ASIG5V.n831 ASIG5V.n830 0.019716
R55576 ASIG5V.n837 ASIG5V.n533 0.019716
R55577 ASIG5V.n838 ASIG5V.n837 0.019716
R55578 ASIG5V.n843 ASIG5V.n532 0.019716
R55579 ASIG5V.n843 ASIG5V.n842 0.019716
R55580 ASIG5V.n849 ASIG5V.n531 0.019716
R55581 ASIG5V.n850 ASIG5V.n849 0.019716
R55582 ASIG5V.n855 ASIG5V.n530 0.019716
R55583 ASIG5V.n855 ASIG5V.n854 0.019716
R55584 ASIG5V.n12298 ASIG5V.n529 0.019716
R55585 ASIG5V.n12299 ASIG5V.n12298 0.019716
R55586 ASIG5V.n969 ASIG5V.n968 0.019716
R55587 ASIG5V.n973 ASIG5V.n970 0.019716
R55588 ASIG5V.n973 ASIG5V.n972 0.019716
R55589 ASIG5V.n979 ASIG5V.n962 0.019716
R55590 ASIG5V.n980 ASIG5V.n979 0.019716
R55591 ASIG5V.n985 ASIG5V.n982 0.019716
R55592 ASIG5V.n985 ASIG5V.n984 0.019716
R55593 ASIG5V.n991 ASIG5V.n958 0.019716
R55594 ASIG5V.n992 ASIG5V.n991 0.019716
R55595 ASIG5V.n997 ASIG5V.n994 0.019716
R55596 ASIG5V.n997 ASIG5V.n996 0.019716
R55597 ASIG5V.n1003 ASIG5V.n954 0.019716
R55598 ASIG5V.n1004 ASIG5V.n1003 0.019716
R55599 ASIG5V.n1009 ASIG5V.n1006 0.019716
R55600 ASIG5V.n1009 ASIG5V.n1008 0.019716
R55601 ASIG5V.n1015 ASIG5V.n950 0.019716
R55602 ASIG5V.n1016 ASIG5V.n1015 0.019716
R55603 ASIG5V.n1021 ASIG5V.n1018 0.019716
R55604 ASIG5V.n1021 ASIG5V.n1020 0.019716
R55605 ASIG5V.n1027 ASIG5V.n946 0.019716
R55606 ASIG5V.n1028 ASIG5V.n1027 0.019716
R55607 ASIG5V.n1033 ASIG5V.n1030 0.019716
R55608 ASIG5V.n1033 ASIG5V.n1032 0.019716
R55609 ASIG5V.n1039 ASIG5V.n942 0.019716
R55610 ASIG5V.n1040 ASIG5V.n1039 0.019716
R55611 ASIG5V.n1045 ASIG5V.n1042 0.019716
R55612 ASIG5V.n1045 ASIG5V.n1044 0.019716
R55613 ASIG5V.n1051 ASIG5V.n938 0.019716
R55614 ASIG5V.n1052 ASIG5V.n1051 0.019716
R55615 ASIG5V.n1057 ASIG5V.n1054 0.019716
R55616 ASIG5V.n1057 ASIG5V.n1056 0.019716
R55617 ASIG5V.n1063 ASIG5V.n934 0.019716
R55618 ASIG5V.n1064 ASIG5V.n1063 0.019716
R55619 ASIG5V.n1069 ASIG5V.n1066 0.019716
R55620 ASIG5V.n1069 ASIG5V.n1068 0.019716
R55621 ASIG5V.n1075 ASIG5V.n930 0.019716
R55622 ASIG5V.n1076 ASIG5V.n1075 0.019716
R55623 ASIG5V.n1081 ASIG5V.n1078 0.019716
R55624 ASIG5V.n1081 ASIG5V.n1080 0.019716
R55625 ASIG5V.n1087 ASIG5V.n926 0.019716
R55626 ASIG5V.n1088 ASIG5V.n1087 0.019716
R55627 ASIG5V.n1093 ASIG5V.n1090 0.019716
R55628 ASIG5V.n1093 ASIG5V.n1092 0.019716
R55629 ASIG5V.n1099 ASIG5V.n922 0.019716
R55630 ASIG5V.n1100 ASIG5V.n1099 0.019716
R55631 ASIG5V.n1105 ASIG5V.n1102 0.019716
R55632 ASIG5V.n1105 ASIG5V.n1104 0.019716
R55633 ASIG5V.n1111 ASIG5V.n918 0.019716
R55634 ASIG5V.n1112 ASIG5V.n1111 0.019716
R55635 ASIG5V.n1117 ASIG5V.n1114 0.019716
R55636 ASIG5V.n1117 ASIG5V.n1116 0.019716
R55637 ASIG5V.n1123 ASIG5V.n914 0.019716
R55638 ASIG5V.n1124 ASIG5V.n1123 0.019716
R55639 ASIG5V.n1129 ASIG5V.n1126 0.019716
R55640 ASIG5V.n1129 ASIG5V.n1128 0.019716
R55641 ASIG5V.n1135 ASIG5V.n910 0.019716
R55642 ASIG5V.n1136 ASIG5V.n1135 0.019716
R55643 ASIG5V.n1141 ASIG5V.n1138 0.019716
R55644 ASIG5V.n1141 ASIG5V.n1140 0.019716
R55645 ASIG5V.n1147 ASIG5V.n906 0.019716
R55646 ASIG5V.n1148 ASIG5V.n1147 0.019716
R55647 ASIG5V.n1153 ASIG5V.n1150 0.019716
R55648 ASIG5V.n1153 ASIG5V.n1152 0.019716
R55649 ASIG5V.n1159 ASIG5V.n902 0.019716
R55650 ASIG5V.n1160 ASIG5V.n1159 0.019716
R55651 ASIG5V.n1165 ASIG5V.n1162 0.019716
R55652 ASIG5V.n1165 ASIG5V.n1164 0.019716
R55653 ASIG5V.n1171 ASIG5V.n898 0.019716
R55654 ASIG5V.n1172 ASIG5V.n1171 0.019716
R55655 ASIG5V.n1177 ASIG5V.n1174 0.019716
R55656 ASIG5V.n1177 ASIG5V.n1176 0.019716
R55657 ASIG5V.n1183 ASIG5V.n894 0.019716
R55658 ASIG5V.n1184 ASIG5V.n1183 0.019716
R55659 ASIG5V.n1189 ASIG5V.n1186 0.019716
R55660 ASIG5V.n1189 ASIG5V.n1188 0.019716
R55661 ASIG5V.n1195 ASIG5V.n890 0.019716
R55662 ASIG5V.n1196 ASIG5V.n1195 0.019716
R55663 ASIG5V.n1201 ASIG5V.n1198 0.019716
R55664 ASIG5V.n1201 ASIG5V.n1200 0.019716
R55665 ASIG5V.n1208 ASIG5V.n886 0.019716
R55666 ASIG5V.n1209 ASIG5V.n1208 0.019716
R55667 ASIG5V.n1212 ASIG5V.n1211 0.019716
R55668 ASIG5V.n1213 ASIG5V.n1212 0.019716
R55669 ASIG5V.n1314 ASIG5V.n1313 0.019716
R55670 ASIG5V.n12025 ASIG5V.n1267 0.019716
R55671 ASIG5V.n12026 ASIG5V.n12025 0.019716
R55672 ASIG5V.n12031 ASIG5V.n1266 0.019716
R55673 ASIG5V.n12031 ASIG5V.n12030 0.019716
R55674 ASIG5V.n12037 ASIG5V.n1265 0.019716
R55675 ASIG5V.n12038 ASIG5V.n12037 0.019716
R55676 ASIG5V.n12043 ASIG5V.n1264 0.019716
R55677 ASIG5V.n12043 ASIG5V.n12042 0.019716
R55678 ASIG5V.n12049 ASIG5V.n1263 0.019716
R55679 ASIG5V.n12050 ASIG5V.n12049 0.019716
R55680 ASIG5V.n12055 ASIG5V.n1262 0.019716
R55681 ASIG5V.n12055 ASIG5V.n12054 0.019716
R55682 ASIG5V.n12061 ASIG5V.n1261 0.019716
R55683 ASIG5V.n12062 ASIG5V.n12061 0.019716
R55684 ASIG5V.n12067 ASIG5V.n1260 0.019716
R55685 ASIG5V.n12067 ASIG5V.n12066 0.019716
R55686 ASIG5V.n12073 ASIG5V.n1259 0.019716
R55687 ASIG5V.n12074 ASIG5V.n12073 0.019716
R55688 ASIG5V.n12079 ASIG5V.n1258 0.019716
R55689 ASIG5V.n12079 ASIG5V.n12078 0.019716
R55690 ASIG5V.n12085 ASIG5V.n1257 0.019716
R55691 ASIG5V.n12086 ASIG5V.n12085 0.019716
R55692 ASIG5V.n12091 ASIG5V.n1256 0.019716
R55693 ASIG5V.n12091 ASIG5V.n12090 0.019716
R55694 ASIG5V.n12097 ASIG5V.n1255 0.019716
R55695 ASIG5V.n12098 ASIG5V.n12097 0.019716
R55696 ASIG5V.n12103 ASIG5V.n1254 0.019716
R55697 ASIG5V.n12103 ASIG5V.n12102 0.019716
R55698 ASIG5V.n12109 ASIG5V.n1253 0.019716
R55699 ASIG5V.n12110 ASIG5V.n12109 0.019716
R55700 ASIG5V.n12115 ASIG5V.n1252 0.019716
R55701 ASIG5V.n12115 ASIG5V.n12114 0.019716
R55702 ASIG5V.n12121 ASIG5V.n1251 0.019716
R55703 ASIG5V.n12122 ASIG5V.n12121 0.019716
R55704 ASIG5V.n12127 ASIG5V.n1250 0.019716
R55705 ASIG5V.n12127 ASIG5V.n12126 0.019716
R55706 ASIG5V.n12133 ASIG5V.n1249 0.019716
R55707 ASIG5V.n12134 ASIG5V.n12133 0.019716
R55708 ASIG5V.n12139 ASIG5V.n1248 0.019716
R55709 ASIG5V.n12139 ASIG5V.n12138 0.019716
R55710 ASIG5V.n12145 ASIG5V.n1247 0.019716
R55711 ASIG5V.n12146 ASIG5V.n12145 0.019716
R55712 ASIG5V.n12151 ASIG5V.n1246 0.019716
R55713 ASIG5V.n12151 ASIG5V.n12150 0.019716
R55714 ASIG5V.n12157 ASIG5V.n1245 0.019716
R55715 ASIG5V.n12158 ASIG5V.n12157 0.019716
R55716 ASIG5V.n12163 ASIG5V.n1244 0.019716
R55717 ASIG5V.n12163 ASIG5V.n12162 0.019716
R55718 ASIG5V.n12169 ASIG5V.n1243 0.019716
R55719 ASIG5V.n12170 ASIG5V.n12169 0.019716
R55720 ASIG5V.n12175 ASIG5V.n1242 0.019716
R55721 ASIG5V.n12175 ASIG5V.n12174 0.019716
R55722 ASIG5V.n12181 ASIG5V.n1241 0.019716
R55723 ASIG5V.n12182 ASIG5V.n12181 0.019716
R55724 ASIG5V.n12187 ASIG5V.n1240 0.019716
R55725 ASIG5V.n12187 ASIG5V.n12186 0.019716
R55726 ASIG5V.n12193 ASIG5V.n1239 0.019716
R55727 ASIG5V.n12194 ASIG5V.n12193 0.019716
R55728 ASIG5V.n12199 ASIG5V.n1238 0.019716
R55729 ASIG5V.n12199 ASIG5V.n12198 0.019716
R55730 ASIG5V.n12205 ASIG5V.n1237 0.019716
R55731 ASIG5V.n12206 ASIG5V.n12205 0.019716
R55732 ASIG5V.n12211 ASIG5V.n1236 0.019716
R55733 ASIG5V.n12211 ASIG5V.n12210 0.019716
R55734 ASIG5V.n12217 ASIG5V.n1235 0.019716
R55735 ASIG5V.n12218 ASIG5V.n12217 0.019716
R55736 ASIG5V.n12223 ASIG5V.n1234 0.019716
R55737 ASIG5V.n12223 ASIG5V.n12222 0.019716
R55738 ASIG5V.n12229 ASIG5V.n1233 0.019716
R55739 ASIG5V.n12230 ASIG5V.n12229 0.019716
R55740 ASIG5V.n12235 ASIG5V.n1232 0.019716
R55741 ASIG5V.n12235 ASIG5V.n12234 0.019716
R55742 ASIG5V.n12241 ASIG5V.n1231 0.019716
R55743 ASIG5V.n12242 ASIG5V.n12241 0.019716
R55744 ASIG5V.n12247 ASIG5V.n1230 0.019716
R55745 ASIG5V.n12247 ASIG5V.n12246 0.019716
R55746 ASIG5V.n12253 ASIG5V.n1229 0.019716
R55747 ASIG5V.n12254 ASIG5V.n12253 0.019716
R55748 ASIG5V.n12259 ASIG5V.n1228 0.019716
R55749 ASIG5V.n12259 ASIG5V.n12258 0.019716
R55750 ASIG5V.n12265 ASIG5V.n1227 0.019716
R55751 ASIG5V.n12266 ASIG5V.n12265 0.019716
R55752 ASIG5V.n12010 ASIG5V.n1371 0.019716
R55753 ASIG5V.n1477 ASIG5V.n1414 0.019716
R55754 ASIG5V.n1477 ASIG5V.n1369 0.019716
R55755 ASIG5V.n1486 ASIG5V.n1413 0.019716
R55756 ASIG5V.n1486 ASIG5V.n1368 0.019716
R55757 ASIG5V.n1474 ASIG5V.n1412 0.019716
R55758 ASIG5V.n1474 ASIG5V.n1367 0.019716
R55759 ASIG5V.n1495 ASIG5V.n1411 0.019716
R55760 ASIG5V.n1495 ASIG5V.n1366 0.019716
R55761 ASIG5V.n1471 ASIG5V.n1410 0.019716
R55762 ASIG5V.n1471 ASIG5V.n1365 0.019716
R55763 ASIG5V.n1504 ASIG5V.n1409 0.019716
R55764 ASIG5V.n1504 ASIG5V.n1364 0.019716
R55765 ASIG5V.n1468 ASIG5V.n1408 0.019716
R55766 ASIG5V.n1468 ASIG5V.n1363 0.019716
R55767 ASIG5V.n1513 ASIG5V.n1407 0.019716
R55768 ASIG5V.n1513 ASIG5V.n1362 0.019716
R55769 ASIG5V.n1465 ASIG5V.n1406 0.019716
R55770 ASIG5V.n1465 ASIG5V.n1361 0.019716
R55771 ASIG5V.n1522 ASIG5V.n1405 0.019716
R55772 ASIG5V.n1522 ASIG5V.n1360 0.019716
R55773 ASIG5V.n1462 ASIG5V.n1404 0.019716
R55774 ASIG5V.n1462 ASIG5V.n1359 0.019716
R55775 ASIG5V.n1531 ASIG5V.n1403 0.019716
R55776 ASIG5V.n1531 ASIG5V.n1358 0.019716
R55777 ASIG5V.n1459 ASIG5V.n1402 0.019716
R55778 ASIG5V.n1459 ASIG5V.n1357 0.019716
R55779 ASIG5V.n1540 ASIG5V.n1401 0.019716
R55780 ASIG5V.n1540 ASIG5V.n1356 0.019716
R55781 ASIG5V.n1456 ASIG5V.n1400 0.019716
R55782 ASIG5V.n1456 ASIG5V.n1355 0.019716
R55783 ASIG5V.n1549 ASIG5V.n1399 0.019716
R55784 ASIG5V.n1549 ASIG5V.n1354 0.019716
R55785 ASIG5V.n1453 ASIG5V.n1398 0.019716
R55786 ASIG5V.n1453 ASIG5V.n1353 0.019716
R55787 ASIG5V.n1558 ASIG5V.n1397 0.019716
R55788 ASIG5V.n1558 ASIG5V.n1352 0.019716
R55789 ASIG5V.n1450 ASIG5V.n1396 0.019716
R55790 ASIG5V.n1450 ASIG5V.n1351 0.019716
R55791 ASIG5V.n1567 ASIG5V.n1395 0.019716
R55792 ASIG5V.n1567 ASIG5V.n1350 0.019716
R55793 ASIG5V.n1447 ASIG5V.n1394 0.019716
R55794 ASIG5V.n1447 ASIG5V.n1349 0.019716
R55795 ASIG5V.n1576 ASIG5V.n1393 0.019716
R55796 ASIG5V.n1576 ASIG5V.n1348 0.019716
R55797 ASIG5V.n1444 ASIG5V.n1392 0.019716
R55798 ASIG5V.n1444 ASIG5V.n1347 0.019716
R55799 ASIG5V.n1585 ASIG5V.n1391 0.019716
R55800 ASIG5V.n1585 ASIG5V.n1346 0.019716
R55801 ASIG5V.n1441 ASIG5V.n1390 0.019716
R55802 ASIG5V.n1441 ASIG5V.n1345 0.019716
R55803 ASIG5V.n1594 ASIG5V.n1389 0.019716
R55804 ASIG5V.n1594 ASIG5V.n1344 0.019716
R55805 ASIG5V.n1438 ASIG5V.n1388 0.019716
R55806 ASIG5V.n1438 ASIG5V.n1343 0.019716
R55807 ASIG5V.n1603 ASIG5V.n1387 0.019716
R55808 ASIG5V.n1603 ASIG5V.n1342 0.019716
R55809 ASIG5V.n1435 ASIG5V.n1386 0.019716
R55810 ASIG5V.n1435 ASIG5V.n1341 0.019716
R55811 ASIG5V.n1612 ASIG5V.n1385 0.019716
R55812 ASIG5V.n1612 ASIG5V.n1340 0.019716
R55813 ASIG5V.n1432 ASIG5V.n1384 0.019716
R55814 ASIG5V.n1432 ASIG5V.n1339 0.019716
R55815 ASIG5V.n1621 ASIG5V.n1383 0.019716
R55816 ASIG5V.n1621 ASIG5V.n1338 0.019716
R55817 ASIG5V.n1429 ASIG5V.n1382 0.019716
R55818 ASIG5V.n1429 ASIG5V.n1337 0.019716
R55819 ASIG5V.n1630 ASIG5V.n1381 0.019716
R55820 ASIG5V.n1630 ASIG5V.n1336 0.019716
R55821 ASIG5V.n1426 ASIG5V.n1380 0.019716
R55822 ASIG5V.n1426 ASIG5V.n1335 0.019716
R55823 ASIG5V.n1639 ASIG5V.n1379 0.019716
R55824 ASIG5V.n1639 ASIG5V.n1334 0.019716
R55825 ASIG5V.n1423 ASIG5V.n1378 0.019716
R55826 ASIG5V.n1423 ASIG5V.n1333 0.019716
R55827 ASIG5V.n1648 ASIG5V.n1377 0.019716
R55828 ASIG5V.n1648 ASIG5V.n1332 0.019716
R55829 ASIG5V.n1420 ASIG5V.n1376 0.019716
R55830 ASIG5V.n1420 ASIG5V.n1331 0.019716
R55831 ASIG5V.n1657 ASIG5V.n1375 0.019716
R55832 ASIG5V.n1657 ASIG5V.n1330 0.019716
R55833 ASIG5V.n1417 ASIG5V.n1374 0.019716
R55834 ASIG5V.n1417 ASIG5V.n1329 0.019716
R55835 ASIG5V.n11996 ASIG5V.n1718 0.019716
R55836 ASIG5V.n1824 ASIG5V.n1762 0.019716
R55837 ASIG5V.n1824 ASIG5V.n1716 0.019716
R55838 ASIG5V.n11814 ASIG5V.n1761 0.019716
R55839 ASIG5V.n11814 ASIG5V.n1715 0.019716
R55840 ASIG5V.n1821 ASIG5V.n1760 0.019716
R55841 ASIG5V.n1821 ASIG5V.n1714 0.019716
R55842 ASIG5V.n11823 ASIG5V.n1759 0.019716
R55843 ASIG5V.n11823 ASIG5V.n1713 0.019716
R55844 ASIG5V.n1818 ASIG5V.n1758 0.019716
R55845 ASIG5V.n1818 ASIG5V.n1712 0.019716
R55846 ASIG5V.n11832 ASIG5V.n1757 0.019716
R55847 ASIG5V.n11832 ASIG5V.n1711 0.019716
R55848 ASIG5V.n1815 ASIG5V.n1756 0.019716
R55849 ASIG5V.n1815 ASIG5V.n1710 0.019716
R55850 ASIG5V.n11841 ASIG5V.n1755 0.019716
R55851 ASIG5V.n11841 ASIG5V.n1709 0.019716
R55852 ASIG5V.n1812 ASIG5V.n1754 0.019716
R55853 ASIG5V.n1812 ASIG5V.n1708 0.019716
R55854 ASIG5V.n11850 ASIG5V.n1753 0.019716
R55855 ASIG5V.n11850 ASIG5V.n1707 0.019716
R55856 ASIG5V.n1809 ASIG5V.n1752 0.019716
R55857 ASIG5V.n1809 ASIG5V.n1706 0.019716
R55858 ASIG5V.n11859 ASIG5V.n1751 0.019716
R55859 ASIG5V.n11859 ASIG5V.n1705 0.019716
R55860 ASIG5V.n1806 ASIG5V.n1750 0.019716
R55861 ASIG5V.n1806 ASIG5V.n1704 0.019716
R55862 ASIG5V.n11868 ASIG5V.n1749 0.019716
R55863 ASIG5V.n11868 ASIG5V.n1703 0.019716
R55864 ASIG5V.n1803 ASIG5V.n1748 0.019716
R55865 ASIG5V.n1803 ASIG5V.n1702 0.019716
R55866 ASIG5V.n11877 ASIG5V.n1747 0.019716
R55867 ASIG5V.n11877 ASIG5V.n1701 0.019716
R55868 ASIG5V.n1800 ASIG5V.n1746 0.019716
R55869 ASIG5V.n1800 ASIG5V.n1700 0.019716
R55870 ASIG5V.n11886 ASIG5V.n1745 0.019716
R55871 ASIG5V.n11886 ASIG5V.n1699 0.019716
R55872 ASIG5V.n1797 ASIG5V.n1744 0.019716
R55873 ASIG5V.n1797 ASIG5V.n1698 0.019716
R55874 ASIG5V.n11895 ASIG5V.n1743 0.019716
R55875 ASIG5V.n11895 ASIG5V.n1697 0.019716
R55876 ASIG5V.n1794 ASIG5V.n1742 0.019716
R55877 ASIG5V.n1794 ASIG5V.n1696 0.019716
R55878 ASIG5V.n11904 ASIG5V.n1741 0.019716
R55879 ASIG5V.n11904 ASIG5V.n1695 0.019716
R55880 ASIG5V.n1791 ASIG5V.n1740 0.019716
R55881 ASIG5V.n1791 ASIG5V.n1694 0.019716
R55882 ASIG5V.n11913 ASIG5V.n1739 0.019716
R55883 ASIG5V.n11913 ASIG5V.n1693 0.019716
R55884 ASIG5V.n1788 ASIG5V.n1738 0.019716
R55885 ASIG5V.n1788 ASIG5V.n1692 0.019716
R55886 ASIG5V.n11922 ASIG5V.n1737 0.019716
R55887 ASIG5V.n11922 ASIG5V.n1691 0.019716
R55888 ASIG5V.n1785 ASIG5V.n1736 0.019716
R55889 ASIG5V.n1785 ASIG5V.n1690 0.019716
R55890 ASIG5V.n11931 ASIG5V.n1735 0.019716
R55891 ASIG5V.n11931 ASIG5V.n1689 0.019716
R55892 ASIG5V.n1782 ASIG5V.n1734 0.019716
R55893 ASIG5V.n1782 ASIG5V.n1688 0.019716
R55894 ASIG5V.n11940 ASIG5V.n1733 0.019716
R55895 ASIG5V.n11940 ASIG5V.n1687 0.019716
R55896 ASIG5V.n1779 ASIG5V.n1732 0.019716
R55897 ASIG5V.n1779 ASIG5V.n1686 0.019716
R55898 ASIG5V.n11949 ASIG5V.n1731 0.019716
R55899 ASIG5V.n11949 ASIG5V.n1685 0.019716
R55900 ASIG5V.n1776 ASIG5V.n1730 0.019716
R55901 ASIG5V.n1776 ASIG5V.n1684 0.019716
R55902 ASIG5V.n11958 ASIG5V.n1729 0.019716
R55903 ASIG5V.n11958 ASIG5V.n1683 0.019716
R55904 ASIG5V.n1773 ASIG5V.n1728 0.019716
R55905 ASIG5V.n1773 ASIG5V.n1682 0.019716
R55906 ASIG5V.n11967 ASIG5V.n1727 0.019716
R55907 ASIG5V.n11967 ASIG5V.n1681 0.019716
R55908 ASIG5V.n1770 ASIG5V.n1726 0.019716
R55909 ASIG5V.n1770 ASIG5V.n1680 0.019716
R55910 ASIG5V.n11976 ASIG5V.n1725 0.019716
R55911 ASIG5V.n11976 ASIG5V.n1679 0.019716
R55912 ASIG5V.n1767 ASIG5V.n1724 0.019716
R55913 ASIG5V.n1767 ASIG5V.n1678 0.019716
R55914 ASIG5V.n11985 ASIG5V.n1723 0.019716
R55915 ASIG5V.n11985 ASIG5V.n1677 0.019716
R55916 ASIG5V.n1764 ASIG5V.n1722 0.019716
R55917 ASIG5V.n1764 ASIG5V.n1676 0.019716
R55918 ASIG5V.n1950 ASIG5V.n1949 0.019716
R55919 ASIG5V.n1955 ASIG5V.n1905 0.019716
R55920 ASIG5V.n1956 ASIG5V.n1955 0.019716
R55921 ASIG5V.n1961 ASIG5V.n1904 0.019716
R55922 ASIG5V.n1961 ASIG5V.n1960 0.019716
R55923 ASIG5V.n1967 ASIG5V.n1903 0.019716
R55924 ASIG5V.n1968 ASIG5V.n1967 0.019716
R55925 ASIG5V.n1973 ASIG5V.n1902 0.019716
R55926 ASIG5V.n1973 ASIG5V.n1972 0.019716
R55927 ASIG5V.n1979 ASIG5V.n1901 0.019716
R55928 ASIG5V.n1980 ASIG5V.n1979 0.019716
R55929 ASIG5V.n1985 ASIG5V.n1900 0.019716
R55930 ASIG5V.n1985 ASIG5V.n1984 0.019716
R55931 ASIG5V.n1991 ASIG5V.n1899 0.019716
R55932 ASIG5V.n1992 ASIG5V.n1991 0.019716
R55933 ASIG5V.n1997 ASIG5V.n1898 0.019716
R55934 ASIG5V.n1997 ASIG5V.n1996 0.019716
R55935 ASIG5V.n2003 ASIG5V.n1897 0.019716
R55936 ASIG5V.n2004 ASIG5V.n2003 0.019716
R55937 ASIG5V.n2009 ASIG5V.n1896 0.019716
R55938 ASIG5V.n2009 ASIG5V.n2008 0.019716
R55939 ASIG5V.n2015 ASIG5V.n1895 0.019716
R55940 ASIG5V.n2016 ASIG5V.n2015 0.019716
R55941 ASIG5V.n2021 ASIG5V.n1894 0.019716
R55942 ASIG5V.n2021 ASIG5V.n2020 0.019716
R55943 ASIG5V.n2027 ASIG5V.n1893 0.019716
R55944 ASIG5V.n2028 ASIG5V.n2027 0.019716
R55945 ASIG5V.n2033 ASIG5V.n1892 0.019716
R55946 ASIG5V.n2033 ASIG5V.n2032 0.019716
R55947 ASIG5V.n2039 ASIG5V.n1891 0.019716
R55948 ASIG5V.n2040 ASIG5V.n2039 0.019716
R55949 ASIG5V.n2045 ASIG5V.n1890 0.019716
R55950 ASIG5V.n2045 ASIG5V.n2044 0.019716
R55951 ASIG5V.n2051 ASIG5V.n1889 0.019716
R55952 ASIG5V.n2052 ASIG5V.n2051 0.019716
R55953 ASIG5V.n2057 ASIG5V.n1888 0.019716
R55954 ASIG5V.n2057 ASIG5V.n2056 0.019716
R55955 ASIG5V.n2063 ASIG5V.n1887 0.019716
R55956 ASIG5V.n2064 ASIG5V.n2063 0.019716
R55957 ASIG5V.n2069 ASIG5V.n1886 0.019716
R55958 ASIG5V.n2069 ASIG5V.n2068 0.019716
R55959 ASIG5V.n2075 ASIG5V.n1885 0.019716
R55960 ASIG5V.n2076 ASIG5V.n2075 0.019716
R55961 ASIG5V.n2081 ASIG5V.n1884 0.019716
R55962 ASIG5V.n2081 ASIG5V.n2080 0.019716
R55963 ASIG5V.n2087 ASIG5V.n1883 0.019716
R55964 ASIG5V.n2088 ASIG5V.n2087 0.019716
R55965 ASIG5V.n2093 ASIG5V.n1882 0.019716
R55966 ASIG5V.n2093 ASIG5V.n2092 0.019716
R55967 ASIG5V.n2099 ASIG5V.n1881 0.019716
R55968 ASIG5V.n2100 ASIG5V.n2099 0.019716
R55969 ASIG5V.n2105 ASIG5V.n1880 0.019716
R55970 ASIG5V.n2105 ASIG5V.n2104 0.019716
R55971 ASIG5V.n2111 ASIG5V.n1879 0.019716
R55972 ASIG5V.n2112 ASIG5V.n2111 0.019716
R55973 ASIG5V.n2117 ASIG5V.n1878 0.019716
R55974 ASIG5V.n2117 ASIG5V.n2116 0.019716
R55975 ASIG5V.n2123 ASIG5V.n1877 0.019716
R55976 ASIG5V.n2124 ASIG5V.n2123 0.019716
R55977 ASIG5V.n2129 ASIG5V.n1876 0.019716
R55978 ASIG5V.n2129 ASIG5V.n2128 0.019716
R55979 ASIG5V.n2135 ASIG5V.n1875 0.019716
R55980 ASIG5V.n2136 ASIG5V.n2135 0.019716
R55981 ASIG5V.n2141 ASIG5V.n1874 0.019716
R55982 ASIG5V.n2141 ASIG5V.n2140 0.019716
R55983 ASIG5V.n2147 ASIG5V.n1873 0.019716
R55984 ASIG5V.n2148 ASIG5V.n2147 0.019716
R55985 ASIG5V.n2153 ASIG5V.n1872 0.019716
R55986 ASIG5V.n2153 ASIG5V.n2152 0.019716
R55987 ASIG5V.n2159 ASIG5V.n1871 0.019716
R55988 ASIG5V.n2160 ASIG5V.n2159 0.019716
R55989 ASIG5V.n2165 ASIG5V.n1870 0.019716
R55990 ASIG5V.n2165 ASIG5V.n2164 0.019716
R55991 ASIG5V.n2171 ASIG5V.n1869 0.019716
R55992 ASIG5V.n2172 ASIG5V.n2171 0.019716
R55993 ASIG5V.n2177 ASIG5V.n1868 0.019716
R55994 ASIG5V.n2177 ASIG5V.n2176 0.019716
R55995 ASIG5V.n2183 ASIG5V.n1867 0.019716
R55996 ASIG5V.n2184 ASIG5V.n2183 0.019716
R55997 ASIG5V.n2189 ASIG5V.n1866 0.019716
R55998 ASIG5V.n2189 ASIG5V.n2188 0.019716
R55999 ASIG5V.n2195 ASIG5V.n1865 0.019716
R56000 ASIG5V.n2196 ASIG5V.n2195 0.019716
R56001 ASIG5V.n2307 ASIG5V.n2306 0.019716
R56002 ASIG5V.n2312 ASIG5V.n2262 0.019716
R56003 ASIG5V.n2313 ASIG5V.n2312 0.019716
R56004 ASIG5V.n2318 ASIG5V.n2261 0.019716
R56005 ASIG5V.n2318 ASIG5V.n2317 0.019716
R56006 ASIG5V.n2324 ASIG5V.n2260 0.019716
R56007 ASIG5V.n2325 ASIG5V.n2324 0.019716
R56008 ASIG5V.n2330 ASIG5V.n2259 0.019716
R56009 ASIG5V.n2330 ASIG5V.n2329 0.019716
R56010 ASIG5V.n2336 ASIG5V.n2258 0.019716
R56011 ASIG5V.n2337 ASIG5V.n2336 0.019716
R56012 ASIG5V.n2342 ASIG5V.n2257 0.019716
R56013 ASIG5V.n2342 ASIG5V.n2341 0.019716
R56014 ASIG5V.n2348 ASIG5V.n2256 0.019716
R56015 ASIG5V.n2349 ASIG5V.n2348 0.019716
R56016 ASIG5V.n2354 ASIG5V.n2255 0.019716
R56017 ASIG5V.n2354 ASIG5V.n2353 0.019716
R56018 ASIG5V.n2360 ASIG5V.n2254 0.019716
R56019 ASIG5V.n2361 ASIG5V.n2360 0.019716
R56020 ASIG5V.n2366 ASIG5V.n2253 0.019716
R56021 ASIG5V.n2366 ASIG5V.n2365 0.019716
R56022 ASIG5V.n2372 ASIG5V.n2252 0.019716
R56023 ASIG5V.n2373 ASIG5V.n2372 0.019716
R56024 ASIG5V.n2378 ASIG5V.n2251 0.019716
R56025 ASIG5V.n2378 ASIG5V.n2377 0.019716
R56026 ASIG5V.n2384 ASIG5V.n2250 0.019716
R56027 ASIG5V.n2385 ASIG5V.n2384 0.019716
R56028 ASIG5V.n2390 ASIG5V.n2249 0.019716
R56029 ASIG5V.n2390 ASIG5V.n2389 0.019716
R56030 ASIG5V.n2396 ASIG5V.n2248 0.019716
R56031 ASIG5V.n2397 ASIG5V.n2396 0.019716
R56032 ASIG5V.n2402 ASIG5V.n2247 0.019716
R56033 ASIG5V.n2402 ASIG5V.n2401 0.019716
R56034 ASIG5V.n2408 ASIG5V.n2246 0.019716
R56035 ASIG5V.n2409 ASIG5V.n2408 0.019716
R56036 ASIG5V.n2414 ASIG5V.n2245 0.019716
R56037 ASIG5V.n2414 ASIG5V.n2413 0.019716
R56038 ASIG5V.n2420 ASIG5V.n2244 0.019716
R56039 ASIG5V.n2421 ASIG5V.n2420 0.019716
R56040 ASIG5V.n2426 ASIG5V.n2243 0.019716
R56041 ASIG5V.n2426 ASIG5V.n2425 0.019716
R56042 ASIG5V.n2432 ASIG5V.n2242 0.019716
R56043 ASIG5V.n2433 ASIG5V.n2432 0.019716
R56044 ASIG5V.n2438 ASIG5V.n2241 0.019716
R56045 ASIG5V.n2438 ASIG5V.n2437 0.019716
R56046 ASIG5V.n2444 ASIG5V.n2240 0.019716
R56047 ASIG5V.n2445 ASIG5V.n2444 0.019716
R56048 ASIG5V.n2450 ASIG5V.n2239 0.019716
R56049 ASIG5V.n2450 ASIG5V.n2449 0.019716
R56050 ASIG5V.n2456 ASIG5V.n2238 0.019716
R56051 ASIG5V.n2457 ASIG5V.n2456 0.019716
R56052 ASIG5V.n2462 ASIG5V.n2237 0.019716
R56053 ASIG5V.n2462 ASIG5V.n2461 0.019716
R56054 ASIG5V.n2468 ASIG5V.n2236 0.019716
R56055 ASIG5V.n2469 ASIG5V.n2468 0.019716
R56056 ASIG5V.n2474 ASIG5V.n2235 0.019716
R56057 ASIG5V.n2474 ASIG5V.n2473 0.019716
R56058 ASIG5V.n2480 ASIG5V.n2234 0.019716
R56059 ASIG5V.n2481 ASIG5V.n2480 0.019716
R56060 ASIG5V.n2486 ASIG5V.n2233 0.019716
R56061 ASIG5V.n2486 ASIG5V.n2485 0.019716
R56062 ASIG5V.n2492 ASIG5V.n2232 0.019716
R56063 ASIG5V.n2493 ASIG5V.n2492 0.019716
R56064 ASIG5V.n2498 ASIG5V.n2231 0.019716
R56065 ASIG5V.n2498 ASIG5V.n2497 0.019716
R56066 ASIG5V.n2504 ASIG5V.n2230 0.019716
R56067 ASIG5V.n2505 ASIG5V.n2504 0.019716
R56068 ASIG5V.n2510 ASIG5V.n2229 0.019716
R56069 ASIG5V.n2510 ASIG5V.n2509 0.019716
R56070 ASIG5V.n2516 ASIG5V.n2228 0.019716
R56071 ASIG5V.n2517 ASIG5V.n2516 0.019716
R56072 ASIG5V.n2522 ASIG5V.n2227 0.019716
R56073 ASIG5V.n2522 ASIG5V.n2521 0.019716
R56074 ASIG5V.n2528 ASIG5V.n2226 0.019716
R56075 ASIG5V.n2529 ASIG5V.n2528 0.019716
R56076 ASIG5V.n2534 ASIG5V.n2225 0.019716
R56077 ASIG5V.n2534 ASIG5V.n2533 0.019716
R56078 ASIG5V.n2540 ASIG5V.n2224 0.019716
R56079 ASIG5V.n2541 ASIG5V.n2540 0.019716
R56080 ASIG5V.n2546 ASIG5V.n2223 0.019716
R56081 ASIG5V.n2546 ASIG5V.n2545 0.019716
R56082 ASIG5V.n2552 ASIG5V.n2222 0.019716
R56083 ASIG5V.n2553 ASIG5V.n2552 0.019716
R56084 ASIG5V.n2659 ASIG5V.n2658 0.019716
R56085 ASIG5V.n2664 ASIG5V.n2610 0.019716
R56086 ASIG5V.n2665 ASIG5V.n2664 0.019716
R56087 ASIG5V.n2670 ASIG5V.n2609 0.019716
R56088 ASIG5V.n2670 ASIG5V.n2669 0.019716
R56089 ASIG5V.n2676 ASIG5V.n2608 0.019716
R56090 ASIG5V.n2677 ASIG5V.n2676 0.019716
R56091 ASIG5V.n2682 ASIG5V.n2607 0.019716
R56092 ASIG5V.n2682 ASIG5V.n2681 0.019716
R56093 ASIG5V.n2688 ASIG5V.n2606 0.019716
R56094 ASIG5V.n2689 ASIG5V.n2688 0.019716
R56095 ASIG5V.n2694 ASIG5V.n2605 0.019716
R56096 ASIG5V.n2694 ASIG5V.n2693 0.019716
R56097 ASIG5V.n2700 ASIG5V.n2604 0.019716
R56098 ASIG5V.n2701 ASIG5V.n2700 0.019716
R56099 ASIG5V.n2706 ASIG5V.n2603 0.019716
R56100 ASIG5V.n2706 ASIG5V.n2705 0.019716
R56101 ASIG5V.n2712 ASIG5V.n2602 0.019716
R56102 ASIG5V.n2713 ASIG5V.n2712 0.019716
R56103 ASIG5V.n2718 ASIG5V.n2601 0.019716
R56104 ASIG5V.n2718 ASIG5V.n2717 0.019716
R56105 ASIG5V.n2724 ASIG5V.n2600 0.019716
R56106 ASIG5V.n2725 ASIG5V.n2724 0.019716
R56107 ASIG5V.n2730 ASIG5V.n2599 0.019716
R56108 ASIG5V.n2730 ASIG5V.n2729 0.019716
R56109 ASIG5V.n2736 ASIG5V.n2598 0.019716
R56110 ASIG5V.n2737 ASIG5V.n2736 0.019716
R56111 ASIG5V.n2742 ASIG5V.n2597 0.019716
R56112 ASIG5V.n2742 ASIG5V.n2741 0.019716
R56113 ASIG5V.n2748 ASIG5V.n2596 0.019716
R56114 ASIG5V.n2749 ASIG5V.n2748 0.019716
R56115 ASIG5V.n2754 ASIG5V.n2595 0.019716
R56116 ASIG5V.n2754 ASIG5V.n2753 0.019716
R56117 ASIG5V.n2760 ASIG5V.n2594 0.019716
R56118 ASIG5V.n2761 ASIG5V.n2760 0.019716
R56119 ASIG5V.n2766 ASIG5V.n2593 0.019716
R56120 ASIG5V.n2766 ASIG5V.n2765 0.019716
R56121 ASIG5V.n2772 ASIG5V.n2592 0.019716
R56122 ASIG5V.n2773 ASIG5V.n2772 0.019716
R56123 ASIG5V.n2778 ASIG5V.n2591 0.019716
R56124 ASIG5V.n2778 ASIG5V.n2777 0.019716
R56125 ASIG5V.n2784 ASIG5V.n2590 0.019716
R56126 ASIG5V.n2785 ASIG5V.n2784 0.019716
R56127 ASIG5V.n2790 ASIG5V.n2589 0.019716
R56128 ASIG5V.n2790 ASIG5V.n2789 0.019716
R56129 ASIG5V.n2796 ASIG5V.n2588 0.019716
R56130 ASIG5V.n2797 ASIG5V.n2796 0.019716
R56131 ASIG5V.n2802 ASIG5V.n2587 0.019716
R56132 ASIG5V.n2802 ASIG5V.n2801 0.019716
R56133 ASIG5V.n2808 ASIG5V.n2586 0.019716
R56134 ASIG5V.n2809 ASIG5V.n2808 0.019716
R56135 ASIG5V.n2814 ASIG5V.n2585 0.019716
R56136 ASIG5V.n2814 ASIG5V.n2813 0.019716
R56137 ASIG5V.n2820 ASIG5V.n2584 0.019716
R56138 ASIG5V.n2821 ASIG5V.n2820 0.019716
R56139 ASIG5V.n2826 ASIG5V.n2583 0.019716
R56140 ASIG5V.n2826 ASIG5V.n2825 0.019716
R56141 ASIG5V.n2832 ASIG5V.n2582 0.019716
R56142 ASIG5V.n2833 ASIG5V.n2832 0.019716
R56143 ASIG5V.n2838 ASIG5V.n2581 0.019716
R56144 ASIG5V.n2838 ASIG5V.n2837 0.019716
R56145 ASIG5V.n2844 ASIG5V.n2580 0.019716
R56146 ASIG5V.n2845 ASIG5V.n2844 0.019716
R56147 ASIG5V.n2850 ASIG5V.n2579 0.019716
R56148 ASIG5V.n2850 ASIG5V.n2849 0.019716
R56149 ASIG5V.n2856 ASIG5V.n2578 0.019716
R56150 ASIG5V.n2857 ASIG5V.n2856 0.019716
R56151 ASIG5V.n2862 ASIG5V.n2577 0.019716
R56152 ASIG5V.n2862 ASIG5V.n2861 0.019716
R56153 ASIG5V.n2868 ASIG5V.n2576 0.019716
R56154 ASIG5V.n2869 ASIG5V.n2868 0.019716
R56155 ASIG5V.n2874 ASIG5V.n2575 0.019716
R56156 ASIG5V.n2874 ASIG5V.n2873 0.019716
R56157 ASIG5V.n2880 ASIG5V.n2574 0.019716
R56158 ASIG5V.n2881 ASIG5V.n2880 0.019716
R56159 ASIG5V.n2886 ASIG5V.n2573 0.019716
R56160 ASIG5V.n2886 ASIG5V.n2885 0.019716
R56161 ASIG5V.n2892 ASIG5V.n2572 0.019716
R56162 ASIG5V.n2893 ASIG5V.n2892 0.019716
R56163 ASIG5V.n2898 ASIG5V.n2571 0.019716
R56164 ASIG5V.n2898 ASIG5V.n2897 0.019716
R56165 ASIG5V.n11768 ASIG5V.n2570 0.019716
R56166 ASIG5V.n11769 ASIG5V.n11768 0.019716
R56167 ASIG5V.n3000 ASIG5V.n2999 0.019716
R56168 ASIG5V.n11508 ASIG5V.n2954 0.019716
R56169 ASIG5V.n11509 ASIG5V.n11508 0.019716
R56170 ASIG5V.n11514 ASIG5V.n2953 0.019716
R56171 ASIG5V.n11514 ASIG5V.n11513 0.019716
R56172 ASIG5V.n11520 ASIG5V.n2952 0.019716
R56173 ASIG5V.n11521 ASIG5V.n11520 0.019716
R56174 ASIG5V.n11526 ASIG5V.n2951 0.019716
R56175 ASIG5V.n11526 ASIG5V.n11525 0.019716
R56176 ASIG5V.n11532 ASIG5V.n2950 0.019716
R56177 ASIG5V.n11533 ASIG5V.n11532 0.019716
R56178 ASIG5V.n11538 ASIG5V.n2949 0.019716
R56179 ASIG5V.n11538 ASIG5V.n11537 0.019716
R56180 ASIG5V.n11544 ASIG5V.n2948 0.019716
R56181 ASIG5V.n11545 ASIG5V.n11544 0.019716
R56182 ASIG5V.n11550 ASIG5V.n2947 0.019716
R56183 ASIG5V.n11550 ASIG5V.n11549 0.019716
R56184 ASIG5V.n11556 ASIG5V.n2946 0.019716
R56185 ASIG5V.n11557 ASIG5V.n11556 0.019716
R56186 ASIG5V.n11562 ASIG5V.n2945 0.019716
R56187 ASIG5V.n11562 ASIG5V.n11561 0.019716
R56188 ASIG5V.n11568 ASIG5V.n2944 0.019716
R56189 ASIG5V.n11569 ASIG5V.n11568 0.019716
R56190 ASIG5V.n11574 ASIG5V.n2943 0.019716
R56191 ASIG5V.n11574 ASIG5V.n11573 0.019716
R56192 ASIG5V.n11580 ASIG5V.n2942 0.019716
R56193 ASIG5V.n11581 ASIG5V.n11580 0.019716
R56194 ASIG5V.n11586 ASIG5V.n2941 0.019716
R56195 ASIG5V.n11586 ASIG5V.n11585 0.019716
R56196 ASIG5V.n11592 ASIG5V.n2940 0.019716
R56197 ASIG5V.n11593 ASIG5V.n11592 0.019716
R56198 ASIG5V.n11598 ASIG5V.n2939 0.019716
R56199 ASIG5V.n11598 ASIG5V.n11597 0.019716
R56200 ASIG5V.n11604 ASIG5V.n2938 0.019716
R56201 ASIG5V.n11605 ASIG5V.n11604 0.019716
R56202 ASIG5V.n11610 ASIG5V.n2937 0.019716
R56203 ASIG5V.n11610 ASIG5V.n11609 0.019716
R56204 ASIG5V.n11616 ASIG5V.n2936 0.019716
R56205 ASIG5V.n11617 ASIG5V.n11616 0.019716
R56206 ASIG5V.n11622 ASIG5V.n2935 0.019716
R56207 ASIG5V.n11622 ASIG5V.n11621 0.019716
R56208 ASIG5V.n11628 ASIG5V.n2934 0.019716
R56209 ASIG5V.n11629 ASIG5V.n11628 0.019716
R56210 ASIG5V.n11634 ASIG5V.n2933 0.019716
R56211 ASIG5V.n11634 ASIG5V.n11633 0.019716
R56212 ASIG5V.n11640 ASIG5V.n2932 0.019716
R56213 ASIG5V.n11641 ASIG5V.n11640 0.019716
R56214 ASIG5V.n11646 ASIG5V.n2931 0.019716
R56215 ASIG5V.n11646 ASIG5V.n11645 0.019716
R56216 ASIG5V.n11652 ASIG5V.n2930 0.019716
R56217 ASIG5V.n11653 ASIG5V.n11652 0.019716
R56218 ASIG5V.n11658 ASIG5V.n2929 0.019716
R56219 ASIG5V.n11658 ASIG5V.n11657 0.019716
R56220 ASIG5V.n11664 ASIG5V.n2928 0.019716
R56221 ASIG5V.n11665 ASIG5V.n11664 0.019716
R56222 ASIG5V.n11670 ASIG5V.n2927 0.019716
R56223 ASIG5V.n11670 ASIG5V.n11669 0.019716
R56224 ASIG5V.n11676 ASIG5V.n2926 0.019716
R56225 ASIG5V.n11677 ASIG5V.n11676 0.019716
R56226 ASIG5V.n11682 ASIG5V.n2925 0.019716
R56227 ASIG5V.n11682 ASIG5V.n11681 0.019716
R56228 ASIG5V.n11688 ASIG5V.n2924 0.019716
R56229 ASIG5V.n11689 ASIG5V.n11688 0.019716
R56230 ASIG5V.n11694 ASIG5V.n2923 0.019716
R56231 ASIG5V.n11694 ASIG5V.n11693 0.019716
R56232 ASIG5V.n11700 ASIG5V.n2922 0.019716
R56233 ASIG5V.n11701 ASIG5V.n11700 0.019716
R56234 ASIG5V.n11706 ASIG5V.n2921 0.019716
R56235 ASIG5V.n11706 ASIG5V.n11705 0.019716
R56236 ASIG5V.n11712 ASIG5V.n2920 0.019716
R56237 ASIG5V.n11713 ASIG5V.n11712 0.019716
R56238 ASIG5V.n11718 ASIG5V.n2919 0.019716
R56239 ASIG5V.n11718 ASIG5V.n11717 0.019716
R56240 ASIG5V.n11724 ASIG5V.n2918 0.019716
R56241 ASIG5V.n11725 ASIG5V.n11724 0.019716
R56242 ASIG5V.n11730 ASIG5V.n2917 0.019716
R56243 ASIG5V.n11730 ASIG5V.n11729 0.019716
R56244 ASIG5V.n11736 ASIG5V.n2916 0.019716
R56245 ASIG5V.n11737 ASIG5V.n11736 0.019716
R56246 ASIG5V.n11742 ASIG5V.n2915 0.019716
R56247 ASIG5V.n11742 ASIG5V.n11741 0.019716
R56248 ASIG5V.n11748 ASIG5V.n2914 0.019716
R56249 ASIG5V.n11749 ASIG5V.n11748 0.019716
R56250 ASIG5V.n11235 ASIG5V.n11234 0.019716
R56251 ASIG5V.n11242 ASIG5V.n10014 0.019716
R56252 ASIG5V.n11243 ASIG5V.n11242 0.019716
R56253 ASIG5V.n11248 ASIG5V.n10013 0.019716
R56254 ASIG5V.n11248 ASIG5V.n11247 0.019716
R56255 ASIG5V.n11254 ASIG5V.n10012 0.019716
R56256 ASIG5V.n11255 ASIG5V.n11254 0.019716
R56257 ASIG5V.n11260 ASIG5V.n10011 0.019716
R56258 ASIG5V.n11260 ASIG5V.n11259 0.019716
R56259 ASIG5V.n11266 ASIG5V.n10010 0.019716
R56260 ASIG5V.n11267 ASIG5V.n11266 0.019716
R56261 ASIG5V.n11272 ASIG5V.n10009 0.019716
R56262 ASIG5V.n11272 ASIG5V.n11271 0.019716
R56263 ASIG5V.n11278 ASIG5V.n10008 0.019716
R56264 ASIG5V.n11279 ASIG5V.n11278 0.019716
R56265 ASIG5V.n11284 ASIG5V.n10007 0.019716
R56266 ASIG5V.n11284 ASIG5V.n11283 0.019716
R56267 ASIG5V.n11290 ASIG5V.n10006 0.019716
R56268 ASIG5V.n11291 ASIG5V.n11290 0.019716
R56269 ASIG5V.n11296 ASIG5V.n10005 0.019716
R56270 ASIG5V.n11296 ASIG5V.n11295 0.019716
R56271 ASIG5V.n11302 ASIG5V.n10004 0.019716
R56272 ASIG5V.n11303 ASIG5V.n11302 0.019716
R56273 ASIG5V.n11308 ASIG5V.n10003 0.019716
R56274 ASIG5V.n11308 ASIG5V.n11307 0.019716
R56275 ASIG5V.n11314 ASIG5V.n10002 0.019716
R56276 ASIG5V.n11315 ASIG5V.n11314 0.019716
R56277 ASIG5V.n11320 ASIG5V.n10001 0.019716
R56278 ASIG5V.n11320 ASIG5V.n11319 0.019716
R56279 ASIG5V.n11326 ASIG5V.n10000 0.019716
R56280 ASIG5V.n11327 ASIG5V.n11326 0.019716
R56281 ASIG5V.n11332 ASIG5V.n9999 0.019716
R56282 ASIG5V.n11332 ASIG5V.n11331 0.019716
R56283 ASIG5V.n11338 ASIG5V.n9998 0.019716
R56284 ASIG5V.n11339 ASIG5V.n11338 0.019716
R56285 ASIG5V.n11344 ASIG5V.n9997 0.019716
R56286 ASIG5V.n11344 ASIG5V.n11343 0.019716
R56287 ASIG5V.n11350 ASIG5V.n9996 0.019716
R56288 ASIG5V.n11351 ASIG5V.n11350 0.019716
R56289 ASIG5V.n11356 ASIG5V.n9995 0.019716
R56290 ASIG5V.n11356 ASIG5V.n11355 0.019716
R56291 ASIG5V.n11362 ASIG5V.n9994 0.019716
R56292 ASIG5V.n11363 ASIG5V.n11362 0.019716
R56293 ASIG5V.n11368 ASIG5V.n9993 0.019716
R56294 ASIG5V.n11368 ASIG5V.n11367 0.019716
R56295 ASIG5V.n11374 ASIG5V.n9992 0.019716
R56296 ASIG5V.n11375 ASIG5V.n11374 0.019716
R56297 ASIG5V.n11380 ASIG5V.n9991 0.019716
R56298 ASIG5V.n11380 ASIG5V.n11379 0.019716
R56299 ASIG5V.n11386 ASIG5V.n9990 0.019716
R56300 ASIG5V.n11387 ASIG5V.n11386 0.019716
R56301 ASIG5V.n11392 ASIG5V.n9989 0.019716
R56302 ASIG5V.n11392 ASIG5V.n11391 0.019716
R56303 ASIG5V.n11398 ASIG5V.n9988 0.019716
R56304 ASIG5V.n11399 ASIG5V.n11398 0.019716
R56305 ASIG5V.n11404 ASIG5V.n9987 0.019716
R56306 ASIG5V.n11404 ASIG5V.n11403 0.019716
R56307 ASIG5V.n11410 ASIG5V.n9986 0.019716
R56308 ASIG5V.n11411 ASIG5V.n11410 0.019716
R56309 ASIG5V.n11416 ASIG5V.n9985 0.019716
R56310 ASIG5V.n11416 ASIG5V.n11415 0.019716
R56311 ASIG5V.n11422 ASIG5V.n9984 0.019716
R56312 ASIG5V.n11423 ASIG5V.n11422 0.019716
R56313 ASIG5V.n11428 ASIG5V.n9983 0.019716
R56314 ASIG5V.n11428 ASIG5V.n11427 0.019716
R56315 ASIG5V.n11434 ASIG5V.n9982 0.019716
R56316 ASIG5V.n11435 ASIG5V.n11434 0.019716
R56317 ASIG5V.n11440 ASIG5V.n9981 0.019716
R56318 ASIG5V.n11440 ASIG5V.n11439 0.019716
R56319 ASIG5V.n11446 ASIG5V.n9980 0.019716
R56320 ASIG5V.n11447 ASIG5V.n11446 0.019716
R56321 ASIG5V.n11452 ASIG5V.n9979 0.019716
R56322 ASIG5V.n11452 ASIG5V.n11451 0.019716
R56323 ASIG5V.n11458 ASIG5V.n9978 0.019716
R56324 ASIG5V.n11459 ASIG5V.n11458 0.019716
R56325 ASIG5V.n11464 ASIG5V.n9977 0.019716
R56326 ASIG5V.n11464 ASIG5V.n11463 0.019716
R56327 ASIG5V.n11470 ASIG5V.n9976 0.019716
R56328 ASIG5V.n11471 ASIG5V.n11470 0.019716
R56329 ASIG5V.n11476 ASIG5V.n9975 0.019716
R56330 ASIG5V.n11476 ASIG5V.n11475 0.019716
R56331 ASIG5V.n11482 ASIG5V.n9974 0.019716
R56332 ASIG5V.n11483 ASIG5V.n11482 0.019716
R56333 ASIG5V.n10355 ASIG5V.n10354 0.019716
R56334 ASIG5V.n10117 ASIG5V.n10066 0.019716
R56335 ASIG5V.n10117 ASIG5V.n10115 0.019716
R56336 ASIG5V.n10346 ASIG5V.n10065 0.019716
R56337 ASIG5V.n10346 ASIG5V.n10114 0.019716
R56338 ASIG5V.n10121 ASIG5V.n10064 0.019716
R56339 ASIG5V.n10121 ASIG5V.n10113 0.019716
R56340 ASIG5V.n10337 ASIG5V.n10063 0.019716
R56341 ASIG5V.n10337 ASIG5V.n10112 0.019716
R56342 ASIG5V.n10124 ASIG5V.n10062 0.019716
R56343 ASIG5V.n10124 ASIG5V.n10111 0.019716
R56344 ASIG5V.n10328 ASIG5V.n10061 0.019716
R56345 ASIG5V.n10328 ASIG5V.n10110 0.019716
R56346 ASIG5V.n10127 ASIG5V.n10060 0.019716
R56347 ASIG5V.n10127 ASIG5V.n10109 0.019716
R56348 ASIG5V.n10319 ASIG5V.n10059 0.019716
R56349 ASIG5V.n10319 ASIG5V.n10108 0.019716
R56350 ASIG5V.n10130 ASIG5V.n10058 0.019716
R56351 ASIG5V.n10130 ASIG5V.n10107 0.019716
R56352 ASIG5V.n10310 ASIG5V.n10057 0.019716
R56353 ASIG5V.n10310 ASIG5V.n10106 0.019716
R56354 ASIG5V.n10133 ASIG5V.n10056 0.019716
R56355 ASIG5V.n10133 ASIG5V.n10105 0.019716
R56356 ASIG5V.n10301 ASIG5V.n10055 0.019716
R56357 ASIG5V.n10301 ASIG5V.n10104 0.019716
R56358 ASIG5V.n10136 ASIG5V.n10054 0.019716
R56359 ASIG5V.n10136 ASIG5V.n10103 0.019716
R56360 ASIG5V.n10292 ASIG5V.n10053 0.019716
R56361 ASIG5V.n10292 ASIG5V.n10102 0.019716
R56362 ASIG5V.n10139 ASIG5V.n10052 0.019716
R56363 ASIG5V.n10139 ASIG5V.n10101 0.019716
R56364 ASIG5V.n10283 ASIG5V.n10051 0.019716
R56365 ASIG5V.n10283 ASIG5V.n10100 0.019716
R56366 ASIG5V.n10142 ASIG5V.n10050 0.019716
R56367 ASIG5V.n10142 ASIG5V.n10099 0.019716
R56368 ASIG5V.n10274 ASIG5V.n10049 0.019716
R56369 ASIG5V.n10274 ASIG5V.n10098 0.019716
R56370 ASIG5V.n10145 ASIG5V.n10048 0.019716
R56371 ASIG5V.n10145 ASIG5V.n10097 0.019716
R56372 ASIG5V.n10265 ASIG5V.n10047 0.019716
R56373 ASIG5V.n10265 ASIG5V.n10096 0.019716
R56374 ASIG5V.n10148 ASIG5V.n10046 0.019716
R56375 ASIG5V.n10148 ASIG5V.n10095 0.019716
R56376 ASIG5V.n10256 ASIG5V.n10045 0.019716
R56377 ASIG5V.n10256 ASIG5V.n10094 0.019716
R56378 ASIG5V.n10151 ASIG5V.n10044 0.019716
R56379 ASIG5V.n10151 ASIG5V.n10093 0.019716
R56380 ASIG5V.n10247 ASIG5V.n10043 0.019716
R56381 ASIG5V.n10247 ASIG5V.n10092 0.019716
R56382 ASIG5V.n10154 ASIG5V.n10042 0.019716
R56383 ASIG5V.n10154 ASIG5V.n10091 0.019716
R56384 ASIG5V.n10238 ASIG5V.n10041 0.019716
R56385 ASIG5V.n10238 ASIG5V.n10090 0.019716
R56386 ASIG5V.n10157 ASIG5V.n10040 0.019716
R56387 ASIG5V.n10157 ASIG5V.n10089 0.019716
R56388 ASIG5V.n10229 ASIG5V.n10039 0.019716
R56389 ASIG5V.n10229 ASIG5V.n10088 0.019716
R56390 ASIG5V.n10160 ASIG5V.n10038 0.019716
R56391 ASIG5V.n10160 ASIG5V.n10087 0.019716
R56392 ASIG5V.n10220 ASIG5V.n10037 0.019716
R56393 ASIG5V.n10220 ASIG5V.n10086 0.019716
R56394 ASIG5V.n10163 ASIG5V.n10036 0.019716
R56395 ASIG5V.n10163 ASIG5V.n10085 0.019716
R56396 ASIG5V.n10211 ASIG5V.n10035 0.019716
R56397 ASIG5V.n10211 ASIG5V.n10084 0.019716
R56398 ASIG5V.n10166 ASIG5V.n10034 0.019716
R56399 ASIG5V.n10166 ASIG5V.n10083 0.019716
R56400 ASIG5V.n10202 ASIG5V.n10033 0.019716
R56401 ASIG5V.n10202 ASIG5V.n10082 0.019716
R56402 ASIG5V.n10169 ASIG5V.n10032 0.019716
R56403 ASIG5V.n10169 ASIG5V.n10081 0.019716
R56404 ASIG5V.n10193 ASIG5V.n10031 0.019716
R56405 ASIG5V.n10193 ASIG5V.n10080 0.019716
R56406 ASIG5V.n10172 ASIG5V.n10030 0.019716
R56407 ASIG5V.n10172 ASIG5V.n10079 0.019716
R56408 ASIG5V.n10184 ASIG5V.n10029 0.019716
R56409 ASIG5V.n10184 ASIG5V.n10078 0.019716
R56410 ASIG5V.n10175 ASIG5V.n10028 0.019716
R56411 ASIG5V.n10175 ASIG5V.n10077 0.019716
R56412 ASIG5V.n10075 ASIG5V.n10027 0.019716
R56413 ASIG5V.n10357 ASIG5V.n10075 0.019716
R56414 ASIG5V.n10071 ASIG5V.n10026 0.019716
R56415 ASIG5V.n10071 ASIG5V.n10070 0.019716
R56416 ASIG5V.n10355 ASIG5V.n10067 0.019716
R56417 ASIG5V.n10354 ASIG5V.n10066 0.019716
R56418 ASIG5V.n10348 ASIG5V.n10065 0.019716
R56419 ASIG5V.n10348 ASIG5V.n10115 0.019716
R56420 ASIG5V.n10344 ASIG5V.n10064 0.019716
R56421 ASIG5V.n10344 ASIG5V.n10114 0.019716
R56422 ASIG5V.n10339 ASIG5V.n10063 0.019716
R56423 ASIG5V.n10339 ASIG5V.n10113 0.019716
R56424 ASIG5V.n10335 ASIG5V.n10062 0.019716
R56425 ASIG5V.n10335 ASIG5V.n10112 0.019716
R56426 ASIG5V.n10330 ASIG5V.n10061 0.019716
R56427 ASIG5V.n10330 ASIG5V.n10111 0.019716
R56428 ASIG5V.n10326 ASIG5V.n10060 0.019716
R56429 ASIG5V.n10326 ASIG5V.n10110 0.019716
R56430 ASIG5V.n10321 ASIG5V.n10059 0.019716
R56431 ASIG5V.n10321 ASIG5V.n10109 0.019716
R56432 ASIG5V.n10317 ASIG5V.n10058 0.019716
R56433 ASIG5V.n10317 ASIG5V.n10108 0.019716
R56434 ASIG5V.n10312 ASIG5V.n10057 0.019716
R56435 ASIG5V.n10312 ASIG5V.n10107 0.019716
R56436 ASIG5V.n10308 ASIG5V.n10056 0.019716
R56437 ASIG5V.n10308 ASIG5V.n10106 0.019716
R56438 ASIG5V.n10303 ASIG5V.n10055 0.019716
R56439 ASIG5V.n10303 ASIG5V.n10105 0.019716
R56440 ASIG5V.n10299 ASIG5V.n10054 0.019716
R56441 ASIG5V.n10299 ASIG5V.n10104 0.019716
R56442 ASIG5V.n10294 ASIG5V.n10053 0.019716
R56443 ASIG5V.n10294 ASIG5V.n10103 0.019716
R56444 ASIG5V.n10290 ASIG5V.n10052 0.019716
R56445 ASIG5V.n10290 ASIG5V.n10102 0.019716
R56446 ASIG5V.n10285 ASIG5V.n10051 0.019716
R56447 ASIG5V.n10285 ASIG5V.n10101 0.019716
R56448 ASIG5V.n10281 ASIG5V.n10050 0.019716
R56449 ASIG5V.n10281 ASIG5V.n10100 0.019716
R56450 ASIG5V.n10276 ASIG5V.n10049 0.019716
R56451 ASIG5V.n10276 ASIG5V.n10099 0.019716
R56452 ASIG5V.n10272 ASIG5V.n10048 0.019716
R56453 ASIG5V.n10272 ASIG5V.n10098 0.019716
R56454 ASIG5V.n10267 ASIG5V.n10047 0.019716
R56455 ASIG5V.n10267 ASIG5V.n10097 0.019716
R56456 ASIG5V.n10263 ASIG5V.n10046 0.019716
R56457 ASIG5V.n10263 ASIG5V.n10096 0.019716
R56458 ASIG5V.n10258 ASIG5V.n10045 0.019716
R56459 ASIG5V.n10258 ASIG5V.n10095 0.019716
R56460 ASIG5V.n10254 ASIG5V.n10044 0.019716
R56461 ASIG5V.n10254 ASIG5V.n10094 0.019716
R56462 ASIG5V.n10249 ASIG5V.n10043 0.019716
R56463 ASIG5V.n10249 ASIG5V.n10093 0.019716
R56464 ASIG5V.n10245 ASIG5V.n10042 0.019716
R56465 ASIG5V.n10245 ASIG5V.n10092 0.019716
R56466 ASIG5V.n10240 ASIG5V.n10041 0.019716
R56467 ASIG5V.n10240 ASIG5V.n10091 0.019716
R56468 ASIG5V.n10236 ASIG5V.n10040 0.019716
R56469 ASIG5V.n10236 ASIG5V.n10090 0.019716
R56470 ASIG5V.n10231 ASIG5V.n10039 0.019716
R56471 ASIG5V.n10231 ASIG5V.n10089 0.019716
R56472 ASIG5V.n10227 ASIG5V.n10038 0.019716
R56473 ASIG5V.n10227 ASIG5V.n10088 0.019716
R56474 ASIG5V.n10222 ASIG5V.n10037 0.019716
R56475 ASIG5V.n10222 ASIG5V.n10087 0.019716
R56476 ASIG5V.n10218 ASIG5V.n10036 0.019716
R56477 ASIG5V.n10218 ASIG5V.n10086 0.019716
R56478 ASIG5V.n10213 ASIG5V.n10035 0.019716
R56479 ASIG5V.n10213 ASIG5V.n10085 0.019716
R56480 ASIG5V.n10209 ASIG5V.n10034 0.019716
R56481 ASIG5V.n10209 ASIG5V.n10084 0.019716
R56482 ASIG5V.n10204 ASIG5V.n10033 0.019716
R56483 ASIG5V.n10204 ASIG5V.n10083 0.019716
R56484 ASIG5V.n10200 ASIG5V.n10032 0.019716
R56485 ASIG5V.n10200 ASIG5V.n10082 0.019716
R56486 ASIG5V.n10195 ASIG5V.n10031 0.019716
R56487 ASIG5V.n10195 ASIG5V.n10081 0.019716
R56488 ASIG5V.n10191 ASIG5V.n10030 0.019716
R56489 ASIG5V.n10191 ASIG5V.n10080 0.019716
R56490 ASIG5V.n10186 ASIG5V.n10029 0.019716
R56491 ASIG5V.n10186 ASIG5V.n10079 0.019716
R56492 ASIG5V.n10182 ASIG5V.n10028 0.019716
R56493 ASIG5V.n10182 ASIG5V.n10078 0.019716
R56494 ASIG5V.n10177 ASIG5V.n10027 0.019716
R56495 ASIG5V.n10177 ASIG5V.n10077 0.019716
R56496 ASIG5V.n10358 ASIG5V.n10026 0.019716
R56497 ASIG5V.n10358 ASIG5V.n10357 0.019716
R56498 ASIG5V.n11182 ASIG5V.n10070 0.019716
R56499 ASIG5V.n11234 ASIG5V.n10015 0.019716
R56500 ASIG5V.n11235 ASIG5V.n10014 0.019716
R56501 ASIG5V.n11244 ASIG5V.n10013 0.019716
R56502 ASIG5V.n11244 ASIG5V.n11243 0.019716
R56503 ASIG5V.n11246 ASIG5V.n10012 0.019716
R56504 ASIG5V.n11247 ASIG5V.n11246 0.019716
R56505 ASIG5V.n11256 ASIG5V.n10011 0.019716
R56506 ASIG5V.n11256 ASIG5V.n11255 0.019716
R56507 ASIG5V.n11258 ASIG5V.n10010 0.019716
R56508 ASIG5V.n11259 ASIG5V.n11258 0.019716
R56509 ASIG5V.n11268 ASIG5V.n10009 0.019716
R56510 ASIG5V.n11268 ASIG5V.n11267 0.019716
R56511 ASIG5V.n11270 ASIG5V.n10008 0.019716
R56512 ASIG5V.n11271 ASIG5V.n11270 0.019716
R56513 ASIG5V.n11280 ASIG5V.n10007 0.019716
R56514 ASIG5V.n11280 ASIG5V.n11279 0.019716
R56515 ASIG5V.n11282 ASIG5V.n10006 0.019716
R56516 ASIG5V.n11283 ASIG5V.n11282 0.019716
R56517 ASIG5V.n11292 ASIG5V.n10005 0.019716
R56518 ASIG5V.n11292 ASIG5V.n11291 0.019716
R56519 ASIG5V.n11294 ASIG5V.n10004 0.019716
R56520 ASIG5V.n11295 ASIG5V.n11294 0.019716
R56521 ASIG5V.n11304 ASIG5V.n10003 0.019716
R56522 ASIG5V.n11304 ASIG5V.n11303 0.019716
R56523 ASIG5V.n11306 ASIG5V.n10002 0.019716
R56524 ASIG5V.n11307 ASIG5V.n11306 0.019716
R56525 ASIG5V.n11316 ASIG5V.n10001 0.019716
R56526 ASIG5V.n11316 ASIG5V.n11315 0.019716
R56527 ASIG5V.n11318 ASIG5V.n10000 0.019716
R56528 ASIG5V.n11319 ASIG5V.n11318 0.019716
R56529 ASIG5V.n11328 ASIG5V.n9999 0.019716
R56530 ASIG5V.n11328 ASIG5V.n11327 0.019716
R56531 ASIG5V.n11330 ASIG5V.n9998 0.019716
R56532 ASIG5V.n11331 ASIG5V.n11330 0.019716
R56533 ASIG5V.n11340 ASIG5V.n9997 0.019716
R56534 ASIG5V.n11340 ASIG5V.n11339 0.019716
R56535 ASIG5V.n11342 ASIG5V.n9996 0.019716
R56536 ASIG5V.n11343 ASIG5V.n11342 0.019716
R56537 ASIG5V.n11352 ASIG5V.n9995 0.019716
R56538 ASIG5V.n11352 ASIG5V.n11351 0.019716
R56539 ASIG5V.n11354 ASIG5V.n9994 0.019716
R56540 ASIG5V.n11355 ASIG5V.n11354 0.019716
R56541 ASIG5V.n11364 ASIG5V.n9993 0.019716
R56542 ASIG5V.n11364 ASIG5V.n11363 0.019716
R56543 ASIG5V.n11366 ASIG5V.n9992 0.019716
R56544 ASIG5V.n11367 ASIG5V.n11366 0.019716
R56545 ASIG5V.n11376 ASIG5V.n9991 0.019716
R56546 ASIG5V.n11376 ASIG5V.n11375 0.019716
R56547 ASIG5V.n11378 ASIG5V.n9990 0.019716
R56548 ASIG5V.n11379 ASIG5V.n11378 0.019716
R56549 ASIG5V.n11388 ASIG5V.n9989 0.019716
R56550 ASIG5V.n11388 ASIG5V.n11387 0.019716
R56551 ASIG5V.n11390 ASIG5V.n9988 0.019716
R56552 ASIG5V.n11391 ASIG5V.n11390 0.019716
R56553 ASIG5V.n11400 ASIG5V.n9987 0.019716
R56554 ASIG5V.n11400 ASIG5V.n11399 0.019716
R56555 ASIG5V.n11402 ASIG5V.n9986 0.019716
R56556 ASIG5V.n11403 ASIG5V.n11402 0.019716
R56557 ASIG5V.n11412 ASIG5V.n9985 0.019716
R56558 ASIG5V.n11412 ASIG5V.n11411 0.019716
R56559 ASIG5V.n11414 ASIG5V.n9984 0.019716
R56560 ASIG5V.n11415 ASIG5V.n11414 0.019716
R56561 ASIG5V.n11424 ASIG5V.n9983 0.019716
R56562 ASIG5V.n11424 ASIG5V.n11423 0.019716
R56563 ASIG5V.n11426 ASIG5V.n9982 0.019716
R56564 ASIG5V.n11427 ASIG5V.n11426 0.019716
R56565 ASIG5V.n11436 ASIG5V.n9981 0.019716
R56566 ASIG5V.n11436 ASIG5V.n11435 0.019716
R56567 ASIG5V.n11438 ASIG5V.n9980 0.019716
R56568 ASIG5V.n11439 ASIG5V.n11438 0.019716
R56569 ASIG5V.n11448 ASIG5V.n9979 0.019716
R56570 ASIG5V.n11448 ASIG5V.n11447 0.019716
R56571 ASIG5V.n11450 ASIG5V.n9978 0.019716
R56572 ASIG5V.n11451 ASIG5V.n11450 0.019716
R56573 ASIG5V.n11460 ASIG5V.n9977 0.019716
R56574 ASIG5V.n11460 ASIG5V.n11459 0.019716
R56575 ASIG5V.n11462 ASIG5V.n9976 0.019716
R56576 ASIG5V.n11463 ASIG5V.n11462 0.019716
R56577 ASIG5V.n11472 ASIG5V.n9975 0.019716
R56578 ASIG5V.n11472 ASIG5V.n11471 0.019716
R56579 ASIG5V.n11474 ASIG5V.n9974 0.019716
R56580 ASIG5V.n11475 ASIG5V.n11474 0.019716
R56581 ASIG5V.n11484 ASIG5V.n11483 0.019716
R56582 ASIG5V.n2999 ASIG5V.n2955 0.019716
R56583 ASIG5V.n3000 ASIG5V.n2954 0.019716
R56584 ASIG5V.n11510 ASIG5V.n2953 0.019716
R56585 ASIG5V.n11510 ASIG5V.n11509 0.019716
R56586 ASIG5V.n11512 ASIG5V.n2952 0.019716
R56587 ASIG5V.n11513 ASIG5V.n11512 0.019716
R56588 ASIG5V.n11522 ASIG5V.n2951 0.019716
R56589 ASIG5V.n11522 ASIG5V.n11521 0.019716
R56590 ASIG5V.n11524 ASIG5V.n2950 0.019716
R56591 ASIG5V.n11525 ASIG5V.n11524 0.019716
R56592 ASIG5V.n11534 ASIG5V.n2949 0.019716
R56593 ASIG5V.n11534 ASIG5V.n11533 0.019716
R56594 ASIG5V.n11536 ASIG5V.n2948 0.019716
R56595 ASIG5V.n11537 ASIG5V.n11536 0.019716
R56596 ASIG5V.n11546 ASIG5V.n2947 0.019716
R56597 ASIG5V.n11546 ASIG5V.n11545 0.019716
R56598 ASIG5V.n11548 ASIG5V.n2946 0.019716
R56599 ASIG5V.n11549 ASIG5V.n11548 0.019716
R56600 ASIG5V.n11558 ASIG5V.n2945 0.019716
R56601 ASIG5V.n11558 ASIG5V.n11557 0.019716
R56602 ASIG5V.n11560 ASIG5V.n2944 0.019716
R56603 ASIG5V.n11561 ASIG5V.n11560 0.019716
R56604 ASIG5V.n11570 ASIG5V.n2943 0.019716
R56605 ASIG5V.n11570 ASIG5V.n11569 0.019716
R56606 ASIG5V.n11572 ASIG5V.n2942 0.019716
R56607 ASIG5V.n11573 ASIG5V.n11572 0.019716
R56608 ASIG5V.n11582 ASIG5V.n2941 0.019716
R56609 ASIG5V.n11582 ASIG5V.n11581 0.019716
R56610 ASIG5V.n11584 ASIG5V.n2940 0.019716
R56611 ASIG5V.n11585 ASIG5V.n11584 0.019716
R56612 ASIG5V.n11594 ASIG5V.n2939 0.019716
R56613 ASIG5V.n11594 ASIG5V.n11593 0.019716
R56614 ASIG5V.n11596 ASIG5V.n2938 0.019716
R56615 ASIG5V.n11597 ASIG5V.n11596 0.019716
R56616 ASIG5V.n11606 ASIG5V.n2937 0.019716
R56617 ASIG5V.n11606 ASIG5V.n11605 0.019716
R56618 ASIG5V.n11608 ASIG5V.n2936 0.019716
R56619 ASIG5V.n11609 ASIG5V.n11608 0.019716
R56620 ASIG5V.n11618 ASIG5V.n2935 0.019716
R56621 ASIG5V.n11618 ASIG5V.n11617 0.019716
R56622 ASIG5V.n11620 ASIG5V.n2934 0.019716
R56623 ASIG5V.n11621 ASIG5V.n11620 0.019716
R56624 ASIG5V.n11630 ASIG5V.n2933 0.019716
R56625 ASIG5V.n11630 ASIG5V.n11629 0.019716
R56626 ASIG5V.n11632 ASIG5V.n2932 0.019716
R56627 ASIG5V.n11633 ASIG5V.n11632 0.019716
R56628 ASIG5V.n11642 ASIG5V.n2931 0.019716
R56629 ASIG5V.n11642 ASIG5V.n11641 0.019716
R56630 ASIG5V.n11644 ASIG5V.n2930 0.019716
R56631 ASIG5V.n11645 ASIG5V.n11644 0.019716
R56632 ASIG5V.n11654 ASIG5V.n2929 0.019716
R56633 ASIG5V.n11654 ASIG5V.n11653 0.019716
R56634 ASIG5V.n11656 ASIG5V.n2928 0.019716
R56635 ASIG5V.n11657 ASIG5V.n11656 0.019716
R56636 ASIG5V.n11666 ASIG5V.n2927 0.019716
R56637 ASIG5V.n11666 ASIG5V.n11665 0.019716
R56638 ASIG5V.n11668 ASIG5V.n2926 0.019716
R56639 ASIG5V.n11669 ASIG5V.n11668 0.019716
R56640 ASIG5V.n11678 ASIG5V.n2925 0.019716
R56641 ASIG5V.n11678 ASIG5V.n11677 0.019716
R56642 ASIG5V.n11680 ASIG5V.n2924 0.019716
R56643 ASIG5V.n11681 ASIG5V.n11680 0.019716
R56644 ASIG5V.n11690 ASIG5V.n2923 0.019716
R56645 ASIG5V.n11690 ASIG5V.n11689 0.019716
R56646 ASIG5V.n11692 ASIG5V.n2922 0.019716
R56647 ASIG5V.n11693 ASIG5V.n11692 0.019716
R56648 ASIG5V.n11702 ASIG5V.n2921 0.019716
R56649 ASIG5V.n11702 ASIG5V.n11701 0.019716
R56650 ASIG5V.n11704 ASIG5V.n2920 0.019716
R56651 ASIG5V.n11705 ASIG5V.n11704 0.019716
R56652 ASIG5V.n11714 ASIG5V.n2919 0.019716
R56653 ASIG5V.n11714 ASIG5V.n11713 0.019716
R56654 ASIG5V.n11716 ASIG5V.n2918 0.019716
R56655 ASIG5V.n11717 ASIG5V.n11716 0.019716
R56656 ASIG5V.n11726 ASIG5V.n2917 0.019716
R56657 ASIG5V.n11726 ASIG5V.n11725 0.019716
R56658 ASIG5V.n11728 ASIG5V.n2916 0.019716
R56659 ASIG5V.n11729 ASIG5V.n11728 0.019716
R56660 ASIG5V.n11738 ASIG5V.n2915 0.019716
R56661 ASIG5V.n11738 ASIG5V.n11737 0.019716
R56662 ASIG5V.n11740 ASIG5V.n2914 0.019716
R56663 ASIG5V.n11741 ASIG5V.n11740 0.019716
R56664 ASIG5V.n11750 ASIG5V.n11749 0.019716
R56665 ASIG5V.n2658 ASIG5V.n2611 0.019716
R56666 ASIG5V.n2659 ASIG5V.n2610 0.019716
R56667 ASIG5V.n2666 ASIG5V.n2609 0.019716
R56668 ASIG5V.n2666 ASIG5V.n2665 0.019716
R56669 ASIG5V.n2668 ASIG5V.n2608 0.019716
R56670 ASIG5V.n2669 ASIG5V.n2668 0.019716
R56671 ASIG5V.n2678 ASIG5V.n2607 0.019716
R56672 ASIG5V.n2678 ASIG5V.n2677 0.019716
R56673 ASIG5V.n2680 ASIG5V.n2606 0.019716
R56674 ASIG5V.n2681 ASIG5V.n2680 0.019716
R56675 ASIG5V.n2690 ASIG5V.n2605 0.019716
R56676 ASIG5V.n2690 ASIG5V.n2689 0.019716
R56677 ASIG5V.n2692 ASIG5V.n2604 0.019716
R56678 ASIG5V.n2693 ASIG5V.n2692 0.019716
R56679 ASIG5V.n2702 ASIG5V.n2603 0.019716
R56680 ASIG5V.n2702 ASIG5V.n2701 0.019716
R56681 ASIG5V.n2704 ASIG5V.n2602 0.019716
R56682 ASIG5V.n2705 ASIG5V.n2704 0.019716
R56683 ASIG5V.n2714 ASIG5V.n2601 0.019716
R56684 ASIG5V.n2714 ASIG5V.n2713 0.019716
R56685 ASIG5V.n2716 ASIG5V.n2600 0.019716
R56686 ASIG5V.n2717 ASIG5V.n2716 0.019716
R56687 ASIG5V.n2726 ASIG5V.n2599 0.019716
R56688 ASIG5V.n2726 ASIG5V.n2725 0.019716
R56689 ASIG5V.n2728 ASIG5V.n2598 0.019716
R56690 ASIG5V.n2729 ASIG5V.n2728 0.019716
R56691 ASIG5V.n2738 ASIG5V.n2597 0.019716
R56692 ASIG5V.n2738 ASIG5V.n2737 0.019716
R56693 ASIG5V.n2740 ASIG5V.n2596 0.019716
R56694 ASIG5V.n2741 ASIG5V.n2740 0.019716
R56695 ASIG5V.n2750 ASIG5V.n2595 0.019716
R56696 ASIG5V.n2750 ASIG5V.n2749 0.019716
R56697 ASIG5V.n2752 ASIG5V.n2594 0.019716
R56698 ASIG5V.n2753 ASIG5V.n2752 0.019716
R56699 ASIG5V.n2762 ASIG5V.n2593 0.019716
R56700 ASIG5V.n2762 ASIG5V.n2761 0.019716
R56701 ASIG5V.n2764 ASIG5V.n2592 0.019716
R56702 ASIG5V.n2765 ASIG5V.n2764 0.019716
R56703 ASIG5V.n2774 ASIG5V.n2591 0.019716
R56704 ASIG5V.n2774 ASIG5V.n2773 0.019716
R56705 ASIG5V.n2776 ASIG5V.n2590 0.019716
R56706 ASIG5V.n2777 ASIG5V.n2776 0.019716
R56707 ASIG5V.n2786 ASIG5V.n2589 0.019716
R56708 ASIG5V.n2786 ASIG5V.n2785 0.019716
R56709 ASIG5V.n2788 ASIG5V.n2588 0.019716
R56710 ASIG5V.n2789 ASIG5V.n2788 0.019716
R56711 ASIG5V.n2798 ASIG5V.n2587 0.019716
R56712 ASIG5V.n2798 ASIG5V.n2797 0.019716
R56713 ASIG5V.n2800 ASIG5V.n2586 0.019716
R56714 ASIG5V.n2801 ASIG5V.n2800 0.019716
R56715 ASIG5V.n2810 ASIG5V.n2585 0.019716
R56716 ASIG5V.n2810 ASIG5V.n2809 0.019716
R56717 ASIG5V.n2812 ASIG5V.n2584 0.019716
R56718 ASIG5V.n2813 ASIG5V.n2812 0.019716
R56719 ASIG5V.n2822 ASIG5V.n2583 0.019716
R56720 ASIG5V.n2822 ASIG5V.n2821 0.019716
R56721 ASIG5V.n2824 ASIG5V.n2582 0.019716
R56722 ASIG5V.n2825 ASIG5V.n2824 0.019716
R56723 ASIG5V.n2834 ASIG5V.n2581 0.019716
R56724 ASIG5V.n2834 ASIG5V.n2833 0.019716
R56725 ASIG5V.n2836 ASIG5V.n2580 0.019716
R56726 ASIG5V.n2837 ASIG5V.n2836 0.019716
R56727 ASIG5V.n2846 ASIG5V.n2579 0.019716
R56728 ASIG5V.n2846 ASIG5V.n2845 0.019716
R56729 ASIG5V.n2848 ASIG5V.n2578 0.019716
R56730 ASIG5V.n2849 ASIG5V.n2848 0.019716
R56731 ASIG5V.n2858 ASIG5V.n2577 0.019716
R56732 ASIG5V.n2858 ASIG5V.n2857 0.019716
R56733 ASIG5V.n2860 ASIG5V.n2576 0.019716
R56734 ASIG5V.n2861 ASIG5V.n2860 0.019716
R56735 ASIG5V.n2870 ASIG5V.n2575 0.019716
R56736 ASIG5V.n2870 ASIG5V.n2869 0.019716
R56737 ASIG5V.n2872 ASIG5V.n2574 0.019716
R56738 ASIG5V.n2873 ASIG5V.n2872 0.019716
R56739 ASIG5V.n2882 ASIG5V.n2573 0.019716
R56740 ASIG5V.n2882 ASIG5V.n2881 0.019716
R56741 ASIG5V.n2884 ASIG5V.n2572 0.019716
R56742 ASIG5V.n2885 ASIG5V.n2884 0.019716
R56743 ASIG5V.n2894 ASIG5V.n2571 0.019716
R56744 ASIG5V.n2894 ASIG5V.n2893 0.019716
R56745 ASIG5V.n2896 ASIG5V.n2570 0.019716
R56746 ASIG5V.n2897 ASIG5V.n2896 0.019716
R56747 ASIG5V.n11770 ASIG5V.n11769 0.019716
R56748 ASIG5V.n2306 ASIG5V.n2263 0.019716
R56749 ASIG5V.n2307 ASIG5V.n2262 0.019716
R56750 ASIG5V.n2314 ASIG5V.n2261 0.019716
R56751 ASIG5V.n2314 ASIG5V.n2313 0.019716
R56752 ASIG5V.n2316 ASIG5V.n2260 0.019716
R56753 ASIG5V.n2317 ASIG5V.n2316 0.019716
R56754 ASIG5V.n2326 ASIG5V.n2259 0.019716
R56755 ASIG5V.n2326 ASIG5V.n2325 0.019716
R56756 ASIG5V.n2328 ASIG5V.n2258 0.019716
R56757 ASIG5V.n2329 ASIG5V.n2328 0.019716
R56758 ASIG5V.n2338 ASIG5V.n2257 0.019716
R56759 ASIG5V.n2338 ASIG5V.n2337 0.019716
R56760 ASIG5V.n2340 ASIG5V.n2256 0.019716
R56761 ASIG5V.n2341 ASIG5V.n2340 0.019716
R56762 ASIG5V.n2350 ASIG5V.n2255 0.019716
R56763 ASIG5V.n2350 ASIG5V.n2349 0.019716
R56764 ASIG5V.n2352 ASIG5V.n2254 0.019716
R56765 ASIG5V.n2353 ASIG5V.n2352 0.019716
R56766 ASIG5V.n2362 ASIG5V.n2253 0.019716
R56767 ASIG5V.n2362 ASIG5V.n2361 0.019716
R56768 ASIG5V.n2364 ASIG5V.n2252 0.019716
R56769 ASIG5V.n2365 ASIG5V.n2364 0.019716
R56770 ASIG5V.n2374 ASIG5V.n2251 0.019716
R56771 ASIG5V.n2374 ASIG5V.n2373 0.019716
R56772 ASIG5V.n2376 ASIG5V.n2250 0.019716
R56773 ASIG5V.n2377 ASIG5V.n2376 0.019716
R56774 ASIG5V.n2386 ASIG5V.n2249 0.019716
R56775 ASIG5V.n2386 ASIG5V.n2385 0.019716
R56776 ASIG5V.n2388 ASIG5V.n2248 0.019716
R56777 ASIG5V.n2389 ASIG5V.n2388 0.019716
R56778 ASIG5V.n2398 ASIG5V.n2247 0.019716
R56779 ASIG5V.n2398 ASIG5V.n2397 0.019716
R56780 ASIG5V.n2400 ASIG5V.n2246 0.019716
R56781 ASIG5V.n2401 ASIG5V.n2400 0.019716
R56782 ASIG5V.n2410 ASIG5V.n2245 0.019716
R56783 ASIG5V.n2410 ASIG5V.n2409 0.019716
R56784 ASIG5V.n2412 ASIG5V.n2244 0.019716
R56785 ASIG5V.n2413 ASIG5V.n2412 0.019716
R56786 ASIG5V.n2422 ASIG5V.n2243 0.019716
R56787 ASIG5V.n2422 ASIG5V.n2421 0.019716
R56788 ASIG5V.n2424 ASIG5V.n2242 0.019716
R56789 ASIG5V.n2425 ASIG5V.n2424 0.019716
R56790 ASIG5V.n2434 ASIG5V.n2241 0.019716
R56791 ASIG5V.n2434 ASIG5V.n2433 0.019716
R56792 ASIG5V.n2436 ASIG5V.n2240 0.019716
R56793 ASIG5V.n2437 ASIG5V.n2436 0.019716
R56794 ASIG5V.n2446 ASIG5V.n2239 0.019716
R56795 ASIG5V.n2446 ASIG5V.n2445 0.019716
R56796 ASIG5V.n2448 ASIG5V.n2238 0.019716
R56797 ASIG5V.n2449 ASIG5V.n2448 0.019716
R56798 ASIG5V.n2458 ASIG5V.n2237 0.019716
R56799 ASIG5V.n2458 ASIG5V.n2457 0.019716
R56800 ASIG5V.n2460 ASIG5V.n2236 0.019716
R56801 ASIG5V.n2461 ASIG5V.n2460 0.019716
R56802 ASIG5V.n2470 ASIG5V.n2235 0.019716
R56803 ASIG5V.n2470 ASIG5V.n2469 0.019716
R56804 ASIG5V.n2472 ASIG5V.n2234 0.019716
R56805 ASIG5V.n2473 ASIG5V.n2472 0.019716
R56806 ASIG5V.n2482 ASIG5V.n2233 0.019716
R56807 ASIG5V.n2482 ASIG5V.n2481 0.019716
R56808 ASIG5V.n2484 ASIG5V.n2232 0.019716
R56809 ASIG5V.n2485 ASIG5V.n2484 0.019716
R56810 ASIG5V.n2494 ASIG5V.n2231 0.019716
R56811 ASIG5V.n2494 ASIG5V.n2493 0.019716
R56812 ASIG5V.n2496 ASIG5V.n2230 0.019716
R56813 ASIG5V.n2497 ASIG5V.n2496 0.019716
R56814 ASIG5V.n2506 ASIG5V.n2229 0.019716
R56815 ASIG5V.n2506 ASIG5V.n2505 0.019716
R56816 ASIG5V.n2508 ASIG5V.n2228 0.019716
R56817 ASIG5V.n2509 ASIG5V.n2508 0.019716
R56818 ASIG5V.n2518 ASIG5V.n2227 0.019716
R56819 ASIG5V.n2518 ASIG5V.n2517 0.019716
R56820 ASIG5V.n2520 ASIG5V.n2226 0.019716
R56821 ASIG5V.n2521 ASIG5V.n2520 0.019716
R56822 ASIG5V.n2530 ASIG5V.n2225 0.019716
R56823 ASIG5V.n2530 ASIG5V.n2529 0.019716
R56824 ASIG5V.n2532 ASIG5V.n2224 0.019716
R56825 ASIG5V.n2533 ASIG5V.n2532 0.019716
R56826 ASIG5V.n2542 ASIG5V.n2223 0.019716
R56827 ASIG5V.n2542 ASIG5V.n2541 0.019716
R56828 ASIG5V.n2544 ASIG5V.n2222 0.019716
R56829 ASIG5V.n2545 ASIG5V.n2544 0.019716
R56830 ASIG5V.n2554 ASIG5V.n2553 0.019716
R56831 ASIG5V.n1949 ASIG5V.n1906 0.019716
R56832 ASIG5V.n1950 ASIG5V.n1905 0.019716
R56833 ASIG5V.n1957 ASIG5V.n1904 0.019716
R56834 ASIG5V.n1957 ASIG5V.n1956 0.019716
R56835 ASIG5V.n1959 ASIG5V.n1903 0.019716
R56836 ASIG5V.n1960 ASIG5V.n1959 0.019716
R56837 ASIG5V.n1969 ASIG5V.n1902 0.019716
R56838 ASIG5V.n1969 ASIG5V.n1968 0.019716
R56839 ASIG5V.n1971 ASIG5V.n1901 0.019716
R56840 ASIG5V.n1972 ASIG5V.n1971 0.019716
R56841 ASIG5V.n1981 ASIG5V.n1900 0.019716
R56842 ASIG5V.n1981 ASIG5V.n1980 0.019716
R56843 ASIG5V.n1983 ASIG5V.n1899 0.019716
R56844 ASIG5V.n1984 ASIG5V.n1983 0.019716
R56845 ASIG5V.n1993 ASIG5V.n1898 0.019716
R56846 ASIG5V.n1993 ASIG5V.n1992 0.019716
R56847 ASIG5V.n1995 ASIG5V.n1897 0.019716
R56848 ASIG5V.n1996 ASIG5V.n1995 0.019716
R56849 ASIG5V.n2005 ASIG5V.n1896 0.019716
R56850 ASIG5V.n2005 ASIG5V.n2004 0.019716
R56851 ASIG5V.n2007 ASIG5V.n1895 0.019716
R56852 ASIG5V.n2008 ASIG5V.n2007 0.019716
R56853 ASIG5V.n2017 ASIG5V.n1894 0.019716
R56854 ASIG5V.n2017 ASIG5V.n2016 0.019716
R56855 ASIG5V.n2019 ASIG5V.n1893 0.019716
R56856 ASIG5V.n2020 ASIG5V.n2019 0.019716
R56857 ASIG5V.n2029 ASIG5V.n1892 0.019716
R56858 ASIG5V.n2029 ASIG5V.n2028 0.019716
R56859 ASIG5V.n2031 ASIG5V.n1891 0.019716
R56860 ASIG5V.n2032 ASIG5V.n2031 0.019716
R56861 ASIG5V.n2041 ASIG5V.n1890 0.019716
R56862 ASIG5V.n2041 ASIG5V.n2040 0.019716
R56863 ASIG5V.n2043 ASIG5V.n1889 0.019716
R56864 ASIG5V.n2044 ASIG5V.n2043 0.019716
R56865 ASIG5V.n2053 ASIG5V.n1888 0.019716
R56866 ASIG5V.n2053 ASIG5V.n2052 0.019716
R56867 ASIG5V.n2055 ASIG5V.n1887 0.019716
R56868 ASIG5V.n2056 ASIG5V.n2055 0.019716
R56869 ASIG5V.n2065 ASIG5V.n1886 0.019716
R56870 ASIG5V.n2065 ASIG5V.n2064 0.019716
R56871 ASIG5V.n2067 ASIG5V.n1885 0.019716
R56872 ASIG5V.n2068 ASIG5V.n2067 0.019716
R56873 ASIG5V.n2077 ASIG5V.n1884 0.019716
R56874 ASIG5V.n2077 ASIG5V.n2076 0.019716
R56875 ASIG5V.n2079 ASIG5V.n1883 0.019716
R56876 ASIG5V.n2080 ASIG5V.n2079 0.019716
R56877 ASIG5V.n2089 ASIG5V.n1882 0.019716
R56878 ASIG5V.n2089 ASIG5V.n2088 0.019716
R56879 ASIG5V.n2091 ASIG5V.n1881 0.019716
R56880 ASIG5V.n2092 ASIG5V.n2091 0.019716
R56881 ASIG5V.n2101 ASIG5V.n1880 0.019716
R56882 ASIG5V.n2101 ASIG5V.n2100 0.019716
R56883 ASIG5V.n2103 ASIG5V.n1879 0.019716
R56884 ASIG5V.n2104 ASIG5V.n2103 0.019716
R56885 ASIG5V.n2113 ASIG5V.n1878 0.019716
R56886 ASIG5V.n2113 ASIG5V.n2112 0.019716
R56887 ASIG5V.n2115 ASIG5V.n1877 0.019716
R56888 ASIG5V.n2116 ASIG5V.n2115 0.019716
R56889 ASIG5V.n2125 ASIG5V.n1876 0.019716
R56890 ASIG5V.n2125 ASIG5V.n2124 0.019716
R56891 ASIG5V.n2127 ASIG5V.n1875 0.019716
R56892 ASIG5V.n2128 ASIG5V.n2127 0.019716
R56893 ASIG5V.n2137 ASIG5V.n1874 0.019716
R56894 ASIG5V.n2137 ASIG5V.n2136 0.019716
R56895 ASIG5V.n2139 ASIG5V.n1873 0.019716
R56896 ASIG5V.n2140 ASIG5V.n2139 0.019716
R56897 ASIG5V.n2149 ASIG5V.n1872 0.019716
R56898 ASIG5V.n2149 ASIG5V.n2148 0.019716
R56899 ASIG5V.n2151 ASIG5V.n1871 0.019716
R56900 ASIG5V.n2152 ASIG5V.n2151 0.019716
R56901 ASIG5V.n2161 ASIG5V.n1870 0.019716
R56902 ASIG5V.n2161 ASIG5V.n2160 0.019716
R56903 ASIG5V.n2163 ASIG5V.n1869 0.019716
R56904 ASIG5V.n2164 ASIG5V.n2163 0.019716
R56905 ASIG5V.n2173 ASIG5V.n1868 0.019716
R56906 ASIG5V.n2173 ASIG5V.n2172 0.019716
R56907 ASIG5V.n2175 ASIG5V.n1867 0.019716
R56908 ASIG5V.n2176 ASIG5V.n2175 0.019716
R56909 ASIG5V.n2185 ASIG5V.n1866 0.019716
R56910 ASIG5V.n2185 ASIG5V.n2184 0.019716
R56911 ASIG5V.n2187 ASIG5V.n1865 0.019716
R56912 ASIG5V.n2188 ASIG5V.n2187 0.019716
R56913 ASIG5V.n2197 ASIG5V.n2196 0.019716
R56914 ASIG5V.n11996 ASIG5V.n11995 0.019716
R56915 ASIG5V.n1762 ASIG5V.n1718 0.019716
R56916 ASIG5V.n11812 ASIG5V.n1761 0.019716
R56917 ASIG5V.n11812 ASIG5V.n1716 0.019716
R56918 ASIG5V.n11816 ASIG5V.n1760 0.019716
R56919 ASIG5V.n11816 ASIG5V.n1715 0.019716
R56920 ASIG5V.n11821 ASIG5V.n1759 0.019716
R56921 ASIG5V.n11821 ASIG5V.n1714 0.019716
R56922 ASIG5V.n11825 ASIG5V.n1758 0.019716
R56923 ASIG5V.n11825 ASIG5V.n1713 0.019716
R56924 ASIG5V.n11830 ASIG5V.n1757 0.019716
R56925 ASIG5V.n11830 ASIG5V.n1712 0.019716
R56926 ASIG5V.n11834 ASIG5V.n1756 0.019716
R56927 ASIG5V.n11834 ASIG5V.n1711 0.019716
R56928 ASIG5V.n11839 ASIG5V.n1755 0.019716
R56929 ASIG5V.n11839 ASIG5V.n1710 0.019716
R56930 ASIG5V.n11843 ASIG5V.n1754 0.019716
R56931 ASIG5V.n11843 ASIG5V.n1709 0.019716
R56932 ASIG5V.n11848 ASIG5V.n1753 0.019716
R56933 ASIG5V.n11848 ASIG5V.n1708 0.019716
R56934 ASIG5V.n11852 ASIG5V.n1752 0.019716
R56935 ASIG5V.n11852 ASIG5V.n1707 0.019716
R56936 ASIG5V.n11857 ASIG5V.n1751 0.019716
R56937 ASIG5V.n11857 ASIG5V.n1706 0.019716
R56938 ASIG5V.n11861 ASIG5V.n1750 0.019716
R56939 ASIG5V.n11861 ASIG5V.n1705 0.019716
R56940 ASIG5V.n11866 ASIG5V.n1749 0.019716
R56941 ASIG5V.n11866 ASIG5V.n1704 0.019716
R56942 ASIG5V.n11870 ASIG5V.n1748 0.019716
R56943 ASIG5V.n11870 ASIG5V.n1703 0.019716
R56944 ASIG5V.n11875 ASIG5V.n1747 0.019716
R56945 ASIG5V.n11875 ASIG5V.n1702 0.019716
R56946 ASIG5V.n11879 ASIG5V.n1746 0.019716
R56947 ASIG5V.n11879 ASIG5V.n1701 0.019716
R56948 ASIG5V.n11884 ASIG5V.n1745 0.019716
R56949 ASIG5V.n11884 ASIG5V.n1700 0.019716
R56950 ASIG5V.n11888 ASIG5V.n1744 0.019716
R56951 ASIG5V.n11888 ASIG5V.n1699 0.019716
R56952 ASIG5V.n11893 ASIG5V.n1743 0.019716
R56953 ASIG5V.n11893 ASIG5V.n1698 0.019716
R56954 ASIG5V.n11897 ASIG5V.n1742 0.019716
R56955 ASIG5V.n11897 ASIG5V.n1697 0.019716
R56956 ASIG5V.n11902 ASIG5V.n1741 0.019716
R56957 ASIG5V.n11902 ASIG5V.n1696 0.019716
R56958 ASIG5V.n11906 ASIG5V.n1740 0.019716
R56959 ASIG5V.n11906 ASIG5V.n1695 0.019716
R56960 ASIG5V.n11911 ASIG5V.n1739 0.019716
R56961 ASIG5V.n11911 ASIG5V.n1694 0.019716
R56962 ASIG5V.n11915 ASIG5V.n1738 0.019716
R56963 ASIG5V.n11915 ASIG5V.n1693 0.019716
R56964 ASIG5V.n11920 ASIG5V.n1737 0.019716
R56965 ASIG5V.n11920 ASIG5V.n1692 0.019716
R56966 ASIG5V.n11924 ASIG5V.n1736 0.019716
R56967 ASIG5V.n11924 ASIG5V.n1691 0.019716
R56968 ASIG5V.n11929 ASIG5V.n1735 0.019716
R56969 ASIG5V.n11929 ASIG5V.n1690 0.019716
R56970 ASIG5V.n11933 ASIG5V.n1734 0.019716
R56971 ASIG5V.n11933 ASIG5V.n1689 0.019716
R56972 ASIG5V.n11938 ASIG5V.n1733 0.019716
R56973 ASIG5V.n11938 ASIG5V.n1688 0.019716
R56974 ASIG5V.n11942 ASIG5V.n1732 0.019716
R56975 ASIG5V.n11942 ASIG5V.n1687 0.019716
R56976 ASIG5V.n11947 ASIG5V.n1731 0.019716
R56977 ASIG5V.n11947 ASIG5V.n1686 0.019716
R56978 ASIG5V.n11951 ASIG5V.n1730 0.019716
R56979 ASIG5V.n11951 ASIG5V.n1685 0.019716
R56980 ASIG5V.n11956 ASIG5V.n1729 0.019716
R56981 ASIG5V.n11956 ASIG5V.n1684 0.019716
R56982 ASIG5V.n11960 ASIG5V.n1728 0.019716
R56983 ASIG5V.n11960 ASIG5V.n1683 0.019716
R56984 ASIG5V.n11965 ASIG5V.n1727 0.019716
R56985 ASIG5V.n11965 ASIG5V.n1682 0.019716
R56986 ASIG5V.n11969 ASIG5V.n1726 0.019716
R56987 ASIG5V.n11969 ASIG5V.n1681 0.019716
R56988 ASIG5V.n11974 ASIG5V.n1725 0.019716
R56989 ASIG5V.n11974 ASIG5V.n1680 0.019716
R56990 ASIG5V.n11978 ASIG5V.n1724 0.019716
R56991 ASIG5V.n11978 ASIG5V.n1679 0.019716
R56992 ASIG5V.n11983 ASIG5V.n1723 0.019716
R56993 ASIG5V.n11983 ASIG5V.n1678 0.019716
R56994 ASIG5V.n11987 ASIG5V.n1722 0.019716
R56995 ASIG5V.n11987 ASIG5V.n1677 0.019716
R56996 ASIG5V.n11993 ASIG5V.n1676 0.019716
R56997 ASIG5V.n12010 ASIG5V.n12009 0.019716
R56998 ASIG5V.n1414 ASIG5V.n1371 0.019716
R56999 ASIG5V.n1484 ASIG5V.n1413 0.019716
R57000 ASIG5V.n1484 ASIG5V.n1369 0.019716
R57001 ASIG5V.n1488 ASIG5V.n1412 0.019716
R57002 ASIG5V.n1488 ASIG5V.n1368 0.019716
R57003 ASIG5V.n1493 ASIG5V.n1411 0.019716
R57004 ASIG5V.n1493 ASIG5V.n1367 0.019716
R57005 ASIG5V.n1497 ASIG5V.n1410 0.019716
R57006 ASIG5V.n1497 ASIG5V.n1366 0.019716
R57007 ASIG5V.n1502 ASIG5V.n1409 0.019716
R57008 ASIG5V.n1502 ASIG5V.n1365 0.019716
R57009 ASIG5V.n1506 ASIG5V.n1408 0.019716
R57010 ASIG5V.n1506 ASIG5V.n1364 0.019716
R57011 ASIG5V.n1511 ASIG5V.n1407 0.019716
R57012 ASIG5V.n1511 ASIG5V.n1363 0.019716
R57013 ASIG5V.n1515 ASIG5V.n1406 0.019716
R57014 ASIG5V.n1515 ASIG5V.n1362 0.019716
R57015 ASIG5V.n1520 ASIG5V.n1405 0.019716
R57016 ASIG5V.n1520 ASIG5V.n1361 0.019716
R57017 ASIG5V.n1524 ASIG5V.n1404 0.019716
R57018 ASIG5V.n1524 ASIG5V.n1360 0.019716
R57019 ASIG5V.n1529 ASIG5V.n1403 0.019716
R57020 ASIG5V.n1529 ASIG5V.n1359 0.019716
R57021 ASIG5V.n1533 ASIG5V.n1402 0.019716
R57022 ASIG5V.n1533 ASIG5V.n1358 0.019716
R57023 ASIG5V.n1538 ASIG5V.n1401 0.019716
R57024 ASIG5V.n1538 ASIG5V.n1357 0.019716
R57025 ASIG5V.n1542 ASIG5V.n1400 0.019716
R57026 ASIG5V.n1542 ASIG5V.n1356 0.019716
R57027 ASIG5V.n1547 ASIG5V.n1399 0.019716
R57028 ASIG5V.n1547 ASIG5V.n1355 0.019716
R57029 ASIG5V.n1551 ASIG5V.n1398 0.019716
R57030 ASIG5V.n1551 ASIG5V.n1354 0.019716
R57031 ASIG5V.n1556 ASIG5V.n1397 0.019716
R57032 ASIG5V.n1556 ASIG5V.n1353 0.019716
R57033 ASIG5V.n1560 ASIG5V.n1396 0.019716
R57034 ASIG5V.n1560 ASIG5V.n1352 0.019716
R57035 ASIG5V.n1565 ASIG5V.n1395 0.019716
R57036 ASIG5V.n1565 ASIG5V.n1351 0.019716
R57037 ASIG5V.n1569 ASIG5V.n1394 0.019716
R57038 ASIG5V.n1569 ASIG5V.n1350 0.019716
R57039 ASIG5V.n1574 ASIG5V.n1393 0.019716
R57040 ASIG5V.n1574 ASIG5V.n1349 0.019716
R57041 ASIG5V.n1578 ASIG5V.n1392 0.019716
R57042 ASIG5V.n1578 ASIG5V.n1348 0.019716
R57043 ASIG5V.n1583 ASIG5V.n1391 0.019716
R57044 ASIG5V.n1583 ASIG5V.n1347 0.019716
R57045 ASIG5V.n1587 ASIG5V.n1390 0.019716
R57046 ASIG5V.n1587 ASIG5V.n1346 0.019716
R57047 ASIG5V.n1592 ASIG5V.n1389 0.019716
R57048 ASIG5V.n1592 ASIG5V.n1345 0.019716
R57049 ASIG5V.n1596 ASIG5V.n1388 0.019716
R57050 ASIG5V.n1596 ASIG5V.n1344 0.019716
R57051 ASIG5V.n1601 ASIG5V.n1387 0.019716
R57052 ASIG5V.n1601 ASIG5V.n1343 0.019716
R57053 ASIG5V.n1605 ASIG5V.n1386 0.019716
R57054 ASIG5V.n1605 ASIG5V.n1342 0.019716
R57055 ASIG5V.n1610 ASIG5V.n1385 0.019716
R57056 ASIG5V.n1610 ASIG5V.n1341 0.019716
R57057 ASIG5V.n1614 ASIG5V.n1384 0.019716
R57058 ASIG5V.n1614 ASIG5V.n1340 0.019716
R57059 ASIG5V.n1619 ASIG5V.n1383 0.019716
R57060 ASIG5V.n1619 ASIG5V.n1339 0.019716
R57061 ASIG5V.n1623 ASIG5V.n1382 0.019716
R57062 ASIG5V.n1623 ASIG5V.n1338 0.019716
R57063 ASIG5V.n1628 ASIG5V.n1381 0.019716
R57064 ASIG5V.n1628 ASIG5V.n1337 0.019716
R57065 ASIG5V.n1632 ASIG5V.n1380 0.019716
R57066 ASIG5V.n1632 ASIG5V.n1336 0.019716
R57067 ASIG5V.n1637 ASIG5V.n1379 0.019716
R57068 ASIG5V.n1637 ASIG5V.n1335 0.019716
R57069 ASIG5V.n1641 ASIG5V.n1378 0.019716
R57070 ASIG5V.n1641 ASIG5V.n1334 0.019716
R57071 ASIG5V.n1646 ASIG5V.n1377 0.019716
R57072 ASIG5V.n1646 ASIG5V.n1333 0.019716
R57073 ASIG5V.n1650 ASIG5V.n1376 0.019716
R57074 ASIG5V.n1650 ASIG5V.n1332 0.019716
R57075 ASIG5V.n1655 ASIG5V.n1375 0.019716
R57076 ASIG5V.n1655 ASIG5V.n1331 0.019716
R57077 ASIG5V.n1659 ASIG5V.n1374 0.019716
R57078 ASIG5V.n1659 ASIG5V.n1330 0.019716
R57079 ASIG5V.n12007 ASIG5V.n1329 0.019716
R57080 ASIG5V.n1313 ASIG5V.n1268 0.019716
R57081 ASIG5V.n1314 ASIG5V.n1267 0.019716
R57082 ASIG5V.n12027 ASIG5V.n1266 0.019716
R57083 ASIG5V.n12027 ASIG5V.n12026 0.019716
R57084 ASIG5V.n12029 ASIG5V.n1265 0.019716
R57085 ASIG5V.n12030 ASIG5V.n12029 0.019716
R57086 ASIG5V.n12039 ASIG5V.n1264 0.019716
R57087 ASIG5V.n12039 ASIG5V.n12038 0.019716
R57088 ASIG5V.n12041 ASIG5V.n1263 0.019716
R57089 ASIG5V.n12042 ASIG5V.n12041 0.019716
R57090 ASIG5V.n12051 ASIG5V.n1262 0.019716
R57091 ASIG5V.n12051 ASIG5V.n12050 0.019716
R57092 ASIG5V.n12053 ASIG5V.n1261 0.019716
R57093 ASIG5V.n12054 ASIG5V.n12053 0.019716
R57094 ASIG5V.n12063 ASIG5V.n1260 0.019716
R57095 ASIG5V.n12063 ASIG5V.n12062 0.019716
R57096 ASIG5V.n12065 ASIG5V.n1259 0.019716
R57097 ASIG5V.n12066 ASIG5V.n12065 0.019716
R57098 ASIG5V.n12075 ASIG5V.n1258 0.019716
R57099 ASIG5V.n12075 ASIG5V.n12074 0.019716
R57100 ASIG5V.n12077 ASIG5V.n1257 0.019716
R57101 ASIG5V.n12078 ASIG5V.n12077 0.019716
R57102 ASIG5V.n12087 ASIG5V.n1256 0.019716
R57103 ASIG5V.n12087 ASIG5V.n12086 0.019716
R57104 ASIG5V.n12089 ASIG5V.n1255 0.019716
R57105 ASIG5V.n12090 ASIG5V.n12089 0.019716
R57106 ASIG5V.n12099 ASIG5V.n1254 0.019716
R57107 ASIG5V.n12099 ASIG5V.n12098 0.019716
R57108 ASIG5V.n12101 ASIG5V.n1253 0.019716
R57109 ASIG5V.n12102 ASIG5V.n12101 0.019716
R57110 ASIG5V.n12111 ASIG5V.n1252 0.019716
R57111 ASIG5V.n12111 ASIG5V.n12110 0.019716
R57112 ASIG5V.n12113 ASIG5V.n1251 0.019716
R57113 ASIG5V.n12114 ASIG5V.n12113 0.019716
R57114 ASIG5V.n12123 ASIG5V.n1250 0.019716
R57115 ASIG5V.n12123 ASIG5V.n12122 0.019716
R57116 ASIG5V.n12125 ASIG5V.n1249 0.019716
R57117 ASIG5V.n12126 ASIG5V.n12125 0.019716
R57118 ASIG5V.n12135 ASIG5V.n1248 0.019716
R57119 ASIG5V.n12135 ASIG5V.n12134 0.019716
R57120 ASIG5V.n12137 ASIG5V.n1247 0.019716
R57121 ASIG5V.n12138 ASIG5V.n12137 0.019716
R57122 ASIG5V.n12147 ASIG5V.n1246 0.019716
R57123 ASIG5V.n12147 ASIG5V.n12146 0.019716
R57124 ASIG5V.n12149 ASIG5V.n1245 0.019716
R57125 ASIG5V.n12150 ASIG5V.n12149 0.019716
R57126 ASIG5V.n12159 ASIG5V.n1244 0.019716
R57127 ASIG5V.n12159 ASIG5V.n12158 0.019716
R57128 ASIG5V.n12161 ASIG5V.n1243 0.019716
R57129 ASIG5V.n12162 ASIG5V.n12161 0.019716
R57130 ASIG5V.n12171 ASIG5V.n1242 0.019716
R57131 ASIG5V.n12171 ASIG5V.n12170 0.019716
R57132 ASIG5V.n12173 ASIG5V.n1241 0.019716
R57133 ASIG5V.n12174 ASIG5V.n12173 0.019716
R57134 ASIG5V.n12183 ASIG5V.n1240 0.019716
R57135 ASIG5V.n12183 ASIG5V.n12182 0.019716
R57136 ASIG5V.n12185 ASIG5V.n1239 0.019716
R57137 ASIG5V.n12186 ASIG5V.n12185 0.019716
R57138 ASIG5V.n12195 ASIG5V.n1238 0.019716
R57139 ASIG5V.n12195 ASIG5V.n12194 0.019716
R57140 ASIG5V.n12197 ASIG5V.n1237 0.019716
R57141 ASIG5V.n12198 ASIG5V.n12197 0.019716
R57142 ASIG5V.n12207 ASIG5V.n1236 0.019716
R57143 ASIG5V.n12207 ASIG5V.n12206 0.019716
R57144 ASIG5V.n12209 ASIG5V.n1235 0.019716
R57145 ASIG5V.n12210 ASIG5V.n12209 0.019716
R57146 ASIG5V.n12219 ASIG5V.n1234 0.019716
R57147 ASIG5V.n12219 ASIG5V.n12218 0.019716
R57148 ASIG5V.n12221 ASIG5V.n1233 0.019716
R57149 ASIG5V.n12222 ASIG5V.n12221 0.019716
R57150 ASIG5V.n12231 ASIG5V.n1232 0.019716
R57151 ASIG5V.n12231 ASIG5V.n12230 0.019716
R57152 ASIG5V.n12233 ASIG5V.n1231 0.019716
R57153 ASIG5V.n12234 ASIG5V.n12233 0.019716
R57154 ASIG5V.n12243 ASIG5V.n1230 0.019716
R57155 ASIG5V.n12243 ASIG5V.n12242 0.019716
R57156 ASIG5V.n12245 ASIG5V.n1229 0.019716
R57157 ASIG5V.n12246 ASIG5V.n12245 0.019716
R57158 ASIG5V.n12255 ASIG5V.n1228 0.019716
R57159 ASIG5V.n12255 ASIG5V.n12254 0.019716
R57160 ASIG5V.n12257 ASIG5V.n1227 0.019716
R57161 ASIG5V.n12258 ASIG5V.n12257 0.019716
R57162 ASIG5V.n12267 ASIG5V.n12266 0.019716
R57163 ASIG5V.n968 ASIG5V.n967 0.019716
R57164 ASIG5V.n970 ASIG5V.n969 0.019716
R57165 ASIG5V.n971 ASIG5V.n962 0.019716
R57166 ASIG5V.n972 ASIG5V.n971 0.019716
R57167 ASIG5V.n982 ASIG5V.n981 0.019716
R57168 ASIG5V.n981 ASIG5V.n980 0.019716
R57169 ASIG5V.n983 ASIG5V.n958 0.019716
R57170 ASIG5V.n984 ASIG5V.n983 0.019716
R57171 ASIG5V.n994 ASIG5V.n993 0.019716
R57172 ASIG5V.n993 ASIG5V.n992 0.019716
R57173 ASIG5V.n995 ASIG5V.n954 0.019716
R57174 ASIG5V.n996 ASIG5V.n995 0.019716
R57175 ASIG5V.n1006 ASIG5V.n1005 0.019716
R57176 ASIG5V.n1005 ASIG5V.n1004 0.019716
R57177 ASIG5V.n1007 ASIG5V.n950 0.019716
R57178 ASIG5V.n1008 ASIG5V.n1007 0.019716
R57179 ASIG5V.n1018 ASIG5V.n1017 0.019716
R57180 ASIG5V.n1017 ASIG5V.n1016 0.019716
R57181 ASIG5V.n1019 ASIG5V.n946 0.019716
R57182 ASIG5V.n1020 ASIG5V.n1019 0.019716
R57183 ASIG5V.n1030 ASIG5V.n1029 0.019716
R57184 ASIG5V.n1029 ASIG5V.n1028 0.019716
R57185 ASIG5V.n1031 ASIG5V.n942 0.019716
R57186 ASIG5V.n1032 ASIG5V.n1031 0.019716
R57187 ASIG5V.n1042 ASIG5V.n1041 0.019716
R57188 ASIG5V.n1041 ASIG5V.n1040 0.019716
R57189 ASIG5V.n1043 ASIG5V.n938 0.019716
R57190 ASIG5V.n1044 ASIG5V.n1043 0.019716
R57191 ASIG5V.n1054 ASIG5V.n1053 0.019716
R57192 ASIG5V.n1053 ASIG5V.n1052 0.019716
R57193 ASIG5V.n1055 ASIG5V.n934 0.019716
R57194 ASIG5V.n1056 ASIG5V.n1055 0.019716
R57195 ASIG5V.n1066 ASIG5V.n1065 0.019716
R57196 ASIG5V.n1065 ASIG5V.n1064 0.019716
R57197 ASIG5V.n1067 ASIG5V.n930 0.019716
R57198 ASIG5V.n1068 ASIG5V.n1067 0.019716
R57199 ASIG5V.n1078 ASIG5V.n1077 0.019716
R57200 ASIG5V.n1077 ASIG5V.n1076 0.019716
R57201 ASIG5V.n1079 ASIG5V.n926 0.019716
R57202 ASIG5V.n1080 ASIG5V.n1079 0.019716
R57203 ASIG5V.n1090 ASIG5V.n1089 0.019716
R57204 ASIG5V.n1089 ASIG5V.n1088 0.019716
R57205 ASIG5V.n1091 ASIG5V.n922 0.019716
R57206 ASIG5V.n1092 ASIG5V.n1091 0.019716
R57207 ASIG5V.n1102 ASIG5V.n1101 0.019716
R57208 ASIG5V.n1101 ASIG5V.n1100 0.019716
R57209 ASIG5V.n1103 ASIG5V.n918 0.019716
R57210 ASIG5V.n1104 ASIG5V.n1103 0.019716
R57211 ASIG5V.n1114 ASIG5V.n1113 0.019716
R57212 ASIG5V.n1113 ASIG5V.n1112 0.019716
R57213 ASIG5V.n1115 ASIG5V.n914 0.019716
R57214 ASIG5V.n1116 ASIG5V.n1115 0.019716
R57215 ASIG5V.n1126 ASIG5V.n1125 0.019716
R57216 ASIG5V.n1125 ASIG5V.n1124 0.019716
R57217 ASIG5V.n1127 ASIG5V.n910 0.019716
R57218 ASIG5V.n1128 ASIG5V.n1127 0.019716
R57219 ASIG5V.n1138 ASIG5V.n1137 0.019716
R57220 ASIG5V.n1137 ASIG5V.n1136 0.019716
R57221 ASIG5V.n1139 ASIG5V.n906 0.019716
R57222 ASIG5V.n1140 ASIG5V.n1139 0.019716
R57223 ASIG5V.n1150 ASIG5V.n1149 0.019716
R57224 ASIG5V.n1149 ASIG5V.n1148 0.019716
R57225 ASIG5V.n1151 ASIG5V.n902 0.019716
R57226 ASIG5V.n1152 ASIG5V.n1151 0.019716
R57227 ASIG5V.n1162 ASIG5V.n1161 0.019716
R57228 ASIG5V.n1161 ASIG5V.n1160 0.019716
R57229 ASIG5V.n1163 ASIG5V.n898 0.019716
R57230 ASIG5V.n1164 ASIG5V.n1163 0.019716
R57231 ASIG5V.n1174 ASIG5V.n1173 0.019716
R57232 ASIG5V.n1173 ASIG5V.n1172 0.019716
R57233 ASIG5V.n1175 ASIG5V.n894 0.019716
R57234 ASIG5V.n1176 ASIG5V.n1175 0.019716
R57235 ASIG5V.n1186 ASIG5V.n1185 0.019716
R57236 ASIG5V.n1185 ASIG5V.n1184 0.019716
R57237 ASIG5V.n1187 ASIG5V.n890 0.019716
R57238 ASIG5V.n1188 ASIG5V.n1187 0.019716
R57239 ASIG5V.n1198 ASIG5V.n1197 0.019716
R57240 ASIG5V.n1197 ASIG5V.n1196 0.019716
R57241 ASIG5V.n1199 ASIG5V.n886 0.019716
R57242 ASIG5V.n1200 ASIG5V.n1199 0.019716
R57243 ASIG5V.n1211 ASIG5V.n1210 0.019716
R57244 ASIG5V.n1210 ASIG5V.n1209 0.019716
R57245 ASIG5V.n1214 ASIG5V.n1213 0.019716
R57246 ASIG5V.n615 ASIG5V.n570 0.019716
R57247 ASIG5V.n616 ASIG5V.n569 0.019716
R57248 ASIG5V.n623 ASIG5V.n568 0.019716
R57249 ASIG5V.n623 ASIG5V.n622 0.019716
R57250 ASIG5V.n625 ASIG5V.n567 0.019716
R57251 ASIG5V.n626 ASIG5V.n625 0.019716
R57252 ASIG5V.n635 ASIG5V.n566 0.019716
R57253 ASIG5V.n635 ASIG5V.n634 0.019716
R57254 ASIG5V.n637 ASIG5V.n565 0.019716
R57255 ASIG5V.n638 ASIG5V.n637 0.019716
R57256 ASIG5V.n647 ASIG5V.n564 0.019716
R57257 ASIG5V.n647 ASIG5V.n646 0.019716
R57258 ASIG5V.n649 ASIG5V.n563 0.019716
R57259 ASIG5V.n650 ASIG5V.n649 0.019716
R57260 ASIG5V.n659 ASIG5V.n562 0.019716
R57261 ASIG5V.n659 ASIG5V.n658 0.019716
R57262 ASIG5V.n661 ASIG5V.n561 0.019716
R57263 ASIG5V.n662 ASIG5V.n661 0.019716
R57264 ASIG5V.n671 ASIG5V.n560 0.019716
R57265 ASIG5V.n671 ASIG5V.n670 0.019716
R57266 ASIG5V.n673 ASIG5V.n559 0.019716
R57267 ASIG5V.n674 ASIG5V.n673 0.019716
R57268 ASIG5V.n683 ASIG5V.n558 0.019716
R57269 ASIG5V.n683 ASIG5V.n682 0.019716
R57270 ASIG5V.n685 ASIG5V.n557 0.019716
R57271 ASIG5V.n686 ASIG5V.n685 0.019716
R57272 ASIG5V.n695 ASIG5V.n556 0.019716
R57273 ASIG5V.n695 ASIG5V.n694 0.019716
R57274 ASIG5V.n697 ASIG5V.n555 0.019716
R57275 ASIG5V.n698 ASIG5V.n697 0.019716
R57276 ASIG5V.n707 ASIG5V.n554 0.019716
R57277 ASIG5V.n707 ASIG5V.n706 0.019716
R57278 ASIG5V.n709 ASIG5V.n553 0.019716
R57279 ASIG5V.n710 ASIG5V.n709 0.019716
R57280 ASIG5V.n719 ASIG5V.n552 0.019716
R57281 ASIG5V.n719 ASIG5V.n718 0.019716
R57282 ASIG5V.n721 ASIG5V.n551 0.019716
R57283 ASIG5V.n722 ASIG5V.n721 0.019716
R57284 ASIG5V.n731 ASIG5V.n550 0.019716
R57285 ASIG5V.n731 ASIG5V.n730 0.019716
R57286 ASIG5V.n733 ASIG5V.n549 0.019716
R57287 ASIG5V.n734 ASIG5V.n733 0.019716
R57288 ASIG5V.n743 ASIG5V.n548 0.019716
R57289 ASIG5V.n743 ASIG5V.n742 0.019716
R57290 ASIG5V.n745 ASIG5V.n547 0.019716
R57291 ASIG5V.n746 ASIG5V.n745 0.019716
R57292 ASIG5V.n755 ASIG5V.n546 0.019716
R57293 ASIG5V.n755 ASIG5V.n754 0.019716
R57294 ASIG5V.n757 ASIG5V.n545 0.019716
R57295 ASIG5V.n758 ASIG5V.n757 0.019716
R57296 ASIG5V.n767 ASIG5V.n544 0.019716
R57297 ASIG5V.n767 ASIG5V.n766 0.019716
R57298 ASIG5V.n769 ASIG5V.n543 0.019716
R57299 ASIG5V.n770 ASIG5V.n769 0.019716
R57300 ASIG5V.n779 ASIG5V.n542 0.019716
R57301 ASIG5V.n779 ASIG5V.n778 0.019716
R57302 ASIG5V.n781 ASIG5V.n541 0.019716
R57303 ASIG5V.n782 ASIG5V.n781 0.019716
R57304 ASIG5V.n791 ASIG5V.n540 0.019716
R57305 ASIG5V.n791 ASIG5V.n790 0.019716
R57306 ASIG5V.n793 ASIG5V.n539 0.019716
R57307 ASIG5V.n794 ASIG5V.n793 0.019716
R57308 ASIG5V.n803 ASIG5V.n538 0.019716
R57309 ASIG5V.n803 ASIG5V.n802 0.019716
R57310 ASIG5V.n805 ASIG5V.n537 0.019716
R57311 ASIG5V.n806 ASIG5V.n805 0.019716
R57312 ASIG5V.n815 ASIG5V.n536 0.019716
R57313 ASIG5V.n815 ASIG5V.n814 0.019716
R57314 ASIG5V.n817 ASIG5V.n535 0.019716
R57315 ASIG5V.n818 ASIG5V.n817 0.019716
R57316 ASIG5V.n827 ASIG5V.n534 0.019716
R57317 ASIG5V.n827 ASIG5V.n826 0.019716
R57318 ASIG5V.n829 ASIG5V.n533 0.019716
R57319 ASIG5V.n830 ASIG5V.n829 0.019716
R57320 ASIG5V.n839 ASIG5V.n532 0.019716
R57321 ASIG5V.n839 ASIG5V.n838 0.019716
R57322 ASIG5V.n841 ASIG5V.n531 0.019716
R57323 ASIG5V.n842 ASIG5V.n841 0.019716
R57324 ASIG5V.n851 ASIG5V.n530 0.019716
R57325 ASIG5V.n851 ASIG5V.n850 0.019716
R57326 ASIG5V.n853 ASIG5V.n529 0.019716
R57327 ASIG5V.n854 ASIG5V.n853 0.019716
R57328 ASIG5V.n12300 ASIG5V.n12299 0.019716
R57329 ASIG5V.n261 ASIG5V.n215 0.019716
R57330 ASIG5V.n262 ASIG5V.n214 0.019716
R57331 ASIG5V.n269 ASIG5V.n213 0.019716
R57332 ASIG5V.n269 ASIG5V.n268 0.019716
R57333 ASIG5V.n271 ASIG5V.n212 0.019716
R57334 ASIG5V.n272 ASIG5V.n271 0.019716
R57335 ASIG5V.n281 ASIG5V.n211 0.019716
R57336 ASIG5V.n281 ASIG5V.n280 0.019716
R57337 ASIG5V.n283 ASIG5V.n210 0.019716
R57338 ASIG5V.n284 ASIG5V.n283 0.019716
R57339 ASIG5V.n293 ASIG5V.n209 0.019716
R57340 ASIG5V.n293 ASIG5V.n292 0.019716
R57341 ASIG5V.n295 ASIG5V.n208 0.019716
R57342 ASIG5V.n296 ASIG5V.n295 0.019716
R57343 ASIG5V.n305 ASIG5V.n207 0.019716
R57344 ASIG5V.n305 ASIG5V.n304 0.019716
R57345 ASIG5V.n307 ASIG5V.n206 0.019716
R57346 ASIG5V.n308 ASIG5V.n307 0.019716
R57347 ASIG5V.n317 ASIG5V.n205 0.019716
R57348 ASIG5V.n317 ASIG5V.n316 0.019716
R57349 ASIG5V.n319 ASIG5V.n204 0.019716
R57350 ASIG5V.n320 ASIG5V.n319 0.019716
R57351 ASIG5V.n329 ASIG5V.n203 0.019716
R57352 ASIG5V.n329 ASIG5V.n328 0.019716
R57353 ASIG5V.n331 ASIG5V.n202 0.019716
R57354 ASIG5V.n332 ASIG5V.n331 0.019716
R57355 ASIG5V.n341 ASIG5V.n201 0.019716
R57356 ASIG5V.n341 ASIG5V.n340 0.019716
R57357 ASIG5V.n343 ASIG5V.n200 0.019716
R57358 ASIG5V.n344 ASIG5V.n343 0.019716
R57359 ASIG5V.n353 ASIG5V.n199 0.019716
R57360 ASIG5V.n353 ASIG5V.n352 0.019716
R57361 ASIG5V.n355 ASIG5V.n198 0.019716
R57362 ASIG5V.n356 ASIG5V.n355 0.019716
R57363 ASIG5V.n365 ASIG5V.n197 0.019716
R57364 ASIG5V.n365 ASIG5V.n364 0.019716
R57365 ASIG5V.n367 ASIG5V.n196 0.019716
R57366 ASIG5V.n368 ASIG5V.n367 0.019716
R57367 ASIG5V.n377 ASIG5V.n195 0.019716
R57368 ASIG5V.n377 ASIG5V.n376 0.019716
R57369 ASIG5V.n379 ASIG5V.n194 0.019716
R57370 ASIG5V.n380 ASIG5V.n379 0.019716
R57371 ASIG5V.n389 ASIG5V.n193 0.019716
R57372 ASIG5V.n389 ASIG5V.n388 0.019716
R57373 ASIG5V.n391 ASIG5V.n192 0.019716
R57374 ASIG5V.n392 ASIG5V.n391 0.019716
R57375 ASIG5V.n401 ASIG5V.n191 0.019716
R57376 ASIG5V.n401 ASIG5V.n400 0.019716
R57377 ASIG5V.n403 ASIG5V.n190 0.019716
R57378 ASIG5V.n404 ASIG5V.n403 0.019716
R57379 ASIG5V.n413 ASIG5V.n189 0.019716
R57380 ASIG5V.n413 ASIG5V.n412 0.019716
R57381 ASIG5V.n415 ASIG5V.n188 0.019716
R57382 ASIG5V.n416 ASIG5V.n415 0.019716
R57383 ASIG5V.n425 ASIG5V.n187 0.019716
R57384 ASIG5V.n425 ASIG5V.n424 0.019716
R57385 ASIG5V.n427 ASIG5V.n186 0.019716
R57386 ASIG5V.n428 ASIG5V.n427 0.019716
R57387 ASIG5V.n437 ASIG5V.n185 0.019716
R57388 ASIG5V.n437 ASIG5V.n436 0.019716
R57389 ASIG5V.n439 ASIG5V.n184 0.019716
R57390 ASIG5V.n440 ASIG5V.n439 0.019716
R57391 ASIG5V.n449 ASIG5V.n183 0.019716
R57392 ASIG5V.n449 ASIG5V.n448 0.019716
R57393 ASIG5V.n451 ASIG5V.n182 0.019716
R57394 ASIG5V.n452 ASIG5V.n451 0.019716
R57395 ASIG5V.n461 ASIG5V.n181 0.019716
R57396 ASIG5V.n461 ASIG5V.n460 0.019716
R57397 ASIG5V.n463 ASIG5V.n180 0.019716
R57398 ASIG5V.n464 ASIG5V.n463 0.019716
R57399 ASIG5V.n473 ASIG5V.n179 0.019716
R57400 ASIG5V.n473 ASIG5V.n472 0.019716
R57401 ASIG5V.n475 ASIG5V.n178 0.019716
R57402 ASIG5V.n476 ASIG5V.n475 0.019716
R57403 ASIG5V.n485 ASIG5V.n177 0.019716
R57404 ASIG5V.n485 ASIG5V.n484 0.019716
R57405 ASIG5V.n487 ASIG5V.n176 0.019716
R57406 ASIG5V.n488 ASIG5V.n487 0.019716
R57407 ASIG5V.n497 ASIG5V.n175 0.019716
R57408 ASIG5V.n497 ASIG5V.n496 0.019716
R57409 ASIG5V.n499 ASIG5V.n174 0.019716
R57410 ASIG5V.n500 ASIG5V.n499 0.019716
R57411 ASIG5V.n12322 ASIG5V.n12321 0.019716
R57412 ASIG5V.n12527 ASIG5V.n12526 0.019716
R57413 ASIG5V.n97 ASIG5V.n53 0.019716
R57414 ASIG5V.n12343 ASIG5V.n96 0.019716
R57415 ASIG5V.n12343 ASIG5V.n51 0.019716
R57416 ASIG5V.n12347 ASIG5V.n95 0.019716
R57417 ASIG5V.n12347 ASIG5V.n50 0.019716
R57418 ASIG5V.n12352 ASIG5V.n94 0.019716
R57419 ASIG5V.n12352 ASIG5V.n49 0.019716
R57420 ASIG5V.n12356 ASIG5V.n93 0.019716
R57421 ASIG5V.n12356 ASIG5V.n48 0.019716
R57422 ASIG5V.n12361 ASIG5V.n92 0.019716
R57423 ASIG5V.n12361 ASIG5V.n47 0.019716
R57424 ASIG5V.n12365 ASIG5V.n91 0.019716
R57425 ASIG5V.n12365 ASIG5V.n46 0.019716
R57426 ASIG5V.n12370 ASIG5V.n90 0.019716
R57427 ASIG5V.n12370 ASIG5V.n45 0.019716
R57428 ASIG5V.n12374 ASIG5V.n89 0.019716
R57429 ASIG5V.n12374 ASIG5V.n44 0.019716
R57430 ASIG5V.n12379 ASIG5V.n88 0.019716
R57431 ASIG5V.n12379 ASIG5V.n43 0.019716
R57432 ASIG5V.n12383 ASIG5V.n87 0.019716
R57433 ASIG5V.n12383 ASIG5V.n42 0.019716
R57434 ASIG5V.n12388 ASIG5V.n86 0.019716
R57435 ASIG5V.n12388 ASIG5V.n41 0.019716
R57436 ASIG5V.n12392 ASIG5V.n85 0.019716
R57437 ASIG5V.n12392 ASIG5V.n40 0.019716
R57438 ASIG5V.n12397 ASIG5V.n84 0.019716
R57439 ASIG5V.n12397 ASIG5V.n39 0.019716
R57440 ASIG5V.n12401 ASIG5V.n83 0.019716
R57441 ASIG5V.n12401 ASIG5V.n38 0.019716
R57442 ASIG5V.n12406 ASIG5V.n82 0.019716
R57443 ASIG5V.n12406 ASIG5V.n37 0.019716
R57444 ASIG5V.n12410 ASIG5V.n81 0.019716
R57445 ASIG5V.n12410 ASIG5V.n36 0.019716
R57446 ASIG5V.n12415 ASIG5V.n80 0.019716
R57447 ASIG5V.n12415 ASIG5V.n35 0.019716
R57448 ASIG5V.n12419 ASIG5V.n79 0.019716
R57449 ASIG5V.n12419 ASIG5V.n34 0.019716
R57450 ASIG5V.n12424 ASIG5V.n78 0.019716
R57451 ASIG5V.n12424 ASIG5V.n33 0.019716
R57452 ASIG5V.n12428 ASIG5V.n77 0.019716
R57453 ASIG5V.n12428 ASIG5V.n32 0.019716
R57454 ASIG5V.n12433 ASIG5V.n76 0.019716
R57455 ASIG5V.n12433 ASIG5V.n31 0.019716
R57456 ASIG5V.n12437 ASIG5V.n75 0.019716
R57457 ASIG5V.n12437 ASIG5V.n30 0.019716
R57458 ASIG5V.n12442 ASIG5V.n74 0.019716
R57459 ASIG5V.n12442 ASIG5V.n29 0.019716
R57460 ASIG5V.n12446 ASIG5V.n73 0.019716
R57461 ASIG5V.n12446 ASIG5V.n28 0.019716
R57462 ASIG5V.n12451 ASIG5V.n72 0.019716
R57463 ASIG5V.n12451 ASIG5V.n27 0.019716
R57464 ASIG5V.n12455 ASIG5V.n71 0.019716
R57465 ASIG5V.n12455 ASIG5V.n26 0.019716
R57466 ASIG5V.n12460 ASIG5V.n70 0.019716
R57467 ASIG5V.n12460 ASIG5V.n25 0.019716
R57468 ASIG5V.n12464 ASIG5V.n69 0.019716
R57469 ASIG5V.n12464 ASIG5V.n24 0.019716
R57470 ASIG5V.n12469 ASIG5V.n68 0.019716
R57471 ASIG5V.n12469 ASIG5V.n23 0.019716
R57472 ASIG5V.n12473 ASIG5V.n67 0.019716
R57473 ASIG5V.n12473 ASIG5V.n22 0.019716
R57474 ASIG5V.n12478 ASIG5V.n66 0.019716
R57475 ASIG5V.n12478 ASIG5V.n21 0.019716
R57476 ASIG5V.n12482 ASIG5V.n65 0.019716
R57477 ASIG5V.n12482 ASIG5V.n20 0.019716
R57478 ASIG5V.n12487 ASIG5V.n64 0.019716
R57479 ASIG5V.n12487 ASIG5V.n19 0.019716
R57480 ASIG5V.n12491 ASIG5V.n63 0.019716
R57481 ASIG5V.n12491 ASIG5V.n18 0.019716
R57482 ASIG5V.n12496 ASIG5V.n62 0.019716
R57483 ASIG5V.n12496 ASIG5V.n17 0.019716
R57484 ASIG5V.n12500 ASIG5V.n61 0.019716
R57485 ASIG5V.n12500 ASIG5V.n16 0.019716
R57486 ASIG5V.n12505 ASIG5V.n60 0.019716
R57487 ASIG5V.n12505 ASIG5V.n15 0.019716
R57488 ASIG5V.n12509 ASIG5V.n59 0.019716
R57489 ASIG5V.n12509 ASIG5V.n14 0.019716
R57490 ASIG5V.n12514 ASIG5V.n58 0.019716
R57491 ASIG5V.n12514 ASIG5V.n13 0.019716
R57492 ASIG5V.n12518 ASIG5V.n57 0.019716
R57493 ASIG5V.n12518 ASIG5V.n12 0.019716
R57494 ASIG5V.n12524 ASIG5V.n11 0.019716
R57495 ASIG5V.n8880 ASIG5V.n8879 0.019716
R57496 ASIG5V.n8589 ASIG5V.n8319 0.019716
R57497 ASIG5V.n8872 ASIG5V.n8871 0.019716
R57498 ASIG5V.n8872 ASIG5V.n8318 0.019716
R57499 ASIG5V.n8867 ASIG5V.n8866 0.019716
R57500 ASIG5V.n8867 ASIG5V.n8317 0.019716
R57501 ASIG5V.n8860 ASIG5V.n8859 0.019716
R57502 ASIG5V.n8860 ASIG5V.n8316 0.019716
R57503 ASIG5V.n8855 ASIG5V.n8854 0.019716
R57504 ASIG5V.n8855 ASIG5V.n8315 0.019716
R57505 ASIG5V.n8848 ASIG5V.n8847 0.019716
R57506 ASIG5V.n8848 ASIG5V.n8314 0.019716
R57507 ASIG5V.n8843 ASIG5V.n8842 0.019716
R57508 ASIG5V.n8843 ASIG5V.n8313 0.019716
R57509 ASIG5V.n8836 ASIG5V.n8835 0.019716
R57510 ASIG5V.n8836 ASIG5V.n8312 0.019716
R57511 ASIG5V.n8831 ASIG5V.n8830 0.019716
R57512 ASIG5V.n8831 ASIG5V.n8311 0.019716
R57513 ASIG5V.n8824 ASIG5V.n8823 0.019716
R57514 ASIG5V.n8824 ASIG5V.n8310 0.019716
R57515 ASIG5V.n8819 ASIG5V.n8818 0.019716
R57516 ASIG5V.n8819 ASIG5V.n8309 0.019716
R57517 ASIG5V.n8812 ASIG5V.n8811 0.019716
R57518 ASIG5V.n8812 ASIG5V.n8308 0.019716
R57519 ASIG5V.n8807 ASIG5V.n8806 0.019716
R57520 ASIG5V.n8807 ASIG5V.n8307 0.019716
R57521 ASIG5V.n8800 ASIG5V.n8799 0.019716
R57522 ASIG5V.n8800 ASIG5V.n8306 0.019716
R57523 ASIG5V.n8795 ASIG5V.n8794 0.019716
R57524 ASIG5V.n8795 ASIG5V.n8305 0.019716
R57525 ASIG5V.n8788 ASIG5V.n8787 0.019716
R57526 ASIG5V.n8788 ASIG5V.n8304 0.019716
R57527 ASIG5V.n8783 ASIG5V.n8782 0.019716
R57528 ASIG5V.n8783 ASIG5V.n8303 0.019716
R57529 ASIG5V.n8776 ASIG5V.n8775 0.019716
R57530 ASIG5V.n8776 ASIG5V.n8302 0.019716
R57531 ASIG5V.n8771 ASIG5V.n8770 0.019716
R57532 ASIG5V.n8771 ASIG5V.n8301 0.019716
R57533 ASIG5V.n8764 ASIG5V.n8763 0.019716
R57534 ASIG5V.n8764 ASIG5V.n8300 0.019716
R57535 ASIG5V.n8759 ASIG5V.n8758 0.019716
R57536 ASIG5V.n8759 ASIG5V.n8299 0.019716
R57537 ASIG5V.n8752 ASIG5V.n8751 0.019716
R57538 ASIG5V.n8752 ASIG5V.n8298 0.019716
R57539 ASIG5V.n8747 ASIG5V.n8746 0.019716
R57540 ASIG5V.n8747 ASIG5V.n8297 0.019716
R57541 ASIG5V.n8740 ASIG5V.n8739 0.019716
R57542 ASIG5V.n8740 ASIG5V.n8296 0.019716
R57543 ASIG5V.n8735 ASIG5V.n8734 0.019716
R57544 ASIG5V.n8735 ASIG5V.n8295 0.019716
R57545 ASIG5V.n8728 ASIG5V.n8727 0.019716
R57546 ASIG5V.n8728 ASIG5V.n8294 0.019716
R57547 ASIG5V.n8723 ASIG5V.n8722 0.019716
R57548 ASIG5V.n8723 ASIG5V.n8293 0.019716
R57549 ASIG5V.n8716 ASIG5V.n8715 0.019716
R57550 ASIG5V.n8716 ASIG5V.n8292 0.019716
R57551 ASIG5V.n8711 ASIG5V.n8710 0.019716
R57552 ASIG5V.n8711 ASIG5V.n8291 0.019716
R57553 ASIG5V.n8704 ASIG5V.n8703 0.019716
R57554 ASIG5V.n8704 ASIG5V.n8290 0.019716
R57555 ASIG5V.n8699 ASIG5V.n8698 0.019716
R57556 ASIG5V.n8699 ASIG5V.n8289 0.019716
R57557 ASIG5V.n8692 ASIG5V.n8691 0.019716
R57558 ASIG5V.n8692 ASIG5V.n8288 0.019716
R57559 ASIG5V.n8687 ASIG5V.n8686 0.019716
R57560 ASIG5V.n8687 ASIG5V.n8287 0.019716
R57561 ASIG5V.n8680 ASIG5V.n8679 0.019716
R57562 ASIG5V.n8680 ASIG5V.n8286 0.019716
R57563 ASIG5V.n8675 ASIG5V.n8674 0.019716
R57564 ASIG5V.n8675 ASIG5V.n8285 0.019716
R57565 ASIG5V.n8668 ASIG5V.n8667 0.019716
R57566 ASIG5V.n8668 ASIG5V.n8284 0.019716
R57567 ASIG5V.n8663 ASIG5V.n8662 0.019716
R57568 ASIG5V.n8663 ASIG5V.n8283 0.019716
R57569 ASIG5V.n8656 ASIG5V.n8655 0.019716
R57570 ASIG5V.n8656 ASIG5V.n8282 0.019716
R57571 ASIG5V.n8651 ASIG5V.n8650 0.019716
R57572 ASIG5V.n8651 ASIG5V.n8281 0.019716
R57573 ASIG5V.n8644 ASIG5V.n8643 0.019716
R57574 ASIG5V.n8644 ASIG5V.n8280 0.019716
R57575 ASIG5V.n8639 ASIG5V.n8638 0.019716
R57576 ASIG5V.n8639 ASIG5V.n8279 0.019716
R57577 ASIG5V.n8632 ASIG5V.n8278 0.019716
R57578 ASIG5V.n8894 ASIG5V.n8893 0.019716
R57579 ASIG5V.n8258 ASIG5V.n8214 0.019716
R57580 ASIG5V.n8562 ASIG5V.n8257 0.019716
R57581 ASIG5V.n8562 ASIG5V.n8212 0.019716
R57582 ASIG5V.n8557 ASIG5V.n8256 0.019716
R57583 ASIG5V.n8557 ASIG5V.n8211 0.019716
R57584 ASIG5V.n8553 ASIG5V.n8255 0.019716
R57585 ASIG5V.n8553 ASIG5V.n8210 0.019716
R57586 ASIG5V.n8548 ASIG5V.n8254 0.019716
R57587 ASIG5V.n8548 ASIG5V.n8209 0.019716
R57588 ASIG5V.n8544 ASIG5V.n8253 0.019716
R57589 ASIG5V.n8544 ASIG5V.n8208 0.019716
R57590 ASIG5V.n8539 ASIG5V.n8252 0.019716
R57591 ASIG5V.n8539 ASIG5V.n8207 0.019716
R57592 ASIG5V.n8535 ASIG5V.n8251 0.019716
R57593 ASIG5V.n8535 ASIG5V.n8206 0.019716
R57594 ASIG5V.n8530 ASIG5V.n8250 0.019716
R57595 ASIG5V.n8530 ASIG5V.n8205 0.019716
R57596 ASIG5V.n8526 ASIG5V.n8249 0.019716
R57597 ASIG5V.n8526 ASIG5V.n8204 0.019716
R57598 ASIG5V.n8521 ASIG5V.n8248 0.019716
R57599 ASIG5V.n8521 ASIG5V.n8203 0.019716
R57600 ASIG5V.n8517 ASIG5V.n8247 0.019716
R57601 ASIG5V.n8517 ASIG5V.n8202 0.019716
R57602 ASIG5V.n8512 ASIG5V.n8246 0.019716
R57603 ASIG5V.n8512 ASIG5V.n8201 0.019716
R57604 ASIG5V.n8508 ASIG5V.n8245 0.019716
R57605 ASIG5V.n8508 ASIG5V.n8200 0.019716
R57606 ASIG5V.n8503 ASIG5V.n8244 0.019716
R57607 ASIG5V.n8503 ASIG5V.n8199 0.019716
R57608 ASIG5V.n8499 ASIG5V.n8243 0.019716
R57609 ASIG5V.n8499 ASIG5V.n8198 0.019716
R57610 ASIG5V.n8494 ASIG5V.n8242 0.019716
R57611 ASIG5V.n8494 ASIG5V.n8197 0.019716
R57612 ASIG5V.n8490 ASIG5V.n8241 0.019716
R57613 ASIG5V.n8490 ASIG5V.n8196 0.019716
R57614 ASIG5V.n8485 ASIG5V.n8240 0.019716
R57615 ASIG5V.n8485 ASIG5V.n8195 0.019716
R57616 ASIG5V.n8481 ASIG5V.n8239 0.019716
R57617 ASIG5V.n8481 ASIG5V.n8194 0.019716
R57618 ASIG5V.n8476 ASIG5V.n8238 0.019716
R57619 ASIG5V.n8476 ASIG5V.n8193 0.019716
R57620 ASIG5V.n8472 ASIG5V.n8237 0.019716
R57621 ASIG5V.n8472 ASIG5V.n8192 0.019716
R57622 ASIG5V.n8467 ASIG5V.n8236 0.019716
R57623 ASIG5V.n8467 ASIG5V.n8191 0.019716
R57624 ASIG5V.n8463 ASIG5V.n8235 0.019716
R57625 ASIG5V.n8463 ASIG5V.n8190 0.019716
R57626 ASIG5V.n8458 ASIG5V.n8234 0.019716
R57627 ASIG5V.n8458 ASIG5V.n8189 0.019716
R57628 ASIG5V.n8454 ASIG5V.n8233 0.019716
R57629 ASIG5V.n8454 ASIG5V.n8188 0.019716
R57630 ASIG5V.n8449 ASIG5V.n8232 0.019716
R57631 ASIG5V.n8449 ASIG5V.n8187 0.019716
R57632 ASIG5V.n8445 ASIG5V.n8231 0.019716
R57633 ASIG5V.n8445 ASIG5V.n8186 0.019716
R57634 ASIG5V.n8440 ASIG5V.n8230 0.019716
R57635 ASIG5V.n8440 ASIG5V.n8185 0.019716
R57636 ASIG5V.n8436 ASIG5V.n8229 0.019716
R57637 ASIG5V.n8436 ASIG5V.n8184 0.019716
R57638 ASIG5V.n8431 ASIG5V.n8228 0.019716
R57639 ASIG5V.n8431 ASIG5V.n8183 0.019716
R57640 ASIG5V.n8427 ASIG5V.n8227 0.019716
R57641 ASIG5V.n8427 ASIG5V.n8182 0.019716
R57642 ASIG5V.n8422 ASIG5V.n8226 0.019716
R57643 ASIG5V.n8422 ASIG5V.n8181 0.019716
R57644 ASIG5V.n8418 ASIG5V.n8225 0.019716
R57645 ASIG5V.n8418 ASIG5V.n8180 0.019716
R57646 ASIG5V.n8413 ASIG5V.n8224 0.019716
R57647 ASIG5V.n8413 ASIG5V.n8179 0.019716
R57648 ASIG5V.n8409 ASIG5V.n8223 0.019716
R57649 ASIG5V.n8409 ASIG5V.n8178 0.019716
R57650 ASIG5V.n8404 ASIG5V.n8222 0.019716
R57651 ASIG5V.n8404 ASIG5V.n8177 0.019716
R57652 ASIG5V.n8400 ASIG5V.n8221 0.019716
R57653 ASIG5V.n8400 ASIG5V.n8176 0.019716
R57654 ASIG5V.n8395 ASIG5V.n8220 0.019716
R57655 ASIG5V.n8395 ASIG5V.n8175 0.019716
R57656 ASIG5V.n8391 ASIG5V.n8219 0.019716
R57657 ASIG5V.n8391 ASIG5V.n8174 0.019716
R57658 ASIG5V.n8386 ASIG5V.n8218 0.019716
R57659 ASIG5V.n8386 ASIG5V.n8173 0.019716
R57660 ASIG5V.n8891 ASIG5V.n8172 0.019716
R57661 ASIG5V.n7229 ASIG5V.n7228 0.019716
R57662 ASIG5V.n7227 ASIG5V.n7226 0.019716
R57663 ASIG5V.n6904 ASIG5V.n6903 0.019716
R57664 ASIG5V.n6903 ASIG5V.n6899 0.019716
R57665 ASIG5V.n7217 ASIG5V.n7216 0.019716
R57666 ASIG5V.n7218 ASIG5V.n7217 0.019716
R57667 ASIG5V.n6910 ASIG5V.n6909 0.019716
R57668 ASIG5V.n6909 ASIG5V.n6905 0.019716
R57669 ASIG5V.n7207 ASIG5V.n7206 0.019716
R57670 ASIG5V.n7208 ASIG5V.n7207 0.019716
R57671 ASIG5V.n6916 ASIG5V.n6915 0.019716
R57672 ASIG5V.n6915 ASIG5V.n6911 0.019716
R57673 ASIG5V.n7197 ASIG5V.n7196 0.019716
R57674 ASIG5V.n7198 ASIG5V.n7197 0.019716
R57675 ASIG5V.n6922 ASIG5V.n6921 0.019716
R57676 ASIG5V.n6921 ASIG5V.n6917 0.019716
R57677 ASIG5V.n7187 ASIG5V.n7186 0.019716
R57678 ASIG5V.n7188 ASIG5V.n7187 0.019716
R57679 ASIG5V.n6928 ASIG5V.n6927 0.019716
R57680 ASIG5V.n6927 ASIG5V.n6923 0.019716
R57681 ASIG5V.n7177 ASIG5V.n7176 0.019716
R57682 ASIG5V.n7178 ASIG5V.n7177 0.019716
R57683 ASIG5V.n6934 ASIG5V.n6933 0.019716
R57684 ASIG5V.n6933 ASIG5V.n6929 0.019716
R57685 ASIG5V.n7167 ASIG5V.n7166 0.019716
R57686 ASIG5V.n7168 ASIG5V.n7167 0.019716
R57687 ASIG5V.n6940 ASIG5V.n6939 0.019716
R57688 ASIG5V.n6939 ASIG5V.n6935 0.019716
R57689 ASIG5V.n7157 ASIG5V.n7156 0.019716
R57690 ASIG5V.n7158 ASIG5V.n7157 0.019716
R57691 ASIG5V.n6946 ASIG5V.n6945 0.019716
R57692 ASIG5V.n6945 ASIG5V.n6941 0.019716
R57693 ASIG5V.n7147 ASIG5V.n7146 0.019716
R57694 ASIG5V.n7148 ASIG5V.n7147 0.019716
R57695 ASIG5V.n6952 ASIG5V.n6951 0.019716
R57696 ASIG5V.n6951 ASIG5V.n6947 0.019716
R57697 ASIG5V.n7137 ASIG5V.n7136 0.019716
R57698 ASIG5V.n7138 ASIG5V.n7137 0.019716
R57699 ASIG5V.n6958 ASIG5V.n6957 0.019716
R57700 ASIG5V.n6957 ASIG5V.n6953 0.019716
R57701 ASIG5V.n7127 ASIG5V.n7126 0.019716
R57702 ASIG5V.n7128 ASIG5V.n7127 0.019716
R57703 ASIG5V.n6964 ASIG5V.n6963 0.019716
R57704 ASIG5V.n6963 ASIG5V.n6959 0.019716
R57705 ASIG5V.n7117 ASIG5V.n7116 0.019716
R57706 ASIG5V.n7118 ASIG5V.n7117 0.019716
R57707 ASIG5V.n6970 ASIG5V.n6969 0.019716
R57708 ASIG5V.n6969 ASIG5V.n6965 0.019716
R57709 ASIG5V.n7107 ASIG5V.n7106 0.019716
R57710 ASIG5V.n7108 ASIG5V.n7107 0.019716
R57711 ASIG5V.n6976 ASIG5V.n6975 0.019716
R57712 ASIG5V.n6975 ASIG5V.n6971 0.019716
R57713 ASIG5V.n7097 ASIG5V.n7096 0.019716
R57714 ASIG5V.n7098 ASIG5V.n7097 0.019716
R57715 ASIG5V.n6982 ASIG5V.n6981 0.019716
R57716 ASIG5V.n6981 ASIG5V.n6977 0.019716
R57717 ASIG5V.n7087 ASIG5V.n7086 0.019716
R57718 ASIG5V.n7088 ASIG5V.n7087 0.019716
R57719 ASIG5V.n6988 ASIG5V.n6987 0.019716
R57720 ASIG5V.n6987 ASIG5V.n6983 0.019716
R57721 ASIG5V.n7077 ASIG5V.n7076 0.019716
R57722 ASIG5V.n7078 ASIG5V.n7077 0.019716
R57723 ASIG5V.n6994 ASIG5V.n6993 0.019716
R57724 ASIG5V.n6993 ASIG5V.n6989 0.019716
R57725 ASIG5V.n7067 ASIG5V.n7066 0.019716
R57726 ASIG5V.n7068 ASIG5V.n7067 0.019716
R57727 ASIG5V.n7000 ASIG5V.n6999 0.019716
R57728 ASIG5V.n6999 ASIG5V.n6995 0.019716
R57729 ASIG5V.n7057 ASIG5V.n7056 0.019716
R57730 ASIG5V.n7058 ASIG5V.n7057 0.019716
R57731 ASIG5V.n7006 ASIG5V.n7005 0.019716
R57732 ASIG5V.n7005 ASIG5V.n7001 0.019716
R57733 ASIG5V.n7047 ASIG5V.n7046 0.019716
R57734 ASIG5V.n7048 ASIG5V.n7047 0.019716
R57735 ASIG5V.n7012 ASIG5V.n7011 0.019716
R57736 ASIG5V.n7011 ASIG5V.n7007 0.019716
R57737 ASIG5V.n7037 ASIG5V.n7036 0.019716
R57738 ASIG5V.n7038 ASIG5V.n7037 0.019716
R57739 ASIG5V.n7018 ASIG5V.n7017 0.019716
R57740 ASIG5V.n7017 ASIG5V.n7013 0.019716
R57741 ASIG5V.n7027 ASIG5V.n7026 0.019716
R57742 ASIG5V.n7028 ASIG5V.n7027 0.019716
R57743 ASIG5V.n7020 ASIG5V.n7019 0.019716
R57744 ASIG5V.n8918 ASIG5V.n8917 0.019716
R57745 ASIG5V.n6631 ASIG5V.n6588 0.019716
R57746 ASIG5V.n6701 ASIG5V.n6630 0.019716
R57747 ASIG5V.n6701 ASIG5V.n6586 0.019716
R57748 ASIG5V.n6705 ASIG5V.n6629 0.019716
R57749 ASIG5V.n6705 ASIG5V.n6585 0.019716
R57750 ASIG5V.n6710 ASIG5V.n6628 0.019716
R57751 ASIG5V.n6710 ASIG5V.n6584 0.019716
R57752 ASIG5V.n6714 ASIG5V.n6627 0.019716
R57753 ASIG5V.n6714 ASIG5V.n6583 0.019716
R57754 ASIG5V.n6719 ASIG5V.n6626 0.019716
R57755 ASIG5V.n6719 ASIG5V.n6582 0.019716
R57756 ASIG5V.n6723 ASIG5V.n6625 0.019716
R57757 ASIG5V.n6723 ASIG5V.n6581 0.019716
R57758 ASIG5V.n6728 ASIG5V.n6624 0.019716
R57759 ASIG5V.n6728 ASIG5V.n6580 0.019716
R57760 ASIG5V.n6732 ASIG5V.n6623 0.019716
R57761 ASIG5V.n6732 ASIG5V.n6579 0.019716
R57762 ASIG5V.n6737 ASIG5V.n6622 0.019716
R57763 ASIG5V.n6737 ASIG5V.n6578 0.019716
R57764 ASIG5V.n6741 ASIG5V.n6621 0.019716
R57765 ASIG5V.n6741 ASIG5V.n6577 0.019716
R57766 ASIG5V.n6746 ASIG5V.n6620 0.019716
R57767 ASIG5V.n6746 ASIG5V.n6576 0.019716
R57768 ASIG5V.n6750 ASIG5V.n6619 0.019716
R57769 ASIG5V.n6750 ASIG5V.n6575 0.019716
R57770 ASIG5V.n6755 ASIG5V.n6618 0.019716
R57771 ASIG5V.n6755 ASIG5V.n6574 0.019716
R57772 ASIG5V.n6759 ASIG5V.n6617 0.019716
R57773 ASIG5V.n6759 ASIG5V.n6573 0.019716
R57774 ASIG5V.n6764 ASIG5V.n6616 0.019716
R57775 ASIG5V.n6764 ASIG5V.n6572 0.019716
R57776 ASIG5V.n6768 ASIG5V.n6615 0.019716
R57777 ASIG5V.n6768 ASIG5V.n6571 0.019716
R57778 ASIG5V.n6773 ASIG5V.n6614 0.019716
R57779 ASIG5V.n6773 ASIG5V.n6570 0.019716
R57780 ASIG5V.n6777 ASIG5V.n6613 0.019716
R57781 ASIG5V.n6777 ASIG5V.n6569 0.019716
R57782 ASIG5V.n6782 ASIG5V.n6612 0.019716
R57783 ASIG5V.n6782 ASIG5V.n6568 0.019716
R57784 ASIG5V.n6786 ASIG5V.n6611 0.019716
R57785 ASIG5V.n6786 ASIG5V.n6567 0.019716
R57786 ASIG5V.n6791 ASIG5V.n6610 0.019716
R57787 ASIG5V.n6791 ASIG5V.n6566 0.019716
R57788 ASIG5V.n6795 ASIG5V.n6609 0.019716
R57789 ASIG5V.n6795 ASIG5V.n6565 0.019716
R57790 ASIG5V.n6800 ASIG5V.n6608 0.019716
R57791 ASIG5V.n6800 ASIG5V.n6564 0.019716
R57792 ASIG5V.n6804 ASIG5V.n6607 0.019716
R57793 ASIG5V.n6804 ASIG5V.n6563 0.019716
R57794 ASIG5V.n6809 ASIG5V.n6606 0.019716
R57795 ASIG5V.n6809 ASIG5V.n6562 0.019716
R57796 ASIG5V.n6813 ASIG5V.n6605 0.019716
R57797 ASIG5V.n6813 ASIG5V.n6561 0.019716
R57798 ASIG5V.n6818 ASIG5V.n6604 0.019716
R57799 ASIG5V.n6818 ASIG5V.n6560 0.019716
R57800 ASIG5V.n6822 ASIG5V.n6603 0.019716
R57801 ASIG5V.n6822 ASIG5V.n6559 0.019716
R57802 ASIG5V.n6827 ASIG5V.n6602 0.019716
R57803 ASIG5V.n6827 ASIG5V.n6558 0.019716
R57804 ASIG5V.n6831 ASIG5V.n6601 0.019716
R57805 ASIG5V.n6831 ASIG5V.n6557 0.019716
R57806 ASIG5V.n6836 ASIG5V.n6600 0.019716
R57807 ASIG5V.n6836 ASIG5V.n6556 0.019716
R57808 ASIG5V.n6840 ASIG5V.n6599 0.019716
R57809 ASIG5V.n6840 ASIG5V.n6555 0.019716
R57810 ASIG5V.n6845 ASIG5V.n6598 0.019716
R57811 ASIG5V.n6845 ASIG5V.n6554 0.019716
R57812 ASIG5V.n6849 ASIG5V.n6597 0.019716
R57813 ASIG5V.n6849 ASIG5V.n6553 0.019716
R57814 ASIG5V.n6854 ASIG5V.n6596 0.019716
R57815 ASIG5V.n6854 ASIG5V.n6552 0.019716
R57816 ASIG5V.n6858 ASIG5V.n6595 0.019716
R57817 ASIG5V.n6858 ASIG5V.n6551 0.019716
R57818 ASIG5V.n6863 ASIG5V.n6594 0.019716
R57819 ASIG5V.n6863 ASIG5V.n6550 0.019716
R57820 ASIG5V.n6867 ASIG5V.n6593 0.019716
R57821 ASIG5V.n6867 ASIG5V.n6549 0.019716
R57822 ASIG5V.n6872 ASIG5V.n6592 0.019716
R57823 ASIG5V.n6872 ASIG5V.n6548 0.019716
R57824 ASIG5V.n6876 ASIG5V.n6591 0.019716
R57825 ASIG5V.n6876 ASIG5V.n6547 0.019716
R57826 ASIG5V.n8915 ASIG5V.n6546 0.019716
R57827 ASIG5V.n6530 ASIG5V.n6487 0.019716
R57828 ASIG5V.n6531 ASIG5V.n6486 0.019716
R57829 ASIG5V.n8935 ASIG5V.n6485 0.019716
R57830 ASIG5V.n8935 ASIG5V.n8934 0.019716
R57831 ASIG5V.n8937 ASIG5V.n6484 0.019716
R57832 ASIG5V.n8938 ASIG5V.n8937 0.019716
R57833 ASIG5V.n8947 ASIG5V.n6483 0.019716
R57834 ASIG5V.n8947 ASIG5V.n8946 0.019716
R57835 ASIG5V.n8949 ASIG5V.n6482 0.019716
R57836 ASIG5V.n8950 ASIG5V.n8949 0.019716
R57837 ASIG5V.n8959 ASIG5V.n6481 0.019716
R57838 ASIG5V.n8959 ASIG5V.n8958 0.019716
R57839 ASIG5V.n8961 ASIG5V.n6480 0.019716
R57840 ASIG5V.n8962 ASIG5V.n8961 0.019716
R57841 ASIG5V.n8971 ASIG5V.n6479 0.019716
R57842 ASIG5V.n8971 ASIG5V.n8970 0.019716
R57843 ASIG5V.n8973 ASIG5V.n6478 0.019716
R57844 ASIG5V.n8974 ASIG5V.n8973 0.019716
R57845 ASIG5V.n8983 ASIG5V.n6477 0.019716
R57846 ASIG5V.n8983 ASIG5V.n8982 0.019716
R57847 ASIG5V.n8985 ASIG5V.n6476 0.019716
R57848 ASIG5V.n8986 ASIG5V.n8985 0.019716
R57849 ASIG5V.n8995 ASIG5V.n6475 0.019716
R57850 ASIG5V.n8995 ASIG5V.n8994 0.019716
R57851 ASIG5V.n8997 ASIG5V.n6474 0.019716
R57852 ASIG5V.n8998 ASIG5V.n8997 0.019716
R57853 ASIG5V.n9007 ASIG5V.n6473 0.019716
R57854 ASIG5V.n9007 ASIG5V.n9006 0.019716
R57855 ASIG5V.n9009 ASIG5V.n6472 0.019716
R57856 ASIG5V.n9010 ASIG5V.n9009 0.019716
R57857 ASIG5V.n9019 ASIG5V.n6471 0.019716
R57858 ASIG5V.n9019 ASIG5V.n9018 0.019716
R57859 ASIG5V.n9021 ASIG5V.n6470 0.019716
R57860 ASIG5V.n9022 ASIG5V.n9021 0.019716
R57861 ASIG5V.n9031 ASIG5V.n6469 0.019716
R57862 ASIG5V.n9031 ASIG5V.n9030 0.019716
R57863 ASIG5V.n9033 ASIG5V.n6468 0.019716
R57864 ASIG5V.n9034 ASIG5V.n9033 0.019716
R57865 ASIG5V.n9043 ASIG5V.n6467 0.019716
R57866 ASIG5V.n9043 ASIG5V.n9042 0.019716
R57867 ASIG5V.n9045 ASIG5V.n6466 0.019716
R57868 ASIG5V.n9046 ASIG5V.n9045 0.019716
R57869 ASIG5V.n9055 ASIG5V.n6465 0.019716
R57870 ASIG5V.n9055 ASIG5V.n9054 0.019716
R57871 ASIG5V.n9057 ASIG5V.n6464 0.019716
R57872 ASIG5V.n9058 ASIG5V.n9057 0.019716
R57873 ASIG5V.n9067 ASIG5V.n6463 0.019716
R57874 ASIG5V.n9067 ASIG5V.n9066 0.019716
R57875 ASIG5V.n9069 ASIG5V.n6462 0.019716
R57876 ASIG5V.n9070 ASIG5V.n9069 0.019716
R57877 ASIG5V.n9079 ASIG5V.n6461 0.019716
R57878 ASIG5V.n9079 ASIG5V.n9078 0.019716
R57879 ASIG5V.n9081 ASIG5V.n6460 0.019716
R57880 ASIG5V.n9082 ASIG5V.n9081 0.019716
R57881 ASIG5V.n9091 ASIG5V.n6459 0.019716
R57882 ASIG5V.n9091 ASIG5V.n9090 0.019716
R57883 ASIG5V.n9093 ASIG5V.n6458 0.019716
R57884 ASIG5V.n9094 ASIG5V.n9093 0.019716
R57885 ASIG5V.n9103 ASIG5V.n6457 0.019716
R57886 ASIG5V.n9103 ASIG5V.n9102 0.019716
R57887 ASIG5V.n9105 ASIG5V.n6456 0.019716
R57888 ASIG5V.n9106 ASIG5V.n9105 0.019716
R57889 ASIG5V.n9115 ASIG5V.n6455 0.019716
R57890 ASIG5V.n9115 ASIG5V.n9114 0.019716
R57891 ASIG5V.n9117 ASIG5V.n6454 0.019716
R57892 ASIG5V.n9118 ASIG5V.n9117 0.019716
R57893 ASIG5V.n9127 ASIG5V.n6453 0.019716
R57894 ASIG5V.n9127 ASIG5V.n9126 0.019716
R57895 ASIG5V.n9129 ASIG5V.n6452 0.019716
R57896 ASIG5V.n9130 ASIG5V.n9129 0.019716
R57897 ASIG5V.n9139 ASIG5V.n6451 0.019716
R57898 ASIG5V.n9139 ASIG5V.n9138 0.019716
R57899 ASIG5V.n9141 ASIG5V.n6450 0.019716
R57900 ASIG5V.n9142 ASIG5V.n9141 0.019716
R57901 ASIG5V.n9151 ASIG5V.n6449 0.019716
R57902 ASIG5V.n9151 ASIG5V.n9150 0.019716
R57903 ASIG5V.n9153 ASIG5V.n6448 0.019716
R57904 ASIG5V.n9154 ASIG5V.n9153 0.019716
R57905 ASIG5V.n9163 ASIG5V.n6447 0.019716
R57906 ASIG5V.n9163 ASIG5V.n9162 0.019716
R57907 ASIG5V.n9165 ASIG5V.n6446 0.019716
R57908 ASIG5V.n9166 ASIG5V.n9165 0.019716
R57909 ASIG5V.n9175 ASIG5V.n9174 0.019716
R57910 ASIG5V.n9381 ASIG5V.n9380 0.019716
R57911 ASIG5V.n6351 ASIG5V.n6307 0.019716
R57912 ASIG5V.n9197 ASIG5V.n6350 0.019716
R57913 ASIG5V.n9197 ASIG5V.n6305 0.019716
R57914 ASIG5V.n9201 ASIG5V.n6349 0.019716
R57915 ASIG5V.n9201 ASIG5V.n6304 0.019716
R57916 ASIG5V.n9206 ASIG5V.n6348 0.019716
R57917 ASIG5V.n9206 ASIG5V.n6303 0.019716
R57918 ASIG5V.n9210 ASIG5V.n6347 0.019716
R57919 ASIG5V.n9210 ASIG5V.n6302 0.019716
R57920 ASIG5V.n9215 ASIG5V.n6346 0.019716
R57921 ASIG5V.n9215 ASIG5V.n6301 0.019716
R57922 ASIG5V.n9219 ASIG5V.n6345 0.019716
R57923 ASIG5V.n9219 ASIG5V.n6300 0.019716
R57924 ASIG5V.n9224 ASIG5V.n6344 0.019716
R57925 ASIG5V.n9224 ASIG5V.n6299 0.019716
R57926 ASIG5V.n9228 ASIG5V.n6343 0.019716
R57927 ASIG5V.n9228 ASIG5V.n6298 0.019716
R57928 ASIG5V.n9233 ASIG5V.n6342 0.019716
R57929 ASIG5V.n9233 ASIG5V.n6297 0.019716
R57930 ASIG5V.n9237 ASIG5V.n6341 0.019716
R57931 ASIG5V.n9237 ASIG5V.n6296 0.019716
R57932 ASIG5V.n9242 ASIG5V.n6340 0.019716
R57933 ASIG5V.n9242 ASIG5V.n6295 0.019716
R57934 ASIG5V.n9246 ASIG5V.n6339 0.019716
R57935 ASIG5V.n9246 ASIG5V.n6294 0.019716
R57936 ASIG5V.n9251 ASIG5V.n6338 0.019716
R57937 ASIG5V.n9251 ASIG5V.n6293 0.019716
R57938 ASIG5V.n9255 ASIG5V.n6337 0.019716
R57939 ASIG5V.n9255 ASIG5V.n6292 0.019716
R57940 ASIG5V.n9260 ASIG5V.n6336 0.019716
R57941 ASIG5V.n9260 ASIG5V.n6291 0.019716
R57942 ASIG5V.n9264 ASIG5V.n6335 0.019716
R57943 ASIG5V.n9264 ASIG5V.n6290 0.019716
R57944 ASIG5V.n9269 ASIG5V.n6334 0.019716
R57945 ASIG5V.n9269 ASIG5V.n6289 0.019716
R57946 ASIG5V.n9273 ASIG5V.n6333 0.019716
R57947 ASIG5V.n9273 ASIG5V.n6288 0.019716
R57948 ASIG5V.n9278 ASIG5V.n6332 0.019716
R57949 ASIG5V.n9278 ASIG5V.n6287 0.019716
R57950 ASIG5V.n9282 ASIG5V.n6331 0.019716
R57951 ASIG5V.n9282 ASIG5V.n6286 0.019716
R57952 ASIG5V.n9287 ASIG5V.n6330 0.019716
R57953 ASIG5V.n9287 ASIG5V.n6285 0.019716
R57954 ASIG5V.n9291 ASIG5V.n6329 0.019716
R57955 ASIG5V.n9291 ASIG5V.n6284 0.019716
R57956 ASIG5V.n9296 ASIG5V.n6328 0.019716
R57957 ASIG5V.n9296 ASIG5V.n6283 0.019716
R57958 ASIG5V.n9300 ASIG5V.n6327 0.019716
R57959 ASIG5V.n9300 ASIG5V.n6282 0.019716
R57960 ASIG5V.n9305 ASIG5V.n6326 0.019716
R57961 ASIG5V.n9305 ASIG5V.n6281 0.019716
R57962 ASIG5V.n9309 ASIG5V.n6325 0.019716
R57963 ASIG5V.n9309 ASIG5V.n6280 0.019716
R57964 ASIG5V.n9314 ASIG5V.n6324 0.019716
R57965 ASIG5V.n9314 ASIG5V.n6279 0.019716
R57966 ASIG5V.n9318 ASIG5V.n6323 0.019716
R57967 ASIG5V.n9318 ASIG5V.n6278 0.019716
R57968 ASIG5V.n9323 ASIG5V.n6322 0.019716
R57969 ASIG5V.n9323 ASIG5V.n6277 0.019716
R57970 ASIG5V.n9327 ASIG5V.n6321 0.019716
R57971 ASIG5V.n9327 ASIG5V.n6276 0.019716
R57972 ASIG5V.n9332 ASIG5V.n6320 0.019716
R57973 ASIG5V.n9332 ASIG5V.n6275 0.019716
R57974 ASIG5V.n9336 ASIG5V.n6319 0.019716
R57975 ASIG5V.n9336 ASIG5V.n6274 0.019716
R57976 ASIG5V.n9341 ASIG5V.n6318 0.019716
R57977 ASIG5V.n9341 ASIG5V.n6273 0.019716
R57978 ASIG5V.n9345 ASIG5V.n6317 0.019716
R57979 ASIG5V.n9345 ASIG5V.n6272 0.019716
R57980 ASIG5V.n9350 ASIG5V.n6316 0.019716
R57981 ASIG5V.n9350 ASIG5V.n6271 0.019716
R57982 ASIG5V.n9354 ASIG5V.n6315 0.019716
R57983 ASIG5V.n9354 ASIG5V.n6270 0.019716
R57984 ASIG5V.n9359 ASIG5V.n6314 0.019716
R57985 ASIG5V.n9359 ASIG5V.n6269 0.019716
R57986 ASIG5V.n9363 ASIG5V.n6313 0.019716
R57987 ASIG5V.n9363 ASIG5V.n6268 0.019716
R57988 ASIG5V.n9368 ASIG5V.n6312 0.019716
R57989 ASIG5V.n9368 ASIG5V.n6267 0.019716
R57990 ASIG5V.n9372 ASIG5V.n6311 0.019716
R57991 ASIG5V.n9372 ASIG5V.n6266 0.019716
R57992 ASIG5V.n9378 ASIG5V.n6265 0.019716
R57993 ASIG5V.n9395 ASIG5V.n9394 0.019716
R57994 ASIG5V.n5998 ASIG5V.n5955 0.019716
R57995 ASIG5V.n6068 ASIG5V.n5997 0.019716
R57996 ASIG5V.n6068 ASIG5V.n5953 0.019716
R57997 ASIG5V.n6072 ASIG5V.n5996 0.019716
R57998 ASIG5V.n6072 ASIG5V.n5952 0.019716
R57999 ASIG5V.n6077 ASIG5V.n5995 0.019716
R58000 ASIG5V.n6077 ASIG5V.n5951 0.019716
R58001 ASIG5V.n6081 ASIG5V.n5994 0.019716
R58002 ASIG5V.n6081 ASIG5V.n5950 0.019716
R58003 ASIG5V.n6086 ASIG5V.n5993 0.019716
R58004 ASIG5V.n6086 ASIG5V.n5949 0.019716
R58005 ASIG5V.n6090 ASIG5V.n5992 0.019716
R58006 ASIG5V.n6090 ASIG5V.n5948 0.019716
R58007 ASIG5V.n6095 ASIG5V.n5991 0.019716
R58008 ASIG5V.n6095 ASIG5V.n5947 0.019716
R58009 ASIG5V.n6099 ASIG5V.n5990 0.019716
R58010 ASIG5V.n6099 ASIG5V.n5946 0.019716
R58011 ASIG5V.n6104 ASIG5V.n5989 0.019716
R58012 ASIG5V.n6104 ASIG5V.n5945 0.019716
R58013 ASIG5V.n6108 ASIG5V.n5988 0.019716
R58014 ASIG5V.n6108 ASIG5V.n5944 0.019716
R58015 ASIG5V.n6113 ASIG5V.n5987 0.019716
R58016 ASIG5V.n6113 ASIG5V.n5943 0.019716
R58017 ASIG5V.n6117 ASIG5V.n5986 0.019716
R58018 ASIG5V.n6117 ASIG5V.n5942 0.019716
R58019 ASIG5V.n6122 ASIG5V.n5985 0.019716
R58020 ASIG5V.n6122 ASIG5V.n5941 0.019716
R58021 ASIG5V.n6126 ASIG5V.n5984 0.019716
R58022 ASIG5V.n6126 ASIG5V.n5940 0.019716
R58023 ASIG5V.n6131 ASIG5V.n5983 0.019716
R58024 ASIG5V.n6131 ASIG5V.n5939 0.019716
R58025 ASIG5V.n6135 ASIG5V.n5982 0.019716
R58026 ASIG5V.n6135 ASIG5V.n5938 0.019716
R58027 ASIG5V.n6140 ASIG5V.n5981 0.019716
R58028 ASIG5V.n6140 ASIG5V.n5937 0.019716
R58029 ASIG5V.n6144 ASIG5V.n5980 0.019716
R58030 ASIG5V.n6144 ASIG5V.n5936 0.019716
R58031 ASIG5V.n6149 ASIG5V.n5979 0.019716
R58032 ASIG5V.n6149 ASIG5V.n5935 0.019716
R58033 ASIG5V.n6153 ASIG5V.n5978 0.019716
R58034 ASIG5V.n6153 ASIG5V.n5934 0.019716
R58035 ASIG5V.n6158 ASIG5V.n5977 0.019716
R58036 ASIG5V.n6158 ASIG5V.n5933 0.019716
R58037 ASIG5V.n6162 ASIG5V.n5976 0.019716
R58038 ASIG5V.n6162 ASIG5V.n5932 0.019716
R58039 ASIG5V.n6167 ASIG5V.n5975 0.019716
R58040 ASIG5V.n6167 ASIG5V.n5931 0.019716
R58041 ASIG5V.n6171 ASIG5V.n5974 0.019716
R58042 ASIG5V.n6171 ASIG5V.n5930 0.019716
R58043 ASIG5V.n6176 ASIG5V.n5973 0.019716
R58044 ASIG5V.n6176 ASIG5V.n5929 0.019716
R58045 ASIG5V.n6180 ASIG5V.n5972 0.019716
R58046 ASIG5V.n6180 ASIG5V.n5928 0.019716
R58047 ASIG5V.n6185 ASIG5V.n5971 0.019716
R58048 ASIG5V.n6185 ASIG5V.n5927 0.019716
R58049 ASIG5V.n6189 ASIG5V.n5970 0.019716
R58050 ASIG5V.n6189 ASIG5V.n5926 0.019716
R58051 ASIG5V.n6194 ASIG5V.n5969 0.019716
R58052 ASIG5V.n6194 ASIG5V.n5925 0.019716
R58053 ASIG5V.n6198 ASIG5V.n5968 0.019716
R58054 ASIG5V.n6198 ASIG5V.n5924 0.019716
R58055 ASIG5V.n6203 ASIG5V.n5967 0.019716
R58056 ASIG5V.n6203 ASIG5V.n5923 0.019716
R58057 ASIG5V.n6207 ASIG5V.n5966 0.019716
R58058 ASIG5V.n6207 ASIG5V.n5922 0.019716
R58059 ASIG5V.n6212 ASIG5V.n5965 0.019716
R58060 ASIG5V.n6212 ASIG5V.n5921 0.019716
R58061 ASIG5V.n6216 ASIG5V.n5964 0.019716
R58062 ASIG5V.n6216 ASIG5V.n5920 0.019716
R58063 ASIG5V.n6221 ASIG5V.n5963 0.019716
R58064 ASIG5V.n6221 ASIG5V.n5919 0.019716
R58065 ASIG5V.n6225 ASIG5V.n5962 0.019716
R58066 ASIG5V.n6225 ASIG5V.n5918 0.019716
R58067 ASIG5V.n6230 ASIG5V.n5961 0.019716
R58068 ASIG5V.n6230 ASIG5V.n5917 0.019716
R58069 ASIG5V.n6234 ASIG5V.n5960 0.019716
R58070 ASIG5V.n6234 ASIG5V.n5916 0.019716
R58071 ASIG5V.n6239 ASIG5V.n5959 0.019716
R58072 ASIG5V.n6239 ASIG5V.n5915 0.019716
R58073 ASIG5V.n6243 ASIG5V.n5958 0.019716
R58074 ASIG5V.n6243 ASIG5V.n5914 0.019716
R58075 ASIG5V.n9392 ASIG5V.n5913 0.019716
R58076 ASIG5V.n5905 ASIG5V.n5904 0.019716
R58077 ASIG5V.n5903 ASIG5V.n5902 0.019716
R58078 ASIG5V.n5580 ASIG5V.n5579 0.019716
R58079 ASIG5V.n5579 ASIG5V.n5575 0.019716
R58080 ASIG5V.n5893 ASIG5V.n5892 0.019716
R58081 ASIG5V.n5894 ASIG5V.n5893 0.019716
R58082 ASIG5V.n5586 ASIG5V.n5585 0.019716
R58083 ASIG5V.n5585 ASIG5V.n5581 0.019716
R58084 ASIG5V.n5883 ASIG5V.n5882 0.019716
R58085 ASIG5V.n5884 ASIG5V.n5883 0.019716
R58086 ASIG5V.n5592 ASIG5V.n5591 0.019716
R58087 ASIG5V.n5591 ASIG5V.n5587 0.019716
R58088 ASIG5V.n5873 ASIG5V.n5872 0.019716
R58089 ASIG5V.n5874 ASIG5V.n5873 0.019716
R58090 ASIG5V.n5598 ASIG5V.n5597 0.019716
R58091 ASIG5V.n5597 ASIG5V.n5593 0.019716
R58092 ASIG5V.n5863 ASIG5V.n5862 0.019716
R58093 ASIG5V.n5864 ASIG5V.n5863 0.019716
R58094 ASIG5V.n5604 ASIG5V.n5603 0.019716
R58095 ASIG5V.n5603 ASIG5V.n5599 0.019716
R58096 ASIG5V.n5853 ASIG5V.n5852 0.019716
R58097 ASIG5V.n5854 ASIG5V.n5853 0.019716
R58098 ASIG5V.n5610 ASIG5V.n5609 0.019716
R58099 ASIG5V.n5609 ASIG5V.n5605 0.019716
R58100 ASIG5V.n5843 ASIG5V.n5842 0.019716
R58101 ASIG5V.n5844 ASIG5V.n5843 0.019716
R58102 ASIG5V.n5616 ASIG5V.n5615 0.019716
R58103 ASIG5V.n5615 ASIG5V.n5611 0.019716
R58104 ASIG5V.n5833 ASIG5V.n5832 0.019716
R58105 ASIG5V.n5834 ASIG5V.n5833 0.019716
R58106 ASIG5V.n5622 ASIG5V.n5621 0.019716
R58107 ASIG5V.n5621 ASIG5V.n5617 0.019716
R58108 ASIG5V.n5823 ASIG5V.n5822 0.019716
R58109 ASIG5V.n5824 ASIG5V.n5823 0.019716
R58110 ASIG5V.n5628 ASIG5V.n5627 0.019716
R58111 ASIG5V.n5627 ASIG5V.n5623 0.019716
R58112 ASIG5V.n5813 ASIG5V.n5812 0.019716
R58113 ASIG5V.n5814 ASIG5V.n5813 0.019716
R58114 ASIG5V.n5634 ASIG5V.n5633 0.019716
R58115 ASIG5V.n5633 ASIG5V.n5629 0.019716
R58116 ASIG5V.n5803 ASIG5V.n5802 0.019716
R58117 ASIG5V.n5804 ASIG5V.n5803 0.019716
R58118 ASIG5V.n5640 ASIG5V.n5639 0.019716
R58119 ASIG5V.n5639 ASIG5V.n5635 0.019716
R58120 ASIG5V.n5793 ASIG5V.n5792 0.019716
R58121 ASIG5V.n5794 ASIG5V.n5793 0.019716
R58122 ASIG5V.n5646 ASIG5V.n5645 0.019716
R58123 ASIG5V.n5645 ASIG5V.n5641 0.019716
R58124 ASIG5V.n5783 ASIG5V.n5782 0.019716
R58125 ASIG5V.n5784 ASIG5V.n5783 0.019716
R58126 ASIG5V.n5652 ASIG5V.n5651 0.019716
R58127 ASIG5V.n5651 ASIG5V.n5647 0.019716
R58128 ASIG5V.n5773 ASIG5V.n5772 0.019716
R58129 ASIG5V.n5774 ASIG5V.n5773 0.019716
R58130 ASIG5V.n5658 ASIG5V.n5657 0.019716
R58131 ASIG5V.n5657 ASIG5V.n5653 0.019716
R58132 ASIG5V.n5763 ASIG5V.n5762 0.019716
R58133 ASIG5V.n5764 ASIG5V.n5763 0.019716
R58134 ASIG5V.n5664 ASIG5V.n5663 0.019716
R58135 ASIG5V.n5663 ASIG5V.n5659 0.019716
R58136 ASIG5V.n5753 ASIG5V.n5752 0.019716
R58137 ASIG5V.n5754 ASIG5V.n5753 0.019716
R58138 ASIG5V.n5670 ASIG5V.n5669 0.019716
R58139 ASIG5V.n5669 ASIG5V.n5665 0.019716
R58140 ASIG5V.n5743 ASIG5V.n5742 0.019716
R58141 ASIG5V.n5744 ASIG5V.n5743 0.019716
R58142 ASIG5V.n5676 ASIG5V.n5675 0.019716
R58143 ASIG5V.n5675 ASIG5V.n5671 0.019716
R58144 ASIG5V.n5733 ASIG5V.n5732 0.019716
R58145 ASIG5V.n5734 ASIG5V.n5733 0.019716
R58146 ASIG5V.n5682 ASIG5V.n5681 0.019716
R58147 ASIG5V.n5681 ASIG5V.n5677 0.019716
R58148 ASIG5V.n5723 ASIG5V.n5722 0.019716
R58149 ASIG5V.n5724 ASIG5V.n5723 0.019716
R58150 ASIG5V.n5688 ASIG5V.n5687 0.019716
R58151 ASIG5V.n5687 ASIG5V.n5683 0.019716
R58152 ASIG5V.n5713 ASIG5V.n5712 0.019716
R58153 ASIG5V.n5714 ASIG5V.n5713 0.019716
R58154 ASIG5V.n5694 ASIG5V.n5693 0.019716
R58155 ASIG5V.n5693 ASIG5V.n5689 0.019716
R58156 ASIG5V.n5703 ASIG5V.n5702 0.019716
R58157 ASIG5V.n5704 ASIG5V.n5703 0.019716
R58158 ASIG5V.n5696 ASIG5V.n5695 0.019716
R58159 ASIG5V.n9418 ASIG5V.n9417 0.019716
R58160 ASIG5V.n5552 ASIG5V.n5507 0.019716
R58161 ASIG5V.n7954 ASIG5V.n5551 0.019716
R58162 ASIG5V.n7954 ASIG5V.n5505 0.019716
R58163 ASIG5V.n7949 ASIG5V.n5550 0.019716
R58164 ASIG5V.n7949 ASIG5V.n5504 0.019716
R58165 ASIG5V.n7945 ASIG5V.n5549 0.019716
R58166 ASIG5V.n7945 ASIG5V.n5503 0.019716
R58167 ASIG5V.n7940 ASIG5V.n5548 0.019716
R58168 ASIG5V.n7940 ASIG5V.n5502 0.019716
R58169 ASIG5V.n7936 ASIG5V.n5547 0.019716
R58170 ASIG5V.n7936 ASIG5V.n5501 0.019716
R58171 ASIG5V.n7931 ASIG5V.n5546 0.019716
R58172 ASIG5V.n7931 ASIG5V.n5500 0.019716
R58173 ASIG5V.n7927 ASIG5V.n5545 0.019716
R58174 ASIG5V.n7927 ASIG5V.n5499 0.019716
R58175 ASIG5V.n7922 ASIG5V.n5544 0.019716
R58176 ASIG5V.n7922 ASIG5V.n5498 0.019716
R58177 ASIG5V.n7918 ASIG5V.n5543 0.019716
R58178 ASIG5V.n7918 ASIG5V.n5497 0.019716
R58179 ASIG5V.n7913 ASIG5V.n5542 0.019716
R58180 ASIG5V.n7913 ASIG5V.n5496 0.019716
R58181 ASIG5V.n7909 ASIG5V.n5541 0.019716
R58182 ASIG5V.n7909 ASIG5V.n5495 0.019716
R58183 ASIG5V.n7904 ASIG5V.n5540 0.019716
R58184 ASIG5V.n7904 ASIG5V.n5494 0.019716
R58185 ASIG5V.n7900 ASIG5V.n5539 0.019716
R58186 ASIG5V.n7900 ASIG5V.n5493 0.019716
R58187 ASIG5V.n7895 ASIG5V.n5538 0.019716
R58188 ASIG5V.n7895 ASIG5V.n5492 0.019716
R58189 ASIG5V.n7891 ASIG5V.n5537 0.019716
R58190 ASIG5V.n7891 ASIG5V.n5491 0.019716
R58191 ASIG5V.n7886 ASIG5V.n5536 0.019716
R58192 ASIG5V.n7886 ASIG5V.n5490 0.019716
R58193 ASIG5V.n7882 ASIG5V.n5535 0.019716
R58194 ASIG5V.n7882 ASIG5V.n5489 0.019716
R58195 ASIG5V.n7877 ASIG5V.n5534 0.019716
R58196 ASIG5V.n7877 ASIG5V.n5488 0.019716
R58197 ASIG5V.n7873 ASIG5V.n5533 0.019716
R58198 ASIG5V.n7873 ASIG5V.n5487 0.019716
R58199 ASIG5V.n7868 ASIG5V.n5532 0.019716
R58200 ASIG5V.n7868 ASIG5V.n5486 0.019716
R58201 ASIG5V.n7864 ASIG5V.n5531 0.019716
R58202 ASIG5V.n7864 ASIG5V.n5485 0.019716
R58203 ASIG5V.n7859 ASIG5V.n5530 0.019716
R58204 ASIG5V.n7859 ASIG5V.n5484 0.019716
R58205 ASIG5V.n7855 ASIG5V.n5529 0.019716
R58206 ASIG5V.n7855 ASIG5V.n5483 0.019716
R58207 ASIG5V.n7850 ASIG5V.n5528 0.019716
R58208 ASIG5V.n7850 ASIG5V.n5482 0.019716
R58209 ASIG5V.n7846 ASIG5V.n5527 0.019716
R58210 ASIG5V.n7846 ASIG5V.n5481 0.019716
R58211 ASIG5V.n7841 ASIG5V.n5526 0.019716
R58212 ASIG5V.n7841 ASIG5V.n5480 0.019716
R58213 ASIG5V.n7837 ASIG5V.n5525 0.019716
R58214 ASIG5V.n7837 ASIG5V.n5479 0.019716
R58215 ASIG5V.n7832 ASIG5V.n5524 0.019716
R58216 ASIG5V.n7832 ASIG5V.n5478 0.019716
R58217 ASIG5V.n7828 ASIG5V.n5523 0.019716
R58218 ASIG5V.n7828 ASIG5V.n5477 0.019716
R58219 ASIG5V.n7823 ASIG5V.n5522 0.019716
R58220 ASIG5V.n7823 ASIG5V.n5476 0.019716
R58221 ASIG5V.n7819 ASIG5V.n5521 0.019716
R58222 ASIG5V.n7819 ASIG5V.n5475 0.019716
R58223 ASIG5V.n7814 ASIG5V.n5520 0.019716
R58224 ASIG5V.n7814 ASIG5V.n5474 0.019716
R58225 ASIG5V.n7810 ASIG5V.n5519 0.019716
R58226 ASIG5V.n7810 ASIG5V.n5473 0.019716
R58227 ASIG5V.n7805 ASIG5V.n5518 0.019716
R58228 ASIG5V.n7805 ASIG5V.n5472 0.019716
R58229 ASIG5V.n7801 ASIG5V.n5517 0.019716
R58230 ASIG5V.n7801 ASIG5V.n5471 0.019716
R58231 ASIG5V.n7796 ASIG5V.n5516 0.019716
R58232 ASIG5V.n7796 ASIG5V.n5470 0.019716
R58233 ASIG5V.n7792 ASIG5V.n5515 0.019716
R58234 ASIG5V.n7792 ASIG5V.n5469 0.019716
R58235 ASIG5V.n7787 ASIG5V.n5514 0.019716
R58236 ASIG5V.n7787 ASIG5V.n5468 0.019716
R58237 ASIG5V.n7783 ASIG5V.n5513 0.019716
R58238 ASIG5V.n7783 ASIG5V.n5467 0.019716
R58239 ASIG5V.n7778 ASIG5V.n5512 0.019716
R58240 ASIG5V.n7778 ASIG5V.n5466 0.019716
R58241 ASIG5V.n9415 ASIG5V.n5465 0.019716
R58242 ASIG5V.n5211 ASIG5V.n5165 0.019716
R58243 ASIG5V.n5212 ASIG5V.n5164 0.019716
R58244 ASIG5V.n5221 ASIG5V.n5163 0.019716
R58245 ASIG5V.n5221 ASIG5V.n5220 0.019716
R58246 ASIG5V.n5223 ASIG5V.n5162 0.019716
R58247 ASIG5V.n5224 ASIG5V.n5223 0.019716
R58248 ASIG5V.n5233 ASIG5V.n5161 0.019716
R58249 ASIG5V.n5233 ASIG5V.n5232 0.019716
R58250 ASIG5V.n5235 ASIG5V.n5160 0.019716
R58251 ASIG5V.n5236 ASIG5V.n5235 0.019716
R58252 ASIG5V.n5245 ASIG5V.n5159 0.019716
R58253 ASIG5V.n5245 ASIG5V.n5244 0.019716
R58254 ASIG5V.n5247 ASIG5V.n5158 0.019716
R58255 ASIG5V.n5248 ASIG5V.n5247 0.019716
R58256 ASIG5V.n5257 ASIG5V.n5157 0.019716
R58257 ASIG5V.n5257 ASIG5V.n5256 0.019716
R58258 ASIG5V.n5259 ASIG5V.n5156 0.019716
R58259 ASIG5V.n5260 ASIG5V.n5259 0.019716
R58260 ASIG5V.n5269 ASIG5V.n5155 0.019716
R58261 ASIG5V.n5269 ASIG5V.n5268 0.019716
R58262 ASIG5V.n5271 ASIG5V.n5154 0.019716
R58263 ASIG5V.n5272 ASIG5V.n5271 0.019716
R58264 ASIG5V.n5281 ASIG5V.n5153 0.019716
R58265 ASIG5V.n5281 ASIG5V.n5280 0.019716
R58266 ASIG5V.n5283 ASIG5V.n5152 0.019716
R58267 ASIG5V.n5284 ASIG5V.n5283 0.019716
R58268 ASIG5V.n5293 ASIG5V.n5151 0.019716
R58269 ASIG5V.n5293 ASIG5V.n5292 0.019716
R58270 ASIG5V.n5295 ASIG5V.n5150 0.019716
R58271 ASIG5V.n5296 ASIG5V.n5295 0.019716
R58272 ASIG5V.n5305 ASIG5V.n5149 0.019716
R58273 ASIG5V.n5305 ASIG5V.n5304 0.019716
R58274 ASIG5V.n5307 ASIG5V.n5148 0.019716
R58275 ASIG5V.n5308 ASIG5V.n5307 0.019716
R58276 ASIG5V.n5317 ASIG5V.n5147 0.019716
R58277 ASIG5V.n5317 ASIG5V.n5316 0.019716
R58278 ASIG5V.n5319 ASIG5V.n5146 0.019716
R58279 ASIG5V.n5320 ASIG5V.n5319 0.019716
R58280 ASIG5V.n5329 ASIG5V.n5145 0.019716
R58281 ASIG5V.n5329 ASIG5V.n5328 0.019716
R58282 ASIG5V.n5331 ASIG5V.n5144 0.019716
R58283 ASIG5V.n5332 ASIG5V.n5331 0.019716
R58284 ASIG5V.n5341 ASIG5V.n5143 0.019716
R58285 ASIG5V.n5341 ASIG5V.n5340 0.019716
R58286 ASIG5V.n5343 ASIG5V.n5142 0.019716
R58287 ASIG5V.n5344 ASIG5V.n5343 0.019716
R58288 ASIG5V.n5353 ASIG5V.n5141 0.019716
R58289 ASIG5V.n5353 ASIG5V.n5352 0.019716
R58290 ASIG5V.n5355 ASIG5V.n5140 0.019716
R58291 ASIG5V.n5356 ASIG5V.n5355 0.019716
R58292 ASIG5V.n5365 ASIG5V.n5139 0.019716
R58293 ASIG5V.n5365 ASIG5V.n5364 0.019716
R58294 ASIG5V.n5367 ASIG5V.n5138 0.019716
R58295 ASIG5V.n5368 ASIG5V.n5367 0.019716
R58296 ASIG5V.n5377 ASIG5V.n5137 0.019716
R58297 ASIG5V.n5377 ASIG5V.n5376 0.019716
R58298 ASIG5V.n5379 ASIG5V.n5136 0.019716
R58299 ASIG5V.n5380 ASIG5V.n5379 0.019716
R58300 ASIG5V.n5389 ASIG5V.n5135 0.019716
R58301 ASIG5V.n5389 ASIG5V.n5388 0.019716
R58302 ASIG5V.n5391 ASIG5V.n5134 0.019716
R58303 ASIG5V.n5392 ASIG5V.n5391 0.019716
R58304 ASIG5V.n5401 ASIG5V.n5133 0.019716
R58305 ASIG5V.n5401 ASIG5V.n5400 0.019716
R58306 ASIG5V.n5403 ASIG5V.n5132 0.019716
R58307 ASIG5V.n5404 ASIG5V.n5403 0.019716
R58308 ASIG5V.n5413 ASIG5V.n5131 0.019716
R58309 ASIG5V.n5413 ASIG5V.n5412 0.019716
R58310 ASIG5V.n5415 ASIG5V.n5130 0.019716
R58311 ASIG5V.n5416 ASIG5V.n5415 0.019716
R58312 ASIG5V.n5425 ASIG5V.n5129 0.019716
R58313 ASIG5V.n5425 ASIG5V.n5424 0.019716
R58314 ASIG5V.n5427 ASIG5V.n5128 0.019716
R58315 ASIG5V.n5428 ASIG5V.n5427 0.019716
R58316 ASIG5V.n5437 ASIG5V.n5127 0.019716
R58317 ASIG5V.n5437 ASIG5V.n5436 0.019716
R58318 ASIG5V.n5439 ASIG5V.n5126 0.019716
R58319 ASIG5V.n5440 ASIG5V.n5439 0.019716
R58320 ASIG5V.n5449 ASIG5V.n5125 0.019716
R58321 ASIG5V.n5449 ASIG5V.n5448 0.019716
R58322 ASIG5V.n5451 ASIG5V.n5124 0.019716
R58323 ASIG5V.n5452 ASIG5V.n5451 0.019716
R58324 ASIG5V.n9431 ASIG5V.n9430 0.019716
R58325 ASIG5V.n9483 ASIG5V.n5116 0.019716
R58326 ASIG5V.n9484 ASIG5V.n5115 0.019716
R58327 ASIG5V.n9493 ASIG5V.n5114 0.019716
R58328 ASIG5V.n9493 ASIG5V.n9492 0.019716
R58329 ASIG5V.n9495 ASIG5V.n5113 0.019716
R58330 ASIG5V.n9496 ASIG5V.n9495 0.019716
R58331 ASIG5V.n9505 ASIG5V.n5112 0.019716
R58332 ASIG5V.n9505 ASIG5V.n9504 0.019716
R58333 ASIG5V.n9507 ASIG5V.n5111 0.019716
R58334 ASIG5V.n9508 ASIG5V.n9507 0.019716
R58335 ASIG5V.n9517 ASIG5V.n5110 0.019716
R58336 ASIG5V.n9517 ASIG5V.n9516 0.019716
R58337 ASIG5V.n9519 ASIG5V.n5109 0.019716
R58338 ASIG5V.n9520 ASIG5V.n9519 0.019716
R58339 ASIG5V.n9529 ASIG5V.n5108 0.019716
R58340 ASIG5V.n9529 ASIG5V.n9528 0.019716
R58341 ASIG5V.n9531 ASIG5V.n5107 0.019716
R58342 ASIG5V.n9532 ASIG5V.n9531 0.019716
R58343 ASIG5V.n9541 ASIG5V.n5106 0.019716
R58344 ASIG5V.n9541 ASIG5V.n9540 0.019716
R58345 ASIG5V.n9543 ASIG5V.n5105 0.019716
R58346 ASIG5V.n9544 ASIG5V.n9543 0.019716
R58347 ASIG5V.n9553 ASIG5V.n5104 0.019716
R58348 ASIG5V.n9553 ASIG5V.n9552 0.019716
R58349 ASIG5V.n9555 ASIG5V.n5103 0.019716
R58350 ASIG5V.n9556 ASIG5V.n9555 0.019716
R58351 ASIG5V.n9565 ASIG5V.n5102 0.019716
R58352 ASIG5V.n9565 ASIG5V.n9564 0.019716
R58353 ASIG5V.n9567 ASIG5V.n5101 0.019716
R58354 ASIG5V.n9568 ASIG5V.n9567 0.019716
R58355 ASIG5V.n9577 ASIG5V.n5100 0.019716
R58356 ASIG5V.n9577 ASIG5V.n9576 0.019716
R58357 ASIG5V.n9579 ASIG5V.n5099 0.019716
R58358 ASIG5V.n9580 ASIG5V.n9579 0.019716
R58359 ASIG5V.n9589 ASIG5V.n5098 0.019716
R58360 ASIG5V.n9589 ASIG5V.n9588 0.019716
R58361 ASIG5V.n9591 ASIG5V.n5097 0.019716
R58362 ASIG5V.n9592 ASIG5V.n9591 0.019716
R58363 ASIG5V.n9601 ASIG5V.n5096 0.019716
R58364 ASIG5V.n9601 ASIG5V.n9600 0.019716
R58365 ASIG5V.n9603 ASIG5V.n5095 0.019716
R58366 ASIG5V.n9604 ASIG5V.n9603 0.019716
R58367 ASIG5V.n9613 ASIG5V.n5094 0.019716
R58368 ASIG5V.n9613 ASIG5V.n9612 0.019716
R58369 ASIG5V.n9615 ASIG5V.n5093 0.019716
R58370 ASIG5V.n9616 ASIG5V.n9615 0.019716
R58371 ASIG5V.n9625 ASIG5V.n5092 0.019716
R58372 ASIG5V.n9625 ASIG5V.n9624 0.019716
R58373 ASIG5V.n9627 ASIG5V.n5091 0.019716
R58374 ASIG5V.n9628 ASIG5V.n9627 0.019716
R58375 ASIG5V.n9637 ASIG5V.n5090 0.019716
R58376 ASIG5V.n9637 ASIG5V.n9636 0.019716
R58377 ASIG5V.n9639 ASIG5V.n5089 0.019716
R58378 ASIG5V.n9640 ASIG5V.n9639 0.019716
R58379 ASIG5V.n9649 ASIG5V.n5088 0.019716
R58380 ASIG5V.n9649 ASIG5V.n9648 0.019716
R58381 ASIG5V.n9651 ASIG5V.n5087 0.019716
R58382 ASIG5V.n9652 ASIG5V.n9651 0.019716
R58383 ASIG5V.n9661 ASIG5V.n5086 0.019716
R58384 ASIG5V.n9661 ASIG5V.n9660 0.019716
R58385 ASIG5V.n9663 ASIG5V.n5085 0.019716
R58386 ASIG5V.n9664 ASIG5V.n9663 0.019716
R58387 ASIG5V.n9673 ASIG5V.n5084 0.019716
R58388 ASIG5V.n9673 ASIG5V.n9672 0.019716
R58389 ASIG5V.n9675 ASIG5V.n5083 0.019716
R58390 ASIG5V.n9676 ASIG5V.n9675 0.019716
R58391 ASIG5V.n9685 ASIG5V.n5082 0.019716
R58392 ASIG5V.n9685 ASIG5V.n9684 0.019716
R58393 ASIG5V.n9687 ASIG5V.n5081 0.019716
R58394 ASIG5V.n9688 ASIG5V.n9687 0.019716
R58395 ASIG5V.n9697 ASIG5V.n5080 0.019716
R58396 ASIG5V.n9697 ASIG5V.n9696 0.019716
R58397 ASIG5V.n9699 ASIG5V.n5079 0.019716
R58398 ASIG5V.n9700 ASIG5V.n9699 0.019716
R58399 ASIG5V.n9709 ASIG5V.n5078 0.019716
R58400 ASIG5V.n9709 ASIG5V.n9708 0.019716
R58401 ASIG5V.n9711 ASIG5V.n5077 0.019716
R58402 ASIG5V.n9712 ASIG5V.n9711 0.019716
R58403 ASIG5V.n9721 ASIG5V.n5076 0.019716
R58404 ASIG5V.n9721 ASIG5V.n9720 0.019716
R58405 ASIG5V.n9723 ASIG5V.n5075 0.019716
R58406 ASIG5V.n9724 ASIG5V.n9723 0.019716
R58407 ASIG5V.n9733 ASIG5V.n9732 0.019716
R58408 ASIG5V.n3264 ASIG5V.n3220 0.019716
R58409 ASIG5V.n3265 ASIG5V.n3219 0.019716
R58410 ASIG5V.n4822 ASIG5V.n3218 0.019716
R58411 ASIG5V.n4822 ASIG5V.n4821 0.019716
R58412 ASIG5V.n4824 ASIG5V.n3217 0.019716
R58413 ASIG5V.n4825 ASIG5V.n4824 0.019716
R58414 ASIG5V.n4834 ASIG5V.n3216 0.019716
R58415 ASIG5V.n4834 ASIG5V.n4833 0.019716
R58416 ASIG5V.n4836 ASIG5V.n3215 0.019716
R58417 ASIG5V.n4837 ASIG5V.n4836 0.019716
R58418 ASIG5V.n4846 ASIG5V.n3214 0.019716
R58419 ASIG5V.n4846 ASIG5V.n4845 0.019716
R58420 ASIG5V.n4848 ASIG5V.n3213 0.019716
R58421 ASIG5V.n4849 ASIG5V.n4848 0.019716
R58422 ASIG5V.n4858 ASIG5V.n3212 0.019716
R58423 ASIG5V.n4858 ASIG5V.n4857 0.019716
R58424 ASIG5V.n4860 ASIG5V.n3211 0.019716
R58425 ASIG5V.n4861 ASIG5V.n4860 0.019716
R58426 ASIG5V.n4870 ASIG5V.n3210 0.019716
R58427 ASIG5V.n4870 ASIG5V.n4869 0.019716
R58428 ASIG5V.n4872 ASIG5V.n3209 0.019716
R58429 ASIG5V.n4873 ASIG5V.n4872 0.019716
R58430 ASIG5V.n4882 ASIG5V.n3208 0.019716
R58431 ASIG5V.n4882 ASIG5V.n4881 0.019716
R58432 ASIG5V.n4884 ASIG5V.n3207 0.019716
R58433 ASIG5V.n4885 ASIG5V.n4884 0.019716
R58434 ASIG5V.n4894 ASIG5V.n3206 0.019716
R58435 ASIG5V.n4894 ASIG5V.n4893 0.019716
R58436 ASIG5V.n4896 ASIG5V.n3205 0.019716
R58437 ASIG5V.n4897 ASIG5V.n4896 0.019716
R58438 ASIG5V.n4906 ASIG5V.n3204 0.019716
R58439 ASIG5V.n4906 ASIG5V.n4905 0.019716
R58440 ASIG5V.n4908 ASIG5V.n3203 0.019716
R58441 ASIG5V.n4909 ASIG5V.n4908 0.019716
R58442 ASIG5V.n4918 ASIG5V.n3202 0.019716
R58443 ASIG5V.n4918 ASIG5V.n4917 0.019716
R58444 ASIG5V.n4920 ASIG5V.n3201 0.019716
R58445 ASIG5V.n4921 ASIG5V.n4920 0.019716
R58446 ASIG5V.n4930 ASIG5V.n3200 0.019716
R58447 ASIG5V.n4930 ASIG5V.n4929 0.019716
R58448 ASIG5V.n4932 ASIG5V.n3199 0.019716
R58449 ASIG5V.n4933 ASIG5V.n4932 0.019716
R58450 ASIG5V.n4942 ASIG5V.n3198 0.019716
R58451 ASIG5V.n4942 ASIG5V.n4941 0.019716
R58452 ASIG5V.n4944 ASIG5V.n3197 0.019716
R58453 ASIG5V.n4945 ASIG5V.n4944 0.019716
R58454 ASIG5V.n4954 ASIG5V.n3196 0.019716
R58455 ASIG5V.n4954 ASIG5V.n4953 0.019716
R58456 ASIG5V.n4956 ASIG5V.n3195 0.019716
R58457 ASIG5V.n4957 ASIG5V.n4956 0.019716
R58458 ASIG5V.n4966 ASIG5V.n3194 0.019716
R58459 ASIG5V.n4966 ASIG5V.n4965 0.019716
R58460 ASIG5V.n4968 ASIG5V.n3193 0.019716
R58461 ASIG5V.n4969 ASIG5V.n4968 0.019716
R58462 ASIG5V.n4978 ASIG5V.n3192 0.019716
R58463 ASIG5V.n4978 ASIG5V.n4977 0.019716
R58464 ASIG5V.n4980 ASIG5V.n3191 0.019716
R58465 ASIG5V.n4981 ASIG5V.n4980 0.019716
R58466 ASIG5V.n4990 ASIG5V.n3190 0.019716
R58467 ASIG5V.n4990 ASIG5V.n4989 0.019716
R58468 ASIG5V.n4992 ASIG5V.n3189 0.019716
R58469 ASIG5V.n4993 ASIG5V.n4992 0.019716
R58470 ASIG5V.n5002 ASIG5V.n3188 0.019716
R58471 ASIG5V.n5002 ASIG5V.n5001 0.019716
R58472 ASIG5V.n5004 ASIG5V.n3187 0.019716
R58473 ASIG5V.n5005 ASIG5V.n5004 0.019716
R58474 ASIG5V.n5014 ASIG5V.n3186 0.019716
R58475 ASIG5V.n5014 ASIG5V.n5013 0.019716
R58476 ASIG5V.n5016 ASIG5V.n3185 0.019716
R58477 ASIG5V.n5017 ASIG5V.n5016 0.019716
R58478 ASIG5V.n5026 ASIG5V.n3184 0.019716
R58479 ASIG5V.n5026 ASIG5V.n5025 0.019716
R58480 ASIG5V.n5028 ASIG5V.n3183 0.019716
R58481 ASIG5V.n5029 ASIG5V.n5028 0.019716
R58482 ASIG5V.n5038 ASIG5V.n3182 0.019716
R58483 ASIG5V.n5038 ASIG5V.n5037 0.019716
R58484 ASIG5V.n5040 ASIG5V.n3181 0.019716
R58485 ASIG5V.n5041 ASIG5V.n5040 0.019716
R58486 ASIG5V.n5050 ASIG5V.n3180 0.019716
R58487 ASIG5V.n5050 ASIG5V.n5049 0.019716
R58488 ASIG5V.n5052 ASIG5V.n3179 0.019716
R58489 ASIG5V.n5053 ASIG5V.n5052 0.019716
R58490 ASIG5V.n5063 ASIG5V.n5062 0.019716
R58491 ASIG5V.n3614 ASIG5V.n3613 0.019716
R58492 ASIG5V.n3612 ASIG5V.n3611 0.019716
R58493 ASIG5V.n3289 ASIG5V.n3288 0.019716
R58494 ASIG5V.n3288 ASIG5V.n3284 0.019716
R58495 ASIG5V.n3602 ASIG5V.n3601 0.019716
R58496 ASIG5V.n3603 ASIG5V.n3602 0.019716
R58497 ASIG5V.n3295 ASIG5V.n3294 0.019716
R58498 ASIG5V.n3294 ASIG5V.n3290 0.019716
R58499 ASIG5V.n3592 ASIG5V.n3591 0.019716
R58500 ASIG5V.n3593 ASIG5V.n3592 0.019716
R58501 ASIG5V.n3301 ASIG5V.n3300 0.019716
R58502 ASIG5V.n3300 ASIG5V.n3296 0.019716
R58503 ASIG5V.n3582 ASIG5V.n3581 0.019716
R58504 ASIG5V.n3583 ASIG5V.n3582 0.019716
R58505 ASIG5V.n3307 ASIG5V.n3306 0.019716
R58506 ASIG5V.n3306 ASIG5V.n3302 0.019716
R58507 ASIG5V.n3572 ASIG5V.n3571 0.019716
R58508 ASIG5V.n3573 ASIG5V.n3572 0.019716
R58509 ASIG5V.n3313 ASIG5V.n3312 0.019716
R58510 ASIG5V.n3312 ASIG5V.n3308 0.019716
R58511 ASIG5V.n3562 ASIG5V.n3561 0.019716
R58512 ASIG5V.n3563 ASIG5V.n3562 0.019716
R58513 ASIG5V.n3319 ASIG5V.n3318 0.019716
R58514 ASIG5V.n3318 ASIG5V.n3314 0.019716
R58515 ASIG5V.n3552 ASIG5V.n3551 0.019716
R58516 ASIG5V.n3553 ASIG5V.n3552 0.019716
R58517 ASIG5V.n3325 ASIG5V.n3324 0.019716
R58518 ASIG5V.n3324 ASIG5V.n3320 0.019716
R58519 ASIG5V.n3542 ASIG5V.n3541 0.019716
R58520 ASIG5V.n3543 ASIG5V.n3542 0.019716
R58521 ASIG5V.n3331 ASIG5V.n3330 0.019716
R58522 ASIG5V.n3330 ASIG5V.n3326 0.019716
R58523 ASIG5V.n3532 ASIG5V.n3531 0.019716
R58524 ASIG5V.n3533 ASIG5V.n3532 0.019716
R58525 ASIG5V.n3337 ASIG5V.n3336 0.019716
R58526 ASIG5V.n3336 ASIG5V.n3332 0.019716
R58527 ASIG5V.n3522 ASIG5V.n3521 0.019716
R58528 ASIG5V.n3523 ASIG5V.n3522 0.019716
R58529 ASIG5V.n3343 ASIG5V.n3342 0.019716
R58530 ASIG5V.n3342 ASIG5V.n3338 0.019716
R58531 ASIG5V.n3512 ASIG5V.n3511 0.019716
R58532 ASIG5V.n3513 ASIG5V.n3512 0.019716
R58533 ASIG5V.n3349 ASIG5V.n3348 0.019716
R58534 ASIG5V.n3348 ASIG5V.n3344 0.019716
R58535 ASIG5V.n3502 ASIG5V.n3501 0.019716
R58536 ASIG5V.n3503 ASIG5V.n3502 0.019716
R58537 ASIG5V.n3355 ASIG5V.n3354 0.019716
R58538 ASIG5V.n3354 ASIG5V.n3350 0.019716
R58539 ASIG5V.n3492 ASIG5V.n3491 0.019716
R58540 ASIG5V.n3493 ASIG5V.n3492 0.019716
R58541 ASIG5V.n3361 ASIG5V.n3360 0.019716
R58542 ASIG5V.n3360 ASIG5V.n3356 0.019716
R58543 ASIG5V.n3482 ASIG5V.n3481 0.019716
R58544 ASIG5V.n3483 ASIG5V.n3482 0.019716
R58545 ASIG5V.n3367 ASIG5V.n3366 0.019716
R58546 ASIG5V.n3366 ASIG5V.n3362 0.019716
R58547 ASIG5V.n3472 ASIG5V.n3471 0.019716
R58548 ASIG5V.n3473 ASIG5V.n3472 0.019716
R58549 ASIG5V.n3373 ASIG5V.n3372 0.019716
R58550 ASIG5V.n3372 ASIG5V.n3368 0.019716
R58551 ASIG5V.n3462 ASIG5V.n3461 0.019716
R58552 ASIG5V.n3463 ASIG5V.n3462 0.019716
R58553 ASIG5V.n3379 ASIG5V.n3378 0.019716
R58554 ASIG5V.n3378 ASIG5V.n3374 0.019716
R58555 ASIG5V.n3452 ASIG5V.n3451 0.019716
R58556 ASIG5V.n3453 ASIG5V.n3452 0.019716
R58557 ASIG5V.n3385 ASIG5V.n3384 0.019716
R58558 ASIG5V.n3384 ASIG5V.n3380 0.019716
R58559 ASIG5V.n3442 ASIG5V.n3441 0.019716
R58560 ASIG5V.n3443 ASIG5V.n3442 0.019716
R58561 ASIG5V.n3391 ASIG5V.n3390 0.019716
R58562 ASIG5V.n3390 ASIG5V.n3386 0.019716
R58563 ASIG5V.n3432 ASIG5V.n3431 0.019716
R58564 ASIG5V.n3433 ASIG5V.n3432 0.019716
R58565 ASIG5V.n3397 ASIG5V.n3396 0.019716
R58566 ASIG5V.n3396 ASIG5V.n3392 0.019716
R58567 ASIG5V.n3422 ASIG5V.n3421 0.019716
R58568 ASIG5V.n3423 ASIG5V.n3422 0.019716
R58569 ASIG5V.n3403 ASIG5V.n3402 0.019716
R58570 ASIG5V.n3402 ASIG5V.n3398 0.019716
R58571 ASIG5V.n3412 ASIG5V.n3411 0.019716
R58572 ASIG5V.n3413 ASIG5V.n3412 0.019716
R58573 ASIG5V.n3405 ASIG5V.n3404 0.019716
R58574 ASIG5V.n4774 ASIG5V.n3671 0.019716
R58575 ASIG5V.n3675 ASIG5V.n3671 0.019716
R58576 ASIG5V.n4590 ASIG5V.n3670 0.019716
R58577 ASIG5V.n4590 ASIG5V.n3676 0.019716
R58578 ASIG5V.n3773 ASIG5V.n3669 0.019716
R58579 ASIG5V.n3773 ASIG5V.n3677 0.019716
R58580 ASIG5V.n4599 ASIG5V.n3668 0.019716
R58581 ASIG5V.n4599 ASIG5V.n3678 0.019716
R58582 ASIG5V.n3770 ASIG5V.n3667 0.019716
R58583 ASIG5V.n3770 ASIG5V.n3679 0.019716
R58584 ASIG5V.n4608 ASIG5V.n3666 0.019716
R58585 ASIG5V.n4608 ASIG5V.n3680 0.019716
R58586 ASIG5V.n3767 ASIG5V.n3665 0.019716
R58587 ASIG5V.n3767 ASIG5V.n3681 0.019716
R58588 ASIG5V.n4617 ASIG5V.n3664 0.019716
R58589 ASIG5V.n4617 ASIG5V.n3682 0.019716
R58590 ASIG5V.n3764 ASIG5V.n3663 0.019716
R58591 ASIG5V.n3764 ASIG5V.n3683 0.019716
R58592 ASIG5V.n4626 ASIG5V.n3662 0.019716
R58593 ASIG5V.n4626 ASIG5V.n3684 0.019716
R58594 ASIG5V.n3761 ASIG5V.n3661 0.019716
R58595 ASIG5V.n3761 ASIG5V.n3685 0.019716
R58596 ASIG5V.n4635 ASIG5V.n3660 0.019716
R58597 ASIG5V.n4635 ASIG5V.n3686 0.019716
R58598 ASIG5V.n3758 ASIG5V.n3659 0.019716
R58599 ASIG5V.n3758 ASIG5V.n3687 0.019716
R58600 ASIG5V.n4644 ASIG5V.n3658 0.019716
R58601 ASIG5V.n4644 ASIG5V.n3688 0.019716
R58602 ASIG5V.n3755 ASIG5V.n3657 0.019716
R58603 ASIG5V.n3755 ASIG5V.n3689 0.019716
R58604 ASIG5V.n4653 ASIG5V.n3656 0.019716
R58605 ASIG5V.n4653 ASIG5V.n3690 0.019716
R58606 ASIG5V.n3752 ASIG5V.n3655 0.019716
R58607 ASIG5V.n3752 ASIG5V.n3691 0.019716
R58608 ASIG5V.n4662 ASIG5V.n3654 0.019716
R58609 ASIG5V.n4662 ASIG5V.n3692 0.019716
R58610 ASIG5V.n3749 ASIG5V.n3653 0.019716
R58611 ASIG5V.n3749 ASIG5V.n3693 0.019716
R58612 ASIG5V.n4671 ASIG5V.n3652 0.019716
R58613 ASIG5V.n4671 ASIG5V.n3694 0.019716
R58614 ASIG5V.n3746 ASIG5V.n3651 0.019716
R58615 ASIG5V.n3746 ASIG5V.n3695 0.019716
R58616 ASIG5V.n4680 ASIG5V.n3650 0.019716
R58617 ASIG5V.n4680 ASIG5V.n3696 0.019716
R58618 ASIG5V.n3743 ASIG5V.n3649 0.019716
R58619 ASIG5V.n3743 ASIG5V.n3697 0.019716
R58620 ASIG5V.n4689 ASIG5V.n3648 0.019716
R58621 ASIG5V.n4689 ASIG5V.n3698 0.019716
R58622 ASIG5V.n3740 ASIG5V.n3647 0.019716
R58623 ASIG5V.n3740 ASIG5V.n3699 0.019716
R58624 ASIG5V.n4698 ASIG5V.n3646 0.019716
R58625 ASIG5V.n4698 ASIG5V.n3700 0.019716
R58626 ASIG5V.n3737 ASIG5V.n3645 0.019716
R58627 ASIG5V.n3737 ASIG5V.n3701 0.019716
R58628 ASIG5V.n4707 ASIG5V.n3644 0.019716
R58629 ASIG5V.n4707 ASIG5V.n3702 0.019716
R58630 ASIG5V.n3734 ASIG5V.n3643 0.019716
R58631 ASIG5V.n3734 ASIG5V.n3703 0.019716
R58632 ASIG5V.n4716 ASIG5V.n3642 0.019716
R58633 ASIG5V.n4716 ASIG5V.n3704 0.019716
R58634 ASIG5V.n3731 ASIG5V.n3641 0.019716
R58635 ASIG5V.n3731 ASIG5V.n3705 0.019716
R58636 ASIG5V.n4725 ASIG5V.n3640 0.019716
R58637 ASIG5V.n4725 ASIG5V.n3706 0.019716
R58638 ASIG5V.n3728 ASIG5V.n3639 0.019716
R58639 ASIG5V.n3728 ASIG5V.n3707 0.019716
R58640 ASIG5V.n4734 ASIG5V.n3638 0.019716
R58641 ASIG5V.n4734 ASIG5V.n3708 0.019716
R58642 ASIG5V.n3725 ASIG5V.n3637 0.019716
R58643 ASIG5V.n3725 ASIG5V.n3709 0.019716
R58644 ASIG5V.n4743 ASIG5V.n3636 0.019716
R58645 ASIG5V.n4743 ASIG5V.n3710 0.019716
R58646 ASIG5V.n3722 ASIG5V.n3635 0.019716
R58647 ASIG5V.n3722 ASIG5V.n3711 0.019716
R58648 ASIG5V.n4752 ASIG5V.n3634 0.019716
R58649 ASIG5V.n4752 ASIG5V.n3712 0.019716
R58650 ASIG5V.n3719 ASIG5V.n3633 0.019716
R58651 ASIG5V.n3719 ASIG5V.n3713 0.019716
R58652 ASIG5V.n4761 ASIG5V.n3632 0.019716
R58653 ASIG5V.n4761 ASIG5V.n3714 0.019716
R58654 ASIG5V.n3716 ASIG5V.n3631 0.019716
R58655 ASIG5V.n3716 ASIG5V.n3715 0.019716
R58656 ASIG5V.n4771 ASIG5V.n3630 0.019716
R58657 ASIG5V.n4774 ASIG5V.n4773 0.019716
R58658 ASIG5V.n4588 ASIG5V.n3670 0.019716
R58659 ASIG5V.n4588 ASIG5V.n3675 0.019716
R58660 ASIG5V.n4592 ASIG5V.n3669 0.019716
R58661 ASIG5V.n4592 ASIG5V.n3676 0.019716
R58662 ASIG5V.n4597 ASIG5V.n3668 0.019716
R58663 ASIG5V.n4597 ASIG5V.n3677 0.019716
R58664 ASIG5V.n4601 ASIG5V.n3667 0.019716
R58665 ASIG5V.n4601 ASIG5V.n3678 0.019716
R58666 ASIG5V.n4606 ASIG5V.n3666 0.019716
R58667 ASIG5V.n4606 ASIG5V.n3679 0.019716
R58668 ASIG5V.n4610 ASIG5V.n3665 0.019716
R58669 ASIG5V.n4610 ASIG5V.n3680 0.019716
R58670 ASIG5V.n4615 ASIG5V.n3664 0.019716
R58671 ASIG5V.n4615 ASIG5V.n3681 0.019716
R58672 ASIG5V.n4619 ASIG5V.n3663 0.019716
R58673 ASIG5V.n4619 ASIG5V.n3682 0.019716
R58674 ASIG5V.n4624 ASIG5V.n3662 0.019716
R58675 ASIG5V.n4624 ASIG5V.n3683 0.019716
R58676 ASIG5V.n4628 ASIG5V.n3661 0.019716
R58677 ASIG5V.n4628 ASIG5V.n3684 0.019716
R58678 ASIG5V.n4633 ASIG5V.n3660 0.019716
R58679 ASIG5V.n4633 ASIG5V.n3685 0.019716
R58680 ASIG5V.n4637 ASIG5V.n3659 0.019716
R58681 ASIG5V.n4637 ASIG5V.n3686 0.019716
R58682 ASIG5V.n4642 ASIG5V.n3658 0.019716
R58683 ASIG5V.n4642 ASIG5V.n3687 0.019716
R58684 ASIG5V.n4646 ASIG5V.n3657 0.019716
R58685 ASIG5V.n4646 ASIG5V.n3688 0.019716
R58686 ASIG5V.n4651 ASIG5V.n3656 0.019716
R58687 ASIG5V.n4651 ASIG5V.n3689 0.019716
R58688 ASIG5V.n4655 ASIG5V.n3655 0.019716
R58689 ASIG5V.n4655 ASIG5V.n3690 0.019716
R58690 ASIG5V.n4660 ASIG5V.n3654 0.019716
R58691 ASIG5V.n4660 ASIG5V.n3691 0.019716
R58692 ASIG5V.n4664 ASIG5V.n3653 0.019716
R58693 ASIG5V.n4664 ASIG5V.n3692 0.019716
R58694 ASIG5V.n4669 ASIG5V.n3652 0.019716
R58695 ASIG5V.n4669 ASIG5V.n3693 0.019716
R58696 ASIG5V.n4673 ASIG5V.n3651 0.019716
R58697 ASIG5V.n4673 ASIG5V.n3694 0.019716
R58698 ASIG5V.n4678 ASIG5V.n3650 0.019716
R58699 ASIG5V.n4678 ASIG5V.n3695 0.019716
R58700 ASIG5V.n4682 ASIG5V.n3649 0.019716
R58701 ASIG5V.n4682 ASIG5V.n3696 0.019716
R58702 ASIG5V.n4687 ASIG5V.n3648 0.019716
R58703 ASIG5V.n4687 ASIG5V.n3697 0.019716
R58704 ASIG5V.n4691 ASIG5V.n3647 0.019716
R58705 ASIG5V.n4691 ASIG5V.n3698 0.019716
R58706 ASIG5V.n4696 ASIG5V.n3646 0.019716
R58707 ASIG5V.n4696 ASIG5V.n3699 0.019716
R58708 ASIG5V.n4700 ASIG5V.n3645 0.019716
R58709 ASIG5V.n4700 ASIG5V.n3700 0.019716
R58710 ASIG5V.n4705 ASIG5V.n3644 0.019716
R58711 ASIG5V.n4705 ASIG5V.n3701 0.019716
R58712 ASIG5V.n4709 ASIG5V.n3643 0.019716
R58713 ASIG5V.n4709 ASIG5V.n3702 0.019716
R58714 ASIG5V.n4714 ASIG5V.n3642 0.019716
R58715 ASIG5V.n4714 ASIG5V.n3703 0.019716
R58716 ASIG5V.n4718 ASIG5V.n3641 0.019716
R58717 ASIG5V.n4718 ASIG5V.n3704 0.019716
R58718 ASIG5V.n4723 ASIG5V.n3640 0.019716
R58719 ASIG5V.n4723 ASIG5V.n3705 0.019716
R58720 ASIG5V.n4727 ASIG5V.n3639 0.019716
R58721 ASIG5V.n4727 ASIG5V.n3706 0.019716
R58722 ASIG5V.n4732 ASIG5V.n3638 0.019716
R58723 ASIG5V.n4732 ASIG5V.n3707 0.019716
R58724 ASIG5V.n4736 ASIG5V.n3637 0.019716
R58725 ASIG5V.n4736 ASIG5V.n3708 0.019716
R58726 ASIG5V.n4741 ASIG5V.n3636 0.019716
R58727 ASIG5V.n4741 ASIG5V.n3709 0.019716
R58728 ASIG5V.n4745 ASIG5V.n3635 0.019716
R58729 ASIG5V.n4745 ASIG5V.n3710 0.019716
R58730 ASIG5V.n4750 ASIG5V.n3634 0.019716
R58731 ASIG5V.n4750 ASIG5V.n3711 0.019716
R58732 ASIG5V.n4754 ASIG5V.n3633 0.019716
R58733 ASIG5V.n4754 ASIG5V.n3712 0.019716
R58734 ASIG5V.n4759 ASIG5V.n3632 0.019716
R58735 ASIG5V.n4759 ASIG5V.n3713 0.019716
R58736 ASIG5V.n4763 ASIG5V.n3631 0.019716
R58737 ASIG5V.n4763 ASIG5V.n3714 0.019716
R58738 ASIG5V.n4768 ASIG5V.n3630 0.019716
R58739 ASIG5V.n4768 ASIG5V.n3715 0.019716
R58740 ASIG5V.n11162 ASIG5V.n10415 0.019716
R58741 ASIG5V.n10464 ASIG5V.n10414 0.019716
R58742 ASIG5V.n10464 ASIG5V.n10462 0.019716
R58743 ASIG5V.n11153 ASIG5V.n10413 0.019716
R58744 ASIG5V.n11153 ASIG5V.n10461 0.019716
R58745 ASIG5V.n10928 ASIG5V.n10412 0.019716
R58746 ASIG5V.n10928 ASIG5V.n10460 0.019716
R58747 ASIG5V.n11145 ASIG5V.n10411 0.019716
R58748 ASIG5V.n11145 ASIG5V.n10459 0.019716
R58749 ASIG5V.n10932 ASIG5V.n10410 0.019716
R58750 ASIG5V.n10932 ASIG5V.n10458 0.019716
R58751 ASIG5V.n11137 ASIG5V.n10409 0.019716
R58752 ASIG5V.n11137 ASIG5V.n10457 0.019716
R58753 ASIG5V.n10936 ASIG5V.n10408 0.019716
R58754 ASIG5V.n10936 ASIG5V.n10456 0.019716
R58755 ASIG5V.n11129 ASIG5V.n10407 0.019716
R58756 ASIG5V.n11129 ASIG5V.n10455 0.019716
R58757 ASIG5V.n10940 ASIG5V.n10406 0.019716
R58758 ASIG5V.n10940 ASIG5V.n10454 0.019716
R58759 ASIG5V.n11121 ASIG5V.n10405 0.019716
R58760 ASIG5V.n11121 ASIG5V.n10453 0.019716
R58761 ASIG5V.n10944 ASIG5V.n10404 0.019716
R58762 ASIG5V.n10944 ASIG5V.n10452 0.019716
R58763 ASIG5V.n11113 ASIG5V.n10403 0.019716
R58764 ASIG5V.n11113 ASIG5V.n10451 0.019716
R58765 ASIG5V.n10948 ASIG5V.n10402 0.019716
R58766 ASIG5V.n10948 ASIG5V.n10450 0.019716
R58767 ASIG5V.n11105 ASIG5V.n10401 0.019716
R58768 ASIG5V.n11105 ASIG5V.n10449 0.019716
R58769 ASIG5V.n10952 ASIG5V.n10400 0.019716
R58770 ASIG5V.n10952 ASIG5V.n10448 0.019716
R58771 ASIG5V.n11097 ASIG5V.n10399 0.019716
R58772 ASIG5V.n11097 ASIG5V.n10447 0.019716
R58773 ASIG5V.n10956 ASIG5V.n10398 0.019716
R58774 ASIG5V.n10956 ASIG5V.n10446 0.019716
R58775 ASIG5V.n11089 ASIG5V.n10397 0.019716
R58776 ASIG5V.n11089 ASIG5V.n10445 0.019716
R58777 ASIG5V.n10960 ASIG5V.n10396 0.019716
R58778 ASIG5V.n10960 ASIG5V.n10444 0.019716
R58779 ASIG5V.n11081 ASIG5V.n10395 0.019716
R58780 ASIG5V.n11081 ASIG5V.n10443 0.019716
R58781 ASIG5V.n10964 ASIG5V.n10394 0.019716
R58782 ASIG5V.n10964 ASIG5V.n10442 0.019716
R58783 ASIG5V.n11073 ASIG5V.n10393 0.019716
R58784 ASIG5V.n11073 ASIG5V.n10441 0.019716
R58785 ASIG5V.n10968 ASIG5V.n10392 0.019716
R58786 ASIG5V.n10968 ASIG5V.n10440 0.019716
R58787 ASIG5V.n11065 ASIG5V.n10391 0.019716
R58788 ASIG5V.n11065 ASIG5V.n10439 0.019716
R58789 ASIG5V.n10972 ASIG5V.n10390 0.019716
R58790 ASIG5V.n10972 ASIG5V.n10438 0.019716
R58791 ASIG5V.n11057 ASIG5V.n10389 0.019716
R58792 ASIG5V.n11057 ASIG5V.n10437 0.019716
R58793 ASIG5V.n10976 ASIG5V.n10388 0.019716
R58794 ASIG5V.n10976 ASIG5V.n10436 0.019716
R58795 ASIG5V.n11049 ASIG5V.n10387 0.019716
R58796 ASIG5V.n11049 ASIG5V.n10435 0.019716
R58797 ASIG5V.n10980 ASIG5V.n10386 0.019716
R58798 ASIG5V.n10980 ASIG5V.n10434 0.019716
R58799 ASIG5V.n11041 ASIG5V.n10385 0.019716
R58800 ASIG5V.n11041 ASIG5V.n10433 0.019716
R58801 ASIG5V.n10984 ASIG5V.n10384 0.019716
R58802 ASIG5V.n10984 ASIG5V.n10432 0.019716
R58803 ASIG5V.n11033 ASIG5V.n10383 0.019716
R58804 ASIG5V.n11033 ASIG5V.n10431 0.019716
R58805 ASIG5V.n10988 ASIG5V.n10382 0.019716
R58806 ASIG5V.n10988 ASIG5V.n10430 0.019716
R58807 ASIG5V.n11025 ASIG5V.n10381 0.019716
R58808 ASIG5V.n11025 ASIG5V.n10429 0.019716
R58809 ASIG5V.n10992 ASIG5V.n10380 0.019716
R58810 ASIG5V.n10992 ASIG5V.n10428 0.019716
R58811 ASIG5V.n11017 ASIG5V.n10379 0.019716
R58812 ASIG5V.n11017 ASIG5V.n10427 0.019716
R58813 ASIG5V.n10996 ASIG5V.n10378 0.019716
R58814 ASIG5V.n10996 ASIG5V.n10426 0.019716
R58815 ASIG5V.n11009 ASIG5V.n10377 0.019716
R58816 ASIG5V.n11009 ASIG5V.n10425 0.019716
R58817 ASIG5V.n11000 ASIG5V.n10376 0.019716
R58818 ASIG5V.n11000 ASIG5V.n10424 0.019716
R58819 ASIG5V.n10422 ASIG5V.n10375 0.019716
R58820 ASIG5V.n11164 ASIG5V.n10422 0.019716
R58821 ASIG5V.n10418 ASIG5V.n10374 0.019716
R58822 ASIG5V.n10418 ASIG5V.n10417 0.019716
R58823 ASIG5V.n11161 ASIG5V.n10414 0.019716
R58824 ASIG5V.n11162 ASIG5V.n11161 0.019716
R58825 ASIG5V.n11155 ASIG5V.n10413 0.019716
R58826 ASIG5V.n11155 ASIG5V.n10462 0.019716
R58827 ASIG5V.n10930 ASIG5V.n10412 0.019716
R58828 ASIG5V.n10930 ASIG5V.n10461 0.019716
R58829 ASIG5V.n11147 ASIG5V.n10411 0.019716
R58830 ASIG5V.n11147 ASIG5V.n10460 0.019716
R58831 ASIG5V.n10934 ASIG5V.n10410 0.019716
R58832 ASIG5V.n10934 ASIG5V.n10459 0.019716
R58833 ASIG5V.n11139 ASIG5V.n10409 0.019716
R58834 ASIG5V.n11139 ASIG5V.n10458 0.019716
R58835 ASIG5V.n10938 ASIG5V.n10408 0.019716
R58836 ASIG5V.n10938 ASIG5V.n10457 0.019716
R58837 ASIG5V.n11131 ASIG5V.n10407 0.019716
R58838 ASIG5V.n11131 ASIG5V.n10456 0.019716
R58839 ASIG5V.n10942 ASIG5V.n10406 0.019716
R58840 ASIG5V.n10942 ASIG5V.n10455 0.019716
R58841 ASIG5V.n11123 ASIG5V.n10405 0.019716
R58842 ASIG5V.n11123 ASIG5V.n10454 0.019716
R58843 ASIG5V.n10946 ASIG5V.n10404 0.019716
R58844 ASIG5V.n10946 ASIG5V.n10453 0.019716
R58845 ASIG5V.n11115 ASIG5V.n10403 0.019716
R58846 ASIG5V.n11115 ASIG5V.n10452 0.019716
R58847 ASIG5V.n10950 ASIG5V.n10402 0.019716
R58848 ASIG5V.n10950 ASIG5V.n10451 0.019716
R58849 ASIG5V.n11107 ASIG5V.n10401 0.019716
R58850 ASIG5V.n11107 ASIG5V.n10450 0.019716
R58851 ASIG5V.n10954 ASIG5V.n10400 0.019716
R58852 ASIG5V.n10954 ASIG5V.n10449 0.019716
R58853 ASIG5V.n11099 ASIG5V.n10399 0.019716
R58854 ASIG5V.n11099 ASIG5V.n10448 0.019716
R58855 ASIG5V.n10958 ASIG5V.n10398 0.019716
R58856 ASIG5V.n10958 ASIG5V.n10447 0.019716
R58857 ASIG5V.n11091 ASIG5V.n10397 0.019716
R58858 ASIG5V.n11091 ASIG5V.n10446 0.019716
R58859 ASIG5V.n10962 ASIG5V.n10396 0.019716
R58860 ASIG5V.n10962 ASIG5V.n10445 0.019716
R58861 ASIG5V.n11083 ASIG5V.n10395 0.019716
R58862 ASIG5V.n11083 ASIG5V.n10444 0.019716
R58863 ASIG5V.n10966 ASIG5V.n10394 0.019716
R58864 ASIG5V.n10966 ASIG5V.n10443 0.019716
R58865 ASIG5V.n11075 ASIG5V.n10393 0.019716
R58866 ASIG5V.n11075 ASIG5V.n10442 0.019716
R58867 ASIG5V.n10970 ASIG5V.n10392 0.019716
R58868 ASIG5V.n10970 ASIG5V.n10441 0.019716
R58869 ASIG5V.n11067 ASIG5V.n10391 0.019716
R58870 ASIG5V.n11067 ASIG5V.n10440 0.019716
R58871 ASIG5V.n10974 ASIG5V.n10390 0.019716
R58872 ASIG5V.n10974 ASIG5V.n10439 0.019716
R58873 ASIG5V.n11059 ASIG5V.n10389 0.019716
R58874 ASIG5V.n11059 ASIG5V.n10438 0.019716
R58875 ASIG5V.n10978 ASIG5V.n10388 0.019716
R58876 ASIG5V.n10978 ASIG5V.n10437 0.019716
R58877 ASIG5V.n11051 ASIG5V.n10387 0.019716
R58878 ASIG5V.n11051 ASIG5V.n10436 0.019716
R58879 ASIG5V.n10982 ASIG5V.n10386 0.019716
R58880 ASIG5V.n10982 ASIG5V.n10435 0.019716
R58881 ASIG5V.n11043 ASIG5V.n10385 0.019716
R58882 ASIG5V.n11043 ASIG5V.n10434 0.019716
R58883 ASIG5V.n10986 ASIG5V.n10384 0.019716
R58884 ASIG5V.n10986 ASIG5V.n10433 0.019716
R58885 ASIG5V.n11035 ASIG5V.n10383 0.019716
R58886 ASIG5V.n11035 ASIG5V.n10432 0.019716
R58887 ASIG5V.n10990 ASIG5V.n10382 0.019716
R58888 ASIG5V.n10990 ASIG5V.n10431 0.019716
R58889 ASIG5V.n11027 ASIG5V.n10381 0.019716
R58890 ASIG5V.n11027 ASIG5V.n10430 0.019716
R58891 ASIG5V.n10994 ASIG5V.n10380 0.019716
R58892 ASIG5V.n10994 ASIG5V.n10429 0.019716
R58893 ASIG5V.n11019 ASIG5V.n10379 0.019716
R58894 ASIG5V.n11019 ASIG5V.n10428 0.019716
R58895 ASIG5V.n10998 ASIG5V.n10378 0.019716
R58896 ASIG5V.n10998 ASIG5V.n10427 0.019716
R58897 ASIG5V.n11011 ASIG5V.n10377 0.019716
R58898 ASIG5V.n11011 ASIG5V.n10426 0.019716
R58899 ASIG5V.n11002 ASIG5V.n10376 0.019716
R58900 ASIG5V.n11002 ASIG5V.n10425 0.019716
R58901 ASIG5V.n11003 ASIG5V.n10375 0.019716
R58902 ASIG5V.n11003 ASIG5V.n10424 0.019716
R58903 ASIG5V.n11165 ASIG5V.n10374 0.019716
R58904 ASIG5V.n11165 ASIG5V.n11164 0.019716
R58905 ASIG5V.n11171 ASIG5V.n10417 0.019716
R58906 ASIG5V.n4553 ASIG5V.n3829 0.019716
R58907 ASIG5V.n4310 ASIG5V.n3828 0.019716
R58908 ASIG5V.n4310 ASIG5V.n4308 0.019716
R58909 ASIG5V.n4544 ASIG5V.n3827 0.019716
R58910 ASIG5V.n4544 ASIG5V.n4307 0.019716
R58911 ASIG5V.n4313 ASIG5V.n3826 0.019716
R58912 ASIG5V.n4313 ASIG5V.n4306 0.019716
R58913 ASIG5V.n4536 ASIG5V.n3825 0.019716
R58914 ASIG5V.n4536 ASIG5V.n4305 0.019716
R58915 ASIG5V.n4317 ASIG5V.n3824 0.019716
R58916 ASIG5V.n4317 ASIG5V.n4304 0.019716
R58917 ASIG5V.n4528 ASIG5V.n3823 0.019716
R58918 ASIG5V.n4528 ASIG5V.n4303 0.019716
R58919 ASIG5V.n4321 ASIG5V.n3822 0.019716
R58920 ASIG5V.n4321 ASIG5V.n4302 0.019716
R58921 ASIG5V.n4520 ASIG5V.n3821 0.019716
R58922 ASIG5V.n4520 ASIG5V.n4301 0.019716
R58923 ASIG5V.n4325 ASIG5V.n3820 0.019716
R58924 ASIG5V.n4325 ASIG5V.n4300 0.019716
R58925 ASIG5V.n4512 ASIG5V.n3819 0.019716
R58926 ASIG5V.n4512 ASIG5V.n4299 0.019716
R58927 ASIG5V.n4329 ASIG5V.n3818 0.019716
R58928 ASIG5V.n4329 ASIG5V.n4298 0.019716
R58929 ASIG5V.n4504 ASIG5V.n3817 0.019716
R58930 ASIG5V.n4504 ASIG5V.n4297 0.019716
R58931 ASIG5V.n4333 ASIG5V.n3816 0.019716
R58932 ASIG5V.n4333 ASIG5V.n4296 0.019716
R58933 ASIG5V.n4496 ASIG5V.n3815 0.019716
R58934 ASIG5V.n4496 ASIG5V.n4295 0.019716
R58935 ASIG5V.n4337 ASIG5V.n3814 0.019716
R58936 ASIG5V.n4337 ASIG5V.n4294 0.019716
R58937 ASIG5V.n4488 ASIG5V.n3813 0.019716
R58938 ASIG5V.n4488 ASIG5V.n4293 0.019716
R58939 ASIG5V.n4341 ASIG5V.n3812 0.019716
R58940 ASIG5V.n4341 ASIG5V.n4292 0.019716
R58941 ASIG5V.n4480 ASIG5V.n3811 0.019716
R58942 ASIG5V.n4480 ASIG5V.n4291 0.019716
R58943 ASIG5V.n4345 ASIG5V.n3810 0.019716
R58944 ASIG5V.n4345 ASIG5V.n4290 0.019716
R58945 ASIG5V.n4472 ASIG5V.n3809 0.019716
R58946 ASIG5V.n4472 ASIG5V.n4289 0.019716
R58947 ASIG5V.n4349 ASIG5V.n3808 0.019716
R58948 ASIG5V.n4349 ASIG5V.n4288 0.019716
R58949 ASIG5V.n4464 ASIG5V.n3807 0.019716
R58950 ASIG5V.n4464 ASIG5V.n4287 0.019716
R58951 ASIG5V.n4353 ASIG5V.n3806 0.019716
R58952 ASIG5V.n4353 ASIG5V.n4286 0.019716
R58953 ASIG5V.n4456 ASIG5V.n3805 0.019716
R58954 ASIG5V.n4456 ASIG5V.n4285 0.019716
R58955 ASIG5V.n4357 ASIG5V.n3804 0.019716
R58956 ASIG5V.n4357 ASIG5V.n4284 0.019716
R58957 ASIG5V.n4448 ASIG5V.n3803 0.019716
R58958 ASIG5V.n4448 ASIG5V.n4283 0.019716
R58959 ASIG5V.n4361 ASIG5V.n3802 0.019716
R58960 ASIG5V.n4361 ASIG5V.n4282 0.019716
R58961 ASIG5V.n4440 ASIG5V.n3801 0.019716
R58962 ASIG5V.n4440 ASIG5V.n4281 0.019716
R58963 ASIG5V.n4365 ASIG5V.n3800 0.019716
R58964 ASIG5V.n4365 ASIG5V.n4280 0.019716
R58965 ASIG5V.n4432 ASIG5V.n3799 0.019716
R58966 ASIG5V.n4432 ASIG5V.n4279 0.019716
R58967 ASIG5V.n4369 ASIG5V.n3798 0.019716
R58968 ASIG5V.n4369 ASIG5V.n4278 0.019716
R58969 ASIG5V.n4424 ASIG5V.n3797 0.019716
R58970 ASIG5V.n4424 ASIG5V.n4277 0.019716
R58971 ASIG5V.n4373 ASIG5V.n3796 0.019716
R58972 ASIG5V.n4373 ASIG5V.n4276 0.019716
R58973 ASIG5V.n4416 ASIG5V.n3795 0.019716
R58974 ASIG5V.n4416 ASIG5V.n4275 0.019716
R58975 ASIG5V.n4377 ASIG5V.n3794 0.019716
R58976 ASIG5V.n4377 ASIG5V.n4274 0.019716
R58977 ASIG5V.n4408 ASIG5V.n3793 0.019716
R58978 ASIG5V.n4408 ASIG5V.n4273 0.019716
R58979 ASIG5V.n4381 ASIG5V.n3792 0.019716
R58980 ASIG5V.n4381 ASIG5V.n4272 0.019716
R58981 ASIG5V.n4400 ASIG5V.n3791 0.019716
R58982 ASIG5V.n4400 ASIG5V.n4271 0.019716
R58983 ASIG5V.n4385 ASIG5V.n3790 0.019716
R58984 ASIG5V.n4385 ASIG5V.n4270 0.019716
R58985 ASIG5V.n4392 ASIG5V.n3789 0.019716
R58986 ASIG5V.n4392 ASIG5V.n4269 0.019716
R58987 ASIG5V.n3833 ASIG5V.n3788 0.019716
R58988 ASIG5V.n3833 ASIG5V.n3832 0.019716
R58989 ASIG5V.n4552 ASIG5V.n3828 0.019716
R58990 ASIG5V.n4553 ASIG5V.n4552 0.019716
R58991 ASIG5V.n4546 ASIG5V.n3827 0.019716
R58992 ASIG5V.n4546 ASIG5V.n4308 0.019716
R58993 ASIG5V.n4315 ASIG5V.n3826 0.019716
R58994 ASIG5V.n4315 ASIG5V.n4307 0.019716
R58995 ASIG5V.n4538 ASIG5V.n3825 0.019716
R58996 ASIG5V.n4538 ASIG5V.n4306 0.019716
R58997 ASIG5V.n4319 ASIG5V.n3824 0.019716
R58998 ASIG5V.n4319 ASIG5V.n4305 0.019716
R58999 ASIG5V.n4530 ASIG5V.n3823 0.019716
R59000 ASIG5V.n4530 ASIG5V.n4304 0.019716
R59001 ASIG5V.n4323 ASIG5V.n3822 0.019716
R59002 ASIG5V.n4323 ASIG5V.n4303 0.019716
R59003 ASIG5V.n4522 ASIG5V.n3821 0.019716
R59004 ASIG5V.n4522 ASIG5V.n4302 0.019716
R59005 ASIG5V.n4327 ASIG5V.n3820 0.019716
R59006 ASIG5V.n4327 ASIG5V.n4301 0.019716
R59007 ASIG5V.n4514 ASIG5V.n3819 0.019716
R59008 ASIG5V.n4514 ASIG5V.n4300 0.019716
R59009 ASIG5V.n4331 ASIG5V.n3818 0.019716
R59010 ASIG5V.n4331 ASIG5V.n4299 0.019716
R59011 ASIG5V.n4506 ASIG5V.n3817 0.019716
R59012 ASIG5V.n4506 ASIG5V.n4298 0.019716
R59013 ASIG5V.n4335 ASIG5V.n3816 0.019716
R59014 ASIG5V.n4335 ASIG5V.n4297 0.019716
R59015 ASIG5V.n4498 ASIG5V.n3815 0.019716
R59016 ASIG5V.n4498 ASIG5V.n4296 0.019716
R59017 ASIG5V.n4339 ASIG5V.n3814 0.019716
R59018 ASIG5V.n4339 ASIG5V.n4295 0.019716
R59019 ASIG5V.n4490 ASIG5V.n3813 0.019716
R59020 ASIG5V.n4490 ASIG5V.n4294 0.019716
R59021 ASIG5V.n4343 ASIG5V.n3812 0.019716
R59022 ASIG5V.n4343 ASIG5V.n4293 0.019716
R59023 ASIG5V.n4482 ASIG5V.n3811 0.019716
R59024 ASIG5V.n4482 ASIG5V.n4292 0.019716
R59025 ASIG5V.n4347 ASIG5V.n3810 0.019716
R59026 ASIG5V.n4347 ASIG5V.n4291 0.019716
R59027 ASIG5V.n4474 ASIG5V.n3809 0.019716
R59028 ASIG5V.n4474 ASIG5V.n4290 0.019716
R59029 ASIG5V.n4351 ASIG5V.n3808 0.019716
R59030 ASIG5V.n4351 ASIG5V.n4289 0.019716
R59031 ASIG5V.n4466 ASIG5V.n3807 0.019716
R59032 ASIG5V.n4466 ASIG5V.n4288 0.019716
R59033 ASIG5V.n4355 ASIG5V.n3806 0.019716
R59034 ASIG5V.n4355 ASIG5V.n4287 0.019716
R59035 ASIG5V.n4458 ASIG5V.n3805 0.019716
R59036 ASIG5V.n4458 ASIG5V.n4286 0.019716
R59037 ASIG5V.n4359 ASIG5V.n3804 0.019716
R59038 ASIG5V.n4359 ASIG5V.n4285 0.019716
R59039 ASIG5V.n4450 ASIG5V.n3803 0.019716
R59040 ASIG5V.n4450 ASIG5V.n4284 0.019716
R59041 ASIG5V.n4363 ASIG5V.n3802 0.019716
R59042 ASIG5V.n4363 ASIG5V.n4283 0.019716
R59043 ASIG5V.n4442 ASIG5V.n3801 0.019716
R59044 ASIG5V.n4442 ASIG5V.n4282 0.019716
R59045 ASIG5V.n4367 ASIG5V.n3800 0.019716
R59046 ASIG5V.n4367 ASIG5V.n4281 0.019716
R59047 ASIG5V.n4434 ASIG5V.n3799 0.019716
R59048 ASIG5V.n4434 ASIG5V.n4280 0.019716
R59049 ASIG5V.n4371 ASIG5V.n3798 0.019716
R59050 ASIG5V.n4371 ASIG5V.n4279 0.019716
R59051 ASIG5V.n4426 ASIG5V.n3797 0.019716
R59052 ASIG5V.n4426 ASIG5V.n4278 0.019716
R59053 ASIG5V.n4375 ASIG5V.n3796 0.019716
R59054 ASIG5V.n4375 ASIG5V.n4277 0.019716
R59055 ASIG5V.n4418 ASIG5V.n3795 0.019716
R59056 ASIG5V.n4418 ASIG5V.n4276 0.019716
R59057 ASIG5V.n4379 ASIG5V.n3794 0.019716
R59058 ASIG5V.n4379 ASIG5V.n4275 0.019716
R59059 ASIG5V.n4410 ASIG5V.n3793 0.019716
R59060 ASIG5V.n4410 ASIG5V.n4274 0.019716
R59061 ASIG5V.n4383 ASIG5V.n3792 0.019716
R59062 ASIG5V.n4383 ASIG5V.n4273 0.019716
R59063 ASIG5V.n4402 ASIG5V.n3791 0.019716
R59064 ASIG5V.n4402 ASIG5V.n4272 0.019716
R59065 ASIG5V.n4387 ASIG5V.n3790 0.019716
R59066 ASIG5V.n4387 ASIG5V.n4271 0.019716
R59067 ASIG5V.n4394 ASIG5V.n3789 0.019716
R59068 ASIG5V.n4394 ASIG5V.n4270 0.019716
R59069 ASIG5V.n4389 ASIG5V.n3788 0.019716
R59070 ASIG5V.n4389 ASIG5V.n4269 0.019716
R59071 ASIG5V.n4567 ASIG5V.n3832 0.019716
R59072 ASIG5V.n12532 ASIG5V.n7 0.019625
R59073 ASIG5V.n11178 ASIG5V.n10368 0.019625
R59074 ASIG5V.n1664 ASIG5V.n1416 0.0195611
R59075 ASIG5V.n1863 ASIG5V.n1850 0.0195611
R59076 ASIG5V.n12005 ASIG5V.n1665 0.0195611
R59077 ASIG5V.n1857 ASIG5V.n1852 0.0195611
R59078 ASIG5V.n12316 ASIG5V.n12315 0.019175
R59079 ASIG5V.n11491 ASIG5V.n11490 0.019175
R59080 ASIG5V.n6884 ASIG5V.n6633 0.0191681
R59081 ASIG5V.n8913 ASIG5V.n8912 0.0191681
R59082 ASIG5V.n8115 ASIG5V.n7467 0.0191
R59083 ASIG5V.n8128 ASIG5V.n7313 0.0191
R59084 ASIG5V.n8141 ASIG5V.n7292 0.0191
R59085 ASIG5V.n8154 ASIG5V.n7272 0.0191
R59086 ASIG5V.n7540 ASIG5V.n7528 0.0191
R59087 ASIG5V.n9753 ASIG5V.n3159 0.0191
R59088 ASIG5V.n4561 ASIG5V.n3831 0.0187751
R59089 ASIG5V.n4562 ASIG5V.n3835 0.0187751
R59090 ASIG5V.n9425 ASIG5V.n9424 0.018725
R59091 ASIG5V.n9742 ASIG5V.n3172 0.0175961
R59092 ASIG5V.n9741 ASIG5V.n3174 0.0175961
R59093 ASIG5V.n4265 ASIG5V.n3784 0.017282
R59094 ASIG5V.n4572 ASIG5V.n3784 0.017282
R59095 ASIG5V.n4575 ASIG5V.n4574 0.017282
R59096 ASIG5V.n4574 ASIG5V.n3777 0.017282
R59097 ASIG5V.n4583 ASIG5V.n3617 0.017282
R59098 ASIG5V.n4791 ASIG5V.n3617 0.017282
R59099 ASIG5V.n4795 ASIG5V.n4794 0.017282
R59100 ASIG5V.n4794 ASIG5V.n4793 0.017282
R59101 ASIG5V.n4812 ASIG5V.n3163 0.017282
R59102 ASIG5V.n9747 ASIG5V.n3164 0.017282
R59103 ASIG5V.n9438 ASIG5V.n3164 0.017282
R59104 ASIG5V.n9438 ASIG5V.n9437 0.017282
R59105 ASIG5V.n9437 ASIG5V.n9436 0.017282
R59106 ASIG5V.n7964 ASIG5V.n7961 0.017282
R59107 ASIG5V.n7970 ASIG5V.n7961 0.017282
R59108 ASIG5V.n7972 ASIG5V.n7714 0.017282
R59109 ASIG5V.n9402 ASIG5V.n9401 0.017282
R59110 ASIG5V.n9401 ASIG5V.n9400 0.017282
R59111 ASIG5V.n6422 ASIG5V.n6420 0.017282
R59112 ASIG5V.n6422 ASIG5V.n6421 0.017282
R59113 ASIG5V.n6421 ASIG5V.n6415 0.017282
R59114 ASIG5V.n6535 ASIG5V.n6534 0.017282
R59115 ASIG5V.n8925 ASIG5V.n8924 0.017282
R59116 ASIG5V.n8924 ASIG5V.n8923 0.017282
R59117 ASIG5V.n7234 ASIG5V.n7232 0.017282
R59118 ASIG5V.n7243 ASIG5V.n7232 0.017282
R59119 ASIG5V.n8900 ASIG5V.n8899 0.017282
R59120 ASIG5V.n8899 ASIG5V.n8168 0.017282
R59121 ASIG5V.n8570 ASIG5V.n8322 0.017282
R59122 ASIG5V.n8576 ASIG5V.n8322 0.017282
R59123 ASIG5V.n8586 ASIG5V.n8577 0.017282
R59124 ASIG5V.n8577 ASIG5V.n161 0.017282
R59125 ASIG5V.n12336 ASIG5V.n162 0.017282
R59126 ASIG5V.n12330 ASIG5V.n162 0.017282
R59127 ASIG5V.n12327 ASIG5V.n170 0.017282
R59128 ASIG5V.n12307 ASIG5V.n170 0.017282
R59129 ASIG5V.n12305 ASIG5V.n525 0.017282
R59130 ASIG5V.n12285 ASIG5V.n525 0.017282
R59131 ASIG5V.n12285 ASIG5V.n12284 0.017282
R59132 ASIG5V.n12282 ASIG5V.n870 0.017282
R59133 ASIG5V.n12017 ASIG5V.n12016 0.017282
R59134 ASIG5V.n12016 ASIG5V.n12015 0.017282
R59135 ASIG5V.n1830 ASIG5V.n1829 0.017282
R59136 ASIG5V.n1829 ASIG5V.n1826 0.017282
R59137 ASIG5V.n11805 ASIG5V.n1827 0.017282
R59138 ASIG5V.n11799 ASIG5V.n1827 0.017282
R59139 ASIG5V.n11795 ASIG5V.n1843 0.017282
R59140 ASIG5V.n2560 ASIG5V.n1843 0.017282
R59141 ASIG5V.n11778 ASIG5V.n2562 0.017282
R59142 ASIG5V.n11778 ASIG5V.n11777 0.017282
R59143 ASIG5V.n11775 ASIG5V.n2564 0.017282
R59144 ASIG5V.n11500 ASIG5V.n11499 0.017282
R59145 ASIG5V.n11499 ASIG5V.n11498 0.017282
R59146 ASIG5V.n11189 ASIG5V.n10021 0.017282
R59147 ASIG5V.n11189 ASIG5V.n11188 0.017282
R59148 ASIG5V.n11188 ASIG5V.n11187 0.017282
R59149 ASIG5V.n10476 ASIG5V.n10475 0.017282
R59150 ASIG5V.n10476 ASIG5V.n10466 0.017282
R59151 ASIG5V.n10924 ASIG5V.n10467 0.017282
R59152 ASIG5V.n10708 ASIG5V.n10467 0.017282
R59153 ASIG5V.n12530 ASIG5V.n9 0.0172031
R59154 ASIG5V.n10366 ASIG5V.n10069 0.0172031
R59155 ASIG5V.n12531 ASIG5V.n8 0.0172031
R59156 ASIG5V.n11180 ASIG5V.n11179 0.0172031
R59157 ASIG5V.n9182 ASIG5V.n9181 0.016925
R59158 ASIG5V.n12313 ASIG5V.n217 0.01681
R59159 ASIG5V.n11493 ASIG5V.n9967 0.01681
R59160 ASIG5V.n12314 ASIG5V.n517 0.01681
R59161 ASIG5V.n11492 ASIG5V.n9968 0.01681
R59162 ASIG5V.n7982 ASIG5V.n7981 0.0167406
R59163 ASIG5V.n8570 ASIG5V.n8569 0.0167406
R59164 ASIG5V.n11498 ASIG5V.n9961 0.0167406
R59165 ASIG5V.n12001 ASIG5V.n1670 0.016475
R59166 ASIG5V.n1858 ASIG5V.n1670 0.016475
R59167 ASIG5V.n10709 ASIG5V.n10708 0.0164699
R59168 ASIG5V.n9422 ASIG5V.n5167 0.016417
R59169 ASIG5V.n9423 ASIG5V.n5461 0.016417
R59170 ASIG5V.n12307 ASIG5V.n12306 0.0161992
R59171 ASIG5V.n7340 ASIG5V.n870 0.0161992
R59172 ASIG5V.n11796 ASIG5V.n11795 0.0161992
R59173 ASIG5V.n9181 ASIG5V.n9180 0.016025
R59174 ASIG5V.n4575 ASIG5V.n4573 0.0156579
R59175 ASIG5V.n9400 ASIG5V.n5909 0.0156579
R59176 ASIG5V.n11798 ASIG5V.n11797 0.0156579
R59177 ASIG5V.n4267 ASIG5V.n3786 0.0154799
R59178 ASIG5V.n4570 ASIG5V.n3786 0.0154799
R59179 ASIG5V.n4578 ASIG5V.n4577 0.0154799
R59180 ASIG5V.n4579 ASIG5V.n4578 0.0154799
R59181 ASIG5V.n4788 ASIG5V.n3619 0.0154799
R59182 ASIG5V.n4789 ASIG5V.n4788 0.0154799
R59183 ASIG5V.n4797 ASIG5V.n3269 0.0154799
R59184 ASIG5V.n4809 ASIG5V.n3269 0.0154799
R59185 ASIG5V.n4811 ASIG5V.n3167 0.0154799
R59186 ASIG5V.n9745 ASIG5V.n3167 0.0154799
R59187 ASIG5V.n9745 ASIG5V.n3168 0.0154799
R59188 ASIG5V.n9440 ASIG5V.n3168 0.0154799
R59189 ASIG5V.n9440 ASIG5V.n5118 0.0154799
R59190 ASIG5V.n9434 ASIG5V.n5118 0.0154799
R59191 ASIG5V.n7967 ASIG5V.n7966 0.0154799
R59192 ASIG5V.n7968 ASIG5V.n7967 0.0154799
R59193 ASIG5V.n7975 ASIG5V.n7974 0.0154799
R59194 ASIG5V.n7979 ASIG5V.n7975 0.0154799
R59195 ASIG5V.n9404 ASIG5V.n5570 0.0154799
R59196 ASIG5V.n9398 ASIG5V.n5570 0.0154799
R59197 ASIG5V.n6424 ASIG5V.n6418 0.0154799
R59198 ASIG5V.n6425 ASIG5V.n6424 0.0154799
R59199 ASIG5V.n6426 ASIG5V.n6425 0.0154799
R59200 ASIG5V.n9188 ASIG5V.n9187 0.0154799
R59201 ASIG5V.n9187 ASIG5V.n6430 0.0154799
R59202 ASIG5V.n6542 ASIG5V.n6539 0.0154799
R59203 ASIG5V.n8921 ASIG5V.n6542 0.0154799
R59204 ASIG5V.n7237 ASIG5V.n7236 0.0154799
R59205 ASIG5V.n7241 ASIG5V.n7237 0.0154799
R59206 ASIG5V.n8904 ASIG5V.n6894 0.0154799
R59207 ASIG5V.n8897 ASIG5V.n6894 0.0154799
R59208 ASIG5V.n8897 ASIG5V.n8170 0.0154799
R59209 ASIG5V.n8573 ASIG5V.n8572 0.0154799
R59210 ASIG5V.n8574 ASIG5V.n8573 0.0154799
R59211 ASIG5V.n8584 ASIG5V.n8581 0.0154799
R59212 ASIG5V.n8581 ASIG5V.n8580 0.0154799
R59213 ASIG5V.n12334 ASIG5V.n12333 0.0154799
R59214 ASIG5V.n12333 ASIG5V.n12332 0.0154799
R59215 ASIG5V.n12325 ASIG5V.n172 0.0154799
R59216 ASIG5V.n12309 ASIG5V.n172 0.0154799
R59217 ASIG5V.n12303 ASIG5V.n527 0.0154799
R59218 ASIG5V.n12287 ASIG5V.n527 0.0154799
R59219 ASIG5V.n12287 ASIG5V.n867 0.0154799
R59220 ASIG5V.n12280 ASIG5V.n874 0.0154799
R59221 ASIG5V.n1319 ASIG5V.n874 0.0154799
R59222 ASIG5V.n1324 ASIG5V.n1321 0.0154799
R59223 ASIG5V.n12013 ASIG5V.n1324 0.0154799
R59224 ASIG5V.n1833 ASIG5V.n1832 0.0154799
R59225 ASIG5V.n1834 ASIG5V.n1833 0.0154799
R59226 ASIG5V.n11803 ASIG5V.n11802 0.0154799
R59227 ASIG5V.n11802 ASIG5V.n11801 0.0154799
R59228 ASIG5V.n11801 ASIG5V.n1838 0.0154799
R59229 ASIG5V.n11793 ASIG5V.n1847 0.0154799
R59230 ASIG5V.n2558 ASIG5V.n1847 0.0154799
R59231 ASIG5V.n11780 ASIG5V.n2214 0.0154799
R59232 ASIG5V.n11780 ASIG5V.n2215 0.0154799
R59233 ASIG5V.n11773 ASIG5V.n2568 0.0154799
R59234 ASIG5V.n9958 ASIG5V.n2568 0.0154799
R59235 ASIG5V.n9963 ASIG5V.n9960 0.0154799
R59236 ASIG5V.n11496 ASIG5V.n9963 0.0154799
R59237 ASIG5V.n11191 ASIG5V.n10017 0.0154799
R59238 ASIG5V.n11191 ASIG5V.n10018 0.0154799
R59239 ASIG5V.n11185 ASIG5V.n10018 0.0154799
R59240 ASIG5V.n10473 ASIG5V.n10470 0.0154799
R59241 ASIG5V.n10479 ASIG5V.n10470 0.0154799
R59242 ASIG5V.n10922 ASIG5V.n10921 0.0154799
R59243 ASIG5V.n10921 ASIG5V.n10481 0.0154799
R59244 ASIG5V.n4266 ASIG5V.n3785 0.0154799
R59245 ASIG5V.n4571 ASIG5V.n3785 0.0154799
R59246 ASIG5V.n4576 ASIG5V.n3778 0.0154799
R59247 ASIG5V.n4580 ASIG5V.n3778 0.0154799
R59248 ASIG5V.n4582 ASIG5V.n3618 0.0154799
R59249 ASIG5V.n4790 ASIG5V.n3618 0.0154799
R59250 ASIG5V.n4796 ASIG5V.n3281 0.0154799
R59251 ASIG5V.n3281 ASIG5V.n3268 0.0154799
R59252 ASIG5V.n4813 ASIG5V.n3165 0.0154799
R59253 ASIG5V.n9746 ASIG5V.n3165 0.0154799
R59254 ASIG5V.n9746 ASIG5V.n3166 0.0154799
R59255 ASIG5V.n9439 ASIG5V.n3166 0.0154799
R59256 ASIG5V.n9439 ASIG5V.n5119 0.0154799
R59257 ASIG5V.n9435 ASIG5V.n5119 0.0154799
R59258 ASIG5V.n7965 ASIG5V.n7962 0.0154799
R59259 ASIG5V.n7969 ASIG5V.n7962 0.0154799
R59260 ASIG5V.n7973 ASIG5V.n7715 0.0154799
R59261 ASIG5V.n7980 ASIG5V.n7715 0.0154799
R59262 ASIG5V.n9403 ASIG5V.n5572 0.0154799
R59263 ASIG5V.n9399 ASIG5V.n5572 0.0154799
R59264 ASIG5V.n6423 ASIG5V.n6419 0.0154799
R59265 ASIG5V.n6423 ASIG5V.n6417 0.0154799
R59266 ASIG5V.n6427 ASIG5V.n6417 0.0154799
R59267 ASIG5V.n9189 ASIG5V.n6429 0.0154799
R59268 ASIG5V.n6536 ASIG5V.n6429 0.0154799
R59269 ASIG5V.n8926 ASIG5V.n6537 0.0154799
R59270 ASIG5V.n8922 ASIG5V.n6537 0.0154799
R59271 ASIG5V.n7235 ASIG5V.n7233 0.0154799
R59272 ASIG5V.n7242 ASIG5V.n7233 0.0154799
R59273 ASIG5V.n8903 ASIG5V.n6896 0.0154799
R59274 ASIG5V.n8898 ASIG5V.n6896 0.0154799
R59275 ASIG5V.n8898 ASIG5V.n8169 0.0154799
R59276 ASIG5V.n8571 ASIG5V.n8323 0.0154799
R59277 ASIG5V.n8575 ASIG5V.n8323 0.0154799
R59278 ASIG5V.n8585 ASIG5V.n8578 0.0154799
R59279 ASIG5V.n8579 ASIG5V.n8578 0.0154799
R59280 ASIG5V.n12335 ASIG5V.n164 0.0154799
R59281 ASIG5V.n12331 ASIG5V.n164 0.0154799
R59282 ASIG5V.n12326 ASIG5V.n171 0.0154799
R59283 ASIG5V.n12308 ASIG5V.n171 0.0154799
R59284 ASIG5V.n12304 ASIG5V.n526 0.0154799
R59285 ASIG5V.n12286 ASIG5V.n526 0.0154799
R59286 ASIG5V.n12286 ASIG5V.n868 0.0154799
R59287 ASIG5V.n12281 ASIG5V.n872 0.0154799
R59288 ASIG5V.n1317 ASIG5V.n872 0.0154799
R59289 ASIG5V.n12018 ASIG5V.n1318 0.0154799
R59290 ASIG5V.n12014 ASIG5V.n1318 0.0154799
R59291 ASIG5V.n1831 ASIG5V.n1828 0.0154799
R59292 ASIG5V.n1835 ASIG5V.n1828 0.0154799
R59293 ASIG5V.n11804 ASIG5V.n1837 0.0154799
R59294 ASIG5V.n11800 ASIG5V.n1837 0.0154799
R59295 ASIG5V.n11800 ASIG5V.n1840 0.0154799
R59296 ASIG5V.n11794 ASIG5V.n1845 0.0154799
R59297 ASIG5V.n2559 ASIG5V.n1845 0.0154799
R59298 ASIG5V.n11779 ASIG5V.n2216 0.0154799
R59299 ASIG5V.n11779 ASIG5V.n2217 0.0154799
R59300 ASIG5V.n11774 ASIG5V.n2566 0.0154799
R59301 ASIG5V.n9955 ASIG5V.n2566 0.0154799
R59302 ASIG5V.n11501 ASIG5V.n9956 0.0154799
R59303 ASIG5V.n11497 ASIG5V.n9956 0.0154799
R59304 ASIG5V.n11190 ASIG5V.n10019 0.0154799
R59305 ASIG5V.n11190 ASIG5V.n10020 0.0154799
R59306 ASIG5V.n11186 ASIG5V.n10020 0.0154799
R59307 ASIG5V.n10477 ASIG5V.n10474 0.0154799
R59308 ASIG5V.n10478 ASIG5V.n10477 0.0154799
R59309 ASIG5V.n10923 ASIG5V.n10469 0.0154799
R59310 ASIG5V.n10707 ASIG5V.n10469 0.0154799
R59311 ASIG5V.n9748 ASIG5V.n3163 0.0151165
R59312 ASIG5V.n9191 ASIG5V.n9190 0.0151165
R59313 ASIG5V.n8572 ASIG5V.n8215 0.0149966
R59314 ASIG5V.n11496 ASIG5V.n9964 0.0149966
R59315 ASIG5V.n8571 ASIG5V.n8324 0.0149966
R59316 ASIG5V.n11497 ASIG5V.n9962 0.0149966
R59317 ASIG5V.n9184 ASIG5V.n6434 0.014845
R59318 ASIG5V.n9183 ASIG5V.n6436 0.014845
R59319 ASIG5V.n10699 ASIG5V.n10481 0.014755
R59320 ASIG5V.n10707 ASIG5V.n10706 0.014755
R59321 ASIG5V.n12283 ASIG5V.n12282 0.0145752
R59322 ASIG5V.n11806 ASIG5V.n1826 0.0145752
R59323 ASIG5V.n12309 ASIG5V.n522 0.0145134
R59324 ASIG5V.n11793 ASIG5V.n1846 0.0145134
R59325 ASIG5V.n12308 ASIG5V.n523 0.0145134
R59326 ASIG5V.n11794 ASIG5V.n1844 0.0145134
R59327 ASIG5V.n11999 ASIG5V.n1673 0.014452
R59328 ASIG5V.n1860 ASIG5V.n1673 0.014452
R59329 ASIG5V.n12000 ASIG5V.n1671 0.014452
R59330 ASIG5V.n1859 ASIG5V.n1671 0.014452
R59331 ASIG5V.n10715 ASIG5V.n10693 0.01445
R59332 ASIG5V.n10717 ASIG5V.n10716 0.01445
R59333 ASIG5V.n10718 ASIG5V.n10717 0.01445
R59334 ASIG5V.n10719 ASIG5V.n10718 0.01445
R59335 ASIG5V.n10720 ASIG5V.n10719 0.01445
R59336 ASIG5V.n10721 ASIG5V.n10720 0.01445
R59337 ASIG5V.n10722 ASIG5V.n10721 0.01445
R59338 ASIG5V.n10723 ASIG5V.n10722 0.01445
R59339 ASIG5V.n10724 ASIG5V.n10723 0.01445
R59340 ASIG5V.n10725 ASIG5V.n10724 0.01445
R59341 ASIG5V.n10726 ASIG5V.n10725 0.01445
R59342 ASIG5V.n10727 ASIG5V.n10726 0.01445
R59343 ASIG5V.n10728 ASIG5V.n10727 0.01445
R59344 ASIG5V.n10729 ASIG5V.n10728 0.01445
R59345 ASIG5V.n10730 ASIG5V.n10729 0.01445
R59346 ASIG5V.n10731 ASIG5V.n10730 0.01445
R59347 ASIG5V.n10732 ASIG5V.n10731 0.01445
R59348 ASIG5V.n10733 ASIG5V.n10732 0.01445
R59349 ASIG5V.n10734 ASIG5V.n10733 0.01445
R59350 ASIG5V.n10735 ASIG5V.n10734 0.01445
R59351 ASIG5V.n10736 ASIG5V.n10735 0.01445
R59352 ASIG5V.n10737 ASIG5V.n10736 0.01445
R59353 ASIG5V.n10738 ASIG5V.n10737 0.01445
R59354 ASIG5V.n10739 ASIG5V.n10738 0.01445
R59355 ASIG5V.n10740 ASIG5V.n10739 0.01445
R59356 ASIG5V.n10741 ASIG5V.n10740 0.01445
R59357 ASIG5V.n10742 ASIG5V.n10741 0.01445
R59358 ASIG5V.n10743 ASIG5V.n10742 0.01445
R59359 ASIG5V.n10744 ASIG5V.n10743 0.01445
R59360 ASIG5V.n10745 ASIG5V.n10744 0.01445
R59361 ASIG5V.n10746 ASIG5V.n10745 0.01445
R59362 ASIG5V.n10747 ASIG5V.n10746 0.01445
R59363 ASIG5V.n10748 ASIG5V.n10747 0.01445
R59364 ASIG5V.n10749 ASIG5V.n10748 0.01445
R59365 ASIG5V.n10750 ASIG5V.n10749 0.01445
R59366 ASIG5V.n10751 ASIG5V.n10750 0.01445
R59367 ASIG5V.n10752 ASIG5V.n10751 0.01445
R59368 ASIG5V.n10753 ASIG5V.n10752 0.01445
R59369 ASIG5V.n10754 ASIG5V.n10753 0.01445
R59370 ASIG5V.n10755 ASIG5V.n10754 0.01445
R59371 ASIG5V.n10756 ASIG5V.n10755 0.01445
R59372 ASIG5V.n10757 ASIG5V.n10756 0.01445
R59373 ASIG5V.n10758 ASIG5V.n10757 0.01445
R59374 ASIG5V.n10759 ASIG5V.n10758 0.01445
R59375 ASIG5V.n10760 ASIG5V.n10759 0.01445
R59376 ASIG5V.n10761 ASIG5V.n10760 0.01445
R59377 ASIG5V.n10762 ASIG5V.n10761 0.01445
R59378 ASIG5V.n10763 ASIG5V.n10762 0.01445
R59379 ASIG5V.n10764 ASIG5V.n10763 0.01445
R59380 ASIG5V.n10765 ASIG5V.n10764 0.01445
R59381 ASIG5V.n10766 ASIG5V.n10765 0.01445
R59382 ASIG5V.n10767 ASIG5V.n10766 0.01445
R59383 ASIG5V.n10768 ASIG5V.n10767 0.01445
R59384 ASIG5V.n10769 ASIG5V.n10768 0.01445
R59385 ASIG5V.n10770 ASIG5V.n10769 0.01445
R59386 ASIG5V.n10771 ASIG5V.n10770 0.01445
R59387 ASIG5V.n10772 ASIG5V.n10771 0.01445
R59388 ASIG5V.n10773 ASIG5V.n10772 0.01445
R59389 ASIG5V.n10774 ASIG5V.n10773 0.01445
R59390 ASIG5V.n10775 ASIG5V.n10774 0.01445
R59391 ASIG5V.n10776 ASIG5V.n10775 0.01445
R59392 ASIG5V.n10777 ASIG5V.n10776 0.01445
R59393 ASIG5V.n10778 ASIG5V.n10777 0.01445
R59394 ASIG5V.n10779 ASIG5V.n10778 0.01445
R59395 ASIG5V.n10780 ASIG5V.n10779 0.01445
R59396 ASIG5V.n10781 ASIG5V.n10780 0.01445
R59397 ASIG5V.n10782 ASIG5V.n10781 0.01445
R59398 ASIG5V.n10783 ASIG5V.n10782 0.01445
R59399 ASIG5V.n10784 ASIG5V.n10783 0.01445
R59400 ASIG5V.n10785 ASIG5V.n10784 0.01445
R59401 ASIG5V.n10786 ASIG5V.n10785 0.01445
R59402 ASIG5V.n10787 ASIG5V.n10786 0.01445
R59403 ASIG5V.n10788 ASIG5V.n10787 0.01445
R59404 ASIG5V.n10789 ASIG5V.n10788 0.01445
R59405 ASIG5V.n10790 ASIG5V.n10789 0.01445
R59406 ASIG5V.n10791 ASIG5V.n10790 0.01445
R59407 ASIG5V.n10792 ASIG5V.n10791 0.01445
R59408 ASIG5V.n10793 ASIG5V.n10792 0.01445
R59409 ASIG5V.n10794 ASIG5V.n10793 0.01445
R59410 ASIG5V.n10795 ASIG5V.n10794 0.01445
R59411 ASIG5V.n10796 ASIG5V.n10795 0.01445
R59412 ASIG5V.n10797 ASIG5V.n10796 0.01445
R59413 ASIG5V.n10798 ASIG5V.n10797 0.01445
R59414 ASIG5V.n10799 ASIG5V.n10798 0.01445
R59415 ASIG5V.n10800 ASIG5V.n10799 0.01445
R59416 ASIG5V.n10801 ASIG5V.n10800 0.01445
R59417 ASIG5V.n10802 ASIG5V.n10801 0.01445
R59418 ASIG5V.n10803 ASIG5V.n10802 0.01445
R59419 ASIG5V.n10804 ASIG5V.n10803 0.01445
R59420 ASIG5V.n10805 ASIG5V.n10804 0.01445
R59421 ASIG5V.n10806 ASIG5V.n10805 0.01445
R59422 ASIG5V.n10807 ASIG5V.n10806 0.01445
R59423 ASIG5V.n10808 ASIG5V.n10807 0.01445
R59424 ASIG5V.n10809 ASIG5V.n10808 0.01445
R59425 ASIG5V.n10810 ASIG5V.n10809 0.01445
R59426 ASIG5V.n10811 ASIG5V.n10810 0.01445
R59427 ASIG5V.n10812 ASIG5V.n10811 0.01445
R59428 ASIG5V.n10812 ASIG5V.n10489 0.01445
R59429 ASIG5V.n10714 ASIG5V.n10694 0.01445
R59430 ASIG5V.n10909 ASIG5V.n10692 0.01445
R59431 ASIG5V.n10909 ASIG5V.n10908 0.01445
R59432 ASIG5V.n10908 ASIG5V.n10907 0.01445
R59433 ASIG5V.n10907 ASIG5V.n10906 0.01445
R59434 ASIG5V.n10906 ASIG5V.n10905 0.01445
R59435 ASIG5V.n10905 ASIG5V.n10904 0.01445
R59436 ASIG5V.n10904 ASIG5V.n10903 0.01445
R59437 ASIG5V.n10903 ASIG5V.n10902 0.01445
R59438 ASIG5V.n10902 ASIG5V.n10901 0.01445
R59439 ASIG5V.n10901 ASIG5V.n10900 0.01445
R59440 ASIG5V.n10900 ASIG5V.n10899 0.01445
R59441 ASIG5V.n10899 ASIG5V.n10898 0.01445
R59442 ASIG5V.n10898 ASIG5V.n10897 0.01445
R59443 ASIG5V.n10897 ASIG5V.n10896 0.01445
R59444 ASIG5V.n10896 ASIG5V.n10895 0.01445
R59445 ASIG5V.n10895 ASIG5V.n10894 0.01445
R59446 ASIG5V.n10894 ASIG5V.n10893 0.01445
R59447 ASIG5V.n10893 ASIG5V.n10892 0.01445
R59448 ASIG5V.n10892 ASIG5V.n10891 0.01445
R59449 ASIG5V.n10891 ASIG5V.n10890 0.01445
R59450 ASIG5V.n10890 ASIG5V.n10889 0.01445
R59451 ASIG5V.n10889 ASIG5V.n10888 0.01445
R59452 ASIG5V.n10888 ASIG5V.n10887 0.01445
R59453 ASIG5V.n10887 ASIG5V.n10886 0.01445
R59454 ASIG5V.n10886 ASIG5V.n10885 0.01445
R59455 ASIG5V.n10885 ASIG5V.n10884 0.01445
R59456 ASIG5V.n10884 ASIG5V.n10883 0.01445
R59457 ASIG5V.n10883 ASIG5V.n10882 0.01445
R59458 ASIG5V.n10882 ASIG5V.n10881 0.01445
R59459 ASIG5V.n10881 ASIG5V.n10880 0.01445
R59460 ASIG5V.n10880 ASIG5V.n10879 0.01445
R59461 ASIG5V.n10879 ASIG5V.n10878 0.01445
R59462 ASIG5V.n10878 ASIG5V.n10877 0.01445
R59463 ASIG5V.n10877 ASIG5V.n10876 0.01445
R59464 ASIG5V.n10876 ASIG5V.n10875 0.01445
R59465 ASIG5V.n10875 ASIG5V.n10874 0.01445
R59466 ASIG5V.n10874 ASIG5V.n10873 0.01445
R59467 ASIG5V.n10873 ASIG5V.n10872 0.01445
R59468 ASIG5V.n10872 ASIG5V.n10871 0.01445
R59469 ASIG5V.n10871 ASIG5V.n10870 0.01445
R59470 ASIG5V.n10870 ASIG5V.n10869 0.01445
R59471 ASIG5V.n10869 ASIG5V.n10868 0.01445
R59472 ASIG5V.n10868 ASIG5V.n10867 0.01445
R59473 ASIG5V.n10867 ASIG5V.n10866 0.01445
R59474 ASIG5V.n10866 ASIG5V.n10865 0.01445
R59475 ASIG5V.n10865 ASIG5V.n10864 0.01445
R59476 ASIG5V.n10864 ASIG5V.n10863 0.01445
R59477 ASIG5V.n10863 ASIG5V.n10862 0.01445
R59478 ASIG5V.n10862 ASIG5V.n10861 0.01445
R59479 ASIG5V.n10861 ASIG5V.n10860 0.01445
R59480 ASIG5V.n10860 ASIG5V.n10859 0.01445
R59481 ASIG5V.n10859 ASIG5V.n10858 0.01445
R59482 ASIG5V.n10858 ASIG5V.n10857 0.01445
R59483 ASIG5V.n10857 ASIG5V.n10856 0.01445
R59484 ASIG5V.n10856 ASIG5V.n10855 0.01445
R59485 ASIG5V.n10855 ASIG5V.n10854 0.01445
R59486 ASIG5V.n10854 ASIG5V.n10853 0.01445
R59487 ASIG5V.n10853 ASIG5V.n10852 0.01445
R59488 ASIG5V.n10852 ASIG5V.n10851 0.01445
R59489 ASIG5V.n10851 ASIG5V.n10850 0.01445
R59490 ASIG5V.n10850 ASIG5V.n10849 0.01445
R59491 ASIG5V.n10849 ASIG5V.n10848 0.01445
R59492 ASIG5V.n10848 ASIG5V.n10847 0.01445
R59493 ASIG5V.n10847 ASIG5V.n10846 0.01445
R59494 ASIG5V.n10846 ASIG5V.n10845 0.01445
R59495 ASIG5V.n10845 ASIG5V.n10844 0.01445
R59496 ASIG5V.n10844 ASIG5V.n10843 0.01445
R59497 ASIG5V.n10843 ASIG5V.n10842 0.01445
R59498 ASIG5V.n10842 ASIG5V.n10841 0.01445
R59499 ASIG5V.n10841 ASIG5V.n10840 0.01445
R59500 ASIG5V.n10840 ASIG5V.n10839 0.01445
R59501 ASIG5V.n10839 ASIG5V.n10838 0.01445
R59502 ASIG5V.n10838 ASIG5V.n10837 0.01445
R59503 ASIG5V.n10837 ASIG5V.n10836 0.01445
R59504 ASIG5V.n10836 ASIG5V.n10835 0.01445
R59505 ASIG5V.n10835 ASIG5V.n10834 0.01445
R59506 ASIG5V.n10834 ASIG5V.n10833 0.01445
R59507 ASIG5V.n10833 ASIG5V.n10832 0.01445
R59508 ASIG5V.n10832 ASIG5V.n10831 0.01445
R59509 ASIG5V.n10831 ASIG5V.n10830 0.01445
R59510 ASIG5V.n10830 ASIG5V.n10829 0.01445
R59511 ASIG5V.n10829 ASIG5V.n10828 0.01445
R59512 ASIG5V.n10828 ASIG5V.n10827 0.01445
R59513 ASIG5V.n10827 ASIG5V.n10826 0.01445
R59514 ASIG5V.n10826 ASIG5V.n10825 0.01445
R59515 ASIG5V.n10825 ASIG5V.n10824 0.01445
R59516 ASIG5V.n10824 ASIG5V.n10823 0.01445
R59517 ASIG5V.n10823 ASIG5V.n10822 0.01445
R59518 ASIG5V.n10822 ASIG5V.n10821 0.01445
R59519 ASIG5V.n10821 ASIG5V.n10820 0.01445
R59520 ASIG5V.n10820 ASIG5V.n10819 0.01445
R59521 ASIG5V.n10819 ASIG5V.n10818 0.01445
R59522 ASIG5V.n10818 ASIG5V.n10817 0.01445
R59523 ASIG5V.n10817 ASIG5V.n10816 0.01445
R59524 ASIG5V.n10816 ASIG5V.n10815 0.01445
R59525 ASIG5V.n10815 ASIG5V.n10814 0.01445
R59526 ASIG5V.n10814 ASIG5V.n10813 0.01445
R59527 ASIG5V.n4263 ASIG5V.n3844 0.01445
R59528 ASIG5V.n4102 ASIG5V.n4101 0.01445
R59529 ASIG5V.n4102 ASIG5V.n4100 0.01445
R59530 ASIG5V.n4106 ASIG5V.n4100 0.01445
R59531 ASIG5V.n4107 ASIG5V.n4106 0.01445
R59532 ASIG5V.n4108 ASIG5V.n4107 0.01445
R59533 ASIG5V.n4108 ASIG5V.n4098 0.01445
R59534 ASIG5V.n4112 ASIG5V.n4098 0.01445
R59535 ASIG5V.n4113 ASIG5V.n4112 0.01445
R59536 ASIG5V.n4114 ASIG5V.n4113 0.01445
R59537 ASIG5V.n4114 ASIG5V.n4096 0.01445
R59538 ASIG5V.n4118 ASIG5V.n4096 0.01445
R59539 ASIG5V.n4119 ASIG5V.n4118 0.01445
R59540 ASIG5V.n4120 ASIG5V.n4119 0.01445
R59541 ASIG5V.n4120 ASIG5V.n4094 0.01445
R59542 ASIG5V.n4124 ASIG5V.n4094 0.01445
R59543 ASIG5V.n4125 ASIG5V.n4124 0.01445
R59544 ASIG5V.n4126 ASIG5V.n4125 0.01445
R59545 ASIG5V.n4126 ASIG5V.n4092 0.01445
R59546 ASIG5V.n4130 ASIG5V.n4092 0.01445
R59547 ASIG5V.n4131 ASIG5V.n4130 0.01445
R59548 ASIG5V.n4132 ASIG5V.n4131 0.01445
R59549 ASIG5V.n4132 ASIG5V.n4090 0.01445
R59550 ASIG5V.n4136 ASIG5V.n4090 0.01445
R59551 ASIG5V.n4137 ASIG5V.n4136 0.01445
R59552 ASIG5V.n4138 ASIG5V.n4137 0.01445
R59553 ASIG5V.n4138 ASIG5V.n4088 0.01445
R59554 ASIG5V.n4142 ASIG5V.n4088 0.01445
R59555 ASIG5V.n4143 ASIG5V.n4142 0.01445
R59556 ASIG5V.n4144 ASIG5V.n4143 0.01445
R59557 ASIG5V.n4144 ASIG5V.n4086 0.01445
R59558 ASIG5V.n4148 ASIG5V.n4086 0.01445
R59559 ASIG5V.n4149 ASIG5V.n4148 0.01445
R59560 ASIG5V.n4150 ASIG5V.n4149 0.01445
R59561 ASIG5V.n4150 ASIG5V.n4084 0.01445
R59562 ASIG5V.n4154 ASIG5V.n4084 0.01445
R59563 ASIG5V.n4155 ASIG5V.n4154 0.01445
R59564 ASIG5V.n4156 ASIG5V.n4155 0.01445
R59565 ASIG5V.n4156 ASIG5V.n4082 0.01445
R59566 ASIG5V.n4160 ASIG5V.n4082 0.01445
R59567 ASIG5V.n4161 ASIG5V.n4160 0.01445
R59568 ASIG5V.n4162 ASIG5V.n4161 0.01445
R59569 ASIG5V.n4162 ASIG5V.n4080 0.01445
R59570 ASIG5V.n4166 ASIG5V.n4080 0.01445
R59571 ASIG5V.n4167 ASIG5V.n4166 0.01445
R59572 ASIG5V.n4168 ASIG5V.n4167 0.01445
R59573 ASIG5V.n4168 ASIG5V.n4078 0.01445
R59574 ASIG5V.n4172 ASIG5V.n4078 0.01445
R59575 ASIG5V.n4173 ASIG5V.n4172 0.01445
R59576 ASIG5V.n4174 ASIG5V.n4173 0.01445
R59577 ASIG5V.n4174 ASIG5V.n4076 0.01445
R59578 ASIG5V.n4178 ASIG5V.n4076 0.01445
R59579 ASIG5V.n4179 ASIG5V.n4178 0.01445
R59580 ASIG5V.n4180 ASIG5V.n4179 0.01445
R59581 ASIG5V.n4180 ASIG5V.n4074 0.01445
R59582 ASIG5V.n4184 ASIG5V.n4074 0.01445
R59583 ASIG5V.n4185 ASIG5V.n4184 0.01445
R59584 ASIG5V.n4186 ASIG5V.n4185 0.01445
R59585 ASIG5V.n4186 ASIG5V.n4072 0.01445
R59586 ASIG5V.n4190 ASIG5V.n4072 0.01445
R59587 ASIG5V.n4191 ASIG5V.n4190 0.01445
R59588 ASIG5V.n4192 ASIG5V.n4191 0.01445
R59589 ASIG5V.n4192 ASIG5V.n4070 0.01445
R59590 ASIG5V.n4196 ASIG5V.n4070 0.01445
R59591 ASIG5V.n4197 ASIG5V.n4196 0.01445
R59592 ASIG5V.n4198 ASIG5V.n4197 0.01445
R59593 ASIG5V.n4198 ASIG5V.n4068 0.01445
R59594 ASIG5V.n4202 ASIG5V.n4068 0.01445
R59595 ASIG5V.n4203 ASIG5V.n4202 0.01445
R59596 ASIG5V.n4204 ASIG5V.n4203 0.01445
R59597 ASIG5V.n4204 ASIG5V.n4066 0.01445
R59598 ASIG5V.n4208 ASIG5V.n4066 0.01445
R59599 ASIG5V.n4209 ASIG5V.n4208 0.01445
R59600 ASIG5V.n4210 ASIG5V.n4209 0.01445
R59601 ASIG5V.n4210 ASIG5V.n4064 0.01445
R59602 ASIG5V.n4214 ASIG5V.n4064 0.01445
R59603 ASIG5V.n4215 ASIG5V.n4214 0.01445
R59604 ASIG5V.n4216 ASIG5V.n4215 0.01445
R59605 ASIG5V.n4216 ASIG5V.n4062 0.01445
R59606 ASIG5V.n4220 ASIG5V.n4062 0.01445
R59607 ASIG5V.n4221 ASIG5V.n4220 0.01445
R59608 ASIG5V.n4222 ASIG5V.n4221 0.01445
R59609 ASIG5V.n4222 ASIG5V.n4060 0.01445
R59610 ASIG5V.n4226 ASIG5V.n4060 0.01445
R59611 ASIG5V.n4227 ASIG5V.n4226 0.01445
R59612 ASIG5V.n4228 ASIG5V.n4227 0.01445
R59613 ASIG5V.n4228 ASIG5V.n4058 0.01445
R59614 ASIG5V.n4232 ASIG5V.n4058 0.01445
R59615 ASIG5V.n4233 ASIG5V.n4232 0.01445
R59616 ASIG5V.n4234 ASIG5V.n4233 0.01445
R59617 ASIG5V.n4234 ASIG5V.n4056 0.01445
R59618 ASIG5V.n4238 ASIG5V.n4056 0.01445
R59619 ASIG5V.n4239 ASIG5V.n4238 0.01445
R59620 ASIG5V.n4240 ASIG5V.n4239 0.01445
R59621 ASIG5V.n4240 ASIG5V.n4054 0.01445
R59622 ASIG5V.n4244 ASIG5V.n4054 0.01445
R59623 ASIG5V.n4245 ASIG5V.n4244 0.01445
R59624 ASIG5V.n4246 ASIG5V.n4245 0.01445
R59625 ASIG5V.n4262 ASIG5V.n3845 0.01445
R59626 ASIG5V.n4103 ASIG5V.n3856 0.01445
R59627 ASIG5V.n4104 ASIG5V.n4103 0.01445
R59628 ASIG5V.n4105 ASIG5V.n4104 0.01445
R59629 ASIG5V.n4105 ASIG5V.n4099 0.01445
R59630 ASIG5V.n4109 ASIG5V.n4099 0.01445
R59631 ASIG5V.n4110 ASIG5V.n4109 0.01445
R59632 ASIG5V.n4111 ASIG5V.n4110 0.01445
R59633 ASIG5V.n4111 ASIG5V.n4097 0.01445
R59634 ASIG5V.n4115 ASIG5V.n4097 0.01445
R59635 ASIG5V.n4116 ASIG5V.n4115 0.01445
R59636 ASIG5V.n4117 ASIG5V.n4116 0.01445
R59637 ASIG5V.n4117 ASIG5V.n4095 0.01445
R59638 ASIG5V.n4121 ASIG5V.n4095 0.01445
R59639 ASIG5V.n4122 ASIG5V.n4121 0.01445
R59640 ASIG5V.n4123 ASIG5V.n4122 0.01445
R59641 ASIG5V.n4123 ASIG5V.n4093 0.01445
R59642 ASIG5V.n4127 ASIG5V.n4093 0.01445
R59643 ASIG5V.n4128 ASIG5V.n4127 0.01445
R59644 ASIG5V.n4129 ASIG5V.n4128 0.01445
R59645 ASIG5V.n4129 ASIG5V.n4091 0.01445
R59646 ASIG5V.n4133 ASIG5V.n4091 0.01445
R59647 ASIG5V.n4134 ASIG5V.n4133 0.01445
R59648 ASIG5V.n4135 ASIG5V.n4134 0.01445
R59649 ASIG5V.n4135 ASIG5V.n4089 0.01445
R59650 ASIG5V.n4139 ASIG5V.n4089 0.01445
R59651 ASIG5V.n4140 ASIG5V.n4139 0.01445
R59652 ASIG5V.n4141 ASIG5V.n4140 0.01445
R59653 ASIG5V.n4141 ASIG5V.n4087 0.01445
R59654 ASIG5V.n4145 ASIG5V.n4087 0.01445
R59655 ASIG5V.n4146 ASIG5V.n4145 0.01445
R59656 ASIG5V.n4147 ASIG5V.n4146 0.01445
R59657 ASIG5V.n4147 ASIG5V.n4085 0.01445
R59658 ASIG5V.n4151 ASIG5V.n4085 0.01445
R59659 ASIG5V.n4152 ASIG5V.n4151 0.01445
R59660 ASIG5V.n4153 ASIG5V.n4152 0.01445
R59661 ASIG5V.n4153 ASIG5V.n4083 0.01445
R59662 ASIG5V.n4157 ASIG5V.n4083 0.01445
R59663 ASIG5V.n4158 ASIG5V.n4157 0.01445
R59664 ASIG5V.n4159 ASIG5V.n4158 0.01445
R59665 ASIG5V.n4159 ASIG5V.n4081 0.01445
R59666 ASIG5V.n4163 ASIG5V.n4081 0.01445
R59667 ASIG5V.n4164 ASIG5V.n4163 0.01445
R59668 ASIG5V.n4165 ASIG5V.n4164 0.01445
R59669 ASIG5V.n4165 ASIG5V.n4079 0.01445
R59670 ASIG5V.n4169 ASIG5V.n4079 0.01445
R59671 ASIG5V.n4170 ASIG5V.n4169 0.01445
R59672 ASIG5V.n4171 ASIG5V.n4170 0.01445
R59673 ASIG5V.n4171 ASIG5V.n4077 0.01445
R59674 ASIG5V.n4175 ASIG5V.n4077 0.01445
R59675 ASIG5V.n4176 ASIG5V.n4175 0.01445
R59676 ASIG5V.n4177 ASIG5V.n4176 0.01445
R59677 ASIG5V.n4177 ASIG5V.n4075 0.01445
R59678 ASIG5V.n4181 ASIG5V.n4075 0.01445
R59679 ASIG5V.n4182 ASIG5V.n4181 0.01445
R59680 ASIG5V.n4183 ASIG5V.n4182 0.01445
R59681 ASIG5V.n4183 ASIG5V.n4073 0.01445
R59682 ASIG5V.n4187 ASIG5V.n4073 0.01445
R59683 ASIG5V.n4188 ASIG5V.n4187 0.01445
R59684 ASIG5V.n4189 ASIG5V.n4188 0.01445
R59685 ASIG5V.n4189 ASIG5V.n4071 0.01445
R59686 ASIG5V.n4193 ASIG5V.n4071 0.01445
R59687 ASIG5V.n4194 ASIG5V.n4193 0.01445
R59688 ASIG5V.n4195 ASIG5V.n4194 0.01445
R59689 ASIG5V.n4195 ASIG5V.n4069 0.01445
R59690 ASIG5V.n4199 ASIG5V.n4069 0.01445
R59691 ASIG5V.n4200 ASIG5V.n4199 0.01445
R59692 ASIG5V.n4201 ASIG5V.n4200 0.01445
R59693 ASIG5V.n4201 ASIG5V.n4067 0.01445
R59694 ASIG5V.n4205 ASIG5V.n4067 0.01445
R59695 ASIG5V.n4206 ASIG5V.n4205 0.01445
R59696 ASIG5V.n4207 ASIG5V.n4206 0.01445
R59697 ASIG5V.n4207 ASIG5V.n4065 0.01445
R59698 ASIG5V.n4211 ASIG5V.n4065 0.01445
R59699 ASIG5V.n4212 ASIG5V.n4211 0.01445
R59700 ASIG5V.n4213 ASIG5V.n4212 0.01445
R59701 ASIG5V.n4213 ASIG5V.n4063 0.01445
R59702 ASIG5V.n4217 ASIG5V.n4063 0.01445
R59703 ASIG5V.n4218 ASIG5V.n4217 0.01445
R59704 ASIG5V.n4219 ASIG5V.n4218 0.01445
R59705 ASIG5V.n4219 ASIG5V.n4061 0.01445
R59706 ASIG5V.n4223 ASIG5V.n4061 0.01445
R59707 ASIG5V.n4224 ASIG5V.n4223 0.01445
R59708 ASIG5V.n4225 ASIG5V.n4224 0.01445
R59709 ASIG5V.n4225 ASIG5V.n4059 0.01445
R59710 ASIG5V.n4229 ASIG5V.n4059 0.01445
R59711 ASIG5V.n4230 ASIG5V.n4229 0.01445
R59712 ASIG5V.n4231 ASIG5V.n4230 0.01445
R59713 ASIG5V.n4231 ASIG5V.n4057 0.01445
R59714 ASIG5V.n4235 ASIG5V.n4057 0.01445
R59715 ASIG5V.n4236 ASIG5V.n4235 0.01445
R59716 ASIG5V.n4237 ASIG5V.n4236 0.01445
R59717 ASIG5V.n4237 ASIG5V.n4055 0.01445
R59718 ASIG5V.n4241 ASIG5V.n4055 0.01445
R59719 ASIG5V.n4242 ASIG5V.n4241 0.01445
R59720 ASIG5V.n4243 ASIG5V.n4242 0.01445
R59721 ASIG5V.n4243 ASIG5V.n4053 0.01445
R59722 ASIG5V.n4252 ASIG5V.n4053 0.01445
R59723 ASIG5V.n4265 ASIG5V.n4264 0.0143045
R59724 ASIG5V.n9425 ASIG5V.n5457 0.014225
R59725 ASIG5V.n9178 ASIG5V.n6434 0.014059
R59726 ASIG5V.n9179 ASIG5V.n6436 0.014059
R59727 ASIG5V.n6534 ASIG5V.n6416 0.0140338
R59728 ASIG5V.n7244 ASIG5V.n7243 0.0140338
R59729 ASIG5V.n10475 ASIG5V.n10022 0.0140338
R59730 ASIG5V.n4577 ASIG5V.n3779 0.0140302
R59731 ASIG5V.n9398 ASIG5V.n5911 0.0140302
R59732 ASIG5V.n4576 ASIG5V.n3782 0.0140302
R59733 ASIG5V.n9399 ASIG5V.n5910 0.0140302
R59734 ASIG5V.n12316 ASIG5V.n505 0.013775
R59735 ASIG5V.n11490 ASIG5V.n11489 0.013775
R59736 ASIG5V.n9188 ASIG5V.n6308 0.013547
R59737 ASIG5V.n9189 ASIG5V.n6428 0.013547
R59738 ASIG5V.n4793 ASIG5V.n3267 0.0134925
R59739 ASIG5V.n7964 ASIG5V.n5120 0.0134925
R59740 ASIG5V.n510 ASIG5V.n7 0.013325
R59741 ASIG5V.n10368 ASIG5V.n10367 0.013325
R59742 ASIG5V.n12280 ASIG5V.n873 0.0130638
R59743 ASIG5V.n1834 ASIG5V.n1719 0.0130638
R59744 ASIG5V.n12281 ASIG5V.n871 0.0130638
R59745 ASIG5V.n1836 ASIG5V.n1835 0.0130638
R59746 ASIG5V.n8587 ASIG5V.n8586 0.0129511
R59747 ASIG5V.n9954 ASIG5V.n9953 0.0129511
R59748 ASIG5V.n9954 ASIG5V.n3002 0.0129511
R59749 ASIG5V.n9739 ASIG5V.n9738 0.012875
R59750 ASIG5V.n4267 ASIG5V.n3841 0.0128221
R59751 ASIG5V.n4266 ASIG5V.n3842 0.0128221
R59752 ASIG5V.n7241 ASIG5V.n6893 0.0125805
R59753 ASIG5V.n10473 ASIG5V.n10024 0.0125805
R59754 ASIG5V.n7242 ASIG5V.n6895 0.0125805
R59755 ASIG5V.n10474 ASIG5V.n10023 0.0125805
R59756 ASIG5V.n5459 ASIG5V.n5167 0.0124869
R59757 ASIG5V.n5461 ASIG5V.n5460 0.0124869
R59758 ASIG5V.n12330 ASIG5V.n12329 0.0124098
R59759 ASIG5V.n2562 ASIG5V.n2561 0.0124098
R59760 ASIG5V.n10706 ASIG5V.n10705 0.0123125
R59761 ASIG5V.n10699 ASIG5V.n10698 0.0123125
R59762 ASIG5V.n3852 ASIG5V.n3842 0.0123125
R59763 ASIG5V.n3853 ASIG5V.n3841 0.0123125
R59764 ASIG5V.n4810 ASIG5V.n4809 0.0120973
R59765 ASIG5V.n7966 ASIG5V.n5122 0.0120973
R59766 ASIG5V.n4814 ASIG5V.n3268 0.0120973
R59767 ASIG5V.n7965 ASIG5V.n5121 0.0120973
R59768 ASIG5V.n515 ASIG5V.n217 0.0120939
R59769 ASIG5V.n11487 ASIG5V.n9967 0.0120939
R59770 ASIG5V.n517 ASIG5V.n516 0.0120939
R59771 ASIG5V.n11488 ASIG5V.n9968 0.0120939
R59772 ASIG5V.n10914 ASIG5V.n10489 0.011975
R59773 ASIG5V.n4248 ASIG5V.n4246 0.011975
R59774 ASIG5V.n9888 ASIG5V.n3080 0.0119575
R59775 ASIG5V.n9884 ASIG5V.n9883 0.0119575
R59776 ASIG5V.n3084 ASIG5V.n3079 0.0119575
R59777 ASIG5V.n9891 ASIG5V.n3082 0.0119575
R59778 ASIG5V.n7472 ASIG5V.n7471 0.0119575
R59779 ASIG5V.n8103 ASIG5V.n8101 0.0119575
R59780 ASIG5V.n8102 ASIG5V.n7470 0.0119575
R59781 ASIG5V.n8107 ASIG5V.n7468 0.0119575
R59782 ASIG5V.n8108 ASIG5V.n7466 0.0119575
R59783 ASIG5V.n8114 ASIG5V.n8112 0.0119575
R59784 ASIG5V.n8113 ASIG5V.n7465 0.0119575
R59785 ASIG5V.n8116 ASIG5V.n7462 0.0119575
R59786 ASIG5V.n8118 ASIG5V.n7461 0.0119575
R59787 ASIG5V.n8120 ASIG5V.n7322 0.0119575
R59788 ASIG5V.n8119 ASIG5V.n7320 0.0119575
R59789 ASIG5V.n8124 ASIG5V.n7323 0.0119575
R59790 ASIG5V.n7326 ASIG5V.n7324 0.0119575
R59791 ASIG5V.n7453 ASIG5V.n7452 0.0119575
R59792 ASIG5V.n7451 ASIG5V.n7325 0.0119575
R59793 ASIG5V.n7450 ASIG5V.n7449 0.0119575
R59794 ASIG5V.n7330 ASIG5V.n7327 0.0119575
R59795 ASIG5V.n7442 ASIG5V.n7441 0.0119575
R59796 ASIG5V.n7440 ASIG5V.n7329 0.0119575
R59797 ASIG5V.n7439 ASIG5V.n7438 0.0119575
R59798 ASIG5V.n7334 ASIG5V.n7331 0.0119575
R59799 ASIG5V.n7431 ASIG5V.n7430 0.0119575
R59800 ASIG5V.n7429 ASIG5V.n7333 0.0119575
R59801 ASIG5V.n7428 ASIG5V.n7427 0.0119575
R59802 ASIG5V.n7416 ASIG5V.n7335 0.0119575
R59803 ASIG5V.n7420 ASIG5V.n7419 0.0119575
R59804 ASIG5V.n7418 ASIG5V.n7415 0.0119575
R59805 ASIG5V.n7417 ASIG5V.n1841 0.0119575
R59806 ASIG5V.n7471 ASIG5V.n3083 0.0119575
R59807 ASIG5V.n8101 ASIG5V.n7472 0.0119575
R59808 ASIG5V.n8103 ASIG5V.n8102 0.0119575
R59809 ASIG5V.n7470 ASIG5V.n7468 0.0119575
R59810 ASIG5V.n9888 ASIG5V.n3081 0.0119575
R59811 ASIG5V.n9884 ASIG5V.n3080 0.0119575
R59812 ASIG5V.n9883 ASIG5V.n3084 0.0119575
R59813 ASIG5V.n3082 ASIG5V.n3079 0.0119575
R59814 ASIG5V.n8109 ASIG5V.n8108 0.0119575
R59815 ASIG5V.n8112 ASIG5V.n7466 0.0119575
R59816 ASIG5V.n8114 ASIG5V.n8113 0.0119575
R59817 ASIG5V.n7465 ASIG5V.n7462 0.0119575
R59818 ASIG5V.n3090 ASIG5V.n3086 0.0119575
R59819 ASIG5V.n9878 ASIG5V.n9877 0.0119575
R59820 ASIG5V.n9880 ASIG5V.n3089 0.0119575
R59821 ASIG5V.n9881 ASIG5V.n3088 0.0119575
R59822 ASIG5V.n7478 ASIG5V.n7474 0.0119575
R59823 ASIG5V.n8094 ASIG5V.n8093 0.0119575
R59824 ASIG5V.n8096 ASIG5V.n7477 0.0119575
R59825 ASIG5V.n8097 ASIG5V.n7476 0.0119575
R59826 ASIG5V.n7632 ASIG5V.n7631 0.0119575
R59827 ASIG5V.n7628 ASIG5V.n7622 0.0119575
R59828 ASIG5V.n7627 ASIG5V.n7626 0.0119575
R59829 ASIG5V.n7624 ASIG5V.n7621 0.0119575
R59830 ASIG5V.n7314 ASIG5V.n7312 0.0119575
R59831 ASIG5V.n8127 ASIG5V.n7316 0.0119575
R59832 ASIG5V.n7317 ASIG5V.n7311 0.0119575
R59833 ASIG5V.n8129 ASIG5V.n7308 0.0119575
R59834 ASIG5V.n7306 ASIG5V.n7305 0.0119575
R59835 ASIG5V.n8133 ASIG5V.n7301 0.0119575
R59836 ASIG5V.n8132 ASIG5V.n7299 0.0119575
R59837 ASIG5V.n8137 ASIG5V.n7302 0.0119575
R59838 ASIG5V.n7370 ASIG5V.n7368 0.0119575
R59839 ASIG5V.n7373 ASIG5V.n7371 0.0119575
R59840 ASIG5V.n7372 ASIG5V.n7367 0.0119575
R59841 ASIG5V.n7377 ASIG5V.n7364 0.0119575
R59842 ASIG5V.n7363 ASIG5V.n7362 0.0119575
R59843 ASIG5V.n7381 ASIG5V.n7359 0.0119575
R59844 ASIG5V.n7380 ASIG5V.n7357 0.0119575
R59845 ASIG5V.n7385 ASIG5V.n7360 0.0119575
R59846 ASIG5V.n7343 ASIG5V.n7337 0.0119575
R59847 ASIG5V.n7409 ASIG5V.n7408 0.0119575
R59848 ASIG5V.n7411 ASIG5V.n7342 0.0119575
R59849 ASIG5V.n7412 ASIG5V.n7341 0.0119575
R59850 ASIG5V.n7633 ASIG5V.n7632 0.0119575
R59851 ASIG5V.n7631 ASIG5V.n7622 0.0119575
R59852 ASIG5V.n7628 ASIG5V.n7627 0.0119575
R59853 ASIG5V.n7626 ASIG5V.n7621 0.0119575
R59854 ASIG5V.n7478 ASIG5V.n7475 0.0119575
R59855 ASIG5V.n8094 ASIG5V.n7474 0.0119575
R59856 ASIG5V.n8093 ASIG5V.n7477 0.0119575
R59857 ASIG5V.n8097 ASIG5V.n8096 0.0119575
R59858 ASIG5V.n3090 ASIG5V.n3087 0.0119575
R59859 ASIG5V.n9878 ASIG5V.n3086 0.0119575
R59860 ASIG5V.n9877 ASIG5V.n3089 0.0119575
R59861 ASIG5V.n9881 ASIG5V.n9880 0.0119575
R59862 ASIG5V.n7315 ASIG5V.n7314 0.0119575
R59863 ASIG5V.n8118 ASIG5V.n8117 0.0119575
R59864 ASIG5V.n7316 ASIG5V.n7312 0.0119575
R59865 ASIG5V.n7461 ASIG5V.n7322 0.0119575
R59866 ASIG5V.n8120 ASIG5V.n8119 0.0119575
R59867 ASIG5V.n8127 ASIG5V.n7317 0.0119575
R59868 ASIG5V.n7323 ASIG5V.n7320 0.0119575
R59869 ASIG5V.n7311 ASIG5V.n7308 0.0119575
R59870 ASIG5V.n3097 ASIG5V.n3093 0.0119575
R59871 ASIG5V.n9869 ASIG5V.n9868 0.0119575
R59872 ASIG5V.n9871 ASIG5V.n3096 0.0119575
R59873 ASIG5V.n9872 ASIG5V.n3095 0.0119575
R59874 ASIG5V.n7485 ASIG5V.n7481 0.0119575
R59875 ASIG5V.n8085 ASIG5V.n8084 0.0119575
R59876 ASIG5V.n8087 ASIG5V.n7484 0.0119575
R59877 ASIG5V.n8088 ASIG5V.n7483 0.0119575
R59878 ASIG5V.n7620 ASIG5V.n7619 0.0119575
R59879 ASIG5V.n7639 ASIG5V.n7572 0.0119575
R59880 ASIG5V.n7638 ASIG5V.n7570 0.0119575
R59881 ASIG5V.n7643 ASIG5V.n7573 0.0119575
R59882 ASIG5V.n7613 ASIG5V.n7574 0.0119575
R59883 ASIG5V.n7614 ASIG5V.n7612 0.0119575
R59884 ASIG5V.n7609 ASIG5V.n7606 0.0119575
R59885 ASIG5V.n7607 ASIG5V.n7605 0.0119575
R59886 ASIG5V.n7293 ASIG5V.n7291 0.0119575
R59887 ASIG5V.n8140 ASIG5V.n7295 0.0119575
R59888 ASIG5V.n7296 ASIG5V.n7290 0.0119575
R59889 ASIG5V.n8142 ASIG5V.n7288 0.0119575
R59890 ASIG5V.n7286 ASIG5V.n7285 0.0119575
R59891 ASIG5V.n8146 ASIG5V.n7281 0.0119575
R59892 ASIG5V.n8145 ASIG5V.n7279 0.0119575
R59893 ASIG5V.n8150 ASIG5V.n7282 0.0119575
R59894 ASIG5V.n7388 ASIG5V.n7352 0.0119575
R59895 ASIG5V.n7389 ASIG5V.n7351 0.0119575
R59896 ASIG5V.n7353 ASIG5V.n7349 0.0119575
R59897 ASIG5V.n7391 ASIG5V.n7347 0.0119575
R59898 ASIG5V.n7394 ASIG5V.n7346 0.0119575
R59899 ASIG5V.n7400 ASIG5V.n7399 0.0119575
R59900 ASIG5V.n7402 ASIG5V.n7393 0.0119575
R59901 ASIG5V.n7403 ASIG5V.n169 0.0119575
R59902 ASIG5V.n7617 ASIG5V.n7574 0.0119575
R59903 ASIG5V.n7614 ASIG5V.n7613 0.0119575
R59904 ASIG5V.n7612 ASIG5V.n7606 0.0119575
R59905 ASIG5V.n7609 ASIG5V.n7605 0.0119575
R59906 ASIG5V.n7636 ASIG5V.n7619 0.0119575
R59907 ASIG5V.n7620 ASIG5V.n7572 0.0119575
R59908 ASIG5V.n7639 ASIG5V.n7638 0.0119575
R59909 ASIG5V.n7573 ASIG5V.n7570 0.0119575
R59910 ASIG5V.n7485 ASIG5V.n7482 0.0119575
R59911 ASIG5V.n8085 ASIG5V.n7481 0.0119575
R59912 ASIG5V.n8084 ASIG5V.n7484 0.0119575
R59913 ASIG5V.n8088 ASIG5V.n8087 0.0119575
R59914 ASIG5V.n3097 ASIG5V.n3094 0.0119575
R59915 ASIG5V.n9869 ASIG5V.n3093 0.0119575
R59916 ASIG5V.n9868 ASIG5V.n3096 0.0119575
R59917 ASIG5V.n9872 ASIG5V.n9871 0.0119575
R59918 ASIG5V.n7294 ASIG5V.n7293 0.0119575
R59919 ASIG5V.n8130 ASIG5V.n7305 0.0119575
R59920 ASIG5V.n7459 ASIG5V.n7324 0.0119575
R59921 ASIG5V.n7295 ASIG5V.n7291 0.0119575
R59922 ASIG5V.n7306 ASIG5V.n7301 0.0119575
R59923 ASIG5V.n7452 ASIG5V.n7326 0.0119575
R59924 ASIG5V.n7453 ASIG5V.n7325 0.0119575
R59925 ASIG5V.n8133 ASIG5V.n8132 0.0119575
R59926 ASIG5V.n8140 ASIG5V.n7296 0.0119575
R59927 ASIG5V.n7451 ASIG5V.n7450 0.0119575
R59928 ASIG5V.n7302 ASIG5V.n7299 0.0119575
R59929 ASIG5V.n7290 ASIG5V.n7288 0.0119575
R59930 ASIG5V.n3104 ASIG5V.n3100 0.0119575
R59931 ASIG5V.n9860 ASIG5V.n9859 0.0119575
R59932 ASIG5V.n9862 ASIG5V.n3103 0.0119575
R59933 ASIG5V.n9863 ASIG5V.n3102 0.0119575
R59934 ASIG5V.n7492 ASIG5V.n7488 0.0119575
R59935 ASIG5V.n8076 ASIG5V.n8075 0.0119575
R59936 ASIG5V.n8078 ASIG5V.n7491 0.0119575
R59937 ASIG5V.n8079 ASIG5V.n7490 0.0119575
R59938 ASIG5V.n7569 ASIG5V.n7568 0.0119575
R59939 ASIG5V.n7648 ASIG5V.n7564 0.0119575
R59940 ASIG5V.n7647 ASIG5V.n7562 0.0119575
R59941 ASIG5V.n7652 ASIG5V.n7565 0.0119575
R59942 ASIG5V.n7600 ASIG5V.n7577 0.0119575
R59943 ASIG5V.n7595 ASIG5V.n7594 0.0119575
R59944 ASIG5V.n7602 ASIG5V.n7596 0.0119575
R59945 ASIG5V.n7603 ASIG5V.n7593 0.0119575
R59946 ASIG5V.n7582 ASIG5V.n7578 0.0119575
R59947 ASIG5V.n7585 ASIG5V.n7584 0.0119575
R59948 ASIG5V.n7586 ASIG5V.n7581 0.0119575
R59949 ASIG5V.n7590 ASIG5V.n7583 0.0119575
R59950 ASIG5V.n7273 ASIG5V.n7271 0.0119575
R59951 ASIG5V.n8153 ASIG5V.n7275 0.0119575
R59952 ASIG5V.n7276 ASIG5V.n7270 0.0119575
R59953 ASIG5V.n8155 ASIG5V.n7267 0.0119575
R59954 ASIG5V.n8158 ASIG5V.n7262 0.0119575
R59955 ASIG5V.n8159 ASIG5V.n7261 0.0119575
R59956 ASIG5V.n7263 ASIG5V.n7259 0.0119575
R59957 ASIG5V.n8161 ASIG5V.n7256 0.0119575
R59958 ASIG5V.n8164 ASIG5V.n7251 0.0119575
R59959 ASIG5V.n8165 ASIG5V.n7250 0.0119575
R59960 ASIG5V.n7252 ASIG5V.n7248 0.0119575
R59961 ASIG5V.n8167 ASIG5V.n7245 0.0119575
R59962 ASIG5V.n7592 ASIG5V.n7578 0.0119575
R59963 ASIG5V.n7584 ASIG5V.n7582 0.0119575
R59964 ASIG5V.n7586 ASIG5V.n7585 0.0119575
R59965 ASIG5V.n7583 ASIG5V.n7581 0.0119575
R59966 ASIG5V.n7600 ASIG5V.n7566 0.0119575
R59967 ASIG5V.n7594 ASIG5V.n7577 0.0119575
R59968 ASIG5V.n7596 ASIG5V.n7595 0.0119575
R59969 ASIG5V.n7603 ASIG5V.n7602 0.0119575
R59970 ASIG5V.n7645 ASIG5V.n7568 0.0119575
R59971 ASIG5V.n7569 ASIG5V.n7564 0.0119575
R59972 ASIG5V.n7648 ASIG5V.n7647 0.0119575
R59973 ASIG5V.n7565 ASIG5V.n7562 0.0119575
R59974 ASIG5V.n7492 ASIG5V.n7489 0.0119575
R59975 ASIG5V.n8076 ASIG5V.n7488 0.0119575
R59976 ASIG5V.n8075 ASIG5V.n7491 0.0119575
R59977 ASIG5V.n8079 ASIG5V.n8078 0.0119575
R59978 ASIG5V.n3104 ASIG5V.n3101 0.0119575
R59979 ASIG5V.n9860 ASIG5V.n3100 0.0119575
R59980 ASIG5V.n9859 ASIG5V.n3103 0.0119575
R59981 ASIG5V.n9863 ASIG5V.n9862 0.0119575
R59982 ASIG5V.n7274 ASIG5V.n7273 0.0119575
R59983 ASIG5V.n8143 ASIG5V.n7285 0.0119575
R59984 ASIG5V.n7368 ASIG5V.n7303 0.0119575
R59985 ASIG5V.n7448 ASIG5V.n7327 0.0119575
R59986 ASIG5V.n7275 ASIG5V.n7271 0.0119575
R59987 ASIG5V.n7286 ASIG5V.n7281 0.0119575
R59988 ASIG5V.n7371 ASIG5V.n7370 0.0119575
R59989 ASIG5V.n7441 ASIG5V.n7330 0.0119575
R59990 ASIG5V.n7442 ASIG5V.n7329 0.0119575
R59991 ASIG5V.n7373 ASIG5V.n7372 0.0119575
R59992 ASIG5V.n8146 ASIG5V.n8145 0.0119575
R59993 ASIG5V.n8153 ASIG5V.n7276 0.0119575
R59994 ASIG5V.n7440 ASIG5V.n7439 0.0119575
R59995 ASIG5V.n7367 ASIG5V.n7364 0.0119575
R59996 ASIG5V.n7282 ASIG5V.n7279 0.0119575
R59997 ASIG5V.n7270 ASIG5V.n7267 0.0119575
R59998 ASIG5V.n3111 ASIG5V.n3107 0.0119575
R59999 ASIG5V.n9851 ASIG5V.n9850 0.0119575
R60000 ASIG5V.n9853 ASIG5V.n3110 0.0119575
R60001 ASIG5V.n9854 ASIG5V.n3109 0.0119575
R60002 ASIG5V.n7499 ASIG5V.n7495 0.0119575
R60003 ASIG5V.n8067 ASIG5V.n8066 0.0119575
R60004 ASIG5V.n8069 ASIG5V.n7498 0.0119575
R60005 ASIG5V.n8070 ASIG5V.n7497 0.0119575
R60006 ASIG5V.n7657 ASIG5V.n7561 0.0119575
R60007 ASIG5V.n7660 ASIG5V.n7658 0.0119575
R60008 ASIG5V.n7659 ASIG5V.n7560 0.0119575
R60009 ASIG5V.n7664 ASIG5V.n7558 0.0119575
R60010 ASIG5V.n7668 ASIG5V.n7556 0.0119575
R60011 ASIG5V.n7671 ASIG5V.n7669 0.0119575
R60012 ASIG5V.n7670 ASIG5V.n7555 0.0119575
R60013 ASIG5V.n7675 ASIG5V.n7553 0.0119575
R60014 ASIG5V.n7679 ASIG5V.n7551 0.0119575
R60015 ASIG5V.n7682 ASIG5V.n7680 0.0119575
R60016 ASIG5V.n7681 ASIG5V.n7550 0.0119575
R60017 ASIG5V.n7686 ASIG5V.n7548 0.0119575
R60018 ASIG5V.n7690 ASIG5V.n7689 0.0119575
R60019 ASIG5V.n7693 ASIG5V.n7691 0.0119575
R60020 ASIG5V.n7692 ASIG5V.n7547 0.0119575
R60021 ASIG5V.n7697 ASIG5V.n7545 0.0119575
R60022 ASIG5V.n7700 ASIG5V.n7699 0.0119575
R60023 ASIG5V.n7701 ASIG5V.n7544 0.0119575
R60024 ASIG5V.n7543 ASIG5V.n7541 0.0119575
R60025 ASIG5V.n7704 ASIG5V.n7539 0.0119575
R60026 ASIG5V.n7706 ASIG5V.n7538 0.0119575
R60027 ASIG5V.n7708 ASIG5V.n7535 0.0119575
R60028 ASIG5V.n7707 ASIG5V.n7533 0.0119575
R60029 ASIG5V.n7712 ASIG5V.n7536 0.0119575
R60030 ASIG5V.n7689 ASIG5V.n7688 0.0119575
R60031 ASIG5V.n7691 ASIG5V.n7690 0.0119575
R60032 ASIG5V.n7693 ASIG5V.n7692 0.0119575
R60033 ASIG5V.n7547 ASIG5V.n7545 0.0119575
R60034 ASIG5V.n7677 ASIG5V.n7551 0.0119575
R60035 ASIG5V.n7680 ASIG5V.n7679 0.0119575
R60036 ASIG5V.n7682 ASIG5V.n7681 0.0119575
R60037 ASIG5V.n7550 ASIG5V.n7548 0.0119575
R60038 ASIG5V.n7666 ASIG5V.n7556 0.0119575
R60039 ASIG5V.n7669 ASIG5V.n7668 0.0119575
R60040 ASIG5V.n7671 ASIG5V.n7670 0.0119575
R60041 ASIG5V.n7555 ASIG5V.n7553 0.0119575
R60042 ASIG5V.n7655 ASIG5V.n7561 0.0119575
R60043 ASIG5V.n7658 ASIG5V.n7657 0.0119575
R60044 ASIG5V.n7660 ASIG5V.n7659 0.0119575
R60045 ASIG5V.n7560 ASIG5V.n7558 0.0119575
R60046 ASIG5V.n7499 ASIG5V.n7496 0.0119575
R60047 ASIG5V.n8067 ASIG5V.n7495 0.0119575
R60048 ASIG5V.n8066 ASIG5V.n7498 0.0119575
R60049 ASIG5V.n8070 ASIG5V.n8069 0.0119575
R60050 ASIG5V.n3111 ASIG5V.n3108 0.0119575
R60051 ASIG5V.n9851 ASIG5V.n3107 0.0119575
R60052 ASIG5V.n9850 ASIG5V.n3110 0.0119575
R60053 ASIG5V.n9854 ASIG5V.n9853 0.0119575
R60054 ASIG5V.n7699 ASIG5V.n7698 0.0119575
R60055 ASIG5V.n8156 ASIG5V.n7262 0.0119575
R60056 ASIG5V.n7352 ASIG5V.n7283 0.0119575
R60057 ASIG5V.n7378 ASIG5V.n7362 0.0119575
R60058 ASIG5V.n7437 ASIG5V.n7331 0.0119575
R60059 ASIG5V.n7701 ASIG5V.n7700 0.0119575
R60060 ASIG5V.n8159 ASIG5V.n8158 0.0119575
R60061 ASIG5V.n7389 ASIG5V.n7388 0.0119575
R60062 ASIG5V.n7363 ASIG5V.n7359 0.0119575
R60063 ASIG5V.n7430 ASIG5V.n7334 0.0119575
R60064 ASIG5V.n7431 ASIG5V.n7333 0.0119575
R60065 ASIG5V.n7381 ASIG5V.n7380 0.0119575
R60066 ASIG5V.n7353 ASIG5V.n7351 0.0119575
R60067 ASIG5V.n7263 ASIG5V.n7261 0.0119575
R60068 ASIG5V.n7544 ASIG5V.n7543 0.0119575
R60069 ASIG5V.n7429 ASIG5V.n7428 0.0119575
R60070 ASIG5V.n7360 ASIG5V.n7357 0.0119575
R60071 ASIG5V.n7349 ASIG5V.n7347 0.0119575
R60072 ASIG5V.n7259 ASIG5V.n7256 0.0119575
R60073 ASIG5V.n7541 ASIG5V.n7539 0.0119575
R60074 ASIG5V.n9827 ASIG5V.n3121 0.0119575
R60075 ASIG5V.n9833 ASIG5V.n9832 0.0119575
R60076 ASIG5V.n9835 ASIG5V.n9826 0.0119575
R60077 ASIG5V.n9836 ASIG5V.n9825 0.0119575
R60078 ASIG5V.n3126 ASIG5V.n3123 0.0119575
R60079 ASIG5V.n9819 ASIG5V.n9818 0.0119575
R60080 ASIG5V.n9821 ASIG5V.n9814 0.0119575
R60081 ASIG5V.n9822 ASIG5V.n9813 0.0119575
R60082 ASIG5V.n3131 ASIG5V.n3128 0.0119575
R60083 ASIG5V.n9807 ASIG5V.n9806 0.0119575
R60084 ASIG5V.n9809 ASIG5V.n9802 0.0119575
R60085 ASIG5V.n9810 ASIG5V.n9801 0.0119575
R60086 ASIG5V.n3136 ASIG5V.n3133 0.0119575
R60087 ASIG5V.n9795 ASIG5V.n9794 0.0119575
R60088 ASIG5V.n9797 ASIG5V.n9790 0.0119575
R60089 ASIG5V.n9798 ASIG5V.n9789 0.0119575
R60090 ASIG5V.n3141 ASIG5V.n3138 0.0119575
R60091 ASIG5V.n9783 ASIG5V.n9782 0.0119575
R60092 ASIG5V.n9785 ASIG5V.n9778 0.0119575
R60093 ASIG5V.n9786 ASIG5V.n9777 0.0119575
R60094 ASIG5V.n3146 ASIG5V.n3143 0.0119575
R60095 ASIG5V.n9771 ASIG5V.n9770 0.0119575
R60096 ASIG5V.n9773 ASIG5V.n9766 0.0119575
R60097 ASIG5V.n9774 ASIG5V.n9765 0.0119575
R60098 ASIG5V.n3152 ASIG5V.n3148 0.0119575
R60099 ASIG5V.n9757 ASIG5V.n9756 0.0119575
R60100 ASIG5V.n9758 ASIG5V.n3151 0.0119575
R60101 ASIG5V.n9762 ASIG5V.n3154 0.0119575
R60102 ASIG5V.n3158 ASIG5V.n3156 0.0119575
R60103 ASIG5V.n9749 ASIG5V.n3161 0.0119575
R60104 ASIG5V.n3160 ASIG5V.n3157 0.0119575
R60105 ASIG5V.n9752 ASIG5V.n3162 0.0119575
R60106 ASIG5V.n9764 ASIG5V.n3148 0.0119575
R60107 ASIG5V.n9756 ASIG5V.n3152 0.0119575
R60108 ASIG5V.n9758 ASIG5V.n9757 0.0119575
R60109 ASIG5V.n3154 ASIG5V.n3151 0.0119575
R60110 ASIG5V.n9776 ASIG5V.n3143 0.0119575
R60111 ASIG5V.n9771 ASIG5V.n3146 0.0119575
R60112 ASIG5V.n9770 ASIG5V.n9766 0.0119575
R60113 ASIG5V.n9774 ASIG5V.n9773 0.0119575
R60114 ASIG5V.n9788 ASIG5V.n3138 0.0119575
R60115 ASIG5V.n9783 ASIG5V.n3141 0.0119575
R60116 ASIG5V.n9782 ASIG5V.n9778 0.0119575
R60117 ASIG5V.n9786 ASIG5V.n9785 0.0119575
R60118 ASIG5V.n9800 ASIG5V.n3133 0.0119575
R60119 ASIG5V.n9795 ASIG5V.n3136 0.0119575
R60120 ASIG5V.n9794 ASIG5V.n9790 0.0119575
R60121 ASIG5V.n9798 ASIG5V.n9797 0.0119575
R60122 ASIG5V.n9812 ASIG5V.n3128 0.0119575
R60123 ASIG5V.n9807 ASIG5V.n3131 0.0119575
R60124 ASIG5V.n9806 ASIG5V.n9802 0.0119575
R60125 ASIG5V.n9810 ASIG5V.n9809 0.0119575
R60126 ASIG5V.n9824 ASIG5V.n3123 0.0119575
R60127 ASIG5V.n9819 ASIG5V.n3126 0.0119575
R60128 ASIG5V.n9818 ASIG5V.n9814 0.0119575
R60129 ASIG5V.n9822 ASIG5V.n9821 0.0119575
R60130 ASIG5V.n9827 ASIG5V.n3122 0.0119575
R60131 ASIG5V.n9833 ASIG5V.n3121 0.0119575
R60132 ASIG5V.n9832 ASIG5V.n9826 0.0119575
R60133 ASIG5V.n9836 ASIG5V.n9835 0.0119575
R60134 ASIG5V.n9754 ASIG5V.n3156 0.0119575
R60135 ASIG5V.n7706 ASIG5V.n7705 0.0119575
R60136 ASIG5V.n8162 ASIG5V.n7251 0.0119575
R60137 ASIG5V.n7394 ASIG5V.n7392 0.0119575
R60138 ASIG5V.n7343 ASIG5V.n7338 0.0119575
R60139 ASIG5V.n7426 ASIG5V.n7335 0.0119575
R60140 ASIG5V.n9749 ASIG5V.n3158 0.0119575
R60141 ASIG5V.n7538 ASIG5V.n7535 0.0119575
R60142 ASIG5V.n8165 ASIG5V.n8164 0.0119575
R60143 ASIG5V.n7400 ASIG5V.n7346 0.0119575
R60144 ASIG5V.n7409 ASIG5V.n7337 0.0119575
R60145 ASIG5V.n7419 ASIG5V.n7416 0.0119575
R60146 ASIG5V.n7420 ASIG5V.n7415 0.0119575
R60147 ASIG5V.n7408 ASIG5V.n7342 0.0119575
R60148 ASIG5V.n7399 ASIG5V.n7393 0.0119575
R60149 ASIG5V.n7252 ASIG5V.n7250 0.0119575
R60150 ASIG5V.n7708 ASIG5V.n7707 0.0119575
R60151 ASIG5V.n3161 ASIG5V.n3160 0.0119575
R60152 ASIG5V.n7418 ASIG5V.n7417 0.0119575
R60153 ASIG5V.n7412 ASIG5V.n7411 0.0119575
R60154 ASIG5V.n7403 ASIG5V.n7402 0.0119575
R60155 ASIG5V.n7248 ASIG5V.n7245 0.0119575
R60156 ASIG5V.n7536 ASIG5V.n7533 0.0119575
R60157 ASIG5V.n3162 ASIG5V.n3157 0.0119575
R60158 ASIG5V.n9903 ASIG5V.n9896 0.0119575
R60159 ASIG5V.n9904 ASIG5V.n9895 0.0119575
R60160 ASIG5V.n9897 ASIG5V.n9893 0.0119575
R60161 ASIG5V.n9906 ASIG5V.n3076 0.0119575
R60162 ASIG5V.n9909 ASIG5V.n3071 0.0119575
R60163 ASIG5V.n9910 ASIG5V.n3070 0.0119575
R60164 ASIG5V.n3072 ASIG5V.n3068 0.0119575
R60165 ASIG5V.n9912 ASIG5V.n3065 0.0119575
R60166 ASIG5V.n9915 ASIG5V.n3060 0.0119575
R60167 ASIG5V.n9916 ASIG5V.n3059 0.0119575
R60168 ASIG5V.n3061 ASIG5V.n3057 0.0119575
R60169 ASIG5V.n9918 ASIG5V.n3054 0.0119575
R60170 ASIG5V.n9921 ASIG5V.n3049 0.0119575
R60171 ASIG5V.n9922 ASIG5V.n3048 0.0119575
R60172 ASIG5V.n3050 ASIG5V.n3046 0.0119575
R60173 ASIG5V.n9924 ASIG5V.n3043 0.0119575
R60174 ASIG5V.n9927 ASIG5V.n3038 0.0119575
R60175 ASIG5V.n9928 ASIG5V.n3037 0.0119575
R60176 ASIG5V.n3039 ASIG5V.n3035 0.0119575
R60177 ASIG5V.n9930 ASIG5V.n3032 0.0119575
R60178 ASIG5V.n9933 ASIG5V.n3027 0.0119575
R60179 ASIG5V.n9934 ASIG5V.n3026 0.0119575
R60180 ASIG5V.n3028 ASIG5V.n3024 0.0119575
R60181 ASIG5V.n9936 ASIG5V.n3021 0.0119575
R60182 ASIG5V.n9939 ASIG5V.n3016 0.0119575
R60183 ASIG5V.n9940 ASIG5V.n3015 0.0119575
R60184 ASIG5V.n3017 ASIG5V.n3013 0.0119575
R60185 ASIG5V.n9942 ASIG5V.n3010 0.0119575
R60186 ASIG5V.n3008 ASIG5V.n3007 0.0119575
R60187 ASIG5V.n9948 ASIG5V.n9946 0.0119575
R60188 ASIG5V.n9947 ASIG5V.n3006 0.0119575
R60189 ASIG5V.n9952 ASIG5V.n3003 0.0119575
R60190 ASIG5V.n9943 ASIG5V.n3007 0.0119575
R60191 ASIG5V.n9946 ASIG5V.n3008 0.0119575
R60192 ASIG5V.n9948 ASIG5V.n9947 0.0119575
R60193 ASIG5V.n3006 ASIG5V.n3003 0.0119575
R60194 ASIG5V.n9937 ASIG5V.n3016 0.0119575
R60195 ASIG5V.n9940 ASIG5V.n9939 0.0119575
R60196 ASIG5V.n3017 ASIG5V.n3015 0.0119575
R60197 ASIG5V.n3013 ASIG5V.n3010 0.0119575
R60198 ASIG5V.n9931 ASIG5V.n3027 0.0119575
R60199 ASIG5V.n9934 ASIG5V.n9933 0.0119575
R60200 ASIG5V.n3028 ASIG5V.n3026 0.0119575
R60201 ASIG5V.n3024 ASIG5V.n3021 0.0119575
R60202 ASIG5V.n9925 ASIG5V.n3038 0.0119575
R60203 ASIG5V.n9928 ASIG5V.n9927 0.0119575
R60204 ASIG5V.n3039 ASIG5V.n3037 0.0119575
R60205 ASIG5V.n3035 ASIG5V.n3032 0.0119575
R60206 ASIG5V.n9919 ASIG5V.n3049 0.0119575
R60207 ASIG5V.n9922 ASIG5V.n9921 0.0119575
R60208 ASIG5V.n3050 ASIG5V.n3048 0.0119575
R60209 ASIG5V.n3046 ASIG5V.n3043 0.0119575
R60210 ASIG5V.n9913 ASIG5V.n3060 0.0119575
R60211 ASIG5V.n9916 ASIG5V.n9915 0.0119575
R60212 ASIG5V.n3061 ASIG5V.n3059 0.0119575
R60213 ASIG5V.n3057 ASIG5V.n3054 0.0119575
R60214 ASIG5V.n9907 ASIG5V.n3071 0.0119575
R60215 ASIG5V.n9910 ASIG5V.n9909 0.0119575
R60216 ASIG5V.n3072 ASIG5V.n3070 0.0119575
R60217 ASIG5V.n3068 ASIG5V.n3065 0.0119575
R60218 ASIG5V.n9901 ASIG5V.n9896 0.0119575
R60219 ASIG5V.n9904 ASIG5V.n9903 0.0119575
R60220 ASIG5V.n9897 ASIG5V.n9895 0.0119575
R60221 ASIG5V.n9893 ASIG5V.n3076 0.0119575
R60222 ASIG5V.n3118 ASIG5V.n3114 0.0119575
R60223 ASIG5V.n9842 ASIG5V.n9841 0.0119575
R60224 ASIG5V.n9844 ASIG5V.n3117 0.0119575
R60225 ASIG5V.n9845 ASIG5V.n3116 0.0119575
R60226 ASIG5V.n8058 ASIG5V.n7502 0.0119575
R60227 ASIG5V.n8053 ASIG5V.n8052 0.0119575
R60228 ASIG5V.n8060 ASIG5V.n8054 0.0119575
R60229 ASIG5V.n8061 ASIG5V.n8051 0.0119575
R60230 ASIG5V.n7507 ASIG5V.n7504 0.0119575
R60231 ASIG5V.n8042 ASIG5V.n8041 0.0119575
R60232 ASIG5V.n8047 ASIG5V.n8043 0.0119575
R60233 ASIG5V.n8048 ASIG5V.n8040 0.0119575
R60234 ASIG5V.n7512 ASIG5V.n7509 0.0119575
R60235 ASIG5V.n8031 ASIG5V.n8030 0.0119575
R60236 ASIG5V.n8036 ASIG5V.n8032 0.0119575
R60237 ASIG5V.n8037 ASIG5V.n8029 0.0119575
R60238 ASIG5V.n7517 ASIG5V.n7514 0.0119575
R60239 ASIG5V.n8020 ASIG5V.n8019 0.0119575
R60240 ASIG5V.n8025 ASIG5V.n8021 0.0119575
R60241 ASIG5V.n8026 ASIG5V.n8018 0.0119575
R60242 ASIG5V.n7522 ASIG5V.n7519 0.0119575
R60243 ASIG5V.n8009 ASIG5V.n8008 0.0119575
R60244 ASIG5V.n8014 ASIG5V.n8010 0.0119575
R60245 ASIG5V.n8015 ASIG5V.n8007 0.0119575
R60246 ASIG5V.n7527 ASIG5V.n7524 0.0119575
R60247 ASIG5V.n7998 ASIG5V.n7997 0.0119575
R60248 ASIG5V.n8003 ASIG5V.n7999 0.0119575
R60249 ASIG5V.n8004 ASIG5V.n7996 0.0119575
R60250 ASIG5V.n7532 ASIG5V.n7529 0.0119575
R60251 ASIG5V.n7990 ASIG5V.n7989 0.0119575
R60252 ASIG5V.n7992 ASIG5V.n7984 0.0119575
R60253 ASIG5V.n7993 ASIG5V.n7983 0.0119575
R60254 ASIG5V.n7995 ASIG5V.n7529 0.0119575
R60255 ASIG5V.n7990 ASIG5V.n7532 0.0119575
R60256 ASIG5V.n7989 ASIG5V.n7984 0.0119575
R60257 ASIG5V.n7993 ASIG5V.n7992 0.0119575
R60258 ASIG5V.n8006 ASIG5V.n7524 0.0119575
R60259 ASIG5V.n7997 ASIG5V.n7527 0.0119575
R60260 ASIG5V.n7999 ASIG5V.n7998 0.0119575
R60261 ASIG5V.n8004 ASIG5V.n8003 0.0119575
R60262 ASIG5V.n8017 ASIG5V.n7519 0.0119575
R60263 ASIG5V.n8008 ASIG5V.n7522 0.0119575
R60264 ASIG5V.n8010 ASIG5V.n8009 0.0119575
R60265 ASIG5V.n8015 ASIG5V.n8014 0.0119575
R60266 ASIG5V.n8028 ASIG5V.n7514 0.0119575
R60267 ASIG5V.n8019 ASIG5V.n7517 0.0119575
R60268 ASIG5V.n8021 ASIG5V.n8020 0.0119575
R60269 ASIG5V.n8026 ASIG5V.n8025 0.0119575
R60270 ASIG5V.n8039 ASIG5V.n7509 0.0119575
R60271 ASIG5V.n8030 ASIG5V.n7512 0.0119575
R60272 ASIG5V.n8032 ASIG5V.n8031 0.0119575
R60273 ASIG5V.n8037 ASIG5V.n8036 0.0119575
R60274 ASIG5V.n8050 ASIG5V.n7504 0.0119575
R60275 ASIG5V.n8041 ASIG5V.n7507 0.0119575
R60276 ASIG5V.n8043 ASIG5V.n8042 0.0119575
R60277 ASIG5V.n8048 ASIG5V.n8047 0.0119575
R60278 ASIG5V.n8058 ASIG5V.n7503 0.0119575
R60279 ASIG5V.n8052 ASIG5V.n7502 0.0119575
R60280 ASIG5V.n8054 ASIG5V.n8053 0.0119575
R60281 ASIG5V.n8061 ASIG5V.n8060 0.0119575
R60282 ASIG5V.n3118 ASIG5V.n3115 0.0119575
R60283 ASIG5V.n9842 ASIG5V.n3114 0.0119575
R60284 ASIG5V.n9841 ASIG5V.n3117 0.0119575
R60285 ASIG5V.n9845 ASIG5V.n9844 0.0119575
R60286 ASIG5V.n4584 ASIG5V.n4583 0.0118684
R60287 ASIG5V.n7981 ASIG5V.n5908 0.0118684
R60288 ASIG5V.n512 ASIG5V.n9 0.0117009
R60289 ASIG5V.n10363 ASIG5V.n10069 0.0117009
R60290 ASIG5V.n511 ASIG5V.n8 0.0117009
R60291 ASIG5V.n11180 ASIG5V.n10364 0.0117009
R60292 ASIG5V.n8584 ASIG5V.n8320 0.0116141
R60293 ASIG5V.n9959 ASIG5V.n9958 0.0116141
R60294 ASIG5V.n8585 ASIG5V.n8321 0.0116141
R60295 ASIG5V.n11502 ASIG5V.n9955 0.0116141
R60296 ASIG5V.n4564 ASIG5V.n4560 0.011525
R60297 ASIG5V.n8925 ASIG5V.n6533 0.0113271
R60298 ASIG5V.n8901 ASIG5V.n8900 0.0113271
R60299 ASIG5V.n9736 ASIG5V.n3172 0.0113079
R60300 ASIG5V.n9737 ASIG5V.n3174 0.0113079
R60301 ASIG5V.n12332 ASIG5V.n165 0.0111309
R60302 ASIG5V.n2220 ASIG5V.n2214 0.0111309
R60303 ASIG5V.n12331 ASIG5V.n167 0.0111309
R60304 ASIG5V.n2219 ASIG5V.n2216 0.0111309
R60305 ASIG5V.n6886 ASIG5V.n6885 0.011075
R60306 ASIG5V.n12017 ASIG5V.n1316 0.0107857
R60307 ASIG5V.n12015 ASIG5V.n1322 0.0107857
R60308 ASIG5V.n3672 ASIG5V.n3619 0.0106477
R60309 ASIG5V.n7979 ASIG5V.n5569 0.0106477
R60310 ASIG5V.n4582 ASIG5V.n4581 0.0106477
R60311 ASIG5V.n7980 ASIG5V.n5571 0.0106477
R60312 ASIG5V.n12003 ASIG5V.n1669 0.010625
R60313 ASIG5V.n2204 ASIG5V.n2203 0.010625
R60314 ASIG5V.n3615 ASIG5V.n3280 0.0105588
R60315 ASIG5V.n3406 ASIG5V.n3274 0.0105588
R60316 ASIG5V.n3614 ASIG5V.n3279 0.0105588
R60317 ASIG5V.n3405 ASIG5V.n3275 0.0105588
R60318 ASIG5V.n4815 ASIG5V.n4814 0.0105588
R60319 ASIG5V.n3222 ASIG5V.n3176 0.0105588
R60320 ASIG5V.n4810 ASIG5V.n3220 0.0105588
R60321 ASIG5V.n5063 ASIG5V.n3177 0.0105588
R60322 ASIG5V.n9486 ASIG5V.n3166 0.0105588
R60323 ASIG5V.n9442 ASIG5V.n3174 0.0105588
R60324 ASIG5V.n5116 ASIG5V.n3168 0.0105588
R60325 ASIG5V.n9733 ASIG5V.n3172 0.0105588
R60326 ASIG5V.n5214 ASIG5V.n5121 0.0105588
R60327 ASIG5V.n5461 ASIG5V.n5168 0.0105588
R60328 ASIG5V.n5165 ASIG5V.n5122 0.0105588
R60329 ASIG5V.n9431 ASIG5V.n5167 0.0105588
R60330 ASIG5V.n7716 ASIG5V.n5509 0.0105588
R60331 ASIG5V.n9414 ASIG5V.n9413 0.0105588
R60332 ASIG5V.n9417 ASIG5V.n5508 0.0105588
R60333 ASIG5V.n9415 ASIG5V.n5554 0.0105588
R60334 ASIG5V.n5906 ASIG5V.n5571 0.0105588
R60335 ASIG5V.n5697 ASIG5V.n5564 0.0105588
R60336 ASIG5V.n5905 ASIG5V.n5569 0.0105588
R60337 ASIG5V.n5696 ASIG5V.n5566 0.0105588
R60338 ASIG5V.n5956 ASIG5V.n5910 0.0105588
R60339 ASIG5V.n9391 ASIG5V.n9390 0.0105588
R60340 ASIG5V.n9394 ASIG5V.n5911 0.0105588
R60341 ASIG5V.n9392 ASIG5V.n6000 0.0105588
R60342 ASIG5V.n6428 ASIG5V.n6309 0.0105588
R60343 ASIG5V.n9377 ASIG5V.n6260 0.0105588
R60344 ASIG5V.n9380 ASIG5V.n6308 0.0105588
R60345 ASIG5V.n9378 ASIG5V.n6262 0.0105588
R60346 ASIG5V.n8928 ASIG5V.n8927 0.0105588
R60347 ASIG5V.n6489 ASIG5V.n6436 0.0105588
R60348 ASIG5V.n6538 ASIG5V.n6487 0.0105588
R60349 ASIG5V.n9175 ASIG5V.n6434 0.0105588
R60350 ASIG5V.n6589 ASIG5V.n6541 0.0105588
R60351 ASIG5V.n8914 ASIG5V.n8913 0.0105588
R60352 ASIG5V.n8917 ASIG5V.n6543 0.0105588
R60353 ASIG5V.n8915 ASIG5V.n6633 0.0105588
R60354 ASIG5V.n7230 ASIG5V.n6895 0.0105588
R60355 ASIG5V.n7021 ASIG5V.n6888 0.0105588
R60356 ASIG5V.n7229 ASIG5V.n6893 0.0105588
R60357 ASIG5V.n7020 ASIG5V.n6890 0.0105588
R60358 ASIG5V.n8324 ASIG5V.n8216 0.0105588
R60359 ASIG5V.n8890 ASIG5V.n8889 0.0105588
R60360 ASIG5V.n8893 ASIG5V.n8215 0.0105588
R60361 ASIG5V.n8891 ASIG5V.n8260 0.0105588
R60362 ASIG5V.n8878 ASIG5V.n8321 0.0105588
R60363 ASIG5V.n8633 ASIG5V.n4 0.0105588
R60364 ASIG5V.n8879 ASIG5V.n8320 0.0105588
R60365 ASIG5V.n8632 ASIG5V.n2 0.0105588
R60366 ASIG5V.n163 ASIG5V.n55 0.0105588
R60367 ASIG5V.n12523 ASIG5V.n8 0.0105588
R60368 ASIG5V.n12526 ASIG5V.n54 0.0105588
R60369 ASIG5V.n12524 ASIG5V.n9 0.0105588
R60370 ASIG5V.n260 ASIG5V.n167 0.0105588
R60371 ASIG5V.n517 ASIG5V.n218 0.0105588
R60372 ASIG5V.n215 ASIG5V.n165 0.0105588
R60373 ASIG5V.n12322 ASIG5V.n217 0.0105588
R60374 ASIG5V.n614 ASIG5V.n523 0.0105588
R60375 ASIG5V.n862 ASIG5V.n573 0.0105588
R60376 ASIG5V.n570 ASIG5V.n522 0.0105588
R60377 ASIG5V.n12300 ASIG5V.n572 0.0105588
R60378 ASIG5V.n966 ASIG5V.n871 0.0105588
R60379 ASIG5V.n1215 ASIG5V.n881 0.0105588
R60380 ASIG5V.n967 ASIG5V.n873 0.0105588
R60381 ASIG5V.n1214 ASIG5V.n879 0.0105588
R60382 ASIG5V.n12020 ASIG5V.n12019 0.0105588
R60383 ASIG5V.n1270 ASIG5V.n1222 0.0105588
R60384 ASIG5V.n1320 ASIG5V.n1268 0.0105588
R60385 ASIG5V.n12267 ASIG5V.n1224 0.0105588
R60386 ASIG5V.n1372 ASIG5V.n1323 0.0105588
R60387 ASIG5V.n12006 ASIG5V.n12005 0.0105588
R60388 ASIG5V.n12009 ASIG5V.n1325 0.0105588
R60389 ASIG5V.n12007 ASIG5V.n1416 0.0105588
R60390 ASIG5V.n1836 ASIG5V.n1720 0.0105588
R60391 ASIG5V.n11992 ASIG5V.n1671 0.0105588
R60392 ASIG5V.n11995 ASIG5V.n1719 0.0105588
R60393 ASIG5V.n11993 ASIG5V.n1673 0.0105588
R60394 ASIG5V.n1948 ASIG5V.n1844 0.0105588
R60395 ASIG5V.n1907 ASIG5V.n1857 0.0105588
R60396 ASIG5V.n1906 ASIG5V.n1846 0.0105588
R60397 ASIG5V.n2197 ASIG5V.n1863 0.0105588
R60398 ASIG5V.n2305 ASIG5V.n2219 0.0105588
R60399 ASIG5V.n2264 ASIG5V.n2208 0.0105588
R60400 ASIG5V.n2263 ASIG5V.n2220 0.0105588
R60401 ASIG5V.n2554 ASIG5V.n2210 0.0105588
R60402 ASIG5V.n2657 ASIG5V.n2565 0.0105588
R60403 ASIG5V.n2903 ASIG5V.n2614 0.0105588
R60404 ASIG5V.n2611 ASIG5V.n2567 0.0105588
R60405 ASIG5V.n11770 ASIG5V.n2613 0.0105588
R60406 ASIG5V.n11503 ASIG5V.n11502 0.0105588
R60407 ASIG5V.n2957 ASIG5V.n2908 0.0105588
R60408 ASIG5V.n9959 ASIG5V.n2955 0.0105588
R60409 ASIG5V.n11750 ASIG5V.n2905 0.0105588
R60410 ASIG5V.n11237 ASIG5V.n9962 0.0105588
R60411 ASIG5V.n11193 ASIG5V.n9968 0.0105588
R60412 ASIG5V.n10015 ASIG5V.n9964 0.0105588
R60413 ASIG5V.n11484 ASIG5V.n9967 0.0105588
R60414 ASIG5V.n10067 ASIG5V.n10024 0.0105588
R60415 ASIG5V.n11182 ASIG5V.n10069 0.0105588
R60416 ASIG5V.n4581 ASIG5V.n3673 0.0105588
R60417 ASIG5V.n4770 ASIG5V.n3626 0.0105588
R60418 ASIG5V.n4773 ASIG5V.n3672 0.0105588
R60419 ASIG5V.n4771 ASIG5V.n3628 0.0105588
R60420 ASIG5V.n10480 ASIG5V.n10415 0.0105588
R60421 ASIG5V.n11171 ASIG5V.n10372 0.0105588
R60422 ASIG5V.n3829 ASIG5V.n3779 0.0105588
R60423 ASIG5V.n4567 ASIG5V.n3831 0.0105588
R60424 ASIG5V.n4309 ASIG5V.n3782 0.0105588
R60425 ASIG5V.n4566 ASIG5V.n3835 0.0105588
R60426 ASIG5V.n10116 ASIG5V.n10023 0.0105588
R60427 ASIG5V.n11181 ASIG5V.n11180 0.0105588
R60428 ASIG5V.n10468 ASIG5V.n10463 0.0105588
R60429 ASIG5V.n11170 ASIG5V.n10370 0.0105588
R60430 ASIG5V ASIG5V.t4 0.0104057
R60431 ASIG5V ASIG5V.t1 0.0104057
R60432 ASIG5V ASIG5V.t0 0.0104057
R60433 ASIG5V ASIG5V.t6 0.0104057
R60434 ASIG5V.n9834 ASIG5V.n9831 0.0102808
R60435 ASIG5V.n9829 ASIG5V.n9828 0.0102808
R60436 ASIG5V.n9837 ASIG5V.n3120 0.0102808
R60437 ASIG5V.n9843 ASIG5V.n9840 0.0102808
R60438 ASIG5V.n9838 ASIG5V.n3119 0.0102808
R60439 ASIG5V.n9846 ASIG5V.n3113 0.0102808
R60440 ASIG5V.n9852 ASIG5V.n9849 0.0102808
R60441 ASIG5V.n9847 ASIG5V.n3112 0.0102808
R60442 ASIG5V.n9855 ASIG5V.n3106 0.0102808
R60443 ASIG5V.n9861 ASIG5V.n9858 0.0102808
R60444 ASIG5V.n9856 ASIG5V.n3105 0.0102808
R60445 ASIG5V.n9864 ASIG5V.n3099 0.0102808
R60446 ASIG5V.n9870 ASIG5V.n9867 0.0102808
R60447 ASIG5V.n9865 ASIG5V.n3098 0.0102808
R60448 ASIG5V.n9873 ASIG5V.n3092 0.0102808
R60449 ASIG5V.n9879 ASIG5V.n9876 0.0102808
R60450 ASIG5V.n9874 ASIG5V.n3091 0.0102808
R60451 ASIG5V.n9882 ASIG5V.n3085 0.0102808
R60452 ASIG5V.n9886 ASIG5V.n9885 0.0102808
R60453 ASIG5V.n9890 ASIG5V.n9889 0.0102808
R60454 ASIG5V.n9892 ASIG5V.n3078 0.0102808
R60455 ASIG5V.n9905 ASIG5V.n9894 0.0102808
R60456 ASIG5V.n9899 ASIG5V.n3077 0.0102808
R60457 ASIG5V.n9902 ASIG5V.n9900 0.0102808
R60458 ASIG5V.n9820 ASIG5V.n3124 0.0102808
R60459 ASIG5V.n9817 ASIG5V.n9816 0.0102808
R60460 ASIG5V.n9823 ASIG5V.n3125 0.0102808
R60461 ASIG5V.n8055 ASIG5V.n3127 0.0102808
R60462 ASIG5V.n8059 ASIG5V.n8057 0.0102808
R60463 ASIG5V.n8062 ASIG5V.n7501 0.0102808
R60464 ASIG5V.n8068 ASIG5V.n8065 0.0102808
R60465 ASIG5V.n8063 ASIG5V.n7500 0.0102808
R60466 ASIG5V.n8071 ASIG5V.n7494 0.0102808
R60467 ASIG5V.n8077 ASIG5V.n8074 0.0102808
R60468 ASIG5V.n8072 ASIG5V.n7493 0.0102808
R60469 ASIG5V.n8080 ASIG5V.n7487 0.0102808
R60470 ASIG5V.n8086 ASIG5V.n8083 0.0102808
R60471 ASIG5V.n8081 ASIG5V.n7486 0.0102808
R60472 ASIG5V.n8089 ASIG5V.n7480 0.0102808
R60473 ASIG5V.n8095 ASIG5V.n8092 0.0102808
R60474 ASIG5V.n8090 ASIG5V.n7479 0.0102808
R60475 ASIG5V.n8098 ASIG5V.n7473 0.0102808
R60476 ASIG5V.n8100 ASIG5V.n8099 0.0102808
R60477 ASIG5V.n8106 ASIG5V.n8105 0.0102808
R60478 ASIG5V.n8104 ASIG5V.n3067 0.0102808
R60479 ASIG5V.n9911 ASIG5V.n3069 0.0102808
R60480 ASIG5V.n3074 ASIG5V.n3066 0.0102808
R60481 ASIG5V.n9908 ASIG5V.n3075 0.0102808
R60482 ASIG5V.n8099 ASIG5V.n7469 0.0102808
R60483 ASIG5V.n8105 ASIG5V.n8104 0.0102808
R60484 ASIG5V.n8106 ASIG5V.n7469 0.0102808
R60485 ASIG5V.n9887 ASIG5V.n9886 0.0102808
R60486 ASIG5V.n9889 ASIG5V.n3078 0.0102808
R60487 ASIG5V.n9890 ASIG5V.n9887 0.0102808
R60488 ASIG5V.n9808 ASIG5V.n3129 0.0102808
R60489 ASIG5V.n9805 ASIG5V.n9804 0.0102808
R60490 ASIG5V.n9811 ASIG5V.n3130 0.0102808
R60491 ASIG5V.n7505 ASIG5V.n3132 0.0102808
R60492 ASIG5V.n8046 ASIG5V.n8045 0.0102808
R60493 ASIG5V.n8049 ASIG5V.n7506 0.0102808
R60494 ASIG5V.n7654 ASIG5V.n7508 0.0102808
R60495 ASIG5V.n7663 ASIG5V.n7662 0.0102808
R60496 ASIG5V.n7661 ASIG5V.n7656 0.0102808
R60497 ASIG5V.n7653 ASIG5V.n7563 0.0102808
R60498 ASIG5V.n7651 ASIG5V.n7650 0.0102808
R60499 ASIG5V.n7649 ASIG5V.n7646 0.0102808
R60500 ASIG5V.n7644 ASIG5V.n7571 0.0102808
R60501 ASIG5V.n7642 ASIG5V.n7641 0.0102808
R60502 ASIG5V.n7640 ASIG5V.n7637 0.0102808
R60503 ASIG5V.n7635 ASIG5V.n7634 0.0102808
R60504 ASIG5V.n7630 ASIG5V.n7625 0.0102808
R60505 ASIG5V.n7629 ASIG5V.n7464 0.0102808
R60506 ASIG5V.n8111 ASIG5V.n7463 0.0102808
R60507 ASIG5V.n8110 ASIG5V.n3056 0.0102808
R60508 ASIG5V.n9917 ASIG5V.n3058 0.0102808
R60509 ASIG5V.n3063 ASIG5V.n3055 0.0102808
R60510 ASIG5V.n9914 ASIG5V.n3064 0.0102808
R60511 ASIG5V.n8111 ASIG5V.n8110 0.0102808
R60512 ASIG5V.n7467 ASIG5V.n7463 0.0102808
R60513 ASIG5V.n7634 ASIG5V.n7623 0.0102808
R60514 ASIG5V.n7630 ASIG5V.n7629 0.0102808
R60515 ASIG5V.n7625 ASIG5V.n7623 0.0102808
R60516 ASIG5V.n8092 ASIG5V.n8091 0.0102808
R60517 ASIG5V.n7479 ASIG5V.n7473 0.0102808
R60518 ASIG5V.n8091 ASIG5V.n8090 0.0102808
R60519 ASIG5V.n9876 ASIG5V.n9875 0.0102808
R60520 ASIG5V.n3091 ASIG5V.n3085 0.0102808
R60521 ASIG5V.n9875 ASIG5V.n9874 0.0102808
R60522 ASIG5V.n9796 ASIG5V.n3134 0.0102808
R60523 ASIG5V.n9793 ASIG5V.n9792 0.0102808
R60524 ASIG5V.n9799 ASIG5V.n3135 0.0102808
R60525 ASIG5V.n7510 ASIG5V.n3137 0.0102808
R60526 ASIG5V.n8035 ASIG5V.n8034 0.0102808
R60527 ASIG5V.n8038 ASIG5V.n7511 0.0102808
R60528 ASIG5V.n7665 ASIG5V.n7513 0.0102808
R60529 ASIG5V.n7674 ASIG5V.n7673 0.0102808
R60530 ASIG5V.n7672 ASIG5V.n7667 0.0102808
R60531 ASIG5V.n7597 ASIG5V.n7557 0.0102808
R60532 ASIG5V.n7601 ASIG5V.n7599 0.0102808
R60533 ASIG5V.n7604 ASIG5V.n7576 0.0102808
R60534 ASIG5V.n7616 ASIG5V.n7615 0.0102808
R60535 ASIG5V.n7610 ASIG5V.n7608 0.0102808
R60536 ASIG5V.n7611 ASIG5V.n7310 0.0102808
R60537 ASIG5V.n7318 ASIG5V.n7309 0.0102808
R60538 ASIG5V.n8126 ASIG5V.n7319 0.0102808
R60539 ASIG5V.n8125 ASIG5V.n7321 0.0102808
R60540 ASIG5V.n8123 ASIG5V.n8122 0.0102808
R60541 ASIG5V.n8121 ASIG5V.n3045 0.0102808
R60542 ASIG5V.n9923 ASIG5V.n3047 0.0102808
R60543 ASIG5V.n3052 ASIG5V.n3044 0.0102808
R60544 ASIG5V.n9920 ASIG5V.n3053 0.0102808
R60545 ASIG5V.n7319 ASIG5V.n7318 0.0102808
R60546 ASIG5V.n7460 ASIG5V.n7321 0.0102808
R60547 ASIG5V.n8122 ASIG5V.n8121 0.0102808
R60548 ASIG5V.n8123 ASIG5V.n7460 0.0102808
R60549 ASIG5V.n7313 ASIG5V.n7309 0.0102808
R60550 ASIG5V.n7616 ASIG5V.n7575 0.0102808
R60551 ASIG5V.n7611 ASIG5V.n7610 0.0102808
R60552 ASIG5V.n7608 ASIG5V.n7575 0.0102808
R60553 ASIG5V.n7618 ASIG5V.n7571 0.0102808
R60554 ASIG5V.n7641 ASIG5V.n7640 0.0102808
R60555 ASIG5V.n7642 ASIG5V.n7618 0.0102808
R60556 ASIG5V.n8083 ASIG5V.n8082 0.0102808
R60557 ASIG5V.n7486 ASIG5V.n7480 0.0102808
R60558 ASIG5V.n8082 ASIG5V.n8081 0.0102808
R60559 ASIG5V.n9867 ASIG5V.n9866 0.0102808
R60560 ASIG5V.n3098 ASIG5V.n3092 0.0102808
R60561 ASIG5V.n9866 ASIG5V.n9865 0.0102808
R60562 ASIG5V.n9784 ASIG5V.n3139 0.0102808
R60563 ASIG5V.n9781 ASIG5V.n9780 0.0102808
R60564 ASIG5V.n9787 ASIG5V.n3140 0.0102808
R60565 ASIG5V.n7515 ASIG5V.n3142 0.0102808
R60566 ASIG5V.n8024 ASIG5V.n8023 0.0102808
R60567 ASIG5V.n8027 ASIG5V.n7516 0.0102808
R60568 ASIG5V.n7676 ASIG5V.n7518 0.0102808
R60569 ASIG5V.n7685 ASIG5V.n7684 0.0102808
R60570 ASIG5V.n7683 ASIG5V.n7678 0.0102808
R60571 ASIG5V.n7579 ASIG5V.n7552 0.0102808
R60572 ASIG5V.n7589 ASIG5V.n7588 0.0102808
R60573 ASIG5V.n7591 ASIG5V.n7580 0.0102808
R60574 ASIG5V.n7297 ASIG5V.n7289 0.0102808
R60575 ASIG5V.n8139 ASIG5V.n7298 0.0102808
R60576 ASIG5V.n8138 ASIG5V.n7300 0.0102808
R60577 ASIG5V.n8136 ASIG5V.n8135 0.0102808
R60578 ASIG5V.n8134 ASIG5V.n8131 0.0102808
R60579 ASIG5V.n7458 ASIG5V.n7307 0.0102808
R60580 ASIG5V.n7456 ASIG5V.n7455 0.0102808
R60581 ASIG5V.n7454 ASIG5V.n3034 0.0102808
R60582 ASIG5V.n9929 ASIG5V.n3036 0.0102808
R60583 ASIG5V.n3041 ASIG5V.n3033 0.0102808
R60584 ASIG5V.n9926 ASIG5V.n3042 0.0102808
R60585 ASIG5V.n7298 ASIG5V.n7297 0.0102808
R60586 ASIG5V.n7304 ASIG5V.n7300 0.0102808
R60587 ASIG5V.n7458 ASIG5V.n7457 0.0102808
R60588 ASIG5V.n7455 ASIG5V.n7454 0.0102808
R60589 ASIG5V.n8135 ASIG5V.n8134 0.0102808
R60590 ASIG5V.n7457 ASIG5V.n7456 0.0102808
R60591 ASIG5V.n8136 ASIG5V.n7304 0.0102808
R60592 ASIG5V.n7292 ASIG5V.n7289 0.0102808
R60593 ASIG5V.n7587 ASIG5V.n7579 0.0102808
R60594 ASIG5V.n7588 ASIG5V.n7580 0.0102808
R60595 ASIG5V.n7589 ASIG5V.n7587 0.0102808
R60596 ASIG5V.n7598 ASIG5V.n7597 0.0102808
R60597 ASIG5V.n7601 ASIG5V.n7576 0.0102808
R60598 ASIG5V.n7599 ASIG5V.n7598 0.0102808
R60599 ASIG5V.n7567 ASIG5V.n7563 0.0102808
R60600 ASIG5V.n7650 ASIG5V.n7649 0.0102808
R60601 ASIG5V.n7651 ASIG5V.n7567 0.0102808
R60602 ASIG5V.n8074 ASIG5V.n8073 0.0102808
R60603 ASIG5V.n7493 ASIG5V.n7487 0.0102808
R60604 ASIG5V.n8073 ASIG5V.n8072 0.0102808
R60605 ASIG5V.n9858 ASIG5V.n9857 0.0102808
R60606 ASIG5V.n3105 ASIG5V.n3099 0.0102808
R60607 ASIG5V.n9857 ASIG5V.n9856 0.0102808
R60608 ASIG5V.n9772 ASIG5V.n3144 0.0102808
R60609 ASIG5V.n9769 ASIG5V.n9768 0.0102808
R60610 ASIG5V.n9775 ASIG5V.n3145 0.0102808
R60611 ASIG5V.n7520 ASIG5V.n3147 0.0102808
R60612 ASIG5V.n8013 ASIG5V.n8012 0.0102808
R60613 ASIG5V.n8016 ASIG5V.n7521 0.0102808
R60614 ASIG5V.n7687 ASIG5V.n7523 0.0102808
R60615 ASIG5V.n7696 ASIG5V.n7695 0.0102808
R60616 ASIG5V.n7694 ASIG5V.n7269 0.0102808
R60617 ASIG5V.n7277 ASIG5V.n7268 0.0102808
R60618 ASIG5V.n8152 ASIG5V.n7278 0.0102808
R60619 ASIG5V.n8151 ASIG5V.n7280 0.0102808
R60620 ASIG5V.n8149 ASIG5V.n8148 0.0102808
R60621 ASIG5V.n8147 ASIG5V.n8144 0.0102808
R60622 ASIG5V.n7365 ASIG5V.n7287 0.0102808
R60623 ASIG5V.n7376 ASIG5V.n7375 0.0102808
R60624 ASIG5V.n7374 ASIG5V.n7369 0.0102808
R60625 ASIG5V.n7447 ASIG5V.n7328 0.0102808
R60626 ASIG5V.n7445 ASIG5V.n7444 0.0102808
R60627 ASIG5V.n7443 ASIG5V.n3023 0.0102808
R60628 ASIG5V.n9935 ASIG5V.n3025 0.0102808
R60629 ASIG5V.n3030 ASIG5V.n3022 0.0102808
R60630 ASIG5V.n9932 ASIG5V.n3031 0.0102808
R60631 ASIG5V.n7278 ASIG5V.n7277 0.0102808
R60632 ASIG5V.n7284 ASIG5V.n7280 0.0102808
R60633 ASIG5V.n7366 ASIG5V.n7365 0.0102808
R60634 ASIG5V.n7447 ASIG5V.n7446 0.0102808
R60635 ASIG5V.n7444 ASIG5V.n7443 0.0102808
R60636 ASIG5V.n7375 ASIG5V.n7374 0.0102808
R60637 ASIG5V.n8148 ASIG5V.n8147 0.0102808
R60638 ASIG5V.n7446 ASIG5V.n7445 0.0102808
R60639 ASIG5V.n7376 ASIG5V.n7366 0.0102808
R60640 ASIG5V.n8149 ASIG5V.n7284 0.0102808
R60641 ASIG5V.n7272 ASIG5V.n7268 0.0102808
R60642 ASIG5V.n7687 ASIG5V.n7546 0.0102808
R60643 ASIG5V.n7695 ASIG5V.n7694 0.0102808
R60644 ASIG5V.n7696 ASIG5V.n7546 0.0102808
R60645 ASIG5V.n7676 ASIG5V.n7549 0.0102808
R60646 ASIG5V.n7684 ASIG5V.n7683 0.0102808
R60647 ASIG5V.n7685 ASIG5V.n7549 0.0102808
R60648 ASIG5V.n7665 ASIG5V.n7554 0.0102808
R60649 ASIG5V.n7673 ASIG5V.n7672 0.0102808
R60650 ASIG5V.n7674 ASIG5V.n7554 0.0102808
R60651 ASIG5V.n7654 ASIG5V.n7559 0.0102808
R60652 ASIG5V.n7662 ASIG5V.n7661 0.0102808
R60653 ASIG5V.n7663 ASIG5V.n7559 0.0102808
R60654 ASIG5V.n8065 ASIG5V.n8064 0.0102808
R60655 ASIG5V.n7500 ASIG5V.n7494 0.0102808
R60656 ASIG5V.n8064 ASIG5V.n8063 0.0102808
R60657 ASIG5V.n9849 ASIG5V.n9848 0.0102808
R60658 ASIG5V.n3112 ASIG5V.n3106 0.0102808
R60659 ASIG5V.n9848 ASIG5V.n9847 0.0102808
R60660 ASIG5V.n9755 ASIG5V.n3149 0.0102808
R60661 ASIG5V.n9761 ASIG5V.n9760 0.0102808
R60662 ASIG5V.n9763 ASIG5V.n3150 0.0102808
R60663 ASIG5V.n7525 ASIG5V.n3153 0.0102808
R60664 ASIG5V.n8002 ASIG5V.n8001 0.0102808
R60665 ASIG5V.n8005 ASIG5V.n7526 0.0102808
R60666 ASIG5V.n7703 ASIG5V.n7702 0.0102808
R60667 ASIG5V.n7542 ASIG5V.n7258 0.0102808
R60668 ASIG5V.n8160 ASIG5V.n7260 0.0102808
R60669 ASIG5V.n7265 ASIG5V.n7257 0.0102808
R60670 ASIG5V.n8157 ASIG5V.n7266 0.0102808
R60671 ASIG5V.n7390 ASIG5V.n7350 0.0102808
R60672 ASIG5V.n7355 ASIG5V.n7348 0.0102808
R60673 ASIG5V.n7387 ASIG5V.n7356 0.0102808
R60674 ASIG5V.n7386 ASIG5V.n7358 0.0102808
R60675 ASIG5V.n7384 ASIG5V.n7383 0.0102808
R60676 ASIG5V.n7382 ASIG5V.n7379 0.0102808
R60677 ASIG5V.n7436 ASIG5V.n7332 0.0102808
R60678 ASIG5V.n7434 ASIG5V.n7433 0.0102808
R60679 ASIG5V.n7432 ASIG5V.n3012 0.0102808
R60680 ASIG5V.n9941 ASIG5V.n3014 0.0102808
R60681 ASIG5V.n3019 ASIG5V.n3011 0.0102808
R60682 ASIG5V.n9938 ASIG5V.n3020 0.0102808
R60683 ASIG5V.n7702 ASIG5V.n7542 0.0102808
R60684 ASIG5V.n7264 ASIG5V.n7260 0.0102808
R60685 ASIG5V.n7354 ASIG5V.n7350 0.0102808
R60686 ASIG5V.n7361 ASIG5V.n7358 0.0102808
R60687 ASIG5V.n7436 ASIG5V.n7435 0.0102808
R60688 ASIG5V.n7433 ASIG5V.n7432 0.0102808
R60689 ASIG5V.n7383 ASIG5V.n7382 0.0102808
R60690 ASIG5V.n7356 ASIG5V.n7355 0.0102808
R60691 ASIG5V.n7266 ASIG5V.n7265 0.0102808
R60692 ASIG5V.n7435 ASIG5V.n7434 0.0102808
R60693 ASIG5V.n7384 ASIG5V.n7361 0.0102808
R60694 ASIG5V.n7354 ASIG5V.n7348 0.0102808
R60695 ASIG5V.n7264 ASIG5V.n7257 0.0102808
R60696 ASIG5V.n7703 ASIG5V.n7540 0.0102808
R60697 ASIG5V.n9759 ASIG5V.n3149 0.0102808
R60698 ASIG5V.n9760 ASIG5V.n3150 0.0102808
R60699 ASIG5V.n9761 ASIG5V.n9759 0.0102808
R60700 ASIG5V.n9767 ASIG5V.n3144 0.0102808
R60701 ASIG5V.n9769 ASIG5V.n3145 0.0102808
R60702 ASIG5V.n9768 ASIG5V.n9767 0.0102808
R60703 ASIG5V.n9779 ASIG5V.n3139 0.0102808
R60704 ASIG5V.n9781 ASIG5V.n3140 0.0102808
R60705 ASIG5V.n9780 ASIG5V.n9779 0.0102808
R60706 ASIG5V.n9791 ASIG5V.n3134 0.0102808
R60707 ASIG5V.n9793 ASIG5V.n3135 0.0102808
R60708 ASIG5V.n9792 ASIG5V.n9791 0.0102808
R60709 ASIG5V.n9803 ASIG5V.n3129 0.0102808
R60710 ASIG5V.n9805 ASIG5V.n3130 0.0102808
R60711 ASIG5V.n9804 ASIG5V.n9803 0.0102808
R60712 ASIG5V.n9815 ASIG5V.n3124 0.0102808
R60713 ASIG5V.n9817 ASIG5V.n3125 0.0102808
R60714 ASIG5V.n9816 ASIG5V.n9815 0.0102808
R60715 ASIG5V.n9831 ASIG5V.n9830 0.0102808
R60716 ASIG5V.n9828 ASIG5V.n3120 0.0102808
R60717 ASIG5V.n9830 ASIG5V.n9829 0.0102808
R60718 ASIG5V.n9751 ASIG5V.n9750 0.0102808
R60719 ASIG5V.n7988 ASIG5V.n3155 0.0102808
R60720 ASIG5V.n7991 ASIG5V.n7530 0.0102808
R60721 ASIG5V.n7987 ASIG5V.n7986 0.0102808
R60722 ASIG5V.n7994 ASIG5V.n7531 0.0102808
R60723 ASIG5V.n7713 ASIG5V.n7534 0.0102808
R60724 ASIG5V.n7711 ASIG5V.n7710 0.0102808
R60725 ASIG5V.n7709 ASIG5V.n7247 0.0102808
R60726 ASIG5V.n8166 ASIG5V.n7249 0.0102808
R60727 ASIG5V.n7254 ASIG5V.n7246 0.0102808
R60728 ASIG5V.n8163 ASIG5V.n7255 0.0102808
R60729 ASIG5V.n7401 ASIG5V.n7398 0.0102808
R60730 ASIG5V.n7396 ASIG5V.n7395 0.0102808
R60731 ASIG5V.n7404 ASIG5V.n7345 0.0102808
R60732 ASIG5V.n7410 ASIG5V.n7407 0.0102808
R60733 ASIG5V.n7405 ASIG5V.n7344 0.0102808
R60734 ASIG5V.n7413 ASIG5V.n7336 0.0102808
R60735 ASIG5V.n7425 ASIG5V.n7414 0.0102808
R60736 ASIG5V.n7423 ASIG5V.n7422 0.0102808
R60737 ASIG5V.n7421 ASIG5V.n3009 0.0102808
R60738 ASIG5V.n9945 ASIG5V.n9944 0.0102808
R60739 ASIG5V.n9951 ASIG5V.n9950 0.0102808
R60740 ASIG5V.n9949 ASIG5V.n3004 0.0102808
R60741 ASIG5V.n9750 ASIG5V.n3155 0.0102808
R60742 ASIG5V.n7537 ASIG5V.n7534 0.0102808
R60743 ASIG5V.n7253 ASIG5V.n7249 0.0102808
R60744 ASIG5V.n7398 ASIG5V.n7397 0.0102808
R60745 ASIG5V.n7407 ASIG5V.n7406 0.0102808
R60746 ASIG5V.n7425 ASIG5V.n7424 0.0102808
R60747 ASIG5V.n7422 ASIG5V.n7421 0.0102808
R60748 ASIG5V.n7344 ASIG5V.n7336 0.0102808
R60749 ASIG5V.n7395 ASIG5V.n7345 0.0102808
R60750 ASIG5V.n7255 ASIG5V.n7254 0.0102808
R60751 ASIG5V.n7710 ASIG5V.n7709 0.0102808
R60752 ASIG5V.n7424 ASIG5V.n7423 0.0102808
R60753 ASIG5V.n7406 ASIG5V.n7405 0.0102808
R60754 ASIG5V.n7397 ASIG5V.n7396 0.0102808
R60755 ASIG5V.n7253 ASIG5V.n7246 0.0102808
R60756 ASIG5V.n7711 ASIG5V.n7537 0.0102808
R60757 ASIG5V.n9751 ASIG5V.n3159 0.0102808
R60758 ASIG5V.n9944 ASIG5V.n3005 0.0102808
R60759 ASIG5V.n9950 ASIG5V.n9949 0.0102808
R60760 ASIG5V.n9951 ASIG5V.n3005 0.0102808
R60761 ASIG5V.n3018 ASIG5V.n3014 0.0102808
R60762 ASIG5V.n3020 ASIG5V.n3019 0.0102808
R60763 ASIG5V.n3018 ASIG5V.n3011 0.0102808
R60764 ASIG5V.n3029 ASIG5V.n3025 0.0102808
R60765 ASIG5V.n3031 ASIG5V.n3030 0.0102808
R60766 ASIG5V.n3029 ASIG5V.n3022 0.0102808
R60767 ASIG5V.n3040 ASIG5V.n3036 0.0102808
R60768 ASIG5V.n3042 ASIG5V.n3041 0.0102808
R60769 ASIG5V.n3040 ASIG5V.n3033 0.0102808
R60770 ASIG5V.n3051 ASIG5V.n3047 0.0102808
R60771 ASIG5V.n3053 ASIG5V.n3052 0.0102808
R60772 ASIG5V.n3051 ASIG5V.n3044 0.0102808
R60773 ASIG5V.n3062 ASIG5V.n3058 0.0102808
R60774 ASIG5V.n3064 ASIG5V.n3063 0.0102808
R60775 ASIG5V.n3062 ASIG5V.n3055 0.0102808
R60776 ASIG5V.n3073 ASIG5V.n3069 0.0102808
R60777 ASIG5V.n3075 ASIG5V.n3074 0.0102808
R60778 ASIG5V.n3073 ASIG5V.n3066 0.0102808
R60779 ASIG5V.n9898 ASIG5V.n9894 0.0102808
R60780 ASIG5V.n9900 ASIG5V.n9899 0.0102808
R60781 ASIG5V.n9898 ASIG5V.n3077 0.0102808
R60782 ASIG5V.n7985 ASIG5V.n7530 0.0102808
R60783 ASIG5V.n7987 ASIG5V.n7531 0.0102808
R60784 ASIG5V.n7986 ASIG5V.n7985 0.0102808
R60785 ASIG5V.n8000 ASIG5V.n7525 0.0102808
R60786 ASIG5V.n8002 ASIG5V.n7526 0.0102808
R60787 ASIG5V.n8001 ASIG5V.n8000 0.0102808
R60788 ASIG5V.n8011 ASIG5V.n7520 0.0102808
R60789 ASIG5V.n8013 ASIG5V.n7521 0.0102808
R60790 ASIG5V.n8012 ASIG5V.n8011 0.0102808
R60791 ASIG5V.n8022 ASIG5V.n7515 0.0102808
R60792 ASIG5V.n8024 ASIG5V.n7516 0.0102808
R60793 ASIG5V.n8023 ASIG5V.n8022 0.0102808
R60794 ASIG5V.n8033 ASIG5V.n7510 0.0102808
R60795 ASIG5V.n8035 ASIG5V.n7511 0.0102808
R60796 ASIG5V.n8034 ASIG5V.n8033 0.0102808
R60797 ASIG5V.n8044 ASIG5V.n7505 0.0102808
R60798 ASIG5V.n8046 ASIG5V.n7506 0.0102808
R60799 ASIG5V.n8045 ASIG5V.n8044 0.0102808
R60800 ASIG5V.n8056 ASIG5V.n8055 0.0102808
R60801 ASIG5V.n8059 ASIG5V.n7501 0.0102808
R60802 ASIG5V.n8057 ASIG5V.n8056 0.0102808
R60803 ASIG5V.n9840 ASIG5V.n9839 0.0102808
R60804 ASIG5V.n3119 ASIG5V.n3113 0.0102808
R60805 ASIG5V.n9839 ASIG5V.n9838 0.0102808
R60806 ASIG5V.n8923 ASIG5V.n6540 0.0102444
R60807 ASIG5V.n10925 ASIG5V.n10924 0.0102444
R60808 ASIG5V.n6439 ASIG5V.n6259 0.010175
R60809 ASIG5V.n10915 ASIG5V.n10914 0.010175
R60810 ASIG5V.n6539 ASIG5V.n6538 0.0101644
R60811 ASIG5V.n8927 ASIG5V.n8926 0.0101644
R60812 ASIG5V.n4558 ASIG5V.n3831 0.0101288
R60813 ASIG5V.n4559 ASIG5V.n3835 0.0101288
R60814 ASIG5V.n6881 ASIG5V.n6633 0.00973581
R60815 ASIG5V.n8913 ASIG5V.n6882 0.00973581
R60816 ASIG5V.n4792 ASIG5V.n4791 0.00970301
R60817 ASIG5V.n7972 ASIG5V.n7971 0.00970301
R60818 ASIG5V.n1321 ASIG5V.n1320 0.00968121
R60819 ASIG5V.n12013 ASIG5V.n1325 0.00968121
R60820 ASIG5V.n12019 ASIG5V.n12018 0.00968121
R60821 ASIG5V.n12014 ASIG5V.n1323 0.00968121
R60822 ASIG5V.n1667 ASIG5V.n1416 0.00934279
R60823 ASIG5V.n2201 ASIG5V.n1863 0.00934279
R60824 ASIG5V.n12005 ASIG5V.n12004 0.00934279
R60825 ASIG5V.n2202 ASIG5V.n1857 0.00934279
R60826 ASIG5V.n8921 ASIG5V.n6543 0.00919799
R60827 ASIG5V.n10922 ASIG5V.n10480 0.00919799
R60828 ASIG5V.n8922 ASIG5V.n6541 0.00919799
R60829 ASIG5V.n10923 ASIG5V.n10468 0.00919799
R60830 ASIG5V.n12337 ASIG5V.n12336 0.00916165
R60831 ASIG5V.n11777 ASIG5V.n11776 0.00916165
R60832 ASIG5V.n6437 ASIG5V.n6262 0.00894978
R60833 ASIG5V.n10491 ASIG5V.n10485 0.00894978
R60834 ASIG5V.n6438 ASIG5V.n6260 0.00894978
R60835 ASIG5V.n10490 ASIG5V.n10487 0.00894978
R60836 ASIG5V.n4789 ASIG5V.n3279 0.00871477
R60837 ASIG5V.n7974 ASIG5V.n5508 0.00871477
R60838 ASIG5V.n4790 ASIG5V.n3280 0.00871477
R60839 ASIG5V.n7973 ASIG5V.n7716 0.00871477
R60840 ASIG5V.n10813 ASIG5V.n10490 0.0087125
R60841 ASIG5V.n10548 ASIG5V.n10491 0.0087125
R60842 ASIG5V.n4252 ASIG5V.n4251 0.0087125
R60843 ASIG5V.n4254 ASIG5V.n4253 0.0087125
R60844 ASIG5V ASIG5V.t7 0.0086761
R60845 ASIG5V ASIG5V.t5 0.0086761
R60846 ASIG5V ASIG5V.t3 0.0086761
R60847 ASIG5V ASIG5V.t2 0.0086761
R60848 ASIG5V.n12337 ASIG5V.n161 0.0086203
R60849 ASIG5V.n11776 ASIG5V.n11775 0.0086203
R60850 ASIG5V.n5562 ASIG5V.n5561 0.008375
R60851 ASIG5V.n12334 ASIG5V.n54 0.00823154
R60852 ASIG5V.n2567 ASIG5V.n2215 0.00823154
R60853 ASIG5V.n12335 ASIG5V.n163 0.00823154
R60854 ASIG5V.n2565 ASIG5V.n2217 0.00823154
R60855 ASIG5V.n4795 ASIG5V.n4792 0.00807895
R60856 ASIG5V.n7971 ASIG5V.n7970 0.00807895
R60857 ASIG5V.n10702 ASIG5V.n10698 0.00796421
R60858 ASIG5V.n10713 ASIG5V.n10695 0.00796421
R60859 ASIG5V.n10910 ASIG5V.n10690 0.00796421
R60860 ASIG5V.n10691 ASIG5V.n10498 0.00796421
R60861 ASIG5V.n10689 ASIG5V.n10687 0.00796421
R60862 ASIG5V.n10688 ASIG5V.n10499 0.00796421
R60863 ASIG5V.n10686 ASIG5V.n10684 0.00796421
R60864 ASIG5V.n10685 ASIG5V.n10500 0.00796421
R60865 ASIG5V.n10683 ASIG5V.n10681 0.00796421
R60866 ASIG5V.n10682 ASIG5V.n10501 0.00796421
R60867 ASIG5V.n10680 ASIG5V.n10678 0.00796421
R60868 ASIG5V.n10679 ASIG5V.n10502 0.00796421
R60869 ASIG5V.n10677 ASIG5V.n10675 0.00796421
R60870 ASIG5V.n10676 ASIG5V.n10503 0.00796421
R60871 ASIG5V.n10674 ASIG5V.n10672 0.00796421
R60872 ASIG5V.n10673 ASIG5V.n10504 0.00796421
R60873 ASIG5V.n10671 ASIG5V.n10669 0.00796421
R60874 ASIG5V.n10670 ASIG5V.n10505 0.00796421
R60875 ASIG5V.n10668 ASIG5V.n10666 0.00796421
R60876 ASIG5V.n10667 ASIG5V.n10506 0.00796421
R60877 ASIG5V.n10665 ASIG5V.n10663 0.00796421
R60878 ASIG5V.n10664 ASIG5V.n10507 0.00796421
R60879 ASIG5V.n10662 ASIG5V.n10660 0.00796421
R60880 ASIG5V.n10661 ASIG5V.n10508 0.00796421
R60881 ASIG5V.n10659 ASIG5V.n10657 0.00796421
R60882 ASIG5V.n10658 ASIG5V.n10509 0.00796421
R60883 ASIG5V.n10656 ASIG5V.n10654 0.00796421
R60884 ASIG5V.n10655 ASIG5V.n10510 0.00796421
R60885 ASIG5V.n10653 ASIG5V.n10651 0.00796421
R60886 ASIG5V.n10652 ASIG5V.n10511 0.00796421
R60887 ASIG5V.n10650 ASIG5V.n10648 0.00796421
R60888 ASIG5V.n10649 ASIG5V.n10512 0.00796421
R60889 ASIG5V.n10647 ASIG5V.n10645 0.00796421
R60890 ASIG5V.n10646 ASIG5V.n10513 0.00796421
R60891 ASIG5V.n10644 ASIG5V.n10642 0.00796421
R60892 ASIG5V.n10643 ASIG5V.n10514 0.00796421
R60893 ASIG5V.n10641 ASIG5V.n10639 0.00796421
R60894 ASIG5V.n10640 ASIG5V.n10515 0.00796421
R60895 ASIG5V.n10638 ASIG5V.n10636 0.00796421
R60896 ASIG5V.n10637 ASIG5V.n10516 0.00796421
R60897 ASIG5V.n10635 ASIG5V.n10633 0.00796421
R60898 ASIG5V.n10634 ASIG5V.n10517 0.00796421
R60899 ASIG5V.n10632 ASIG5V.n10630 0.00796421
R60900 ASIG5V.n10631 ASIG5V.n10518 0.00796421
R60901 ASIG5V.n10629 ASIG5V.n10627 0.00796421
R60902 ASIG5V.n10628 ASIG5V.n10519 0.00796421
R60903 ASIG5V.n10626 ASIG5V.n10624 0.00796421
R60904 ASIG5V.n10625 ASIG5V.n10520 0.00796421
R60905 ASIG5V.n10623 ASIG5V.n10621 0.00796421
R60906 ASIG5V.n10622 ASIG5V.n10521 0.00796421
R60907 ASIG5V.n10620 ASIG5V.n10618 0.00796421
R60908 ASIG5V.n10619 ASIG5V.n10522 0.00796421
R60909 ASIG5V.n10617 ASIG5V.n10615 0.00796421
R60910 ASIG5V.n10616 ASIG5V.n10523 0.00796421
R60911 ASIG5V.n10614 ASIG5V.n10612 0.00796421
R60912 ASIG5V.n10613 ASIG5V.n10524 0.00796421
R60913 ASIG5V.n10611 ASIG5V.n10609 0.00796421
R60914 ASIG5V.n10610 ASIG5V.n10525 0.00796421
R60915 ASIG5V.n10608 ASIG5V.n10606 0.00796421
R60916 ASIG5V.n10607 ASIG5V.n10526 0.00796421
R60917 ASIG5V.n10605 ASIG5V.n10603 0.00796421
R60918 ASIG5V.n10604 ASIG5V.n10527 0.00796421
R60919 ASIG5V.n10602 ASIG5V.n10600 0.00796421
R60920 ASIG5V.n10601 ASIG5V.n10528 0.00796421
R60921 ASIG5V.n10599 ASIG5V.n10597 0.00796421
R60922 ASIG5V.n10598 ASIG5V.n10529 0.00796421
R60923 ASIG5V.n10596 ASIG5V.n10594 0.00796421
R60924 ASIG5V.n10595 ASIG5V.n10530 0.00796421
R60925 ASIG5V.n10593 ASIG5V.n10591 0.00796421
R60926 ASIG5V.n10592 ASIG5V.n10531 0.00796421
R60927 ASIG5V.n10590 ASIG5V.n10588 0.00796421
R60928 ASIG5V.n10589 ASIG5V.n10532 0.00796421
R60929 ASIG5V.n10587 ASIG5V.n10585 0.00796421
R60930 ASIG5V.n10586 ASIG5V.n10533 0.00796421
R60931 ASIG5V.n10584 ASIG5V.n10582 0.00796421
R60932 ASIG5V.n10583 ASIG5V.n10534 0.00796421
R60933 ASIG5V.n10581 ASIG5V.n10579 0.00796421
R60934 ASIG5V.n10580 ASIG5V.n10535 0.00796421
R60935 ASIG5V.n10578 ASIG5V.n10576 0.00796421
R60936 ASIG5V.n10577 ASIG5V.n10536 0.00796421
R60937 ASIG5V.n10575 ASIG5V.n10573 0.00796421
R60938 ASIG5V.n10574 ASIG5V.n10537 0.00796421
R60939 ASIG5V.n10572 ASIG5V.n10570 0.00796421
R60940 ASIG5V.n10571 ASIG5V.n10538 0.00796421
R60941 ASIG5V.n10569 ASIG5V.n10567 0.00796421
R60942 ASIG5V.n10568 ASIG5V.n10539 0.00796421
R60943 ASIG5V.n10566 ASIG5V.n10564 0.00796421
R60944 ASIG5V.n10565 ASIG5V.n10540 0.00796421
R60945 ASIG5V.n10563 ASIG5V.n10561 0.00796421
R60946 ASIG5V.n10562 ASIG5V.n10541 0.00796421
R60947 ASIG5V.n10560 ASIG5V.n10558 0.00796421
R60948 ASIG5V.n10559 ASIG5V.n10542 0.00796421
R60949 ASIG5V.n10557 ASIG5V.n10555 0.00796421
R60950 ASIG5V.n10556 ASIG5V.n10543 0.00796421
R60951 ASIG5V.n10554 ASIG5V.n10552 0.00796421
R60952 ASIG5V.n10553 ASIG5V.n10544 0.00796421
R60953 ASIG5V.n10551 ASIG5V.n10549 0.00796421
R60954 ASIG5V.n10550 ASIG5V.n10545 0.00796421
R60955 ASIG5V.n10548 ASIG5V.n10547 0.00796421
R60956 ASIG5V.n4258 ASIG5V.n3853 0.00796421
R60957 ASIG5V.n4257 ASIG5V.n3846 0.00796421
R60958 ASIG5V.n3906 ASIG5V.n3854 0.00796421
R60959 ASIG5V.n3911 ASIG5V.n3910 0.00796421
R60960 ASIG5V.n4050 ASIG5V.n3905 0.00796421
R60961 ASIG5V.n3913 ASIG5V.n3912 0.00796421
R60962 ASIG5V.n4049 ASIG5V.n3904 0.00796421
R60963 ASIG5V.n3915 ASIG5V.n3914 0.00796421
R60964 ASIG5V.n4048 ASIG5V.n3903 0.00796421
R60965 ASIG5V.n3917 ASIG5V.n3916 0.00796421
R60966 ASIG5V.n4047 ASIG5V.n3902 0.00796421
R60967 ASIG5V.n3919 ASIG5V.n3918 0.00796421
R60968 ASIG5V.n4046 ASIG5V.n3901 0.00796421
R60969 ASIG5V.n3921 ASIG5V.n3920 0.00796421
R60970 ASIG5V.n4045 ASIG5V.n3900 0.00796421
R60971 ASIG5V.n3923 ASIG5V.n3922 0.00796421
R60972 ASIG5V.n4044 ASIG5V.n3899 0.00796421
R60973 ASIG5V.n3925 ASIG5V.n3924 0.00796421
R60974 ASIG5V.n4043 ASIG5V.n3898 0.00796421
R60975 ASIG5V.n3927 ASIG5V.n3926 0.00796421
R60976 ASIG5V.n4042 ASIG5V.n3897 0.00796421
R60977 ASIG5V.n3929 ASIG5V.n3928 0.00796421
R60978 ASIG5V.n4041 ASIG5V.n3896 0.00796421
R60979 ASIG5V.n3931 ASIG5V.n3930 0.00796421
R60980 ASIG5V.n4040 ASIG5V.n3895 0.00796421
R60981 ASIG5V.n3933 ASIG5V.n3932 0.00796421
R60982 ASIG5V.n4039 ASIG5V.n3894 0.00796421
R60983 ASIG5V.n3935 ASIG5V.n3934 0.00796421
R60984 ASIG5V.n4038 ASIG5V.n3893 0.00796421
R60985 ASIG5V.n3937 ASIG5V.n3936 0.00796421
R60986 ASIG5V.n4037 ASIG5V.n3892 0.00796421
R60987 ASIG5V.n3939 ASIG5V.n3938 0.00796421
R60988 ASIG5V.n4036 ASIG5V.n3891 0.00796421
R60989 ASIG5V.n3941 ASIG5V.n3940 0.00796421
R60990 ASIG5V.n4035 ASIG5V.n3890 0.00796421
R60991 ASIG5V.n3943 ASIG5V.n3942 0.00796421
R60992 ASIG5V.n4034 ASIG5V.n3889 0.00796421
R60993 ASIG5V.n3945 ASIG5V.n3944 0.00796421
R60994 ASIG5V.n4033 ASIG5V.n3888 0.00796421
R60995 ASIG5V.n3947 ASIG5V.n3946 0.00796421
R60996 ASIG5V.n4032 ASIG5V.n3887 0.00796421
R60997 ASIG5V.n3949 ASIG5V.n3948 0.00796421
R60998 ASIG5V.n4031 ASIG5V.n3886 0.00796421
R60999 ASIG5V.n3951 ASIG5V.n3950 0.00796421
R61000 ASIG5V.n4030 ASIG5V.n3885 0.00796421
R61001 ASIG5V.n3953 ASIG5V.n3952 0.00796421
R61002 ASIG5V.n4029 ASIG5V.n3884 0.00796421
R61003 ASIG5V.n3955 ASIG5V.n3954 0.00796421
R61004 ASIG5V.n4028 ASIG5V.n3883 0.00796421
R61005 ASIG5V.n3957 ASIG5V.n3956 0.00796421
R61006 ASIG5V.n4027 ASIG5V.n3882 0.00796421
R61007 ASIG5V.n3959 ASIG5V.n3958 0.00796421
R61008 ASIG5V.n4026 ASIG5V.n3881 0.00796421
R61009 ASIG5V.n3961 ASIG5V.n3960 0.00796421
R61010 ASIG5V.n4025 ASIG5V.n3880 0.00796421
R61011 ASIG5V.n3963 ASIG5V.n3962 0.00796421
R61012 ASIG5V.n4024 ASIG5V.n3879 0.00796421
R61013 ASIG5V.n3965 ASIG5V.n3964 0.00796421
R61014 ASIG5V.n4023 ASIG5V.n3878 0.00796421
R61015 ASIG5V.n3967 ASIG5V.n3966 0.00796421
R61016 ASIG5V.n4022 ASIG5V.n3877 0.00796421
R61017 ASIG5V.n3969 ASIG5V.n3968 0.00796421
R61018 ASIG5V.n4021 ASIG5V.n3876 0.00796421
R61019 ASIG5V.n3971 ASIG5V.n3970 0.00796421
R61020 ASIG5V.n4020 ASIG5V.n3875 0.00796421
R61021 ASIG5V.n3973 ASIG5V.n3972 0.00796421
R61022 ASIG5V.n4019 ASIG5V.n3874 0.00796421
R61023 ASIG5V.n3975 ASIG5V.n3974 0.00796421
R61024 ASIG5V.n4018 ASIG5V.n3873 0.00796421
R61025 ASIG5V.n3977 ASIG5V.n3976 0.00796421
R61026 ASIG5V.n4017 ASIG5V.n3872 0.00796421
R61027 ASIG5V.n3979 ASIG5V.n3978 0.00796421
R61028 ASIG5V.n4016 ASIG5V.n3871 0.00796421
R61029 ASIG5V.n3981 ASIG5V.n3980 0.00796421
R61030 ASIG5V.n4015 ASIG5V.n3870 0.00796421
R61031 ASIG5V.n3983 ASIG5V.n3982 0.00796421
R61032 ASIG5V.n4014 ASIG5V.n3869 0.00796421
R61033 ASIG5V.n3985 ASIG5V.n3984 0.00796421
R61034 ASIG5V.n4013 ASIG5V.n3868 0.00796421
R61035 ASIG5V.n3987 ASIG5V.n3986 0.00796421
R61036 ASIG5V.n4012 ASIG5V.n3867 0.00796421
R61037 ASIG5V.n3989 ASIG5V.n3988 0.00796421
R61038 ASIG5V.n4011 ASIG5V.n3866 0.00796421
R61039 ASIG5V.n3991 ASIG5V.n3990 0.00796421
R61040 ASIG5V.n4010 ASIG5V.n3865 0.00796421
R61041 ASIG5V.n3993 ASIG5V.n3992 0.00796421
R61042 ASIG5V.n4009 ASIG5V.n3864 0.00796421
R61043 ASIG5V.n3995 ASIG5V.n3994 0.00796421
R61044 ASIG5V.n4008 ASIG5V.n3863 0.00796421
R61045 ASIG5V.n3997 ASIG5V.n3996 0.00796421
R61046 ASIG5V.n4007 ASIG5V.n3862 0.00796421
R61047 ASIG5V.n3999 ASIG5V.n3998 0.00796421
R61048 ASIG5V.n4006 ASIG5V.n3861 0.00796421
R61049 ASIG5V.n4001 ASIG5V.n4000 0.00796421
R61050 ASIG5V.n4005 ASIG5V.n3860 0.00796421
R61051 ASIG5V.n4003 ASIG5V.n4002 0.00796421
R61052 ASIG5V.n4004 ASIG5V.n3859 0.00796421
R61053 ASIG5V.n3908 ASIG5V.n3907 0.00796421
R61054 ASIG5V.n4254 ASIG5V.n4052 0.00796421
R61055 ASIG5V.n4052 ASIG5V.n3908 0.00796421
R61056 ASIG5V.n10547 ASIG5V.n10545 0.00796421
R61057 ASIG5V.n10551 ASIG5V.n10550 0.00796421
R61058 ASIG5V.n10549 ASIG5V.n10544 0.00796421
R61059 ASIG5V.n10554 ASIG5V.n10553 0.00796421
R61060 ASIG5V.n10552 ASIG5V.n10543 0.00796421
R61061 ASIG5V.n10557 ASIG5V.n10556 0.00796421
R61062 ASIG5V.n10555 ASIG5V.n10542 0.00796421
R61063 ASIG5V.n10560 ASIG5V.n10559 0.00796421
R61064 ASIG5V.n10558 ASIG5V.n10541 0.00796421
R61065 ASIG5V.n10563 ASIG5V.n10562 0.00796421
R61066 ASIG5V.n10561 ASIG5V.n10540 0.00796421
R61067 ASIG5V.n10566 ASIG5V.n10565 0.00796421
R61068 ASIG5V.n10564 ASIG5V.n10539 0.00796421
R61069 ASIG5V.n10569 ASIG5V.n10568 0.00796421
R61070 ASIG5V.n10567 ASIG5V.n10538 0.00796421
R61071 ASIG5V.n10572 ASIG5V.n10571 0.00796421
R61072 ASIG5V.n10570 ASIG5V.n10537 0.00796421
R61073 ASIG5V.n10575 ASIG5V.n10574 0.00796421
R61074 ASIG5V.n10573 ASIG5V.n10536 0.00796421
R61075 ASIG5V.n10578 ASIG5V.n10577 0.00796421
R61076 ASIG5V.n10576 ASIG5V.n10535 0.00796421
R61077 ASIG5V.n10581 ASIG5V.n10580 0.00796421
R61078 ASIG5V.n10579 ASIG5V.n10534 0.00796421
R61079 ASIG5V.n10584 ASIG5V.n10583 0.00796421
R61080 ASIG5V.n10582 ASIG5V.n10533 0.00796421
R61081 ASIG5V.n10587 ASIG5V.n10586 0.00796421
R61082 ASIG5V.n10585 ASIG5V.n10532 0.00796421
R61083 ASIG5V.n10590 ASIG5V.n10589 0.00796421
R61084 ASIG5V.n10588 ASIG5V.n10531 0.00796421
R61085 ASIG5V.n10593 ASIG5V.n10592 0.00796421
R61086 ASIG5V.n10591 ASIG5V.n10530 0.00796421
R61087 ASIG5V.n10596 ASIG5V.n10595 0.00796421
R61088 ASIG5V.n10594 ASIG5V.n10529 0.00796421
R61089 ASIG5V.n10599 ASIG5V.n10598 0.00796421
R61090 ASIG5V.n10597 ASIG5V.n10528 0.00796421
R61091 ASIG5V.n10602 ASIG5V.n10601 0.00796421
R61092 ASIG5V.n10600 ASIG5V.n10527 0.00796421
R61093 ASIG5V.n10605 ASIG5V.n10604 0.00796421
R61094 ASIG5V.n10603 ASIG5V.n10526 0.00796421
R61095 ASIG5V.n10608 ASIG5V.n10607 0.00796421
R61096 ASIG5V.n10606 ASIG5V.n10525 0.00796421
R61097 ASIG5V.n10611 ASIG5V.n10610 0.00796421
R61098 ASIG5V.n10609 ASIG5V.n10524 0.00796421
R61099 ASIG5V.n10614 ASIG5V.n10613 0.00796421
R61100 ASIG5V.n10612 ASIG5V.n10523 0.00796421
R61101 ASIG5V.n10617 ASIG5V.n10616 0.00796421
R61102 ASIG5V.n10615 ASIG5V.n10522 0.00796421
R61103 ASIG5V.n10620 ASIG5V.n10619 0.00796421
R61104 ASIG5V.n10618 ASIG5V.n10521 0.00796421
R61105 ASIG5V.n10623 ASIG5V.n10622 0.00796421
R61106 ASIG5V.n10621 ASIG5V.n10520 0.00796421
R61107 ASIG5V.n10626 ASIG5V.n10625 0.00796421
R61108 ASIG5V.n10624 ASIG5V.n10519 0.00796421
R61109 ASIG5V.n10629 ASIG5V.n10628 0.00796421
R61110 ASIG5V.n10627 ASIG5V.n10518 0.00796421
R61111 ASIG5V.n10632 ASIG5V.n10631 0.00796421
R61112 ASIG5V.n10630 ASIG5V.n10517 0.00796421
R61113 ASIG5V.n10635 ASIG5V.n10634 0.00796421
R61114 ASIG5V.n10633 ASIG5V.n10516 0.00796421
R61115 ASIG5V.n10638 ASIG5V.n10637 0.00796421
R61116 ASIG5V.n10636 ASIG5V.n10515 0.00796421
R61117 ASIG5V.n10641 ASIG5V.n10640 0.00796421
R61118 ASIG5V.n10639 ASIG5V.n10514 0.00796421
R61119 ASIG5V.n10644 ASIG5V.n10643 0.00796421
R61120 ASIG5V.n10642 ASIG5V.n10513 0.00796421
R61121 ASIG5V.n10647 ASIG5V.n10646 0.00796421
R61122 ASIG5V.n10645 ASIG5V.n10512 0.00796421
R61123 ASIG5V.n10650 ASIG5V.n10649 0.00796421
R61124 ASIG5V.n10648 ASIG5V.n10511 0.00796421
R61125 ASIG5V.n10653 ASIG5V.n10652 0.00796421
R61126 ASIG5V.n10651 ASIG5V.n10510 0.00796421
R61127 ASIG5V.n10656 ASIG5V.n10655 0.00796421
R61128 ASIG5V.n10654 ASIG5V.n10509 0.00796421
R61129 ASIG5V.n10659 ASIG5V.n10658 0.00796421
R61130 ASIG5V.n10657 ASIG5V.n10508 0.00796421
R61131 ASIG5V.n10662 ASIG5V.n10661 0.00796421
R61132 ASIG5V.n10660 ASIG5V.n10507 0.00796421
R61133 ASIG5V.n10665 ASIG5V.n10664 0.00796421
R61134 ASIG5V.n10663 ASIG5V.n10506 0.00796421
R61135 ASIG5V.n10668 ASIG5V.n10667 0.00796421
R61136 ASIG5V.n10666 ASIG5V.n10505 0.00796421
R61137 ASIG5V.n10671 ASIG5V.n10670 0.00796421
R61138 ASIG5V.n10669 ASIG5V.n10504 0.00796421
R61139 ASIG5V.n10674 ASIG5V.n10673 0.00796421
R61140 ASIG5V.n10672 ASIG5V.n10503 0.00796421
R61141 ASIG5V.n10677 ASIG5V.n10676 0.00796421
R61142 ASIG5V.n10675 ASIG5V.n10502 0.00796421
R61143 ASIG5V.n10680 ASIG5V.n10679 0.00796421
R61144 ASIG5V.n10678 ASIG5V.n10501 0.00796421
R61145 ASIG5V.n10683 ASIG5V.n10682 0.00796421
R61146 ASIG5V.n10681 ASIG5V.n10500 0.00796421
R61147 ASIG5V.n10686 ASIG5V.n10685 0.00796421
R61148 ASIG5V.n10684 ASIG5V.n10499 0.00796421
R61149 ASIG5V.n10689 ASIG5V.n10688 0.00796421
R61150 ASIG5V.n10687 ASIG5V.n10498 0.00796421
R61151 ASIG5V.n10910 ASIG5V.n10691 0.00796421
R61152 ASIG5V.n10690 ASIG5V.n10497 0.00796421
R61153 ASIG5V.n4261 ASIG5V.n3846 0.00796421
R61154 ASIG5V.n10700 ASIG5V.n10695 0.00796421
R61155 ASIG5V.n4259 ASIG5V.n4258 0.00796421
R61156 ASIG5V.n10711 ASIG5V.n10702 0.00796421
R61157 ASIG5V.n4256 ASIG5V.n3854 0.00796421
R61158 ASIG5V.n3910 ASIG5V.n3906 0.00796421
R61159 ASIG5V.n4050 ASIG5V.n3911 0.00796421
R61160 ASIG5V.n3912 ASIG5V.n3905 0.00796421
R61161 ASIG5V.n4049 ASIG5V.n3913 0.00796421
R61162 ASIG5V.n3914 ASIG5V.n3904 0.00796421
R61163 ASIG5V.n4048 ASIG5V.n3915 0.00796421
R61164 ASIG5V.n3916 ASIG5V.n3903 0.00796421
R61165 ASIG5V.n4047 ASIG5V.n3917 0.00796421
R61166 ASIG5V.n3918 ASIG5V.n3902 0.00796421
R61167 ASIG5V.n4046 ASIG5V.n3919 0.00796421
R61168 ASIG5V.n3920 ASIG5V.n3901 0.00796421
R61169 ASIG5V.n4045 ASIG5V.n3921 0.00796421
R61170 ASIG5V.n3922 ASIG5V.n3900 0.00796421
R61171 ASIG5V.n4044 ASIG5V.n3923 0.00796421
R61172 ASIG5V.n3924 ASIG5V.n3899 0.00796421
R61173 ASIG5V.n4043 ASIG5V.n3925 0.00796421
R61174 ASIG5V.n3926 ASIG5V.n3898 0.00796421
R61175 ASIG5V.n4042 ASIG5V.n3927 0.00796421
R61176 ASIG5V.n3928 ASIG5V.n3897 0.00796421
R61177 ASIG5V.n4041 ASIG5V.n3929 0.00796421
R61178 ASIG5V.n3930 ASIG5V.n3896 0.00796421
R61179 ASIG5V.n4040 ASIG5V.n3931 0.00796421
R61180 ASIG5V.n3932 ASIG5V.n3895 0.00796421
R61181 ASIG5V.n4039 ASIG5V.n3933 0.00796421
R61182 ASIG5V.n3934 ASIG5V.n3894 0.00796421
R61183 ASIG5V.n4038 ASIG5V.n3935 0.00796421
R61184 ASIG5V.n3936 ASIG5V.n3893 0.00796421
R61185 ASIG5V.n4037 ASIG5V.n3937 0.00796421
R61186 ASIG5V.n3938 ASIG5V.n3892 0.00796421
R61187 ASIG5V.n4036 ASIG5V.n3939 0.00796421
R61188 ASIG5V.n3940 ASIG5V.n3891 0.00796421
R61189 ASIG5V.n4035 ASIG5V.n3941 0.00796421
R61190 ASIG5V.n3942 ASIG5V.n3890 0.00796421
R61191 ASIG5V.n4034 ASIG5V.n3943 0.00796421
R61192 ASIG5V.n3944 ASIG5V.n3889 0.00796421
R61193 ASIG5V.n4033 ASIG5V.n3945 0.00796421
R61194 ASIG5V.n3946 ASIG5V.n3888 0.00796421
R61195 ASIG5V.n4032 ASIG5V.n3947 0.00796421
R61196 ASIG5V.n3948 ASIG5V.n3887 0.00796421
R61197 ASIG5V.n4031 ASIG5V.n3949 0.00796421
R61198 ASIG5V.n3950 ASIG5V.n3886 0.00796421
R61199 ASIG5V.n4030 ASIG5V.n3951 0.00796421
R61200 ASIG5V.n3952 ASIG5V.n3885 0.00796421
R61201 ASIG5V.n4029 ASIG5V.n3953 0.00796421
R61202 ASIG5V.n3954 ASIG5V.n3884 0.00796421
R61203 ASIG5V.n4028 ASIG5V.n3955 0.00796421
R61204 ASIG5V.n3956 ASIG5V.n3883 0.00796421
R61205 ASIG5V.n4027 ASIG5V.n3957 0.00796421
R61206 ASIG5V.n3958 ASIG5V.n3882 0.00796421
R61207 ASIG5V.n4026 ASIG5V.n3959 0.00796421
R61208 ASIG5V.n3960 ASIG5V.n3881 0.00796421
R61209 ASIG5V.n4025 ASIG5V.n3961 0.00796421
R61210 ASIG5V.n3962 ASIG5V.n3880 0.00796421
R61211 ASIG5V.n4024 ASIG5V.n3963 0.00796421
R61212 ASIG5V.n3964 ASIG5V.n3879 0.00796421
R61213 ASIG5V.n4023 ASIG5V.n3965 0.00796421
R61214 ASIG5V.n3966 ASIG5V.n3878 0.00796421
R61215 ASIG5V.n4022 ASIG5V.n3967 0.00796421
R61216 ASIG5V.n3968 ASIG5V.n3877 0.00796421
R61217 ASIG5V.n4021 ASIG5V.n3969 0.00796421
R61218 ASIG5V.n3970 ASIG5V.n3876 0.00796421
R61219 ASIG5V.n4020 ASIG5V.n3971 0.00796421
R61220 ASIG5V.n3972 ASIG5V.n3875 0.00796421
R61221 ASIG5V.n4019 ASIG5V.n3973 0.00796421
R61222 ASIG5V.n3974 ASIG5V.n3874 0.00796421
R61223 ASIG5V.n4018 ASIG5V.n3975 0.00796421
R61224 ASIG5V.n3976 ASIG5V.n3873 0.00796421
R61225 ASIG5V.n4017 ASIG5V.n3977 0.00796421
R61226 ASIG5V.n3978 ASIG5V.n3872 0.00796421
R61227 ASIG5V.n4016 ASIG5V.n3979 0.00796421
R61228 ASIG5V.n3980 ASIG5V.n3871 0.00796421
R61229 ASIG5V.n4015 ASIG5V.n3981 0.00796421
R61230 ASIG5V.n3982 ASIG5V.n3870 0.00796421
R61231 ASIG5V.n4014 ASIG5V.n3983 0.00796421
R61232 ASIG5V.n3984 ASIG5V.n3869 0.00796421
R61233 ASIG5V.n4013 ASIG5V.n3985 0.00796421
R61234 ASIG5V.n3986 ASIG5V.n3868 0.00796421
R61235 ASIG5V.n4012 ASIG5V.n3987 0.00796421
R61236 ASIG5V.n3988 ASIG5V.n3867 0.00796421
R61237 ASIG5V.n4011 ASIG5V.n3989 0.00796421
R61238 ASIG5V.n3990 ASIG5V.n3866 0.00796421
R61239 ASIG5V.n4010 ASIG5V.n3991 0.00796421
R61240 ASIG5V.n3992 ASIG5V.n3865 0.00796421
R61241 ASIG5V.n4009 ASIG5V.n3993 0.00796421
R61242 ASIG5V.n3994 ASIG5V.n3864 0.00796421
R61243 ASIG5V.n4008 ASIG5V.n3995 0.00796421
R61244 ASIG5V.n3996 ASIG5V.n3863 0.00796421
R61245 ASIG5V.n4007 ASIG5V.n3997 0.00796421
R61246 ASIG5V.n3998 ASIG5V.n3862 0.00796421
R61247 ASIG5V.n4006 ASIG5V.n3999 0.00796421
R61248 ASIG5V.n4000 ASIG5V.n3861 0.00796421
R61249 ASIG5V.n4005 ASIG5V.n4001 0.00796421
R61250 ASIG5V.n4002 ASIG5V.n3860 0.00796421
R61251 ASIG5V.n4004 ASIG5V.n4003 0.00796421
R61252 ASIG5V.n3907 ASIG5V.n3859 0.00796421
R61253 ASIG5V.n12294 ASIG5V.n859 0.007925
R61254 ASIG5V.n11756 ASIG5V.n11755 0.007925
R61255 ASIG5V.n10710 ASIG5V.n10705 0.00784763
R61256 ASIG5V.n3852 ASIG5V.n3843 0.00784763
R61257 ASIG5V.n8580 ASIG5V.n54 0.00774832
R61258 ASIG5V.n11773 ASIG5V.n2567 0.00774832
R61259 ASIG5V.n8579 ASIG5V.n163 0.00774832
R61260 ASIG5V.n11774 ASIG5V.n2565 0.00774832
R61261 ASIG5V.n7234 ASIG5V.n6540 0.00753759
R61262 ASIG5V.n10925 ASIG5V.n10466 0.00753759
R61263 ASIG5V.n12534 ASIG5V.n6 0.007475
R61264 ASIG5V.n11176 ASIG5V.n10369 0.007475
R61265 ASIG5V.n5554 ASIG5V.n5463 0.00737773
R61266 ASIG5V.n9413 ASIG5V.n5558 0.00737773
R61267 ASIG5V.n4797 ASIG5V.n3279 0.0072651
R61268 ASIG5V.n7968 ASIG5V.n5508 0.0072651
R61269 ASIG5V.n4796 ASIG5V.n3280 0.0072651
R61270 ASIG5V.n7969 ASIG5V.n7716 0.0072651
R61271 ASIG5V.n10709 ASIG5V.n10693 0.0071375
R61272 ASIG5V.n4264 ASIG5V.n4263 0.0071375
R61273 ASIG5V.n4249 ASIG5V.n4248 0.007025
R61274 ASIG5V.n5068 ASIG5V.n3175 0.007025
R61275 ASIG5V.n7339 ASIG5V.n1316 0.00699624
R61276 ASIG5V.n1830 ASIG5V.n1322 0.00699624
R61277 ASIG5V.n572 ASIG5V.n519 0.00698472
R61278 ASIG5V.n11753 ASIG5V.n2905 0.00698472
R61279 ASIG5V.n862 ASIG5V.n861 0.00698472
R61280 ASIG5V.n11754 ASIG5V.n2908 0.00698472
R61281 ASIG5V.n7236 ASIG5V.n6543 0.00678188
R61282 ASIG5V.n10480 ASIG5V.n10479 0.00678188
R61283 ASIG5V.n7235 ASIG5V.n6541 0.00678188
R61284 ASIG5V.n10478 ASIG5V.n10468 0.00678188
R61285 ASIG5V.n12536 ASIG5V.n2 0.0065917
R61286 ASIG5V.n11174 ASIG5V.n10372 0.0065917
R61287 ASIG5V.n12535 ASIG5V.n4 0.0065917
R61288 ASIG5V.n11175 ASIG5V.n10370 0.0065917
R61289 ASIG5V.n6535 ASIG5V.n6533 0.00645489
R61290 ASIG5V.n8902 ASIG5V.n8901 0.00645489
R61291 ASIG5V.n1320 ASIG5V.n1319 0.00629866
R61292 ASIG5V.n1832 ASIG5V.n1325 0.00629866
R61293 ASIG5V.n12019 ASIG5V.n1317 0.00629866
R61294 ASIG5V.n1831 ASIG5V.n1323 0.00629866
R61295 ASIG5V.n10913 ASIG5V.n10490 0.0062375
R61296 ASIG5V.n10912 ASIG5V.n10491 0.0062375
R61297 ASIG5V.n4251 ASIG5V.n4247 0.0062375
R61298 ASIG5V.n4253 ASIG5V.n3909 0.0062375
R61299 ASIG5V.n4253 ASIG5V.n3839 0.00619869
R61300 ASIG5V.n5066 ASIG5V.n3177 0.00619869
R61301 ASIG5V.n4251 ASIG5V.n4250 0.00619869
R61302 ASIG5V.n5067 ASIG5V.n3176 0.00619869
R61303 ASIG5V.n4584 ASIG5V.n3777 0.00591353
R61304 ASIG5V.n9402 ASIG5V.n5908 0.00591353
R61305 ASIG5V.n6538 ASIG5V.n6430 0.00581544
R61306 ASIG5V.n8927 ASIG5V.n6536 0.00581544
R61307 ASIG5V.n4781 ASIG5V.n4780 0.005675
R61308 ASIG5V.n2561 ASIG5V.n2560 0.00537218
R61309 ASIG5V.n4579 ASIG5V.n3672 0.00533221
R61310 ASIG5V.n9404 ASIG5V.n5569 0.00533221
R61311 ASIG5V.n4581 ASIG5V.n4580 0.00533221
R61312 ASIG5V.n9403 ASIG5V.n5571 0.00533221
R61313 ASIG5V.n8909 ASIG5V.n6887 0.005225
R61314 ASIG5V.n4778 ASIG5V.n3628 0.00501965
R61315 ASIG5V.n4779 ASIG5V.n3626 0.00501965
R61316 ASIG5V.n12325 ASIG5V.n165 0.00484899
R61317 ASIG5V.n2558 ASIG5V.n2220 0.00484899
R61318 ASIG5V.n12326 ASIG5V.n167 0.00484899
R61319 ASIG5V.n2559 ASIG5V.n2219 0.00484899
R61320 ASIG5V.n8587 ASIG5V.n8576 0.00483083
R61321 ASIG5V.n9953 ASIG5V.n2564 0.00483083
R61322 ASIG5V.n11500 ASIG5V.n3002 0.00483083
R61323 ASIG5V.n12273 ASIG5V.n12272 0.004775
R61324 ASIG5V.n11787 ASIG5V.n11786 0.004775
R61325 ASIG5V.n8907 ASIG5V.n6890 0.00462664
R61326 ASIG5V.n8908 ASIG5V.n6888 0.00462664
R61327 ASIG5V.n8574 ASIG5V.n8320 0.00436577
R61328 ASIG5V.n9960 ASIG5V.n9959 0.00436577
R61329 ASIG5V.n8575 ASIG5V.n8321 0.00436577
R61330 ASIG5V.n11502 ASIG5V.n11501 0.00436577
R61331 ASIG5V.n9388 ASIG5V.n6258 0.004325
R61332 ASIG5V.n4812 ASIG5V.n3267 0.00428947
R61333 ASIG5V.n9436 ASIG5V.n5120 0.00428947
R61334 ASIG5V.n12328 ASIG5V.n12327 0.00428947
R61335 ASIG5V.n12270 ASIG5V.n1224 0.00423362
R61336 ASIG5V.n2210 ASIG5V.n1851 0.00423362
R61337 ASIG5V.n12271 ASIG5V.n1222 0.00423362
R61338 ASIG5V.n2208 ASIG5V.n1853 0.00423362
R61339 ASIG5V.n4811 ASIG5V.n4810 0.00388255
R61340 ASIG5V.n9434 ASIG5V.n5122 0.00388255
R61341 ASIG5V.n4814 ASIG5V.n4813 0.00388255
R61342 ASIG5V.n9435 ASIG5V.n5121 0.00388255
R61343 ASIG5V.n6250 ASIG5V.n6000 0.00384061
R61344 ASIG5V.n9390 ASIG5V.n9389 0.00384061
R61345 ASIG5V.n9190 ASIG5V.n6416 0.00374812
R61346 ASIG5V.n8902 ASIG5V.n7244 0.00374812
R61347 ASIG5V.n11187 ASIG5V.n10022 0.00374812
R61348 ASIG5V.n8904 ASIG5V.n6893 0.00339933
R61349 ASIG5V.n11185 ASIG5V.n10024 0.00339933
R61350 ASIG5V.n8903 ASIG5V.n6895 0.00339933
R61351 ASIG5V.n11186 ASIG5V.n10023 0.00339933
R61352 ASIG5V.n12284 ASIG5V.n12283 0.00320677
R61353 ASIG5V.n11806 ASIG5V.n11805 0.00320677
R61354 ASIG5V.n873 ASIG5V.n867 0.00291611
R61355 ASIG5V.n11803 ASIG5V.n1719 0.00291611
R61356 ASIG5V.n871 ASIG5V.n868 0.00291611
R61357 ASIG5V.n11804 ASIG5V.n1836 0.00291611
R61358 ASIG5V.n9748 ASIG5V.n9747 0.00266541
R61359 ASIG5V.n9191 ASIG5V.n6415 0.00266541
R61360 ASIG5V.n10706 ASIG5V.n10694 0.0026375
R61361 ASIG5V.n10700 ASIG5V.n10699 0.0026375
R61362 ASIG5V.n4262 ASIG5V.n3842 0.0026375
R61363 ASIG5V.n4261 ASIG5V.n3841 0.0026375
R61364 ASIG5V.n9409 ASIG5V.n5563 0.002525
R61365 ASIG5V.n6426 ASIG5V.n6308 0.00243289
R61366 ASIG5V.n6428 ASIG5V.n6427 0.00243289
R61367 ASIG5V.n9407 ASIG5V.n5566 0.00226856
R61368 ASIG5V.n9408 ASIG5V.n5564 0.00226856
R61369 ASIG5V.n4573 ASIG5V.n4572 0.00212406
R61370 ASIG5V.n6420 ASIG5V.n5909 0.00212406
R61371 ASIG5V.n11799 ASIG5V.n11798 0.00212406
R61372 ASIG5V.n1219 ASIG5V.n1218 0.002075
R61373 ASIG5V.n11764 ASIG5V.n11763 0.002075
R61374 ASIG5V.n4570 ASIG5V.n3779 0.00194966
R61375 ASIG5V.n6418 ASIG5V.n5911 0.00194966
R61376 ASIG5V.n4571 ASIG5V.n3782 0.00194966
R61377 ASIG5V.n6419 ASIG5V.n5910 0.00194966
R61378 ASIG5V.n879 ASIG5V.n864 0.00187555
R61379 ASIG5V.n11761 ASIG5V.n2613 0.00187555
R61380 ASIG5V.n1217 ASIG5V.n881 0.00187555
R61381 ASIG5V.n11762 ASIG5V.n2903 0.00187555
R61382 ASIG5V.n8887 ASIG5V.n8274 0.001625
R61383 ASIG5V.n12329 ASIG5V.n12328 0.00158271
R61384 ASIG5V.n12306 ASIG5V.n12305 0.00158271
R61385 ASIG5V.n7340 ASIG5V.n7339 0.00158271
R61386 ASIG5V.n11797 ASIG5V.n11796 0.00158271
R61387 ASIG5V.n8266 ASIG5V.n8260 0.00148253
R61388 ASIG5V.n8889 ASIG5V.n8888 0.00148253
R61389 ASIG5V.n12303 ASIG5V.n522 0.00146644
R61390 ASIG5V.n1846 ASIG5V.n1838 0.00146644
R61391 ASIG5V.n12304 ASIG5V.n523 0.00146644
R61392 ASIG5V.n1844 ASIG5V.n1840 0.00146644
R61393 ASIG5V.n10704 ASIG5V.n10696 0.00128471
R61394 ASIG5V.n10696 ASIG5V.n10496 0.00128471
R61395 ASIG5V.n4802 ASIG5V.n3273 0.001175
R61396 ASIG5V.n4800 ASIG5V.n3275 0.00108952
R61397 ASIG5V.n4801 ASIG5V.n3274 0.00108952
R61398 ASIG5V.n4260 ASIG5V.n3851 0.00106946
R61399 ASIG5V.n7963 ASIG5V.n5464 0.00106946
R61400 ASIG5V.n6544 ASIG5V.n6488 0.00106946
R61401 ASIG5V.n10472 ASIG5V.n10471 0.00106946
R61402 ASIG5V.n3781 ASIG5V.n3780 0.00106487
R61403 ASIG5V.n11792 ASIG5V.n11791 0.00106487
R61404 ASIG5V.n12289 ASIG5V.n865 0.0010465
R61405 ASIG5V.n7982 ASIG5V.n7714 0.00104135
R61406 ASIG5V.n8569 ASIG5V.n8168 0.00104135
R61407 ASIG5V.n10021 ASIG5V.n9961 0.00104135
R61408 ASIG5V.n8920 ASIG5V.n6545 0.00103731
R61409 ASIG5V.n508 ASIG5V.n52 0.00103731
R61410 ASIG5V.n4051 ASIG5V.n3848 0.00103272
R61411 ASIG5V.n3858 ASIG5V.n3849 0.00103272
R61412 ASIG5V.n3855 ASIG5V.n3847 0.00103272
R61413 ASIG5V.n3857 ASIG5V.n3850 0.00103272
R61414 ASIG5V.n8268 ASIG5V.n8171 0.00102813
R61415 ASIG5V.n12525 ASIG5V.n98 0.00102813
R61416 ASIG5V.n9177 ASIG5V.n6445 0.00101894
R61417 ASIG5V.n513 ASIG5V.n166 0.00101894
R61418 ASIG5V.n6252 ASIG5V.n5912 0.00100976
R61419 ASIG5V.n12011 ASIG5V.n1370 0.00100517
R61420 ASIG5V.n1675 ASIG5V.n1674 0.00100057
R61421 ASIG5V.n4807 ASIG5V.n3270 0.000991389
R61422 ASIG5V.n9420 ASIG5V.n9419 0.000991389
R61423 ASIG5V.n2907 ASIG5V.n2906 0.000991389
R61424 ASIG5V.n8215 ASIG5V.n8170 0.000983221
R61425 ASIG5V.n10017 ASIG5V.n9964 0.000983221
R61426 ASIG5V.n8324 ASIG5V.n8169 0.000983221
R61427 ASIG5V.n10019 ASIG5V.n9962 0.000983221
R61428 ASIG5V.n9744 ASIG5V.n3169 0.000982204
R61429 ASIG5V.n11495 ASIG5V.n9965 0.000982204
R61430 ASIG5V.n9433 ASIG5V.n9432 0.000977612
R61431 ASIG5V.n5511 ASIG5V.n5510 0.00097302
R61432 ASIG5V.n1328 ASIG5V.n1327 0.00097302
R61433 ASIG5V.n2958 ASIG5V.n2913 0.00097302
R61434 ASIG5V.n6264 ASIG5V.n6263 0.000963835
R61435 ASIG5V.n11163 ASIG5V.n10423 0.000959242
R61436 ASIG5V.n11173 ASIG5V.n11172 0.000959242
R61437 ASIG5V.n6590 ASIG5V.n6587 0.00095465
R61438 ASIG5V.n12529 ASIG5V.n10 0.00095465
R61439 ASIG5V.n4777 ASIG5V.n4776 0.000945465
R61440 ASIG5V.n8277 ASIG5V.n8276 0.000945465
R61441 ASIG5V.n4772 ASIG5V.n3674 0.000940873
R61442 ASIG5V.n9186 ASIG5V.n9185 0.00093628
R61443 ASIG5V.n12324 ASIG5V.n173 0.00093628
R61444 ASIG5V.n12008 ASIG5V.n1415 0.00093628
R61445 ASIG5V.n12278 ASIG5V.n878 0.000927095
R61446 ASIG5V.n11184 ASIG5V.n11183 0.000922503
R61447 ASIG5V.n10911 ASIG5V.n10546 0.000922503
R61448 ASIG5V.n10697 ASIG5V.n10492 0.000922503
R61449 ASIG5V.n10701 ASIG5V.n10495 0.000922503
R61450 ASIG5V.n10712 ASIG5V.n10493 0.000922503
R61451 ASIG5V.n3223 ASIG5V.n3178 0.00091791
R61452 ASIG5V.n4787 ASIG5V.n3620 0.000908726
R61453 ASIG5V.n2556 ASIG5V.n2555 0.000908726
R61454 ASIG5V.n11782 ASIG5V.n11781 0.000908726
R61455 ASIG5V.n11997 ASIG5V.n1717 0.000904133
R61456 ASIG5V.n2221 ASIG5V.n1849 0.000904133
R61457 ASIG5V.n5170 ASIG5V.n5169 0.000894948
R61458 ASIG5V.n7976 ASIG5V.n5553 0.000890356
R61459 ASIG5V.n1326 ASIG5V.n1269 0.000890356
R61460 ASIG5V.n11751 ASIG5V.n2956 0.000890356
R61461 ASIG5V.n10920 ASIG5V.n10482 0.000890356
R61462 ASIG5V.n2199 ASIG5V.n2198 0.000876579
R61463 ASIG5V.n4569 ASIG5V.n4568 0.000871986
R61464 ASIG5V.n9396 ASIG5V.n5954 0.000871986
R61465 ASIG5V.n7238 ASIG5V.n6632 0.000871986
R61466 ASIG5V.n8583 ASIG5V.n8582 0.000871986
R61467 ASIG5V.n877 ASIG5V.n876 0.000862801
R61468 ASIG5V.n9973 ASIG5V.n9966 0.000858209
R61469 ASIG5V.n6431 ASIG5V.n6352 0.000853617
R61470 ASIG5V.n520 ASIG5V.n216 0.000853617
R61471 ASIG5V.n11771 ASIG5V.n2612 0.000844432
R61472 ASIG5V.n10703 ASIG5V.n10483 0.000844432
R61473 ASIG5V.n12288 ASIG5V.n866 0.000839839
R61474 ASIG5V.n10356 ASIG5V.n10076 0.000839839
R61475 ASIG5V.n4268 ASIG5V.n3840 0.000835247
R61476 ASIG5V.n5064 ASIG5V.n3221 0.000835247
R61477 ASIG5V.n9441 ASIG5V.n5117 0.000835247
R61478 ASIG5V.n11192 ASIG5V.n10016 0.000835247
R61479 ASIG5V.n4786 ASIG5V.n3276 0.000826062
R61480 ASIG5V.n4799 ASIG5V.n3276 0.000826062
R61481 ASIG5V.n3278 ASIG5V.n3277 0.000826062
R61482 ASIG5V.n2615 ASIG5V.n2569 0.000826062
R61483 ASIG5V.n8895 ASIG5V.n8213 0.00082147
R61484 ASIG5V.n11994 ASIG5V.n1763 0.00082147
R61485 ASIG5V.n4556 ASIG5V.n4268 0.000816877
R61486 ASIG5V.n1861 ASIG5V.n1763 0.000816877
R61487 ASIG5V.n7978 ASIG5V.n7977 0.000807692
R61488 ASIG5V.n12269 ASIG5V.n1226 0.000807692
R61489 ASIG5V.n2616 ASIG5V.n2213 0.000807692
R61490 ASIG5V.n10919 ASIG5V.n10483 0.000807692
R61491 ASIG5V.n5074 ASIG5V.n3170 0.0008031
R61492 ASIG5V.n12311 ASIG5V.n520 0.000798507
R61493 ASIG5V.n1864 ASIG5V.n1839 0.000793915
R61494 ASIG5V.n4555 ASIG5V.n4554 0.000789323
R61495 ASIG5V.n9393 ASIG5V.n5999 0.000789323
R61496 ASIG5V.n7240 ASIG5V.n7239 0.000789323
R61497 ASIG5V.n8892 ASIG5V.n8217 0.000789323
R61498 ASIG5V.n7239 ASIG5V.n7238 0.000780138
R61499 ASIG5V.n11485 ASIG5V.n11192 0.000775545
R61500 ASIG5V.n6310 ASIG5V.n6306 0.000770953
R61501 ASIG5V.n12311 ASIG5V.n12310 0.000770953
R61502 ASIG5V.n12302 ASIG5V.n12301 0.000770953
R61503 ASIG5V.n7977 ASIG5V.n7976 0.000761768
R61504 ASIG5V.n9406 ASIG5V.n5567 0.000761768
R61505 ASIG5V.n6253 ASIG5V.n5568 0.000761768
R61506 ASIG5V.n10920 ASIG5V.n10919 0.000761768
R61507 ASIG5V.n9393 ASIG5V.n5957 0.000757176
R61508 ASIG5V.n9382 ASIG5V.n6306 0.000757176
R61509 ASIG5V.n8906 ASIG5V.n6891 0.000757176
R61510 ASIG5V.n8269 ASIG5V.n6892 0.000757176
R61511 ASIG5V.n4556 ASIG5V.n4555 0.000752583
R61512 ASIG5V.n9735 ASIG5V.n5074 0.000752583
R61513 ASIG5V.n1861 ASIG5V.n1839 0.000752583
R61514 ASIG5V.n11486 ASIG5V.n9973 0.000752583
R61515 ASIG5V.n8896 ASIG5V.n8895 0.000747991
R61516 ASIG5V.n4787 ASIG5V.n4786 0.000743398
R61517 ASIG5V.n4799 ASIG5V.n4798 0.000743398
R61518 ASIG5V.n1272 ASIG5V.n1271 0.000743398
R61519 ASIG5V.n12269 ASIG5V.n12268 0.000743398
R61520 ASIG5V.n11781 ASIG5V.n2213 0.000743398
R61521 ASIG5V.n11772 ASIG5V.n2569 0.000743398
R61522 ASIG5V.n8892 ASIG5V.n8259 0.000738806
R61523 ASIG5V.n4260 ASIG5V.n3840 0.000734214
R61524 ASIG5V.n5169 ASIG5V.n5117 0.000734214
R61525 ASIG5V ASIG5V.n0 0.000734214
R61526 ASIG5V.n1721 ASIG5V.n1717 0.000734214
R61527 ASIG5V.n10076 ASIG5V.n10016 0.000734214
R61528 ASIG5V.n5065 ASIG5V.n5064 0.000729621
R61529 ASIG5V.n875 ASIG5V.n866 0.000729621
R61530 ASIG5V.n9406 ASIG5V.n9405 0.000725029
R61531 ASIG5V.n1271 ASIG5V.n878 0.000725029
R61532 ASIG5V.n10704 ASIG5V.n10703 0.000725029
R61533 ASIG5V.n9734 ASIG5V.n9441 0.000720436
R61534 ASIG5V.n9186 ASIG5V.n6431 0.000715844
R61535 ASIG5V.n8906 ASIG5V.n8905 0.000706659
R61536 ASIG5V.n8882 ASIG5V.n8277 0.000706659
R61537 ASIG5V.n9397 ASIG5V.n9396 0.000697474
R61538 ASIG5V.n8582 ASIG5V.n10 0.000697474
R61539 ASIG5V.n528 ASIG5V.n521 0.000692882
R61540 ASIG5V.n12301 ASIG5V.n571 0.000692882
R61541 ASIG5V.n9383 ASIG5V.n6264 0.000688289
R61542 ASIG5V.n8905 ASIG5V.n6892 0.000688289
R61543 ASIG5V.n12310 ASIG5V.n521 0.000688289
R61544 ASIG5V.n12302 ASIG5V.n528 0.000688289
R61545 ASIG5V.n8881 ASIG5V.n0 0.000683697
R61546 ASIG5V.n8882 ASIG5V.n8881 0.000679104
R61547 ASIG5V.n12537 ASIG5V.n1 0.000679104
R61548 ASIG5V.n1327 ASIG5V.n1326 0.000679104
R61549 ASIG5V.n10482 ASIG5V.n10416 0.000679104
R61550 ASIG5V.n9379 ASIG5V.n6352 0.000674512
R61551 ASIG5V.n11752 ASIG5V.n11751 0.000674512
R61552 ASIG5V.n4569 ASIG5V.n3787 0.00066992
R61553 ASIG5V.n9744 ASIG5V.n9743 0.00066992
R61554 ASIG5V.n2200 ASIG5V.n2199 0.00066992
R61555 ASIG5V.n11495 ASIG5V.n11494 0.00066992
R61556 ASIG5V.n9405 ASIG5V.n5568 0.000665327
R61557 ASIG5V.n2557 ASIG5V.n2221 0.000665327
R61558 ASIG5V.n4775 ASIG5V.n3620 0.000660735
R61559 ASIG5V.n3277 ASIG5V.n3270 0.000660735
R61560 ASIG5V.n9416 ASIG5V.n5553 0.000660735
R61561 ASIG5V.n11782 ASIG5V.n2212 0.000660735
R61562 ASIG5V.n2906 ASIG5V.n2612 0.000660735
R61563 ASIG5V.n12324 ASIG5V.n12323 0.000656142
R61564 ASIG5V.n4808 ASIG5V.n3223 0.00065155
R61565 ASIG5V.n9433 ASIG5V.n5123 0.00065155
R61566 ASIG5V.n11998 ASIG5V.n1675 0.00065155
R61567 ASIG5V.n11184 ASIG5V.n10025 0.00065155
R61568 ASIG5V.n12279 ASIG5V.n877 0.000646958
R61569 ASIG5V.n10911 ASIG5V.n10496 0.000646958
R61570 ASIG5V.n10546 ASIG5V.n10492 0.000646958
R61571 ASIG5V.n10697 ASIG5V.n10495 0.000646958
R61572 ASIG5V.n10701 ASIG5V.n10493 0.000646958
R61573 ASIG5V.n10712 ASIG5V.n10494 0.000646958
R61574 ASIG5V.n6253 ASIG5V.n6252 0.000642365
R61575 ASIG5V.n12279 ASIG5V.n12278 0.000642365
R61576 ASIG5V.n12008 ASIG5V.n1373 0.00063318
R61577 ASIG5V.n4772 ASIG5V.n3629 0.000628588
R61578 ASIG5V.n6445 ASIG5V.n6432 0.000628588
R61579 ASIG5V.n9383 ASIG5V.n9382 0.000623995
R61580 ASIG5V.n9379 ASIG5V.n6310 0.000623995
R61581 ASIG5V.n8269 ASIG5V.n8268 0.000623995
R61582 ASIG5V.n8276 ASIG5V.n8259 0.000623995
R61583 ASIG5V.n4554 ASIG5V.n3787 0.000610218
R61584 ASIG5V.n4568 ASIG5V.n3830 0.000610218
R61585 ASIG5V.n8919 ASIG5V.n6587 0.000610218
R61586 ASIG5V.n8916 ASIG5V.n6632 0.000610218
R61587 ASIG5V.n6263 ASIG5V.n5999 0.000605626
R61588 ASIG5V.n7240 ASIG5V.n6891 0.000605626
R61589 ASIG5V.n865 ASIG5V.n571 0.000605626
R61590 ASIG5V.n2200 ASIG5V.n1864 0.000605626
R61591 ASIG5V.n2198 ASIG5V.n1848 0.000605626
R61592 ASIG5V.n8583 ASIG5V.n1 0.000601033
R61593 ASIG5V.n1272 ASIG5V.n1226 0.000601033
R61594 ASIG5V.n9743 ASIG5V.n3170 0.000596441
R61595 ASIG5V.n9735 ASIG5V.n9734 0.000596441
R61596 ASIG5V.n5510 ASIG5V.n5506 0.000596441
R61597 ASIG5V.n12012 ASIG5V.n1328 0.000596441
R61598 ASIG5V.n9957 ASIG5V.n2958 0.000596441
R61599 ASIG5V.n11163 ASIG5V.n10373 0.000596441
R61600 ASIG5V.n11173 ASIG5V.n10373 0.000596441
R61601 ASIG5V.n3830 ASIG5V.n3781 0.000587256
R61602 ASIG5V.n3221 ASIG5V.n3169 0.000587256
R61603 ASIG5V.n8916 ASIG5V.n6590 0.000587256
R61604 ASIG5V.n11792 ASIG5V.n1848 0.000587256
R61605 ASIG5V.n9965 ASIG5V.n2956 0.000587256
R61606 ASIG5V.n4798 ASIG5V.n3278 0.000582664
R61607 ASIG5V.n7978 ASIG5V.n5567 0.000582664
R61608 ASIG5V.n2555 ASIG5V.n2212 0.000582664
R61609 ASIG5V.n4777 ASIG5V.n3629 0.000578071
R61610 ASIG5V.n4808 ASIG5V.n4807 0.000578071
R61611 ASIG5V.n2557 ASIG5V.n2556 0.000578071
R61612 ASIG5V.n9957 ASIG5V.n2907 0.000578071
R61613 ASIG5V.n10356 ASIG5V.n10025 0.000578071
R61614 ASIG5V.n11183 ASIG5V.n10068 0.000578071
R61615 ASIG5V.n12529 ASIG5V.n12528 0.000573479
R61616 ASIG5V.n219 ASIG5V.n166 0.000573479
R61617 ASIG5V.n7963 ASIG5V.n5166 0.000568886
R61618 ASIG5V.n1674 ASIG5V.n1415 0.000568886
R61619 ASIG5V.n10472 ASIG5V.n10068 0.000568886
R61620 ASIG5V.n9419 ASIG5V.n5506 0.000564294
R61621 ASIG5V.n11772 ASIG5V.n11771 0.000564294
R61622 ASIG5V.n9397 ASIG5V.n5912 0.000559702
R61623 ASIG5V.n219 ASIG5V.n173 0.000559702
R61624 ASIG5V.n12323 ASIG5V.n216 0.000559702
R61625 ASIG5V.n876 ASIG5V.n875 0.000559702
R61626 ASIG5V ASIG5V.n12537 0.000555109
R61627 ASIG5V.n513 ASIG5V.n98 0.000550517
R61628 ASIG5V.n12012 ASIG5V.n12011 0.000550517
R61629 ASIG5V.n4776 ASIG5V.n4775 0.000545924
R61630 ASIG5V.n9176 ASIG5V.n6488 0.000545924
R61631 ASIG5V.n8896 ASIG5V.n8171 0.000541332
R61632 ASIG5V.n8217 ASIG5V.n8213 0.000541332
R61633 ASIG5V.n12528 ASIG5V.n52 0.000541332
R61634 ASIG5V.n12525 ASIG5V.n56 0.000541332
R61635 ASIG5V.n11494 ASIG5V.n9966 0.000541332
R61636 ASIG5V.n11486 ASIG5V.n11485 0.000541332
R61637 ASIG5V.n4255 ASIG5V.n3848 0.000536739
R61638 ASIG5V.n4051 ASIG5V.n3849 0.000536739
R61639 ASIG5V.n3858 ASIG5V.n3847 0.000536739
R61640 ASIG5V.n3855 ASIG5V.n3850 0.000536739
R61641 ASIG5V.n3857 ASIG5V.n3851 0.000536739
R61642 ASIG5V.n6545 ASIG5V.n6544 0.000532147
R61643 ASIG5V.n508 ASIG5V.n56 0.000532147
R61644 ASIG5V.n5170 ASIG5V.n5123 0.000522962
R61645 ASIG5V.n9432 ASIG5V.n5166 0.000522962
R61646 ASIG5V.n5957 ASIG5V.n5954 0.000522962
R61647 ASIG5V.n12289 ASIG5V.n12288 0.000522962
R61648 ASIG5V.n9416 ASIG5V.n5511 0.00051837
R61649 ASIG5V.n12268 ASIG5V.n1269 0.00051837
R61650 ASIG5V.n2616 ASIG5V.n2615 0.00051837
R61651 ASIG5V.n9420 ASIG5V.n5464 0.000513777
R61652 ASIG5V.n1373 ASIG5V.n1370 0.000513777
R61653 ASIG5V.n11998 ASIG5V.n11997 0.000513777
R61654 ASIG5V.n11994 ASIG5V.n1721 0.000513777
R61655 ASIG5V.n10471 ASIG5V.n10423 0.000513777
R61656 ASIG5V.n11172 ASIG5V.n10416 0.000513777
R61657 ASIG5V.n3780 ASIG5V.n3674 0.000504592
R61658 ASIG5V.n5065 ASIG5V.n3178 0.000504592
R61659 ASIG5V.n9185 ASIG5V.n6432 0.000504592
R61660 ASIG5V.n9177 ASIG5V.n9176 0.000504592
R61661 ASIG5V.n8920 ASIG5V.n8919 0.000504592
R61662 ASIG5V.n11791 ASIG5V.n1849 0.000504592
R61663 ASIG5V.n11752 ASIG5V.n2913 0.000504592
R61664 VDD.n11 VDD.n10 4.78206
R61665 VDD.n7 VDD.n6 0.4505
R61666 VDD.n4 VDD.n3 0.4505
R61667 VDD.n17 VDD.n16 0.4505
R61668 VDD.n13 VDD.n0 0.4505
R61669 VDD.n10 VDD.n2 0.412128
R61670 VDD.n12 VDD.n11 0.412128
R61671 VDD.n10 VDD.n9 0.411993
R61672 VDD.n14 VDD.n11 0.411993
R61673 VDD.n8 VDD 0.130161
R61674 VDD VDD.n1 0.130161
R61675 VDD VDD.n8 0.101206
R61676 VDD VDD.n1 0.101206
R61677 VDD.n5 VDD.n2 0.0718563
R61678 VDD.n15 VDD.n14 0.0718563
R61679 VDD.n16 VDD.n15 0.0581272
R61680 VDD VDD.n5 0.0569273
R61681 VDD.n5 VDD.n4 0.026764
R61682 VDD.n15 VDD.n0 0.026764
R61683 VDD.n8 VDD.n7 0.0142814
R61684 VDD.n17 VDD.n1 0.0142814
R61685 VDD.n4 VDD 0.00782857
R61686 VDD VDD.n0 0.00782857
R61687 VDD.n9 VDD.n3 0.00467857
R61688 VDD.n13 VDD.n12 0.00467857
R61689 VDD.n3 VDD.n2 0.00429286
R61690 VDD.n14 VDD.n13 0.00429286
R61691 VDD.n9 VDD 0.00365
R61692 VDD.n12 VDD 0.00365
R61693 VDD.n7 VDD 0.0023
R61694 VDD VDD.n17 0.0023
R61695 VDD.n6 VDD 0.0017
R61696 VDD.n6 VDD 0.000671429
R61697 VDD.n16 VDD 0.000671429
R61698 VSS.n7887 VSS.n2467 20126
R61699 VSS.n2467 VSS.n760 20126
R61700 VSS.n7881 VSS.n7271 17859.7
R61701 VSS.n7886 VSS.n7271 17859.7
R61702 VSS.n7887 VSS.n7886 6553.98
R61703 VSS.n7881 VSS.n760 6553.98
R61704 VSS.n9454 VSS.n9453 6266.18
R61705 VSS.n7888 VSS.n761 6258.6
R61706 VSS.n7888 VSS.n7887 5490.26
R61707 VSS.n9454 VSS.n760 5490.26
R61708 VSS.n7251 VSS.n2499 3474.96
R61709 VSS.n7227 VSS.n2499 3474.96
R61710 VSS.n8569 VSS.n1358 2918.55
R61711 VSS.n8827 VSS.n1358 2918.55
R61712 VSS.n9903 VSS.n9 2402.48
R61713 VSS.n7883 VSS.n9 2401.2
R61714 VSS.n9903 VSS.n8 2400.01
R61715 VSS.n7883 VSS.n8 2398.73
R61716 VSS.n9902 VSS.n10 851.766
R61717 VSS.n4073 VSS.n10 851.766
R61718 VSS.n5730 VSS.n4073 851.766
R61719 VSS.n5898 VSS.n5730 851.766
R61720 VSS.n5895 VSS.n5894 851.766
R61721 VSS.n5894 VSS.n5893 851.766
R61722 VSS.n7270 VSS.n2468 851.766
R61723 VSS.n5732 VSS.n2468 794.593
R61724 VSS.n7271 VSS.n7270 496.031
R61725 VSS.n5898 VSS.n5897 425.884
R61726 VSS.n5897 VSS.n5895 425.884
R61727 VSS.n8571 VSS.n1360 167.197
R61728 VSS.n8571 VSS.n8570 167.197
R61729 VSS.n8568 VSS.n1556 167.197
R61730 VSS.n1556 VSS.n1359 167.197
R61731 VSS.n2520 VSS.n2501 130.218
R61732 VSS.n7250 VSS.n2501 130.218
R61733 VSS.n7252 VSS.n2494 130.218
R61734 VSS.n2523 VSS.n2494 130.218
R61735 VSS.n7251 VSS.n2496 127.05
R61736 VSS.n7227 VSS.n2524 127.05
R61737 VSS.n9903 VSS.n9902 96.6714
R61738 VSS.n8058 VSS.n1551 93.6563
R61739 VSS.n8058 VSS.n1357 93.6563
R61740 VSS.n1615 VSS.n1614 93.6563
R61741 VSS.n1615 VSS.n1356 93.6563
R61742 VSS.n8824 VSS.n1361 93.6563
R61743 VSS.n8825 VSS.n8824 93.6563
R61744 VSS.n8569 VSS.n1553 85.7351
R61745 VSS.n8827 VSS.n1354 85.7351
R61746 VSS.n7230 VSS.n2500 75.5231
R61747 VSS.n7230 VSS.n7229 75.5231
R61748 VSS.n7206 VSS.n7205 75.5231
R61749 VSS.n7206 VSS.n2521 75.5231
R61750 VSS.n7174 VSS.n2495 75.5231
R61751 VSS.n7174 VSS.n2525 75.5231
R61752 VSS.n5893 VSS.n5732 57.1732
R61753 VSS.n1360 VSS.n1357 14.4308
R61754 VSS.n1614 VSS.n1555 14.4308
R61755 VSS.n1555 VSS.n1551 14.4308
R61756 VSS.n8570 VSS.n1551 14.4308
R61757 VSS.n8826 VSS.n8825 14.4308
R61758 VSS.n8826 VSS.n1356 14.4308
R61759 VSS.n8828 VSS.n1356 14.4308
R61760 VSS.n8828 VSS.n1357 14.4308
R61761 VSS.n8568 VSS.n1361 14.4308
R61762 VSS.n1554 VSS.n1361 14.4308
R61763 VSS.n1614 VSS.n1554 14.4308
R61764 VSS.n8825 VSS.n1359 14.4308
R61765 VSS.n3820 VSS.n3290 12.7299
R61766 VSS.n9906 VSS.n9905 10.4832
R61767 VSS.n7879 VSS.n7 10.4832
R61768 VSS.n9905 VSS.n9904 7.99992
R61769 VSS.n9904 VSS.n7 7.96398
R61770 VSS.n9453 VSS.n761 7.57947
R61771 VSS.n7885 VSS.n7880 7.08357
R61772 VSS.n7882 VSS.n5 7.08357
R61773 VSS.n7229 VSS.n2520 6.79968
R61774 VSS.n7205 VSS.n2498 6.79968
R61775 VSS.n2500 VSS.n2498 6.79968
R61776 VSS.n7250 VSS.n2500 6.79968
R61777 VSS.n7226 VSS.n2525 6.79968
R61778 VSS.n7226 VSS.n2521 6.79968
R61779 VSS.n7228 VSS.n2521 6.79968
R61780 VSS.n7229 VSS.n7228 6.79968
R61781 VSS.n7252 VSS.n2495 6.79968
R61782 VSS.n2497 VSS.n2495 6.79968
R61783 VSS.n7205 VSS.n2497 6.79968
R61784 VSS.n2525 VSS.n2523 6.79968
R61785 VSS.n7597 VSS.n7596 6.22202
R61786 VSS.n7880 VSS.n7879 6.10967
R61787 VSS.n9906 VSS.n5 6.10909
R61788 VSS.n7884 VSS.n7882 5.11349
R61789 VSS.n7885 VSS.n7884 5.07814
R61790 VSS.n5522 VSS.n5386 4.5005
R61791 VSS.n5525 VSS.n5386 4.5005
R61792 VSS.n5527 VSS.n5386 4.5005
R61793 VSS.n5386 VSS.n5379 4.5005
R61794 VSS.n5522 VSS.n5384 4.5005
R61795 VSS.n5525 VSS.n5384 4.5005
R61796 VSS.n5527 VSS.n5384 4.5005
R61797 VSS.n5384 VSS.n5379 4.5005
R61798 VSS.n5522 VSS.n5387 4.5005
R61799 VSS.n5525 VSS.n5387 4.5005
R61800 VSS.n5527 VSS.n5387 4.5005
R61801 VSS.n5387 VSS.n5379 4.5005
R61802 VSS.n5522 VSS.n5383 4.5005
R61803 VSS.n5525 VSS.n5383 4.5005
R61804 VSS.n5527 VSS.n5383 4.5005
R61805 VSS.n5383 VSS.n5379 4.5005
R61806 VSS.n5522 VSS.n5393 4.5005
R61807 VSS.n5525 VSS.n5393 4.5005
R61808 VSS.n5393 VSS.n5379 4.5005
R61809 VSS.n5525 VSS.n5391 4.5005
R61810 VSS.n5391 VSS.n5379 4.5005
R61811 VSS.n5525 VSS.n5394 4.5005
R61812 VSS.n5394 VSS.n5379 4.5005
R61813 VSS.n5525 VSS.n5390 4.5005
R61814 VSS.n5390 VSS.n5379 4.5005
R61815 VSS.n5525 VSS.n5524 4.5005
R61816 VSS.n5524 VSS.n5379 4.5005
R61817 VSS.n5525 VSS.n5389 4.5005
R61818 VSS.n5389 VSS.n5379 4.5005
R61819 VSS.n5526 VSS.n5525 4.5005
R61820 VSS.n5527 VSS.n5526 4.5005
R61821 VSS.n5526 VSS.n5379 4.5005
R61822 VSS.n358 VSS.n352 4.5005
R61823 VSS.n362 VSS.n352 4.5005
R61824 VSS.n9646 VSS.n352 4.5005
R61825 VSS.n358 VSS.n350 4.5005
R61826 VSS.n9646 VSS.n350 4.5005
R61827 VSS.n358 VSS.n353 4.5005
R61828 VSS.n9646 VSS.n353 4.5005
R61829 VSS.n358 VSS.n349 4.5005
R61830 VSS.n9646 VSS.n349 4.5005
R61831 VSS.n358 VSS.n354 4.5005
R61832 VSS.n9646 VSS.n354 4.5005
R61833 VSS.n358 VSS.n348 4.5005
R61834 VSS.n362 VSS.n348 4.5005
R61835 VSS.n9646 VSS.n348 4.5005
R61836 VSS.n9646 VSS.n355 4.5005
R61837 VSS.n362 VSS.n355 4.5005
R61838 VSS.n358 VSS.n355 4.5005
R61839 VSS.n9644 VSS.n355 4.5005
R61840 VSS.n9646 VSS.n347 4.5005
R61841 VSS.n362 VSS.n347 4.5005
R61842 VSS.n358 VSS.n347 4.5005
R61843 VSS.n9644 VSS.n347 4.5005
R61844 VSS.n9646 VSS.n356 4.5005
R61845 VSS.n362 VSS.n356 4.5005
R61846 VSS.n358 VSS.n356 4.5005
R61847 VSS.n9644 VSS.n356 4.5005
R61848 VSS.n9646 VSS.n346 4.5005
R61849 VSS.n362 VSS.n346 4.5005
R61850 VSS.n358 VSS.n346 4.5005
R61851 VSS.n9644 VSS.n346 4.5005
R61852 VSS.n9646 VSS.n9645 4.5005
R61853 VSS.n9645 VSS.n362 4.5005
R61854 VSS.n9645 VSS.n358 4.5005
R61855 VSS.n9645 VSS.n9644 4.5005
R61856 VSS.n3081 VSS.n3064 4.5005
R61857 VSS.n6715 VSS.n3064 4.5005
R61858 VSS.n6717 VSS.n3064 4.5005
R61859 VSS.n6715 VSS.n3062 4.5005
R61860 VSS.n6717 VSS.n3062 4.5005
R61861 VSS.n6715 VSS.n3065 4.5005
R61862 VSS.n6717 VSS.n3065 4.5005
R61863 VSS.n6715 VSS.n3061 4.5005
R61864 VSS.n6717 VSS.n3061 4.5005
R61865 VSS.n6715 VSS.n3066 4.5005
R61866 VSS.n6717 VSS.n3066 4.5005
R61867 VSS.n6715 VSS.n3060 4.5005
R61868 VSS.n6717 VSS.n3060 4.5005
R61869 VSS.n6715 VSS.n3067 4.5005
R61870 VSS.n6717 VSS.n3067 4.5005
R61871 VSS.n6715 VSS.n3059 4.5005
R61872 VSS.n6717 VSS.n3059 4.5005
R61873 VSS.n6715 VSS.n3068 4.5005
R61874 VSS.n6717 VSS.n3068 4.5005
R61875 VSS.n6715 VSS.n3058 4.5005
R61876 VSS.n6717 VSS.n3058 4.5005
R61877 VSS.n6716 VSS.n6715 4.5005
R61878 VSS.n6716 VSS.n3075 4.5005
R61879 VSS.n6717 VSS.n6716 4.5005
R61880 VSS.n1296 VSS.n1284 4.5005
R61881 VSS.n8861 VSS.n1296 4.5005
R61882 VSS.n8859 VSS.n1296 4.5005
R61883 VSS.n8861 VSS.n1293 4.5005
R61884 VSS.n8859 VSS.n1293 4.5005
R61885 VSS.n8861 VSS.n1299 4.5005
R61886 VSS.n8859 VSS.n1299 4.5005
R61887 VSS.n8861 VSS.n1292 4.5005
R61888 VSS.n8859 VSS.n1292 4.5005
R61889 VSS.n8861 VSS.n1301 4.5005
R61890 VSS.n1301 VSS.n1288 4.5005
R61891 VSS.n8859 VSS.n1301 4.5005
R61892 VSS.n1291 VSS.n1284 4.5005
R61893 VSS.n8861 VSS.n1291 4.5005
R61894 VSS.n1291 VSS.n1288 4.5005
R61895 VSS.n8859 VSS.n1291 4.5005
R61896 VSS.n8859 VSS.n8858 4.5005
R61897 VSS.n8858 VSS.n1288 4.5005
R61898 VSS.n8858 VSS.n1284 4.5005
R61899 VSS.n1308 VSS.n1288 4.5005
R61900 VSS.n8859 VSS.n1308 4.5005
R61901 VSS.n8861 VSS.n1303 4.5005
R61902 VSS.n8859 VSS.n1303 4.5005
R61903 VSS.n8861 VSS.n1289 4.5005
R61904 VSS.n8859 VSS.n1289 4.5005
R61905 VSS.n8861 VSS.n8860 4.5005
R61906 VSS.n8860 VSS.n1288 4.5005
R61907 VSS.n8860 VSS.n8859 4.5005
R61908 VSS.n1352 VSS.n1099 4.5005
R61909 VSS.n1352 VSS.n1101 4.5005
R61910 VSS.n1352 VSS.n1100 4.5005
R61911 VSS.n8040 VSS.n1099 4.5005
R61912 VSS.n8040 VSS.n1101 4.5005
R61913 VSS.n8040 VSS.n1100 4.5005
R61914 VSS.n1137 VSS.n1100 4.5005
R61915 VSS.n1137 VSS.n1101 4.5005
R61916 VSS.n1137 VSS.n1099 4.5005
R61917 VSS.n8962 VSS.n1137 4.5005
R61918 VSS.n8036 VSS.n1100 4.5005
R61919 VSS.n8036 VSS.n1101 4.5005
R61920 VSS.n8036 VSS.n1099 4.5005
R61921 VSS.n1135 VSS.n1099 4.5005
R61922 VSS.n1135 VSS.n1100 4.5005
R61923 VSS.n1133 VSS.n1099 4.5005
R61924 VSS.n1133 VSS.n1100 4.5005
R61925 VSS.n1131 VSS.n1099 4.5005
R61926 VSS.n1131 VSS.n1100 4.5005
R61927 VSS.n1129 VSS.n1099 4.5005
R61928 VSS.n1129 VSS.n1100 4.5005
R61929 VSS.n1127 VSS.n1099 4.5005
R61930 VSS.n1127 VSS.n1100 4.5005
R61931 VSS.n1125 VSS.n1099 4.5005
R61932 VSS.n1125 VSS.n1100 4.5005
R61933 VSS.n1123 VSS.n1099 4.5005
R61934 VSS.n1123 VSS.n1100 4.5005
R61935 VSS.n1121 VSS.n1099 4.5005
R61936 VSS.n1121 VSS.n1100 4.5005
R61937 VSS.n8578 VSS.n1099 4.5005
R61938 VSS.n8578 VSS.n1101 4.5005
R61939 VSS.n8578 VSS.n1100 4.5005
R61940 VSS.n8962 VSS.n1119 4.5005
R61941 VSS.n1119 VSS.n1099 4.5005
R61942 VSS.n1119 VSS.n1101 4.5005
R61943 VSS.n1119 VSS.n1100 4.5005
R61944 VSS.n8962 VSS.n1118 4.5005
R61945 VSS.n1118 VSS.n1099 4.5005
R61946 VSS.n1118 VSS.n1100 4.5005
R61947 VSS.n1116 VSS.n1099 4.5005
R61948 VSS.n1116 VSS.n1100 4.5005
R61949 VSS.n1114 VSS.n1099 4.5005
R61950 VSS.n1114 VSS.n1100 4.5005
R61951 VSS.n1112 VSS.n1099 4.5005
R61952 VSS.n1112 VSS.n1100 4.5005
R61953 VSS.n1110 VSS.n1099 4.5005
R61954 VSS.n1110 VSS.n1100 4.5005
R61955 VSS.n1108 VSS.n1099 4.5005
R61956 VSS.n1108 VSS.n1100 4.5005
R61957 VSS.n1106 VSS.n1099 4.5005
R61958 VSS.n1106 VSS.n1100 4.5005
R61959 VSS.n1104 VSS.n1099 4.5005
R61960 VSS.n1104 VSS.n1100 4.5005
R61961 VSS.n1099 VSS.n1096 4.5005
R61962 VSS.n1101 VSS.n1096 4.5005
R61963 VSS.n1100 VSS.n1096 4.5005
R61964 VSS.n8963 VSS.n1100 4.5005
R61965 VSS.n8963 VSS.n1101 4.5005
R61966 VSS.n8963 VSS.n1099 4.5005
R61967 VSS.n8963 VSS.n8962 4.5005
R61968 VSS.n8971 VSS.n1075 4.5005
R61969 VSS.n9016 VSS.n8971 4.5005
R61970 VSS.n9011 VSS.n8971 4.5005
R61971 VSS.n9011 VSS.n9001 4.5005
R61972 VSS.n9001 VSS.n1075 4.5005
R61973 VSS.n9014 VSS.n8984 4.5005
R61974 VSS.n8984 VSS.n1075 4.5005
R61975 VSS.n9014 VSS.n8987 4.5005
R61976 VSS.n8987 VSS.n1075 4.5005
R61977 VSS.n9014 VSS.n8983 4.5005
R61978 VSS.n8983 VSS.n1075 4.5005
R61979 VSS.n9014 VSS.n8988 4.5005
R61980 VSS.n8988 VSS.n1075 4.5005
R61981 VSS.n9014 VSS.n8982 4.5005
R61982 VSS.n8982 VSS.n1075 4.5005
R61983 VSS.n9014 VSS.n8989 4.5005
R61984 VSS.n8989 VSS.n1075 4.5005
R61985 VSS.n9014 VSS.n8981 4.5005
R61986 VSS.n8981 VSS.n1075 4.5005
R61987 VSS.n9014 VSS.n8990 4.5005
R61988 VSS.n8990 VSS.n1075 4.5005
R61989 VSS.n9014 VSS.n8980 4.5005
R61990 VSS.n8980 VSS.n1075 4.5005
R61991 VSS.n9014 VSS.n8991 4.5005
R61992 VSS.n8991 VSS.n1075 4.5005
R61993 VSS.n9014 VSS.n8979 4.5005
R61994 VSS.n8979 VSS.n1075 4.5005
R61995 VSS.n9014 VSS.n8992 4.5005
R61996 VSS.n8992 VSS.n1075 4.5005
R61997 VSS.n9014 VSS.n8978 4.5005
R61998 VSS.n8978 VSS.n1075 4.5005
R61999 VSS.n9014 VSS.n8993 4.5005
R62000 VSS.n8993 VSS.n1075 4.5005
R62001 VSS.n9014 VSS.n8977 4.5005
R62002 VSS.n8977 VSS.n1075 4.5005
R62003 VSS.n9014 VSS.n8994 4.5005
R62004 VSS.n8994 VSS.n1075 4.5005
R62005 VSS.n9014 VSS.n8976 4.5005
R62006 VSS.n8976 VSS.n1075 4.5005
R62007 VSS.n9014 VSS.n8995 4.5005
R62008 VSS.n8995 VSS.n1075 4.5005
R62009 VSS.n9014 VSS.n8975 4.5005
R62010 VSS.n8975 VSS.n1075 4.5005
R62011 VSS.n9014 VSS.n9013 4.5005
R62012 VSS.n9013 VSS.n1075 4.5005
R62013 VSS.n9014 VSS.n8974 4.5005
R62014 VSS.n8974 VSS.n1075 4.5005
R62015 VSS.n9015 VSS.n9014 4.5005
R62016 VSS.n9016 VSS.n9015 4.5005
R62017 VSS.n9015 VSS.n1075 4.5005
R62018 VSS.n794 VSS.n780 4.5005
R62019 VSS.n794 VSS.n781 4.5005
R62020 VSS.n9367 VSS.n794 4.5005
R62021 VSS.n797 VSS.n781 4.5005
R62022 VSS.n9367 VSS.n797 4.5005
R62023 VSS.n793 VSS.n781 4.5005
R62024 VSS.n9367 VSS.n793 4.5005
R62025 VSS.n799 VSS.n781 4.5005
R62026 VSS.n9367 VSS.n799 4.5005
R62027 VSS.n792 VSS.n781 4.5005
R62028 VSS.n9367 VSS.n792 4.5005
R62029 VSS.n801 VSS.n781 4.5005
R62030 VSS.n9367 VSS.n801 4.5005
R62031 VSS.n791 VSS.n781 4.5005
R62032 VSS.n9367 VSS.n791 4.5005
R62033 VSS.n803 VSS.n781 4.5005
R62034 VSS.n9367 VSS.n803 4.5005
R62035 VSS.n790 VSS.n781 4.5005
R62036 VSS.n9367 VSS.n790 4.5005
R62037 VSS.n805 VSS.n781 4.5005
R62038 VSS.n9367 VSS.n805 4.5005
R62039 VSS.n789 VSS.n781 4.5005
R62040 VSS.n9367 VSS.n789 4.5005
R62041 VSS.n807 VSS.n781 4.5005
R62042 VSS.n9367 VSS.n807 4.5005
R62043 VSS.n788 VSS.n781 4.5005
R62044 VSS.n9367 VSS.n788 4.5005
R62045 VSS.n809 VSS.n781 4.5005
R62046 VSS.n9367 VSS.n809 4.5005
R62047 VSS.n787 VSS.n781 4.5005
R62048 VSS.n9367 VSS.n787 4.5005
R62049 VSS.n811 VSS.n781 4.5005
R62050 VSS.n9367 VSS.n811 4.5005
R62051 VSS.n786 VSS.n781 4.5005
R62052 VSS.n9367 VSS.n786 4.5005
R62053 VSS.n813 VSS.n781 4.5005
R62054 VSS.n9367 VSS.n813 4.5005
R62055 VSS.n785 VSS.n781 4.5005
R62056 VSS.n9367 VSS.n785 4.5005
R62057 VSS.n815 VSS.n781 4.5005
R62058 VSS.n9367 VSS.n815 4.5005
R62059 VSS.n784 VSS.n781 4.5005
R62060 VSS.n9367 VSS.n784 4.5005
R62061 VSS.n9366 VSS.n781 4.5005
R62062 VSS.n9367 VSS.n9366 4.5005
R62063 VSS.n783 VSS.n781 4.5005
R62064 VSS.n9367 VSS.n783 4.5005
R62065 VSS.n9368 VSS.n780 4.5005
R62066 VSS.n9368 VSS.n781 4.5005
R62067 VSS.n9368 VSS.n9367 4.5005
R62068 VSS.n6424 VSS.n3624 4.5005
R62069 VSS.n6426 VSS.n3624 4.5005
R62070 VSS.n3624 VSS.n3622 4.5005
R62071 VSS.n6425 VSS.n6424 4.5005
R62072 VSS.n6426 VSS.n6425 4.5005
R62073 VSS.n6426 VSS.n3598 4.5005
R62074 VSS.n6428 VSS.n3598 4.5005
R62075 VSS.n6426 VSS.n3601 4.5005
R62076 VSS.n6428 VSS.n3601 4.5005
R62077 VSS.n6426 VSS.n3597 4.5005
R62078 VSS.n6428 VSS.n3597 4.5005
R62079 VSS.n6426 VSS.n3602 4.5005
R62080 VSS.n6428 VSS.n3602 4.5005
R62081 VSS.n6426 VSS.n3596 4.5005
R62082 VSS.n6428 VSS.n3596 4.5005
R62083 VSS.n6426 VSS.n3603 4.5005
R62084 VSS.n6428 VSS.n3603 4.5005
R62085 VSS.n6426 VSS.n3595 4.5005
R62086 VSS.n6428 VSS.n3595 4.5005
R62087 VSS.n6426 VSS.n3604 4.5005
R62088 VSS.n6428 VSS.n3604 4.5005
R62089 VSS.n6426 VSS.n3594 4.5005
R62090 VSS.n6428 VSS.n3594 4.5005
R62091 VSS.n6426 VSS.n3605 4.5005
R62092 VSS.n6428 VSS.n3605 4.5005
R62093 VSS.n6426 VSS.n3593 4.5005
R62094 VSS.n6428 VSS.n3593 4.5005
R62095 VSS.n6426 VSS.n3606 4.5005
R62096 VSS.n6428 VSS.n3606 4.5005
R62097 VSS.n6426 VSS.n3592 4.5005
R62098 VSS.n6428 VSS.n3592 4.5005
R62099 VSS.n6426 VSS.n3607 4.5005
R62100 VSS.n6428 VSS.n3607 4.5005
R62101 VSS.n6426 VSS.n3591 4.5005
R62102 VSS.n6428 VSS.n3591 4.5005
R62103 VSS.n6426 VSS.n3608 4.5005
R62104 VSS.n6428 VSS.n3608 4.5005
R62105 VSS.n6426 VSS.n3590 4.5005
R62106 VSS.n6428 VSS.n3590 4.5005
R62107 VSS.n6426 VSS.n3609 4.5005
R62108 VSS.n6428 VSS.n3609 4.5005
R62109 VSS.n6426 VSS.n3589 4.5005
R62110 VSS.n6428 VSS.n3589 4.5005
R62111 VSS.n6426 VSS.n3610 4.5005
R62112 VSS.n6428 VSS.n3610 4.5005
R62113 VSS.n6426 VSS.n3588 4.5005
R62114 VSS.n6428 VSS.n3588 4.5005
R62115 VSS.n6427 VSS.n6426 4.5005
R62116 VSS.n6427 VSS.n3622 4.5005
R62117 VSS.n6428 VSS.n6427 4.5005
R62118 VSS.n6543 VSS.n3290 4.5005
R62119 VSS.n3315 VSS.n3290 4.5005
R62120 VSS.n6545 VSS.n3290 4.5005
R62121 VSS.n6543 VSS.n3292 4.5005
R62122 VSS.n6545 VSS.n3292 4.5005
R62123 VSS.n6543 VSS.n3289 4.5005
R62124 VSS.n6545 VSS.n3289 4.5005
R62125 VSS.n6543 VSS.n3293 4.5005
R62126 VSS.n6545 VSS.n3293 4.5005
R62127 VSS.n6543 VSS.n3288 4.5005
R62128 VSS.n6545 VSS.n3288 4.5005
R62129 VSS.n6543 VSS.n3294 4.5005
R62130 VSS.n6545 VSS.n3294 4.5005
R62131 VSS.n6543 VSS.n3287 4.5005
R62132 VSS.n6545 VSS.n3287 4.5005
R62133 VSS.n6543 VSS.n3295 4.5005
R62134 VSS.n6545 VSS.n3295 4.5005
R62135 VSS.n6543 VSS.n3286 4.5005
R62136 VSS.n6545 VSS.n3286 4.5005
R62137 VSS.n6543 VSS.n3296 4.5005
R62138 VSS.n6545 VSS.n3296 4.5005
R62139 VSS.n6543 VSS.n3285 4.5005
R62140 VSS.n6545 VSS.n3285 4.5005
R62141 VSS.n6543 VSS.n3297 4.5005
R62142 VSS.n6545 VSS.n3297 4.5005
R62143 VSS.n6543 VSS.n3284 4.5005
R62144 VSS.n6545 VSS.n3284 4.5005
R62145 VSS.n6543 VSS.n3298 4.5005
R62146 VSS.n6545 VSS.n3298 4.5005
R62147 VSS.n6543 VSS.n3283 4.5005
R62148 VSS.n6545 VSS.n3283 4.5005
R62149 VSS.n6543 VSS.n3299 4.5005
R62150 VSS.n6545 VSS.n3299 4.5005
R62151 VSS.n6543 VSS.n3282 4.5005
R62152 VSS.n6545 VSS.n3282 4.5005
R62153 VSS.n6543 VSS.n3300 4.5005
R62154 VSS.n6545 VSS.n3300 4.5005
R62155 VSS.n6543 VSS.n3281 4.5005
R62156 VSS.n6545 VSS.n3281 4.5005
R62157 VSS.n6543 VSS.n3301 4.5005
R62158 VSS.n6545 VSS.n3301 4.5005
R62159 VSS.n6543 VSS.n3280 4.5005
R62160 VSS.n6545 VSS.n3280 4.5005
R62161 VSS.n6543 VSS.n3302 4.5005
R62162 VSS.n6545 VSS.n3302 4.5005
R62163 VSS.n6543 VSS.n3279 4.5005
R62164 VSS.n6545 VSS.n3279 4.5005
R62165 VSS.n6544 VSS.n6543 4.5005
R62166 VSS.n6544 VSS.n3315 4.5005
R62167 VSS.n6545 VSS.n6544 4.5005
R62168 VSS.n6938 VSS.n2838 4.5005
R62169 VSS.n6941 VSS.n2838 4.5005
R62170 VSS.n2838 VSS.n2825 4.5005
R62171 VSS.n6941 VSS.n2835 4.5005
R62172 VSS.n2835 VSS.n2825 4.5005
R62173 VSS.n6941 VSS.n2840 4.5005
R62174 VSS.n2840 VSS.n2825 4.5005
R62175 VSS.n6941 VSS.n2834 4.5005
R62176 VSS.n2834 VSS.n2825 4.5005
R62177 VSS.n6941 VSS.n2842 4.5005
R62178 VSS.n2842 VSS.n2825 4.5005
R62179 VSS.n6941 VSS.n2833 4.5005
R62180 VSS.n2833 VSS.n2825 4.5005
R62181 VSS.n6941 VSS.n2844 4.5005
R62182 VSS.n2844 VSS.n2825 4.5005
R62183 VSS.n6941 VSS.n2832 4.5005
R62184 VSS.n2832 VSS.n2825 4.5005
R62185 VSS.n6941 VSS.n2846 4.5005
R62186 VSS.n2846 VSS.n2825 4.5005
R62187 VSS.n6941 VSS.n2831 4.5005
R62188 VSS.n2831 VSS.n2825 4.5005
R62189 VSS.n6941 VSS.n6940 4.5005
R62190 VSS.n6940 VSS.n2830 4.5005
R62191 VSS.n6940 VSS.n2825 4.5005
R62192 VSS.n8330 VSS.n1687 4.5005
R62193 VSS.n1687 VSS.n1686 4.5005
R62194 VSS.n8327 VSS.n1687 4.5005
R62195 VSS.n1698 VSS.n1686 4.5005
R62196 VSS.n8327 VSS.n1698 4.5005
R62197 VSS.n8317 VSS.n1686 4.5005
R62198 VSS.n8327 VSS.n8317 4.5005
R62199 VSS.n1697 VSS.n1686 4.5005
R62200 VSS.n8327 VSS.n1697 4.5005
R62201 VSS.n8318 VSS.n1686 4.5005
R62202 VSS.n8327 VSS.n8318 4.5005
R62203 VSS.n1696 VSS.n1686 4.5005
R62204 VSS.n8327 VSS.n1696 4.5005
R62205 VSS.n8325 VSS.n1686 4.5005
R62206 VSS.n8327 VSS.n8325 4.5005
R62207 VSS.n1695 VSS.n1686 4.5005
R62208 VSS.n8327 VSS.n1695 4.5005
R62209 VSS.n8326 VSS.n1686 4.5005
R62210 VSS.n8327 VSS.n8326 4.5005
R62211 VSS.n8328 VSS.n1686 4.5005
R62212 VSS.n8328 VSS.n8327 4.5005
R62213 VSS.n1692 VSS.n1686 4.5005
R62214 VSS.n8323 VSS.n1692 4.5005
R62215 VSS.n8327 VSS.n1692 4.5005
R62216 VSS.n2269 VSS.n2221 4.5005
R62217 VSS.n2221 VSS.n2174 4.5005
R62218 VSS.n2221 VSS.n2176 4.5005
R62219 VSS.n2219 VSS.n2174 4.5005
R62220 VSS.n2219 VSS.n2176 4.5005
R62221 VSS.n2217 VSS.n2174 4.5005
R62222 VSS.n2217 VSS.n2176 4.5005
R62223 VSS.n2215 VSS.n2174 4.5005
R62224 VSS.n2215 VSS.n2176 4.5005
R62225 VSS.n2213 VSS.n2174 4.5005
R62226 VSS.n2213 VSS.n2176 4.5005
R62227 VSS.n2211 VSS.n2174 4.5005
R62228 VSS.n2211 VSS.n2176 4.5005
R62229 VSS.n2209 VSS.n2174 4.5005
R62230 VSS.n2209 VSS.n2176 4.5005
R62231 VSS.n2207 VSS.n2174 4.5005
R62232 VSS.n2207 VSS.n2176 4.5005
R62233 VSS.n2205 VSS.n2174 4.5005
R62234 VSS.n2205 VSS.n2176 4.5005
R62235 VSS.n2203 VSS.n2174 4.5005
R62236 VSS.n2203 VSS.n2176 4.5005
R62237 VSS.n2201 VSS.n2174 4.5005
R62238 VSS.n2201 VSS.n2176 4.5005
R62239 VSS.n2199 VSS.n2174 4.5005
R62240 VSS.n2199 VSS.n2176 4.5005
R62241 VSS.n2197 VSS.n2174 4.5005
R62242 VSS.n2197 VSS.n2176 4.5005
R62243 VSS.n2195 VSS.n2174 4.5005
R62244 VSS.n2195 VSS.n2176 4.5005
R62245 VSS.n2193 VSS.n2174 4.5005
R62246 VSS.n2193 VSS.n2176 4.5005
R62247 VSS.n2191 VSS.n2174 4.5005
R62248 VSS.n2191 VSS.n2176 4.5005
R62249 VSS.n2189 VSS.n2174 4.5005
R62250 VSS.n2189 VSS.n2176 4.5005
R62251 VSS.n2187 VSS.n2174 4.5005
R62252 VSS.n2187 VSS.n2176 4.5005
R62253 VSS.n2185 VSS.n2174 4.5005
R62254 VSS.n2185 VSS.n2176 4.5005
R62255 VSS.n2183 VSS.n2174 4.5005
R62256 VSS.n2183 VSS.n2176 4.5005
R62257 VSS.n2181 VSS.n2174 4.5005
R62258 VSS.n2181 VSS.n2176 4.5005
R62259 VSS.n2179 VSS.n2174 4.5005
R62260 VSS.n2179 VSS.n2176 4.5005
R62261 VSS.n2174 VSS.n2173 4.5005
R62262 VSS.n2175 VSS.n2173 4.5005
R62263 VSS.n2176 VSS.n2173 4.5005
R62264 VSS.n2270 VSS.n2175 4.5005
R62265 VSS.n2270 VSS.n2176 4.5005
R62266 VSS.n2270 VSS.n2174 4.5005
R62267 VSS.n2270 VSS.n2269 4.5005
R62268 VSS.n2168 VSS.n2154 4.5005
R62269 VSS.n7929 VSS.n2154 4.5005
R62270 VSS.n2154 VSS.n2142 4.5005
R62271 VSS.n7931 VSS.n2154 4.5005
R62272 VSS.n7931 VSS.n2155 4.5005
R62273 VSS.n2155 VSS.n2142 4.5005
R62274 VSS.n2168 VSS.n2155 4.5005
R62275 VSS.n7929 VSS.n2155 4.5005
R62276 VSS.n7931 VSS.n2153 4.5005
R62277 VSS.n2153 VSS.n2142 4.5005
R62278 VSS.n2168 VSS.n2153 4.5005
R62279 VSS.n7929 VSS.n2153 4.5005
R62280 VSS.n7931 VSS.n2156 4.5005
R62281 VSS.n2156 VSS.n2142 4.5005
R62282 VSS.n2168 VSS.n2156 4.5005
R62283 VSS.n7929 VSS.n2156 4.5005
R62284 VSS.n7931 VSS.n2152 4.5005
R62285 VSS.n2152 VSS.n2142 4.5005
R62286 VSS.n2168 VSS.n2152 4.5005
R62287 VSS.n7929 VSS.n2152 4.5005
R62288 VSS.n2168 VSS.n2157 4.5005
R62289 VSS.n7929 VSS.n2157 4.5005
R62290 VSS.n2157 VSS.n2142 4.5005
R62291 VSS.n7931 VSS.n2157 4.5005
R62292 VSS.n2168 VSS.n2151 4.5005
R62293 VSS.n7929 VSS.n2151 4.5005
R62294 VSS.n2151 VSS.n2142 4.5005
R62295 VSS.n7931 VSS.n2151 4.5005
R62296 VSS.n2168 VSS.n2158 4.5005
R62297 VSS.n7929 VSS.n2158 4.5005
R62298 VSS.n2158 VSS.n2142 4.5005
R62299 VSS.n7931 VSS.n2158 4.5005
R62300 VSS.n7931 VSS.n2150 4.5005
R62301 VSS.n2150 VSS.n2142 4.5005
R62302 VSS.n2168 VSS.n2150 4.5005
R62303 VSS.n7929 VSS.n2150 4.5005
R62304 VSS.n7931 VSS.n2159 4.5005
R62305 VSS.n2159 VSS.n2142 4.5005
R62306 VSS.n2168 VSS.n2159 4.5005
R62307 VSS.n7929 VSS.n2159 4.5005
R62308 VSS.n7931 VSS.n2149 4.5005
R62309 VSS.n2149 VSS.n2142 4.5005
R62310 VSS.n2168 VSS.n2149 4.5005
R62311 VSS.n7929 VSS.n2149 4.5005
R62312 VSS.n7931 VSS.n2160 4.5005
R62313 VSS.n2160 VSS.n2142 4.5005
R62314 VSS.n2168 VSS.n2160 4.5005
R62315 VSS.n7929 VSS.n2160 4.5005
R62316 VSS.n2168 VSS.n2148 4.5005
R62317 VSS.n7929 VSS.n2148 4.5005
R62318 VSS.n2148 VSS.n2142 4.5005
R62319 VSS.n7931 VSS.n2148 4.5005
R62320 VSS.n2168 VSS.n2161 4.5005
R62321 VSS.n7929 VSS.n2161 4.5005
R62322 VSS.n2161 VSS.n2142 4.5005
R62323 VSS.n7931 VSS.n2161 4.5005
R62324 VSS.n2168 VSS.n2147 4.5005
R62325 VSS.n7929 VSS.n2147 4.5005
R62326 VSS.n2147 VSS.n2142 4.5005
R62327 VSS.n7931 VSS.n2147 4.5005
R62328 VSS.n7931 VSS.n2162 4.5005
R62329 VSS.n2162 VSS.n2142 4.5005
R62330 VSS.n2168 VSS.n2162 4.5005
R62331 VSS.n7929 VSS.n2162 4.5005
R62332 VSS.n7931 VSS.n2146 4.5005
R62333 VSS.n2146 VSS.n2142 4.5005
R62334 VSS.n2168 VSS.n2146 4.5005
R62335 VSS.n7929 VSS.n2146 4.5005
R62336 VSS.n7931 VSS.n2163 4.5005
R62337 VSS.n2163 VSS.n2142 4.5005
R62338 VSS.n2168 VSS.n2163 4.5005
R62339 VSS.n7929 VSS.n2163 4.5005
R62340 VSS.n2168 VSS.n2145 4.5005
R62341 VSS.n7929 VSS.n2145 4.5005
R62342 VSS.n2145 VSS.n2142 4.5005
R62343 VSS.n7931 VSS.n2145 4.5005
R62344 VSS.n2168 VSS.n2164 4.5005
R62345 VSS.n7929 VSS.n2164 4.5005
R62346 VSS.n2164 VSS.n2142 4.5005
R62347 VSS.n7931 VSS.n2164 4.5005
R62348 VSS.n2168 VSS.n2144 4.5005
R62349 VSS.n7929 VSS.n2144 4.5005
R62350 VSS.n2144 VSS.n2142 4.5005
R62351 VSS.n7931 VSS.n2144 4.5005
R62352 VSS.n2168 VSS.n2165 4.5005
R62353 VSS.n7929 VSS.n2165 4.5005
R62354 VSS.n2165 VSS.n2142 4.5005
R62355 VSS.n7931 VSS.n2165 4.5005
R62356 VSS.n7931 VSS.n2143 4.5005
R62357 VSS.n2143 VSS.n2142 4.5005
R62358 VSS.n2168 VSS.n2143 4.5005
R62359 VSS.n7929 VSS.n2143 4.5005
R62360 VSS.n7931 VSS.n7930 4.5005
R62361 VSS.n7930 VSS.n2142 4.5005
R62362 VSS.n7930 VSS.n2168 4.5005
R62363 VSS.n7930 VSS.n7929 4.5005
R62364 VSS.n8243 VSS.n1850 4.5005
R62365 VSS.n1864 VSS.n1850 4.5005
R62366 VSS.n1865 VSS.n1850 4.5005
R62367 VSS.n8245 VSS.n1850 4.5005
R62368 VSS.n1865 VSS.n1852 4.5005
R62369 VSS.n8245 VSS.n1852 4.5005
R62370 VSS.n1864 VSS.n1852 4.5005
R62371 VSS.n8243 VSS.n1852 4.5005
R62372 VSS.n1865 VSS.n1849 4.5005
R62373 VSS.n8245 VSS.n1849 4.5005
R62374 VSS.n1864 VSS.n1849 4.5005
R62375 VSS.n8243 VSS.n1849 4.5005
R62376 VSS.n1865 VSS.n1853 4.5005
R62377 VSS.n8245 VSS.n1853 4.5005
R62378 VSS.n1864 VSS.n1853 4.5005
R62379 VSS.n8243 VSS.n1853 4.5005
R62380 VSS.n8243 VSS.n1848 4.5005
R62381 VSS.n1864 VSS.n1848 4.5005
R62382 VSS.n1865 VSS.n1848 4.5005
R62383 VSS.n8245 VSS.n1848 4.5005
R62384 VSS.n8243 VSS.n1854 4.5005
R62385 VSS.n1864 VSS.n1854 4.5005
R62386 VSS.n1865 VSS.n1854 4.5005
R62387 VSS.n8245 VSS.n1854 4.5005
R62388 VSS.n8243 VSS.n1847 4.5005
R62389 VSS.n1864 VSS.n1847 4.5005
R62390 VSS.n1865 VSS.n1847 4.5005
R62391 VSS.n8245 VSS.n1847 4.5005
R62392 VSS.n1865 VSS.n1855 4.5005
R62393 VSS.n8245 VSS.n1855 4.5005
R62394 VSS.n1864 VSS.n1855 4.5005
R62395 VSS.n8243 VSS.n1855 4.5005
R62396 VSS.n1865 VSS.n1846 4.5005
R62397 VSS.n8245 VSS.n1846 4.5005
R62398 VSS.n1864 VSS.n1846 4.5005
R62399 VSS.n8243 VSS.n1846 4.5005
R62400 VSS.n1865 VSS.n1856 4.5005
R62401 VSS.n8245 VSS.n1856 4.5005
R62402 VSS.n1864 VSS.n1856 4.5005
R62403 VSS.n8243 VSS.n1856 4.5005
R62404 VSS.n1865 VSS.n1845 4.5005
R62405 VSS.n8245 VSS.n1845 4.5005
R62406 VSS.n1864 VSS.n1845 4.5005
R62407 VSS.n8243 VSS.n1845 4.5005
R62408 VSS.n8243 VSS.n1857 4.5005
R62409 VSS.n1864 VSS.n1857 4.5005
R62410 VSS.n1865 VSS.n1857 4.5005
R62411 VSS.n8245 VSS.n1857 4.5005
R62412 VSS.n8243 VSS.n1844 4.5005
R62413 VSS.n1864 VSS.n1844 4.5005
R62414 VSS.n1865 VSS.n1844 4.5005
R62415 VSS.n8245 VSS.n1844 4.5005
R62416 VSS.n8243 VSS.n1858 4.5005
R62417 VSS.n1864 VSS.n1858 4.5005
R62418 VSS.n1865 VSS.n1858 4.5005
R62419 VSS.n8245 VSS.n1858 4.5005
R62420 VSS.n1865 VSS.n1843 4.5005
R62421 VSS.n8245 VSS.n1843 4.5005
R62422 VSS.n1864 VSS.n1843 4.5005
R62423 VSS.n8243 VSS.n1843 4.5005
R62424 VSS.n1865 VSS.n1859 4.5005
R62425 VSS.n8245 VSS.n1859 4.5005
R62426 VSS.n1864 VSS.n1859 4.5005
R62427 VSS.n8243 VSS.n1859 4.5005
R62428 VSS.n1865 VSS.n1842 4.5005
R62429 VSS.n8245 VSS.n1842 4.5005
R62430 VSS.n1864 VSS.n1842 4.5005
R62431 VSS.n8243 VSS.n1842 4.5005
R62432 VSS.n8243 VSS.n1860 4.5005
R62433 VSS.n1864 VSS.n1860 4.5005
R62434 VSS.n1865 VSS.n1860 4.5005
R62435 VSS.n8245 VSS.n1860 4.5005
R62436 VSS.n8243 VSS.n1841 4.5005
R62437 VSS.n1864 VSS.n1841 4.5005
R62438 VSS.n1865 VSS.n1841 4.5005
R62439 VSS.n8245 VSS.n1841 4.5005
R62440 VSS.n8243 VSS.n1861 4.5005
R62441 VSS.n1864 VSS.n1861 4.5005
R62442 VSS.n1865 VSS.n1861 4.5005
R62443 VSS.n8245 VSS.n1861 4.5005
R62444 VSS.n8243 VSS.n1840 4.5005
R62445 VSS.n1864 VSS.n1840 4.5005
R62446 VSS.n1865 VSS.n1840 4.5005
R62447 VSS.n8245 VSS.n1840 4.5005
R62448 VSS.n1865 VSS.n1862 4.5005
R62449 VSS.n8245 VSS.n1862 4.5005
R62450 VSS.n1864 VSS.n1862 4.5005
R62451 VSS.n8243 VSS.n1862 4.5005
R62452 VSS.n1865 VSS.n1839 4.5005
R62453 VSS.n8245 VSS.n1839 4.5005
R62454 VSS.n1864 VSS.n1839 4.5005
R62455 VSS.n8243 VSS.n1839 4.5005
R62456 VSS.n8244 VSS.n1865 4.5005
R62457 VSS.n8245 VSS.n8244 4.5005
R62458 VSS.n8244 VSS.n1864 4.5005
R62459 VSS.n8244 VSS.n8243 4.5005
R62460 VSS.n6218 VSS.n3888 4.5005
R62461 VSS.n6221 VSS.n3888 4.5005
R62462 VSS.n6218 VSS.n3886 4.5005
R62463 VSS.n6221 VSS.n3886 4.5005
R62464 VSS.n6218 VSS.n3889 4.5005
R62465 VSS.n6221 VSS.n3889 4.5005
R62466 VSS.n6218 VSS.n3885 4.5005
R62467 VSS.n6221 VSS.n3885 4.5005
R62468 VSS.n6221 VSS.n6220 4.5005
R62469 VSS.n6218 VSS.n6217 4.5005
R62470 VSS.n6216 VSS.n6215 4.5005
R62471 VSS.n6215 VSS.n3898 4.5005
R62472 VSS.n6215 VSS.n3902 4.5005
R62473 VSS.n6213 VSS.n3902 4.5005
R62474 VSS.n6215 VSS.n3897 4.5005
R62475 VSS.n6213 VSS.n3897 4.5005
R62476 VSS.n6215 VSS.n3903 4.5005
R62477 VSS.n6213 VSS.n3903 4.5005
R62478 VSS.n6215 VSS.n3896 4.5005
R62479 VSS.n6213 VSS.n3896 4.5005
R62480 VSS.n6215 VSS.n6214 4.5005
R62481 VSS.n6214 VSS.n6213 4.5005
R62482 VSS.n4786 VSS.n4558 4.5005
R62483 VSS.n4558 VSS.n4552 4.5005
R62484 VSS.n4563 VSS.n4558 4.5005
R62485 VSS.n4786 VSS.n4557 4.5005
R62486 VSS.n4557 VSS.n4552 4.5005
R62487 VSS.n4781 VSS.n4552 4.5005
R62488 VSS.n4784 VSS.n4781 4.5005
R62489 VSS.n4575 VSS.n4552 4.5005
R62490 VSS.n4784 VSS.n4575 4.5005
R62491 VSS.n4783 VSS.n4552 4.5005
R62492 VSS.n4784 VSS.n4783 4.5005
R62493 VSS.n4574 VSS.n4552 4.5005
R62494 VSS.n4784 VSS.n4574 4.5005
R62495 VSS.n4786 VSS.n4559 4.5005
R62496 VSS.n4559 VSS.n4552 4.5005
R62497 VSS.n4784 VSS.n4559 4.5005
R62498 VSS.n4786 VSS.n4554 4.5005
R62499 VSS.n4554 VSS.n4552 4.5005
R62500 VSS.n4563 VSS.n4554 4.5005
R62501 VSS.n4784 VSS.n4554 4.5005
R62502 VSS.n4786 VSS.n4560 4.5005
R62503 VSS.n4560 VSS.n4552 4.5005
R62504 VSS.n4563 VSS.n4560 4.5005
R62505 VSS.n4784 VSS.n4560 4.5005
R62506 VSS.n4786 VSS.n4553 4.5005
R62507 VSS.n4553 VSS.n4552 4.5005
R62508 VSS.n4563 VSS.n4553 4.5005
R62509 VSS.n4784 VSS.n4553 4.5005
R62510 VSS.n4786 VSS.n4785 4.5005
R62511 VSS.n4785 VSS.n4552 4.5005
R62512 VSS.n4785 VSS.n4563 4.5005
R62513 VSS.n4785 VSS.n4784 4.5005
R62514 VSS.n9749 VSS.n227 4.5005
R62515 VSS.n9749 VSS.n228 4.5005
R62516 VSS.n9758 VSS.n9749 4.5005
R62517 VSS.n232 VSS.n228 4.5005
R62518 VSS.n9758 VSS.n232 4.5005
R62519 VSS.n9752 VSS.n228 4.5005
R62520 VSS.n9758 VSS.n9752 4.5005
R62521 VSS.n231 VSS.n228 4.5005
R62522 VSS.n9758 VSS.n231 4.5005
R62523 VSS.n9755 VSS.n228 4.5005
R62524 VSS.n9758 VSS.n9755 4.5005
R62525 VSS.n230 VSS.n228 4.5005
R62526 VSS.n9758 VSS.n230 4.5005
R62527 VSS.n9757 VSS.n228 4.5005
R62528 VSS.n9757 VSS.n226 4.5005
R62529 VSS.n9758 VSS.n9757 4.5005
R62530 VSS.n227 VSS.n221 4.5005
R62531 VSS.n228 VSS.n221 4.5005
R62532 VSS.n226 VSS.n221 4.5005
R62533 VSS.n9758 VSS.n221 4.5005
R62534 VSS.n227 VSS.n224 4.5005
R62535 VSS.n228 VSS.n224 4.5005
R62536 VSS.n226 VSS.n224 4.5005
R62537 VSS.n9758 VSS.n224 4.5005
R62538 VSS.n227 VSS.n225 4.5005
R62539 VSS.n228 VSS.n225 4.5005
R62540 VSS.n226 VSS.n225 4.5005
R62541 VSS.n9758 VSS.n225 4.5005
R62542 VSS.n9759 VSS.n227 4.5005
R62543 VSS.n9759 VSS.n228 4.5005
R62544 VSS.n9759 VSS.n226 4.5005
R62545 VSS.n9759 VSS.n9758 4.5005
R62546 VSS.n7153 VSS.n2566 4.5005
R62547 VSS.n2570 VSS.n2569 4.5005
R62548 VSS.n2570 VSS.n2566 4.5005
R62549 VSS.n7156 VSS.n2566 4.5005
R62550 VSS.n7156 VSS.n7155 4.5005
R62551 VSS.n9696 VSS.n9695 4.5005
R62552 VSS.n9695 VSS.n250 4.5005
R62553 VSS.n9695 VSS.n9694 4.5005
R62554 VSS.n262 VSS.n250 4.5005
R62555 VSS.n9694 VSS.n262 4.5005
R62556 VSS.n264 VSS.n250 4.5005
R62557 VSS.n9694 VSS.n264 4.5005
R62558 VSS.n261 VSS.n250 4.5005
R62559 VSS.n9694 VSS.n261 4.5005
R62560 VSS.n265 VSS.n250 4.5005
R62561 VSS.n9694 VSS.n265 4.5005
R62562 VSS.n260 VSS.n250 4.5005
R62563 VSS.n9694 VSS.n260 4.5005
R62564 VSS.n9693 VSS.n250 4.5005
R62565 VSS.n9693 VSS.n269 4.5005
R62566 VSS.n9694 VSS.n9693 4.5005
R62567 VSS.n9696 VSS.n254 4.5005
R62568 VSS.n254 VSS.n250 4.5005
R62569 VSS.n269 VSS.n254 4.5005
R62570 VSS.n9694 VSS.n254 4.5005
R62571 VSS.n9696 VSS.n253 4.5005
R62572 VSS.n253 VSS.n250 4.5005
R62573 VSS.n269 VSS.n253 4.5005
R62574 VSS.n9694 VSS.n253 4.5005
R62575 VSS.n9696 VSS.n252 4.5005
R62576 VSS.n252 VSS.n250 4.5005
R62577 VSS.n269 VSS.n252 4.5005
R62578 VSS.n9694 VSS.n252 4.5005
R62579 VSS.n9696 VSS.n251 4.5005
R62580 VSS.n251 VSS.n250 4.5005
R62581 VSS.n269 VSS.n251 4.5005
R62582 VSS.n9694 VSS.n251 4.5005
R62583 VSS.n288 VSS.n280 4.5005
R62584 VSS.n289 VSS.n280 4.5005
R62585 VSS.n287 VSS.n280 4.5005
R62586 VSS.n9683 VSS.n280 4.5005
R62587 VSS.n9684 VSS.n288 4.5005
R62588 VSS.n9684 VSS.n289 4.5005
R62589 VSS.n9684 VSS.n287 4.5005
R62590 VSS.n9684 VSS.n9683 4.5005
R62591 VSS.n298 VSS.n288 4.5005
R62592 VSS.n298 VSS.n289 4.5005
R62593 VSS.n298 VSS.n287 4.5005
R62594 VSS.n9683 VSS.n298 4.5005
R62595 VSS.n294 VSS.n288 4.5005
R62596 VSS.n294 VSS.n289 4.5005
R62597 VSS.n294 VSS.n287 4.5005
R62598 VSS.n9683 VSS.n294 4.5005
R62599 VSS.n300 VSS.n288 4.5005
R62600 VSS.n300 VSS.n289 4.5005
R62601 VSS.n9683 VSS.n300 4.5005
R62602 VSS.n293 VSS.n289 4.5005
R62603 VSS.n9683 VSS.n293 4.5005
R62604 VSS.n303 VSS.n289 4.5005
R62605 VSS.n9683 VSS.n303 4.5005
R62606 VSS.n292 VSS.n289 4.5005
R62607 VSS.n9683 VSS.n292 4.5005
R62608 VSS.n306 VSS.n289 4.5005
R62609 VSS.n9683 VSS.n306 4.5005
R62610 VSS.n291 VSS.n289 4.5005
R62611 VSS.n9683 VSS.n291 4.5005
R62612 VSS.n9682 VSS.n289 4.5005
R62613 VSS.n9682 VSS.n287 4.5005
R62614 VSS.n9683 VSS.n9682 4.5005
R62615 VSS.n9681 VSS.n309 4.5005
R62616 VSS.n9681 VSS.n310 4.5005
R62617 VSS.n9681 VSS.n9680 4.5005
R62618 VSS.n316 VSS.n310 4.5005
R62619 VSS.n9680 VSS.n316 4.5005
R62620 VSS.n319 VSS.n310 4.5005
R62621 VSS.n9680 VSS.n319 4.5005
R62622 VSS.n315 VSS.n310 4.5005
R62623 VSS.n9680 VSS.n315 4.5005
R62624 VSS.n321 VSS.n310 4.5005
R62625 VSS.n9680 VSS.n321 4.5005
R62626 VSS.n314 VSS.n309 4.5005
R62627 VSS.n314 VSS.n310 4.5005
R62628 VSS.n9680 VSS.n314 4.5005
R62629 VSS.n9680 VSS.n322 4.5005
R62630 VSS.n9678 VSS.n322 4.5005
R62631 VSS.n322 VSS.n310 4.5005
R62632 VSS.n322 VSS.n309 4.5005
R62633 VSS.n9680 VSS.n313 4.5005
R62634 VSS.n9678 VSS.n313 4.5005
R62635 VSS.n313 VSS.n310 4.5005
R62636 VSS.n313 VSS.n309 4.5005
R62637 VSS.n9680 VSS.n323 4.5005
R62638 VSS.n9678 VSS.n323 4.5005
R62639 VSS.n323 VSS.n310 4.5005
R62640 VSS.n323 VSS.n309 4.5005
R62641 VSS.n9680 VSS.n312 4.5005
R62642 VSS.n9678 VSS.n312 4.5005
R62643 VSS.n312 VSS.n310 4.5005
R62644 VSS.n312 VSS.n309 4.5005
R62645 VSS.n9680 VSS.n9679 4.5005
R62646 VSS.n9679 VSS.n9678 4.5005
R62647 VSS.n9679 VSS.n310 4.5005
R62648 VSS.n9679 VSS.n309 4.5005
R62649 VSS.n3550 VSS.n3525 4.5005
R62650 VSS.n6451 VSS.n3525 4.5005
R62651 VSS.n6453 VSS.n3525 4.5005
R62652 VSS.n6451 VSS.n3527 4.5005
R62653 VSS.n6453 VSS.n3527 4.5005
R62654 VSS.n6451 VSS.n3524 4.5005
R62655 VSS.n6453 VSS.n3524 4.5005
R62656 VSS.n6451 VSS.n3528 4.5005
R62657 VSS.n6453 VSS.n3528 4.5005
R62658 VSS.n6451 VSS.n3523 4.5005
R62659 VSS.n6453 VSS.n3523 4.5005
R62660 VSS.n6451 VSS.n3529 4.5005
R62661 VSS.n6453 VSS.n3529 4.5005
R62662 VSS.n6451 VSS.n3522 4.5005
R62663 VSS.n6453 VSS.n3522 4.5005
R62664 VSS.n6451 VSS.n3530 4.5005
R62665 VSS.n6453 VSS.n3530 4.5005
R62666 VSS.n6451 VSS.n3521 4.5005
R62667 VSS.n6453 VSS.n3521 4.5005
R62668 VSS.n6451 VSS.n3531 4.5005
R62669 VSS.n6453 VSS.n3531 4.5005
R62670 VSS.n6451 VSS.n3520 4.5005
R62671 VSS.n6453 VSS.n3520 4.5005
R62672 VSS.n6451 VSS.n3532 4.5005
R62673 VSS.n6453 VSS.n3532 4.5005
R62674 VSS.n6451 VSS.n3519 4.5005
R62675 VSS.n6453 VSS.n3519 4.5005
R62676 VSS.n6451 VSS.n3533 4.5005
R62677 VSS.n6453 VSS.n3533 4.5005
R62678 VSS.n6451 VSS.n3518 4.5005
R62679 VSS.n6453 VSS.n3518 4.5005
R62680 VSS.n6451 VSS.n3534 4.5005
R62681 VSS.n6453 VSS.n3534 4.5005
R62682 VSS.n6451 VSS.n3517 4.5005
R62683 VSS.n6453 VSS.n3517 4.5005
R62684 VSS.n6451 VSS.n3535 4.5005
R62685 VSS.n6453 VSS.n3535 4.5005
R62686 VSS.n6451 VSS.n3516 4.5005
R62687 VSS.n6453 VSS.n3516 4.5005
R62688 VSS.n6451 VSS.n3536 4.5005
R62689 VSS.n6453 VSS.n3536 4.5005
R62690 VSS.n6451 VSS.n3515 4.5005
R62691 VSS.n6453 VSS.n3515 4.5005
R62692 VSS.n6451 VSS.n3537 4.5005
R62693 VSS.n6453 VSS.n3537 4.5005
R62694 VSS.n6451 VSS.n3514 4.5005
R62695 VSS.n6453 VSS.n3514 4.5005
R62696 VSS.n6452 VSS.n3550 4.5005
R62697 VSS.n6452 VSS.n6451 4.5005
R62698 VSS.n6453 VSS.n6452 4.5005
R62699 VSS.n6752 VSS.n2973 4.5005
R62700 VSS.n6752 VSS.n2974 4.5005
R62701 VSS.n6752 VSS.n6751 4.5005
R62702 VSS.n2980 VSS.n2974 4.5005
R62703 VSS.n6751 VSS.n2980 4.5005
R62704 VSS.n2983 VSS.n2974 4.5005
R62705 VSS.n6751 VSS.n2983 4.5005
R62706 VSS.n2979 VSS.n2974 4.5005
R62707 VSS.n6751 VSS.n2979 4.5005
R62708 VSS.n2985 VSS.n2974 4.5005
R62709 VSS.n6751 VSS.n2985 4.5005
R62710 VSS.n2978 VSS.n2974 4.5005
R62711 VSS.n6751 VSS.n2978 4.5005
R62712 VSS.n2987 VSS.n2974 4.5005
R62713 VSS.n6751 VSS.n2987 4.5005
R62714 VSS.n2977 VSS.n2974 4.5005
R62715 VSS.n6751 VSS.n2977 4.5005
R62716 VSS.n2989 VSS.n2974 4.5005
R62717 VSS.n6751 VSS.n2989 4.5005
R62718 VSS.n2976 VSS.n2974 4.5005
R62719 VSS.n6751 VSS.n2976 4.5005
R62720 VSS.n6750 VSS.n2974 4.5005
R62721 VSS.n6750 VSS.n6749 4.5005
R62722 VSS.n6751 VSS.n6750 4.5005
R62723 VSS.n1333 VSS.n1323 4.5005
R62724 VSS.n1333 VSS.n1324 4.5005
R62725 VSS.n8842 VSS.n1333 4.5005
R62726 VSS.n1330 VSS.n1324 4.5005
R62727 VSS.n8842 VSS.n1330 4.5005
R62728 VSS.n1336 VSS.n1324 4.5005
R62729 VSS.n8842 VSS.n1336 4.5005
R62730 VSS.n1329 VSS.n1324 4.5005
R62731 VSS.n8842 VSS.n1329 4.5005
R62732 VSS.n1338 VSS.n1324 4.5005
R62733 VSS.n1338 VSS.n1322 4.5005
R62734 VSS.n8842 VSS.n1338 4.5005
R62735 VSS.n8843 VSS.n1323 4.5005
R62736 VSS.n8843 VSS.n1324 4.5005
R62737 VSS.n8843 VSS.n1322 4.5005
R62738 VSS.n8843 VSS.n8842 4.5005
R62739 VSS.n8842 VSS.n1318 4.5005
R62740 VSS.n1322 VSS.n1318 4.5005
R62741 VSS.n1323 VSS.n1318 4.5005
R62742 VSS.n1328 VSS.n1323 4.5005
R62743 VSS.n8842 VSS.n1328 4.5005
R62744 VSS.n1341 VSS.n1324 4.5005
R62745 VSS.n8842 VSS.n1341 4.5005
R62746 VSS.n1326 VSS.n1324 4.5005
R62747 VSS.n8842 VSS.n1326 4.5005
R62748 VSS.n8841 VSS.n1323 4.5005
R62749 VSS.n8841 VSS.n1324 4.5005
R62750 VSS.n8842 VSS.n8841 4.5005
R62751 VSS.n8806 VSS.n1393 4.5005
R62752 VSS.n8806 VSS.n1394 4.5005
R62753 VSS.n8806 VSS.n8805 4.5005
R62754 VSS.n1408 VSS.n1393 4.5005
R62755 VSS.n1408 VSS.n1394 4.5005
R62756 VSS.n8805 VSS.n1408 4.5005
R62757 VSS.n8805 VSS.n1406 4.5005
R62758 VSS.n8803 VSS.n1406 4.5005
R62759 VSS.n1406 VSS.n1394 4.5005
R62760 VSS.n1406 VSS.n1393 4.5005
R62761 VSS.n8805 VSS.n1410 4.5005
R62762 VSS.n8803 VSS.n1410 4.5005
R62763 VSS.n1410 VSS.n1393 4.5005
R62764 VSS.n1405 VSS.n1393 4.5005
R62765 VSS.n8805 VSS.n1405 4.5005
R62766 VSS.n1412 VSS.n1394 4.5005
R62767 VSS.n8805 VSS.n1412 4.5005
R62768 VSS.n1404 VSS.n1394 4.5005
R62769 VSS.n8805 VSS.n1404 4.5005
R62770 VSS.n1414 VSS.n1394 4.5005
R62771 VSS.n8805 VSS.n1414 4.5005
R62772 VSS.n1403 VSS.n1394 4.5005
R62773 VSS.n8805 VSS.n1403 4.5005
R62774 VSS.n1416 VSS.n1394 4.5005
R62775 VSS.n8805 VSS.n1416 4.5005
R62776 VSS.n1402 VSS.n1394 4.5005
R62777 VSS.n8805 VSS.n1402 4.5005
R62778 VSS.n1418 VSS.n1394 4.5005
R62779 VSS.n8805 VSS.n1418 4.5005
R62780 VSS.n1401 VSS.n1394 4.5005
R62781 VSS.n8803 VSS.n1401 4.5005
R62782 VSS.n8805 VSS.n1401 4.5005
R62783 VSS.n1419 VSS.n1393 4.5005
R62784 VSS.n1419 VSS.n1394 4.5005
R62785 VSS.n8803 VSS.n1419 4.5005
R62786 VSS.n8805 VSS.n1419 4.5005
R62787 VSS.n1400 VSS.n1393 4.5005
R62788 VSS.n1400 VSS.n1394 4.5005
R62789 VSS.n8805 VSS.n1400 4.5005
R62790 VSS.n1421 VSS.n1394 4.5005
R62791 VSS.n8805 VSS.n1421 4.5005
R62792 VSS.n1399 VSS.n1394 4.5005
R62793 VSS.n8805 VSS.n1399 4.5005
R62794 VSS.n1423 VSS.n1394 4.5005
R62795 VSS.n8805 VSS.n1423 4.5005
R62796 VSS.n1398 VSS.n1394 4.5005
R62797 VSS.n8805 VSS.n1398 4.5005
R62798 VSS.n1425 VSS.n1394 4.5005
R62799 VSS.n8805 VSS.n1425 4.5005
R62800 VSS.n1397 VSS.n1394 4.5005
R62801 VSS.n8805 VSS.n1397 4.5005
R62802 VSS.n1427 VSS.n1394 4.5005
R62803 VSS.n8805 VSS.n1427 4.5005
R62804 VSS.n1396 VSS.n1394 4.5005
R62805 VSS.n8803 VSS.n1396 4.5005
R62806 VSS.n8805 VSS.n1396 4.5005
R62807 VSS.n8805 VSS.n8804 4.5005
R62808 VSS.n8804 VSS.n8803 4.5005
R62809 VSS.n8804 VSS.n1394 4.5005
R62810 VSS.n8804 VSS.n1393 4.5005
R62811 VSS.n1032 VSS.n1020 4.5005
R62812 VSS.n9055 VSS.n1032 4.5005
R62813 VSS.n9050 VSS.n1032 4.5005
R62814 VSS.n9050 VSS.n9039 4.5005
R62815 VSS.n9039 VSS.n1020 4.5005
R62816 VSS.n9053 VSS.n1043 4.5005
R62817 VSS.n1043 VSS.n1020 4.5005
R62818 VSS.n9053 VSS.n1046 4.5005
R62819 VSS.n1046 VSS.n1020 4.5005
R62820 VSS.n9053 VSS.n1042 4.5005
R62821 VSS.n1042 VSS.n1020 4.5005
R62822 VSS.n9053 VSS.n1047 4.5005
R62823 VSS.n1047 VSS.n1020 4.5005
R62824 VSS.n9053 VSS.n1041 4.5005
R62825 VSS.n1041 VSS.n1020 4.5005
R62826 VSS.n9053 VSS.n1048 4.5005
R62827 VSS.n1048 VSS.n1020 4.5005
R62828 VSS.n9053 VSS.n1040 4.5005
R62829 VSS.n1040 VSS.n1020 4.5005
R62830 VSS.n9053 VSS.n1049 4.5005
R62831 VSS.n1049 VSS.n1020 4.5005
R62832 VSS.n9053 VSS.n1039 4.5005
R62833 VSS.n1039 VSS.n1020 4.5005
R62834 VSS.n9053 VSS.n1050 4.5005
R62835 VSS.n1050 VSS.n1020 4.5005
R62836 VSS.n9053 VSS.n1038 4.5005
R62837 VSS.n1038 VSS.n1020 4.5005
R62838 VSS.n9053 VSS.n1051 4.5005
R62839 VSS.n1051 VSS.n1020 4.5005
R62840 VSS.n9053 VSS.n1037 4.5005
R62841 VSS.n1037 VSS.n1020 4.5005
R62842 VSS.n9053 VSS.n1052 4.5005
R62843 VSS.n1052 VSS.n1020 4.5005
R62844 VSS.n9053 VSS.n1036 4.5005
R62845 VSS.n1036 VSS.n1020 4.5005
R62846 VSS.n9053 VSS.n1053 4.5005
R62847 VSS.n1053 VSS.n1020 4.5005
R62848 VSS.n9053 VSS.n1035 4.5005
R62849 VSS.n1035 VSS.n1020 4.5005
R62850 VSS.n9053 VSS.n1054 4.5005
R62851 VSS.n1054 VSS.n1020 4.5005
R62852 VSS.n9053 VSS.n1034 4.5005
R62853 VSS.n1034 VSS.n1020 4.5005
R62854 VSS.n9053 VSS.n9052 4.5005
R62855 VSS.n9052 VSS.n1020 4.5005
R62856 VSS.n9053 VSS.n1033 4.5005
R62857 VSS.n1033 VSS.n1020 4.5005
R62858 VSS.n9053 VSS.n843 4.5005
R62859 VSS.n9055 VSS.n843 4.5005
R62860 VSS.n1020 VSS.n843 4.5005
R62861 VSS.n9314 VSS.n9313 4.5005
R62862 VSS.n9313 VSS.n831 4.5005
R62863 VSS.n9313 VSS.n9312 4.5005
R62864 VSS.n9288 VSS.n831 4.5005
R62865 VSS.n9312 VSS.n9288 4.5005
R62866 VSS.n856 VSS.n831 4.5005
R62867 VSS.n9312 VSS.n856 4.5005
R62868 VSS.n9289 VSS.n831 4.5005
R62869 VSS.n9312 VSS.n9289 4.5005
R62870 VSS.n855 VSS.n831 4.5005
R62871 VSS.n9312 VSS.n855 4.5005
R62872 VSS.n9290 VSS.n831 4.5005
R62873 VSS.n9312 VSS.n9290 4.5005
R62874 VSS.n854 VSS.n831 4.5005
R62875 VSS.n9312 VSS.n854 4.5005
R62876 VSS.n9291 VSS.n831 4.5005
R62877 VSS.n9312 VSS.n9291 4.5005
R62878 VSS.n853 VSS.n831 4.5005
R62879 VSS.n9312 VSS.n853 4.5005
R62880 VSS.n9292 VSS.n831 4.5005
R62881 VSS.n9312 VSS.n9292 4.5005
R62882 VSS.n852 VSS.n831 4.5005
R62883 VSS.n9312 VSS.n852 4.5005
R62884 VSS.n9293 VSS.n831 4.5005
R62885 VSS.n9312 VSS.n9293 4.5005
R62886 VSS.n851 VSS.n831 4.5005
R62887 VSS.n9312 VSS.n851 4.5005
R62888 VSS.n9294 VSS.n831 4.5005
R62889 VSS.n9312 VSS.n9294 4.5005
R62890 VSS.n850 VSS.n831 4.5005
R62891 VSS.n9312 VSS.n850 4.5005
R62892 VSS.n9295 VSS.n831 4.5005
R62893 VSS.n9312 VSS.n9295 4.5005
R62894 VSS.n849 VSS.n831 4.5005
R62895 VSS.n9312 VSS.n849 4.5005
R62896 VSS.n9296 VSS.n831 4.5005
R62897 VSS.n9312 VSS.n9296 4.5005
R62898 VSS.n848 VSS.n831 4.5005
R62899 VSS.n9312 VSS.n848 4.5005
R62900 VSS.n9297 VSS.n831 4.5005
R62901 VSS.n9312 VSS.n9297 4.5005
R62902 VSS.n847 VSS.n831 4.5005
R62903 VSS.n9312 VSS.n847 4.5005
R62904 VSS.n9311 VSS.n831 4.5005
R62905 VSS.n9312 VSS.n9311 4.5005
R62906 VSS.n846 VSS.n831 4.5005
R62907 VSS.n9312 VSS.n846 4.5005
R62908 VSS.n9314 VSS.n771 4.5005
R62909 VSS.n831 VSS.n771 4.5005
R62910 VSS.n9312 VSS.n771 4.5005
R62911 VSS.n7101 VSS.n7057 4.5005
R62912 VSS.n7101 VSS.n7055 4.5005
R62913 VSS.n7079 VSS.n7074 4.5005
R62914 VSS.n7079 VSS.n7076 4.5005
R62915 VSS.n7079 VSS.n7078 4.5005
R62916 VSS.n7078 VSS.n2599 4.5005
R62917 VSS.n7002 VSS.n7001 4.5005
R62918 VSS.n6770 VSS.n6769 4.5005
R62919 VSS.n6768 VSS.n2954 4.5005
R62920 VSS.n6774 VSS.n2955 4.5005
R62921 VSS.n6777 VSS.n6775 4.5005
R62922 VSS.n6780 VSS.n6778 4.5005
R62923 VSS.n6783 VSS.n6781 4.5005
R62924 VSS.n6786 VSS.n6784 4.5005
R62925 VSS.n6788 VSS.n6787 4.5005
R62926 VSS.n6792 VSS.n6789 4.5005
R62927 VSS.n6795 VSS.n6793 4.5005
R62928 VSS.n6798 VSS.n6796 4.5005
R62929 VSS.n6800 VSS.n2953 4.5005
R62930 VSS.n6803 VSS.n6802 4.5005
R62931 VSS.n2939 VSS.n2938 4.5005
R62932 VSS.n6837 VSS.n6807 4.5005
R62933 VSS.n6836 VSS.n6808 4.5005
R62934 VSS.n6835 VSS.n6809 4.5005
R62935 VSS.n6812 VSS.n6810 4.5005
R62936 VSS.n6831 VSS.n6813 4.5005
R62937 VSS.n6830 VSS.n6814 4.5005
R62938 VSS.n6829 VSS.n6815 4.5005
R62939 VSS.n6818 VSS.n6816 4.5005
R62940 VSS.n6825 VSS.n6819 4.5005
R62941 VSS.n6824 VSS.n6820 4.5005
R62942 VSS.n6823 VSS.n6821 4.5005
R62943 VSS.n2651 VSS.n2650 4.5005
R62944 VSS.n6767 VSS.n2957 4.5005
R62945 VSS.n5880 VSS.n5733 4.5005
R62946 VSS.n5828 VSS.n5824 4.5005
R62947 VSS.n5830 VSS.n5829 4.5005
R62948 VSS.n5822 VSS.n5821 4.5005
R62949 VSS.n5835 VSS.n5834 4.5005
R62950 VSS.n5836 VSS.n5820 4.5005
R62951 VSS.n5838 VSS.n5837 4.5005
R62952 VSS.n5818 VSS.n5817 4.5005
R62953 VSS.n5843 VSS.n5842 4.5005
R62954 VSS.n5844 VSS.n5816 4.5005
R62955 VSS.n5846 VSS.n5845 4.5005
R62956 VSS.n5814 VSS.n5813 4.5005
R62957 VSS.n5852 VSS.n5851 4.5005
R62958 VSS.n5853 VSS.n5812 4.5005
R62959 VSS.n5855 VSS.n5854 4.5005
R62960 VSS.n5856 VSS.n5810 4.5005
R62961 VSS.n5860 VSS.n5859 4.5005
R62962 VSS.n5861 VSS.n5809 4.5005
R62963 VSS.n5863 VSS.n5862 4.5005
R62964 VSS.n5807 VSS.n5806 4.5005
R62965 VSS.n5868 VSS.n5867 4.5005
R62966 VSS.n5869 VSS.n5805 4.5005
R62967 VSS.n5871 VSS.n5870 4.5005
R62968 VSS.n5803 VSS.n5802 4.5005
R62969 VSS.n5876 VSS.n5875 4.5005
R62970 VSS.n5877 VSS.n5801 4.5005
R62971 VSS.n5882 VSS.n5881 4.5005
R62972 VSS.n5827 VSS.n5826 4.5005
R62973 VSS.n6613 VSS.n6612 4.5005
R62974 VSS.n3795 VSS.n3722 4.5005
R62975 VSS.n3794 VSS.n3723 4.5005
R62976 VSS.n3792 VSS.n3724 4.5005
R62977 VSS.n3790 VSS.n3725 4.5005
R62978 VSS.n3788 VSS.n3726 4.5005
R62979 VSS.n3786 VSS.n3727 4.5005
R62980 VSS.n3784 VSS.n3728 4.5005
R62981 VSS.n3782 VSS.n3729 4.5005
R62982 VSS.n3779 VSS.n3730 4.5005
R62983 VSS.n3778 VSS.n3731 4.5005
R62984 VSS.n3776 VSS.n3732 4.5005
R62985 VSS.n3774 VSS.n3733 4.5005
R62986 VSS.n3772 VSS.n3734 4.5005
R62987 VSS.n3770 VSS.n3735 4.5005
R62988 VSS.n3768 VSS.n3736 4.5005
R62989 VSS.n3765 VSS.n3737 4.5005
R62990 VSS.n3764 VSS.n3738 4.5005
R62991 VSS.n3762 VSS.n3739 4.5005
R62992 VSS.n3760 VSS.n3740 4.5005
R62993 VSS.n3758 VSS.n3741 4.5005
R62994 VSS.n3756 VSS.n3742 4.5005
R62995 VSS.n3754 VSS.n3743 4.5005
R62996 VSS.n3752 VSS.n3744 4.5005
R62997 VSS.n3749 VSS.n3745 4.5005
R62998 VSS.n3748 VSS.n3746 4.5005
R62999 VSS.n3162 VSS.n3160 4.5005
R63000 VSS.n3796 VSS.n3721 4.5005
R63001 VSS.n6310 VSS.n6309 4.5005
R63002 VSS.n6033 VSS.n5960 4.5005
R63003 VSS.n6032 VSS.n5961 4.5005
R63004 VSS.n5964 VSS.n5962 4.5005
R63005 VSS.n6028 VSS.n5965 4.5005
R63006 VSS.n6027 VSS.n5966 4.5005
R63007 VSS.n6026 VSS.n5967 4.5005
R63008 VSS.n5970 VSS.n5968 4.5005
R63009 VSS.n6022 VSS.n5971 4.5005
R63010 VSS.n6021 VSS.n5972 4.5005
R63011 VSS.n6020 VSS.n5973 4.5005
R63012 VSS.n5976 VSS.n5974 4.5005
R63013 VSS.n6016 VSS.n5977 4.5005
R63014 VSS.n6015 VSS.n5978 4.5005
R63015 VSS.n6014 VSS.n5979 4.5005
R63016 VSS.n5982 VSS.n5980 4.5005
R63017 VSS.n6010 VSS.n5983 4.5005
R63018 VSS.n6009 VSS.n5984 4.5005
R63019 VSS.n6008 VSS.n5985 4.5005
R63020 VSS.n5988 VSS.n5986 4.5005
R63021 VSS.n6004 VSS.n5989 4.5005
R63022 VSS.n6003 VSS.n5990 4.5005
R63023 VSS.n6002 VSS.n5991 4.5005
R63024 VSS.n5994 VSS.n5992 4.5005
R63025 VSS.n5998 VSS.n5995 4.5005
R63026 VSS.n5997 VSS.n5996 4.5005
R63027 VSS.n3713 VSS.n3712 4.5005
R63028 VSS.n6034 VSS.n5959 4.5005
R63029 VSS.n5905 VSS.n4068 4.5005
R63030 VSS.n6121 VSS.n4030 4.5005
R63031 VSS.n6120 VSS.n4031 4.5005
R63032 VSS.n4034 VSS.n4032 4.5005
R63033 VSS.n6116 VSS.n4035 4.5005
R63034 VSS.n6115 VSS.n4036 4.5005
R63035 VSS.n6114 VSS.n4037 4.5005
R63036 VSS.n4040 VSS.n4038 4.5005
R63037 VSS.n6110 VSS.n4041 4.5005
R63038 VSS.n6109 VSS.n4042 4.5005
R63039 VSS.n6108 VSS.n4043 4.5005
R63040 VSS.n4046 VSS.n4044 4.5005
R63041 VSS.n6104 VSS.n4047 4.5005
R63042 VSS.n6103 VSS.n4048 4.5005
R63043 VSS.n6102 VSS.n4049 4.5005
R63044 VSS.n4052 VSS.n4050 4.5005
R63045 VSS.n6098 VSS.n4053 4.5005
R63046 VSS.n6097 VSS.n4054 4.5005
R63047 VSS.n6096 VSS.n4055 4.5005
R63048 VSS.n4058 VSS.n4056 4.5005
R63049 VSS.n6092 VSS.n4059 4.5005
R63050 VSS.n6091 VSS.n4060 4.5005
R63051 VSS.n6090 VSS.n4061 4.5005
R63052 VSS.n4064 VSS.n4062 4.5005
R63053 VSS.n6086 VSS.n4065 4.5005
R63054 VSS.n6085 VSS.n4066 4.5005
R63055 VSS.n6084 VSS.n4067 4.5005
R63056 VSS.n6122 VSS.n4029 4.5005
R63057 VSS.n5719 VSS.n4075 4.5005
R63058 VSS.n5660 VSS.n5659 4.5005
R63059 VSS.n4260 VSS.n4259 4.5005
R63060 VSS.n5667 VSS.n5666 4.5005
R63061 VSS.n4244 VSS.n4243 4.5005
R63062 VSS.n5672 VSS.n5671 4.5005
R63063 VSS.n4241 VSS.n4240 4.5005
R63064 VSS.n5677 VSS.n5676 4.5005
R63065 VSS.n5678 VSS.n4239 4.5005
R63066 VSS.n5680 VSS.n5679 4.5005
R63067 VSS.n4237 VSS.n4236 4.5005
R63068 VSS.n5685 VSS.n5684 4.5005
R63069 VSS.n5686 VSS.n4235 4.5005
R63070 VSS.n5688 VSS.n5687 4.5005
R63071 VSS.n4233 VSS.n4232 4.5005
R63072 VSS.n5693 VSS.n5692 4.5005
R63073 VSS.n5694 VSS.n4231 4.5005
R63074 VSS.n5696 VSS.n5695 4.5005
R63075 VSS.n4229 VSS.n4228 4.5005
R63076 VSS.n5701 VSS.n5700 4.5005
R63077 VSS.n5702 VSS.n4227 4.5005
R63078 VSS.n5705 VSS.n5704 4.5005
R63079 VSS.n5703 VSS.n4224 4.5005
R63080 VSS.n5709 VSS.n4225 4.5005
R63081 VSS.n5712 VSS.n5710 4.5005
R63082 VSS.n5714 VSS.n4223 4.5005
R63083 VSS.n5717 VSS.n5716 4.5005
R63084 VSS.n5658 VSS.n5657 4.5005
R63085 VSS.n4924 VSS.n4923 4.5005
R63086 VSS.n4964 VSS.n4874 4.5005
R63087 VSS.n4877 VSS.n4875 4.5005
R63088 VSS.n4960 VSS.n4878 4.5005
R63089 VSS.n4959 VSS.n4879 4.5005
R63090 VSS.n4958 VSS.n4880 4.5005
R63091 VSS.n4883 VSS.n4881 4.5005
R63092 VSS.n4954 VSS.n4884 4.5005
R63093 VSS.n4953 VSS.n4885 4.5005
R63094 VSS.n4952 VSS.n4886 4.5005
R63095 VSS.n4889 VSS.n4887 4.5005
R63096 VSS.n4948 VSS.n4890 4.5005
R63097 VSS.n4947 VSS.n4891 4.5005
R63098 VSS.n4946 VSS.n4892 4.5005
R63099 VSS.n4895 VSS.n4893 4.5005
R63100 VSS.n4942 VSS.n4896 4.5005
R63101 VSS.n4941 VSS.n4897 4.5005
R63102 VSS.n4940 VSS.n4898 4.5005
R63103 VSS.n4901 VSS.n4899 4.5005
R63104 VSS.n4936 VSS.n4902 4.5005
R63105 VSS.n4935 VSS.n4903 4.5005
R63106 VSS.n4934 VSS.n4904 4.5005
R63107 VSS.n4907 VSS.n4905 4.5005
R63108 VSS.n4930 VSS.n4908 4.5005
R63109 VSS.n4929 VSS.n4909 4.5005
R63110 VSS.n4928 VSS.n4910 4.5005
R63111 VSS.n4912 VSS.n4911 4.5005
R63112 VSS.n4966 VSS.n4965 4.5005
R63113 VSS.n4866 VSS.n4865 4.5005
R63114 VSS.n5122 VSS.n4457 4.5005
R63115 VSS.n5120 VSS.n4458 4.5005
R63116 VSS.n5118 VSS.n4459 4.5005
R63117 VSS.n5116 VSS.n4460 4.5005
R63118 VSS.n4463 VSS.n4461 4.5005
R63119 VSS.n5112 VSS.n4464 4.5005
R63120 VSS.n5111 VSS.n4465 4.5005
R63121 VSS.n5110 VSS.n4466 4.5005
R63122 VSS.n4469 VSS.n4467 4.5005
R63123 VSS.n5106 VSS.n4470 4.5005
R63124 VSS.n5105 VSS.n4471 4.5005
R63125 VSS.n5104 VSS.n4472 4.5005
R63126 VSS.n4475 VSS.n4473 4.5005
R63127 VSS.n5100 VSS.n4476 4.5005
R63128 VSS.n5099 VSS.n4477 4.5005
R63129 VSS.n5098 VSS.n4478 4.5005
R63130 VSS.n4481 VSS.n4479 4.5005
R63131 VSS.n5094 VSS.n4482 4.5005
R63132 VSS.n5093 VSS.n4483 4.5005
R63133 VSS.n5092 VSS.n4484 4.5005
R63134 VSS.n4487 VSS.n4485 4.5005
R63135 VSS.n5088 VSS.n4488 4.5005
R63136 VSS.n5087 VSS.n4489 4.5005
R63137 VSS.n4856 VSS.n4490 4.5005
R63138 VSS.n4861 VSS.n4859 4.5005
R63139 VSS.n4863 VSS.n4858 4.5005
R63140 VSS.n5125 VSS.n5124 4.5005
R63141 VSS.n7146 VSS.n2470 4.5005
R63142 VSS.n5020 VSS.n4855 4.5005
R63143 VSS.n4872 VSS.n4855 4.5005
R63144 VSS.n5018 VSS.n4855 4.5005
R63145 VSS.n5020 VSS.n4853 4.5005
R63146 VSS.n4872 VSS.n4853 4.5005
R63147 VSS.n5018 VSS.n4853 4.5005
R63148 VSS.n5020 VSS.n4857 4.5005
R63149 VSS.n4872 VSS.n4857 4.5005
R63150 VSS.n5018 VSS.n4857 4.5005
R63151 VSS.n5018 VSS.n4852 4.5005
R63152 VSS.n4872 VSS.n4852 4.5005
R63153 VSS.n5020 VSS.n4852 4.5005
R63154 VSS.n5018 VSS.n4867 4.5005
R63155 VSS.n4872 VSS.n4867 4.5005
R63156 VSS.n5020 VSS.n4867 4.5005
R63157 VSS.n5018 VSS.n4851 4.5005
R63158 VSS.n5020 VSS.n4851 4.5005
R63159 VSS.n5018 VSS.n4868 4.5005
R63160 VSS.n5020 VSS.n4868 4.5005
R63161 VSS.n5018 VSS.n4850 4.5005
R63162 VSS.n4872 VSS.n4850 4.5005
R63163 VSS.n5020 VSS.n4850 4.5005
R63164 VSS.n5018 VSS.n4869 4.5005
R63165 VSS.n4872 VSS.n4869 4.5005
R63166 VSS.n5020 VSS.n4869 4.5005
R63167 VSS.n5018 VSS.n4849 4.5005
R63168 VSS.n4872 VSS.n4849 4.5005
R63169 VSS.n5020 VSS.n4849 4.5005
R63170 VSS.n5019 VSS.n5018 4.5005
R63171 VSS.n5019 VSS.n4872 4.5005
R63172 VSS.n5020 VSS.n5019 4.5005
R63173 VSS.n4254 VSS.n4246 4.5005
R63174 VSS.n4254 VSS.n4245 4.5005
R63175 VSS.n5669 VSS.n4254 4.5005
R63176 VSS.n4252 VSS.n4246 4.5005
R63177 VSS.n4252 VSS.n4245 4.5005
R63178 VSS.n5669 VSS.n4252 4.5005
R63179 VSS.n4255 VSS.n4246 4.5005
R63180 VSS.n4255 VSS.n4245 4.5005
R63181 VSS.n5669 VSS.n4255 4.5005
R63182 VSS.n4251 VSS.n4246 4.5005
R63183 VSS.n4251 VSS.n4245 4.5005
R63184 VSS.n5669 VSS.n4251 4.5005
R63185 VSS.n4257 VSS.n4246 4.5005
R63186 VSS.n5669 VSS.n4257 4.5005
R63187 VSS.n4250 VSS.n4246 4.5005
R63188 VSS.n5669 VSS.n4250 4.5005
R63189 VSS.n5669 VSS.n4258 4.5005
R63190 VSS.n4258 VSS.n4245 4.5005
R63191 VSS.n4258 VSS.n4246 4.5005
R63192 VSS.n5669 VSS.n4249 4.5005
R63193 VSS.n4249 VSS.n4245 4.5005
R63194 VSS.n4249 VSS.n4246 4.5005
R63195 VSS.n5668 VSS.n4246 4.5005
R63196 VSS.n5668 VSS.n4245 4.5005
R63197 VSS.n5669 VSS.n5668 4.5005
R63198 VSS.n4248 VSS.n4246 4.5005
R63199 VSS.n4248 VSS.n4245 4.5005
R63200 VSS.n5669 VSS.n4248 4.5005
R63201 VSS.n5670 VSS.n4246 4.5005
R63202 VSS.n5670 VSS.n4245 4.5005
R63203 VSS.n5670 VSS.n5669 4.5005
R63204 VSS.n4222 VSS.n4171 4.5005
R63205 VSS.n4222 VSS.n4170 4.5005
R63206 VSS.n5723 VSS.n4222 4.5005
R63207 VSS.n4175 VSS.n4171 4.5005
R63208 VSS.n4175 VSS.n4170 4.5005
R63209 VSS.n5723 VSS.n4175 4.5005
R63210 VSS.n5718 VSS.n4171 4.5005
R63211 VSS.n5718 VSS.n4170 4.5005
R63212 VSS.n5723 VSS.n5718 4.5005
R63213 VSS.n5723 VSS.n4174 4.5005
R63214 VSS.n4174 VSS.n4170 4.5005
R63215 VSS.n4174 VSS.n4171 4.5005
R63216 VSS.n5723 VSS.n5721 4.5005
R63217 VSS.n5721 VSS.n4171 4.5005
R63218 VSS.n5723 VSS.n4173 4.5005
R63219 VSS.n4173 VSS.n4171 4.5005
R63220 VSS.n4171 VSS.n4120 4.5005
R63221 VSS.n4170 VSS.n4120 4.5005
R63222 VSS.n5723 VSS.n4120 4.5005
R63223 VSS.n4171 VSS.n4122 4.5005
R63224 VSS.n4170 VSS.n4122 4.5005
R63225 VSS.n5723 VSS.n4122 4.5005
R63226 VSS.n5722 VSS.n4171 4.5005
R63227 VSS.n5722 VSS.n4170 4.5005
R63228 VSS.n5723 VSS.n5722 4.5005
R63229 VSS.n4171 VSS.n4169 4.5005
R63230 VSS.n4170 VSS.n4169 4.5005
R63231 VSS.n5723 VSS.n4169 4.5005
R63232 VSS.n5724 VSS.n4171 4.5005
R63233 VSS.n5724 VSS.n4170 4.5005
R63234 VSS.n5724 VSS.n5723 4.5005
R63235 VSS.n6615 VSS.n3148 4.5005
R63236 VSS.n3161 VSS.n3148 4.5005
R63237 VSS.n3148 VSS.n3135 4.5005
R63238 VSS.n6615 VSS.n3150 4.5005
R63239 VSS.n3161 VSS.n3150 4.5005
R63240 VSS.n3150 VSS.n3135 4.5005
R63241 VSS.n3147 VSS.n3135 4.5005
R63242 VSS.n3161 VSS.n3147 4.5005
R63243 VSS.n6615 VSS.n3147 4.5005
R63244 VSS.n3151 VSS.n3135 4.5005
R63245 VSS.n3161 VSS.n3151 4.5005
R63246 VSS.n6615 VSS.n3151 4.5005
R63247 VSS.n3146 VSS.n3135 4.5005
R63248 VSS.n3161 VSS.n3146 4.5005
R63249 VSS.n6615 VSS.n3146 4.5005
R63250 VSS.n3152 VSS.n3135 4.5005
R63251 VSS.n3161 VSS.n3152 4.5005
R63252 VSS.n6615 VSS.n3152 4.5005
R63253 VSS.n6615 VSS.n3145 4.5005
R63254 VSS.n3161 VSS.n3145 4.5005
R63255 VSS.n3145 VSS.n3135 4.5005
R63256 VSS.n6615 VSS.n3153 4.5005
R63257 VSS.n3161 VSS.n3153 4.5005
R63258 VSS.n3153 VSS.n3135 4.5005
R63259 VSS.n6615 VSS.n3144 4.5005
R63260 VSS.n3161 VSS.n3144 4.5005
R63261 VSS.n3144 VSS.n3135 4.5005
R63262 VSS.n3154 VSS.n3135 4.5005
R63263 VSS.n3161 VSS.n3154 4.5005
R63264 VSS.n6615 VSS.n3154 4.5005
R63265 VSS.n3143 VSS.n3135 4.5005
R63266 VSS.n3161 VSS.n3143 4.5005
R63267 VSS.n6615 VSS.n3143 4.5005
R63268 VSS.n3155 VSS.n3135 4.5005
R63269 VSS.n3161 VSS.n3155 4.5005
R63270 VSS.n6615 VSS.n3155 4.5005
R63271 VSS.n6615 VSS.n3142 4.5005
R63272 VSS.n3161 VSS.n3142 4.5005
R63273 VSS.n3142 VSS.n3135 4.5005
R63274 VSS.n6615 VSS.n3156 4.5005
R63275 VSS.n3161 VSS.n3156 4.5005
R63276 VSS.n3156 VSS.n3135 4.5005
R63277 VSS.n6615 VSS.n3141 4.5005
R63278 VSS.n3161 VSS.n3141 4.5005
R63279 VSS.n3141 VSS.n3135 4.5005
R63280 VSS.n6615 VSS.n3157 4.5005
R63281 VSS.n3161 VSS.n3157 4.5005
R63282 VSS.n3157 VSS.n3135 4.5005
R63283 VSS.n3140 VSS.n3135 4.5005
R63284 VSS.n3161 VSS.n3140 4.5005
R63285 VSS.n6615 VSS.n3140 4.5005
R63286 VSS.n3158 VSS.n3135 4.5005
R63287 VSS.n3161 VSS.n3158 4.5005
R63288 VSS.n6615 VSS.n3158 4.5005
R63289 VSS.n3139 VSS.n3135 4.5005
R63290 VSS.n3161 VSS.n3139 4.5005
R63291 VSS.n6615 VSS.n3139 4.5005
R63292 VSS.n6615 VSS.n3159 4.5005
R63293 VSS.n3161 VSS.n3159 4.5005
R63294 VSS.n3159 VSS.n3135 4.5005
R63295 VSS.n6615 VSS.n3138 4.5005
R63296 VSS.n3161 VSS.n3138 4.5005
R63297 VSS.n3138 VSS.n3135 4.5005
R63298 VSS.n6615 VSS.n6614 4.5005
R63299 VSS.n6614 VSS.n3161 4.5005
R63300 VSS.n6614 VSS.n3135 4.5005
R63301 VSS.n3137 VSS.n3135 4.5005
R63302 VSS.n6615 VSS.n3137 4.5005
R63303 VSS.n6616 VSS.n3135 4.5005
R63304 VSS.n6616 VSS.n6615 4.5005
R63305 VSS.n6805 VSS.n2949 4.5005
R63306 VSS.n2949 VSS.n2940 4.5005
R63307 VSS.n2949 VSS.n2941 4.5005
R63308 VSS.n6805 VSS.n2947 4.5005
R63309 VSS.n2947 VSS.n2940 4.5005
R63310 VSS.n2947 VSS.n2941 4.5005
R63311 VSS.n2950 VSS.n2941 4.5005
R63312 VSS.n2950 VSS.n2940 4.5005
R63313 VSS.n6805 VSS.n2950 4.5005
R63314 VSS.n2946 VSS.n2941 4.5005
R63315 VSS.n2946 VSS.n2940 4.5005
R63316 VSS.n6805 VSS.n2946 4.5005
R63317 VSS.n2951 VSS.n2941 4.5005
R63318 VSS.n2951 VSS.n2940 4.5005
R63319 VSS.n6805 VSS.n2951 4.5005
R63320 VSS.n2945 VSS.n2941 4.5005
R63321 VSS.n2945 VSS.n2940 4.5005
R63322 VSS.n6805 VSS.n2945 4.5005
R63323 VSS.n6805 VSS.n2952 4.5005
R63324 VSS.n2952 VSS.n2940 4.5005
R63325 VSS.n2952 VSS.n2941 4.5005
R63326 VSS.n6805 VSS.n2944 4.5005
R63327 VSS.n2944 VSS.n2940 4.5005
R63328 VSS.n2944 VSS.n2941 4.5005
R63329 VSS.n6805 VSS.n6804 4.5005
R63330 VSS.n6804 VSS.n2940 4.5005
R63331 VSS.n6804 VSS.n2941 4.5005
R63332 VSS.n2943 VSS.n2941 4.5005
R63333 VSS.n2943 VSS.n2940 4.5005
R63334 VSS.n6805 VSS.n2943 4.5005
R63335 VSS.n6806 VSS.n2941 4.5005
R63336 VSS.n6806 VSS.n2940 4.5005
R63337 VSS.n6806 VSS.n6805 4.5005
R63338 VSS.n8816 VSS.n8815 4.5005
R63339 VSS.n8815 VSS.n1368 4.5005
R63340 VSS.n8813 VSS.n1368 4.5005
R63341 VSS.n1383 VSS.n1368 4.5005
R63342 VSS.n1382 VSS.n1368 4.5005
R63343 VSS.n8812 VSS.n1385 4.5005
R63344 VSS.n1385 VSS.n1368 4.5005
R63345 VSS.n8816 VSS.n1373 4.5005
R63346 VSS.n8812 VSS.n1373 4.5005
R63347 VSS.n1373 VSS.n1368 4.5005
R63348 VSS.n8817 VSS.n1368 4.5005
R63349 VSS.n8817 VSS.n8816 4.5005
R63350 VSS.n1371 VSS.n1368 4.5005
R63351 VSS.n1380 VSS.n1368 4.5005
R63352 VSS.n1379 VSS.n1368 4.5005
R63353 VSS.n8812 VSS.n8811 4.5005
R63354 VSS.n8811 VSS.n1368 4.5005
R63355 VSS.n8712 VSS.n1452 4.5005
R63356 VSS.n8710 VSS.n1452 4.5005
R63357 VSS.n8712 VSS.n1453 4.5005
R63358 VSS.n8710 VSS.n1453 4.5005
R63359 VSS.n8710 VSS.n1451 4.5005
R63360 VSS.n1462 VSS.n1451 4.5005
R63361 VSS.n8712 VSS.n1451 4.5005
R63362 VSS.n8710 VSS.n1454 4.5005
R63363 VSS.n8712 VSS.n1454 4.5005
R63364 VSS.n8710 VSS.n1473 4.5005
R63365 VSS.n8710 VSS.n8695 4.5005
R63366 VSS.n8710 VSS.n1471 4.5005
R63367 VSS.n8710 VSS.n8697 4.5005
R63368 VSS.n8710 VSS.n1470 4.5005
R63369 VSS.n8710 VSS.n8699 4.5005
R63370 VSS.n8710 VSS.n1469 4.5005
R63371 VSS.n8710 VSS.n8701 4.5005
R63372 VSS.n8712 VSS.n1446 4.5005
R63373 VSS.n8710 VSS.n1446 4.5005
R63374 VSS.n8712 VSS.n1455 4.5005
R63375 VSS.n1462 VSS.n1455 4.5005
R63376 VSS.n8710 VSS.n1455 4.5005
R63377 VSS.n8712 VSS.n1445 4.5005
R63378 VSS.n8710 VSS.n1445 4.5005
R63379 VSS.n8710 VSS.n8703 4.5005
R63380 VSS.n8710 VSS.n1468 4.5005
R63381 VSS.n8710 VSS.n8705 4.5005
R63382 VSS.n8710 VSS.n1467 4.5005
R63383 VSS.n8710 VSS.n8707 4.5005
R63384 VSS.n8710 VSS.n1466 4.5005
R63385 VSS.n8710 VSS.n8709 4.5005
R63386 VSS.n1465 VSS.n1462 4.5005
R63387 VSS.n8710 VSS.n1465 4.5005
R63388 VSS.n8711 VSS.n8710 4.5005
R63389 VSS.n8711 VSS.n1462 4.5005
R63390 VSS.n8712 VSS.n8711 4.5005
R63391 VSS.n995 VSS.n981 4.5005
R63392 VSS.n9109 VSS.n995 4.5005
R63393 VSS.n9080 VSS.n981 4.5005
R63394 VSS.n9079 VSS.n981 4.5005
R63395 VSS.n9083 VSS.n981 4.5005
R63396 VSS.n9082 VSS.n981 4.5005
R63397 VSS.n9086 VSS.n981 4.5005
R63398 VSS.n9085 VSS.n981 4.5005
R63399 VSS.n9089 VSS.n981 4.5005
R63400 VSS.n9088 VSS.n981 4.5005
R63401 VSS.n9092 VSS.n981 4.5005
R63402 VSS.n9091 VSS.n981 4.5005
R63403 VSS.n9095 VSS.n981 4.5005
R63404 VSS.n9094 VSS.n981 4.5005
R63405 VSS.n9098 VSS.n981 4.5005
R63406 VSS.n9097 VSS.n981 4.5005
R63407 VSS.n9101 VSS.n981 4.5005
R63408 VSS.n9100 VSS.n981 4.5005
R63409 VSS.n9104 VSS.n981 4.5005
R63410 VSS.n9103 VSS.n981 4.5005
R63411 VSS.n9107 VSS.n981 4.5005
R63412 VSS.n9106 VSS.n981 4.5005
R63413 VSS.n9110 VSS.n981 4.5005
R63414 VSS.n9112 VSS.n981 4.5005
R63415 VSS.n9109 VSS.n994 4.5005
R63416 VSS.n994 VSS.n981 4.5005
R63417 VSS.n9256 VSS.n874 4.5005
R63418 VSS.n9253 VSS.n874 4.5005
R63419 VSS.n9253 VSS.n9231 4.5005
R63420 VSS.n9253 VSS.n897 4.5005
R63421 VSS.n9253 VSS.n9232 4.5005
R63422 VSS.n9253 VSS.n896 4.5005
R63423 VSS.n9253 VSS.n9233 4.5005
R63424 VSS.n9253 VSS.n895 4.5005
R63425 VSS.n9253 VSS.n9234 4.5005
R63426 VSS.n9253 VSS.n894 4.5005
R63427 VSS.n9253 VSS.n9235 4.5005
R63428 VSS.n9253 VSS.n893 4.5005
R63429 VSS.n9253 VSS.n9236 4.5005
R63430 VSS.n9253 VSS.n892 4.5005
R63431 VSS.n9253 VSS.n9237 4.5005
R63432 VSS.n9253 VSS.n891 4.5005
R63433 VSS.n9253 VSS.n9238 4.5005
R63434 VSS.n9253 VSS.n890 4.5005
R63435 VSS.n9253 VSS.n9239 4.5005
R63436 VSS.n9253 VSS.n889 4.5005
R63437 VSS.n9253 VSS.n9252 4.5005
R63438 VSS.n9253 VSS.n888 4.5005
R63439 VSS.n9254 VSS.n9253 4.5005
R63440 VSS.n9253 VSS.n885 4.5005
R63441 VSS.n9256 VSS.n766 4.5005
R63442 VSS.n9253 VSS.n766 4.5005
R63443 VSS.n7217 VSS.n2530 4.5005
R63444 VSS.n7220 VSS.n2530 4.5005
R63445 VSS.n7223 VSS.n2530 4.5005
R63446 VSS.n7214 VSS.n7213 4.5005
R63447 VSS.n7220 VSS.n2528 4.5005
R63448 VSS.n7223 VSS.n2528 4.5005
R63449 VSS.n7211 VSS.n2534 4.5005
R63450 VSS.n7222 VSS.n7217 4.5005
R63451 VSS.n7223 VSS.n7222 4.5005
R63452 VSS.n7081 VSS.n7063 4.5005
R63453 VSS.n7084 VSS.n7063 4.5005
R63454 VSS.n7094 VSS.n7085 4.5005
R63455 VSS.n7094 VSS.n7093 4.5005
R63456 VSS.n7095 VSS.n7094 4.5005
R63457 VSS.n7084 VSS.n7061 4.5005
R63458 VSS.n7093 VSS.n2532 4.5005
R63459 VSS.n7095 VSS.n2532 4.5005
R63460 VSS.n7084 VSS.n7083 4.5005
R63461 VSS.n7096 VSS.n7085 4.5005
R63462 VSS.n7096 VSS.n7095 4.5005
R63463 VSS.n7171 VSS.n2543 4.5005
R63464 VSS.n7171 VSS.n7170 4.5005
R63465 VSS.n7169 VSS.n2548 4.5005
R63466 VSS.n7165 VSS.n2548 4.5005
R63467 VSS.n7167 VSS.n2548 4.5005
R63468 VSS.n7170 VSS.n2546 4.5005
R63469 VSS.n7166 VSS.n7165 4.5005
R63470 VSS.n7167 VSS.n7166 4.5005
R63471 VSS.n7170 VSS.n2536 4.5005
R63472 VSS.n7169 VSS.n7168 4.5005
R63473 VSS.n7168 VSS.n7167 4.5005
R63474 VSS.n2563 VSS.n2557 4.5005
R63475 VSS.n7159 VSS.n7158 4.5005
R63476 VSS.n7159 VSS.n2554 4.5005
R63477 VSS.n7162 VSS.n2554 4.5005
R63478 VSS.n7162 VSS.n7161 4.5005
R63479 VSS.n2563 VSS.n2562 4.5005
R63480 VSS.n2562 VSS.n2559 4.5005
R63481 VSS.n2562 VSS.n2561 4.5005
R63482 VSS.n2493 VSS.n2480 4.5005
R63483 VSS.n7263 VSS.n2480 4.5005
R63484 VSS.n7263 VSS.n7262 4.5005
R63485 VSS.n7262 VSS.n7261 4.5005
R63486 VSS.n7245 VSS.n7243 4.5005
R63487 VSS.n7243 VSS.n2506 4.5005
R63488 VSS.n7240 VSS.n2508 4.5005
R63489 VSS.n7240 VSS.n7239 4.5005
R63490 VSS.n7241 VSS.n7240 4.5005
R63491 VSS.n7239 VSS.n2511 4.5005
R63492 VSS.n7241 VSS.n2511 4.5005
R63493 VSS.n7192 VSS.n7188 4.5005
R63494 VSS.n7195 VSS.n7188 4.5005
R63495 VSS.n7198 VSS.n7188 4.5005
R63496 VSS.n7195 VSS.n2491 4.5005
R63497 VSS.n7198 VSS.n2491 4.5005
R63498 VSS.n7255 VSS.n2488 4.5005
R63499 VSS.n2488 VSS.n2485 4.5005
R63500 VSS.n7258 VSS.n2488 4.5005
R63501 VSS.n7259 VSS.n2485 4.5005
R63502 VSS.n7259 VSS.n7258 4.5005
R63503 VSS.n7257 VSS.n7255 4.5005
R63504 VSS.n7258 VSS.n7257 4.5005
R63505 VSS.n7197 VSS.n7192 4.5005
R63506 VSS.n7198 VSS.n7197 4.5005
R63507 VSS.n7242 VSS.n2508 4.5005
R63508 VSS.n7242 VSS.n7241 4.5005
R63509 VSS.n7247 VSS.n2506 4.5005
R63510 VSS.n7248 VSS.n7247 4.5005
R63511 VSS.n5062 VSS.n4523 4.5005
R63512 VSS.n5062 VSS.n4524 4.5005
R63513 VSS.n5071 VSS.n5062 4.5005
R63514 VSS.n4528 VSS.n4524 4.5005
R63515 VSS.n5071 VSS.n4528 4.5005
R63516 VSS.n5065 VSS.n4524 4.5005
R63517 VSS.n5071 VSS.n5065 4.5005
R63518 VSS.n4527 VSS.n4524 4.5005
R63519 VSS.n5071 VSS.n4527 4.5005
R63520 VSS.n5068 VSS.n4524 4.5005
R63521 VSS.n5071 VSS.n5068 4.5005
R63522 VSS.n4526 VSS.n4524 4.5005
R63523 VSS.n5071 VSS.n4526 4.5005
R63524 VSS.n5070 VSS.n4524 4.5005
R63525 VSS.n5070 VSS.n4522 4.5005
R63526 VSS.n5071 VSS.n5070 4.5005
R63527 VSS.n4523 VSS.n4517 4.5005
R63528 VSS.n4524 VSS.n4517 4.5005
R63529 VSS.n4522 VSS.n4517 4.5005
R63530 VSS.n5071 VSS.n4517 4.5005
R63531 VSS.n4523 VSS.n4520 4.5005
R63532 VSS.n4524 VSS.n4520 4.5005
R63533 VSS.n4522 VSS.n4520 4.5005
R63534 VSS.n5071 VSS.n4520 4.5005
R63535 VSS.n4523 VSS.n4521 4.5005
R63536 VSS.n4524 VSS.n4521 4.5005
R63537 VSS.n4522 VSS.n4521 4.5005
R63538 VSS.n5071 VSS.n4521 4.5005
R63539 VSS.n5072 VSS.n4523 4.5005
R63540 VSS.n5072 VSS.n4524 4.5005
R63541 VSS.n5072 VSS.n4522 4.5005
R63542 VSS.n5072 VSS.n5071 4.5005
R63543 VSS.n4290 VSS.n4284 4.5005
R63544 VSS.n4291 VSS.n4284 4.5005
R63545 VSS.n4289 VSS.n4284 4.5005
R63546 VSS.n5641 VSS.n4284 4.5005
R63547 VSS.n4290 VSS.n4287 4.5005
R63548 VSS.n4291 VSS.n4287 4.5005
R63549 VSS.n4289 VSS.n4287 4.5005
R63550 VSS.n5641 VSS.n4287 4.5005
R63551 VSS.n4290 VSS.n4288 4.5005
R63552 VSS.n4291 VSS.n4288 4.5005
R63553 VSS.n4289 VSS.n4288 4.5005
R63554 VSS.n5641 VSS.n4288 4.5005
R63555 VSS.n5642 VSS.n4290 4.5005
R63556 VSS.n5642 VSS.n4291 4.5005
R63557 VSS.n5642 VSS.n4289 4.5005
R63558 VSS.n5642 VSS.n5641 4.5005
R63559 VSS.n5632 VSS.n4290 4.5005
R63560 VSS.n5632 VSS.n4291 4.5005
R63561 VSS.n5641 VSS.n5632 4.5005
R63562 VSS.n4295 VSS.n4291 4.5005
R63563 VSS.n5641 VSS.n4295 4.5005
R63564 VSS.n5635 VSS.n4291 4.5005
R63565 VSS.n5641 VSS.n5635 4.5005
R63566 VSS.n4294 VSS.n4291 4.5005
R63567 VSS.n5641 VSS.n4294 4.5005
R63568 VSS.n5638 VSS.n4291 4.5005
R63569 VSS.n5641 VSS.n5638 4.5005
R63570 VSS.n4293 VSS.n4291 4.5005
R63571 VSS.n5641 VSS.n4293 4.5005
R63572 VSS.n5640 VSS.n4291 4.5005
R63573 VSS.n5640 VSS.n4289 4.5005
R63574 VSS.n5641 VSS.n5640 4.5005
R63575 VSS.n6159 VSS.n3988 4.5005
R63576 VSS.n6161 VSS.n3988 4.5005
R63577 VSS.n3988 VSS.n3975 4.5005
R63578 VSS.n6161 VSS.n3985 4.5005
R63579 VSS.n3985 VSS.n3975 4.5005
R63580 VSS.n6161 VSS.n3990 4.5005
R63581 VSS.n3990 VSS.n3975 4.5005
R63582 VSS.n6161 VSS.n3984 4.5005
R63583 VSS.n3984 VSS.n3975 4.5005
R63584 VSS.n6161 VSS.n3992 4.5005
R63585 VSS.n3992 VSS.n3975 4.5005
R63586 VSS.n6159 VSS.n3983 4.5005
R63587 VSS.n6161 VSS.n3983 4.5005
R63588 VSS.n3983 VSS.n3975 4.5005
R63589 VSS.n3993 VSS.n3975 4.5005
R63590 VSS.n3993 VSS.n3980 4.5005
R63591 VSS.n6161 VSS.n3993 4.5005
R63592 VSS.n6159 VSS.n3993 4.5005
R63593 VSS.n3982 VSS.n3975 4.5005
R63594 VSS.n3982 VSS.n3980 4.5005
R63595 VSS.n6161 VSS.n3982 4.5005
R63596 VSS.n6159 VSS.n3982 4.5005
R63597 VSS.n3994 VSS.n3975 4.5005
R63598 VSS.n3994 VSS.n3980 4.5005
R63599 VSS.n6161 VSS.n3994 4.5005
R63600 VSS.n6159 VSS.n3994 4.5005
R63601 VSS.n3981 VSS.n3975 4.5005
R63602 VSS.n3981 VSS.n3980 4.5005
R63603 VSS.n6161 VSS.n3981 4.5005
R63604 VSS.n6159 VSS.n3981 4.5005
R63605 VSS.n6160 VSS.n3975 4.5005
R63606 VSS.n6160 VSS.n3980 4.5005
R63607 VSS.n6161 VSS.n6160 4.5005
R63608 VSS.n6160 VSS.n6159 4.5005
R63609 VSS.n3451 VSS.n3426 4.5005
R63610 VSS.n6505 VSS.n3426 4.5005
R63611 VSS.n6507 VSS.n3426 4.5005
R63612 VSS.n6505 VSS.n3428 4.5005
R63613 VSS.n6507 VSS.n3428 4.5005
R63614 VSS.n6505 VSS.n3425 4.5005
R63615 VSS.n6507 VSS.n3425 4.5005
R63616 VSS.n6505 VSS.n3429 4.5005
R63617 VSS.n6507 VSS.n3429 4.5005
R63618 VSS.n6505 VSS.n3424 4.5005
R63619 VSS.n6507 VSS.n3424 4.5005
R63620 VSS.n6505 VSS.n3430 4.5005
R63621 VSS.n6507 VSS.n3430 4.5005
R63622 VSS.n6505 VSS.n3423 4.5005
R63623 VSS.n6507 VSS.n3423 4.5005
R63624 VSS.n6505 VSS.n3431 4.5005
R63625 VSS.n6507 VSS.n3431 4.5005
R63626 VSS.n6505 VSS.n3422 4.5005
R63627 VSS.n6507 VSS.n3422 4.5005
R63628 VSS.n6505 VSS.n3432 4.5005
R63629 VSS.n6507 VSS.n3432 4.5005
R63630 VSS.n6505 VSS.n3421 4.5005
R63631 VSS.n6507 VSS.n3421 4.5005
R63632 VSS.n6505 VSS.n3433 4.5005
R63633 VSS.n6507 VSS.n3433 4.5005
R63634 VSS.n6505 VSS.n3420 4.5005
R63635 VSS.n6507 VSS.n3420 4.5005
R63636 VSS.n6505 VSS.n3434 4.5005
R63637 VSS.n6507 VSS.n3434 4.5005
R63638 VSS.n6505 VSS.n3419 4.5005
R63639 VSS.n6507 VSS.n3419 4.5005
R63640 VSS.n6505 VSS.n3435 4.5005
R63641 VSS.n6507 VSS.n3435 4.5005
R63642 VSS.n6505 VSS.n3418 4.5005
R63643 VSS.n6507 VSS.n3418 4.5005
R63644 VSS.n6505 VSS.n3436 4.5005
R63645 VSS.n6507 VSS.n3436 4.5005
R63646 VSS.n6505 VSS.n3417 4.5005
R63647 VSS.n6507 VSS.n3417 4.5005
R63648 VSS.n6505 VSS.n3437 4.5005
R63649 VSS.n6507 VSS.n3437 4.5005
R63650 VSS.n6505 VSS.n3416 4.5005
R63651 VSS.n6507 VSS.n3416 4.5005
R63652 VSS.n6505 VSS.n3438 4.5005
R63653 VSS.n6507 VSS.n3438 4.5005
R63654 VSS.n6505 VSS.n3415 4.5005
R63655 VSS.n6507 VSS.n3415 4.5005
R63656 VSS.n6506 VSS.n3451 4.5005
R63657 VSS.n6506 VSS.n6505 4.5005
R63658 VSS.n6507 VSS.n6506 4.5005
R63659 VSS.n6876 VSS.n2898 4.5005
R63660 VSS.n6879 VSS.n2898 4.5005
R63661 VSS.n2898 VSS.n2885 4.5005
R63662 VSS.n6879 VSS.n2895 4.5005
R63663 VSS.n2895 VSS.n2885 4.5005
R63664 VSS.n6879 VSS.n2900 4.5005
R63665 VSS.n2900 VSS.n2885 4.5005
R63666 VSS.n6879 VSS.n2894 4.5005
R63667 VSS.n2894 VSS.n2885 4.5005
R63668 VSS.n6879 VSS.n2902 4.5005
R63669 VSS.n2902 VSS.n2885 4.5005
R63670 VSS.n6879 VSS.n2893 4.5005
R63671 VSS.n2893 VSS.n2885 4.5005
R63672 VSS.n6879 VSS.n2904 4.5005
R63673 VSS.n2904 VSS.n2885 4.5005
R63674 VSS.n6879 VSS.n2892 4.5005
R63675 VSS.n2892 VSS.n2885 4.5005
R63676 VSS.n6879 VSS.n2906 4.5005
R63677 VSS.n2906 VSS.n2885 4.5005
R63678 VSS.n6879 VSS.n2891 4.5005
R63679 VSS.n2891 VSS.n2885 4.5005
R63680 VSS.n6879 VSS.n6878 4.5005
R63681 VSS.n6878 VSS.n2890 4.5005
R63682 VSS.n6878 VSS.n2885 4.5005
R63683 VSS.n8412 VSS.n1659 4.5005
R63684 VSS.n1659 VSS.n1655 4.5005
R63685 VSS.n1664 VSS.n1659 4.5005
R63686 VSS.n8382 VSS.n1655 4.5005
R63687 VSS.n8382 VSS.n1664 4.5005
R63688 VSS.n8380 VSS.n1655 4.5005
R63689 VSS.n8380 VSS.n1664 4.5005
R63690 VSS.n8379 VSS.n1655 4.5005
R63691 VSS.n8379 VSS.n1664 4.5005
R63692 VSS.n8405 VSS.n1655 4.5005
R63693 VSS.n8410 VSS.n8405 4.5005
R63694 VSS.n8405 VSS.n1664 4.5005
R63695 VSS.n8412 VSS.n1658 4.5005
R63696 VSS.n1658 VSS.n1655 4.5005
R63697 VSS.n8410 VSS.n1658 4.5005
R63698 VSS.n1664 VSS.n1658 4.5005
R63699 VSS.n8411 VSS.n1664 4.5005
R63700 VSS.n8411 VSS.n8410 4.5005
R63701 VSS.n8412 VSS.n8411 4.5005
R63702 VSS.n8412 VSS.n1657 4.5005
R63703 VSS.n1664 VSS.n1657 4.5005
R63704 VSS.n8406 VSS.n1655 4.5005
R63705 VSS.n8406 VSS.n1664 4.5005
R63706 VSS.n8408 VSS.n1655 4.5005
R63707 VSS.n8408 VSS.n1664 4.5005
R63708 VSS.n8412 VSS.n1602 4.5005
R63709 VSS.n1655 VSS.n1602 4.5005
R63710 VSS.n1664 VSS.n1602 4.5005
R63711 VSS.n8635 VSS.n1535 4.5005
R63712 VSS.n1535 VSS.n1523 4.5005
R63713 VSS.n1541 VSS.n1535 4.5005
R63714 VSS.n8635 VSS.n1536 4.5005
R63715 VSS.n1536 VSS.n1523 4.5005
R63716 VSS.n1541 VSS.n1536 4.5005
R63717 VSS.n1541 VSS.n1534 4.5005
R63718 VSS.n8633 VSS.n1534 4.5005
R63719 VSS.n1534 VSS.n1523 4.5005
R63720 VSS.n8635 VSS.n1534 4.5005
R63721 VSS.n1541 VSS.n1538 4.5005
R63722 VSS.n8633 VSS.n1538 4.5005
R63723 VSS.n8635 VSS.n1538 4.5005
R63724 VSS.n8635 VSS.n1533 4.5005
R63725 VSS.n1541 VSS.n1533 4.5005
R63726 VSS.n8611 VSS.n1523 4.5005
R63727 VSS.n8611 VSS.n1541 4.5005
R63728 VSS.n8614 VSS.n1523 4.5005
R63729 VSS.n8614 VSS.n1541 4.5005
R63730 VSS.n8613 VSS.n1523 4.5005
R63731 VSS.n8613 VSS.n1541 4.5005
R63732 VSS.n8617 VSS.n1523 4.5005
R63733 VSS.n8617 VSS.n1541 4.5005
R63734 VSS.n8616 VSS.n1523 4.5005
R63735 VSS.n8616 VSS.n1541 4.5005
R63736 VSS.n8620 VSS.n1523 4.5005
R63737 VSS.n8620 VSS.n1541 4.5005
R63738 VSS.n8619 VSS.n1523 4.5005
R63739 VSS.n8619 VSS.n1541 4.5005
R63740 VSS.n8608 VSS.n1523 4.5005
R63741 VSS.n8633 VSS.n8608 4.5005
R63742 VSS.n8608 VSS.n1541 4.5005
R63743 VSS.n8635 VSS.n1539 4.5005
R63744 VSS.n1539 VSS.n1523 4.5005
R63745 VSS.n8633 VSS.n1539 4.5005
R63746 VSS.n1541 VSS.n1539 4.5005
R63747 VSS.n8635 VSS.n1528 4.5005
R63748 VSS.n1528 VSS.n1523 4.5005
R63749 VSS.n1541 VSS.n1528 4.5005
R63750 VSS.n8622 VSS.n1523 4.5005
R63751 VSS.n8622 VSS.n1541 4.5005
R63752 VSS.n8625 VSS.n1523 4.5005
R63753 VSS.n8625 VSS.n1541 4.5005
R63754 VSS.n8624 VSS.n1523 4.5005
R63755 VSS.n8624 VSS.n1541 4.5005
R63756 VSS.n8628 VSS.n1523 4.5005
R63757 VSS.n8628 VSS.n1541 4.5005
R63758 VSS.n8627 VSS.n1523 4.5005
R63759 VSS.n8627 VSS.n1541 4.5005
R63760 VSS.n8631 VSS.n1523 4.5005
R63761 VSS.n8631 VSS.n1541 4.5005
R63762 VSS.n8630 VSS.n1523 4.5005
R63763 VSS.n8630 VSS.n1541 4.5005
R63764 VSS.n1544 VSS.n1523 4.5005
R63765 VSS.n8633 VSS.n1544 4.5005
R63766 VSS.n1544 VSS.n1541 4.5005
R63767 VSS.n8634 VSS.n1541 4.5005
R63768 VSS.n8634 VSS.n8633 4.5005
R63769 VSS.n8634 VSS.n1523 4.5005
R63770 VSS.n8635 VSS.n8634 4.5005
R63771 VSS.n8163 VSS.n1993 4.5005
R63772 VSS.n1993 VSS.n1979 4.5005
R63773 VSS.n8159 VSS.n1993 4.5005
R63774 VSS.n8159 VSS.n1997 4.5005
R63775 VSS.n8163 VSS.n1997 4.5005
R63776 VSS.n1992 VSS.n1980 4.5005
R63777 VSS.n8163 VSS.n1992 4.5005
R63778 VSS.n1999 VSS.n1980 4.5005
R63779 VSS.n8163 VSS.n1999 4.5005
R63780 VSS.n1991 VSS.n1980 4.5005
R63781 VSS.n8163 VSS.n1991 4.5005
R63782 VSS.n2001 VSS.n1980 4.5005
R63783 VSS.n8163 VSS.n2001 4.5005
R63784 VSS.n1990 VSS.n1980 4.5005
R63785 VSS.n8163 VSS.n1990 4.5005
R63786 VSS.n2003 VSS.n1980 4.5005
R63787 VSS.n8163 VSS.n2003 4.5005
R63788 VSS.n1989 VSS.n1980 4.5005
R63789 VSS.n8163 VSS.n1989 4.5005
R63790 VSS.n2005 VSS.n1980 4.5005
R63791 VSS.n8163 VSS.n2005 4.5005
R63792 VSS.n1988 VSS.n1980 4.5005
R63793 VSS.n8163 VSS.n1988 4.5005
R63794 VSS.n2007 VSS.n1980 4.5005
R63795 VSS.n8163 VSS.n2007 4.5005
R63796 VSS.n1987 VSS.n1980 4.5005
R63797 VSS.n8163 VSS.n1987 4.5005
R63798 VSS.n2009 VSS.n1980 4.5005
R63799 VSS.n8163 VSS.n2009 4.5005
R63800 VSS.n1986 VSS.n1980 4.5005
R63801 VSS.n8163 VSS.n1986 4.5005
R63802 VSS.n2011 VSS.n1980 4.5005
R63803 VSS.n8163 VSS.n2011 4.5005
R63804 VSS.n1985 VSS.n1980 4.5005
R63805 VSS.n8163 VSS.n1985 4.5005
R63806 VSS.n2013 VSS.n1980 4.5005
R63807 VSS.n8163 VSS.n2013 4.5005
R63808 VSS.n1984 VSS.n1980 4.5005
R63809 VSS.n8163 VSS.n1984 4.5005
R63810 VSS.n2015 VSS.n1980 4.5005
R63811 VSS.n8163 VSS.n2015 4.5005
R63812 VSS.n1983 VSS.n1980 4.5005
R63813 VSS.n8163 VSS.n1983 4.5005
R63814 VSS.n8162 VSS.n1980 4.5005
R63815 VSS.n8163 VSS.n8162 4.5005
R63816 VSS.n1982 VSS.n1980 4.5005
R63817 VSS.n8163 VSS.n1982 4.5005
R63818 VSS.n8164 VSS.n1980 4.5005
R63819 VSS.n8164 VSS.n1979 4.5005
R63820 VSS.n8164 VSS.n8163 4.5005
R63821 VSS.n8194 VSS.n8165 4.5005
R63822 VSS.n8198 VSS.n8165 4.5005
R63823 VSS.n8165 VSS.n1949 4.5005
R63824 VSS.n8198 VSS.n8167 4.5005
R63825 VSS.n8167 VSS.n1949 4.5005
R63826 VSS.n8198 VSS.n1977 4.5005
R63827 VSS.n1977 VSS.n1949 4.5005
R63828 VSS.n8198 VSS.n8168 4.5005
R63829 VSS.n8168 VSS.n1949 4.5005
R63830 VSS.n8198 VSS.n1976 4.5005
R63831 VSS.n1976 VSS.n1949 4.5005
R63832 VSS.n8198 VSS.n8169 4.5005
R63833 VSS.n8169 VSS.n1949 4.5005
R63834 VSS.n8198 VSS.n1975 4.5005
R63835 VSS.n1975 VSS.n1949 4.5005
R63836 VSS.n8198 VSS.n8170 4.5005
R63837 VSS.n8170 VSS.n1949 4.5005
R63838 VSS.n8198 VSS.n1974 4.5005
R63839 VSS.n1974 VSS.n1949 4.5005
R63840 VSS.n8198 VSS.n8171 4.5005
R63841 VSS.n8171 VSS.n1949 4.5005
R63842 VSS.n8198 VSS.n1973 4.5005
R63843 VSS.n1973 VSS.n1949 4.5005
R63844 VSS.n8198 VSS.n8172 4.5005
R63845 VSS.n8172 VSS.n1949 4.5005
R63846 VSS.n8198 VSS.n1972 4.5005
R63847 VSS.n1972 VSS.n1949 4.5005
R63848 VSS.n8198 VSS.n8173 4.5005
R63849 VSS.n8173 VSS.n1949 4.5005
R63850 VSS.n8198 VSS.n1971 4.5005
R63851 VSS.n1971 VSS.n1949 4.5005
R63852 VSS.n8198 VSS.n8174 4.5005
R63853 VSS.n8174 VSS.n1949 4.5005
R63854 VSS.n8198 VSS.n1970 4.5005
R63855 VSS.n1970 VSS.n1949 4.5005
R63856 VSS.n8198 VSS.n8175 4.5005
R63857 VSS.n8175 VSS.n1949 4.5005
R63858 VSS.n8198 VSS.n1969 4.5005
R63859 VSS.n1969 VSS.n1949 4.5005
R63860 VSS.n8198 VSS.n8196 4.5005
R63861 VSS.n8196 VSS.n1949 4.5005
R63862 VSS.n8198 VSS.n1968 4.5005
R63863 VSS.n1968 VSS.n1949 4.5005
R63864 VSS.n8198 VSS.n8197 4.5005
R63865 VSS.n8197 VSS.n1949 4.5005
R63866 VSS.n8199 VSS.n8198 4.5005
R63867 VSS.n8199 VSS.n1949 4.5005
R63868 VSS.n8194 VSS.n1966 4.5005
R63869 VSS.n8198 VSS.n1966 4.5005
R63870 VSS.n1966 VSS.n1949 4.5005
R63871 VSS.n8607 VSS.n8606 4.5005
R63872 VSS.n8596 VSS.n8572 4.5005
R63873 VSS.n8592 VSS.n8572 4.5005
R63874 VSS.n8587 VSS.n8586 4.5005
R63875 VSS.n8581 VSS.n8580 4.5005
R63876 VSS.n8585 VSS.n8584 4.5005
R63877 VSS.n8591 VSS.n8590 4.5005
R63878 VSS.n8604 VSS.n8603 4.5005
R63879 VSS.n8080 VSS.n8079 4.5005
R63880 VSS.n8083 VSS.n8079 4.5005
R63881 VSS.n8079 VSS.n1547 4.5005
R63882 VSS.n8086 VSS.n8085 4.5005
R63883 VSS.n5236 VSS.n4331 4.5005
R63884 VSS.n5236 VSS.n4332 4.5005
R63885 VSS.n5245 VSS.n5236 4.5005
R63886 VSS.n4336 VSS.n4332 4.5005
R63887 VSS.n5245 VSS.n4336 4.5005
R63888 VSS.n5239 VSS.n4332 4.5005
R63889 VSS.n5245 VSS.n5239 4.5005
R63890 VSS.n4335 VSS.n4332 4.5005
R63891 VSS.n5245 VSS.n4335 4.5005
R63892 VSS.n5242 VSS.n4332 4.5005
R63893 VSS.n5245 VSS.n5242 4.5005
R63894 VSS.n4334 VSS.n4332 4.5005
R63895 VSS.n5245 VSS.n4334 4.5005
R63896 VSS.n5244 VSS.n4332 4.5005
R63897 VSS.n5244 VSS.n4330 4.5005
R63898 VSS.n5245 VSS.n5244 4.5005
R63899 VSS.n4331 VSS.n4327 4.5005
R63900 VSS.n4332 VSS.n4327 4.5005
R63901 VSS.n4330 VSS.n4327 4.5005
R63902 VSS.n5245 VSS.n4327 4.5005
R63903 VSS.n4331 VSS.n4329 4.5005
R63904 VSS.n4332 VSS.n4329 4.5005
R63905 VSS.n4330 VSS.n4329 4.5005
R63906 VSS.n5245 VSS.n4329 4.5005
R63907 VSS.n5246 VSS.n4331 4.5005
R63908 VSS.n5246 VSS.n4332 4.5005
R63909 VSS.n5246 VSS.n4330 4.5005
R63910 VSS.n5246 VSS.n5245 4.5005
R63911 VSS.n4331 VSS.n4320 4.5005
R63912 VSS.n4332 VSS.n4320 4.5005
R63913 VSS.n4330 VSS.n4320 4.5005
R63914 VSS.n5245 VSS.n4320 4.5005
R63915 VSS.n5303 VSS.n4316 4.5005
R63916 VSS.n4316 VSS.n4313 4.5005
R63917 VSS.n5296 VSS.n4316 4.5005
R63918 VSS.n5300 VSS.n4316 4.5005
R63919 VSS.n5303 VSS.n4315 4.5005
R63920 VSS.n4315 VSS.n4313 4.5005
R63921 VSS.n5296 VSS.n4315 4.5005
R63922 VSS.n5300 VSS.n4315 4.5005
R63923 VSS.n5303 VSS.n4317 4.5005
R63924 VSS.n4317 VSS.n4313 4.5005
R63925 VSS.n5296 VSS.n4317 4.5005
R63926 VSS.n5300 VSS.n4317 4.5005
R63927 VSS.n5303 VSS.n4314 4.5005
R63928 VSS.n4314 VSS.n4313 4.5005
R63929 VSS.n5296 VSS.n4314 4.5005
R63930 VSS.n5300 VSS.n4314 4.5005
R63931 VSS.n5303 VSS.n5264 4.5005
R63932 VSS.n5264 VSS.n4313 4.5005
R63933 VSS.n5300 VSS.n5264 4.5005
R63934 VSS.n5271 VSS.n4313 4.5005
R63935 VSS.n5300 VSS.n5271 4.5005
R63936 VSS.n5298 VSS.n4313 4.5005
R63937 VSS.n5300 VSS.n5298 4.5005
R63938 VSS.n5270 VSS.n4313 4.5005
R63939 VSS.n5300 VSS.n5270 4.5005
R63940 VSS.n5299 VSS.n4313 4.5005
R63941 VSS.n5300 VSS.n5299 4.5005
R63942 VSS.n5301 VSS.n4313 4.5005
R63943 VSS.n5301 VSS.n5300 4.5005
R63944 VSS.n5267 VSS.n4313 4.5005
R63945 VSS.n5296 VSS.n5267 4.5005
R63946 VSS.n5300 VSS.n5267 4.5005
R63947 VSS.n6195 VSS.n3945 4.5005
R63948 VSS.n3951 VSS.n3945 4.5005
R63949 VSS.n6197 VSS.n3945 4.5005
R63950 VSS.n3951 VSS.n3943 4.5005
R63951 VSS.n6197 VSS.n3943 4.5005
R63952 VSS.n3951 VSS.n3946 4.5005
R63953 VSS.n6197 VSS.n3946 4.5005
R63954 VSS.n3951 VSS.n3942 4.5005
R63955 VSS.n6197 VSS.n3942 4.5005
R63956 VSS.n3951 VSS.n3947 4.5005
R63957 VSS.n6197 VSS.n3947 4.5005
R63958 VSS.n6195 VSS.n3941 4.5005
R63959 VSS.n3951 VSS.n3941 4.5005
R63960 VSS.n6197 VSS.n3941 4.5005
R63961 VSS.n6197 VSS.n3948 4.5005
R63962 VSS.n3956 VSS.n3948 4.5005
R63963 VSS.n3951 VSS.n3948 4.5005
R63964 VSS.n6195 VSS.n3948 4.5005
R63965 VSS.n6197 VSS.n3940 4.5005
R63966 VSS.n3956 VSS.n3940 4.5005
R63967 VSS.n3951 VSS.n3940 4.5005
R63968 VSS.n6195 VSS.n3940 4.5005
R63969 VSS.n6197 VSS.n3949 4.5005
R63970 VSS.n3956 VSS.n3949 4.5005
R63971 VSS.n3951 VSS.n3949 4.5005
R63972 VSS.n6195 VSS.n3949 4.5005
R63973 VSS.n6197 VSS.n3939 4.5005
R63974 VSS.n3956 VSS.n3939 4.5005
R63975 VSS.n3951 VSS.n3939 4.5005
R63976 VSS.n6195 VSS.n3939 4.5005
R63977 VSS.n6197 VSS.n6196 4.5005
R63978 VSS.n6196 VSS.n3956 4.5005
R63979 VSS.n6196 VSS.n3951 4.5005
R63980 VSS.n6196 VSS.n6195 4.5005
R63981 VSS.n3377 VSS.n3352 4.5005
R63982 VSS.n6530 VSS.n3352 4.5005
R63983 VSS.n6532 VSS.n3352 4.5005
R63984 VSS.n6530 VSS.n3354 4.5005
R63985 VSS.n6532 VSS.n3354 4.5005
R63986 VSS.n6530 VSS.n3351 4.5005
R63987 VSS.n6532 VSS.n3351 4.5005
R63988 VSS.n6530 VSS.n3355 4.5005
R63989 VSS.n6532 VSS.n3355 4.5005
R63990 VSS.n6530 VSS.n3350 4.5005
R63991 VSS.n6532 VSS.n3350 4.5005
R63992 VSS.n6530 VSS.n3356 4.5005
R63993 VSS.n6532 VSS.n3356 4.5005
R63994 VSS.n6530 VSS.n3349 4.5005
R63995 VSS.n6532 VSS.n3349 4.5005
R63996 VSS.n6530 VSS.n3357 4.5005
R63997 VSS.n6532 VSS.n3357 4.5005
R63998 VSS.n6530 VSS.n3348 4.5005
R63999 VSS.n6532 VSS.n3348 4.5005
R64000 VSS.n6530 VSS.n3358 4.5005
R64001 VSS.n6532 VSS.n3358 4.5005
R64002 VSS.n6530 VSS.n3347 4.5005
R64003 VSS.n6532 VSS.n3347 4.5005
R64004 VSS.n6530 VSS.n3359 4.5005
R64005 VSS.n6532 VSS.n3359 4.5005
R64006 VSS.n6530 VSS.n3346 4.5005
R64007 VSS.n6532 VSS.n3346 4.5005
R64008 VSS.n6530 VSS.n3360 4.5005
R64009 VSS.n6532 VSS.n3360 4.5005
R64010 VSS.n6530 VSS.n3345 4.5005
R64011 VSS.n6532 VSS.n3345 4.5005
R64012 VSS.n6530 VSS.n3361 4.5005
R64013 VSS.n6532 VSS.n3361 4.5005
R64014 VSS.n6530 VSS.n3344 4.5005
R64015 VSS.n6532 VSS.n3344 4.5005
R64016 VSS.n6530 VSS.n3362 4.5005
R64017 VSS.n6532 VSS.n3362 4.5005
R64018 VSS.n6530 VSS.n3343 4.5005
R64019 VSS.n6532 VSS.n3343 4.5005
R64020 VSS.n6530 VSS.n3363 4.5005
R64021 VSS.n6532 VSS.n3363 4.5005
R64022 VSS.n6530 VSS.n3342 4.5005
R64023 VSS.n6532 VSS.n3342 4.5005
R64024 VSS.n6530 VSS.n3364 4.5005
R64025 VSS.n6532 VSS.n3364 4.5005
R64026 VSS.n6530 VSS.n3341 4.5005
R64027 VSS.n6532 VSS.n3341 4.5005
R64028 VSS.n6531 VSS.n3377 4.5005
R64029 VSS.n6531 VSS.n6530 4.5005
R64030 VSS.n6532 VSS.n6531 4.5005
R64031 VSS.n6915 VSS.n2864 4.5005
R64032 VSS.n6918 VSS.n2864 4.5005
R64033 VSS.n2864 VSS.n2851 4.5005
R64034 VSS.n6918 VSS.n2861 4.5005
R64035 VSS.n2861 VSS.n2851 4.5005
R64036 VSS.n6918 VSS.n2866 4.5005
R64037 VSS.n2866 VSS.n2851 4.5005
R64038 VSS.n6918 VSS.n2860 4.5005
R64039 VSS.n2860 VSS.n2851 4.5005
R64040 VSS.n6918 VSS.n2868 4.5005
R64041 VSS.n2868 VSS.n2851 4.5005
R64042 VSS.n6918 VSS.n2859 4.5005
R64043 VSS.n2859 VSS.n2851 4.5005
R64044 VSS.n6918 VSS.n2870 4.5005
R64045 VSS.n2870 VSS.n2851 4.5005
R64046 VSS.n6918 VSS.n2858 4.5005
R64047 VSS.n2858 VSS.n2851 4.5005
R64048 VSS.n6918 VSS.n2872 4.5005
R64049 VSS.n2872 VSS.n2851 4.5005
R64050 VSS.n6918 VSS.n2857 4.5005
R64051 VSS.n2857 VSS.n2851 4.5005
R64052 VSS.n6918 VSS.n6917 4.5005
R64053 VSS.n6917 VSS.n2856 4.5005
R64054 VSS.n6917 VSS.n2851 4.5005
R64055 VSS.n1580 VSS.n1569 4.5005
R64056 VSS.n1580 VSS.n1570 4.5005
R64057 VSS.n8559 VSS.n1580 4.5005
R64058 VSS.n1577 VSS.n1570 4.5005
R64059 VSS.n8559 VSS.n1577 4.5005
R64060 VSS.n1583 VSS.n1570 4.5005
R64061 VSS.n8559 VSS.n1583 4.5005
R64062 VSS.n1576 VSS.n1570 4.5005
R64063 VSS.n8559 VSS.n1576 4.5005
R64064 VSS.n1570 VSS.n1567 4.5005
R64065 VSS.n1568 VSS.n1567 4.5005
R64066 VSS.n8559 VSS.n1567 4.5005
R64067 VSS.n8560 VSS.n1569 4.5005
R64068 VSS.n8560 VSS.n1570 4.5005
R64069 VSS.n8560 VSS.n1568 4.5005
R64070 VSS.n8560 VSS.n8559 4.5005
R64071 VSS.n8559 VSS.n1563 4.5005
R64072 VSS.n1568 VSS.n1563 4.5005
R64073 VSS.n1569 VSS.n1563 4.5005
R64074 VSS.n1574 VSS.n1569 4.5005
R64075 VSS.n8559 VSS.n1574 4.5005
R64076 VSS.n1586 VSS.n1570 4.5005
R64077 VSS.n8559 VSS.n1586 4.5005
R64078 VSS.n1572 VSS.n1570 4.5005
R64079 VSS.n8559 VSS.n1572 4.5005
R64080 VSS.n8558 VSS.n1569 4.5005
R64081 VSS.n8558 VSS.n1570 4.5005
R64082 VSS.n8559 VSS.n8558 4.5005
R64083 VSS.n8088 VSS.n1595 4.5005
R64084 VSS.n2089 VSS.n1595 4.5005
R64085 VSS.n2090 VSS.n1595 4.5005
R64086 VSS.n8088 VSS.n8001 4.5005
R64087 VSS.n8001 VSS.n2089 4.5005
R64088 VSS.n8001 VSS.n2090 4.5005
R64089 VSS.n2125 VSS.n2090 4.5005
R64090 VSS.n2125 VSS.n2091 4.5005
R64091 VSS.n2125 VSS.n2089 4.5005
R64092 VSS.n8088 VSS.n2125 4.5005
R64093 VSS.n8077 VSS.n2090 4.5005
R64094 VSS.n8077 VSS.n2091 4.5005
R64095 VSS.n8088 VSS.n8077 4.5005
R64096 VSS.n8088 VSS.n2124 4.5005
R64097 VSS.n2124 VSS.n2090 4.5005
R64098 VSS.n2122 VSS.n2089 4.5005
R64099 VSS.n2122 VSS.n2090 4.5005
R64100 VSS.n2120 VSS.n2089 4.5005
R64101 VSS.n2120 VSS.n2090 4.5005
R64102 VSS.n2118 VSS.n2089 4.5005
R64103 VSS.n2118 VSS.n2090 4.5005
R64104 VSS.n2116 VSS.n2089 4.5005
R64105 VSS.n2116 VSS.n2090 4.5005
R64106 VSS.n2114 VSS.n2089 4.5005
R64107 VSS.n2114 VSS.n2090 4.5005
R64108 VSS.n2112 VSS.n2089 4.5005
R64109 VSS.n2112 VSS.n2090 4.5005
R64110 VSS.n2110 VSS.n2089 4.5005
R64111 VSS.n2110 VSS.n2090 4.5005
R64112 VSS.n8078 VSS.n2089 4.5005
R64113 VSS.n8078 VSS.n2091 4.5005
R64114 VSS.n8078 VSS.n2090 4.5005
R64115 VSS.n8088 VSS.n8087 4.5005
R64116 VSS.n8087 VSS.n2089 4.5005
R64117 VSS.n8087 VSS.n2091 4.5005
R64118 VSS.n8087 VSS.n2090 4.5005
R64119 VSS.n8088 VSS.n2108 4.5005
R64120 VSS.n2108 VSS.n2089 4.5005
R64121 VSS.n2108 VSS.n2090 4.5005
R64122 VSS.n2106 VSS.n2089 4.5005
R64123 VSS.n2106 VSS.n2090 4.5005
R64124 VSS.n2104 VSS.n2089 4.5005
R64125 VSS.n2104 VSS.n2090 4.5005
R64126 VSS.n2102 VSS.n2089 4.5005
R64127 VSS.n2102 VSS.n2090 4.5005
R64128 VSS.n2100 VSS.n2089 4.5005
R64129 VSS.n2100 VSS.n2090 4.5005
R64130 VSS.n2098 VSS.n2089 4.5005
R64131 VSS.n2098 VSS.n2090 4.5005
R64132 VSS.n2096 VSS.n2089 4.5005
R64133 VSS.n2096 VSS.n2090 4.5005
R64134 VSS.n2094 VSS.n2089 4.5005
R64135 VSS.n2094 VSS.n2090 4.5005
R64136 VSS.n2089 VSS.n2086 4.5005
R64137 VSS.n2091 VSS.n2086 4.5005
R64138 VSS.n2090 VSS.n2086 4.5005
R64139 VSS.n8089 VSS.n2090 4.5005
R64140 VSS.n8089 VSS.n2091 4.5005
R64141 VSS.n8089 VSS.n2089 4.5005
R64142 VSS.n8089 VSS.n8088 4.5005
R64143 VSS.n8101 VSS.n8097 4.5005
R64144 VSS.n8097 VSS.n2035 4.5005
R64145 VSS.n8097 VSS.n2031 4.5005
R64146 VSS.n8100 VSS.n2031 4.5005
R64147 VSS.n8101 VSS.n8100 4.5005
R64148 VSS.n8103 VSS.n2046 4.5005
R64149 VSS.n8101 VSS.n2046 4.5005
R64150 VSS.n8103 VSS.n2051 4.5005
R64151 VSS.n8101 VSS.n2051 4.5005
R64152 VSS.n8103 VSS.n2045 4.5005
R64153 VSS.n8101 VSS.n2045 4.5005
R64154 VSS.n8103 VSS.n2054 4.5005
R64155 VSS.n8101 VSS.n2054 4.5005
R64156 VSS.n8103 VSS.n2044 4.5005
R64157 VSS.n8101 VSS.n2044 4.5005
R64158 VSS.n8103 VSS.n2057 4.5005
R64159 VSS.n8101 VSS.n2057 4.5005
R64160 VSS.n8103 VSS.n2043 4.5005
R64161 VSS.n8101 VSS.n2043 4.5005
R64162 VSS.n8103 VSS.n2060 4.5005
R64163 VSS.n8101 VSS.n2060 4.5005
R64164 VSS.n8103 VSS.n2042 4.5005
R64165 VSS.n8101 VSS.n2042 4.5005
R64166 VSS.n8103 VSS.n2063 4.5005
R64167 VSS.n8101 VSS.n2063 4.5005
R64168 VSS.n8103 VSS.n2041 4.5005
R64169 VSS.n8101 VSS.n2041 4.5005
R64170 VSS.n8103 VSS.n2066 4.5005
R64171 VSS.n8101 VSS.n2066 4.5005
R64172 VSS.n8103 VSS.n2040 4.5005
R64173 VSS.n8101 VSS.n2040 4.5005
R64174 VSS.n8103 VSS.n2069 4.5005
R64175 VSS.n8101 VSS.n2069 4.5005
R64176 VSS.n8103 VSS.n2039 4.5005
R64177 VSS.n8101 VSS.n2039 4.5005
R64178 VSS.n8103 VSS.n2072 4.5005
R64179 VSS.n8101 VSS.n2072 4.5005
R64180 VSS.n8103 VSS.n2038 4.5005
R64181 VSS.n8101 VSS.n2038 4.5005
R64182 VSS.n8103 VSS.n2075 4.5005
R64183 VSS.n8101 VSS.n2075 4.5005
R64184 VSS.n8103 VSS.n2037 4.5005
R64185 VSS.n8101 VSS.n2037 4.5005
R64186 VSS.n8103 VSS.n2078 4.5005
R64187 VSS.n8101 VSS.n2078 4.5005
R64188 VSS.n8103 VSS.n2036 4.5005
R64189 VSS.n8101 VSS.n2036 4.5005
R64190 VSS.n8103 VSS.n8102 4.5005
R64191 VSS.n8102 VSS.n2035 4.5005
R64192 VSS.n8102 VSS.n8101 4.5005
R64193 VSS.n8224 VSS.n1909 4.5005
R64194 VSS.n8228 VSS.n1909 4.5005
R64195 VSS.n1909 VSS.n1880 4.5005
R64196 VSS.n8228 VSS.n1911 4.5005
R64197 VSS.n1911 VSS.n1880 4.5005
R64198 VSS.n8228 VSS.n1908 4.5005
R64199 VSS.n1908 VSS.n1880 4.5005
R64200 VSS.n8228 VSS.n1912 4.5005
R64201 VSS.n1912 VSS.n1880 4.5005
R64202 VSS.n8228 VSS.n1907 4.5005
R64203 VSS.n1907 VSS.n1880 4.5005
R64204 VSS.n8228 VSS.n1913 4.5005
R64205 VSS.n1913 VSS.n1880 4.5005
R64206 VSS.n8228 VSS.n1906 4.5005
R64207 VSS.n1906 VSS.n1880 4.5005
R64208 VSS.n8228 VSS.n1914 4.5005
R64209 VSS.n1914 VSS.n1880 4.5005
R64210 VSS.n8228 VSS.n1905 4.5005
R64211 VSS.n1905 VSS.n1880 4.5005
R64212 VSS.n8228 VSS.n1915 4.5005
R64213 VSS.n1915 VSS.n1880 4.5005
R64214 VSS.n8228 VSS.n1904 4.5005
R64215 VSS.n1904 VSS.n1880 4.5005
R64216 VSS.n8228 VSS.n1916 4.5005
R64217 VSS.n1916 VSS.n1880 4.5005
R64218 VSS.n8228 VSS.n1903 4.5005
R64219 VSS.n1903 VSS.n1880 4.5005
R64220 VSS.n8228 VSS.n1917 4.5005
R64221 VSS.n1917 VSS.n1880 4.5005
R64222 VSS.n8228 VSS.n1902 4.5005
R64223 VSS.n1902 VSS.n1880 4.5005
R64224 VSS.n8228 VSS.n1918 4.5005
R64225 VSS.n1918 VSS.n1880 4.5005
R64226 VSS.n8228 VSS.n1901 4.5005
R64227 VSS.n1901 VSS.n1880 4.5005
R64228 VSS.n8228 VSS.n1919 4.5005
R64229 VSS.n1919 VSS.n1880 4.5005
R64230 VSS.n8228 VSS.n1900 4.5005
R64231 VSS.n1900 VSS.n1880 4.5005
R64232 VSS.n8228 VSS.n8226 4.5005
R64233 VSS.n8226 VSS.n1880 4.5005
R64234 VSS.n8228 VSS.n1899 4.5005
R64235 VSS.n1899 VSS.n1880 4.5005
R64236 VSS.n8228 VSS.n8227 4.5005
R64237 VSS.n8227 VSS.n1880 4.5005
R64238 VSS.n8229 VSS.n8228 4.5005
R64239 VSS.n8229 VSS.n1880 4.5005
R64240 VSS.n8224 VSS.n1897 4.5005
R64241 VSS.n8228 VSS.n1897 4.5005
R64242 VSS.n1897 VSS.n1880 4.5005
R64243 VSS.n8548 VSS.n8547 4.5005
R64244 VSS.n8547 VSS.n8546 4.5005
R64245 VSS.n8810 VSS.n8809 4.5005
R64246 VSS.n8840 VSS.n1345 4.5005
R64247 VSS.n8840 VSS.n8839 4.5005
R64248 VSS.n8836 VSS.n1305 4.5005
R64249 VSS.n8831 VSS.n1305 4.5005
R64250 VSS.n8831 VSS.n1349 4.5005
R64251 VSS.n8836 VSS.n1349 4.5005
R64252 VSS.n8838 VSS.n1349 4.5005
R64253 VSS.n8839 VSS.n1348 4.5005
R64254 VSS.n1348 VSS.n1345 4.5005
R64255 VSS.n8808 VSS.n1348 4.5005
R64256 VSS.n8809 VSS.n1389 4.5005
R64257 VSS.n1613 VSS.n1389 4.5005
R64258 VSS.n8546 VSS.n1596 4.5005
R64259 VSS.n8548 VSS.n1596 4.5005
R64260 VSS.n8550 VSS.n1596 4.5005
R64261 VSS.n8551 VSS.n1590 4.5005
R64262 VSS.n8837 VSS.n8836 4.5005
R64263 VSS.n8838 VSS.n8837 4.5005
R64264 VSS.n8807 VSS.n1345 4.5005
R64265 VSS.n8808 VSS.n8807 4.5005
R64266 VSS.n1613 VSS.n1612 4.5005
R64267 VSS.n8549 VSS.n8548 4.5005
R64268 VSS.n8550 VSS.n8549 4.5005
R64269 VSS.n8554 VSS.n8551 4.5005
R64270 VSS.n8554 VSS.n1594 4.5005
R64271 VSS.n8554 VSS.n8553 4.5005
R64272 VSS.n8555 VSS.n8554 4.5005
R64273 VSS.n8072 VSS.n8004 4.5005
R64274 VSS.n8072 VSS.n8071 4.5005
R64275 VSS.n8068 VSS.n8067 4.5005
R64276 VSS.n8067 VSS.n8066 4.5005
R64277 VSS.n8054 VSS.n8053 4.5005
R64278 VSS.n8049 VSS.n8048 4.5005
R64279 VSS.n8048 VSS.n8047 4.5005
R64280 VSS.n8044 VSS.n8043 4.5005
R64281 VSS.n8043 VSS.n8042 4.5005
R64282 VSS.n8042 VSS.n8033 4.5005
R64283 VSS.n8046 VSS.n8033 4.5005
R64284 VSS.n8047 VSS.n8026 4.5005
R64285 VSS.n8051 VSS.n8026 4.5005
R64286 VSS.n8054 VSS.n8022 4.5005
R64287 VSS.n8024 VSS.n8022 4.5005
R64288 VSS.n8057 VSS.n8022 4.5005
R64289 VSS.n8066 VSS.n8011 4.5005
R64290 VSS.n8070 VSS.n8011 4.5005
R64291 VSS.n8071 VSS.n8008 4.5005
R64292 VSS.n8074 VSS.n8008 4.5005
R64293 VSS.n8045 VSS.n8044 4.5005
R64294 VSS.n8045 VSS.n8035 4.5005
R64295 VSS.n8046 VSS.n8045 4.5005
R64296 VSS.n8050 VSS.n8049 4.5005
R64297 VSS.n8050 VSS.n8028 4.5005
R64298 VSS.n8051 VSS.n8050 4.5005
R64299 VSS.n8056 VSS.n8024 4.5005
R64300 VSS.n8057 VSS.n8056 4.5005
R64301 VSS.n8069 VSS.n8068 4.5005
R64302 VSS.n8069 VSS.n8013 4.5005
R64303 VSS.n8070 VSS.n8069 4.5005
R64304 VSS.n8075 VSS.n8004 4.5005
R64305 VSS.n8075 VSS.n8002 4.5005
R64306 VSS.n8075 VSS.n8074 4.5005
R64307 VSS.n8561 VSS.n1565 4.5005
R64308 VSS.n8404 VSS.n8403 4.5005
R64309 VSS.n8822 VSS.n1365 4.5005
R64310 VSS.n1365 VSS.n1321 4.5005
R64311 VSS.n8849 VSS.n1315 4.5005
R64312 VSS.n8854 VSS.n1312 4.5005
R64313 VSS.n8851 VSS.n1313 4.5005
R64314 VSS.n8856 VSS.n8851 4.5005
R64315 VSS.n8844 VSS.n1320 4.5005
R64316 VSS.n8847 VSS.n8844 4.5005
R64317 VSS.n8822 VSS.n1363 4.5005
R64318 VSS.n8392 VSS.n8390 4.5005
R64319 VSS.n8392 VSS.n8391 4.5005
R64320 VSS.n8563 VSS.n1559 4.5005
R64321 VSS.n8565 VSS.n1559 4.5005
R64322 VSS.n8857 VSS.n1312 4.5005
R64323 VSS.n8857 VSS.n1311 4.5005
R64324 VSS.n8857 VSS.n1313 4.5005
R64325 VSS.n8857 VSS.n8856 4.5005
R64326 VSS.n8849 VSS.n8848 4.5005
R64327 VSS.n8848 VSS.n1317 4.5005
R64328 VSS.n8848 VSS.n1320 4.5005
R64329 VSS.n8848 VSS.n8847 4.5005
R64330 VSS.n8821 VSS.n1321 4.5005
R64331 VSS.n8821 VSS.n8820 4.5005
R64332 VSS.n8822 VSS.n8821 4.5005
R64333 VSS.n8403 VSS.n1662 4.5005
R64334 VSS.n8387 VSS.n1662 4.5005
R64335 VSS.n8390 VSS.n1662 4.5005
R64336 VSS.n8391 VSS.n1662 4.5005
R64337 VSS.n8564 VSS.n1565 4.5005
R64338 VSS.n8564 VSS.n1562 4.5005
R64339 VSS.n8564 VSS.n8563 4.5005
R64340 VSS.n8565 VSS.n8564 4.5005
R64341 VSS.n7126 VSS.n2589 4.5005
R64342 VSS.n7126 VSS.n7125 4.5005
R64343 VSS.n7119 VSS.n2505 4.5005
R64344 VSS.n7117 VSS.n2505 4.5005
R64345 VSS.n7109 VSS.n7108 4.5005
R64346 VSS.n7104 VSS.n7102 4.5005
R64347 VSS.n7102 VSS.n7054 4.5005
R64348 VSS.n7050 VSS.n7048 4.5005
R64349 VSS.n7048 VSS.n2608 4.5005
R64350 VSS.n7052 VSS.n2608 4.5005
R64351 VSS.n7053 VSS.n7052 4.5005
R64352 VSS.n7106 VSS.n7054 4.5005
R64353 VSS.n7107 VSS.n7106 4.5005
R64354 VSS.n7108 VSS.n1377 4.5005
R64355 VSS.n2598 VSS.n1377 4.5005
R64356 VSS.n7111 VSS.n1377 4.5005
R64357 VSS.n7121 VSS.n7117 4.5005
R64358 VSS.n7122 VSS.n7121 4.5005
R64359 VSS.n7125 VSS.n7124 4.5005
R64360 VSS.n7124 VSS.n1557 4.5005
R64361 VSS.n7116 VSS.n7115 4.5005
R64362 VSS.n7115 VSS.n2596 4.5005
R64363 VSS.n7115 VSS.n7114 4.5005
R64364 VSS.n7114 VSS.n7113 4.5005
R64365 VSS.n8602 VSS.n1549 4.5005
R64366 VSS.n8598 VSS.n1549 4.5005
R64367 VSS.n8402 VSS.n8396 4.5005
R64368 VSS.n8396 VSS.n1362 4.5005
R64369 VSS.n8402 VSS.n8394 4.5005
R64370 VSS.n8401 VSS.n1362 4.5005
R64371 VSS.n8401 VSS.n8400 4.5005
R64372 VSS.n8402 VSS.n8401 4.5005
R64373 VSS.n8542 VSS.n8541 4.5005
R64374 VSS.n8542 VSS.n1604 4.5005
R64375 VSS.n8545 VSS.n1604 4.5005
R64376 VSS.n8545 VSS.n8544 4.5005
R64377 VSS.n8062 VSS.n8061 4.5005
R64378 VSS.n8062 VSS.n8018 4.5005
R64379 VSS.n8020 VSS.n8018 4.5005
R64380 VSS.n8065 VSS.n8018 4.5005
R64381 VSS.n8064 VSS.n8020 4.5005
R64382 VSS.n8065 VSS.n8064 4.5005
R64383 VSS.n7267 VSS.n7266 4.5005
R64384 VSS.n7266 VSS.n7265 4.5005
R64385 VSS.n7265 VSS.n2477 4.5005
R64386 VSS.n7265 VSS.n7264 4.5005
R64387 VSS.n7072 VSS.n7071 4.5005
R64388 VSS.n7233 VSS.n2515 4.5005
R64389 VSS.n7233 VSS.n7232 4.5005
R64390 VSS.n7232 VSS.n2518 4.5005
R64391 VSS.n7201 VSS.n7184 4.5005
R64392 VSS.n7204 VSS.n7184 4.5005
R64393 VSS.n7204 VSS.n7182 4.5005
R64394 VSS.n7179 VSS.n7178 4.5005
R64395 VSS.n7180 VSS.n7179 4.5005
R64396 VSS.n7180 VSS.n2478 4.5005
R64397 VSS.n7181 VSS.n7180 4.5005
R64398 VSS.n7204 VSS.n7203 4.5005
R64399 VSS.n7232 VSS.n2513 4.5005
R64400 VSS.n7072 VSS.n2594 4.5005
R64401 VSS.n7069 VSS.n2594 4.5005
R64402 VSS.n7068 VSS.n2594 4.5005
R64403 VSS.n7001 VSS.n7000 4.5005
R64404 VSS.n2652 VSS.n2651 4.5005
R64405 VSS.n6823 VSS.n6822 4.5005
R64406 VSS.n6824 VSS.n6817 4.5005
R64407 VSS.n6826 VSS.n6825 4.5005
R64408 VSS.n6827 VSS.n6816 4.5005
R64409 VSS.n6829 VSS.n6828 4.5005
R64410 VSS.n6830 VSS.n6811 4.5005
R64411 VSS.n6832 VSS.n6831 4.5005
R64412 VSS.n6833 VSS.n6810 4.5005
R64413 VSS.n6835 VSS.n6834 4.5005
R64414 VSS.n6836 VSS.n2937 4.5005
R64415 VSS.n6838 VSS.n6837 4.5005
R64416 VSS.n2938 VSS.n2936 4.5005
R64417 VSS.n6802 VSS.n6801 4.5005
R64418 VSS.n6800 VSS.n6799 4.5005
R64419 VSS.n6798 VSS.n6797 4.5005
R64420 VSS.n6795 VSS.n6794 4.5005
R64421 VSS.n6792 VSS.n6791 4.5005
R64422 VSS.n6790 VSS.n6787 4.5005
R64423 VSS.n6786 VSS.n6785 4.5005
R64424 VSS.n6783 VSS.n6782 4.5005
R64425 VSS.n6780 VSS.n6779 4.5005
R64426 VSS.n6777 VSS.n6776 4.5005
R64427 VSS.n6774 VSS.n6773 4.5005
R64428 VSS.n6772 VSS.n2954 4.5005
R64429 VSS.n6771 VSS.n6770 4.5005
R64430 VSS.n2957 VSS.n2956 4.5005
R64431 VSS.n5884 VSS.n5733 4.5005
R64432 VSS.n5883 VSS.n5882 4.5005
R64433 VSS.n5801 VSS.n5800 4.5005
R64434 VSS.n5875 VSS.n5874 4.5005
R64435 VSS.n5873 VSS.n5803 4.5005
R64436 VSS.n5872 VSS.n5871 4.5005
R64437 VSS.n5805 VSS.n5804 4.5005
R64438 VSS.n5867 VSS.n5866 4.5005
R64439 VSS.n5865 VSS.n5807 4.5005
R64440 VSS.n5864 VSS.n5863 4.5005
R64441 VSS.n5809 VSS.n5808 4.5005
R64442 VSS.n5859 VSS.n5858 4.5005
R64443 VSS.n5857 VSS.n5856 4.5005
R64444 VSS.n5855 VSS.n5811 4.5005
R64445 VSS.n5849 VSS.n5812 4.5005
R64446 VSS.n5851 VSS.n5850 4.5005
R64447 VSS.n5848 VSS.n5814 4.5005
R64448 VSS.n5847 VSS.n5846 4.5005
R64449 VSS.n5816 VSS.n5815 4.5005
R64450 VSS.n5842 VSS.n5841 4.5005
R64451 VSS.n5840 VSS.n5818 4.5005
R64452 VSS.n5839 VSS.n5838 4.5005
R64453 VSS.n5820 VSS.n5819 4.5005
R64454 VSS.n5834 VSS.n5833 4.5005
R64455 VSS.n5832 VSS.n5822 4.5005
R64456 VSS.n5831 VSS.n5830 4.5005
R64457 VSS.n5824 VSS.n5823 4.5005
R64458 VSS.n5826 VSS.n5825 4.5005
R64459 VSS.n6612 VSS.n6611 4.5005
R64460 VSS.n3167 VSS.n3162 4.5005
R64461 VSS.n3748 VSS.n3747 4.5005
R64462 VSS.n3750 VSS.n3749 4.5005
R64463 VSS.n3752 VSS.n3751 4.5005
R64464 VSS.n3754 VSS.n3753 4.5005
R64465 VSS.n3756 VSS.n3755 4.5005
R64466 VSS.n3758 VSS.n3757 4.5005
R64467 VSS.n3760 VSS.n3759 4.5005
R64468 VSS.n3762 VSS.n3761 4.5005
R64469 VSS.n3764 VSS.n3763 4.5005
R64470 VSS.n3766 VSS.n3765 4.5005
R64471 VSS.n3768 VSS.n3767 4.5005
R64472 VSS.n3770 VSS.n3769 4.5005
R64473 VSS.n3772 VSS.n3771 4.5005
R64474 VSS.n3774 VSS.n3773 4.5005
R64475 VSS.n3776 VSS.n3775 4.5005
R64476 VSS.n3778 VSS.n3777 4.5005
R64477 VSS.n3780 VSS.n3779 4.5005
R64478 VSS.n3782 VSS.n3781 4.5005
R64479 VSS.n3784 VSS.n3783 4.5005
R64480 VSS.n3786 VSS.n3785 4.5005
R64481 VSS.n3788 VSS.n3787 4.5005
R64482 VSS.n3790 VSS.n3789 4.5005
R64483 VSS.n3792 VSS.n3791 4.5005
R64484 VSS.n3794 VSS.n3793 4.5005
R64485 VSS.n3795 VSS.n3720 4.5005
R64486 VSS.n3797 VSS.n3796 4.5005
R64487 VSS.n6309 VSS.n6308 4.5005
R64488 VSS.n3714 VSS.n3713 4.5005
R64489 VSS.n5997 VSS.n5993 4.5005
R64490 VSS.n5999 VSS.n5998 4.5005
R64491 VSS.n6000 VSS.n5992 4.5005
R64492 VSS.n6002 VSS.n6001 4.5005
R64493 VSS.n6003 VSS.n5987 4.5005
R64494 VSS.n6005 VSS.n6004 4.5005
R64495 VSS.n6006 VSS.n5986 4.5005
R64496 VSS.n6008 VSS.n6007 4.5005
R64497 VSS.n6009 VSS.n5981 4.5005
R64498 VSS.n6011 VSS.n6010 4.5005
R64499 VSS.n6012 VSS.n5980 4.5005
R64500 VSS.n6014 VSS.n6013 4.5005
R64501 VSS.n6015 VSS.n5975 4.5005
R64502 VSS.n6017 VSS.n6016 4.5005
R64503 VSS.n6018 VSS.n5974 4.5005
R64504 VSS.n6020 VSS.n6019 4.5005
R64505 VSS.n6021 VSS.n5969 4.5005
R64506 VSS.n6023 VSS.n6022 4.5005
R64507 VSS.n6024 VSS.n5968 4.5005
R64508 VSS.n6026 VSS.n6025 4.5005
R64509 VSS.n6027 VSS.n5963 4.5005
R64510 VSS.n6029 VSS.n6028 4.5005
R64511 VSS.n6030 VSS.n5962 4.5005
R64512 VSS.n6032 VSS.n6031 4.5005
R64513 VSS.n6033 VSS.n5901 4.5005
R64514 VSS.n6035 VSS.n6034 4.5005
R64515 VSS.n6082 VSS.n4068 4.5005
R64516 VSS.n6084 VSS.n6083 4.5005
R64517 VSS.n6085 VSS.n4063 4.5005
R64518 VSS.n6087 VSS.n6086 4.5005
R64519 VSS.n6088 VSS.n4062 4.5005
R64520 VSS.n6090 VSS.n6089 4.5005
R64521 VSS.n6091 VSS.n4057 4.5005
R64522 VSS.n6093 VSS.n6092 4.5005
R64523 VSS.n6094 VSS.n4056 4.5005
R64524 VSS.n6096 VSS.n6095 4.5005
R64525 VSS.n6097 VSS.n4051 4.5005
R64526 VSS.n6099 VSS.n6098 4.5005
R64527 VSS.n6100 VSS.n4050 4.5005
R64528 VSS.n6102 VSS.n6101 4.5005
R64529 VSS.n6103 VSS.n4045 4.5005
R64530 VSS.n6105 VSS.n6104 4.5005
R64531 VSS.n6106 VSS.n4044 4.5005
R64532 VSS.n6108 VSS.n6107 4.5005
R64533 VSS.n6109 VSS.n4039 4.5005
R64534 VSS.n6111 VSS.n6110 4.5005
R64535 VSS.n6112 VSS.n4038 4.5005
R64536 VSS.n6114 VSS.n6113 4.5005
R64537 VSS.n6115 VSS.n4033 4.5005
R64538 VSS.n6117 VSS.n6116 4.5005
R64539 VSS.n6118 VSS.n4032 4.5005
R64540 VSS.n6120 VSS.n6119 4.5005
R64541 VSS.n6121 VSS.n4028 4.5005
R64542 VSS.n6123 VSS.n6122 4.5005
R64543 VSS.n4075 VSS.n4074 4.5005
R64544 VSS.n5716 VSS.n5715 4.5005
R64545 VSS.n5714 VSS.n5713 4.5005
R64546 VSS.n5712 VSS.n5711 4.5005
R64547 VSS.n5709 VSS.n5708 4.5005
R64548 VSS.n5707 VSS.n4224 4.5005
R64549 VSS.n5706 VSS.n5705 4.5005
R64550 VSS.n4227 VSS.n4226 4.5005
R64551 VSS.n5700 VSS.n5699 4.5005
R64552 VSS.n5698 VSS.n4229 4.5005
R64553 VSS.n5697 VSS.n5696 4.5005
R64554 VSS.n4231 VSS.n4230 4.5005
R64555 VSS.n5692 VSS.n5691 4.5005
R64556 VSS.n5690 VSS.n4233 4.5005
R64557 VSS.n5689 VSS.n5688 4.5005
R64558 VSS.n4235 VSS.n4234 4.5005
R64559 VSS.n5684 VSS.n5683 4.5005
R64560 VSS.n5682 VSS.n4237 4.5005
R64561 VSS.n5681 VSS.n5680 4.5005
R64562 VSS.n4239 VSS.n4238 4.5005
R64563 VSS.n5676 VSS.n5675 4.5005
R64564 VSS.n5674 VSS.n4241 4.5005
R64565 VSS.n5673 VSS.n5672 4.5005
R64566 VSS.n4263 VSS.n4243 4.5005
R64567 VSS.n5666 VSS.n5665 4.5005
R64568 VSS.n4266 VSS.n4260 4.5005
R64569 VSS.n5661 VSS.n5660 4.5005
R64570 VSS.n5658 VSS.n5656 4.5005
R64571 VSS.n4925 VSS.n4924 4.5005
R64572 VSS.n4926 VSS.n4911 4.5005
R64573 VSS.n4928 VSS.n4927 4.5005
R64574 VSS.n4929 VSS.n4906 4.5005
R64575 VSS.n4931 VSS.n4930 4.5005
R64576 VSS.n4932 VSS.n4905 4.5005
R64577 VSS.n4934 VSS.n4933 4.5005
R64578 VSS.n4935 VSS.n4900 4.5005
R64579 VSS.n4937 VSS.n4936 4.5005
R64580 VSS.n4938 VSS.n4899 4.5005
R64581 VSS.n4940 VSS.n4939 4.5005
R64582 VSS.n4941 VSS.n4894 4.5005
R64583 VSS.n4943 VSS.n4942 4.5005
R64584 VSS.n4944 VSS.n4893 4.5005
R64585 VSS.n4946 VSS.n4945 4.5005
R64586 VSS.n4947 VSS.n4888 4.5005
R64587 VSS.n4949 VSS.n4948 4.5005
R64588 VSS.n4950 VSS.n4887 4.5005
R64589 VSS.n4952 VSS.n4951 4.5005
R64590 VSS.n4953 VSS.n4882 4.5005
R64591 VSS.n4955 VSS.n4954 4.5005
R64592 VSS.n4956 VSS.n4881 4.5005
R64593 VSS.n4958 VSS.n4957 4.5005
R64594 VSS.n4959 VSS.n4876 4.5005
R64595 VSS.n4961 VSS.n4960 4.5005
R64596 VSS.n4962 VSS.n4875 4.5005
R64597 VSS.n4964 VSS.n4963 4.5005
R64598 VSS.n4965 VSS.n4507 4.5005
R64599 VSS.n4865 VSS.n4864 4.5005
R64600 VSS.n4863 VSS.n4862 4.5005
R64601 VSS.n4861 VSS.n4860 4.5005
R64602 VSS.n4492 VSS.n4490 4.5005
R64603 VSS.n5087 VSS.n5086 4.5005
R64604 VSS.n5089 VSS.n5088 4.5005
R64605 VSS.n5090 VSS.n4485 4.5005
R64606 VSS.n5092 VSS.n5091 4.5005
R64607 VSS.n5093 VSS.n4480 4.5005
R64608 VSS.n5095 VSS.n5094 4.5005
R64609 VSS.n5096 VSS.n4479 4.5005
R64610 VSS.n5098 VSS.n5097 4.5005
R64611 VSS.n5099 VSS.n4474 4.5005
R64612 VSS.n5101 VSS.n5100 4.5005
R64613 VSS.n5102 VSS.n4473 4.5005
R64614 VSS.n5104 VSS.n5103 4.5005
R64615 VSS.n5105 VSS.n4468 4.5005
R64616 VSS.n5107 VSS.n5106 4.5005
R64617 VSS.n5108 VSS.n4467 4.5005
R64618 VSS.n5110 VSS.n5109 4.5005
R64619 VSS.n5111 VSS.n4462 4.5005
R64620 VSS.n5113 VSS.n5112 4.5005
R64621 VSS.n5114 VSS.n4461 4.5005
R64622 VSS.n5116 VSS.n5115 4.5005
R64623 VSS.n5118 VSS.n5117 4.5005
R64624 VSS.n5120 VSS.n5119 4.5005
R64625 VSS.n5122 VSS.n5121 4.5005
R64626 VSS.n5124 VSS.n5123 4.5005
R64627 VSS.n4493 VSS.n4486 4.5005
R64628 VSS.n4491 VSS.n4486 4.5005
R64629 VSS.n5084 VSS.n4486 4.5005
R64630 VSS.n5085 VSS.n4493 4.5005
R64631 VSS.n5085 VSS.n4491 4.5005
R64632 VSS.n5085 VSS.n5084 4.5005
R64633 VSS.n4500 VSS.n4493 4.5005
R64634 VSS.n4500 VSS.n4491 4.5005
R64635 VSS.n5084 VSS.n4500 4.5005
R64636 VSS.n4498 VSS.n4493 4.5005
R64637 VSS.n4498 VSS.n4491 4.5005
R64638 VSS.n5084 VSS.n4498 4.5005
R64639 VSS.n4501 VSS.n4493 4.5005
R64640 VSS.n4501 VSS.n4491 4.5005
R64641 VSS.n5084 VSS.n4501 4.5005
R64642 VSS.n4497 VSS.n4493 4.5005
R64643 VSS.n5084 VSS.n4497 4.5005
R64644 VSS.n4503 VSS.n4493 4.5005
R64645 VSS.n5084 VSS.n4503 4.5005
R64646 VSS.n4496 VSS.n4493 4.5005
R64647 VSS.n4496 VSS.n4491 4.5005
R64648 VSS.n5084 VSS.n4496 4.5005
R64649 VSS.n4504 VSS.n4493 4.5005
R64650 VSS.n4504 VSS.n4491 4.5005
R64651 VSS.n5084 VSS.n4504 4.5005
R64652 VSS.n4495 VSS.n4493 4.5005
R64653 VSS.n4495 VSS.n4491 4.5005
R64654 VSS.n5084 VSS.n4495 4.5005
R64655 VSS.n5083 VSS.n4493 4.5005
R64656 VSS.n5083 VSS.n4491 4.5005
R64657 VSS.n5084 VSS.n5083 4.5005
R64658 VSS.n4272 VSS.n4264 4.5005
R64659 VSS.n4272 VSS.n4262 4.5005
R64660 VSS.n5663 VSS.n4272 4.5005
R64661 VSS.n4270 VSS.n4264 4.5005
R64662 VSS.n4270 VSS.n4262 4.5005
R64663 VSS.n5663 VSS.n4270 4.5005
R64664 VSS.n4273 VSS.n4264 4.5005
R64665 VSS.n4273 VSS.n4262 4.5005
R64666 VSS.n5663 VSS.n4273 4.5005
R64667 VSS.n4269 VSS.n4264 4.5005
R64668 VSS.n4269 VSS.n4262 4.5005
R64669 VSS.n5663 VSS.n4269 4.5005
R64670 VSS.n5655 VSS.n4264 4.5005
R64671 VSS.n5663 VSS.n5655 4.5005
R64672 VSS.n4268 VSS.n4264 4.5005
R64673 VSS.n5663 VSS.n4268 4.5005
R64674 VSS.n5662 VSS.n4264 4.5005
R64675 VSS.n5662 VSS.n4262 4.5005
R64676 VSS.n5663 VSS.n5662 4.5005
R64677 VSS.n4267 VSS.n4264 4.5005
R64678 VSS.n4267 VSS.n4262 4.5005
R64679 VSS.n5663 VSS.n4267 4.5005
R64680 VSS.n4264 VSS.n4261 4.5005
R64681 VSS.n4262 VSS.n4261 4.5005
R64682 VSS.n5663 VSS.n4261 4.5005
R64683 VSS.n5664 VSS.n4264 4.5005
R64684 VSS.n5664 VSS.n4262 4.5005
R64685 VSS.n5664 VSS.n5663 4.5005
R64686 VSS.n4264 VSS.n4242 4.5005
R64687 VSS.n4262 VSS.n4242 4.5005
R64688 VSS.n5663 VSS.n4242 4.5005
R64689 VSS.n6125 VSS.n4021 4.5005
R64690 VSS.n4021 VSS.n4014 4.5005
R64691 VSS.n4021 VSS.n4009 4.5005
R64692 VSS.n6125 VSS.n4019 4.5005
R64693 VSS.n4019 VSS.n4014 4.5005
R64694 VSS.n4019 VSS.n4009 4.5005
R64695 VSS.n6125 VSS.n4022 4.5005
R64696 VSS.n4022 VSS.n4014 4.5005
R64697 VSS.n4022 VSS.n4009 4.5005
R64698 VSS.n6125 VSS.n4018 4.5005
R64699 VSS.n4018 VSS.n4014 4.5005
R64700 VSS.n4018 VSS.n4009 4.5005
R64701 VSS.n6125 VSS.n4024 4.5005
R64702 VSS.n4024 VSS.n4009 4.5005
R64703 VSS.n6125 VSS.n4017 4.5005
R64704 VSS.n4017 VSS.n4009 4.5005
R64705 VSS.n4025 VSS.n4009 4.5005
R64706 VSS.n4025 VSS.n4014 4.5005
R64707 VSS.n6125 VSS.n4025 4.5005
R64708 VSS.n4016 VSS.n4009 4.5005
R64709 VSS.n4016 VSS.n4014 4.5005
R64710 VSS.n6125 VSS.n4016 4.5005
R64711 VSS.n4026 VSS.n4009 4.5005
R64712 VSS.n4026 VSS.n4014 4.5005
R64713 VSS.n6125 VSS.n4026 4.5005
R64714 VSS.n4015 VSS.n4009 4.5005
R64715 VSS.n4015 VSS.n4014 4.5005
R64716 VSS.n6125 VSS.n4015 4.5005
R64717 VSS.n6124 VSS.n4009 4.5005
R64718 VSS.n6124 VSS.n4014 4.5005
R64719 VSS.n6125 VSS.n6124 4.5005
R64720 VSS.n3178 VSS.n3165 4.5005
R64721 VSS.n6480 VSS.n3178 4.5005
R64722 VSS.n6609 VSS.n3178 4.5005
R64723 VSS.n3180 VSS.n3165 4.5005
R64724 VSS.n6480 VSS.n3180 4.5005
R64725 VSS.n6609 VSS.n3180 4.5005
R64726 VSS.n3177 VSS.n3165 4.5005
R64727 VSS.n6480 VSS.n3177 4.5005
R64728 VSS.n6609 VSS.n3177 4.5005
R64729 VSS.n3181 VSS.n3165 4.5005
R64730 VSS.n6480 VSS.n3181 4.5005
R64731 VSS.n6609 VSS.n3181 4.5005
R64732 VSS.n3176 VSS.n3165 4.5005
R64733 VSS.n6480 VSS.n3176 4.5005
R64734 VSS.n6609 VSS.n3176 4.5005
R64735 VSS.n3182 VSS.n3165 4.5005
R64736 VSS.n6480 VSS.n3182 4.5005
R64737 VSS.n6609 VSS.n3182 4.5005
R64738 VSS.n3175 VSS.n3165 4.5005
R64739 VSS.n6480 VSS.n3175 4.5005
R64740 VSS.n6609 VSS.n3175 4.5005
R64741 VSS.n3183 VSS.n3165 4.5005
R64742 VSS.n6480 VSS.n3183 4.5005
R64743 VSS.n6609 VSS.n3183 4.5005
R64744 VSS.n3174 VSS.n3165 4.5005
R64745 VSS.n6480 VSS.n3174 4.5005
R64746 VSS.n6609 VSS.n3174 4.5005
R64747 VSS.n3184 VSS.n3165 4.5005
R64748 VSS.n6480 VSS.n3184 4.5005
R64749 VSS.n6609 VSS.n3184 4.5005
R64750 VSS.n3173 VSS.n3165 4.5005
R64751 VSS.n6480 VSS.n3173 4.5005
R64752 VSS.n6609 VSS.n3173 4.5005
R64753 VSS.n3185 VSS.n3165 4.5005
R64754 VSS.n6480 VSS.n3185 4.5005
R64755 VSS.n6609 VSS.n3185 4.5005
R64756 VSS.n3172 VSS.n3165 4.5005
R64757 VSS.n6480 VSS.n3172 4.5005
R64758 VSS.n6609 VSS.n3172 4.5005
R64759 VSS.n3186 VSS.n3165 4.5005
R64760 VSS.n6480 VSS.n3186 4.5005
R64761 VSS.n6609 VSS.n3186 4.5005
R64762 VSS.n3171 VSS.n3165 4.5005
R64763 VSS.n6480 VSS.n3171 4.5005
R64764 VSS.n6609 VSS.n3171 4.5005
R64765 VSS.n3187 VSS.n3165 4.5005
R64766 VSS.n6480 VSS.n3187 4.5005
R64767 VSS.n6609 VSS.n3187 4.5005
R64768 VSS.n3170 VSS.n3165 4.5005
R64769 VSS.n6480 VSS.n3170 4.5005
R64770 VSS.n6609 VSS.n3170 4.5005
R64771 VSS.n3188 VSS.n3165 4.5005
R64772 VSS.n6480 VSS.n3188 4.5005
R64773 VSS.n6609 VSS.n3188 4.5005
R64774 VSS.n3169 VSS.n3165 4.5005
R64775 VSS.n6480 VSS.n3169 4.5005
R64776 VSS.n6609 VSS.n3169 4.5005
R64777 VSS.n3189 VSS.n3165 4.5005
R64778 VSS.n6480 VSS.n3189 4.5005
R64779 VSS.n6609 VSS.n3189 4.5005
R64780 VSS.n3168 VSS.n3165 4.5005
R64781 VSS.n6480 VSS.n3168 4.5005
R64782 VSS.n6609 VSS.n3168 4.5005
R64783 VSS.n3165 VSS.n3163 4.5005
R64784 VSS.n6480 VSS.n3163 4.5005
R64785 VSS.n6609 VSS.n3163 4.5005
R64786 VSS.n6610 VSS.n3165 4.5005
R64787 VSS.n6610 VSS.n6609 4.5005
R64788 VSS.n6608 VSS.n3165 4.5005
R64789 VSS.n6609 VSS.n6608 4.5005
R64790 VSS.n6840 VSS.n2931 4.5005
R64791 VSS.n2931 VSS.n2924 4.5005
R64792 VSS.n2931 VSS.n2919 4.5005
R64793 VSS.n6840 VSS.n2929 4.5005
R64794 VSS.n2929 VSS.n2924 4.5005
R64795 VSS.n2929 VSS.n2919 4.5005
R64796 VSS.n6840 VSS.n2932 4.5005
R64797 VSS.n2932 VSS.n2924 4.5005
R64798 VSS.n2932 VSS.n2919 4.5005
R64799 VSS.n6840 VSS.n2928 4.5005
R64800 VSS.n2928 VSS.n2924 4.5005
R64801 VSS.n2928 VSS.n2919 4.5005
R64802 VSS.n6840 VSS.n2933 4.5005
R64803 VSS.n2933 VSS.n2924 4.5005
R64804 VSS.n2933 VSS.n2919 4.5005
R64805 VSS.n6840 VSS.n2927 4.5005
R64806 VSS.n2927 VSS.n2924 4.5005
R64807 VSS.n2927 VSS.n2919 4.5005
R64808 VSS.n6840 VSS.n2934 4.5005
R64809 VSS.n2934 VSS.n2924 4.5005
R64810 VSS.n2934 VSS.n2919 4.5005
R64811 VSS.n6840 VSS.n2926 4.5005
R64812 VSS.n2926 VSS.n2924 4.5005
R64813 VSS.n2926 VSS.n2919 4.5005
R64814 VSS.n6840 VSS.n2935 4.5005
R64815 VSS.n2935 VSS.n2924 4.5005
R64816 VSS.n2935 VSS.n2919 4.5005
R64817 VSS.n6840 VSS.n2925 4.5005
R64818 VSS.n2925 VSS.n2924 4.5005
R64819 VSS.n2925 VSS.n2919 4.5005
R64820 VSS.n6840 VSS.n6839 4.5005
R64821 VSS.n6839 VSS.n2924 4.5005
R64822 VSS.n6839 VSS.n2919 4.5005
R64823 VSS.n8535 VSS.n1627 4.5005
R64824 VSS.n8538 VSS.n1627 4.5005
R64825 VSS.n8538 VSS.n1624 4.5005
R64826 VSS.n8538 VSS.n1629 4.5005
R64827 VSS.n8538 VSS.n1623 4.5005
R64828 VSS.n1630 VSS.n1617 4.5005
R64829 VSS.n8538 VSS.n1630 4.5005
R64830 VSS.n8535 VSS.n1622 4.5005
R64831 VSS.n1622 VSS.n1617 4.5005
R64832 VSS.n8538 VSS.n1622 4.5005
R64833 VSS.n8538 VSS.n1632 4.5005
R64834 VSS.n8535 VSS.n1632 4.5005
R64835 VSS.n8538 VSS.n1621 4.5005
R64836 VSS.n8538 VSS.n8537 4.5005
R64837 VSS.n8538 VSS.n1620 4.5005
R64838 VSS.n8539 VSS.n1617 4.5005
R64839 VSS.n8539 VSS.n8538 4.5005
R64840 VSS.n8686 VSS.n1485 4.5005
R64841 VSS.n8684 VSS.n1485 4.5005
R64842 VSS.n8686 VSS.n1486 4.5005
R64843 VSS.n8684 VSS.n1486 4.5005
R64844 VSS.n8684 VSS.n1484 4.5005
R64845 VSS.n1495 VSS.n1484 4.5005
R64846 VSS.n8686 VSS.n1484 4.5005
R64847 VSS.n8684 VSS.n1487 4.5005
R64848 VSS.n8686 VSS.n1487 4.5005
R64849 VSS.n8684 VSS.n1506 4.5005
R64850 VSS.n8684 VSS.n8669 4.5005
R64851 VSS.n8684 VSS.n1504 4.5005
R64852 VSS.n8684 VSS.n8671 4.5005
R64853 VSS.n8684 VSS.n1503 4.5005
R64854 VSS.n8684 VSS.n8673 4.5005
R64855 VSS.n8684 VSS.n1502 4.5005
R64856 VSS.n8684 VSS.n8675 4.5005
R64857 VSS.n8686 VSS.n1479 4.5005
R64858 VSS.n8684 VSS.n1479 4.5005
R64859 VSS.n8686 VSS.n1488 4.5005
R64860 VSS.n1495 VSS.n1488 4.5005
R64861 VSS.n8684 VSS.n1488 4.5005
R64862 VSS.n8686 VSS.n1478 4.5005
R64863 VSS.n8684 VSS.n1478 4.5005
R64864 VSS.n8684 VSS.n8677 4.5005
R64865 VSS.n8684 VSS.n1501 4.5005
R64866 VSS.n8684 VSS.n8679 4.5005
R64867 VSS.n8684 VSS.n1500 4.5005
R64868 VSS.n8684 VSS.n8681 4.5005
R64869 VSS.n8684 VSS.n1499 4.5005
R64870 VSS.n8684 VSS.n8683 4.5005
R64871 VSS.n1498 VSS.n1495 4.5005
R64872 VSS.n8684 VSS.n1498 4.5005
R64873 VSS.n8685 VSS.n8684 4.5005
R64874 VSS.n8685 VSS.n1495 4.5005
R64875 VSS.n8686 VSS.n8685 4.5005
R64876 VSS.n974 VSS.n956 4.5005
R64877 VSS.n9150 VSS.n974 4.5005
R64878 VSS.n9121 VSS.n956 4.5005
R64879 VSS.n9120 VSS.n956 4.5005
R64880 VSS.n9124 VSS.n956 4.5005
R64881 VSS.n9123 VSS.n956 4.5005
R64882 VSS.n9127 VSS.n956 4.5005
R64883 VSS.n9126 VSS.n956 4.5005
R64884 VSS.n9130 VSS.n956 4.5005
R64885 VSS.n9129 VSS.n956 4.5005
R64886 VSS.n9133 VSS.n956 4.5005
R64887 VSS.n9132 VSS.n956 4.5005
R64888 VSS.n9136 VSS.n956 4.5005
R64889 VSS.n9135 VSS.n956 4.5005
R64890 VSS.n9139 VSS.n956 4.5005
R64891 VSS.n9138 VSS.n956 4.5005
R64892 VSS.n9142 VSS.n956 4.5005
R64893 VSS.n9141 VSS.n956 4.5005
R64894 VSS.n9145 VSS.n956 4.5005
R64895 VSS.n9144 VSS.n956 4.5005
R64896 VSS.n9148 VSS.n956 4.5005
R64897 VSS.n9147 VSS.n956 4.5005
R64898 VSS.n9151 VSS.n956 4.5005
R64899 VSS.n9153 VSS.n956 4.5005
R64900 VSS.n9150 VSS.n973 4.5005
R64901 VSS.n973 VSS.n956 4.5005
R64902 VSS.n9223 VSS.n902 4.5005
R64903 VSS.n9221 VSS.n902 4.5005
R64904 VSS.n9221 VSS.n9198 4.5005
R64905 VSS.n9221 VSS.n927 4.5005
R64906 VSS.n9221 VSS.n9199 4.5005
R64907 VSS.n9221 VSS.n926 4.5005
R64908 VSS.n9221 VSS.n9200 4.5005
R64909 VSS.n9221 VSS.n925 4.5005
R64910 VSS.n9221 VSS.n9201 4.5005
R64911 VSS.n9221 VSS.n924 4.5005
R64912 VSS.n9221 VSS.n9202 4.5005
R64913 VSS.n9221 VSS.n923 4.5005
R64914 VSS.n9221 VSS.n9203 4.5005
R64915 VSS.n9221 VSS.n922 4.5005
R64916 VSS.n9221 VSS.n9204 4.5005
R64917 VSS.n9221 VSS.n921 4.5005
R64918 VSS.n9221 VSS.n9205 4.5005
R64919 VSS.n9221 VSS.n920 4.5005
R64920 VSS.n9221 VSS.n9206 4.5005
R64921 VSS.n9221 VSS.n919 4.5005
R64922 VSS.n9221 VSS.n9207 4.5005
R64923 VSS.n9221 VSS.n918 4.5005
R64924 VSS.n9221 VSS.n9220 4.5005
R64925 VSS.n9221 VSS.n917 4.5005
R64926 VSS.n9223 VSS.n9222 4.5005
R64927 VSS.n9222 VSS.n9221 4.5005
R64928 VSS.n2574 VSS.n2573 4.5005
R64929 VSS.n2573 VSS.n2572 4.5005
R64930 VSS.n2735 VSS.n2659 4.5005
R64931 VSS.n2734 VSS.n2733 4.5005
R64932 VSS.n2661 VSS.n2660 4.5005
R64933 VSS.n2729 VSS.n2663 4.5005
R64934 VSS.n2728 VSS.n2664 4.5005
R64935 VSS.n2727 VSS.n2665 4.5005
R64936 VSS.n2668 VSS.n2666 4.5005
R64937 VSS.n2723 VSS.n2669 4.5005
R64938 VSS.n2722 VSS.n2670 4.5005
R64939 VSS.n2721 VSS.n2671 4.5005
R64940 VSS.n2674 VSS.n2672 4.5005
R64941 VSS.n2717 VSS.n2675 4.5005
R64942 VSS.n2716 VSS.n2676 4.5005
R64943 VSS.n2715 VSS.n2677 4.5005
R64944 VSS.n2680 VSS.n2678 4.5005
R64945 VSS.n2711 VSS.n2681 4.5005
R64946 VSS.n2710 VSS.n2682 4.5005
R64947 VSS.n2709 VSS.n2683 4.5005
R64948 VSS.n2686 VSS.n2684 4.5005
R64949 VSS.n2705 VSS.n2687 4.5005
R64950 VSS.n2704 VSS.n2688 4.5005
R64951 VSS.n2703 VSS.n2689 4.5005
R64952 VSS.n2692 VSS.n2690 4.5005
R64953 VSS.n2699 VSS.n2693 4.5005
R64954 VSS.n2698 VSS.n2694 4.5005
R64955 VSS.n2697 VSS.n2695 4.5005
R64956 VSS.n2697 VSS.n2696 4.5005
R64957 VSS.n2698 VSS.n2691 4.5005
R64958 VSS.n2700 VSS.n2699 4.5005
R64959 VSS.n2701 VSS.n2690 4.5005
R64960 VSS.n2703 VSS.n2702 4.5005
R64961 VSS.n2704 VSS.n2685 4.5005
R64962 VSS.n2706 VSS.n2705 4.5005
R64963 VSS.n2707 VSS.n2684 4.5005
R64964 VSS.n2709 VSS.n2708 4.5005
R64965 VSS.n2710 VSS.n2679 4.5005
R64966 VSS.n2712 VSS.n2711 4.5005
R64967 VSS.n2713 VSS.n2678 4.5005
R64968 VSS.n2715 VSS.n2714 4.5005
R64969 VSS.n2716 VSS.n2673 4.5005
R64970 VSS.n2718 VSS.n2717 4.5005
R64971 VSS.n2719 VSS.n2672 4.5005
R64972 VSS.n2721 VSS.n2720 4.5005
R64973 VSS.n2722 VSS.n2667 4.5005
R64974 VSS.n2724 VSS.n2723 4.5005
R64975 VSS.n2725 VSS.n2666 4.5005
R64976 VSS.n2727 VSS.n2726 4.5005
R64977 VSS.n2728 VSS.n2662 4.5005
R64978 VSS.n2730 VSS.n2729 4.5005
R64979 VSS.n2731 VSS.n2661 4.5005
R64980 VSS.n2733 VSS.n2732 4.5005
R64981 VSS.n2659 VSS.n2658 4.5005
R64982 VSS.n2738 VSS.n2737 4.5005
R64983 VSS.n2737 VSS.n2736 4.5005
R64984 VSS.n7138 VSS.n7132 4.5005
R64985 VSS.n7138 VSS.n7137 4.5005
R64986 VSS.n7139 VSS.n7138 4.5005
R64987 VSS.n7137 VSS.n2576 4.5005
R64988 VSS.n7139 VSS.n2576 4.5005
R64989 VSS.n7143 VSS.n7140 4.5005
R64990 VSS.n7268 VSS.n2472 4.5005
R64991 VSS.n7137 VSS.n7136 4.5005
R64992 VSS.n7136 VSS.n7132 4.5005
R64993 VSS.n2788 VSS.n2778 4.5005
R64994 VSS.n2786 VSS.n2778 4.5005
R64995 VSS.n2782 VSS.n2778 4.5005
R64996 VSS.n7129 VSS.n2583 4.5005
R64997 VSS.n7129 VSS.n7128 4.5005
R64998 VSS.n7130 VSS.n7129 4.5005
R64999 VSS.n2786 VSS.n2783 4.5005
R65000 VSS.n2783 VSS.n2782 4.5005
R65001 VSS.n7128 VSS.n2580 4.5005
R65002 VSS.n7130 VSS.n2580 4.5005
R65003 VSS.n7128 VSS.n7127 4.5005
R65004 VSS.n7127 VSS.n2583 4.5005
R65005 VSS.n2787 VSS.n2786 4.5005
R65006 VSS.n2788 VSS.n2787 4.5005
R65007 VSS.n2775 VSS.n2773 4.5005
R65008 VSS.n2790 VSS.n2773 4.5005
R65009 VSS.n2791 VSS.n2790 4.5005
R65010 VSS.n4764 VSS.n4722 4.5005
R65011 VSS.n4722 VSS.n4584 4.5005
R65012 VSS.n4762 VSS.n4722 4.5005
R65013 VSS.n4735 VSS.n4584 4.5005
R65014 VSS.n4762 VSS.n4735 4.5005
R65015 VSS.n4739 VSS.n4584 4.5005
R65016 VSS.n4762 VSS.n4739 4.5005
R65017 VSS.n4733 VSS.n4584 4.5005
R65018 VSS.n4762 VSS.n4733 4.5005
R65019 VSS.n4741 VSS.n4584 4.5005
R65020 VSS.n4762 VSS.n4741 4.5005
R65021 VSS.n4732 VSS.n4584 4.5005
R65022 VSS.n4762 VSS.n4732 4.5005
R65023 VSS.n4761 VSS.n4584 4.5005
R65024 VSS.n4761 VSS.n4729 4.5005
R65025 VSS.n4762 VSS.n4761 4.5005
R65026 VSS.n4729 VSS.n4586 4.5005
R65027 VSS.n4762 VSS.n4586 4.5005
R65028 VSS.n4586 VSS.n4584 4.5005
R65029 VSS.n4764 VSS.n4586 4.5005
R65030 VSS.n4764 VSS.n4726 4.5005
R65031 VSS.n4726 VSS.n4584 4.5005
R65032 VSS.n4729 VSS.n4726 4.5005
R65033 VSS.n4762 VSS.n4726 4.5005
R65034 VSS.n4764 VSS.n4585 4.5005
R65035 VSS.n4585 VSS.n4584 4.5005
R65036 VSS.n4729 VSS.n4585 4.5005
R65037 VSS.n4762 VSS.n4585 4.5005
R65038 VSS.n4764 VSS.n4763 4.5005
R65039 VSS.n4763 VSS.n4584 4.5005
R65040 VSS.n4763 VSS.n4729 4.5005
R65041 VSS.n4763 VSS.n4762 4.5005
R65042 VSS.n6239 VSS.n3866 4.5005
R65043 VSS.n6248 VSS.n6239 4.5005
R65044 VSS.n6239 VSS.n3868 4.5005
R65045 VSS.n6239 VSS.n3867 4.5005
R65046 VSS.n3866 VSS.n3865 4.5005
R65047 VSS.n6248 VSS.n3865 4.5005
R65048 VSS.n3868 VSS.n3865 4.5005
R65049 VSS.n3867 VSS.n3865 4.5005
R65050 VSS.n6249 VSS.n3867 4.5005
R65051 VSS.n6249 VSS.n3868 4.5005
R65052 VSS.n6249 VSS.n3866 4.5005
R65053 VSS.n6249 VSS.n6248 4.5005
R65054 VSS.n3867 VSS.n3860 4.5005
R65055 VSS.n3868 VSS.n3860 4.5005
R65056 VSS.n3866 VSS.n3860 4.5005
R65057 VSS.n6248 VSS.n3860 4.5005
R65058 VSS.n3867 VSS.n3862 4.5005
R65059 VSS.n3868 VSS.n3862 4.5005
R65060 VSS.n6248 VSS.n3862 4.5005
R65061 VSS.n3873 VSS.n3868 4.5005
R65062 VSS.n6248 VSS.n3873 4.5005
R65063 VSS.n6242 VSS.n3868 4.5005
R65064 VSS.n6248 VSS.n6242 4.5005
R65065 VSS.n3871 VSS.n3868 4.5005
R65066 VSS.n6248 VSS.n3871 4.5005
R65067 VSS.n6245 VSS.n3868 4.5005
R65068 VSS.n6248 VSS.n6245 4.5005
R65069 VSS.n3870 VSS.n3868 4.5005
R65070 VSS.n6248 VSS.n3870 4.5005
R65071 VSS.n6247 VSS.n3868 4.5005
R65072 VSS.n6247 VSS.n3866 4.5005
R65073 VSS.n6248 VSS.n6247 4.5005
R65074 VSS.n3844 VSS.n3834 4.5005
R65075 VSS.n3844 VSS.n3835 4.5005
R65076 VSS.n6263 VSS.n3844 4.5005
R65077 VSS.n3841 VSS.n3835 4.5005
R65078 VSS.n6263 VSS.n3841 4.5005
R65079 VSS.n3847 VSS.n3835 4.5005
R65080 VSS.n6263 VSS.n3847 4.5005
R65081 VSS.n3840 VSS.n3835 4.5005
R65082 VSS.n6263 VSS.n3840 4.5005
R65083 VSS.n3850 VSS.n3835 4.5005
R65084 VSS.n6263 VSS.n3850 4.5005
R65085 VSS.n3839 VSS.n3834 4.5005
R65086 VSS.n3839 VSS.n3835 4.5005
R65087 VSS.n6263 VSS.n3839 4.5005
R65088 VSS.n3851 VSS.n3833 4.5005
R65089 VSS.n6263 VSS.n3851 4.5005
R65090 VSS.n3851 VSS.n3835 4.5005
R65091 VSS.n3851 VSS.n3834 4.5005
R65092 VSS.n3838 VSS.n3833 4.5005
R65093 VSS.n6263 VSS.n3838 4.5005
R65094 VSS.n3838 VSS.n3835 4.5005
R65095 VSS.n3838 VSS.n3834 4.5005
R65096 VSS.n6262 VSS.n3833 4.5005
R65097 VSS.n6263 VSS.n6262 4.5005
R65098 VSS.n6262 VSS.n3835 4.5005
R65099 VSS.n6262 VSS.n3834 4.5005
R65100 VSS.n3837 VSS.n3834 4.5005
R65101 VSS.n3837 VSS.n3835 4.5005
R65102 VSS.n3837 VSS.n3833 4.5005
R65103 VSS.n6263 VSS.n3837 4.5005
R65104 VSS.n6264 VSS.n3834 4.5005
R65105 VSS.n6264 VSS.n3835 4.5005
R65106 VSS.n6264 VSS.n3833 4.5005
R65107 VSS.n6264 VSS.n6263 4.5005
R65108 VSS.n3246 VSS.n3232 4.5005
R65109 VSS.n3246 VSS.n3233 4.5005
R65110 VSS.n6572 VSS.n3246 4.5005
R65111 VSS.n3249 VSS.n3233 4.5005
R65112 VSS.n6572 VSS.n3249 4.5005
R65113 VSS.n3245 VSS.n3233 4.5005
R65114 VSS.n6572 VSS.n3245 4.5005
R65115 VSS.n3251 VSS.n3233 4.5005
R65116 VSS.n6572 VSS.n3251 4.5005
R65117 VSS.n3244 VSS.n3233 4.5005
R65118 VSS.n6572 VSS.n3244 4.5005
R65119 VSS.n3253 VSS.n3233 4.5005
R65120 VSS.n6572 VSS.n3253 4.5005
R65121 VSS.n3243 VSS.n3233 4.5005
R65122 VSS.n6572 VSS.n3243 4.5005
R65123 VSS.n3255 VSS.n3233 4.5005
R65124 VSS.n6572 VSS.n3255 4.5005
R65125 VSS.n3242 VSS.n3233 4.5005
R65126 VSS.n6572 VSS.n3242 4.5005
R65127 VSS.n3257 VSS.n3233 4.5005
R65128 VSS.n6572 VSS.n3257 4.5005
R65129 VSS.n3241 VSS.n3233 4.5005
R65130 VSS.n6572 VSS.n3241 4.5005
R65131 VSS.n3259 VSS.n3233 4.5005
R65132 VSS.n6572 VSS.n3259 4.5005
R65133 VSS.n3240 VSS.n3233 4.5005
R65134 VSS.n6572 VSS.n3240 4.5005
R65135 VSS.n3261 VSS.n3233 4.5005
R65136 VSS.n6572 VSS.n3261 4.5005
R65137 VSS.n3239 VSS.n3233 4.5005
R65138 VSS.n6572 VSS.n3239 4.5005
R65139 VSS.n3263 VSS.n3233 4.5005
R65140 VSS.n6572 VSS.n3263 4.5005
R65141 VSS.n3238 VSS.n3233 4.5005
R65142 VSS.n6572 VSS.n3238 4.5005
R65143 VSS.n3265 VSS.n3233 4.5005
R65144 VSS.n6572 VSS.n3265 4.5005
R65145 VSS.n3237 VSS.n3233 4.5005
R65146 VSS.n6572 VSS.n3237 4.5005
R65147 VSS.n3267 VSS.n3233 4.5005
R65148 VSS.n6572 VSS.n3267 4.5005
R65149 VSS.n3236 VSS.n3233 4.5005
R65150 VSS.n6572 VSS.n3236 4.5005
R65151 VSS.n6571 VSS.n3233 4.5005
R65152 VSS.n6572 VSS.n6571 4.5005
R65153 VSS.n3235 VSS.n3233 4.5005
R65154 VSS.n6572 VSS.n3235 4.5005
R65155 VSS.n6573 VSS.n3232 4.5005
R65156 VSS.n6573 VSS.n3233 4.5005
R65157 VSS.n6573 VSS.n6572 4.5005
R65158 VSS.n6960 VSS.n2807 4.5005
R65159 VSS.n2807 VSS.n2798 4.5005
R65160 VSS.n6964 VSS.n2807 4.5005
R65161 VSS.n2804 VSS.n2798 4.5005
R65162 VSS.n6964 VSS.n2804 4.5005
R65163 VSS.n2809 VSS.n2798 4.5005
R65164 VSS.n6964 VSS.n2809 4.5005
R65165 VSS.n2803 VSS.n2798 4.5005
R65166 VSS.n6964 VSS.n2803 4.5005
R65167 VSS.n2811 VSS.n2798 4.5005
R65168 VSS.n6964 VSS.n2811 4.5005
R65169 VSS.n2802 VSS.n2798 4.5005
R65170 VSS.n6964 VSS.n2802 4.5005
R65171 VSS.n2813 VSS.n2798 4.5005
R65172 VSS.n6964 VSS.n2813 4.5005
R65173 VSS.n2801 VSS.n2798 4.5005
R65174 VSS.n6964 VSS.n2801 4.5005
R65175 VSS.n6963 VSS.n2798 4.5005
R65176 VSS.n6964 VSS.n6963 4.5005
R65177 VSS.n2800 VSS.n2798 4.5005
R65178 VSS.n6964 VSS.n2800 4.5005
R65179 VSS.n6965 VSS.n2798 4.5005
R65180 VSS.n6965 VSS.n2797 4.5005
R65181 VSS.n6965 VSS.n6964 4.5005
R65182 VSS.n8301 VSS.n1707 4.5005
R65183 VSS.n1707 VSS.n1706 4.5005
R65184 VSS.n8298 VSS.n1707 4.5005
R65185 VSS.n8285 VSS.n1706 4.5005
R65186 VSS.n8298 VSS.n8285 4.5005
R65187 VSS.n8288 VSS.n1706 4.5005
R65188 VSS.n8298 VSS.n8288 4.5005
R65189 VSS.n8284 VSS.n1706 4.5005
R65190 VSS.n8298 VSS.n8284 4.5005
R65191 VSS.n8289 VSS.n1706 4.5005
R65192 VSS.n8298 VSS.n8289 4.5005
R65193 VSS.n8283 VSS.n1706 4.5005
R65194 VSS.n8298 VSS.n8283 4.5005
R65195 VSS.n8296 VSS.n1706 4.5005
R65196 VSS.n8298 VSS.n8296 4.5005
R65197 VSS.n8282 VSS.n1706 4.5005
R65198 VSS.n8298 VSS.n8282 4.5005
R65199 VSS.n8297 VSS.n1706 4.5005
R65200 VSS.n8298 VSS.n8297 4.5005
R65201 VSS.n8299 VSS.n1706 4.5005
R65202 VSS.n8299 VSS.n8298 4.5005
R65203 VSS.n8279 VSS.n1706 4.5005
R65204 VSS.n8294 VSS.n8279 4.5005
R65205 VSS.n8298 VSS.n8279 4.5005
R65206 VSS.n8278 VSS.n1713 4.5005
R65207 VSS.n8278 VSS.n1714 4.5005
R65208 VSS.n8278 VSS.n8277 4.5005
R65209 VSS.n1729 VSS.n1714 4.5005
R65210 VSS.n8277 VSS.n1729 4.5005
R65211 VSS.n1726 VSS.n1714 4.5005
R65212 VSS.n8277 VSS.n1726 4.5005
R65213 VSS.n1731 VSS.n1714 4.5005
R65214 VSS.n8277 VSS.n1731 4.5005
R65215 VSS.n1725 VSS.n1714 4.5005
R65216 VSS.n8277 VSS.n1725 4.5005
R65217 VSS.n1733 VSS.n1714 4.5005
R65218 VSS.n8277 VSS.n1733 4.5005
R65219 VSS.n1724 VSS.n1714 4.5005
R65220 VSS.n8277 VSS.n1724 4.5005
R65221 VSS.n1735 VSS.n1714 4.5005
R65222 VSS.n8277 VSS.n1735 4.5005
R65223 VSS.n1723 VSS.n1714 4.5005
R65224 VSS.n8277 VSS.n1723 4.5005
R65225 VSS.n1737 VSS.n1714 4.5005
R65226 VSS.n8277 VSS.n1737 4.5005
R65227 VSS.n1722 VSS.n1714 4.5005
R65228 VSS.n8277 VSS.n1722 4.5005
R65229 VSS.n1739 VSS.n1714 4.5005
R65230 VSS.n8277 VSS.n1739 4.5005
R65231 VSS.n1721 VSS.n1714 4.5005
R65232 VSS.n8277 VSS.n1721 4.5005
R65233 VSS.n1741 VSS.n1714 4.5005
R65234 VSS.n8277 VSS.n1741 4.5005
R65235 VSS.n1720 VSS.n1714 4.5005
R65236 VSS.n8277 VSS.n1720 4.5005
R65237 VSS.n1743 VSS.n1714 4.5005
R65238 VSS.n8277 VSS.n1743 4.5005
R65239 VSS.n1719 VSS.n1714 4.5005
R65240 VSS.n8277 VSS.n1719 4.5005
R65241 VSS.n1745 VSS.n1714 4.5005
R65242 VSS.n8277 VSS.n1745 4.5005
R65243 VSS.n1718 VSS.n1714 4.5005
R65244 VSS.n8277 VSS.n1718 4.5005
R65245 VSS.n1747 VSS.n1714 4.5005
R65246 VSS.n8277 VSS.n1747 4.5005
R65247 VSS.n1717 VSS.n1714 4.5005
R65248 VSS.n8277 VSS.n1717 4.5005
R65249 VSS.n1749 VSS.n1714 4.5005
R65250 VSS.n8277 VSS.n1749 4.5005
R65251 VSS.n1716 VSS.n1714 4.5005
R65252 VSS.n8277 VSS.n1716 4.5005
R65253 VSS.n8276 VSS.n1713 4.5005
R65254 VSS.n8276 VSS.n1714 4.5005
R65255 VSS.n8277 VSS.n8276 4.5005
R65256 VSS.n8275 VSS.n1752 4.5005
R65257 VSS.n8275 VSS.n1753 4.5005
R65258 VSS.n8275 VSS.n8274 4.5005
R65259 VSS.n1768 VSS.n1753 4.5005
R65260 VSS.n8274 VSS.n1768 4.5005
R65261 VSS.n1765 VSS.n1753 4.5005
R65262 VSS.n8274 VSS.n1765 4.5005
R65263 VSS.n1770 VSS.n1753 4.5005
R65264 VSS.n8274 VSS.n1770 4.5005
R65265 VSS.n1764 VSS.n1753 4.5005
R65266 VSS.n8274 VSS.n1764 4.5005
R65267 VSS.n1772 VSS.n1753 4.5005
R65268 VSS.n8274 VSS.n1772 4.5005
R65269 VSS.n1763 VSS.n1753 4.5005
R65270 VSS.n8274 VSS.n1763 4.5005
R65271 VSS.n1774 VSS.n1753 4.5005
R65272 VSS.n8274 VSS.n1774 4.5005
R65273 VSS.n1762 VSS.n1753 4.5005
R65274 VSS.n8274 VSS.n1762 4.5005
R65275 VSS.n1776 VSS.n1753 4.5005
R65276 VSS.n8274 VSS.n1776 4.5005
R65277 VSS.n1761 VSS.n1753 4.5005
R65278 VSS.n8274 VSS.n1761 4.5005
R65279 VSS.n1778 VSS.n1753 4.5005
R65280 VSS.n8274 VSS.n1778 4.5005
R65281 VSS.n1760 VSS.n1753 4.5005
R65282 VSS.n8274 VSS.n1760 4.5005
R65283 VSS.n1780 VSS.n1753 4.5005
R65284 VSS.n8274 VSS.n1780 4.5005
R65285 VSS.n1759 VSS.n1753 4.5005
R65286 VSS.n8274 VSS.n1759 4.5005
R65287 VSS.n1782 VSS.n1753 4.5005
R65288 VSS.n8274 VSS.n1782 4.5005
R65289 VSS.n1758 VSS.n1753 4.5005
R65290 VSS.n8274 VSS.n1758 4.5005
R65291 VSS.n1784 VSS.n1753 4.5005
R65292 VSS.n8274 VSS.n1784 4.5005
R65293 VSS.n1757 VSS.n1753 4.5005
R65294 VSS.n8274 VSS.n1757 4.5005
R65295 VSS.n1786 VSS.n1753 4.5005
R65296 VSS.n8274 VSS.n1786 4.5005
R65297 VSS.n1756 VSS.n1753 4.5005
R65298 VSS.n8274 VSS.n1756 4.5005
R65299 VSS.n1788 VSS.n1753 4.5005
R65300 VSS.n8274 VSS.n1788 4.5005
R65301 VSS.n1755 VSS.n1753 4.5005
R65302 VSS.n8274 VSS.n1755 4.5005
R65303 VSS.n8273 VSS.n1752 4.5005
R65304 VSS.n8273 VSS.n1753 4.5005
R65305 VSS.n8274 VSS.n8273 4.5005
R65306 VSS.n8272 VSS.n1791 4.5005
R65307 VSS.n8272 VSS.n1792 4.5005
R65308 VSS.n8272 VSS.n8271 4.5005
R65309 VSS.n1807 VSS.n1792 4.5005
R65310 VSS.n8271 VSS.n1807 4.5005
R65311 VSS.n1804 VSS.n1792 4.5005
R65312 VSS.n8271 VSS.n1804 4.5005
R65313 VSS.n1809 VSS.n1792 4.5005
R65314 VSS.n8271 VSS.n1809 4.5005
R65315 VSS.n1803 VSS.n1792 4.5005
R65316 VSS.n8271 VSS.n1803 4.5005
R65317 VSS.n1811 VSS.n1792 4.5005
R65318 VSS.n8271 VSS.n1811 4.5005
R65319 VSS.n1802 VSS.n1792 4.5005
R65320 VSS.n8271 VSS.n1802 4.5005
R65321 VSS.n1813 VSS.n1792 4.5005
R65322 VSS.n8271 VSS.n1813 4.5005
R65323 VSS.n1801 VSS.n1792 4.5005
R65324 VSS.n8271 VSS.n1801 4.5005
R65325 VSS.n1815 VSS.n1792 4.5005
R65326 VSS.n8271 VSS.n1815 4.5005
R65327 VSS.n1800 VSS.n1792 4.5005
R65328 VSS.n8271 VSS.n1800 4.5005
R65329 VSS.n1817 VSS.n1792 4.5005
R65330 VSS.n8271 VSS.n1817 4.5005
R65331 VSS.n1799 VSS.n1792 4.5005
R65332 VSS.n8271 VSS.n1799 4.5005
R65333 VSS.n1819 VSS.n1792 4.5005
R65334 VSS.n8271 VSS.n1819 4.5005
R65335 VSS.n1798 VSS.n1792 4.5005
R65336 VSS.n8271 VSS.n1798 4.5005
R65337 VSS.n1821 VSS.n1792 4.5005
R65338 VSS.n8271 VSS.n1821 4.5005
R65339 VSS.n1797 VSS.n1792 4.5005
R65340 VSS.n8271 VSS.n1797 4.5005
R65341 VSS.n1823 VSS.n1792 4.5005
R65342 VSS.n8271 VSS.n1823 4.5005
R65343 VSS.n1796 VSS.n1792 4.5005
R65344 VSS.n8271 VSS.n1796 4.5005
R65345 VSS.n1825 VSS.n1792 4.5005
R65346 VSS.n8271 VSS.n1825 4.5005
R65347 VSS.n1795 VSS.n1792 4.5005
R65348 VSS.n8271 VSS.n1795 4.5005
R65349 VSS.n1827 VSS.n1792 4.5005
R65350 VSS.n8271 VSS.n1827 4.5005
R65351 VSS.n1794 VSS.n1792 4.5005
R65352 VSS.n8271 VSS.n1794 4.5005
R65353 VSS.n8270 VSS.n1791 4.5005
R65354 VSS.n8270 VSS.n1792 4.5005
R65355 VSS.n8271 VSS.n8270 4.5005
R65356 VSS.n4594 VSS.n4588 4.5005
R65357 VSS.n4594 VSS.n4589 4.5005
R65358 VSS.n4718 VSS.n4594 4.5005
R65359 VSS.n4720 VSS.n4594 4.5005
R65360 VSS.n4596 VSS.n4588 4.5005
R65361 VSS.n4596 VSS.n4589 4.5005
R65362 VSS.n4720 VSS.n4596 4.5005
R65363 VSS.n4593 VSS.n4589 4.5005
R65364 VSS.n4720 VSS.n4593 4.5005
R65365 VSS.n4598 VSS.n4589 4.5005
R65366 VSS.n4720 VSS.n4598 4.5005
R65367 VSS.n4592 VSS.n4589 4.5005
R65368 VSS.n4720 VSS.n4592 4.5005
R65369 VSS.n4600 VSS.n4589 4.5005
R65370 VSS.n4720 VSS.n4600 4.5005
R65371 VSS.n4721 VSS.n4588 4.5005
R65372 VSS.n4721 VSS.n4589 4.5005
R65373 VSS.n4721 VSS.n4720 4.5005
R65374 VSS.n4720 VSS.n4602 4.5005
R65375 VSS.n4718 VSS.n4602 4.5005
R65376 VSS.n4602 VSS.n4588 4.5005
R65377 VSS.n4720 VSS.n4591 4.5005
R65378 VSS.n4718 VSS.n4591 4.5005
R65379 VSS.n4591 VSS.n4588 4.5005
R65380 VSS.n4720 VSS.n4719 4.5005
R65381 VSS.n4719 VSS.n4718 4.5005
R65382 VSS.n4719 VSS.n4589 4.5005
R65383 VSS.n4719 VSS.n4588 4.5005
R65384 VSS.n4631 VSS.n4622 4.5005
R65385 VSS.n4677 VSS.n4622 4.5005
R65386 VSS.n4703 VSS.n4622 4.5005
R65387 VSS.n4705 VSS.n4622 4.5005
R65388 VSS.n4631 VSS.n4624 4.5005
R65389 VSS.n4677 VSS.n4624 4.5005
R65390 VSS.n4705 VSS.n4624 4.5005
R65391 VSS.n4677 VSS.n4621 4.5005
R65392 VSS.n4705 VSS.n4621 4.5005
R65393 VSS.n4677 VSS.n4625 4.5005
R65394 VSS.n4705 VSS.n4625 4.5005
R65395 VSS.n4677 VSS.n4620 4.5005
R65396 VSS.n4705 VSS.n4620 4.5005
R65397 VSS.n4677 VSS.n4626 4.5005
R65398 VSS.n4705 VSS.n4626 4.5005
R65399 VSS.n4631 VSS.n4619 4.5005
R65400 VSS.n4677 VSS.n4619 4.5005
R65401 VSS.n4705 VSS.n4619 4.5005
R65402 VSS.n4705 VSS.n4627 4.5005
R65403 VSS.n4703 VSS.n4627 4.5005
R65404 VSS.n4631 VSS.n4627 4.5005
R65405 VSS.n4705 VSS.n4618 4.5005
R65406 VSS.n4703 VSS.n4618 4.5005
R65407 VSS.n4631 VSS.n4618 4.5005
R65408 VSS.n4704 VSS.n4631 4.5005
R65409 VSS.n4704 VSS.n4677 4.5005
R65410 VSS.n4705 VSS.n4704 4.5005
R65411 VSS.n4704 VSS.n4703 4.5005
R65412 VSS.n4345 VSS.n4339 4.5005
R65413 VSS.n4345 VSS.n4340 4.5005
R65414 VSS.n5231 VSS.n4345 4.5005
R65415 VSS.n5233 VSS.n4345 4.5005
R65416 VSS.n4347 VSS.n4339 4.5005
R65417 VSS.n4347 VSS.n4340 4.5005
R65418 VSS.n5233 VSS.n4347 4.5005
R65419 VSS.n4344 VSS.n4340 4.5005
R65420 VSS.n5233 VSS.n4344 4.5005
R65421 VSS.n4349 VSS.n4340 4.5005
R65422 VSS.n5233 VSS.n4349 4.5005
R65423 VSS.n4343 VSS.n4340 4.5005
R65424 VSS.n5233 VSS.n4343 4.5005
R65425 VSS.n4351 VSS.n4340 4.5005
R65426 VSS.n5233 VSS.n4351 4.5005
R65427 VSS.n5234 VSS.n4339 4.5005
R65428 VSS.n5234 VSS.n4340 4.5005
R65429 VSS.n5234 VSS.n5233 4.5005
R65430 VSS.n5233 VSS.n4353 4.5005
R65431 VSS.n5231 VSS.n4353 4.5005
R65432 VSS.n4353 VSS.n4339 4.5005
R65433 VSS.n5233 VSS.n4342 4.5005
R65434 VSS.n5231 VSS.n4342 4.5005
R65435 VSS.n4342 VSS.n4339 4.5005
R65436 VSS.n5232 VSS.n4339 4.5005
R65437 VSS.n5232 VSS.n4340 4.5005
R65438 VSS.n5233 VSS.n5232 4.5005
R65439 VSS.n5232 VSS.n5231 4.5005
R65440 VSS.n4394 VSS.n4385 4.5005
R65441 VSS.n4397 VSS.n4385 4.5005
R65442 VSS.n5204 VSS.n4385 4.5005
R65443 VSS.n5206 VSS.n4385 4.5005
R65444 VSS.n4394 VSS.n4387 4.5005
R65445 VSS.n4397 VSS.n4387 4.5005
R65446 VSS.n5206 VSS.n4387 4.5005
R65447 VSS.n4397 VSS.n4384 4.5005
R65448 VSS.n5206 VSS.n4384 4.5005
R65449 VSS.n4397 VSS.n4388 4.5005
R65450 VSS.n5206 VSS.n4388 4.5005
R65451 VSS.n4397 VSS.n4383 4.5005
R65452 VSS.n5206 VSS.n4383 4.5005
R65453 VSS.n4397 VSS.n4389 4.5005
R65454 VSS.n5206 VSS.n4389 4.5005
R65455 VSS.n4394 VSS.n4382 4.5005
R65456 VSS.n4397 VSS.n4382 4.5005
R65457 VSS.n5206 VSS.n4382 4.5005
R65458 VSS.n5206 VSS.n4390 4.5005
R65459 VSS.n5204 VSS.n4390 4.5005
R65460 VSS.n4394 VSS.n4390 4.5005
R65461 VSS.n5206 VSS.n4381 4.5005
R65462 VSS.n5204 VSS.n4381 4.5005
R65463 VSS.n4394 VSS.n4381 4.5005
R65464 VSS.n5205 VSS.n4394 4.5005
R65465 VSS.n5205 VSS.n4397 4.5005
R65466 VSS.n5206 VSS.n5205 4.5005
R65467 VSS.n5205 VSS.n5204 4.5005
R65468 VSS.n5177 VSS.n4428 4.5005
R65469 VSS.n4437 VSS.n4428 4.5005
R65470 VSS.n5179 VSS.n4428 4.5005
R65471 VSS.n5177 VSS.n4430 4.5005
R65472 VSS.n5179 VSS.n4430 4.5005
R65473 VSS.n5177 VSS.n4427 4.5005
R65474 VSS.n5179 VSS.n4427 4.5005
R65475 VSS.n5177 VSS.n4431 4.5005
R65476 VSS.n4437 VSS.n4431 4.5005
R65477 VSS.n5179 VSS.n4431 4.5005
R65478 VSS.n5177 VSS.n4426 4.5005
R65479 VSS.n4437 VSS.n4426 4.5005
R65480 VSS.n5179 VSS.n4426 4.5005
R65481 VSS.n5177 VSS.n4432 4.5005
R65482 VSS.n4437 VSS.n4432 4.5005
R65483 VSS.n5179 VSS.n4432 4.5005
R65484 VSS.n5177 VSS.n4425 4.5005
R65485 VSS.n4437 VSS.n4425 4.5005
R65486 VSS.n5179 VSS.n4425 4.5005
R65487 VSS.n5179 VSS.n4433 4.5005
R65488 VSS.n5177 VSS.n4433 4.5005
R65489 VSS.n5179 VSS.n4424 4.5005
R65490 VSS.n5177 VSS.n4424 4.5005
R65491 VSS.n5178 VSS.n5177 4.5005
R65492 VSS.n5178 VSS.n4437 4.5005
R65493 VSS.n5179 VSS.n5178 4.5005
R65494 VSS.n5168 VSS.n4453 4.5005
R65495 VSS.n5171 VSS.n4453 4.5005
R65496 VSS.n4453 VSS.n4448 4.5005
R65497 VSS.n5168 VSS.n5167 4.5005
R65498 VSS.n5167 VSS.n4448 4.5005
R65499 VSS.n5168 VSS.n5126 4.5005
R65500 VSS.n5126 VSS.n4448 4.5005
R65501 VSS.n5168 VSS.n4455 4.5005
R65502 VSS.n5171 VSS.n4455 4.5005
R65503 VSS.n4455 VSS.n4448 4.5005
R65504 VSS.n5168 VSS.n4450 4.5005
R65505 VSS.n5171 VSS.n4450 4.5005
R65506 VSS.n4450 VSS.n4448 4.5005
R65507 VSS.n5168 VSS.n4456 4.5005
R65508 VSS.n5171 VSS.n4456 4.5005
R65509 VSS.n4456 VSS.n4448 4.5005
R65510 VSS.n5168 VSS.n4449 4.5005
R65511 VSS.n5171 VSS.n4449 4.5005
R65512 VSS.n4449 VSS.n4448 4.5005
R65513 VSS.n4448 VSS.n14 4.5005
R65514 VSS.n5168 VSS.n14 4.5005
R65515 VSS.n5169 VSS.n4448 4.5005
R65516 VSS.n5169 VSS.n5168 4.5005
R65517 VSS.n5168 VSS.n16 4.5005
R65518 VSS.n5171 VSS.n16 4.5005
R65519 VSS.n4448 VSS.n16 4.5005
R65520 VSS.n33 VSS.n30 4.5005
R65521 VSS.n34 VSS.n30 4.5005
R65522 VSS.n9889 VSS.n30 4.5005
R65523 VSS.n9892 VSS.n30 4.5005
R65524 VSS.n9893 VSS.n33 4.5005
R65525 VSS.n9893 VSS.n34 4.5005
R65526 VSS.n9893 VSS.n9892 4.5005
R65527 VSS.n40 VSS.n34 4.5005
R65528 VSS.n9892 VSS.n40 4.5005
R65529 VSS.n43 VSS.n34 4.5005
R65530 VSS.n9892 VSS.n43 4.5005
R65531 VSS.n39 VSS.n34 4.5005
R65532 VSS.n9892 VSS.n39 4.5005
R65533 VSS.n9891 VSS.n34 4.5005
R65534 VSS.n9892 VSS.n9891 4.5005
R65535 VSS.n38 VSS.n33 4.5005
R65536 VSS.n38 VSS.n34 4.5005
R65537 VSS.n9892 VSS.n38 4.5005
R65538 VSS.n9892 VSS.n22 4.5005
R65539 VSS.n9889 VSS.n22 4.5005
R65540 VSS.n33 VSS.n22 4.5005
R65541 VSS.n9892 VSS.n37 4.5005
R65542 VSS.n9889 VSS.n37 4.5005
R65543 VSS.n37 VSS.n33 4.5005
R65544 VSS.n33 VSS.n25 4.5005
R65545 VSS.n34 VSS.n25 4.5005
R65546 VSS.n9892 VSS.n25 4.5005
R65547 VSS.n9889 VSS.n25 4.5005
R65548 VSS.n82 VSS.n73 4.5005
R65549 VSS.n85 VSS.n73 4.5005
R65550 VSS.n9862 VSS.n73 4.5005
R65551 VSS.n9864 VSS.n73 4.5005
R65552 VSS.n82 VSS.n75 4.5005
R65553 VSS.n85 VSS.n75 4.5005
R65554 VSS.n9864 VSS.n75 4.5005
R65555 VSS.n85 VSS.n72 4.5005
R65556 VSS.n9864 VSS.n72 4.5005
R65557 VSS.n85 VSS.n76 4.5005
R65558 VSS.n9864 VSS.n76 4.5005
R65559 VSS.n85 VSS.n71 4.5005
R65560 VSS.n9864 VSS.n71 4.5005
R65561 VSS.n85 VSS.n77 4.5005
R65562 VSS.n9864 VSS.n77 4.5005
R65563 VSS.n82 VSS.n70 4.5005
R65564 VSS.n85 VSS.n70 4.5005
R65565 VSS.n9864 VSS.n70 4.5005
R65566 VSS.n9864 VSS.n78 4.5005
R65567 VSS.n9862 VSS.n78 4.5005
R65568 VSS.n82 VSS.n78 4.5005
R65569 VSS.n9864 VSS.n69 4.5005
R65570 VSS.n9862 VSS.n69 4.5005
R65571 VSS.n82 VSS.n69 4.5005
R65572 VSS.n9863 VSS.n82 4.5005
R65573 VSS.n9863 VSS.n85 4.5005
R65574 VSS.n9864 VSS.n9863 4.5005
R65575 VSS.n9863 VSS.n9862 4.5005
R65576 VSS.n146 VSS.n135 4.5005
R65577 VSS.n9822 VSS.n135 4.5005
R65578 VSS.n9832 VSS.n135 4.5005
R65579 VSS.n9834 VSS.n135 4.5005
R65580 VSS.n9822 VSS.n137 4.5005
R65581 VSS.n9832 VSS.n137 4.5005
R65582 VSS.n9834 VSS.n137 4.5005
R65583 VSS.n9822 VSS.n134 4.5005
R65584 VSS.n9834 VSS.n134 4.5005
R65585 VSS.n9822 VSS.n138 4.5005
R65586 VSS.n9834 VSS.n138 4.5005
R65587 VSS.n9822 VSS.n133 4.5005
R65588 VSS.n9834 VSS.n133 4.5005
R65589 VSS.n9822 VSS.n139 4.5005
R65590 VSS.n9834 VSS.n139 4.5005
R65591 VSS.n9822 VSS.n132 4.5005
R65592 VSS.n9832 VSS.n132 4.5005
R65593 VSS.n9834 VSS.n132 4.5005
R65594 VSS.n9799 VSS.n178 4.5005
R65595 VSS.n9799 VSS.n179 4.5005
R65596 VSS.n9809 VSS.n9799 4.5005
R65597 VSS.n184 VSS.n179 4.5005
R65598 VSS.n9809 VSS.n184 4.5005
R65599 VSS.n9802 VSS.n179 4.5005
R65600 VSS.n9809 VSS.n9802 4.5005
R65601 VSS.n183 VSS.n179 4.5005
R65602 VSS.n9809 VSS.n183 4.5005
R65603 VSS.n9805 VSS.n179 4.5005
R65604 VSS.n9809 VSS.n9805 4.5005
R65605 VSS.n182 VSS.n179 4.5005
R65606 VSS.n9809 VSS.n182 4.5005
R65607 VSS.n9807 VSS.n179 4.5005
R65608 VSS.n9807 VSS.n177 4.5005
R65609 VSS.n9809 VSS.n9807 4.5005
R65610 VSS.n9809 VSS.n181 4.5005
R65611 VSS.n181 VSS.n177 4.5005
R65612 VSS.n181 VSS.n179 4.5005
R65613 VSS.n181 VSS.n178 4.5005
R65614 VSS.n9808 VSS.n178 4.5005
R65615 VSS.n9808 VSS.n179 4.5005
R65616 VSS.n9808 VSS.n177 4.5005
R65617 VSS.n9809 VSS.n9808 4.5005
R65618 VSS.n9810 VSS.n178 4.5005
R65619 VSS.n9810 VSS.n179 4.5005
R65620 VSS.n9810 VSS.n177 4.5005
R65621 VSS.n9810 VSS.n9809 4.5005
R65622 VSS.n178 VSS.n172 4.5005
R65623 VSS.n179 VSS.n172 4.5005
R65624 VSS.n177 VSS.n172 4.5005
R65625 VSS.n9809 VSS.n172 4.5005
R65626 VSS.n5438 VSS.n5426 4.5005
R65627 VSS.n5438 VSS.n5431 4.5005
R65628 VSS.n5485 VSS.n5438 4.5005
R65629 VSS.n5482 VSS.n5438 4.5005
R65630 VSS.n5436 VSS.n5426 4.5005
R65631 VSS.n5436 VSS.n5431 4.5005
R65632 VSS.n5485 VSS.n5436 4.5005
R65633 VSS.n5482 VSS.n5436 4.5005
R65634 VSS.n5482 VSS.n5439 4.5005
R65635 VSS.n5485 VSS.n5439 4.5005
R65636 VSS.n5439 VSS.n5431 4.5005
R65637 VSS.n5439 VSS.n5426 4.5005
R65638 VSS.n5482 VSS.n5435 4.5005
R65639 VSS.n5485 VSS.n5435 4.5005
R65640 VSS.n5435 VSS.n5431 4.5005
R65641 VSS.n5435 VSS.n5426 4.5005
R65642 VSS.n5482 VSS.n5475 4.5005
R65643 VSS.n5485 VSS.n5475 4.5005
R65644 VSS.n5475 VSS.n5426 4.5005
R65645 VSS.n5485 VSS.n5434 4.5005
R65646 VSS.n5434 VSS.n5426 4.5005
R65647 VSS.n5485 VSS.n5477 4.5005
R65648 VSS.n5477 VSS.n5426 4.5005
R65649 VSS.n5485 VSS.n5433 4.5005
R65650 VSS.n5433 VSS.n5426 4.5005
R65651 VSS.n5485 VSS.n5479 4.5005
R65652 VSS.n5479 VSS.n5426 4.5005
R65653 VSS.n5485 VSS.n5432 4.5005
R65654 VSS.n5432 VSS.n5426 4.5005
R65655 VSS.n5485 VSS.n5484 4.5005
R65656 VSS.n5484 VSS.n5431 4.5005
R65657 VSS.n5484 VSS.n5426 4.5005
R65658 VSS.n425 VSS.n415 4.5005
R65659 VSS.n9608 VSS.n415 4.5005
R65660 VSS.n415 VSS.n402 4.5005
R65661 VSS.n9608 VSS.n412 4.5005
R65662 VSS.n412 VSS.n402 4.5005
R65663 VSS.n9608 VSS.n417 4.5005
R65664 VSS.n417 VSS.n402 4.5005
R65665 VSS.n9608 VSS.n411 4.5005
R65666 VSS.n411 VSS.n402 4.5005
R65667 VSS.n9608 VSS.n419 4.5005
R65668 VSS.n419 VSS.n402 4.5005
R65669 VSS.n425 VSS.n410 4.5005
R65670 VSS.n9608 VSS.n410 4.5005
R65671 VSS.n410 VSS.n402 4.5005
R65672 VSS.n420 VSS.n402 4.5005
R65673 VSS.n420 VSS.n407 4.5005
R65674 VSS.n9608 VSS.n420 4.5005
R65675 VSS.n425 VSS.n420 4.5005
R65676 VSS.n409 VSS.n402 4.5005
R65677 VSS.n409 VSS.n407 4.5005
R65678 VSS.n9608 VSS.n409 4.5005
R65679 VSS.n425 VSS.n409 4.5005
R65680 VSS.n421 VSS.n402 4.5005
R65681 VSS.n421 VSS.n407 4.5005
R65682 VSS.n9608 VSS.n421 4.5005
R65683 VSS.n425 VSS.n421 4.5005
R65684 VSS.n425 VSS.n408 4.5005
R65685 VSS.n9608 VSS.n408 4.5005
R65686 VSS.n408 VSS.n407 4.5005
R65687 VSS.n408 VSS.n402 4.5005
R65688 VSS.n9607 VSS.n425 4.5005
R65689 VSS.n9608 VSS.n9607 4.5005
R65690 VSS.n9607 VSS.n407 4.5005
R65691 VSS.n9607 VSS.n402 4.5005
R65692 VSS.n9596 VSS.n445 4.5005
R65693 VSS.n9596 VSS.n446 4.5005
R65694 VSS.n9596 VSS.n9595 4.5005
R65695 VSS.n461 VSS.n446 4.5005
R65696 VSS.n9595 VSS.n461 4.5005
R65697 VSS.n458 VSS.n446 4.5005
R65698 VSS.n9595 VSS.n458 4.5005
R65699 VSS.n463 VSS.n446 4.5005
R65700 VSS.n9595 VSS.n463 4.5005
R65701 VSS.n457 VSS.n446 4.5005
R65702 VSS.n9595 VSS.n457 4.5005
R65703 VSS.n465 VSS.n446 4.5005
R65704 VSS.n9595 VSS.n465 4.5005
R65705 VSS.n456 VSS.n446 4.5005
R65706 VSS.n9595 VSS.n456 4.5005
R65707 VSS.n467 VSS.n446 4.5005
R65708 VSS.n9595 VSS.n467 4.5005
R65709 VSS.n455 VSS.n446 4.5005
R65710 VSS.n9595 VSS.n455 4.5005
R65711 VSS.n469 VSS.n446 4.5005
R65712 VSS.n9595 VSS.n469 4.5005
R65713 VSS.n454 VSS.n446 4.5005
R65714 VSS.n9595 VSS.n454 4.5005
R65715 VSS.n471 VSS.n446 4.5005
R65716 VSS.n9595 VSS.n471 4.5005
R65717 VSS.n453 VSS.n446 4.5005
R65718 VSS.n9595 VSS.n453 4.5005
R65719 VSS.n473 VSS.n446 4.5005
R65720 VSS.n9595 VSS.n473 4.5005
R65721 VSS.n452 VSS.n446 4.5005
R65722 VSS.n9595 VSS.n452 4.5005
R65723 VSS.n475 VSS.n446 4.5005
R65724 VSS.n9595 VSS.n475 4.5005
R65725 VSS.n451 VSS.n446 4.5005
R65726 VSS.n9595 VSS.n451 4.5005
R65727 VSS.n477 VSS.n446 4.5005
R65728 VSS.n9595 VSS.n477 4.5005
R65729 VSS.n450 VSS.n446 4.5005
R65730 VSS.n9595 VSS.n450 4.5005
R65731 VSS.n479 VSS.n446 4.5005
R65732 VSS.n9595 VSS.n479 4.5005
R65733 VSS.n449 VSS.n446 4.5005
R65734 VSS.n9595 VSS.n449 4.5005
R65735 VSS.n481 VSS.n446 4.5005
R65736 VSS.n9595 VSS.n481 4.5005
R65737 VSS.n448 VSS.n446 4.5005
R65738 VSS.n9595 VSS.n448 4.5005
R65739 VSS.n9594 VSS.n445 4.5005
R65740 VSS.n9594 VSS.n446 4.5005
R65741 VSS.n9595 VSS.n9594 4.5005
R65742 VSS.n9583 VSS.n502 4.5005
R65743 VSS.n9583 VSS.n503 4.5005
R65744 VSS.n9583 VSS.n9582 4.5005
R65745 VSS.n509 VSS.n503 4.5005
R65746 VSS.n9582 VSS.n509 4.5005
R65747 VSS.n512 VSS.n503 4.5005
R65748 VSS.n9582 VSS.n512 4.5005
R65749 VSS.n508 VSS.n503 4.5005
R65750 VSS.n9582 VSS.n508 4.5005
R65751 VSS.n514 VSS.n503 4.5005
R65752 VSS.n9582 VSS.n514 4.5005
R65753 VSS.n507 VSS.n503 4.5005
R65754 VSS.n9582 VSS.n507 4.5005
R65755 VSS.n516 VSS.n503 4.5005
R65756 VSS.n9582 VSS.n516 4.5005
R65757 VSS.n506 VSS.n503 4.5005
R65758 VSS.n9582 VSS.n506 4.5005
R65759 VSS.n518 VSS.n503 4.5005
R65760 VSS.n9582 VSS.n518 4.5005
R65761 VSS.n505 VSS.n503 4.5005
R65762 VSS.n9582 VSS.n505 4.5005
R65763 VSS.n9581 VSS.n503 4.5005
R65764 VSS.n9581 VSS.n524 4.5005
R65765 VSS.n9582 VSS.n9581 4.5005
R65766 VSS.n9570 VSS.n540 4.5005
R65767 VSS.n9570 VSS.n541 4.5005
R65768 VSS.n9570 VSS.n9569 4.5005
R65769 VSS.n547 VSS.n541 4.5005
R65770 VSS.n9569 VSS.n547 4.5005
R65771 VSS.n550 VSS.n541 4.5005
R65772 VSS.n9569 VSS.n550 4.5005
R65773 VSS.n546 VSS.n541 4.5005
R65774 VSS.n9569 VSS.n546 4.5005
R65775 VSS.n552 VSS.n541 4.5005
R65776 VSS.n9569 VSS.n552 4.5005
R65777 VSS.n545 VSS.n541 4.5005
R65778 VSS.n9569 VSS.n545 4.5005
R65779 VSS.n554 VSS.n541 4.5005
R65780 VSS.n9569 VSS.n554 4.5005
R65781 VSS.n544 VSS.n541 4.5005
R65782 VSS.n9569 VSS.n544 4.5005
R65783 VSS.n556 VSS.n541 4.5005
R65784 VSS.n9569 VSS.n556 4.5005
R65785 VSS.n543 VSS.n541 4.5005
R65786 VSS.n9569 VSS.n543 4.5005
R65787 VSS.n9568 VSS.n541 4.5005
R65788 VSS.n9568 VSS.n562 4.5005
R65789 VSS.n9569 VSS.n9568 4.5005
R65790 VSS.n9567 VSS.n564 4.5005
R65791 VSS.n9567 VSS.n565 4.5005
R65792 VSS.n9567 VSS.n9566 4.5005
R65793 VSS.n580 VSS.n565 4.5005
R65794 VSS.n9566 VSS.n580 4.5005
R65795 VSS.n577 VSS.n565 4.5005
R65796 VSS.n9566 VSS.n577 4.5005
R65797 VSS.n582 VSS.n565 4.5005
R65798 VSS.n9566 VSS.n582 4.5005
R65799 VSS.n576 VSS.n565 4.5005
R65800 VSS.n9566 VSS.n576 4.5005
R65801 VSS.n584 VSS.n565 4.5005
R65802 VSS.n9566 VSS.n584 4.5005
R65803 VSS.n575 VSS.n565 4.5005
R65804 VSS.n9566 VSS.n575 4.5005
R65805 VSS.n586 VSS.n565 4.5005
R65806 VSS.n9566 VSS.n586 4.5005
R65807 VSS.n574 VSS.n565 4.5005
R65808 VSS.n9566 VSS.n574 4.5005
R65809 VSS.n588 VSS.n565 4.5005
R65810 VSS.n9566 VSS.n588 4.5005
R65811 VSS.n573 VSS.n565 4.5005
R65812 VSS.n9566 VSS.n573 4.5005
R65813 VSS.n590 VSS.n565 4.5005
R65814 VSS.n9566 VSS.n590 4.5005
R65815 VSS.n572 VSS.n565 4.5005
R65816 VSS.n9566 VSS.n572 4.5005
R65817 VSS.n592 VSS.n565 4.5005
R65818 VSS.n9566 VSS.n592 4.5005
R65819 VSS.n571 VSS.n565 4.5005
R65820 VSS.n9566 VSS.n571 4.5005
R65821 VSS.n594 VSS.n565 4.5005
R65822 VSS.n9566 VSS.n594 4.5005
R65823 VSS.n570 VSS.n565 4.5005
R65824 VSS.n9566 VSS.n570 4.5005
R65825 VSS.n596 VSS.n565 4.5005
R65826 VSS.n9566 VSS.n596 4.5005
R65827 VSS.n569 VSS.n565 4.5005
R65828 VSS.n9566 VSS.n569 4.5005
R65829 VSS.n598 VSS.n565 4.5005
R65830 VSS.n9566 VSS.n598 4.5005
R65831 VSS.n568 VSS.n565 4.5005
R65832 VSS.n9566 VSS.n568 4.5005
R65833 VSS.n600 VSS.n565 4.5005
R65834 VSS.n9566 VSS.n600 4.5005
R65835 VSS.n567 VSS.n565 4.5005
R65836 VSS.n9566 VSS.n567 4.5005
R65837 VSS.n9565 VSS.n564 4.5005
R65838 VSS.n9565 VSS.n565 4.5005
R65839 VSS.n9566 VSS.n9565 4.5005
R65840 VSS.n9564 VSS.n603 4.5005
R65841 VSS.n9564 VSS.n604 4.5005
R65842 VSS.n9564 VSS.n9563 4.5005
R65843 VSS.n618 VSS.n604 4.5005
R65844 VSS.n9563 VSS.n618 4.5005
R65845 VSS.n615 VSS.n604 4.5005
R65846 VSS.n9563 VSS.n615 4.5005
R65847 VSS.n620 VSS.n604 4.5005
R65848 VSS.n9563 VSS.n620 4.5005
R65849 VSS.n614 VSS.n604 4.5005
R65850 VSS.n9563 VSS.n614 4.5005
R65851 VSS.n622 VSS.n604 4.5005
R65852 VSS.n9563 VSS.n622 4.5005
R65853 VSS.n613 VSS.n604 4.5005
R65854 VSS.n9563 VSS.n613 4.5005
R65855 VSS.n624 VSS.n604 4.5005
R65856 VSS.n9563 VSS.n624 4.5005
R65857 VSS.n612 VSS.n604 4.5005
R65858 VSS.n9563 VSS.n612 4.5005
R65859 VSS.n626 VSS.n604 4.5005
R65860 VSS.n9563 VSS.n626 4.5005
R65861 VSS.n611 VSS.n604 4.5005
R65862 VSS.n9563 VSS.n611 4.5005
R65863 VSS.n628 VSS.n604 4.5005
R65864 VSS.n9563 VSS.n628 4.5005
R65865 VSS.n610 VSS.n604 4.5005
R65866 VSS.n9563 VSS.n610 4.5005
R65867 VSS.n630 VSS.n604 4.5005
R65868 VSS.n9563 VSS.n630 4.5005
R65869 VSS.n609 VSS.n604 4.5005
R65870 VSS.n9563 VSS.n609 4.5005
R65871 VSS.n632 VSS.n604 4.5005
R65872 VSS.n9563 VSS.n632 4.5005
R65873 VSS.n608 VSS.n604 4.5005
R65874 VSS.n9563 VSS.n608 4.5005
R65875 VSS.n634 VSS.n604 4.5005
R65876 VSS.n9563 VSS.n634 4.5005
R65877 VSS.n607 VSS.n604 4.5005
R65878 VSS.n9563 VSS.n607 4.5005
R65879 VSS.n636 VSS.n604 4.5005
R65880 VSS.n9563 VSS.n636 4.5005
R65881 VSS.n606 VSS.n604 4.5005
R65882 VSS.n9563 VSS.n606 4.5005
R65883 VSS.n638 VSS.n604 4.5005
R65884 VSS.n9563 VSS.n638 4.5005
R65885 VSS.n605 VSS.n604 4.5005
R65886 VSS.n9563 VSS.n605 4.5005
R65887 VSS.n9562 VSS.n603 4.5005
R65888 VSS.n9562 VSS.n604 4.5005
R65889 VSS.n9563 VSS.n9562 4.5005
R65890 VSS.n9561 VSS.n641 4.5005
R65891 VSS.n9561 VSS.n642 4.5005
R65892 VSS.n9561 VSS.n9560 4.5005
R65893 VSS.n657 VSS.n642 4.5005
R65894 VSS.n9560 VSS.n657 4.5005
R65895 VSS.n654 VSS.n642 4.5005
R65896 VSS.n9560 VSS.n654 4.5005
R65897 VSS.n659 VSS.n642 4.5005
R65898 VSS.n9560 VSS.n659 4.5005
R65899 VSS.n653 VSS.n642 4.5005
R65900 VSS.n9560 VSS.n653 4.5005
R65901 VSS.n661 VSS.n642 4.5005
R65902 VSS.n9560 VSS.n661 4.5005
R65903 VSS.n652 VSS.n642 4.5005
R65904 VSS.n9560 VSS.n652 4.5005
R65905 VSS.n663 VSS.n642 4.5005
R65906 VSS.n9560 VSS.n663 4.5005
R65907 VSS.n651 VSS.n642 4.5005
R65908 VSS.n9560 VSS.n651 4.5005
R65909 VSS.n665 VSS.n642 4.5005
R65910 VSS.n9560 VSS.n665 4.5005
R65911 VSS.n650 VSS.n642 4.5005
R65912 VSS.n9560 VSS.n650 4.5005
R65913 VSS.n667 VSS.n642 4.5005
R65914 VSS.n9560 VSS.n667 4.5005
R65915 VSS.n649 VSS.n642 4.5005
R65916 VSS.n9560 VSS.n649 4.5005
R65917 VSS.n669 VSS.n642 4.5005
R65918 VSS.n9560 VSS.n669 4.5005
R65919 VSS.n648 VSS.n642 4.5005
R65920 VSS.n9560 VSS.n648 4.5005
R65921 VSS.n671 VSS.n642 4.5005
R65922 VSS.n9560 VSS.n671 4.5005
R65923 VSS.n647 VSS.n642 4.5005
R65924 VSS.n9560 VSS.n647 4.5005
R65925 VSS.n673 VSS.n642 4.5005
R65926 VSS.n9560 VSS.n673 4.5005
R65927 VSS.n646 VSS.n642 4.5005
R65928 VSS.n9560 VSS.n646 4.5005
R65929 VSS.n675 VSS.n642 4.5005
R65930 VSS.n9560 VSS.n675 4.5005
R65931 VSS.n645 VSS.n642 4.5005
R65932 VSS.n9560 VSS.n645 4.5005
R65933 VSS.n677 VSS.n642 4.5005
R65934 VSS.n9560 VSS.n677 4.5005
R65935 VSS.n644 VSS.n642 4.5005
R65936 VSS.n9560 VSS.n644 4.5005
R65937 VSS.n9559 VSS.n641 4.5005
R65938 VSS.n9559 VSS.n642 4.5005
R65939 VSS.n9560 VSS.n9559 4.5005
R65940 VSS.n9834 VSS.n140 4.5005
R65941 VSS.n9832 VSS.n140 4.5005
R65942 VSS.n9822 VSS.n140 4.5005
R65943 VSS.n9834 VSS.n131 4.5005
R65944 VSS.n9832 VSS.n131 4.5005
R65945 VSS.n9822 VSS.n131 4.5005
R65946 VSS.n9833 VSS.n146 4.5005
R65947 VSS.n9833 VSS.n9822 4.5005
R65948 VSS.n9834 VSS.n9833 4.5005
R65949 VSS.n9833 VSS.n9832 4.5005
R65950 VSS.n9816 VSS.n141 4.5005
R65951 VSS.n4639 VSS.n4638 4.5005
R65952 VSS.n4672 VSS.n4671 4.5005
R65953 VSS.n4668 VSS.n4667 4.5005
R65954 VSS.n4664 VSS.n4663 4.5005
R65955 VSS.n4662 VSS.n4661 4.5005
R65956 VSS.n4661 VSS.n11 4.5005
R65957 VSS.n9900 VSS.n13 4.5005
R65958 VSS.n9898 VSS.n13 4.5005
R65959 VSS.n9895 VSS.n9894 4.5005
R65960 VSS.n162 VSS.n161 4.5005
R65961 VSS.n9820 VSS.n9817 4.5005
R65962 VSS.n9818 VSS.n9817 4.5005
R65963 VSS.n4636 VSS.n4604 4.5005
R65964 VSS.n4675 VSS.n4674 4.5005
R65965 VSS.n4670 VSS.n4355 4.5005
R65966 VSS.n4666 VSS.n4395 4.5005
R65967 VSS.n9897 VSS.n20 4.5005
R65968 VSS.n83 VSS.n29 4.5005
R65969 VSS.n9821 VSS.n9820 4.5005
R65970 VSS.n9817 VSS.n9816 4.5005
R65971 VSS.n4636 VSS.n4603 4.5005
R65972 VSS.n4635 VSS.n4603 4.5005
R65973 VSS.n4639 VSS.n4603 4.5005
R65974 VSS.n4674 VSS.n4628 4.5005
R65975 VSS.n4640 VSS.n4628 4.5005
R65976 VSS.n4642 VSS.n4628 4.5005
R65977 VSS.n4641 VSS.n4628 4.5005
R65978 VSS.n4671 VSS.n4628 4.5005
R65979 VSS.n4670 VSS.n4354 4.5005
R65980 VSS.n4644 VSS.n4354 4.5005
R65981 VSS.n4646 VSS.n4354 4.5005
R65982 VSS.n4648 VSS.n4354 4.5005
R65983 VSS.n4667 VSS.n4354 4.5005
R65984 VSS.n4666 VSS.n4391 4.5005
R65985 VSS.n4650 VSS.n4391 4.5005
R65986 VSS.n4652 VSS.n4391 4.5005
R65987 VSS.n4654 VSS.n4391 4.5005
R65988 VSS.n4663 VSS.n4391 4.5005
R65989 VSS.n4662 VSS.n4434 4.5005
R65990 VSS.n4659 VSS.n4434 4.5005
R65991 VSS.n4658 VSS.n4434 4.5005
R65992 VSS.n4434 VSS.n11 4.5005
R65993 VSS.n9900 VSS.n9899 4.5005
R65994 VSS.n9899 VSS.n18 4.5005
R65995 VSS.n9899 VSS.n15 4.5005
R65996 VSS.n9899 VSS.n9898 4.5005
R65997 VSS.n9897 VSS.n9896 4.5005
R65998 VSS.n9896 VSS.n24 4.5005
R65999 VSS.n9896 VSS.n27 4.5005
R66000 VSS.n9896 VSS.n23 4.5005
R66001 VSS.n9896 VSS.n9895 4.5005
R66002 VSS.n79 VSS.n29 4.5005
R66003 VSS.n159 VSS.n79 4.5005
R66004 VSS.n157 VSS.n79 4.5005
R66005 VSS.n155 VSS.n79 4.5005
R66006 VSS.n162 VSS.n79 4.5005
R66007 VSS.n4755 VSS.n4571 4.5005
R66008 VSS.n4753 VSS.n4571 4.5005
R66009 VSS.n5252 VSS.n4322 4.5005
R66010 VSS.n5252 VSS.n5251 4.5005
R66011 VSS.n4519 VSS.n4515 4.5005
R66012 VSS.n5078 VSS.n4515 4.5005
R66013 VSS.n5082 VSS.n5081 4.5005
R66014 VSS.n4974 VSS.n4973 4.5005
R66015 VSS.n9688 VSS.n271 4.5005
R66016 VSS.n9691 VSS.n9688 4.5005
R66017 VSS.n223 VSS.n219 4.5005
R66018 VSS.n9765 VSS.n219 4.5005
R66019 VSS.n9813 VSS.n9812 4.5005
R66020 VSS.n9813 VSS.n173 4.5005
R66021 VSS.n5079 VSS.n4505 4.5005
R66022 VSS.n4971 VSS.n4870 4.5005
R66023 VSS.n9812 VSS.n9811 4.5005
R66024 VSS.n4759 VSS.n4758 4.5005
R66025 VSS.n4755 VSS.n4748 4.5005
R66026 VSS.n4751 VSS.n4748 4.5005
R66027 VSS.n4749 VSS.n4748 4.5005
R66028 VSS.n4753 VSS.n4748 4.5005
R66029 VSS.n4326 VSS.n4322 4.5005
R66030 VSS.n5249 VSS.n4326 4.5005
R66031 VSS.n4328 VSS.n4326 4.5005
R66032 VSS.n5251 VSS.n4326 4.5005
R66033 VSS.n4519 VSS.n4516 4.5005
R66034 VSS.n5076 VSS.n4516 4.5005
R66035 VSS.n4518 VSS.n4516 4.5005
R66036 VSS.n5078 VSS.n4516 4.5005
R66037 VSS.n5079 VSS.n4511 4.5005
R66038 VSS.n4512 VSS.n4511 4.5005
R66039 VSS.n5081 VSS.n4511 4.5005
R66040 VSS.n4971 VSS.n4969 4.5005
R66041 VSS.n4970 VSS.n4969 4.5005
R66042 VSS.n4973 VSS.n4969 4.5005
R66043 VSS.n9689 VSS.n271 4.5005
R66044 VSS.n9689 VSS.n272 4.5005
R66045 VSS.n9689 VSS.n270 4.5005
R66046 VSS.n9691 VSS.n9689 4.5005
R66047 VSS.n223 VSS.n220 4.5005
R66048 VSS.n9763 VSS.n220 4.5005
R66049 VSS.n222 VSS.n220 4.5005
R66050 VSS.n9765 VSS.n220 4.5005
R66051 VSS.n9812 VSS.n171 4.5005
R66052 VSS.n173 VSS.n171 4.5005
R66053 VSS.n4744 VSS.n4743 4.5005
R66054 VSS.n4760 VSS.n4743 4.5005
R66055 VSS.n4760 VSS.n4742 4.5005
R66056 VSS.n4760 VSS.n4759 4.5005
R66057 VSS.n9812 VSS.n170 4.5005
R66058 VSS.n173 VSS.n170 4.5005
R66059 VSS.n4755 VSS.n4746 4.5005
R66060 VSS.n4751 VSS.n4746 4.5005
R66061 VSS.n4749 VSS.n4746 4.5005
R66062 VSS.n4753 VSS.n4746 4.5005
R66063 VSS.n4323 VSS.n4322 4.5005
R66064 VSS.n5249 VSS.n4323 4.5005
R66065 VSS.n4328 VSS.n4323 4.5005
R66066 VSS.n5251 VSS.n4323 4.5005
R66067 VSS.n4519 VSS.n4513 4.5005
R66068 VSS.n5076 VSS.n4513 4.5005
R66069 VSS.n4518 VSS.n4513 4.5005
R66070 VSS.n5078 VSS.n4513 4.5005
R66071 VSS.n5079 VSS.n4508 4.5005
R66072 VSS.n4512 VSS.n4508 4.5005
R66073 VSS.n5081 VSS.n4508 4.5005
R66074 VSS.n4971 VSS.n4967 4.5005
R66075 VSS.n4970 VSS.n4967 4.5005
R66076 VSS.n4973 VSS.n4967 4.5005
R66077 VSS.n9692 VSS.n271 4.5005
R66078 VSS.n9692 VSS.n272 4.5005
R66079 VSS.n9692 VSS.n270 4.5005
R66080 VSS.n9692 VSS.n9691 4.5005
R66081 VSS.n223 VSS.n217 4.5005
R66082 VSS.n9763 VSS.n217 4.5005
R66083 VSS.n222 VSS.n217 4.5005
R66084 VSS.n9765 VSS.n217 4.5005
R66085 VSS.n9814 VSS.n170 4.5005
R66086 VSS.n4755 VSS.n4754 4.5005
R66087 VSS.n4754 VSS.n4751 4.5005
R66088 VSS.n4754 VSS.n4749 4.5005
R66089 VSS.n4754 VSS.n4753 4.5005
R66090 VSS.n5250 VSS.n4322 4.5005
R66091 VSS.n5250 VSS.n5249 4.5005
R66092 VSS.n5250 VSS.n4328 4.5005
R66093 VSS.n5251 VSS.n5250 4.5005
R66094 VSS.n5077 VSS.n4519 4.5005
R66095 VSS.n5077 VSS.n5076 4.5005
R66096 VSS.n5077 VSS.n4518 4.5005
R66097 VSS.n5078 VSS.n5077 4.5005
R66098 VSS.n5080 VSS.n5079 4.5005
R66099 VSS.n5080 VSS.n4512 4.5005
R66100 VSS.n5081 VSS.n5080 4.5005
R66101 VSS.n4972 VSS.n4971 4.5005
R66102 VSS.n4972 VSS.n4970 4.5005
R66103 VSS.n4973 VSS.n4972 4.5005
R66104 VSS.n9690 VSS.n271 4.5005
R66105 VSS.n9690 VSS.n272 4.5005
R66106 VSS.n9690 VSS.n270 4.5005
R66107 VSS.n9691 VSS.n9690 4.5005
R66108 VSS.n9764 VSS.n223 4.5005
R66109 VSS.n9764 VSS.n9763 4.5005
R66110 VSS.n9764 VSS.n222 4.5005
R66111 VSS.n9765 VSS.n9764 4.5005
R66112 VSS.n9814 VSS.n169 4.5005
R66113 VSS.n9814 VSS.n171 4.5005
R66114 VSS.n4759 VSS.n4727 4.5005
R66115 VSS.n4742 VSS.n4727 4.5005
R66116 VSS.n4743 VSS.n4727 4.5005
R66117 VSS.n4759 VSS.n4730 4.5005
R66118 VSS.n4742 VSS.n4730 4.5005
R66119 VSS.n4743 VSS.n4730 4.5005
R66120 VSS.n9814 VSS.n9813 4.5005
R66121 VSS.n5263 VSS.n4319 4.5005
R66122 VSS.n5263 VSS.n5262 4.5005
R66123 VSS.n4286 VSS.n4282 4.5005
R66124 VSS.n5648 VSS.n4282 4.5005
R66125 VSS.n5653 VSS.n5652 4.5005
R66126 VSS.n4921 VSS.n4918 4.5005
R66127 VSS.n285 VSS.n279 4.5005
R66128 VSS.n9686 VSS.n285 4.5005
R66129 VSS.n5451 VSS.n5448 4.5005
R66130 VSS.n5457 VSS.n5448 4.5005
R66131 VSS.n5473 VSS.n5466 4.5005
R66132 VSS.n5473 VSS.n5440 4.5005
R66133 VSS.n4565 VSS.n4564 4.5005
R66134 VSS.n4569 VSS.n4565 4.5005
R66135 VSS.n5650 VSS.n5649 4.5005
R66136 VSS.n4915 VSS.n4914 4.5005
R66137 VSS.n5467 VSS.n5466 4.5005
R66138 VSS.n6251 VSS.n6250 4.5005
R66139 VSS.n4567 VSS.n4564 4.5005
R66140 VSS.n4569 VSS.n4567 4.5005
R66141 VSS.n5256 VSS.n4319 4.5005
R66142 VSS.n5260 VSS.n5256 4.5005
R66143 VSS.n5257 VSS.n5256 4.5005
R66144 VSS.n5262 VSS.n5256 4.5005
R66145 VSS.n4286 VSS.n4283 4.5005
R66146 VSS.n5646 VSS.n4283 4.5005
R66147 VSS.n4285 VSS.n4283 4.5005
R66148 VSS.n5648 VSS.n4283 4.5005
R66149 VSS.n5650 VSS.n4278 4.5005
R66150 VSS.n4279 VSS.n4278 4.5005
R66151 VSS.n5652 VSS.n4278 4.5005
R66152 VSS.n4919 VSS.n4914 4.5005
R66153 VSS.n4919 VSS.n4913 4.5005
R66154 VSS.n4921 VSS.n4919 4.5005
R66155 VSS.n286 VSS.n279 4.5005
R66156 VSS.n286 VSS.n281 4.5005
R66157 VSS.n286 VSS.n278 4.5005
R66158 VSS.n9686 VSS.n286 4.5005
R66159 VSS.n5451 VSS.n5449 4.5005
R66160 VSS.n5455 VSS.n5449 4.5005
R66161 VSS.n5450 VSS.n5449 4.5005
R66162 VSS.n5457 VSS.n5449 4.5005
R66163 VSS.n5471 VSS.n5466 4.5005
R66164 VSS.n5471 VSS.n5440 4.5005
R66165 VSS.n6253 VSS.n3857 4.5005
R66166 VSS.n6253 VSS.n3859 4.5005
R66167 VSS.n3861 VSS.n3859 4.5005
R66168 VSS.n6251 VSS.n3859 4.5005
R66169 VSS.n5466 VSS.n174 4.5005
R66170 VSS.n5440 VSS.n174 4.5005
R66171 VSS.n4570 VSS.n4564 4.5005
R66172 VSS.n4570 VSS.n4569 4.5005
R66173 VSS.n5253 VSS.n4319 4.5005
R66174 VSS.n5260 VSS.n5253 4.5005
R66175 VSS.n5257 VSS.n5253 4.5005
R66176 VSS.n5262 VSS.n5253 4.5005
R66177 VSS.n4286 VSS.n4280 4.5005
R66178 VSS.n5646 VSS.n4280 4.5005
R66179 VSS.n4285 VSS.n4280 4.5005
R66180 VSS.n5648 VSS.n4280 4.5005
R66181 VSS.n5650 VSS.n4275 4.5005
R66182 VSS.n4279 VSS.n4275 4.5005
R66183 VSS.n5652 VSS.n4275 4.5005
R66184 VSS.n4922 VSS.n4914 4.5005
R66185 VSS.n4922 VSS.n4913 4.5005
R66186 VSS.n4922 VSS.n4921 4.5005
R66187 VSS.n9687 VSS.n279 4.5005
R66188 VSS.n9687 VSS.n281 4.5005
R66189 VSS.n9687 VSS.n278 4.5005
R66190 VSS.n9687 VSS.n9686 4.5005
R66191 VSS.n5451 VSS.n5446 4.5005
R66192 VSS.n5455 VSS.n5446 4.5005
R66193 VSS.n5450 VSS.n5446 4.5005
R66194 VSS.n5457 VSS.n5446 4.5005
R66195 VSS.n5472 VSS.n174 4.5005
R66196 VSS.n4568 VSS.n4564 4.5005
R66197 VSS.n4569 VSS.n4568 4.5005
R66198 VSS.n5261 VSS.n4319 4.5005
R66199 VSS.n5261 VSS.n5260 4.5005
R66200 VSS.n5261 VSS.n5257 4.5005
R66201 VSS.n5262 VSS.n5261 4.5005
R66202 VSS.n5647 VSS.n4286 4.5005
R66203 VSS.n5647 VSS.n5646 4.5005
R66204 VSS.n5647 VSS.n4285 4.5005
R66205 VSS.n5648 VSS.n5647 4.5005
R66206 VSS.n5651 VSS.n5650 4.5005
R66207 VSS.n5651 VSS.n4279 4.5005
R66208 VSS.n5652 VSS.n5651 4.5005
R66209 VSS.n4920 VSS.n4914 4.5005
R66210 VSS.n4920 VSS.n4913 4.5005
R66211 VSS.n4921 VSS.n4920 4.5005
R66212 VSS.n9685 VSS.n279 4.5005
R66213 VSS.n9685 VSS.n281 4.5005
R66214 VSS.n9685 VSS.n278 4.5005
R66215 VSS.n9686 VSS.n9685 4.5005
R66216 VSS.n5456 VSS.n5451 4.5005
R66217 VSS.n5456 VSS.n5455 4.5005
R66218 VSS.n5456 VSS.n5450 4.5005
R66219 VSS.n5457 VSS.n5456 4.5005
R66220 VSS.n5472 VSS.n5470 4.5005
R66221 VSS.n5472 VSS.n5471 4.5005
R66222 VSS.n6251 VSS.n3856 4.5005
R66223 VSS.n3861 VSS.n3856 4.5005
R66224 VSS.n6253 VSS.n3856 4.5005
R66225 VSS.n6252 VSS.n6251 4.5005
R66226 VSS.n6252 VSS.n3861 4.5005
R66227 VSS.n6253 VSS.n6252 4.5005
R66228 VSS.n5473 VSS.n5472 4.5005
R66229 VSS.n4096 VSS.n3950 4.5005
R66230 VSS.n4102 VSS.n3950 4.5005
R66231 VSS.n4104 VSS.n3995 4.5005
R66232 VSS.n4110 VSS.n3995 4.5005
R66233 VSS.n4115 VSS.n4027 4.5005
R66234 VSS.n5726 VSS.n5725 4.5005
R66235 VSS.n4168 VSS.n324 4.5005
R66236 VSS.n4166 VSS.n324 4.5005
R66237 VSS.n4164 VSS.n357 4.5005
R66238 VSS.n4162 VSS.n357 4.5005
R66239 VSS.n4157 VSS.n422 4.5005
R66240 VSS.n4151 VSS.n422 4.5005
R66241 VSS.n4093 VSS.n4089 4.5005
R66242 VSS.n4095 VSS.n4089 4.5005
R66243 VSS.n4113 VSS.n4111 4.5005
R66244 VSS.n5728 VSS.n4117 4.5005
R66245 VSS.n4157 VSS.n4149 4.5005
R66246 VSS.n3854 VSS.n3852 4.5005
R66247 VSS.n4093 VSS.n4091 4.5005
R66248 VSS.n4095 VSS.n4091 4.5005
R66249 VSS.n4096 VSS.n4086 4.5005
R66250 VSS.n4100 VSS.n4086 4.5005
R66251 VSS.n4087 VSS.n4086 4.5005
R66252 VSS.n4102 VSS.n4086 4.5005
R66253 VSS.n4104 VSS.n4082 4.5005
R66254 VSS.n4108 VSS.n4082 4.5005
R66255 VSS.n4083 VSS.n4082 4.5005
R66256 VSS.n4110 VSS.n4082 4.5005
R66257 VSS.n4113 VSS.n4078 4.5005
R66258 VSS.n4079 VSS.n4078 4.5005
R66259 VSS.n4115 VSS.n4078 4.5005
R66260 VSS.n5728 VSS.n4119 4.5005
R66261 VSS.n4121 VSS.n4119 4.5005
R66262 VSS.n5726 VSS.n4119 4.5005
R66263 VSS.n4168 VSS.n4126 4.5005
R66264 VSS.n4129 VSS.n4126 4.5005
R66265 VSS.n4127 VSS.n4126 4.5005
R66266 VSS.n4166 VSS.n4126 4.5005
R66267 VSS.n4164 VSS.n4134 4.5005
R66268 VSS.n4137 VSS.n4134 4.5005
R66269 VSS.n4135 VSS.n4134 4.5005
R66270 VSS.n4162 VSS.n4134 4.5005
R66271 VSS.n4157 VSS.n4150 4.5005
R66272 VSS.n4151 VSS.n4150 4.5005
R66273 VSS.n6260 VSS.n6257 4.5005
R66274 VSS.n6260 VSS.n6259 4.5005
R66275 VSS.n6259 VSS.n3853 4.5005
R66276 VSS.n6259 VSS.n3854 4.5005
R66277 VSS.n4157 VSS.n4156 4.5005
R66278 VSS.n4156 VSS.n4151 4.5005
R66279 VSS.n4093 VSS.n4088 4.5005
R66280 VSS.n4095 VSS.n4088 4.5005
R66281 VSS.n4096 VSS.n4084 4.5005
R66282 VSS.n4100 VSS.n4084 4.5005
R66283 VSS.n4087 VSS.n4084 4.5005
R66284 VSS.n4102 VSS.n4084 4.5005
R66285 VSS.n4104 VSS.n4080 4.5005
R66286 VSS.n4108 VSS.n4080 4.5005
R66287 VSS.n4083 VSS.n4080 4.5005
R66288 VSS.n4110 VSS.n4080 4.5005
R66289 VSS.n4113 VSS.n4076 4.5005
R66290 VSS.n4079 VSS.n4076 4.5005
R66291 VSS.n4115 VSS.n4076 4.5005
R66292 VSS.n5728 VSS.n4116 4.5005
R66293 VSS.n4121 VSS.n4116 4.5005
R66294 VSS.n5726 VSS.n4116 4.5005
R66295 VSS.n4168 VSS.n4124 4.5005
R66296 VSS.n4129 VSS.n4124 4.5005
R66297 VSS.n4127 VSS.n4124 4.5005
R66298 VSS.n4166 VSS.n4124 4.5005
R66299 VSS.n4164 VSS.n4132 4.5005
R66300 VSS.n4137 VSS.n4132 4.5005
R66301 VSS.n4135 VSS.n4132 4.5005
R66302 VSS.n4162 VSS.n4132 4.5005
R66303 VSS.n4156 VSS.n4155 4.5005
R66304 VSS.n4094 VSS.n4093 4.5005
R66305 VSS.n4095 VSS.n4094 4.5005
R66306 VSS.n4101 VSS.n4096 4.5005
R66307 VSS.n4101 VSS.n4100 4.5005
R66308 VSS.n4101 VSS.n4087 4.5005
R66309 VSS.n4102 VSS.n4101 4.5005
R66310 VSS.n4109 VSS.n4104 4.5005
R66311 VSS.n4109 VSS.n4108 4.5005
R66312 VSS.n4109 VSS.n4083 4.5005
R66313 VSS.n4110 VSS.n4109 4.5005
R66314 VSS.n4114 VSS.n4113 4.5005
R66315 VSS.n4114 VSS.n4079 4.5005
R66316 VSS.n4115 VSS.n4114 4.5005
R66317 VSS.n5728 VSS.n5727 4.5005
R66318 VSS.n5727 VSS.n4121 4.5005
R66319 VSS.n5727 VSS.n5726 4.5005
R66320 VSS.n4168 VSS.n4167 4.5005
R66321 VSS.n4167 VSS.n4129 4.5005
R66322 VSS.n4167 VSS.n4127 4.5005
R66323 VSS.n4167 VSS.n4166 4.5005
R66324 VSS.n4164 VSS.n4163 4.5005
R66325 VSS.n4163 VSS.n4137 4.5005
R66326 VSS.n4163 VSS.n4135 4.5005
R66327 VSS.n4163 VSS.n4162 4.5005
R66328 VSS.n4155 VSS.n4153 4.5005
R66329 VSS.n4155 VSS.n4150 4.5005
R66330 VSS.n6261 VSS.n3854 4.5005
R66331 VSS.n6261 VSS.n3853 4.5005
R66332 VSS.n6261 VSS.n6260 4.5005
R66333 VSS.n3854 VSS.n3832 4.5005
R66334 VSS.n3853 VSS.n3832 4.5005
R66335 VSS.n6260 VSS.n3832 4.5005
R66336 VSS.n4155 VSS.n422 4.5005
R66337 VSS.n6062 VSS.n6056 4.5005
R66338 VSS.n6068 VSS.n6049 4.5005
R66339 VSS.n6075 VSS.n6041 4.5005
R66340 VSS.n6076 VSS.n6036 4.5005
R66341 VSS.n6079 VSS.n6036 4.5005
R66342 VSS.n5958 VSS.n5903 4.5005
R66343 VSS.n5958 VSS.n5957 4.5005
R66344 VSS.n5949 VSS.n5947 4.5005
R66345 VSS.n5941 VSS.n5939 4.5005
R66346 VSS.n9602 VSS.n426 4.5005
R66347 VSS.n6066 VSS.n6047 4.5005
R66348 VSS.n6068 VSS.n6047 4.5005
R66349 VSS.n6073 VSS.n6039 4.5005
R66350 VSS.n6075 VSS.n6039 4.5005
R66351 VSS.n6079 VSS.n4072 4.5005
R66352 VSS.n5957 VSS.n5909 4.5005
R66353 VSS.n5916 VSS.n5913 4.5005
R66354 VSS.n5949 VSS.n5916 4.5005
R66355 VSS.n5923 VSS.n5920 4.5005
R66356 VSS.n5941 VSS.n5923 4.5005
R66357 VSS.n6271 VSS.n3829 4.5005
R66358 VSS.n6066 VSS.n6050 4.5005
R66359 VSS.n6068 VSS.n6050 4.5005
R66360 VSS.n6073 VSS.n6042 4.5005
R66361 VSS.n6075 VSS.n6042 4.5005
R66362 VSS.n6079 VSS.n6078 4.5005
R66363 VSS.n5957 VSS.n5956 4.5005
R66364 VSS.n5948 VSS.n5913 4.5005
R66365 VSS.n5949 VSS.n5948 4.5005
R66366 VSS.n5940 VSS.n5920 4.5005
R66367 VSS.n5941 VSS.n5940 4.5005
R66368 VSS.n9605 VSS.n9604 4.5005
R66369 VSS.n9604 VSS.n426 4.5005
R66370 VSS.n6269 VSS.n3829 4.5005
R66371 VSS.n9606 VSS.n9605 4.5005
R66372 VSS.n9606 VSS.n426 4.5005
R66373 VSS.n6068 VSS.n3952 4.5005
R66374 VSS.n6075 VSS.n3996 4.5005
R66375 VSS.n5949 VSS.n325 4.5005
R66376 VSS.n5941 VSS.n359 4.5005
R66377 VSS.n6062 VSS.n6061 4.5005
R66378 VSS.n6067 VSS.n6066 4.5005
R66379 VSS.n6068 VSS.n6067 4.5005
R66380 VSS.n6074 VSS.n6073 4.5005
R66381 VSS.n6075 VSS.n6074 4.5005
R66382 VSS.n6076 VSS.n4070 4.5005
R66383 VSS.n5953 VSS.n5903 4.5005
R66384 VSS.n5950 VSS.n5913 4.5005
R66385 VSS.n5950 VSS.n5949 4.5005
R66386 VSS.n5942 VSS.n5920 4.5005
R66387 VSS.n5942 VSS.n5941 4.5005
R66388 VSS.n9604 VSS.n9603 4.5005
R66389 VSS.n6268 VSS.n3829 4.5005
R66390 VSS.n6274 VSS.n3829 4.5005
R66391 VSS.n6274 VSS.n6273 4.5005
R66392 VSS.n9603 VSS.n9602 4.5005
R66393 VSS.n6288 VSS.n3820 4.5005
R66394 VSS.n6294 VSS.n3813 4.5005
R66395 VSS.n6301 VSS.n3804 4.5005
R66396 VSS.n6302 VSS.n3798 4.5005
R66397 VSS.n6305 VSS.n3798 4.5005
R66398 VSS.n6314 VSS.n3709 4.5005
R66399 VSS.n6317 VSS.n3709 4.5005
R66400 VSS.n6323 VSS.n3700 4.5005
R66401 VSS.n6330 VSS.n3691 4.5005
R66402 VSS.n9597 VSS.n435 4.5005
R66403 VSS.n6292 VSS.n3811 4.5005
R66404 VSS.n6294 VSS.n3811 4.5005
R66405 VSS.n6299 VSS.n3802 4.5005
R66406 VSS.n6301 VSS.n3802 4.5005
R66407 VSS.n6305 VSS.n3718 4.5005
R66408 VSS.n6317 VSS.n3707 4.5005
R66409 VSS.n6321 VSS.n3698 4.5005
R66410 VSS.n6323 VSS.n3698 4.5005
R66411 VSS.n6328 VSS.n3689 4.5005
R66412 VSS.n6330 VSS.n3689 4.5005
R66413 VSS.n6282 VSS.n3824 4.5005
R66414 VSS.n6292 VSS.n3814 4.5005
R66415 VSS.n6294 VSS.n3814 4.5005
R66416 VSS.n6299 VSS.n3805 4.5005
R66417 VSS.n6301 VSS.n3805 4.5005
R66418 VSS.n6305 VSS.n6304 4.5005
R66419 VSS.n6317 VSS.n6316 4.5005
R66420 VSS.n6321 VSS.n3701 4.5005
R66421 VSS.n6323 VSS.n3701 4.5005
R66422 VSS.n6328 VSS.n3692 4.5005
R66423 VSS.n6330 VSS.n3692 4.5005
R66424 VSS.n9600 VSS.n9599 4.5005
R66425 VSS.n9599 VSS.n435 4.5005
R66426 VSS.n6282 VSS.n3823 4.5005
R66427 VSS.n9601 VSS.n9600 4.5005
R66428 VSS.n9601 VSS.n435 4.5005
R66429 VSS.n6294 VSS.n3810 4.5005
R66430 VSS.n6301 VSS.n3801 4.5005
R66431 VSS.n6323 VSS.n3697 4.5005
R66432 VSS.n6330 VSS.n3688 4.5005
R66433 VSS.n6288 VSS.n6287 4.5005
R66434 VSS.n6293 VSS.n6292 4.5005
R66435 VSS.n6294 VSS.n6293 4.5005
R66436 VSS.n6300 VSS.n6299 4.5005
R66437 VSS.n6301 VSS.n6300 4.5005
R66438 VSS.n6302 VSS.n3716 4.5005
R66439 VSS.n6314 VSS.n6313 4.5005
R66440 VSS.n6322 VSS.n6321 4.5005
R66441 VSS.n6323 VSS.n6322 4.5005
R66442 VSS.n6329 VSS.n6328 4.5005
R66443 VSS.n6330 VSS.n6329 4.5005
R66444 VSS.n9599 VSS.n9598 4.5005
R66445 VSS.n6282 VSS.n3822 4.5005
R66446 VSS.n6282 VSS.n6281 4.5005
R66447 VSS.n6281 VSS.n6280 4.5005
R66448 VSS.n9598 VSS.n9597 4.5005
R66449 VSS.n6588 VSS.n3219 4.5005
R66450 VSS.n6594 VSS.n3210 4.5005
R66451 VSS.n6601 VSS.n3201 4.5005
R66452 VSS.n6602 VSS.n3195 4.5005
R66453 VSS.n6605 VSS.n3195 4.5005
R66454 VSS.n6620 VSS.n3131 4.5005
R66455 VSS.n6623 VSS.n3131 4.5005
R66456 VSS.n6629 VSS.n2966 4.5005
R66457 VSS.n6639 VSS.n6638 4.5005
R66458 VSS.n9589 VSS.n483 4.5005
R66459 VSS.n6586 VSS.n3217 4.5005
R66460 VSS.n6588 VSS.n3217 4.5005
R66461 VSS.n6592 VSS.n3208 4.5005
R66462 VSS.n6594 VSS.n3208 4.5005
R66463 VSS.n6599 VSS.n3199 4.5005
R66464 VSS.n6601 VSS.n3199 4.5005
R66465 VSS.n6605 VSS.n3193 4.5005
R66466 VSS.n6623 VSS.n3129 4.5005
R66467 VSS.n6627 VSS.n3122 4.5005
R66468 VSS.n6629 VSS.n3122 4.5005
R66469 VSS.n6636 VSS.n3117 4.5005
R66470 VSS.n6638 VSS.n3117 4.5005
R66471 VSS.n6581 VSS.n3226 4.5005
R66472 VSS.n6586 VSS.n3220 4.5005
R66473 VSS.n6588 VSS.n3220 4.5005
R66474 VSS.n6592 VSS.n3211 4.5005
R66475 VSS.n6594 VSS.n3211 4.5005
R66476 VSS.n6599 VSS.n3202 4.5005
R66477 VSS.n6601 VSS.n3202 4.5005
R66478 VSS.n6605 VSS.n6604 4.5005
R66479 VSS.n6623 VSS.n6622 4.5005
R66480 VSS.n6627 VSS.n3123 4.5005
R66481 VSS.n6629 VSS.n3123 4.5005
R66482 VSS.n6636 VSS.n3118 4.5005
R66483 VSS.n6638 VSS.n3118 4.5005
R66484 VSS.n9592 VSS.n9591 4.5005
R66485 VSS.n9591 VSS.n483 4.5005
R66486 VSS.n6581 VSS.n3225 4.5005
R66487 VSS.n9593 VSS.n9592 4.5005
R66488 VSS.n9593 VSS.n483 4.5005
R66489 VSS.n6588 VSS.n3216 4.5005
R66490 VSS.n6594 VSS.n3207 4.5005
R66491 VSS.n6601 VSS.n3198 4.5005
R66492 VSS.n6629 VSS.n3120 4.5005
R66493 VSS.n6638 VSS.n3116 4.5005
R66494 VSS.n6587 VSS.n6586 4.5005
R66495 VSS.n6588 VSS.n6587 4.5005
R66496 VSS.n6593 VSS.n6592 4.5005
R66497 VSS.n6594 VSS.n6593 4.5005
R66498 VSS.n6600 VSS.n6599 4.5005
R66499 VSS.n6601 VSS.n6600 4.5005
R66500 VSS.n6602 VSS.n3191 4.5005
R66501 VSS.n6620 VSS.n6619 4.5005
R66502 VSS.n6628 VSS.n6627 4.5005
R66503 VSS.n6629 VSS.n6628 4.5005
R66504 VSS.n6637 VSS.n6636 4.5005
R66505 VSS.n6638 VSS.n6637 4.5005
R66506 VSS.n9591 VSS.n9590 4.5005
R66507 VSS.n6581 VSS.n3224 4.5005
R66508 VSS.n6581 VSS.n6580 4.5005
R66509 VSS.n6580 VSS.n6579 4.5005
R66510 VSS.n9590 VSS.n9589 4.5005
R66511 VSS.n5786 VSS.n5762 4.5005
R66512 VSS.n5792 VSS.n5753 4.5005
R66513 VSS.n5799 VSS.n5744 4.5005
R66514 VSS.n5888 VSS.n5738 4.5005
R66515 VSS.n5891 VSS.n5738 4.5005
R66516 VSS.n6766 VSS.n2959 4.5005
R66517 VSS.n6766 VSS.n6765 4.5005
R66518 VSS.n6757 VSS.n6753 4.5005
R66519 VSS.n6653 VSS.n6643 4.5005
R66520 VSS.n9584 VSS.n492 4.5005
R66521 VSS.n5784 VSS.n5760 4.5005
R66522 VSS.n5786 VSS.n5760 4.5005
R66523 VSS.n5790 VSS.n5751 4.5005
R66524 VSS.n5792 VSS.n5751 4.5005
R66525 VSS.n5797 VSS.n5742 4.5005
R66526 VSS.n5799 VSS.n5742 4.5005
R66527 VSS.n5891 VSS.n5736 4.5005
R66528 VSS.n6765 VSS.n2962 4.5005
R66529 VSS.n6755 VSS.n2969 4.5005
R66530 VSS.n6757 VSS.n2969 4.5005
R66531 VSS.n6651 VSS.n6641 4.5005
R66532 VSS.n6653 VSS.n6641 4.5005
R66533 VSS.n5779 VSS.n5769 4.5005
R66534 VSS.n5784 VSS.n5763 4.5005
R66535 VSS.n5786 VSS.n5763 4.5005
R66536 VSS.n5790 VSS.n5754 4.5005
R66537 VSS.n5792 VSS.n5754 4.5005
R66538 VSS.n5797 VSS.n5745 4.5005
R66539 VSS.n5799 VSS.n5745 4.5005
R66540 VSS.n5891 VSS.n5890 4.5005
R66541 VSS.n6765 VSS.n6764 4.5005
R66542 VSS.n6756 VSS.n6755 4.5005
R66543 VSS.n6757 VSS.n6756 4.5005
R66544 VSS.n6651 VSS.n6644 4.5005
R66545 VSS.n6653 VSS.n6644 4.5005
R66546 VSS.n9587 VSS.n9586 4.5005
R66547 VSS.n9586 VSS.n492 4.5005
R66548 VSS.n5779 VSS.n5768 4.5005
R66549 VSS.n9588 VSS.n9587 4.5005
R66550 VSS.n9588 VSS.n492 4.5005
R66551 VSS.n5786 VSS.n5759 4.5005
R66552 VSS.n5792 VSS.n5750 4.5005
R66553 VSS.n5799 VSS.n5741 4.5005
R66554 VSS.n6758 VSS.n6757 4.5005
R66555 VSS.n6653 VSS.n6640 4.5005
R66556 VSS.n5785 VSS.n5784 4.5005
R66557 VSS.n5786 VSS.n5785 4.5005
R66558 VSS.n5791 VSS.n5790 4.5005
R66559 VSS.n5792 VSS.n5791 4.5005
R66560 VSS.n5798 VSS.n5797 4.5005
R66561 VSS.n5799 VSS.n5798 4.5005
R66562 VSS.n5888 VSS.n5887 4.5005
R66563 VSS.n6761 VSS.n2959 4.5005
R66564 VSS.n6755 VSS.n2965 4.5005
R66565 VSS.n6757 VSS.n2965 4.5005
R66566 VSS.n6652 VSS.n6651 4.5005
R66567 VSS.n6653 VSS.n6652 4.5005
R66568 VSS.n9586 VSS.n9585 4.5005
R66569 VSS.n5779 VSS.n5767 4.5005
R66570 VSS.n5779 VSS.n5778 4.5005
R66571 VSS.n5778 VSS.n5777 4.5005
R66572 VSS.n9585 VSS.n9584 4.5005
R66573 VSS.n6980 VSS.n2763 4.5005
R66574 VSS.n6986 VSS.n2754 4.5005
R66575 VSS.n6993 VSS.n2745 4.5005
R66576 VSS.n6994 VSS.n2739 4.5005
R66577 VSS.n6997 VSS.n2739 4.5005
R66578 VSS.n7006 VSS.n2647 4.5005
R66579 VSS.n7009 VSS.n2647 4.5005
R66580 VSS.n7015 VSS.n2638 4.5005
R66581 VSS.n7022 VSS.n2629 4.5005
R66582 VSS.n9576 VSS.n525 4.5005
R66583 VSS.n6978 VSS.n2761 4.5005
R66584 VSS.n6980 VSS.n2761 4.5005
R66585 VSS.n6984 VSS.n2752 4.5005
R66586 VSS.n6986 VSS.n2752 4.5005
R66587 VSS.n6991 VSS.n2743 4.5005
R66588 VSS.n6993 VSS.n2743 4.5005
R66589 VSS.n6997 VSS.n2656 4.5005
R66590 VSS.n7009 VSS.n2645 4.5005
R66591 VSS.n7013 VSS.n2636 4.5005
R66592 VSS.n7015 VSS.n2636 4.5005
R66593 VSS.n7020 VSS.n2627 4.5005
R66594 VSS.n7022 VSS.n2627 4.5005
R66595 VSS.n6973 VSS.n2770 4.5005
R66596 VSS.n6978 VSS.n2764 4.5005
R66597 VSS.n6980 VSS.n2764 4.5005
R66598 VSS.n6984 VSS.n2755 4.5005
R66599 VSS.n6986 VSS.n2755 4.5005
R66600 VSS.n6991 VSS.n2746 4.5005
R66601 VSS.n6993 VSS.n2746 4.5005
R66602 VSS.n6997 VSS.n6996 4.5005
R66603 VSS.n7009 VSS.n7008 4.5005
R66604 VSS.n7013 VSS.n2639 4.5005
R66605 VSS.n7015 VSS.n2639 4.5005
R66606 VSS.n7020 VSS.n2630 4.5005
R66607 VSS.n7022 VSS.n2630 4.5005
R66608 VSS.n9579 VSS.n9578 4.5005
R66609 VSS.n9578 VSS.n525 4.5005
R66610 VSS.n6973 VSS.n2769 4.5005
R66611 VSS.n9580 VSS.n9579 4.5005
R66612 VSS.n9580 VSS.n525 4.5005
R66613 VSS.n6980 VSS.n2760 4.5005
R66614 VSS.n6986 VSS.n2751 4.5005
R66615 VSS.n6993 VSS.n2742 4.5005
R66616 VSS.n7015 VSS.n2635 4.5005
R66617 VSS.n7022 VSS.n2626 4.5005
R66618 VSS.n6979 VSS.n6978 4.5005
R66619 VSS.n6980 VSS.n6979 4.5005
R66620 VSS.n6985 VSS.n6984 4.5005
R66621 VSS.n6986 VSS.n6985 4.5005
R66622 VSS.n6992 VSS.n6991 4.5005
R66623 VSS.n6993 VSS.n6992 4.5005
R66624 VSS.n6994 VSS.n2654 4.5005
R66625 VSS.n7006 VSS.n7005 4.5005
R66626 VSS.n7014 VSS.n7013 4.5005
R66627 VSS.n7015 VSS.n7014 4.5005
R66628 VSS.n7021 VSS.n7020 4.5005
R66629 VSS.n7022 VSS.n7021 4.5005
R66630 VSS.n9578 VSS.n9577 4.5005
R66631 VSS.n6973 VSS.n2768 4.5005
R66632 VSS.n6973 VSS.n6972 4.5005
R66633 VSS.n6972 VSS.n6971 4.5005
R66634 VSS.n9577 VSS.n9576 4.5005
R66635 VSS.n7046 VSS.n7045 4.5005
R66636 VSS.n7045 VSS.n2611 4.5005
R66637 VSS.n7045 VSS.n7044 4.5005
R66638 VSS.n2617 VSS.n2611 4.5005
R66639 VSS.n7044 VSS.n2617 4.5005
R66640 VSS.n9575 VSS.n9574 4.5005
R66641 VSS.n9575 VSS.n534 4.5005
R66642 VSS.n9574 VSS.n9573 4.5005
R66643 VSS.n7047 VSS.n2611 4.5005
R66644 VSS.n7047 VSS.n7046 4.5005
R66645 VSS.n7041 VSS.n7040 4.5005
R66646 VSS.n7034 VSS.n7032 4.5005
R66647 VSS.n7040 VSS.n7032 4.5005
R66648 VSS.n7031 VSS.n7030 4.5005
R66649 VSS.n7028 VSS.n2623 4.5005
R66650 VSS.n7030 VSS.n2623 4.5005
R66651 VSS.n7028 VSS.n2624 4.5005
R66652 VSS.n7030 VSS.n2624 4.5005
R66653 VSS.n6662 VSS.n6661 4.5005
R66654 VSS.n6659 VSS.n3110 4.5005
R66655 VSS.n6661 VSS.n3110 4.5005
R66656 VSS.n6659 VSS.n3111 4.5005
R66657 VSS.n6661 VSS.n3111 4.5005
R66658 VSS.n3667 VSS.n3659 4.5005
R66659 VSS.n3665 VSS.n3657 4.5005
R66660 VSS.n3667 VSS.n3657 4.5005
R66661 VSS.n3665 VSS.n3660 4.5005
R66662 VSS.n3667 VSS.n3660 4.5005
R66663 VSS.n6339 VSS.n6338 4.5005
R66664 VSS.n6336 VSS.n3685 4.5005
R66665 VSS.n6338 VSS.n3685 4.5005
R66666 VSS.n6336 VSS.n3686 4.5005
R66667 VSS.n6338 VSS.n3686 4.5005
R66668 VSS.n5934 VSS.n5932 4.5005
R66669 VSS.n5930 VSS.n5927 4.5005
R66670 VSS.n5934 VSS.n5930 4.5005
R66671 VSS.n5933 VSS.n5927 4.5005
R66672 VSS.n5934 VSS.n5933 4.5005
R66673 VSS.n4161 VSS.n396 4.5005
R66674 VSS.n4159 VSS.n396 4.5005
R66675 VSS.n4161 VSS.n4142 4.5005
R66676 VSS.n4145 VSS.n4142 4.5005
R66677 VSS.n4143 VSS.n4142 4.5005
R66678 VSS.n4159 VSS.n4142 4.5005
R66679 VSS.n5458 VSS.n5443 4.5005
R66680 VSS.n5464 VSS.n5443 4.5005
R66681 VSS.n5458 VSS.n5444 4.5005
R66682 VSS.n5462 VSS.n5444 4.5005
R66683 VSS.n5445 VSS.n5444 4.5005
R66684 VSS.n5464 VSS.n5444 4.5005
R66685 VSS.n9766 VSS.n205 4.5005
R66686 VSS.n9773 VSS.n205 4.5005
R66687 VSS.n9771 VSS.n9766 4.5005
R66688 VSS.n9771 VSS.n9769 4.5005
R66689 VSS.n9771 VSS.n216 4.5005
R66690 VSS.n9773 VSS.n9771 4.5005
R66691 VSS.n166 VSS.n165 4.5005
R66692 VSS.n163 VSS.n114 4.5005
R66693 VSS.n9774 VSS.n9766 4.5005
R66694 VSS.n9774 VSS.n9769 4.5005
R66695 VSS.n9774 VSS.n216 4.5005
R66696 VSS.n9774 VSS.n9773 4.5005
R66697 VSS.n9772 VSS.n9766 4.5005
R66698 VSS.n9772 VSS.n9769 4.5005
R66699 VSS.n9772 VSS.n216 4.5005
R66700 VSS.n9773 VSS.n9772 4.5005
R66701 VSS.n5458 VSS.n5441 4.5005
R66702 VSS.n5462 VSS.n5441 4.5005
R66703 VSS.n5445 VSS.n5441 4.5005
R66704 VSS.n5464 VSS.n5441 4.5005
R66705 VSS.n5463 VSS.n5458 4.5005
R66706 VSS.n5463 VSS.n5462 4.5005
R66707 VSS.n5463 VSS.n5445 4.5005
R66708 VSS.n5464 VSS.n5463 4.5005
R66709 VSS.n4161 VSS.n4140 4.5005
R66710 VSS.n4145 VSS.n4140 4.5005
R66711 VSS.n4143 VSS.n4140 4.5005
R66712 VSS.n4159 VSS.n4140 4.5005
R66713 VSS.n4161 VSS.n4160 4.5005
R66714 VSS.n4160 VSS.n4145 4.5005
R66715 VSS.n4160 VSS.n4143 4.5005
R66716 VSS.n4160 VSS.n4159 4.5005
R66717 VSS.n5934 VSS.n397 4.5005
R66718 VSS.n5935 VSS.n5927 4.5005
R66719 VSS.n5935 VSS.n5934 4.5005
R66720 VSS.n6338 VSS.n3684 4.5005
R66721 VSS.n6337 VSS.n6336 4.5005
R66722 VSS.n6338 VSS.n6337 4.5005
R66723 VSS.n3668 VSS.n3667 4.5005
R66724 VSS.n3666 VSS.n3665 4.5005
R66725 VSS.n3667 VSS.n3666 4.5005
R66726 VSS.n6661 VSS.n3109 4.5005
R66727 VSS.n6660 VSS.n6659 4.5005
R66728 VSS.n6661 VSS.n6660 4.5005
R66729 VSS.n7030 VSS.n2622 4.5005
R66730 VSS.n7029 VSS.n7028 4.5005
R66731 VSS.n7030 VSS.n7029 4.5005
R66732 VSS.n7040 VSS.n7039 4.5005
R66733 VSS.n7039 VSS.n7038 4.5005
R66734 VSS.n163 VSS.n110 4.5005
R66735 VSS.n113 VSS.n104 4.5005
R66736 VSS.n116 VSS.n104 4.5005
R66737 VSS.n9847 VSS.n104 4.5005
R66738 VSS.n9849 VSS.n104 4.5005
R66739 VSS.n113 VSS.n106 4.5005
R66740 VSS.n116 VSS.n106 4.5005
R66741 VSS.n9849 VSS.n106 4.5005
R66742 VSS.n116 VSS.n103 4.5005
R66743 VSS.n9849 VSS.n103 4.5005
R66744 VSS.n116 VSS.n107 4.5005
R66745 VSS.n9849 VSS.n107 4.5005
R66746 VSS.n116 VSS.n102 4.5005
R66747 VSS.n9849 VSS.n102 4.5005
R66748 VSS.n116 VSS.n108 4.5005
R66749 VSS.n9849 VSS.n108 4.5005
R66750 VSS.n113 VSS.n101 4.5005
R66751 VSS.n116 VSS.n101 4.5005
R66752 VSS.n9849 VSS.n101 4.5005
R66753 VSS.n9778 VSS.n197 4.5005
R66754 VSS.n197 VSS.n194 4.5005
R66755 VSS.n9776 VSS.n197 4.5005
R66756 VSS.n210 VSS.n194 4.5005
R66757 VSS.n9776 VSS.n210 4.5005
R66758 VSS.n213 VSS.n194 4.5005
R66759 VSS.n9776 VSS.n213 4.5005
R66760 VSS.n208 VSS.n194 4.5005
R66761 VSS.n9776 VSS.n208 4.5005
R66762 VSS.n215 VSS.n194 4.5005
R66763 VSS.n9776 VSS.n215 4.5005
R66764 VSS.n207 VSS.n194 4.5005
R66765 VSS.n9776 VSS.n207 4.5005
R66766 VSS.n9775 VSS.n194 4.5005
R66767 VSS.n9775 VSS.n204 4.5005
R66768 VSS.n9776 VSS.n9775 4.5005
R66769 VSS.n9778 VSS.n196 4.5005
R66770 VSS.n196 VSS.n194 4.5005
R66771 VSS.n204 VSS.n196 4.5005
R66772 VSS.n9776 VSS.n196 4.5005
R66773 VSS.n9778 VSS.n201 4.5005
R66774 VSS.n201 VSS.n194 4.5005
R66775 VSS.n204 VSS.n201 4.5005
R66776 VSS.n9776 VSS.n201 4.5005
R66777 VSS.n9778 VSS.n195 4.5005
R66778 VSS.n195 VSS.n194 4.5005
R66779 VSS.n204 VSS.n195 4.5005
R66780 VSS.n9776 VSS.n195 4.5005
R66781 VSS.n9778 VSS.n9777 4.5005
R66782 VSS.n9777 VSS.n194 4.5005
R66783 VSS.n9777 VSS.n204 4.5005
R66784 VSS.n9777 VSS.n9776 4.5005
R66785 VSS.n5503 VSS.n5414 4.5005
R66786 VSS.n5506 VSS.n5414 4.5005
R66787 VSS.n5414 VSS.n5407 4.5005
R66788 VSS.n5414 VSS.n5402 4.5005
R66789 VSS.n5503 VSS.n5412 4.5005
R66790 VSS.n5506 VSS.n5412 4.5005
R66791 VSS.n5412 VSS.n5407 4.5005
R66792 VSS.n5412 VSS.n5402 4.5005
R66793 VSS.n5503 VSS.n5415 4.5005
R66794 VSS.n5506 VSS.n5415 4.5005
R66795 VSS.n5415 VSS.n5407 4.5005
R66796 VSS.n5415 VSS.n5402 4.5005
R66797 VSS.n5503 VSS.n5411 4.5005
R66798 VSS.n5506 VSS.n5411 4.5005
R66799 VSS.n5411 VSS.n5407 4.5005
R66800 VSS.n5411 VSS.n5402 4.5005
R66801 VSS.n5503 VSS.n5417 4.5005
R66802 VSS.n5506 VSS.n5417 4.5005
R66803 VSS.n5417 VSS.n5402 4.5005
R66804 VSS.n5506 VSS.n5410 4.5005
R66805 VSS.n5410 VSS.n5402 4.5005
R66806 VSS.n5506 VSS.n5419 4.5005
R66807 VSS.n5419 VSS.n5402 4.5005
R66808 VSS.n5506 VSS.n5409 4.5005
R66809 VSS.n5409 VSS.n5402 4.5005
R66810 VSS.n5506 VSS.n5421 4.5005
R66811 VSS.n5421 VSS.n5402 4.5005
R66812 VSS.n5506 VSS.n5408 4.5005
R66813 VSS.n5408 VSS.n5402 4.5005
R66814 VSS.n5506 VSS.n5505 4.5005
R66815 VSS.n5505 VSS.n5407 4.5005
R66816 VSS.n5505 VSS.n5402 4.5005
R66817 VSS.n9626 VSS.n389 4.5005
R66818 VSS.n9628 VSS.n389 4.5005
R66819 VSS.n389 VSS.n376 4.5005
R66820 VSS.n9628 VSS.n386 4.5005
R66821 VSS.n386 VSS.n376 4.5005
R66822 VSS.n9628 VSS.n391 4.5005
R66823 VSS.n391 VSS.n376 4.5005
R66824 VSS.n9628 VSS.n385 4.5005
R66825 VSS.n385 VSS.n376 4.5005
R66826 VSS.n9628 VSS.n393 4.5005
R66827 VSS.n393 VSS.n376 4.5005
R66828 VSS.n9626 VSS.n384 4.5005
R66829 VSS.n9628 VSS.n384 4.5005
R66830 VSS.n384 VSS.n376 4.5005
R66831 VSS.n394 VSS.n376 4.5005
R66832 VSS.n394 VSS.n381 4.5005
R66833 VSS.n9628 VSS.n394 4.5005
R66834 VSS.n9626 VSS.n394 4.5005
R66835 VSS.n383 VSS.n376 4.5005
R66836 VSS.n383 VSS.n381 4.5005
R66837 VSS.n9628 VSS.n383 4.5005
R66838 VSS.n9626 VSS.n383 4.5005
R66839 VSS.n395 VSS.n376 4.5005
R66840 VSS.n395 VSS.n381 4.5005
R66841 VSS.n9628 VSS.n395 4.5005
R66842 VSS.n9626 VSS.n395 4.5005
R66843 VSS.n382 VSS.n376 4.5005
R66844 VSS.n382 VSS.n381 4.5005
R66845 VSS.n9628 VSS.n382 4.5005
R66846 VSS.n9626 VSS.n382 4.5005
R66847 VSS.n9627 VSS.n376 4.5005
R66848 VSS.n9627 VSS.n381 4.5005
R66849 VSS.n9628 VSS.n9627 4.5005
R66850 VSS.n9627 VSS.n9626 4.5005
R66851 VSS.n6396 VSS.n6340 4.5005
R66852 VSS.n6400 VSS.n6340 4.5005
R66853 VSS.n6340 VSS.n3637 4.5005
R66854 VSS.n6400 VSS.n6342 4.5005
R66855 VSS.n6342 VSS.n3637 4.5005
R66856 VSS.n6400 VSS.n3680 4.5005
R66857 VSS.n3680 VSS.n3637 4.5005
R66858 VSS.n6400 VSS.n6343 4.5005
R66859 VSS.n6343 VSS.n3637 4.5005
R66860 VSS.n6400 VSS.n3679 4.5005
R66861 VSS.n3679 VSS.n3637 4.5005
R66862 VSS.n6400 VSS.n6344 4.5005
R66863 VSS.n6344 VSS.n3637 4.5005
R66864 VSS.n6400 VSS.n3678 4.5005
R66865 VSS.n3678 VSS.n3637 4.5005
R66866 VSS.n6400 VSS.n6345 4.5005
R66867 VSS.n6345 VSS.n3637 4.5005
R66868 VSS.n6400 VSS.n3677 4.5005
R66869 VSS.n3677 VSS.n3637 4.5005
R66870 VSS.n6400 VSS.n6346 4.5005
R66871 VSS.n6346 VSS.n3637 4.5005
R66872 VSS.n6400 VSS.n3676 4.5005
R66873 VSS.n3676 VSS.n3637 4.5005
R66874 VSS.n6400 VSS.n6347 4.5005
R66875 VSS.n6347 VSS.n3637 4.5005
R66876 VSS.n6400 VSS.n3675 4.5005
R66877 VSS.n3675 VSS.n3637 4.5005
R66878 VSS.n6400 VSS.n6348 4.5005
R66879 VSS.n6348 VSS.n3637 4.5005
R66880 VSS.n6400 VSS.n3674 4.5005
R66881 VSS.n3674 VSS.n3637 4.5005
R66882 VSS.n6400 VSS.n6349 4.5005
R66883 VSS.n6349 VSS.n3637 4.5005
R66884 VSS.n6400 VSS.n3673 4.5005
R66885 VSS.n3673 VSS.n3637 4.5005
R66886 VSS.n6400 VSS.n6350 4.5005
R66887 VSS.n6350 VSS.n3637 4.5005
R66888 VSS.n6400 VSS.n3672 4.5005
R66889 VSS.n3672 VSS.n3637 4.5005
R66890 VSS.n6400 VSS.n6398 4.5005
R66891 VSS.n6398 VSS.n3637 4.5005
R66892 VSS.n6400 VSS.n3671 4.5005
R66893 VSS.n3671 VSS.n3637 4.5005
R66894 VSS.n6400 VSS.n6399 4.5005
R66895 VSS.n6399 VSS.n3637 4.5005
R66896 VSS.n6401 VSS.n6400 4.5005
R66897 VSS.n6401 VSS.n3637 4.5005
R66898 VSS.n6396 VSS.n3669 4.5005
R66899 VSS.n6400 VSS.n3669 4.5005
R66900 VSS.n3669 VSS.n3637 4.5005
R66901 VSS.n6694 VSS.n6663 4.5005
R66902 VSS.n6697 VSS.n6663 4.5005
R66903 VSS.n6663 VSS.n3092 4.5005
R66904 VSS.n6697 VSS.n3104 4.5005
R66905 VSS.n3104 VSS.n3092 4.5005
R66906 VSS.n6697 VSS.n6664 4.5005
R66907 VSS.n6664 VSS.n3092 4.5005
R66908 VSS.n6697 VSS.n3103 4.5005
R66909 VSS.n3103 VSS.n3092 4.5005
R66910 VSS.n6697 VSS.n6665 4.5005
R66911 VSS.n6665 VSS.n3092 4.5005
R66912 VSS.n6697 VSS.n3102 4.5005
R66913 VSS.n3102 VSS.n3092 4.5005
R66914 VSS.n6697 VSS.n6666 4.5005
R66915 VSS.n6666 VSS.n3092 4.5005
R66916 VSS.n6697 VSS.n3101 4.5005
R66917 VSS.n3101 VSS.n3092 4.5005
R66918 VSS.n6697 VSS.n6696 4.5005
R66919 VSS.n6696 VSS.n3092 4.5005
R66920 VSS.n6697 VSS.n3100 4.5005
R66921 VSS.n3100 VSS.n3092 4.5005
R66922 VSS.n6698 VSS.n6697 4.5005
R66923 VSS.n6699 VSS.n6698 4.5005
R66924 VSS.n6698 VSS.n3092 4.5005
R66925 VSS.n8905 VSS.n1269 4.5005
R66926 VSS.n1269 VSS.n1260 4.5005
R66927 VSS.n8909 VSS.n1269 4.5005
R66928 VSS.n1266 VSS.n1260 4.5005
R66929 VSS.n8909 VSS.n1266 4.5005
R66930 VSS.n1271 VSS.n1260 4.5005
R66931 VSS.n8909 VSS.n1271 4.5005
R66932 VSS.n1265 VSS.n1260 4.5005
R66933 VSS.n8909 VSS.n1265 4.5005
R66934 VSS.n1273 VSS.n1260 4.5005
R66935 VSS.n8909 VSS.n1273 4.5005
R66936 VSS.n1264 VSS.n1260 4.5005
R66937 VSS.n8909 VSS.n1264 4.5005
R66938 VSS.n1275 VSS.n1260 4.5005
R66939 VSS.n8909 VSS.n1275 4.5005
R66940 VSS.n1263 VSS.n1260 4.5005
R66941 VSS.n8909 VSS.n1263 4.5005
R66942 VSS.n8908 VSS.n1260 4.5005
R66943 VSS.n8909 VSS.n8908 4.5005
R66944 VSS.n1262 VSS.n1260 4.5005
R66945 VSS.n8909 VSS.n1262 4.5005
R66946 VSS.n8910 VSS.n1260 4.5005
R66947 VSS.n8910 VSS.n1259 4.5005
R66948 VSS.n8910 VSS.n8909 4.5005
R66949 VSS.n8948 VSS.n8911 4.5005
R66950 VSS.n8911 VSS.n1165 4.5005
R66951 VSS.n8911 VSS.n1150 4.5005
R66952 VSS.n1256 VSS.n1165 4.5005
R66953 VSS.n1256 VSS.n1150 4.5005
R66954 VSS.n1255 VSS.n1165 4.5005
R66955 VSS.n1255 VSS.n1150 4.5005
R66956 VSS.n1253 VSS.n1165 4.5005
R66957 VSS.n1253 VSS.n1150 4.5005
R66958 VSS.n1252 VSS.n1165 4.5005
R66959 VSS.n1252 VSS.n1150 4.5005
R66960 VSS.n1250 VSS.n1165 4.5005
R66961 VSS.n1250 VSS.n1150 4.5005
R66962 VSS.n1249 VSS.n1165 4.5005
R66963 VSS.n1249 VSS.n1150 4.5005
R66964 VSS.n1247 VSS.n1165 4.5005
R66965 VSS.n1247 VSS.n1150 4.5005
R66966 VSS.n1246 VSS.n1165 4.5005
R66967 VSS.n1246 VSS.n1150 4.5005
R66968 VSS.n1244 VSS.n1165 4.5005
R66969 VSS.n1244 VSS.n1150 4.5005
R66970 VSS.n1243 VSS.n1165 4.5005
R66971 VSS.n1243 VSS.n1150 4.5005
R66972 VSS.n1241 VSS.n1165 4.5005
R66973 VSS.n1241 VSS.n1150 4.5005
R66974 VSS.n1240 VSS.n1165 4.5005
R66975 VSS.n1240 VSS.n1150 4.5005
R66976 VSS.n1238 VSS.n1165 4.5005
R66977 VSS.n1238 VSS.n1150 4.5005
R66978 VSS.n1237 VSS.n1165 4.5005
R66979 VSS.n1237 VSS.n1150 4.5005
R66980 VSS.n1235 VSS.n1165 4.5005
R66981 VSS.n1235 VSS.n1150 4.5005
R66982 VSS.n1234 VSS.n1165 4.5005
R66983 VSS.n1234 VSS.n1150 4.5005
R66984 VSS.n1232 VSS.n1165 4.5005
R66985 VSS.n1232 VSS.n1150 4.5005
R66986 VSS.n1231 VSS.n1165 4.5005
R66987 VSS.n1231 VSS.n1150 4.5005
R66988 VSS.n1229 VSS.n1165 4.5005
R66989 VSS.n1229 VSS.n1150 4.5005
R66990 VSS.n1228 VSS.n1165 4.5005
R66991 VSS.n1228 VSS.n1150 4.5005
R66992 VSS.n1226 VSS.n1165 4.5005
R66993 VSS.n1226 VSS.n1150 4.5005
R66994 VSS.n1165 VSS.n1151 4.5005
R66995 VSS.n8950 VSS.n1151 4.5005
R66996 VSS.n1151 VSS.n1150 4.5005
R66997 VSS.n8949 VSS.n1150 4.5005
R66998 VSS.n8950 VSS.n8949 4.5005
R66999 VSS.n8949 VSS.n1165 4.5005
R67000 VSS.n8949 VSS.n8948 4.5005
R67001 VSS.n741 VSS.n729 4.5005
R67002 VSS.n9499 VSS.n741 4.5005
R67003 VSS.n9497 VSS.n741 4.5005
R67004 VSS.n755 VSS.n741 4.5005
R67005 VSS.n755 VSS.n743 4.5005
R67006 VSS.n9497 VSS.n743 4.5005
R67007 VSS.n9499 VSS.n743 4.5005
R67008 VSS.n743 VSS.n729 4.5005
R67009 VSS.n755 VSS.n740 4.5005
R67010 VSS.n9497 VSS.n740 4.5005
R67011 VSS.n9499 VSS.n740 4.5005
R67012 VSS.n740 VSS.n729 4.5005
R67013 VSS.n755 VSS.n744 4.5005
R67014 VSS.n9497 VSS.n744 4.5005
R67015 VSS.n9499 VSS.n744 4.5005
R67016 VSS.n744 VSS.n729 4.5005
R67017 VSS.n755 VSS.n739 4.5005
R67018 VSS.n9497 VSS.n739 4.5005
R67019 VSS.n9499 VSS.n739 4.5005
R67020 VSS.n739 VSS.n729 4.5005
R67021 VSS.n745 VSS.n729 4.5005
R67022 VSS.n9499 VSS.n745 4.5005
R67023 VSS.n9497 VSS.n745 4.5005
R67024 VSS.n755 VSS.n745 4.5005
R67025 VSS.n738 VSS.n729 4.5005
R67026 VSS.n9499 VSS.n738 4.5005
R67027 VSS.n9497 VSS.n738 4.5005
R67028 VSS.n755 VSS.n738 4.5005
R67029 VSS.n746 VSS.n729 4.5005
R67030 VSS.n9499 VSS.n746 4.5005
R67031 VSS.n9497 VSS.n746 4.5005
R67032 VSS.n755 VSS.n746 4.5005
R67033 VSS.n755 VSS.n737 4.5005
R67034 VSS.n9497 VSS.n737 4.5005
R67035 VSS.n9499 VSS.n737 4.5005
R67036 VSS.n737 VSS.n729 4.5005
R67037 VSS.n755 VSS.n747 4.5005
R67038 VSS.n9497 VSS.n747 4.5005
R67039 VSS.n9499 VSS.n747 4.5005
R67040 VSS.n747 VSS.n729 4.5005
R67041 VSS.n755 VSS.n736 4.5005
R67042 VSS.n9497 VSS.n736 4.5005
R67043 VSS.n9499 VSS.n736 4.5005
R67044 VSS.n736 VSS.n729 4.5005
R67045 VSS.n755 VSS.n748 4.5005
R67046 VSS.n9497 VSS.n748 4.5005
R67047 VSS.n9499 VSS.n748 4.5005
R67048 VSS.n748 VSS.n729 4.5005
R67049 VSS.n735 VSS.n729 4.5005
R67050 VSS.n9499 VSS.n735 4.5005
R67051 VSS.n9497 VSS.n735 4.5005
R67052 VSS.n755 VSS.n735 4.5005
R67053 VSS.n749 VSS.n729 4.5005
R67054 VSS.n9499 VSS.n749 4.5005
R67055 VSS.n9497 VSS.n749 4.5005
R67056 VSS.n755 VSS.n749 4.5005
R67057 VSS.n734 VSS.n729 4.5005
R67058 VSS.n9499 VSS.n734 4.5005
R67059 VSS.n9497 VSS.n734 4.5005
R67060 VSS.n755 VSS.n734 4.5005
R67061 VSS.n755 VSS.n750 4.5005
R67062 VSS.n9497 VSS.n750 4.5005
R67063 VSS.n9499 VSS.n750 4.5005
R67064 VSS.n750 VSS.n729 4.5005
R67065 VSS.n755 VSS.n733 4.5005
R67066 VSS.n9497 VSS.n733 4.5005
R67067 VSS.n9499 VSS.n733 4.5005
R67068 VSS.n733 VSS.n729 4.5005
R67069 VSS.n755 VSS.n751 4.5005
R67070 VSS.n9497 VSS.n751 4.5005
R67071 VSS.n9499 VSS.n751 4.5005
R67072 VSS.n751 VSS.n729 4.5005
R67073 VSS.n732 VSS.n729 4.5005
R67074 VSS.n9499 VSS.n732 4.5005
R67075 VSS.n9497 VSS.n732 4.5005
R67076 VSS.n755 VSS.n732 4.5005
R67077 VSS.n752 VSS.n729 4.5005
R67078 VSS.n9499 VSS.n752 4.5005
R67079 VSS.n9497 VSS.n752 4.5005
R67080 VSS.n755 VSS.n752 4.5005
R67081 VSS.n731 VSS.n729 4.5005
R67082 VSS.n9499 VSS.n731 4.5005
R67083 VSS.n9497 VSS.n731 4.5005
R67084 VSS.n755 VSS.n731 4.5005
R67085 VSS.n753 VSS.n729 4.5005
R67086 VSS.n9499 VSS.n753 4.5005
R67087 VSS.n9497 VSS.n753 4.5005
R67088 VSS.n755 VSS.n753 4.5005
R67089 VSS.n755 VSS.n730 4.5005
R67090 VSS.n9497 VSS.n730 4.5005
R67091 VSS.n9499 VSS.n730 4.5005
R67092 VSS.n730 VSS.n729 4.5005
R67093 VSS.n9498 VSS.n755 4.5005
R67094 VSS.n9498 VSS.n9497 4.5005
R67095 VSS.n9499 VSS.n9498 4.5005
R67096 VSS.n9498 VSS.n729 4.5005
R67097 VSS.n9526 VSS.n697 4.5005
R67098 VSS.n697 VSS.n685 4.5005
R67099 VSS.n9524 VSS.n697 4.5005
R67100 VSS.n710 VSS.n697 4.5005
R67101 VSS.n710 VSS.n698 4.5005
R67102 VSS.n9524 VSS.n698 4.5005
R67103 VSS.n698 VSS.n685 4.5005
R67104 VSS.n9526 VSS.n698 4.5005
R67105 VSS.n710 VSS.n696 4.5005
R67106 VSS.n9524 VSS.n696 4.5005
R67107 VSS.n696 VSS.n685 4.5005
R67108 VSS.n9526 VSS.n696 4.5005
R67109 VSS.n710 VSS.n699 4.5005
R67110 VSS.n9524 VSS.n699 4.5005
R67111 VSS.n699 VSS.n685 4.5005
R67112 VSS.n9526 VSS.n699 4.5005
R67113 VSS.n9526 VSS.n695 4.5005
R67114 VSS.n695 VSS.n685 4.5005
R67115 VSS.n9524 VSS.n695 4.5005
R67116 VSS.n710 VSS.n695 4.5005
R67117 VSS.n9526 VSS.n700 4.5005
R67118 VSS.n700 VSS.n685 4.5005
R67119 VSS.n9524 VSS.n700 4.5005
R67120 VSS.n710 VSS.n700 4.5005
R67121 VSS.n9526 VSS.n694 4.5005
R67122 VSS.n694 VSS.n685 4.5005
R67123 VSS.n9524 VSS.n694 4.5005
R67124 VSS.n710 VSS.n694 4.5005
R67125 VSS.n710 VSS.n701 4.5005
R67126 VSS.n9524 VSS.n701 4.5005
R67127 VSS.n701 VSS.n685 4.5005
R67128 VSS.n9526 VSS.n701 4.5005
R67129 VSS.n710 VSS.n693 4.5005
R67130 VSS.n9524 VSS.n693 4.5005
R67131 VSS.n693 VSS.n685 4.5005
R67132 VSS.n9526 VSS.n693 4.5005
R67133 VSS.n710 VSS.n702 4.5005
R67134 VSS.n9524 VSS.n702 4.5005
R67135 VSS.n702 VSS.n685 4.5005
R67136 VSS.n9526 VSS.n702 4.5005
R67137 VSS.n710 VSS.n692 4.5005
R67138 VSS.n9524 VSS.n692 4.5005
R67139 VSS.n692 VSS.n685 4.5005
R67140 VSS.n9526 VSS.n692 4.5005
R67141 VSS.n9526 VSS.n703 4.5005
R67142 VSS.n703 VSS.n685 4.5005
R67143 VSS.n9524 VSS.n703 4.5005
R67144 VSS.n710 VSS.n703 4.5005
R67145 VSS.n9526 VSS.n691 4.5005
R67146 VSS.n691 VSS.n685 4.5005
R67147 VSS.n9524 VSS.n691 4.5005
R67148 VSS.n710 VSS.n691 4.5005
R67149 VSS.n9526 VSS.n704 4.5005
R67150 VSS.n704 VSS.n685 4.5005
R67151 VSS.n9524 VSS.n704 4.5005
R67152 VSS.n710 VSS.n704 4.5005
R67153 VSS.n710 VSS.n690 4.5005
R67154 VSS.n9524 VSS.n690 4.5005
R67155 VSS.n690 VSS.n685 4.5005
R67156 VSS.n9526 VSS.n690 4.5005
R67157 VSS.n710 VSS.n705 4.5005
R67158 VSS.n9524 VSS.n705 4.5005
R67159 VSS.n705 VSS.n685 4.5005
R67160 VSS.n9526 VSS.n705 4.5005
R67161 VSS.n710 VSS.n689 4.5005
R67162 VSS.n9524 VSS.n689 4.5005
R67163 VSS.n689 VSS.n685 4.5005
R67164 VSS.n9526 VSS.n689 4.5005
R67165 VSS.n9526 VSS.n706 4.5005
R67166 VSS.n706 VSS.n685 4.5005
R67167 VSS.n9524 VSS.n706 4.5005
R67168 VSS.n710 VSS.n706 4.5005
R67169 VSS.n9526 VSS.n688 4.5005
R67170 VSS.n688 VSS.n685 4.5005
R67171 VSS.n9524 VSS.n688 4.5005
R67172 VSS.n710 VSS.n688 4.5005
R67173 VSS.n9526 VSS.n707 4.5005
R67174 VSS.n707 VSS.n685 4.5005
R67175 VSS.n9524 VSS.n707 4.5005
R67176 VSS.n710 VSS.n707 4.5005
R67177 VSS.n9526 VSS.n687 4.5005
R67178 VSS.n687 VSS.n685 4.5005
R67179 VSS.n9524 VSS.n687 4.5005
R67180 VSS.n710 VSS.n687 4.5005
R67181 VSS.n710 VSS.n708 4.5005
R67182 VSS.n9524 VSS.n708 4.5005
R67183 VSS.n708 VSS.n685 4.5005
R67184 VSS.n9526 VSS.n708 4.5005
R67185 VSS.n710 VSS.n686 4.5005
R67186 VSS.n9524 VSS.n686 4.5005
R67187 VSS.n686 VSS.n685 4.5005
R67188 VSS.n9526 VSS.n686 4.5005
R67189 VSS.n9525 VSS.n710 4.5005
R67190 VSS.n9525 VSS.n9524 4.5005
R67191 VSS.n9525 VSS.n685 4.5005
R67192 VSS.n9526 VSS.n9525 4.5005
R67193 VSS.n9849 VSS.n109 4.5005
R67194 VSS.n9847 VSS.n109 4.5005
R67195 VSS.n113 VSS.n109 4.5005
R67196 VSS.n9849 VSS.n100 4.5005
R67197 VSS.n9847 VSS.n100 4.5005
R67198 VSS.n113 VSS.n100 4.5005
R67199 VSS.n9848 VSS.n113 4.5005
R67200 VSS.n9848 VSS.n116 4.5005
R67201 VSS.n9849 VSS.n9848 4.5005
R67202 VSS.n9848 VSS.n9847 4.5005
R67203 VSS.n153 VSS.n110 4.5005
R67204 VSS.n151 VSS.n110 4.5005
R67205 VSS.n149 VSS.n110 4.5005
R67206 VSS.n166 VSS.n110 4.5005
R67207 VSS.n2334 VSS.n2330 4.5005
R67208 VSS.n2369 VSS.n2334 4.5005
R67209 VSS.n2369 VSS.n2368 4.5005
R67210 VSS.n2369 VSS.n2333 4.5005
R67211 VSS.n2330 VSS.n1866 4.5005
R67212 VSS.n2369 VSS.n1866 4.5005
R67213 VSS.n2364 VSS.n2341 4.5005
R67214 VSS.n2359 VSS.n2348 4.5005
R67215 VSS.n2356 VSS.n2349 4.5005
R67216 VSS.n2349 VSS.n762 4.5005
R67217 VSS.n9451 VSS.n763 4.5005
R67218 VSS.n9449 VSS.n763 4.5005
R67219 VSS.n9444 VSS.n776 4.5005
R67220 VSS.n9439 VSS.n9373 4.5005
R67221 VSS.n2363 VSS.n2338 4.5005
R67222 VSS.n2364 VSS.n2363 4.5005
R67223 VSS.n2358 VSS.n2345 4.5005
R67224 VSS.n2359 VSS.n2358 4.5005
R67225 VSS.n2354 VSS.n762 4.5005
R67226 VSS.n9449 VSS.n9448 4.5005
R67227 VSS.n9443 VSS.n773 4.5005
R67228 VSS.n9444 VSS.n9443 4.5005
R67229 VSS.n9438 VSS.n9370 4.5005
R67230 VSS.n9439 VSS.n9438 4.5005
R67231 VSS.n2340 VSS.n2338 4.5005
R67232 VSS.n2364 VSS.n2340 4.5005
R67233 VSS.n2347 VSS.n2345 4.5005
R67234 VSS.n2359 VSS.n2347 4.5005
R67235 VSS.n2352 VSS.n762 4.5005
R67236 VSS.n9449 VSS.n768 4.5005
R67237 VSS.n775 VSS.n773 4.5005
R67238 VSS.n9444 VSS.n775 4.5005
R67239 VSS.n9372 VSS.n9370 4.5005
R67240 VSS.n9439 VSS.n9372 4.5005
R67241 VSS.n2366 VSS.n2365 4.5005
R67242 VSS.n2365 VSS.n2338 4.5005
R67243 VSS.n2365 VSS.n2364 4.5005
R67244 VSS.n2361 VSS.n2360 4.5005
R67245 VSS.n2360 VSS.n2345 4.5005
R67246 VSS.n2360 VSS.n2359 4.5005
R67247 VSS.n2356 VSS.n915 4.5005
R67248 VSS.n915 VSS.n762 4.5005
R67249 VSS.n9451 VSS.n9450 4.5005
R67250 VSS.n9450 VSS.n9449 4.5005
R67251 VSS.n9446 VSS.n9445 4.5005
R67252 VSS.n9445 VSS.n773 4.5005
R67253 VSS.n9445 VSS.n9444 4.5005
R67254 VSS.n9441 VSS.n9440 4.5005
R67255 VSS.n9440 VSS.n9370 4.5005
R67256 VSS.n9440 VSS.n9439 4.5005
R67257 VSS.n9436 VSS.n9374 4.5005
R67258 VSS.n9433 VSS.n9374 4.5005
R67259 VSS.n9434 VSS.n9433 4.5005
R67260 VSS.n9433 VSS.n9377 4.5005
R67261 VSS.n9436 VSS.n711 4.5005
R67262 VSS.n9433 VSS.n711 4.5005
R67263 VSS.n2271 VSS.n2170 4.5005
R67264 VSS.n2275 VSS.n2271 4.5005
R67265 VSS.n2275 VSS.n2274 4.5005
R67266 VSS.n2276 VSS.n2170 4.5005
R67267 VSS.n2277 VSS.n2276 4.5005
R67268 VSS.n2276 VSS.n2275 4.5005
R67269 VSS.n8096 VSS.n8095 4.5005
R67270 VSS.n2439 VSS.n2430 4.5005
R67271 VSS.n2440 VSS.n2428 4.5005
R67272 VSS.n2445 VSS.n2428 4.5005
R67273 VSS.n2465 VSS.n2446 4.5005
R67274 VSS.n2462 VSS.n2446 4.5005
R67275 VSS.n2458 VSS.n2454 4.5005
R67276 VSS.n8970 VSS.n8969 4.5005
R67277 VSS.n8091 VSS.n2085 4.5005
R67278 VSS.n8095 VSS.n2085 4.5005
R67279 VSS.n2434 VSS.n2432 4.5005
R67280 VSS.n2439 VSS.n2432 4.5005
R67281 VSS.n2445 VSS.n2444 4.5005
R67282 VSS.n2463 VSS.n2462 4.5005
R67283 VSS.n2459 VSS.n2453 4.5005
R67284 VSS.n2459 VSS.n2458 4.5005
R67285 VSS.n8965 VSS.n1095 4.5005
R67286 VSS.n8969 VSS.n1095 4.5005
R67287 VSS.n8095 VSS.n2083 4.5005
R67288 VSS.n2439 VSS.n1542 4.5005
R67289 VSS.n2458 VSS.n1429 4.5005
R67290 VSS.n8969 VSS.n1093 4.5005
R67291 VSS.n8090 VSS.n2088 4.5005
R67292 VSS.n8091 VSS.n8090 4.5005
R67293 VSS.n2084 VSS.n1540 4.5005
R67294 VSS.n2434 VSS.n1540 4.5005
R67295 VSS.n2445 VSS.n1493 4.5005
R67296 VSS.n2462 VSS.n1460 4.5005
R67297 VSS.n2461 VSS.n1428 4.5005
R67298 VSS.n2453 VSS.n1428 4.5005
R67299 VSS.n8964 VSS.n1098 4.5005
R67300 VSS.n8965 VSS.n8964 4.5005
R67301 VSS.n1220 VSS.n1094 4.5005
R67302 VSS.n1223 VSS.n1220 4.5005
R67303 VSS.n1223 VSS.n1222 4.5005
R67304 VSS.n1224 VSS.n1167 4.5005
R67305 VSS.n1224 VSS.n1223 4.5005
R67306 VSS.n1223 VSS.n1164 4.5005
R67307 VSS.n2795 VSS.n2794 4.38021
R67308 VSS.n4636 VSS.n3855 4.38021
R67309 VSS.n9816 VSS.n9815 4.38021
R67310 VSS.n9571 VSS.n533 4.38021
R67311 VSS.n9815 VSS.n167 4.36815
R67312 VSS.n6254 VSS.n3855 4.36815
R67313 VSS.n6255 VSS.n6254 4.36815
R67314 VSS.n4154 VSS.n167 4.36815
R67315 VSS.n4154 VSS.n434 4.36815
R67316 VSS.n6255 VSS.n3830 4.36815
R67317 VSS.n491 VSS.n443 4.36815
R67318 VSS.n3827 VSS.n3230 4.36815
R67319 VSS.n5772 VSS.n3230 4.36815
R67320 VSS.n500 VSS.n491 4.36815
R67321 VSS.n533 VSS.n500 4.36815
R67322 VSS.n5772 VSS.n2795 4.36815
R67323 VSS.n7141 VSS.n2469 2.2505
R67324 VSS.n7144 VSS.n7143 2.2505
R67325 VSS.n7145 VSS.n7144 2.2505
R67326 VSS.n7269 VSS.n2470 2.2505
R67327 VSS.n7269 VSS.n7268 2.2505
R67328 VSS.n4758 VSS.n4757 2.24726
R67329 VSS.n4745 VSS.n4744 2.24726
R67330 VSS.n176 VSS.n169 2.24726
R67331 VSS.n9811 VSS.n168 2.24726
R67332 VSS.n6250 VSS.n3858 2.24726
R67333 VSS.n3863 VSS.n3857 2.24726
R67334 VSS.n5470 VSS.n5469 2.24726
R67335 VSS.n5468 VSS.n5467 2.24726
R67336 VSS.n6258 VSS.n3852 2.24726
R67337 VSS.n6257 VSS.n6256 2.24726
R67338 VSS.n4153 VSS.n4148 2.24726
R67339 VSS.n4152 VSS.n4149 2.24726
R67340 VSS.n431 VSS.n429 2.24726
R67341 VSS.n6266 VSS.n6265 2.24726
R67342 VSS.n433 VSS.n432 2.24726
R67343 VSS.n440 VSS.n438 2.24726
R67344 VSS.n6275 VSS.n3825 2.24726
R67345 VSS.n442 VSS.n441 2.24726
R67346 VSS.n488 VSS.n486 2.24726
R67347 VSS.n6574 VSS.n3227 2.24726
R67348 VSS.n490 VSS.n489 2.24726
R67349 VSS.n497 VSS.n495 2.24726
R67350 VSS.n5770 VSS.n3229 2.24726
R67351 VSS.n499 VSS.n498 2.24726
R67352 VSS.n530 VSS.n528 2.24726
R67353 VSS.n6966 VSS.n2771 2.24726
R67354 VSS.n532 VSS.n531 2.24726
R67355 VSS.n4750 VSS.n4571 2.2467
R67356 VSS.n5252 VSS.n4321 2.2467
R67357 VSS.n5075 VSS.n4515 2.2467
R67358 VSS.n5082 VSS.n4506 2.2467
R67359 VSS.n4974 VSS.n4873 2.2467
R67360 VSS.n9688 VSS.n277 2.2467
R67361 VSS.n9762 VSS.n219 2.2467
R67362 VSS.n4747 VSS.n4561 2.2467
R67363 VSS.n4752 VSS.n4561 2.2467
R67364 VSS.n5248 VSS.n5247 2.2467
R67365 VSS.n5247 VSS.n4324 2.2467
R67366 VSS.n5074 VSS.n5073 2.2467
R67367 VSS.n5073 VSS.n4514 2.2467
R67368 VSS.n4509 VSS.n4505 2.2467
R67369 VSS.n4968 VSS.n4870 2.2467
R67370 VSS.n274 VSS.n273 2.2467
R67371 VSS.n275 VSS.n274 2.2467
R67372 VSS.n9761 VSS.n9760 2.2467
R67373 VSS.n9760 VSS.n218 2.2467
R67374 VSS.n4566 VSS.n3890 2.2467
R67375 VSS.n5263 VSS.n4318 2.2467
R67376 VSS.n5645 VSS.n4282 2.2467
R67377 VSS.n5653 VSS.n4274 2.2467
R67378 VSS.n4918 VSS.n4917 2.2467
R67379 VSS.n285 VSS.n284 2.2467
R67380 VSS.n5454 VSS.n5448 2.2467
R67381 VSS.n5259 VSS.n5258 2.2467
R67382 VSS.n5258 VSS.n5254 2.2467
R67383 VSS.n5644 VSS.n5643 2.2467
R67384 VSS.n5643 VSS.n4281 2.2467
R67385 VSS.n5649 VSS.n4276 2.2467
R67386 VSS.n4916 VSS.n4915 2.2467
R67387 VSS.n297 VSS.n296 2.2467
R67388 VSS.n297 VSS.n282 2.2467
R67389 VSS.n5453 VSS.n5452 2.2467
R67390 VSS.n5452 VSS.n5447 2.2467
R67391 VSS.n4090 VSS.n3904 2.2467
R67392 VSS.n4099 VSS.n3950 2.2467
R67393 VSS.n4107 VSS.n3995 2.2467
R67394 VSS.n4112 VSS.n4027 2.2467
R67395 VSS.n5725 VSS.n4118 2.2467
R67396 VSS.n4128 VSS.n324 2.2467
R67397 VSS.n4136 VSS.n357 2.2467
R67398 VSS.n4098 VSS.n4097 2.2467
R67399 VSS.n4097 VSS.n4085 2.2467
R67400 VSS.n4106 VSS.n4105 2.2467
R67401 VSS.n4105 VSS.n4081 2.2467
R67402 VSS.n4111 VSS.n4077 2.2467
R67403 VSS.n4123 VSS.n4117 2.2467
R67404 VSS.n4130 VSS.n4125 2.2467
R67405 VSS.n4131 VSS.n4130 2.2467
R67406 VSS.n4138 VSS.n4133 2.2467
R67407 VSS.n4139 VSS.n4138 2.2467
R67408 VSS.n6065 VSS.n6049 2.2467
R67409 VSS.n6072 VSS.n6041 2.2467
R67410 VSS.n5947 VSS.n5911 2.2467
R67411 VSS.n5939 VSS.n5918 2.2467
R67412 VSS.n6054 VSS.n3905 2.2467
R67413 VSS.n6053 VSS.n3952 2.2467
R67414 VSS.n6045 VSS.n3996 2.2467
R67415 VSS.n6081 VSS.n4069 2.2467
R67416 VSS.n5907 VSS.n5906 2.2467
R67417 VSS.n5914 VSS.n325 2.2467
R67418 VSS.n5921 VSS.n359 2.2467
R67419 VSS.n6291 VSS.n3813 2.2467
R67420 VSS.n6298 VSS.n3804 2.2467
R67421 VSS.n6320 VSS.n3700 2.2467
R67422 VSS.n6327 VSS.n3691 2.2467
R67423 VSS.n3821 VSS.n3818 2.2467
R67424 VSS.n3817 VSS.n3810 2.2467
R67425 VSS.n3808 VSS.n3801 2.2467
R67426 VSS.n6307 VSS.n3715 2.2467
R67427 VSS.n6312 VSS.n6311 2.2467
R67428 VSS.n3704 VSS.n3697 2.2467
R67429 VSS.n3695 VSS.n3688 2.2467
R67430 VSS.n6585 VSS.n3219 2.2467
R67431 VSS.n6591 VSS.n3210 2.2467
R67432 VSS.n6598 VSS.n3201 2.2467
R67433 VSS.n6626 VSS.n2966 2.2467
R67434 VSS.n6639 VSS.n3114 2.2467
R67435 VSS.n3223 VSS.n3216 2.2467
R67436 VSS.n3214 VSS.n3207 2.2467
R67437 VSS.n3205 VSS.n3198 2.2467
R67438 VSS.n6607 VSS.n3190 2.2467
R67439 VSS.n6618 VSS.n6617 2.2467
R67440 VSS.n3126 VSS.n3120 2.2467
R67441 VSS.n6635 VSS.n3116 2.2467
R67442 VSS.n5783 VSS.n5762 2.2467
R67443 VSS.n5789 VSS.n5753 2.2467
R67444 VSS.n5796 VSS.n5744 2.2467
R67445 VSS.n6753 VSS.n2964 2.2467
R67446 VSS.n6650 VSS.n6643 2.2467
R67447 VSS.n5766 VSS.n5759 2.2467
R67448 VSS.n5757 VSS.n5750 2.2467
R67449 VSS.n5748 VSS.n5741 2.2467
R67450 VSS.n5886 VSS.n5885 2.2467
R67451 VSS.n5879 VSS.n5878 2.2467
R67452 VSS.n6758 VSS.n2967 2.2467
R67453 VSS.n6647 VSS.n6640 2.2467
R67454 VSS.n6977 VSS.n2763 2.2467
R67455 VSS.n6983 VSS.n2754 2.2467
R67456 VSS.n6990 VSS.n2745 2.2467
R67457 VSS.n7012 VSS.n2638 2.2467
R67458 VSS.n7019 VSS.n2629 2.2467
R67459 VSS.n2767 VSS.n2760 2.2467
R67460 VSS.n2758 VSS.n2751 2.2467
R67461 VSS.n2749 VSS.n2742 2.2467
R67462 VSS.n6999 VSS.n2653 2.2467
R67463 VSS.n7004 VSS.n7003 2.2467
R67464 VSS.n2642 VSS.n2635 2.2467
R67465 VSS.n2633 VSS.n2626 2.2467
R67466 VSS.n7031 VSS.n2620 2.2467
R67467 VSS.n6662 VSS.n3107 2.2467
R67468 VSS.n3664 VSS.n3659 2.2467
R67469 VSS.n6339 VSS.n3682 2.2467
R67470 VSS.n5932 VSS.n5925 2.2467
R67471 VSS.n4144 VSS.n396 2.2467
R67472 VSS.n4146 VSS.n4141 2.2467
R67473 VSS.n4147 VSS.n4146 2.2467
R67474 VSS.n5461 VSS.n5443 2.2467
R67475 VSS.n5460 VSS.n5459 2.2467
R67476 VSS.n5459 VSS.n5442 2.2467
R67477 VSS.n9768 VSS.n205 2.2467
R67478 VSS.n9767 VSS.n202 2.2467
R67479 VSS.n9770 VSS.n202 2.2467
R67480 VSS.n5928 VSS.n397 2.2467
R67481 VSS.n6335 VSS.n3684 2.2467
R67482 VSS.n3668 VSS.n3654 2.2467
R67483 VSS.n6658 VSS.n3109 2.2467
R67484 VSS.n7027 VSS.n2622 2.2467
R67485 VSS.n7152 VSS.n7151 2.24623
R67486 VSS.n2567 VSS.n2564 2.24623
R67487 VSS.n7100 VSS.n7058 2.24623
R67488 VSS.n2529 VSS.n2527 2.24623
R67489 VSS.n7219 VSS.n2531 2.24623
R67490 VSS.n7090 VSS.n7087 2.24623
R67491 VSS.n7092 VSS.n7059 2.24623
R67492 VSS.n7163 VSS.n2551 2.24623
R67493 VSS.n7164 VSS.n2549 2.24623
R67494 VSS.n7157 VSS.n2552 2.24623
R67495 VSS.n2481 VSS.n2479 2.24623
R67496 VSS.n7236 VSS.n2510 2.24623
R67497 VSS.n7187 VSS.n7186 2.24623
R67498 VSS.n2486 VSS.n2483 2.24623
R67499 VSS.n2490 VSS.n2489 2.24623
R67500 VSS.n7194 VSS.n7189 2.24623
R67501 VSS.n7238 VSS.n2507 2.24623
R67502 VSS.n7244 VSS.n2504 2.24623
R67503 VSS.n8556 VSS.n8555 2.24623
R67504 VSS.n8835 VSS.n8834 2.24623
R67505 VSS.n1346 VSS.n1343 2.24623
R67506 VSS.n1603 VSS.n1601 2.24623
R67507 VSS.n8833 VSS.n1351 2.24623
R67508 VSS.n1391 VSS.n1390 2.24623
R67509 VSS.n1600 VSS.n1598 2.24623
R67510 VSS.n1593 VSS.n1592 2.24623
R67511 VSS.n8041 VSS.n8039 2.24623
R67512 VSS.n8032 VSS.n8031 2.24623
R67513 VSS.n8017 VSS.n8016 2.24623
R67514 VSS.n8010 VSS.n8009 2.24623
R67515 VSS.n8852 VSS.n1310 2.24623
R67516 VSS.n8845 VSS.n1316 2.24623
R67517 VSS.n8389 VSS.n8388 2.24623
R67518 VSS.n1566 VSS.n1561 2.24623
R67519 VSS.n7049 VSS.n2605 2.24623
R67520 VSS.n7103 VSS.n2603 2.24623
R67521 VSS.n7118 VSS.n2592 2.24623
R67522 VSS.n2590 VSS.n2587 2.24623
R67523 VSS.n7135 VSS.n2577 2.24623
R67524 VSS.n7134 VSS.n2578 2.24623
R67525 VSS.n2785 VSS.n2784 2.24623
R67526 VSS.n2586 VSS.n2581 2.24623
R67527 VSS.n2585 VSS.n2582 2.24623
R67528 VSS.n2781 VSS.n2779 2.24623
R67529 VSS.n2794 VSS.n2793 2.24623
R67530 VSS.n9605 VSS.n430 2.24623
R67531 VSS.n6273 VSS.n6272 2.24623
R67532 VSS.n6270 VSS.n6267 2.24623
R67533 VSS.n6273 VSS.n3831 2.24623
R67534 VSS.n9603 VSS.n427 2.24623
R67535 VSS.n6267 VSS.n3828 2.24623
R67536 VSS.n9600 VSS.n439 2.24623
R67537 VSS.n6280 VSS.n6279 2.24623
R67538 VSS.n6278 VSS.n6277 2.24623
R67539 VSS.n6280 VSS.n6276 2.24623
R67540 VSS.n9598 VSS.n436 2.24623
R67541 VSS.n6278 VSS.n3826 2.24623
R67542 VSS.n9592 VSS.n487 2.24623
R67543 VSS.n6579 VSS.n6578 2.24623
R67544 VSS.n6577 VSS.n6576 2.24623
R67545 VSS.n6579 VSS.n6575 2.24623
R67546 VSS.n9590 VSS.n484 2.24623
R67547 VSS.n6577 VSS.n3228 2.24623
R67548 VSS.n9587 VSS.n496 2.24623
R67549 VSS.n5777 VSS.n5776 2.24623
R67550 VSS.n5775 VSS.n5774 2.24623
R67551 VSS.n5777 VSS.n5773 2.24623
R67552 VSS.n9585 VSS.n493 2.24623
R67553 VSS.n5775 VSS.n5771 2.24623
R67554 VSS.n9579 VSS.n529 2.24623
R67555 VSS.n6971 VSS.n6970 2.24623
R67556 VSS.n6969 VSS.n6968 2.24623
R67557 VSS.n6971 VSS.n6967 2.24623
R67558 VSS.n9577 VSS.n526 2.24623
R67559 VSS.n6969 VSS.n2772 2.24623
R67560 VSS.n2616 VSS.n2615 2.24623
R67561 VSS.n9571 VSS.n535 2.24623
R67562 VSS.n2613 VSS.n2609 2.24623
R67563 VSS.n7043 VSS.n7042 2.24623
R67564 VSS.n7036 VSS.n7033 2.24623
R67565 VSS.n2370 VSS.n2332 2.24623
R67566 VSS.n2367 VSS.n2330 2.24623
R67567 VSS.n2370 VSS.n2331 2.24623
R67568 VSS.n9378 VSS.n9375 2.24623
R67569 VSS.n9436 VSS.n9435 2.24623
R67570 VSS.n9376 VSS.n9375 2.24623
R67571 VSS.n2277 VSS.n2171 2.24623
R67572 VSS.n2273 VSS.n2170 2.24623
R67573 VSS.n1221 VSS.n1167 2.24623
R67574 VSS.n1168 VSS.n1094 2.24623
R67575 VSS.n2272 VSS.n2172 2.24582
R67576 VSS.n1166 VSS.n1164 2.24582
R67577 VSS.n5527 VSS.n5382 2.24552
R67578 VSS.n5522 VSS.n5395 2.24552
R67579 VSS.n5527 VSS.n5381 2.24552
R67580 VSS.n5523 VSS.n5522 2.24552
R67581 VSS.n5527 VSS.n5380 2.24552
R67582 VSS.n5522 VSS.n5388 2.24552
R67583 VSS.n9644 VSS.n366 2.24552
R67584 VSS.n362 VSS.n360 2.24552
R67585 VSS.n9644 VSS.n365 2.24552
R67586 VSS.n362 VSS.n361 2.24552
R67587 VSS.n9644 VSS.n364 2.24552
R67588 VSS.n3075 VSS.n3074 2.24552
R67589 VSS.n3081 VSS.n3080 2.24552
R67590 VSS.n3075 VSS.n3073 2.24552
R67591 VSS.n3081 VSS.n3079 2.24552
R67592 VSS.n3075 VSS.n3072 2.24552
R67593 VSS.n3081 VSS.n3078 2.24552
R67594 VSS.n3075 VSS.n3071 2.24552
R67595 VSS.n3081 VSS.n3077 2.24552
R67596 VSS.n3075 VSS.n3070 2.24552
R67597 VSS.n3081 VSS.n3069 2.24552
R67598 VSS.n1295 VSS.n1288 2.24552
R67599 VSS.n1297 VSS.n1284 2.24552
R67600 VSS.n1298 VSS.n1288 2.24552
R67601 VSS.n1300 VSS.n1284 2.24552
R67602 VSS.n8861 VSS.n1290 2.24552
R67603 VSS.n1307 VSS.n1284 2.24552
R67604 VSS.n1302 VSS.n1288 2.24552
R67605 VSS.n1304 VSS.n1284 2.24552
R67606 VSS.n8962 VSS.n1138 2.24552
R67607 VSS.n8962 VSS.n1136 2.24552
R67608 VSS.n1134 VSS.n1101 2.24552
R67609 VSS.n8962 VSS.n1132 2.24552
R67610 VSS.n1130 VSS.n1101 2.24552
R67611 VSS.n8962 VSS.n1128 2.24552
R67612 VSS.n1126 VSS.n1101 2.24552
R67613 VSS.n8962 VSS.n1124 2.24552
R67614 VSS.n1122 VSS.n1101 2.24552
R67615 VSS.n8962 VSS.n1120 2.24552
R67616 VSS.n1117 VSS.n1101 2.24552
R67617 VSS.n8962 VSS.n1115 2.24552
R67618 VSS.n1113 VSS.n1101 2.24552
R67619 VSS.n8962 VSS.n1111 2.24552
R67620 VSS.n1109 VSS.n1101 2.24552
R67621 VSS.n8962 VSS.n1107 2.24552
R67622 VSS.n1105 VSS.n1101 2.24552
R67623 VSS.n8962 VSS.n1103 2.24552
R67624 VSS.n9014 VSS.n8986 2.24552
R67625 VSS.n9016 VSS.n1090 2.24552
R67626 VSS.n9011 VSS.n9002 2.24552
R67627 VSS.n9016 VSS.n1089 2.24552
R67628 VSS.n9011 VSS.n9003 2.24552
R67629 VSS.n9016 VSS.n1088 2.24552
R67630 VSS.n9011 VSS.n9004 2.24552
R67631 VSS.n9016 VSS.n1087 2.24552
R67632 VSS.n9011 VSS.n9005 2.24552
R67633 VSS.n9016 VSS.n1086 2.24552
R67634 VSS.n9011 VSS.n9006 2.24552
R67635 VSS.n9016 VSS.n1085 2.24552
R67636 VSS.n9011 VSS.n9007 2.24552
R67637 VSS.n9016 VSS.n1084 2.24552
R67638 VSS.n9011 VSS.n9008 2.24552
R67639 VSS.n9016 VSS.n1083 2.24552
R67640 VSS.n9011 VSS.n9009 2.24552
R67641 VSS.n9016 VSS.n1082 2.24552
R67642 VSS.n9011 VSS.n9010 2.24552
R67643 VSS.n9016 VSS.n1081 2.24552
R67644 VSS.n9012 VSS.n9011 2.24552
R67645 VSS.n9016 VSS.n1080 2.24552
R67646 VSS.n9011 VSS.n8973 2.24552
R67647 VSS.n9363 VSS.n9353 2.24552
R67648 VSS.n796 VSS.n780 2.24552
R67649 VSS.n9363 VSS.n9354 2.24552
R67650 VSS.n798 VSS.n780 2.24552
R67651 VSS.n9363 VSS.n9355 2.24552
R67652 VSS.n800 VSS.n780 2.24552
R67653 VSS.n9363 VSS.n9356 2.24552
R67654 VSS.n802 VSS.n780 2.24552
R67655 VSS.n9363 VSS.n9357 2.24552
R67656 VSS.n804 VSS.n780 2.24552
R67657 VSS.n9363 VSS.n9358 2.24552
R67658 VSS.n806 VSS.n780 2.24552
R67659 VSS.n9363 VSS.n9359 2.24552
R67660 VSS.n808 VSS.n780 2.24552
R67661 VSS.n9363 VSS.n9360 2.24552
R67662 VSS.n810 VSS.n780 2.24552
R67663 VSS.n9363 VSS.n9361 2.24552
R67664 VSS.n812 VSS.n780 2.24552
R67665 VSS.n9363 VSS.n9362 2.24552
R67666 VSS.n814 VSS.n780 2.24552
R67667 VSS.n9364 VSS.n9363 2.24552
R67668 VSS.n9365 VSS.n780 2.24552
R67669 VSS.n9363 VSS.n779 2.24552
R67670 VSS.n6428 VSS.n3600 2.24552
R67671 VSS.n3626 VSS.n3622 2.24552
R67672 VSS.n6424 VSS.n6414 2.24552
R67673 VSS.n3622 VSS.n3621 2.24552
R67674 VSS.n6424 VSS.n6415 2.24552
R67675 VSS.n3622 VSS.n3620 2.24552
R67676 VSS.n6424 VSS.n6416 2.24552
R67677 VSS.n3622 VSS.n3619 2.24552
R67678 VSS.n6424 VSS.n6417 2.24552
R67679 VSS.n3622 VSS.n3618 2.24552
R67680 VSS.n6424 VSS.n6418 2.24552
R67681 VSS.n3622 VSS.n3617 2.24552
R67682 VSS.n6424 VSS.n6419 2.24552
R67683 VSS.n3622 VSS.n3616 2.24552
R67684 VSS.n6424 VSS.n6420 2.24552
R67685 VSS.n3622 VSS.n3615 2.24552
R67686 VSS.n6424 VSS.n6421 2.24552
R67687 VSS.n3622 VSS.n3614 2.24552
R67688 VSS.n6424 VSS.n6422 2.24552
R67689 VSS.n3622 VSS.n3613 2.24552
R67690 VSS.n6424 VSS.n6423 2.24552
R67691 VSS.n3622 VSS.n3612 2.24552
R67692 VSS.n6424 VSS.n3611 2.24552
R67693 VSS.n3328 VSS.n3327 2.24552
R67694 VSS.n3315 VSS.n3314 2.24552
R67695 VSS.n3328 VSS.n3326 2.24552
R67696 VSS.n3315 VSS.n3313 2.24552
R67697 VSS.n3328 VSS.n3325 2.24552
R67698 VSS.n3315 VSS.n3312 2.24552
R67699 VSS.n3328 VSS.n3324 2.24552
R67700 VSS.n3315 VSS.n3311 2.24552
R67701 VSS.n3328 VSS.n3323 2.24552
R67702 VSS.n3315 VSS.n3310 2.24552
R67703 VSS.n3328 VSS.n3322 2.24552
R67704 VSS.n3315 VSS.n3309 2.24552
R67705 VSS.n3328 VSS.n3321 2.24552
R67706 VSS.n3315 VSS.n3308 2.24552
R67707 VSS.n3328 VSS.n3320 2.24552
R67708 VSS.n3315 VSS.n3307 2.24552
R67709 VSS.n3328 VSS.n3319 2.24552
R67710 VSS.n3315 VSS.n3306 2.24552
R67711 VSS.n3328 VSS.n3318 2.24552
R67712 VSS.n3315 VSS.n3305 2.24552
R67713 VSS.n3328 VSS.n3317 2.24552
R67714 VSS.n3315 VSS.n3304 2.24552
R67715 VSS.n3328 VSS.n3303 2.24552
R67716 VSS.n2837 VSS.n2830 2.24552
R67717 VSS.n6938 VSS.n6934 2.24552
R67718 VSS.n2839 VSS.n2830 2.24552
R67719 VSS.n6938 VSS.n6935 2.24552
R67720 VSS.n2841 VSS.n2830 2.24552
R67721 VSS.n6938 VSS.n6936 2.24552
R67722 VSS.n2843 VSS.n2830 2.24552
R67723 VSS.n6938 VSS.n6937 2.24552
R67724 VSS.n2845 VSS.n2830 2.24552
R67725 VSS.n6939 VSS.n6938 2.24552
R67726 VSS.n8323 VSS.n8321 2.24552
R67727 VSS.n8330 VSS.n1688 2.24552
R67728 VSS.n8323 VSS.n8320 2.24552
R67729 VSS.n8330 VSS.n1689 2.24552
R67730 VSS.n8323 VSS.n8319 2.24552
R67731 VSS.n8330 VSS.n1690 2.24552
R67732 VSS.n8324 VSS.n8323 2.24552
R67733 VSS.n8330 VSS.n1691 2.24552
R67734 VSS.n8323 VSS.n1693 2.24552
R67735 VSS.n8330 VSS.n8329 2.24552
R67736 VSS.n2220 VSS.n2175 2.24552
R67737 VSS.n2269 VSS.n2218 2.24552
R67738 VSS.n2216 VSS.n2175 2.24552
R67739 VSS.n2269 VSS.n2214 2.24552
R67740 VSS.n2212 VSS.n2175 2.24552
R67741 VSS.n2269 VSS.n2210 2.24552
R67742 VSS.n2208 VSS.n2175 2.24552
R67743 VSS.n2269 VSS.n2206 2.24552
R67744 VSS.n2204 VSS.n2175 2.24552
R67745 VSS.n2269 VSS.n2202 2.24552
R67746 VSS.n2200 VSS.n2175 2.24552
R67747 VSS.n2269 VSS.n2198 2.24552
R67748 VSS.n2196 VSS.n2175 2.24552
R67749 VSS.n2269 VSS.n2194 2.24552
R67750 VSS.n2192 VSS.n2175 2.24552
R67751 VSS.n2269 VSS.n2190 2.24552
R67752 VSS.n2188 VSS.n2175 2.24552
R67753 VSS.n2269 VSS.n2186 2.24552
R67754 VSS.n2184 VSS.n2175 2.24552
R67755 VSS.n2269 VSS.n2182 2.24552
R67756 VSS.n2180 VSS.n2175 2.24552
R67757 VSS.n2269 VSS.n2178 2.24552
R67758 VSS.n4784 VSS.n4576 2.24552
R67759 VSS.n4780 VSS.n4563 2.24552
R67760 VSS.n4786 VSS.n4556 2.24552
R67761 VSS.n4782 VSS.n4563 2.24552
R67762 VSS.n4786 VSS.n4555 2.24552
R67763 VSS.n4573 VSS.n4563 2.24552
R67764 VSS.n9748 VSS.n226 2.24552
R67765 VSS.n9750 VSS.n227 2.24552
R67766 VSS.n9751 VSS.n226 2.24552
R67767 VSS.n9753 VSS.n227 2.24552
R67768 VSS.n9754 VSS.n226 2.24552
R67769 VSS.n9756 VSS.n227 2.24552
R67770 VSS.n269 VSS.n258 2.24552
R67771 VSS.n9696 VSS.n257 2.24552
R67772 VSS.n269 VSS.n267 2.24552
R67773 VSS.n9696 VSS.n256 2.24552
R67774 VSS.n269 VSS.n266 2.24552
R67775 VSS.n9696 VSS.n255 2.24552
R67776 VSS.n299 VSS.n287 2.24552
R67777 VSS.n301 VSS.n288 2.24552
R67778 VSS.n302 VSS.n287 2.24552
R67779 VSS.n304 VSS.n288 2.24552
R67780 VSS.n305 VSS.n287 2.24552
R67781 VSS.n307 VSS.n288 2.24552
R67782 VSS.n9678 VSS.n308 2.24552
R67783 VSS.n318 VSS.n309 2.24552
R67784 VSS.n9678 VSS.n327 2.24552
R67785 VSS.n320 VSS.n309 2.24552
R67786 VSS.n9678 VSS.n326 2.24552
R67787 VSS.n3562 VSS.n3551 2.24552
R67788 VSS.n3550 VSS.n3549 2.24552
R67789 VSS.n3562 VSS.n3552 2.24552
R67790 VSS.n3550 VSS.n3548 2.24552
R67791 VSS.n3562 VSS.n3553 2.24552
R67792 VSS.n3550 VSS.n3547 2.24552
R67793 VSS.n3562 VSS.n3554 2.24552
R67794 VSS.n3550 VSS.n3546 2.24552
R67795 VSS.n3562 VSS.n3555 2.24552
R67796 VSS.n3550 VSS.n3545 2.24552
R67797 VSS.n3562 VSS.n3556 2.24552
R67798 VSS.n3550 VSS.n3544 2.24552
R67799 VSS.n3562 VSS.n3557 2.24552
R67800 VSS.n3550 VSS.n3543 2.24552
R67801 VSS.n3562 VSS.n3558 2.24552
R67802 VSS.n3550 VSS.n3542 2.24552
R67803 VSS.n3562 VSS.n3559 2.24552
R67804 VSS.n3550 VSS.n3541 2.24552
R67805 VSS.n3562 VSS.n3560 2.24552
R67806 VSS.n3550 VSS.n3540 2.24552
R67807 VSS.n3562 VSS.n3561 2.24552
R67808 VSS.n3550 VSS.n3539 2.24552
R67809 VSS.n3562 VSS.n3538 2.24552
R67810 VSS.n6749 VSS.n2972 2.24552
R67811 VSS.n2982 VSS.n2973 2.24552
R67812 VSS.n6749 VSS.n2994 2.24552
R67813 VSS.n2984 VSS.n2973 2.24552
R67814 VSS.n6749 VSS.n2993 2.24552
R67815 VSS.n2986 VSS.n2973 2.24552
R67816 VSS.n6749 VSS.n2992 2.24552
R67817 VSS.n2988 VSS.n2973 2.24552
R67818 VSS.n6749 VSS.n2991 2.24552
R67819 VSS.n2990 VSS.n2973 2.24552
R67820 VSS.n1332 VSS.n1322 2.24552
R67821 VSS.n1334 VSS.n1323 2.24552
R67822 VSS.n1335 VSS.n1322 2.24552
R67823 VSS.n1337 VSS.n1323 2.24552
R67824 VSS.n1327 VSS.n1324 2.24552
R67825 VSS.n1339 VSS.n1322 2.24552
R67826 VSS.n1340 VSS.n1323 2.24552
R67827 VSS.n1342 VSS.n1322 2.24552
R67828 VSS.n8803 VSS.n1392 2.24552
R67829 VSS.n1409 VSS.n1394 2.24552
R67830 VSS.n8803 VSS.n8795 2.24552
R67831 VSS.n1411 VSS.n1393 2.24552
R67832 VSS.n8803 VSS.n8796 2.24552
R67833 VSS.n1413 VSS.n1393 2.24552
R67834 VSS.n8803 VSS.n8797 2.24552
R67835 VSS.n1415 VSS.n1393 2.24552
R67836 VSS.n8803 VSS.n8798 2.24552
R67837 VSS.n1417 VSS.n1393 2.24552
R67838 VSS.n8803 VSS.n8799 2.24552
R67839 VSS.n1420 VSS.n1393 2.24552
R67840 VSS.n8803 VSS.n8800 2.24552
R67841 VSS.n1422 VSS.n1393 2.24552
R67842 VSS.n8803 VSS.n8801 2.24552
R67843 VSS.n1424 VSS.n1393 2.24552
R67844 VSS.n8803 VSS.n8802 2.24552
R67845 VSS.n1426 VSS.n1393 2.24552
R67846 VSS.n9053 VSS.n1045 2.24552
R67847 VSS.n9055 VSS.n1031 2.24552
R67848 VSS.n9050 VSS.n9040 2.24552
R67849 VSS.n9055 VSS.n1030 2.24552
R67850 VSS.n9050 VSS.n9041 2.24552
R67851 VSS.n9055 VSS.n1029 2.24552
R67852 VSS.n9050 VSS.n9042 2.24552
R67853 VSS.n9055 VSS.n1028 2.24552
R67854 VSS.n9050 VSS.n9043 2.24552
R67855 VSS.n9055 VSS.n1027 2.24552
R67856 VSS.n9050 VSS.n9044 2.24552
R67857 VSS.n9055 VSS.n1026 2.24552
R67858 VSS.n9050 VSS.n9045 2.24552
R67859 VSS.n9055 VSS.n1025 2.24552
R67860 VSS.n9050 VSS.n9046 2.24552
R67861 VSS.n9055 VSS.n1024 2.24552
R67862 VSS.n9050 VSS.n9047 2.24552
R67863 VSS.n9055 VSS.n1023 2.24552
R67864 VSS.n9050 VSS.n9048 2.24552
R67865 VSS.n9055 VSS.n1022 2.24552
R67866 VSS.n9051 VSS.n9050 2.24552
R67867 VSS.n9055 VSS.n1021 2.24552
R67868 VSS.n9050 VSS.n9049 2.24552
R67869 VSS.n9309 VSS.n844 2.24552
R67870 VSS.n9314 VSS.n842 2.24552
R67871 VSS.n9309 VSS.n9299 2.24552
R67872 VSS.n9314 VSS.n841 2.24552
R67873 VSS.n9309 VSS.n9300 2.24552
R67874 VSS.n9314 VSS.n840 2.24552
R67875 VSS.n9309 VSS.n9301 2.24552
R67876 VSS.n9314 VSS.n839 2.24552
R67877 VSS.n9309 VSS.n9302 2.24552
R67878 VSS.n9314 VSS.n838 2.24552
R67879 VSS.n9309 VSS.n9303 2.24552
R67880 VSS.n9314 VSS.n837 2.24552
R67881 VSS.n9309 VSS.n9304 2.24552
R67882 VSS.n9314 VSS.n836 2.24552
R67883 VSS.n9309 VSS.n9305 2.24552
R67884 VSS.n9314 VSS.n835 2.24552
R67885 VSS.n9309 VSS.n9306 2.24552
R67886 VSS.n9314 VSS.n834 2.24552
R67887 VSS.n9309 VSS.n9307 2.24552
R67888 VSS.n9314 VSS.n833 2.24552
R67889 VSS.n9310 VSS.n9309 2.24552
R67890 VSS.n9314 VSS.n832 2.24552
R67891 VSS.n9309 VSS.n9308 2.24552
R67892 VSS.n5061 VSS.n4522 2.24552
R67893 VSS.n5063 VSS.n4523 2.24552
R67894 VSS.n5064 VSS.n4522 2.24552
R67895 VSS.n5066 VSS.n4523 2.24552
R67896 VSS.n5067 VSS.n4522 2.24552
R67897 VSS.n5069 VSS.n4523 2.24552
R67898 VSS.n5631 VSS.n4289 2.24552
R67899 VSS.n5633 VSS.n4290 2.24552
R67900 VSS.n5634 VSS.n4289 2.24552
R67901 VSS.n5636 VSS.n4290 2.24552
R67902 VSS.n5637 VSS.n4289 2.24552
R67903 VSS.n5639 VSS.n4290 2.24552
R67904 VSS.n3987 VSS.n3980 2.24552
R67905 VSS.n6159 VSS.n6157 2.24552
R67906 VSS.n3989 VSS.n3980 2.24552
R67907 VSS.n6159 VSS.n6158 2.24552
R67908 VSS.n3991 VSS.n3980 2.24552
R67909 VSS.n3463 VSS.n3452 2.24552
R67910 VSS.n3451 VSS.n3450 2.24552
R67911 VSS.n3463 VSS.n3453 2.24552
R67912 VSS.n3451 VSS.n3449 2.24552
R67913 VSS.n3463 VSS.n3454 2.24552
R67914 VSS.n3451 VSS.n3448 2.24552
R67915 VSS.n3463 VSS.n3455 2.24552
R67916 VSS.n3451 VSS.n3447 2.24552
R67917 VSS.n3463 VSS.n3456 2.24552
R67918 VSS.n3451 VSS.n3446 2.24552
R67919 VSS.n3463 VSS.n3457 2.24552
R67920 VSS.n3451 VSS.n3445 2.24552
R67921 VSS.n3463 VSS.n3458 2.24552
R67922 VSS.n3451 VSS.n3444 2.24552
R67923 VSS.n3463 VSS.n3459 2.24552
R67924 VSS.n3451 VSS.n3443 2.24552
R67925 VSS.n3463 VSS.n3460 2.24552
R67926 VSS.n3451 VSS.n3442 2.24552
R67927 VSS.n3463 VSS.n3461 2.24552
R67928 VSS.n3451 VSS.n3441 2.24552
R67929 VSS.n3463 VSS.n3462 2.24552
R67930 VSS.n3451 VSS.n3440 2.24552
R67931 VSS.n3463 VSS.n3439 2.24552
R67932 VSS.n2897 VSS.n2890 2.24552
R67933 VSS.n6876 VSS.n6872 2.24552
R67934 VSS.n2899 VSS.n2890 2.24552
R67935 VSS.n6876 VSS.n6873 2.24552
R67936 VSS.n2901 VSS.n2890 2.24552
R67937 VSS.n6876 VSS.n6874 2.24552
R67938 VSS.n2903 VSS.n2890 2.24552
R67939 VSS.n6876 VSS.n6875 2.24552
R67940 VSS.n2905 VSS.n2890 2.24552
R67941 VSS.n6877 VSS.n6876 2.24552
R67942 VSS.n8410 VSS.n8383 2.24552
R67943 VSS.n8412 VSS.n1660 2.24552
R67944 VSS.n8410 VSS.n8381 2.24552
R67945 VSS.n8412 VSS.n1661 2.24552
R67946 VSS.n1663 VSS.n1655 2.24552
R67947 VSS.n8410 VSS.n8407 2.24552
R67948 VSS.n8412 VSS.n1656 2.24552
R67949 VSS.n8410 VSS.n8409 2.24552
R67950 VSS.n8633 VSS.n8610 2.24552
R67951 VSS.n1537 VSS.n1523 2.24552
R67952 VSS.n8633 VSS.n8612 2.24552
R67953 VSS.n8635 VSS.n1532 2.24552
R67954 VSS.n8633 VSS.n8615 2.24552
R67955 VSS.n8635 VSS.n1531 2.24552
R67956 VSS.n8633 VSS.n8618 2.24552
R67957 VSS.n8635 VSS.n1530 2.24552
R67958 VSS.n8633 VSS.n8621 2.24552
R67959 VSS.n8635 VSS.n1529 2.24552
R67960 VSS.n8633 VSS.n8623 2.24552
R67961 VSS.n8635 VSS.n1527 2.24552
R67962 VSS.n8633 VSS.n8626 2.24552
R67963 VSS.n8635 VSS.n1526 2.24552
R67964 VSS.n8633 VSS.n8629 2.24552
R67965 VSS.n8635 VSS.n1525 2.24552
R67966 VSS.n8633 VSS.n8632 2.24552
R67967 VSS.n8635 VSS.n1524 2.24552
R67968 VSS.n1995 VSS.n1980 2.24552
R67969 VSS.n1996 VSS.n1979 2.24552
R67970 VSS.n8159 VSS.n8150 2.24552
R67971 VSS.n1998 VSS.n1979 2.24552
R67972 VSS.n8159 VSS.n8151 2.24552
R67973 VSS.n2000 VSS.n1979 2.24552
R67974 VSS.n8159 VSS.n8152 2.24552
R67975 VSS.n2002 VSS.n1979 2.24552
R67976 VSS.n8159 VSS.n8153 2.24552
R67977 VSS.n2004 VSS.n1979 2.24552
R67978 VSS.n8159 VSS.n8154 2.24552
R67979 VSS.n2006 VSS.n1979 2.24552
R67980 VSS.n8159 VSS.n8155 2.24552
R67981 VSS.n2008 VSS.n1979 2.24552
R67982 VSS.n8159 VSS.n8156 2.24552
R67983 VSS.n2010 VSS.n1979 2.24552
R67984 VSS.n8159 VSS.n8157 2.24552
R67985 VSS.n2012 VSS.n1979 2.24552
R67986 VSS.n8159 VSS.n8158 2.24552
R67987 VSS.n2014 VSS.n1979 2.24552
R67988 VSS.n8160 VSS.n8159 2.24552
R67989 VSS.n8161 VSS.n1979 2.24552
R67990 VSS.n8159 VSS.n1978 2.24552
R67991 VSS.n8201 VSS.n1955 2.24552
R67992 VSS.n8194 VSS.n8184 2.24552
R67993 VSS.n8201 VSS.n1956 2.24552
R67994 VSS.n8194 VSS.n8183 2.24552
R67995 VSS.n8201 VSS.n1957 2.24552
R67996 VSS.n8194 VSS.n8182 2.24552
R67997 VSS.n8201 VSS.n1958 2.24552
R67998 VSS.n8194 VSS.n8181 2.24552
R67999 VSS.n8201 VSS.n1959 2.24552
R68000 VSS.n8194 VSS.n8180 2.24552
R68001 VSS.n8201 VSS.n1960 2.24552
R68002 VSS.n8194 VSS.n8179 2.24552
R68003 VSS.n8201 VSS.n1961 2.24552
R68004 VSS.n8194 VSS.n8178 2.24552
R68005 VSS.n8201 VSS.n1962 2.24552
R68006 VSS.n8194 VSS.n8177 2.24552
R68007 VSS.n8201 VSS.n1963 2.24552
R68008 VSS.n8194 VSS.n8176 2.24552
R68009 VSS.n8201 VSS.n1964 2.24552
R68010 VSS.n8195 VSS.n8194 2.24552
R68011 VSS.n8201 VSS.n1965 2.24552
R68012 VSS.n8194 VSS.n1967 2.24552
R68013 VSS.n8201 VSS.n8200 2.24552
R68014 VSS.n5235 VSS.n4330 2.24552
R68015 VSS.n5237 VSS.n4331 2.24552
R68016 VSS.n5238 VSS.n4330 2.24552
R68017 VSS.n5240 VSS.n4331 2.24552
R68018 VSS.n5241 VSS.n4330 2.24552
R68019 VSS.n5243 VSS.n4331 2.24552
R68020 VSS.n5296 VSS.n5294 2.24552
R68021 VSS.n5303 VSS.n5265 2.24552
R68022 VSS.n5297 VSS.n5296 2.24552
R68023 VSS.n5303 VSS.n5266 2.24552
R68024 VSS.n5296 VSS.n5268 2.24552
R68025 VSS.n5303 VSS.n5302 2.24552
R68026 VSS.n3956 VSS.n3955 2.24552
R68027 VSS.n6195 VSS.n6193 2.24552
R68028 VSS.n3956 VSS.n3954 2.24552
R68029 VSS.n6195 VSS.n6194 2.24552
R68030 VSS.n3956 VSS.n3953 2.24552
R68031 VSS.n3389 VSS.n3378 2.24552
R68032 VSS.n3377 VSS.n3376 2.24552
R68033 VSS.n3389 VSS.n3379 2.24552
R68034 VSS.n3377 VSS.n3375 2.24552
R68035 VSS.n3389 VSS.n3380 2.24552
R68036 VSS.n3377 VSS.n3374 2.24552
R68037 VSS.n3389 VSS.n3381 2.24552
R68038 VSS.n3377 VSS.n3373 2.24552
R68039 VSS.n3389 VSS.n3382 2.24552
R68040 VSS.n3377 VSS.n3372 2.24552
R68041 VSS.n3389 VSS.n3383 2.24552
R68042 VSS.n3377 VSS.n3371 2.24552
R68043 VSS.n3389 VSS.n3384 2.24552
R68044 VSS.n3377 VSS.n3370 2.24552
R68045 VSS.n3389 VSS.n3385 2.24552
R68046 VSS.n3377 VSS.n3369 2.24552
R68047 VSS.n3389 VSS.n3386 2.24552
R68048 VSS.n3377 VSS.n3368 2.24552
R68049 VSS.n3389 VSS.n3387 2.24552
R68050 VSS.n3377 VSS.n3367 2.24552
R68051 VSS.n3389 VSS.n3388 2.24552
R68052 VSS.n3377 VSS.n3366 2.24552
R68053 VSS.n3389 VSS.n3365 2.24552
R68054 VSS.n2863 VSS.n2856 2.24552
R68055 VSS.n6915 VSS.n6911 2.24552
R68056 VSS.n2865 VSS.n2856 2.24552
R68057 VSS.n6915 VSS.n6912 2.24552
R68058 VSS.n2867 VSS.n2856 2.24552
R68059 VSS.n6915 VSS.n6913 2.24552
R68060 VSS.n2869 VSS.n2856 2.24552
R68061 VSS.n6915 VSS.n6914 2.24552
R68062 VSS.n2871 VSS.n2856 2.24552
R68063 VSS.n6916 VSS.n6915 2.24552
R68064 VSS.n1579 VSS.n1568 2.24552
R68065 VSS.n1581 VSS.n1569 2.24552
R68066 VSS.n1582 VSS.n1568 2.24552
R68067 VSS.n1575 VSS.n1569 2.24552
R68068 VSS.n1573 VSS.n1570 2.24552
R68069 VSS.n1584 VSS.n1568 2.24552
R68070 VSS.n1585 VSS.n1569 2.24552
R68071 VSS.n1587 VSS.n1568 2.24552
R68072 VSS.n8000 VSS.n2091 2.24552
R68073 VSS.n8076 VSS.n2089 2.24552
R68074 VSS.n2123 VSS.n2091 2.24552
R68075 VSS.n8088 VSS.n2121 2.24552
R68076 VSS.n2119 VSS.n2091 2.24552
R68077 VSS.n8088 VSS.n2117 2.24552
R68078 VSS.n2115 VSS.n2091 2.24552
R68079 VSS.n8088 VSS.n2113 2.24552
R68080 VSS.n2111 VSS.n2091 2.24552
R68081 VSS.n8088 VSS.n2109 2.24552
R68082 VSS.n2107 VSS.n2091 2.24552
R68083 VSS.n8088 VSS.n2105 2.24552
R68084 VSS.n2103 VSS.n2091 2.24552
R68085 VSS.n8088 VSS.n2101 2.24552
R68086 VSS.n2099 VSS.n2091 2.24552
R68087 VSS.n8088 VSS.n2097 2.24552
R68088 VSS.n2095 VSS.n2091 2.24552
R68089 VSS.n8088 VSS.n2093 2.24552
R68090 VSS.n8103 VSS.n2048 2.24552
R68091 VSS.n8099 VSS.n2035 2.24552
R68092 VSS.n2049 VSS.n2031 2.24552
R68093 VSS.n2050 VSS.n2035 2.24552
R68094 VSS.n2052 VSS.n2031 2.24552
R68095 VSS.n2053 VSS.n2035 2.24552
R68096 VSS.n2055 VSS.n2031 2.24552
R68097 VSS.n2056 VSS.n2035 2.24552
R68098 VSS.n2058 VSS.n2031 2.24552
R68099 VSS.n2059 VSS.n2035 2.24552
R68100 VSS.n2061 VSS.n2031 2.24552
R68101 VSS.n2062 VSS.n2035 2.24552
R68102 VSS.n2064 VSS.n2031 2.24552
R68103 VSS.n2065 VSS.n2035 2.24552
R68104 VSS.n2067 VSS.n2031 2.24552
R68105 VSS.n2068 VSS.n2035 2.24552
R68106 VSS.n2070 VSS.n2031 2.24552
R68107 VSS.n2071 VSS.n2035 2.24552
R68108 VSS.n2073 VSS.n2031 2.24552
R68109 VSS.n2074 VSS.n2035 2.24552
R68110 VSS.n2076 VSS.n2031 2.24552
R68111 VSS.n2077 VSS.n2035 2.24552
R68112 VSS.n2079 VSS.n2031 2.24552
R68113 VSS.n8231 VSS.n1886 2.24552
R68114 VSS.n8224 VSS.n1928 2.24552
R68115 VSS.n8231 VSS.n1887 2.24552
R68116 VSS.n8224 VSS.n1927 2.24552
R68117 VSS.n8231 VSS.n1888 2.24552
R68118 VSS.n8224 VSS.n1926 2.24552
R68119 VSS.n8231 VSS.n1889 2.24552
R68120 VSS.n8224 VSS.n1925 2.24552
R68121 VSS.n8231 VSS.n1890 2.24552
R68122 VSS.n8224 VSS.n1924 2.24552
R68123 VSS.n8231 VSS.n1891 2.24552
R68124 VSS.n8224 VSS.n1923 2.24552
R68125 VSS.n8231 VSS.n1892 2.24552
R68126 VSS.n8224 VSS.n1922 2.24552
R68127 VSS.n8231 VSS.n1893 2.24552
R68128 VSS.n8224 VSS.n1921 2.24552
R68129 VSS.n8231 VSS.n1894 2.24552
R68130 VSS.n8224 VSS.n1920 2.24552
R68131 VSS.n8231 VSS.n1895 2.24552
R68132 VSS.n8225 VSS.n8224 2.24552
R68133 VSS.n8231 VSS.n1896 2.24552
R68134 VSS.n8224 VSS.n1898 2.24552
R68135 VSS.n8231 VSS.n8230 2.24552
R68136 VSS.n4734 VSS.n4729 2.24552
R68137 VSS.n4764 VSS.n4723 2.24552
R68138 VSS.n4738 VSS.n4729 2.24552
R68139 VSS.n4764 VSS.n4724 2.24552
R68140 VSS.n4740 VSS.n4729 2.24552
R68141 VSS.n4764 VSS.n4725 2.24552
R68142 VSS.n3872 VSS.n3866 2.24552
R68143 VSS.n6240 VSS.n3867 2.24552
R68144 VSS.n6241 VSS.n3866 2.24552
R68145 VSS.n6243 VSS.n3867 2.24552
R68146 VSS.n6244 VSS.n3866 2.24552
R68147 VSS.n6246 VSS.n3867 2.24552
R68148 VSS.n3843 VSS.n3833 2.24552
R68149 VSS.n3845 VSS.n3834 2.24552
R68150 VSS.n3846 VSS.n3833 2.24552
R68151 VSS.n3848 VSS.n3834 2.24552
R68152 VSS.n3849 VSS.n3833 2.24552
R68153 VSS.n6568 VSS.n6558 2.24552
R68154 VSS.n3248 VSS.n3232 2.24552
R68155 VSS.n6568 VSS.n6559 2.24552
R68156 VSS.n3250 VSS.n3232 2.24552
R68157 VSS.n6568 VSS.n6560 2.24552
R68158 VSS.n3252 VSS.n3232 2.24552
R68159 VSS.n6568 VSS.n6561 2.24552
R68160 VSS.n3254 VSS.n3232 2.24552
R68161 VSS.n6568 VSS.n6562 2.24552
R68162 VSS.n3256 VSS.n3232 2.24552
R68163 VSS.n6568 VSS.n6563 2.24552
R68164 VSS.n3258 VSS.n3232 2.24552
R68165 VSS.n6568 VSS.n6564 2.24552
R68166 VSS.n3260 VSS.n3232 2.24552
R68167 VSS.n6568 VSS.n6565 2.24552
R68168 VSS.n3262 VSS.n3232 2.24552
R68169 VSS.n6568 VSS.n6566 2.24552
R68170 VSS.n3264 VSS.n3232 2.24552
R68171 VSS.n6568 VSS.n6567 2.24552
R68172 VSS.n3266 VSS.n3232 2.24552
R68173 VSS.n6569 VSS.n6568 2.24552
R68174 VSS.n6570 VSS.n3232 2.24552
R68175 VSS.n6568 VSS.n3231 2.24552
R68176 VSS.n2806 VSS.n2797 2.24552
R68177 VSS.n6960 VSS.n6957 2.24552
R68178 VSS.n2808 VSS.n2797 2.24552
R68179 VSS.n6960 VSS.n6958 2.24552
R68180 VSS.n2810 VSS.n2797 2.24552
R68181 VSS.n6960 VSS.n6959 2.24552
R68182 VSS.n2812 VSS.n2797 2.24552
R68183 VSS.n6961 VSS.n6960 2.24552
R68184 VSS.n6962 VSS.n2797 2.24552
R68185 VSS.n6960 VSS.n2796 2.24552
R68186 VSS.n8294 VSS.n8292 2.24552
R68187 VSS.n8301 VSS.n1708 2.24552
R68188 VSS.n8294 VSS.n8291 2.24552
R68189 VSS.n8301 VSS.n1709 2.24552
R68190 VSS.n8294 VSS.n8290 2.24552
R68191 VSS.n8301 VSS.n1710 2.24552
R68192 VSS.n8295 VSS.n8294 2.24552
R68193 VSS.n8301 VSS.n1711 2.24552
R68194 VSS.n8294 VSS.n8280 2.24552
R68195 VSS.n8301 VSS.n8300 2.24552
R68196 VSS.n2242 VSS.n1712 2.24552
R68197 VSS.n1728 VSS.n1713 2.24552
R68198 VSS.n2242 VSS.n2232 2.24552
R68199 VSS.n1730 VSS.n1713 2.24552
R68200 VSS.n2242 VSS.n2233 2.24552
R68201 VSS.n1732 VSS.n1713 2.24552
R68202 VSS.n2242 VSS.n2234 2.24552
R68203 VSS.n1734 VSS.n1713 2.24552
R68204 VSS.n2242 VSS.n2235 2.24552
R68205 VSS.n1736 VSS.n1713 2.24552
R68206 VSS.n2242 VSS.n2236 2.24552
R68207 VSS.n1738 VSS.n1713 2.24552
R68208 VSS.n2242 VSS.n2237 2.24552
R68209 VSS.n1740 VSS.n1713 2.24552
R68210 VSS.n2242 VSS.n2238 2.24552
R68211 VSS.n1742 VSS.n1713 2.24552
R68212 VSS.n2242 VSS.n2239 2.24552
R68213 VSS.n1744 VSS.n1713 2.24552
R68214 VSS.n2242 VSS.n2240 2.24552
R68215 VSS.n1746 VSS.n1713 2.24552
R68216 VSS.n2242 VSS.n2241 2.24552
R68217 VSS.n1748 VSS.n1713 2.24552
R68218 VSS.n2242 VSS.n1750 2.24552
R68219 VSS.n7911 VSS.n1751 2.24552
R68220 VSS.n1767 VSS.n1752 2.24552
R68221 VSS.n7911 VSS.n7901 2.24552
R68222 VSS.n1769 VSS.n1752 2.24552
R68223 VSS.n7911 VSS.n7902 2.24552
R68224 VSS.n1771 VSS.n1752 2.24552
R68225 VSS.n7911 VSS.n7903 2.24552
R68226 VSS.n1773 VSS.n1752 2.24552
R68227 VSS.n7911 VSS.n7904 2.24552
R68228 VSS.n1775 VSS.n1752 2.24552
R68229 VSS.n7911 VSS.n7905 2.24552
R68230 VSS.n1777 VSS.n1752 2.24552
R68231 VSS.n7911 VSS.n7906 2.24552
R68232 VSS.n1779 VSS.n1752 2.24552
R68233 VSS.n7911 VSS.n7907 2.24552
R68234 VSS.n1781 VSS.n1752 2.24552
R68235 VSS.n7911 VSS.n7908 2.24552
R68236 VSS.n1783 VSS.n1752 2.24552
R68237 VSS.n7911 VSS.n7909 2.24552
R68238 VSS.n1785 VSS.n1752 2.24552
R68239 VSS.n7911 VSS.n7910 2.24552
R68240 VSS.n1787 VSS.n1752 2.24552
R68241 VSS.n7911 VSS.n1789 2.24552
R68242 VSS.n8268 VSS.n1790 2.24552
R68243 VSS.n1806 VSS.n1791 2.24552
R68244 VSS.n8268 VSS.n8258 2.24552
R68245 VSS.n1808 VSS.n1791 2.24552
R68246 VSS.n8268 VSS.n8259 2.24552
R68247 VSS.n1810 VSS.n1791 2.24552
R68248 VSS.n8268 VSS.n8260 2.24552
R68249 VSS.n1812 VSS.n1791 2.24552
R68250 VSS.n8268 VSS.n8261 2.24552
R68251 VSS.n1814 VSS.n1791 2.24552
R68252 VSS.n8268 VSS.n8262 2.24552
R68253 VSS.n1816 VSS.n1791 2.24552
R68254 VSS.n8268 VSS.n8263 2.24552
R68255 VSS.n1818 VSS.n1791 2.24552
R68256 VSS.n8268 VSS.n8264 2.24552
R68257 VSS.n1820 VSS.n1791 2.24552
R68258 VSS.n8268 VSS.n8265 2.24552
R68259 VSS.n1822 VSS.n1791 2.24552
R68260 VSS.n8268 VSS.n8266 2.24552
R68261 VSS.n1824 VSS.n1791 2.24552
R68262 VSS.n8268 VSS.n8267 2.24552
R68263 VSS.n1826 VSS.n1791 2.24552
R68264 VSS.n8269 VSS.n8268 2.24552
R68265 VSS.n4718 VSS.n4606 2.24552
R68266 VSS.n4597 VSS.n4588 2.24552
R68267 VSS.n4718 VSS.n4605 2.24552
R68268 VSS.n4599 VSS.n4588 2.24552
R68269 VSS.n4718 VSS.n4587 2.24552
R68270 VSS.n4601 VSS.n4589 2.24552
R68271 VSS.n4703 VSS.n4680 2.24552
R68272 VSS.n4631 VSS.n4629 2.24552
R68273 VSS.n4703 VSS.n4679 2.24552
R68274 VSS.n4631 VSS.n4630 2.24552
R68275 VSS.n4703 VSS.n4678 2.24552
R68276 VSS.n4677 VSS.n4676 2.24552
R68277 VSS.n5231 VSS.n4357 2.24552
R68278 VSS.n4348 VSS.n4339 2.24552
R68279 VSS.n5231 VSS.n4356 2.24552
R68280 VSS.n4350 VSS.n4339 2.24552
R68281 VSS.n5231 VSS.n4338 2.24552
R68282 VSS.n4352 VSS.n4340 2.24552
R68283 VSS.n5204 VSS.n4400 2.24552
R68284 VSS.n4394 VSS.n4392 2.24552
R68285 VSS.n5204 VSS.n4399 2.24552
R68286 VSS.n4394 VSS.n4393 2.24552
R68287 VSS.n5204 VSS.n4398 2.24552
R68288 VSS.n4397 VSS.n4396 2.24552
R68289 VSS.n9889 VSS.n32 2.24552
R68290 VSS.n42 VSS.n33 2.24552
R68291 VSS.n9889 VSS.n45 2.24552
R68292 VSS.n44 VSS.n33 2.24552
R68293 VSS.n9890 VSS.n9889 2.24552
R68294 VSS.n36 VSS.n34 2.24552
R68295 VSS.n9862 VSS.n88 2.24552
R68296 VSS.n82 VSS.n80 2.24552
R68297 VSS.n9862 VSS.n87 2.24552
R68298 VSS.n82 VSS.n81 2.24552
R68299 VSS.n9862 VSS.n86 2.24552
R68300 VSS.n85 VSS.n84 2.24552
R68301 VSS.n146 VSS.n145 2.24552
R68302 VSS.n9832 VSS.n9830 2.24552
R68303 VSS.n146 VSS.n144 2.24552
R68304 VSS.n9832 VSS.n9831 2.24552
R68305 VSS.n146 VSS.n143 2.24552
R68306 VSS.n9798 VSS.n177 2.24552
R68307 VSS.n9800 VSS.n178 2.24552
R68308 VSS.n9801 VSS.n177 2.24552
R68309 VSS.n9803 VSS.n178 2.24552
R68310 VSS.n9804 VSS.n177 2.24552
R68311 VSS.n9806 VSS.n178 2.24552
R68312 VSS.n5474 VSS.n5431 2.24552
R68313 VSS.n5482 VSS.n5480 2.24552
R68314 VSS.n5476 VSS.n5431 2.24552
R68315 VSS.n5482 VSS.n5481 2.24552
R68316 VSS.n5478 VSS.n5431 2.24552
R68317 VSS.n5483 VSS.n5482 2.24552
R68318 VSS.n414 VSS.n407 2.24552
R68319 VSS.n425 VSS.n423 2.24552
R68320 VSS.n416 VSS.n407 2.24552
R68321 VSS.n425 VSS.n424 2.24552
R68322 VSS.n418 VSS.n407 2.24552
R68323 VSS.n6384 VSS.n444 2.24552
R68324 VSS.n460 VSS.n445 2.24552
R68325 VSS.n6384 VSS.n6374 2.24552
R68326 VSS.n462 VSS.n445 2.24552
R68327 VSS.n6384 VSS.n6375 2.24552
R68328 VSS.n464 VSS.n445 2.24552
R68329 VSS.n6384 VSS.n6376 2.24552
R68330 VSS.n466 VSS.n445 2.24552
R68331 VSS.n6384 VSS.n6377 2.24552
R68332 VSS.n468 VSS.n445 2.24552
R68333 VSS.n6384 VSS.n6378 2.24552
R68334 VSS.n470 VSS.n445 2.24552
R68335 VSS.n6384 VSS.n6379 2.24552
R68336 VSS.n472 VSS.n445 2.24552
R68337 VSS.n6384 VSS.n6380 2.24552
R68338 VSS.n474 VSS.n445 2.24552
R68339 VSS.n6384 VSS.n6381 2.24552
R68340 VSS.n476 VSS.n445 2.24552
R68341 VSS.n6384 VSS.n6382 2.24552
R68342 VSS.n478 VSS.n445 2.24552
R68343 VSS.n6384 VSS.n6383 2.24552
R68344 VSS.n480 VSS.n445 2.24552
R68345 VSS.n6384 VSS.n482 2.24552
R68346 VSS.n524 VSS.n501 2.24552
R68347 VSS.n511 VSS.n502 2.24552
R68348 VSS.n524 VSS.n523 2.24552
R68349 VSS.n513 VSS.n502 2.24552
R68350 VSS.n524 VSS.n522 2.24552
R68351 VSS.n515 VSS.n502 2.24552
R68352 VSS.n524 VSS.n521 2.24552
R68353 VSS.n517 VSS.n502 2.24552
R68354 VSS.n524 VSS.n520 2.24552
R68355 VSS.n519 VSS.n502 2.24552
R68356 VSS.n562 VSS.n539 2.24552
R68357 VSS.n549 VSS.n540 2.24552
R68358 VSS.n562 VSS.n561 2.24552
R68359 VSS.n551 VSS.n540 2.24552
R68360 VSS.n562 VSS.n560 2.24552
R68361 VSS.n553 VSS.n540 2.24552
R68362 VSS.n562 VSS.n559 2.24552
R68363 VSS.n555 VSS.n540 2.24552
R68364 VSS.n562 VSS.n558 2.24552
R68365 VSS.n557 VSS.n540 2.24552
R68366 VSS.n8936 VSS.n563 2.24552
R68367 VSS.n579 VSS.n564 2.24552
R68368 VSS.n8936 VSS.n8926 2.24552
R68369 VSS.n581 VSS.n564 2.24552
R68370 VSS.n8936 VSS.n8927 2.24552
R68371 VSS.n583 VSS.n564 2.24552
R68372 VSS.n8936 VSS.n8928 2.24552
R68373 VSS.n585 VSS.n564 2.24552
R68374 VSS.n8936 VSS.n8929 2.24552
R68375 VSS.n587 VSS.n564 2.24552
R68376 VSS.n8936 VSS.n8930 2.24552
R68377 VSS.n589 VSS.n564 2.24552
R68378 VSS.n8936 VSS.n8931 2.24552
R68379 VSS.n591 VSS.n564 2.24552
R68380 VSS.n8936 VSS.n8932 2.24552
R68381 VSS.n593 VSS.n564 2.24552
R68382 VSS.n8936 VSS.n8933 2.24552
R68383 VSS.n595 VSS.n564 2.24552
R68384 VSS.n8936 VSS.n8934 2.24552
R68385 VSS.n597 VSS.n564 2.24552
R68386 VSS.n8936 VSS.n8935 2.24552
R68387 VSS.n599 VSS.n564 2.24552
R68388 VSS.n8936 VSS.n601 2.24552
R68389 VSS.n9483 VSS.n602 2.24552
R68390 VSS.n617 VSS.n603 2.24552
R68391 VSS.n9483 VSS.n9473 2.24552
R68392 VSS.n619 VSS.n603 2.24552
R68393 VSS.n9483 VSS.n9474 2.24552
R68394 VSS.n621 VSS.n603 2.24552
R68395 VSS.n9483 VSS.n9475 2.24552
R68396 VSS.n623 VSS.n603 2.24552
R68397 VSS.n9483 VSS.n9476 2.24552
R68398 VSS.n625 VSS.n603 2.24552
R68399 VSS.n9483 VSS.n9477 2.24552
R68400 VSS.n627 VSS.n603 2.24552
R68401 VSS.n9483 VSS.n9478 2.24552
R68402 VSS.n629 VSS.n603 2.24552
R68403 VSS.n9483 VSS.n9479 2.24552
R68404 VSS.n631 VSS.n603 2.24552
R68405 VSS.n9483 VSS.n9480 2.24552
R68406 VSS.n633 VSS.n603 2.24552
R68407 VSS.n9483 VSS.n9481 2.24552
R68408 VSS.n635 VSS.n603 2.24552
R68409 VSS.n9483 VSS.n9482 2.24552
R68410 VSS.n637 VSS.n603 2.24552
R68411 VSS.n9483 VSS.n639 2.24552
R68412 VSS.n9557 VSS.n640 2.24552
R68413 VSS.n656 VSS.n641 2.24552
R68414 VSS.n9557 VSS.n9547 2.24552
R68415 VSS.n658 VSS.n641 2.24552
R68416 VSS.n9557 VSS.n9548 2.24552
R68417 VSS.n660 VSS.n641 2.24552
R68418 VSS.n9557 VSS.n9549 2.24552
R68419 VSS.n662 VSS.n641 2.24552
R68420 VSS.n9557 VSS.n9550 2.24552
R68421 VSS.n664 VSS.n641 2.24552
R68422 VSS.n9557 VSS.n9551 2.24552
R68423 VSS.n666 VSS.n641 2.24552
R68424 VSS.n9557 VSS.n9552 2.24552
R68425 VSS.n668 VSS.n641 2.24552
R68426 VSS.n9557 VSS.n9553 2.24552
R68427 VSS.n670 VSS.n641 2.24552
R68428 VSS.n9557 VSS.n9554 2.24552
R68429 VSS.n672 VSS.n641 2.24552
R68430 VSS.n9557 VSS.n9555 2.24552
R68431 VSS.n674 VSS.n641 2.24552
R68432 VSS.n9557 VSS.n9556 2.24552
R68433 VSS.n676 VSS.n641 2.24552
R68434 VSS.n9558 VSS.n9557 2.24552
R68435 VSS.n146 VSS.n142 2.24552
R68436 VSS.n6048 VSS.n6046 2.24552
R68437 VSS.n6040 VSS.n6038 2.24552
R68438 VSS.n5946 VSS.n5915 2.24552
R68439 VSS.n5938 VSS.n5922 2.24552
R68440 VSS.n6064 VSS.n6063 2.24552
R68441 VSS.n6071 VSS.n6070 2.24552
R68442 VSS.n5952 VSS.n5910 2.24552
R68443 VSS.n5944 VSS.n5917 2.24552
R68444 VSS.n6052 VSS.n6046 2.24552
R68445 VSS.n6044 VSS.n6038 2.24552
R68446 VSS.n5915 VSS.n5912 2.24552
R68447 VSS.n5922 VSS.n5919 2.24552
R68448 VSS.n6064 VSS.n6051 2.24552
R68449 VSS.n6071 VSS.n6043 2.24552
R68450 VSS.n5952 VSS.n5951 2.24552
R68451 VSS.n5944 VSS.n5943 2.24552
R68452 VSS.n3812 VSS.n3809 2.24552
R68453 VSS.n3803 VSS.n3800 2.24552
R68454 VSS.n3699 VSS.n3696 2.24552
R68455 VSS.n3690 VSS.n3687 2.24552
R68456 VSS.n6290 VSS.n6289 2.24552
R68457 VSS.n6297 VSS.n6296 2.24552
R68458 VSS.n6319 VSS.n6318 2.24552
R68459 VSS.n6326 VSS.n6325 2.24552
R68460 VSS.n3816 VSS.n3809 2.24552
R68461 VSS.n3807 VSS.n3800 2.24552
R68462 VSS.n3703 VSS.n3696 2.24552
R68463 VSS.n3694 VSS.n3687 2.24552
R68464 VSS.n6290 VSS.n3815 2.24552
R68465 VSS.n6297 VSS.n3806 2.24552
R68466 VSS.n6319 VSS.n3702 2.24552
R68467 VSS.n6326 VSS.n3693 2.24552
R68468 VSS.n3218 VSS.n3215 2.24552
R68469 VSS.n3209 VSS.n3206 2.24552
R68470 VSS.n3200 VSS.n3197 2.24552
R68471 VSS.n3121 VSS.n3119 2.24552
R68472 VSS.n3115 VSS.n3113 2.24552
R68473 VSS.n6584 VSS.n6583 2.24552
R68474 VSS.n6590 VSS.n6589 2.24552
R68475 VSS.n6597 VSS.n6596 2.24552
R68476 VSS.n6625 VSS.n6624 2.24552
R68477 VSS.n6632 VSS.n6631 2.24552
R68478 VSS.n3222 VSS.n3215 2.24552
R68479 VSS.n3213 VSS.n3206 2.24552
R68480 VSS.n3204 VSS.n3197 2.24552
R68481 VSS.n3125 VSS.n3119 2.24552
R68482 VSS.n6634 VSS.n3115 2.24552
R68483 VSS.n6584 VSS.n3221 2.24552
R68484 VSS.n6590 VSS.n3212 2.24552
R68485 VSS.n6597 VSS.n3203 2.24552
R68486 VSS.n6625 VSS.n3124 2.24552
R68487 VSS.n6633 VSS.n6632 2.24552
R68488 VSS.n5761 VSS.n5758 2.24552
R68489 VSS.n5752 VSS.n5749 2.24552
R68490 VSS.n5743 VSS.n5740 2.24552
R68491 VSS.n2971 VSS.n2968 2.24552
R68492 VSS.n6642 VSS.n3112 2.24552
R68493 VSS.n5782 VSS.n5781 2.24552
R68494 VSS.n5788 VSS.n5787 2.24552
R68495 VSS.n5795 VSS.n5794 2.24552
R68496 VSS.n6760 VSS.n2963 2.24552
R68497 VSS.n6649 VSS.n6648 2.24552
R68498 VSS.n5765 VSS.n5758 2.24552
R68499 VSS.n5756 VSS.n5749 2.24552
R68500 VSS.n5747 VSS.n5740 2.24552
R68501 VSS.n6754 VSS.n2968 2.24552
R68502 VSS.n6646 VSS.n3112 2.24552
R68503 VSS.n5782 VSS.n5764 2.24552
R68504 VSS.n5788 VSS.n5755 2.24552
R68505 VSS.n5795 VSS.n5746 2.24552
R68506 VSS.n6760 VSS.n6759 2.24552
R68507 VSS.n6649 VSS.n6645 2.24552
R68508 VSS.n2762 VSS.n2759 2.24552
R68509 VSS.n2753 VSS.n2750 2.24552
R68510 VSS.n2744 VSS.n2741 2.24552
R68511 VSS.n2637 VSS.n2634 2.24552
R68512 VSS.n2628 VSS.n2625 2.24552
R68513 VSS.n6976 VSS.n6975 2.24552
R68514 VSS.n6982 VSS.n6981 2.24552
R68515 VSS.n6989 VSS.n6988 2.24552
R68516 VSS.n7011 VSS.n7010 2.24552
R68517 VSS.n7018 VSS.n7017 2.24552
R68518 VSS.n2766 VSS.n2759 2.24552
R68519 VSS.n2757 VSS.n2750 2.24552
R68520 VSS.n2748 VSS.n2741 2.24552
R68521 VSS.n2641 VSS.n2634 2.24552
R68522 VSS.n2632 VSS.n2625 2.24552
R68523 VSS.n6976 VSS.n2765 2.24552
R68524 VSS.n6982 VSS.n2756 2.24552
R68525 VSS.n6989 VSS.n2747 2.24552
R68526 VSS.n7011 VSS.n2640 2.24552
R68527 VSS.n7018 VSS.n2631 2.24552
R68528 VSS.n2621 VSS.n2619 2.24552
R68529 VSS.n7024 VSS.n7023 2.24552
R68530 VSS.n7026 VSS.n2621 2.24552
R68531 VSS.n3108 VSS.n3106 2.24552
R68532 VSS.n6655 VSS.n6654 2.24552
R68533 VSS.n6657 VSS.n3108 2.24552
R68534 VSS.n3658 VSS.n3656 2.24552
R68535 VSS.n3663 VSS.n3662 2.24552
R68536 VSS.n3661 VSS.n3656 2.24552
R68537 VSS.n3683 VSS.n3681 2.24552
R68538 VSS.n6332 VSS.n6331 2.24552
R68539 VSS.n6334 VSS.n3683 2.24552
R68540 VSS.n5931 VSS.n5929 2.24552
R68541 VSS.n5937 VSS.n5924 2.24552
R68542 VSS.n5929 VSS.n5926 2.24552
R68543 VSS.n5937 VSS.n5936 2.24552
R68544 VSS.n6333 VSS.n6332 2.24552
R68545 VSS.n3663 VSS.n3655 2.24552
R68546 VSS.n6656 VSS.n6655 2.24552
R68547 VSS.n7025 VSS.n7024 2.24552
R68548 VSS.n9847 VSS.n119 2.24552
R68549 VSS.n113 VSS.n111 2.24552
R68550 VSS.n9847 VSS.n118 2.24552
R68551 VSS.n113 VSS.n112 2.24552
R68552 VSS.n9847 VSS.n117 2.24552
R68553 VSS.n209 VSS.n204 2.24552
R68554 VSS.n9778 VSS.n198 2.24552
R68555 VSS.n212 VSS.n204 2.24552
R68556 VSS.n9778 VSS.n199 2.24552
R68557 VSS.n214 VSS.n204 2.24552
R68558 VSS.n9778 VSS.n200 2.24552
R68559 VSS.n5416 VSS.n5407 2.24552
R68560 VSS.n5503 VSS.n5501 2.24552
R68561 VSS.n5418 VSS.n5407 2.24552
R68562 VSS.n5503 VSS.n5502 2.24552
R68563 VSS.n5420 VSS.n5407 2.24552
R68564 VSS.n5504 VSS.n5503 2.24552
R68565 VSS.n388 VSS.n381 2.24552
R68566 VSS.n9626 VSS.n9624 2.24552
R68567 VSS.n390 VSS.n381 2.24552
R68568 VSS.n9626 VSS.n9625 2.24552
R68569 VSS.n392 VSS.n381 2.24552
R68570 VSS.n6403 VSS.n3643 2.24552
R68571 VSS.n6396 VSS.n6359 2.24552
R68572 VSS.n6403 VSS.n3644 2.24552
R68573 VSS.n6396 VSS.n6358 2.24552
R68574 VSS.n6403 VSS.n3645 2.24552
R68575 VSS.n6396 VSS.n6357 2.24552
R68576 VSS.n6403 VSS.n3646 2.24552
R68577 VSS.n6396 VSS.n6356 2.24552
R68578 VSS.n6403 VSS.n3647 2.24552
R68579 VSS.n6396 VSS.n6355 2.24552
R68580 VSS.n6403 VSS.n3648 2.24552
R68581 VSS.n6396 VSS.n6354 2.24552
R68582 VSS.n6403 VSS.n3649 2.24552
R68583 VSS.n6396 VSS.n6353 2.24552
R68584 VSS.n6403 VSS.n3650 2.24552
R68585 VSS.n6396 VSS.n6352 2.24552
R68586 VSS.n6403 VSS.n3651 2.24552
R68587 VSS.n6396 VSS.n6351 2.24552
R68588 VSS.n6403 VSS.n3652 2.24552
R68589 VSS.n6397 VSS.n6396 2.24552
R68590 VSS.n6403 VSS.n3653 2.24552
R68591 VSS.n6396 VSS.n3670 2.24552
R68592 VSS.n6403 VSS.n6402 2.24552
R68593 VSS.n6699 VSS.n3097 2.24552
R68594 VSS.n6694 VSS.n6691 2.24552
R68595 VSS.n6699 VSS.n3096 2.24552
R68596 VSS.n6694 VSS.n6692 2.24552
R68597 VSS.n6699 VSS.n3095 2.24552
R68598 VSS.n6694 VSS.n6693 2.24552
R68599 VSS.n6699 VSS.n3094 2.24552
R68600 VSS.n6695 VSS.n6694 2.24552
R68601 VSS.n6699 VSS.n3093 2.24552
R68602 VSS.n6694 VSS.n3099 2.24552
R68603 VSS.n1268 VSS.n1259 2.24552
R68604 VSS.n8905 VSS.n8902 2.24552
R68605 VSS.n1270 VSS.n1259 2.24552
R68606 VSS.n8905 VSS.n8903 2.24552
R68607 VSS.n1272 VSS.n1259 2.24552
R68608 VSS.n8905 VSS.n8904 2.24552
R68609 VSS.n1274 VSS.n1259 2.24552
R68610 VSS.n8906 VSS.n8905 2.24552
R68611 VSS.n8907 VSS.n1259 2.24552
R68612 VSS.n8905 VSS.n1258 2.24552
R68613 VSS.n8950 VSS.n1153 2.24552
R68614 VSS.n8948 VSS.n1257 2.24552
R68615 VSS.n8950 VSS.n1154 2.24552
R68616 VSS.n8948 VSS.n1254 2.24552
R68617 VSS.n8950 VSS.n1155 2.24552
R68618 VSS.n8948 VSS.n1251 2.24552
R68619 VSS.n8950 VSS.n1156 2.24552
R68620 VSS.n8948 VSS.n1248 2.24552
R68621 VSS.n8950 VSS.n1157 2.24552
R68622 VSS.n8948 VSS.n1245 2.24552
R68623 VSS.n8950 VSS.n1158 2.24552
R68624 VSS.n8948 VSS.n1242 2.24552
R68625 VSS.n8950 VSS.n1159 2.24552
R68626 VSS.n8948 VSS.n1239 2.24552
R68627 VSS.n8950 VSS.n1160 2.24552
R68628 VSS.n8948 VSS.n1236 2.24552
R68629 VSS.n8950 VSS.n1161 2.24552
R68630 VSS.n8948 VSS.n1233 2.24552
R68631 VSS.n8950 VSS.n1162 2.24552
R68632 VSS.n8948 VSS.n1230 2.24552
R68633 VSS.n8950 VSS.n1163 2.24552
R68634 VSS.n8948 VSS.n1227 2.24552
R68635 VSS.n116 VSS.n115 2.24552
R68636 VSS.n2362 VSS.n2339 2.24552
R68637 VSS.n2357 VSS.n2346 2.24552
R68638 VSS.n9442 VSS.n774 2.24552
R68639 VSS.n9437 VSS.n9371 2.24552
R68640 VSS.n2366 VSS.n2336 2.24552
R68641 VSS.n2361 VSS.n2343 2.24552
R68642 VSS.n9446 VSS.n770 2.24552
R68643 VSS.n9441 VSS.n778 2.24552
R68644 VSS.n2339 VSS.n2337 2.24552
R68645 VSS.n2346 VSS.n2344 2.24552
R68646 VSS.n774 VSS.n772 2.24552
R68647 VSS.n9371 VSS.n9369 2.24552
R68648 VSS.n8093 VSS.n2081 2.24552
R68649 VSS.n2437 VSS.n2436 2.24552
R68650 VSS.n2456 VSS.n2452 2.24552
R68651 VSS.n8967 VSS.n1091 2.24552
R68652 VSS.n2088 VSS.n2087 2.24552
R68653 VSS.n2431 VSS.n2084 2.24552
R68654 VSS.n2461 VSS.n2460 2.24552
R68655 VSS.n1098 VSS.n1097 2.24552
R68656 VSS.n7077 VSS.n7065 2.24531
R68657 VSS.n7210 VSS.n7209 2.24531
R68658 VSS.n7216 VSS.n2533 2.24531
R68659 VSS.n7062 VSS.n7060 2.24531
R68660 VSS.n7064 VSS.n2519 2.24531
R68661 VSS.n2545 VSS.n2542 2.24531
R68662 VSS.n7173 VSS.n7172 2.24531
R68663 VSS.n2558 VSS.n2556 2.24531
R68664 VSS.n1609 VSS.n1386 2.24531
R68665 VSS.n1611 VSS.n1610 2.24531
R68666 VSS.n8052 VSS.n8025 2.24531
R68667 VSS.n1366 VSS.n1364 2.24531
R68668 VSS.n2601 VSS.n2600 2.24531
R68669 VSS.n2597 VSS.n2595 2.24531
R68670 VSS.n8397 VSS.n8395 2.24531
R68671 VSS.n8540 VSS.n1608 2.24531
R68672 VSS.n1607 VSS.n1606 2.24531
R68673 VSS.n8060 VSS.n8021 2.24531
R68674 VSS.n2475 VSS.n2473 2.24531
R68675 VSS.n2517 VSS.n2514 2.24531
R68676 VSS.n7183 VSS.n2537 2.24531
R68677 VSS.n7176 VSS.n2540 2.24531
R68678 VSS.n2538 VSS.n2487 2.24531
R68679 VSS.n7199 VSS.n7185 2.24531
R68680 VSS.n7235 VSS.n7234 2.24531
R68681 VSS.n7067 VSS.n7066 2.24531
R68682 VSS.n7142 VSS.n2472 2.24531
R68683 VSS.n7140 VSS.n2471 2.24531
R68684 VSS.n7150 VSS.n7149 2.24531
R68685 VSS.n2341 VSS.n2335 2.24505
R68686 VSS.n2348 VSS.n2342 2.24505
R68687 VSS.n776 VSS.n769 2.24505
R68688 VSS.n9373 VSS.n777 2.24505
R68689 VSS.n8096 VSS.n2082 2.24505
R68690 VSS.n2433 VSS.n2430 2.24505
R68691 VSS.n2454 VSS.n2451 2.24505
R68692 VSS.n8970 VSS.n1092 2.24505
R68693 VSS.n8092 VSS.n2083 2.24505
R68694 VSS.n2435 VSS.n1542 2.24505
R68695 VSS.n2427 VSS.n1496 2.24505
R68696 VSS.n2450 VSS.n1463 2.24505
R68697 VSS.n2455 VSS.n1429 2.24505
R68698 VSS.n8966 VSS.n1093 2.24505
R68699 VSS.n8094 VSS.n8090 2.24505
R68700 VSS.n2438 VSS.n1540 2.24505
R68701 VSS.n2441 VSS.n1493 2.24505
R68702 VSS.n2447 VSS.n1460 2.24505
R68703 VSS.n2457 VSS.n1428 2.24505
R68704 VSS.n8968 VSS.n8964 2.24505
R68705 VSS.n7208 VSS.n2535 2.24456
R68706 VSS.n7213 VSS.n7212 2.24456
R68707 VSS.n7218 VSS.n2528 2.24456
R68708 VSS.n7080 VSS.n7061 2.24456
R68709 VSS.n7091 VSS.n2532 2.24456
R68710 VSS.n2546 VSS.n2541 2.24456
R68711 VSS.n7166 VSS.n2547 2.24456
R68712 VSS.n7237 VSS.n2511 2.24456
R68713 VSS.n7193 VSS.n2491 2.24456
R68714 VSS.n7259 VSS.n2484 2.24456
R68715 VSS.n8557 VSS.n1589 2.24456
R68716 VSS.n8557 VSS.n1588 2.24456
R68717 VSS.n8547 VSS.n1597 2.24456
R68718 VSS.n8810 VSS.n1387 2.24456
R68719 VSS.n8840 VSS.n1344 2.24456
R68720 VSS.n1350 VSS.n1305 2.24456
R68721 VSS.n8552 VSS.n1590 2.24456
R68722 VSS.n8073 VSS.n8072 2.24456
R68723 VSS.n8067 VSS.n8012 2.24456
R68724 VSS.n8053 VSS.n8023 2.24456
R68725 VSS.n8048 VSS.n8027 2.24456
R68726 VSS.n8043 VSS.n8034 2.24456
R68727 VSS.n8038 VSS.n8033 2.24456
R68728 VSS.n8030 VSS.n8026 2.24456
R68729 VSS.n8015 VSS.n8011 2.24456
R68730 VSS.n8008 VSS.n8007 2.24456
R68731 VSS.n8561 VSS.n1560 2.24456
R68732 VSS.n8562 VSS.n8561 2.24456
R68733 VSS.n8404 VSS.n8386 2.24456
R68734 VSS.n8404 VSS.n8385 2.24456
R68735 VSS.n8818 VSS.n1365 2.24456
R68736 VSS.n8846 VSS.n1315 2.24456
R68737 VSS.n1319 VSS.n1315 2.24456
R68738 VSS.n8855 VSS.n8854 2.24456
R68739 VSS.n8854 VSS.n8853 2.24456
R68740 VSS.n8851 VSS.n8850 2.24456
R68741 VSS.n8844 VSS.n1314 2.24456
R68742 VSS.n8819 VSS.n1363 2.24456
R68743 VSS.n8393 VSS.n8392 2.24456
R68744 VSS.n1564 VSS.n1559 2.24456
R68745 VSS.n8398 VSS.n8396 2.24456
R68746 VSS.n8399 VSS.n8394 2.24456
R68747 VSS.n8541 VSS.n1605 2.24456
R68748 VSS.n8061 VSS.n8019 2.24456
R68749 VSS.n2518 VSS.n2512 2.24456
R68750 VSS.n7200 VSS.n7182 2.24456
R68751 VSS.n7177 VSS.n2478 2.24456
R68752 VSS.n7215 VSS.n2534 2.24456
R68753 VSS.n7222 VSS.n7221 2.24456
R68754 VSS.n7083 VSS.n7082 2.24456
R68755 VSS.n7096 VSS.n7086 2.24456
R68756 VSS.n2544 VSS.n2536 2.24456
R68757 VSS.n7168 VSS.n2550 2.24456
R68758 VSS.n7257 VSS.n7256 2.24456
R68759 VSS.n7197 VSS.n7196 2.24456
R68760 VSS.n7242 VSS.n2509 2.24456
R68761 VSS.n8837 VSS.n8832 2.24456
R68762 VSS.n8807 VSS.n1347 2.24456
R68763 VSS.n1612 VSS.n1388 2.24456
R68764 VSS.n8549 VSS.n1599 2.24456
R68765 VSS.n8045 VSS.n8037 2.24456
R68766 VSS.n8050 VSS.n8029 2.24456
R68767 VSS.n8056 VSS.n8055 2.24456
R68768 VSS.n8069 VSS.n8014 2.24456
R68769 VSS.n8075 VSS.n8003 2.24456
R68770 VSS.n8544 VSS.n8543 2.24456
R68771 VSS.n8064 VSS.n8063 2.24456
R68772 VSS.n7181 VSS.n2539 2.24456
R68773 VSS.n7203 VSS.n7202 2.24456
R68774 VSS.n2516 VSS.n2513 2.24456
R68775 VSS.n4872 VSS.n4871 2.24447
R68776 VSS.n4256 VSS.n4245 2.24447
R68777 VSS.n5720 VSS.n4170 2.24447
R68778 VSS.n3161 VSS.n3134 2.24447
R68779 VSS.n8816 VSS.n1375 2.24447
R68780 VSS.n8814 VSS.n8812 2.24447
R68781 VSS.n8816 VSS.n1374 2.24447
R68782 VSS.n8812 VSS.n1384 2.24447
R68783 VSS.n8816 VSS.n1372 2.24447
R68784 VSS.n8812 VSS.n1367 2.24447
R68785 VSS.n8816 VSS.n1370 2.24447
R68786 VSS.n8812 VSS.n1381 2.24447
R68787 VSS.n1462 VSS.n1461 2.24447
R68788 VSS.n8712 VSS.n1450 2.24447
R68789 VSS.n1472 VSS.n1462 2.24447
R68790 VSS.n8712 VSS.n1449 2.24447
R68791 VSS.n8694 VSS.n1462 2.24447
R68792 VSS.n8712 VSS.n1448 2.24447
R68793 VSS.n8696 VSS.n1462 2.24447
R68794 VSS.n8712 VSS.n1447 2.24447
R68795 VSS.n8698 VSS.n1462 2.24447
R68796 VSS.n8700 VSS.n1462 2.24447
R68797 VSS.n8712 VSS.n1456 2.24447
R68798 VSS.n8702 VSS.n1462 2.24447
R68799 VSS.n8712 VSS.n1457 2.24447
R68800 VSS.n8704 VSS.n1462 2.24447
R68801 VSS.n8712 VSS.n1458 2.24447
R68802 VSS.n8706 VSS.n1462 2.24447
R68803 VSS.n8712 VSS.n1459 2.24447
R68804 VSS.n8708 VSS.n1462 2.24447
R68805 VSS.n9109 VSS.n9081 2.24447
R68806 VSS.n9114 VSS.n983 2.24447
R68807 VSS.n9109 VSS.n9084 2.24447
R68808 VSS.n9114 VSS.n984 2.24447
R68809 VSS.n9109 VSS.n9087 2.24447
R68810 VSS.n9114 VSS.n985 2.24447
R68811 VSS.n9109 VSS.n9090 2.24447
R68812 VSS.n9114 VSS.n986 2.24447
R68813 VSS.n9109 VSS.n9093 2.24447
R68814 VSS.n9114 VSS.n987 2.24447
R68815 VSS.n9109 VSS.n9096 2.24447
R68816 VSS.n9114 VSS.n988 2.24447
R68817 VSS.n9109 VSS.n9099 2.24447
R68818 VSS.n9114 VSS.n989 2.24447
R68819 VSS.n9109 VSS.n9102 2.24447
R68820 VSS.n9114 VSS.n990 2.24447
R68821 VSS.n9109 VSS.n9105 2.24447
R68822 VSS.n9114 VSS.n991 2.24447
R68823 VSS.n9109 VSS.n9108 2.24447
R68824 VSS.n9114 VSS.n992 2.24447
R68825 VSS.n9111 VSS.n9109 2.24447
R68826 VSS.n9114 VSS.n993 2.24447
R68827 VSS.n9114 VSS.n9113 2.24447
R68828 VSS.n9256 VSS.n875 2.24447
R68829 VSS.n9250 VSS.n9240 2.24447
R68830 VSS.n9256 VSS.n876 2.24447
R68831 VSS.n9250 VSS.n9241 2.24447
R68832 VSS.n9256 VSS.n877 2.24447
R68833 VSS.n9250 VSS.n9242 2.24447
R68834 VSS.n9256 VSS.n878 2.24447
R68835 VSS.n9250 VSS.n9243 2.24447
R68836 VSS.n9256 VSS.n879 2.24447
R68837 VSS.n9250 VSS.n9244 2.24447
R68838 VSS.n9256 VSS.n880 2.24447
R68839 VSS.n9250 VSS.n9245 2.24447
R68840 VSS.n9256 VSS.n881 2.24447
R68841 VSS.n9250 VSS.n9246 2.24447
R68842 VSS.n9256 VSS.n882 2.24447
R68843 VSS.n9250 VSS.n9247 2.24447
R68844 VSS.n9256 VSS.n883 2.24447
R68845 VSS.n9250 VSS.n9248 2.24447
R68846 VSS.n9256 VSS.n884 2.24447
R68847 VSS.n9251 VSS.n9250 2.24447
R68848 VSS.n9256 VSS.n9255 2.24447
R68849 VSS.n9250 VSS.n886 2.24447
R68850 VSS.n9250 VSS.n9249 2.24447
R68851 VSS.n4502 VSS.n4491 2.24447
R68852 VSS.n5654 VSS.n4262 2.24447
R68853 VSS.n4023 VSS.n4014 2.24447
R68854 VSS.n6480 VSS.n3164 2.24447
R68855 VSS.n8535 VSS.n1636 2.24447
R68856 VSS.n1626 VSS.n1617 2.24447
R68857 VSS.n8535 VSS.n1635 2.24447
R68858 VSS.n1628 VSS.n1617 2.24447
R68859 VSS.n8536 VSS.n8535 2.24447
R68860 VSS.n1631 VSS.n1617 2.24447
R68861 VSS.n8535 VSS.n1618 2.24447
R68862 VSS.n1633 VSS.n1617 2.24447
R68863 VSS.n1495 VSS.n1494 2.24447
R68864 VSS.n8686 VSS.n1483 2.24447
R68865 VSS.n1505 VSS.n1495 2.24447
R68866 VSS.n8686 VSS.n1482 2.24447
R68867 VSS.n8668 VSS.n1495 2.24447
R68868 VSS.n8686 VSS.n1481 2.24447
R68869 VSS.n8670 VSS.n1495 2.24447
R68870 VSS.n8686 VSS.n1480 2.24447
R68871 VSS.n8672 VSS.n1495 2.24447
R68872 VSS.n8674 VSS.n1495 2.24447
R68873 VSS.n8686 VSS.n1489 2.24447
R68874 VSS.n8676 VSS.n1495 2.24447
R68875 VSS.n8686 VSS.n1490 2.24447
R68876 VSS.n8678 VSS.n1495 2.24447
R68877 VSS.n8686 VSS.n1491 2.24447
R68878 VSS.n8680 VSS.n1495 2.24447
R68879 VSS.n8686 VSS.n1492 2.24447
R68880 VSS.n8682 VSS.n1495 2.24447
R68881 VSS.n9150 VSS.n9122 2.24447
R68882 VSS.n9155 VSS.n962 2.24447
R68883 VSS.n9150 VSS.n9125 2.24447
R68884 VSS.n9155 VSS.n963 2.24447
R68885 VSS.n9150 VSS.n9128 2.24447
R68886 VSS.n9155 VSS.n964 2.24447
R68887 VSS.n9150 VSS.n9131 2.24447
R68888 VSS.n9155 VSS.n965 2.24447
R68889 VSS.n9150 VSS.n9134 2.24447
R68890 VSS.n9155 VSS.n966 2.24447
R68891 VSS.n9150 VSS.n9137 2.24447
R68892 VSS.n9155 VSS.n967 2.24447
R68893 VSS.n9150 VSS.n9140 2.24447
R68894 VSS.n9155 VSS.n968 2.24447
R68895 VSS.n9150 VSS.n9143 2.24447
R68896 VSS.n9155 VSS.n969 2.24447
R68897 VSS.n9150 VSS.n9146 2.24447
R68898 VSS.n9155 VSS.n970 2.24447
R68899 VSS.n9150 VSS.n9149 2.24447
R68900 VSS.n9155 VSS.n971 2.24447
R68901 VSS.n9152 VSS.n9150 2.24447
R68902 VSS.n9155 VSS.n972 2.24447
R68903 VSS.n9155 VSS.n9154 2.24447
R68904 VSS.n9223 VSS.n903 2.24447
R68905 VSS.n9218 VSS.n9208 2.24447
R68906 VSS.n9223 VSS.n904 2.24447
R68907 VSS.n9218 VSS.n9209 2.24447
R68908 VSS.n9223 VSS.n905 2.24447
R68909 VSS.n9218 VSS.n9210 2.24447
R68910 VSS.n9223 VSS.n906 2.24447
R68911 VSS.n9218 VSS.n9211 2.24447
R68912 VSS.n9223 VSS.n907 2.24447
R68913 VSS.n9218 VSS.n9212 2.24447
R68914 VSS.n9223 VSS.n908 2.24447
R68915 VSS.n9218 VSS.n9213 2.24447
R68916 VSS.n9223 VSS.n909 2.24447
R68917 VSS.n9218 VSS.n9214 2.24447
R68918 VSS.n9223 VSS.n910 2.24447
R68919 VSS.n9218 VSS.n9215 2.24447
R68920 VSS.n9223 VSS.n911 2.24447
R68921 VSS.n9218 VSS.n9216 2.24447
R68922 VSS.n9223 VSS.n912 2.24447
R68923 VSS.n9218 VSS.n9217 2.24447
R68924 VSS.n9223 VSS.n913 2.24447
R68925 VSS.n9219 VSS.n9218 2.24447
R68926 VSS.n9218 VSS.n914 2.24447
R68927 VSS.n4437 VSS.n4435 2.24447
R68928 VSS.n4437 VSS.n4436 2.24447
R68929 VSS.n5171 VSS.n4451 2.24447
R68930 VSS.n5171 VSS.n5170 2.24447
R68931 VSS.n5900 VSS.n4071 2.24447
R68932 VSS.n5904 VSS.n5902 2.24447
R68933 VSS.n6077 VSS.n6076 2.24447
R68934 VSS.n5955 VSS.n5903 2.24447
R68935 VSS.n6037 VSS.n4071 2.24447
R68936 VSS.n5954 VSS.n5904 2.24447
R68937 VSS.n6080 VSS.n6079 2.24447
R68938 VSS.n5957 VSS.n5908 2.24447
R68939 VSS.n3719 VSS.n3717 2.24447
R68940 VSS.n3708 VSS.n3705 2.24447
R68941 VSS.n6303 VSS.n6302 2.24447
R68942 VSS.n6315 VSS.n6314 2.24447
R68943 VSS.n3799 VSS.n3717 2.24447
R68944 VSS.n3710 VSS.n3705 2.24447
R68945 VSS.n6306 VSS.n6305 2.24447
R68946 VSS.n6317 VSS.n3706 2.24447
R68947 VSS.n3194 VSS.n3192 2.24447
R68948 VSS.n3130 VSS.n3127 2.24447
R68949 VSS.n6603 VSS.n6602 2.24447
R68950 VSS.n6621 VSS.n6620 2.24447
R68951 VSS.n3196 VSS.n3192 2.24447
R68952 VSS.n3132 VSS.n3127 2.24447
R68953 VSS.n6606 VSS.n6605 2.24447
R68954 VSS.n6623 VSS.n3128 2.24447
R68955 VSS.n5737 VSS.n5734 2.24447
R68956 VSS.n2960 VSS.n2958 2.24447
R68957 VSS.n5889 VSS.n5888 2.24447
R68958 VSS.n6763 VSS.n2959 2.24447
R68959 VSS.n5739 VSS.n5734 2.24447
R68960 VSS.n6762 VSS.n2960 2.24447
R68961 VSS.n5891 VSS.n5735 2.24447
R68962 VSS.n6765 VSS.n2961 2.24447
R68963 VSS.n2657 VSS.n2655 2.24447
R68964 VSS.n2646 VSS.n2643 2.24447
R68965 VSS.n6995 VSS.n6994 2.24447
R68966 VSS.n7007 VSS.n7006 2.24447
R68967 VSS.n2740 VSS.n2655 2.24447
R68968 VSS.n2648 VSS.n2643 2.24447
R68969 VSS.n6998 VSS.n6997 2.24447
R68970 VSS.n7009 VSS.n2644 2.24447
R68971 VSS.n2353 VSS.n2350 2.24447
R68972 VSS.n9447 VSS.n764 2.24447
R68973 VSS.n2356 VSS.n2355 2.24447
R68974 VSS.n9451 VSS.n765 2.24447
R68975 VSS.n2351 VSS.n2350 2.24447
R68976 VSS.n767 VSS.n764 2.24447
R68977 VSS.n2443 VSS.n2442 2.24447
R68978 VSS.n2449 VSS.n2448 2.24447
R68979 VSS.n2440 VSS.n2429 2.24447
R68980 VSS.n2465 VSS.n2464 2.24447
R68981 VSS.n7154 VSS.n7153 2.24423
R68982 VSS.n2570 VSS.n2568 2.24423
R68983 VSS.n7156 VSS.n2565 2.24423
R68984 VSS.n7145 VSS.n2571 2.24423
R68985 VSS.n7133 VSS.n2576 2.24423
R68986 VSS.n7136 VSS.n2575 2.24423
R68987 VSS.n2783 VSS.n2777 2.24423
R68988 VSS.n2584 VSS.n2580 2.24423
R68989 VSS.n7127 VSS.n2579 2.24423
R68990 VSS.n2787 VSS.n2780 2.24423
R68991 VSS.n2792 VSS.n2776 2.24423
R68992 VSS.n2791 VSS.n2774 2.24423
R68993 VSS.n4638 VSS.n4637 2.24423
R68994 VSS.n4673 VSS.n4672 2.24423
R68995 VSS.n4672 VSS.n4643 2.24423
R68996 VSS.n4669 VSS.n4668 2.24423
R68997 VSS.n4668 VSS.n4647 2.24423
R68998 VSS.n4665 VSS.n4664 2.24423
R68999 VSS.n4664 VSS.n4653 2.24423
R69000 VSS.n4661 VSS.n4660 2.24423
R69001 VSS.n17 VSS.n13 2.24423
R69002 VSS.n9894 VSS.n21 2.24423
R69003 VSS.n9894 VSS.n31 2.24423
R69004 VSS.n161 VSS.n160 2.24423
R69005 VSS.n161 VSS.n156 2.24423
R69006 VSS.n4634 VSS.n4604 2.24423
R69007 VSS.n4675 VSS.n4633 2.24423
R69008 VSS.n4675 VSS.n4632 2.24423
R69009 VSS.n4645 VSS.n4355 2.24423
R69010 VSS.n4649 VSS.n4355 2.24423
R69011 VSS.n4651 VSS.n4395 2.24423
R69012 VSS.n4655 VSS.n4395 2.24423
R69013 VSS.n4656 VSS.n4438 2.24423
R69014 VSS.n4657 VSS.n4438 2.24423
R69015 VSS.n4452 VSS.n12 2.24423
R69016 VSS.n4452 VSS.n19 2.24423
R69017 VSS.n26 VSS.n20 2.24423
R69018 VSS.n28 VSS.n20 2.24423
R69019 VSS.n158 VSS.n83 2.24423
R69020 VSS.n154 VSS.n83 2.24423
R69021 VSS.n9821 VSS.n147 2.24423
R69022 VSS.n9819 VSS.n141 2.24423
R69023 VSS.n9573 VSS.n9572 2.24423
R69024 VSS.n538 VSS.n537 2.24423
R69025 VSS.n2617 VSS.n2614 2.24423
R69026 VSS.n7047 VSS.n2610 2.24423
R69027 VSS.n7041 VSS.n7035 2.24423
R69028 VSS.n7037 VSS.n7032 2.24423
R69029 VSS.n165 VSS.n164 2.24423
R69030 VSS.n165 VSS.n150 2.24423
R69031 VSS.n152 VSS.n114 2.24423
R69032 VSS.n148 VSS.n114 2.24423
R69033 VSS.n7039 VSS.n2618 2.24423
R69034 VSS.n7101 VSS.n7056 2.24011
R69035 VSS.n7075 VSS.n2599 2.24011
R69036 VSS.n7162 VSS.n2555 2.24011
R69037 VSS.n7262 VSS.n2482 2.24011
R69038 VSS.n7247 VSS.n7246 2.24011
R69039 VSS.n8584 VSS.n8577 2.24011
R69040 VSS.n8584 VSS.n8583 2.24011
R69041 VSS.n8590 VSS.n8575 2.24011
R69042 VSS.n8590 VSS.n8589 2.24011
R69043 VSS.n8593 VSS.n8573 2.24011
R69044 VSS.n8595 VSS.n8573 2.24011
R69045 VSS.n8604 VSS.n1548 2.24011
R69046 VSS.n8605 VSS.n8604 2.24011
R69047 VSS.n8086 VSS.n8082 2.24011
R69048 VSS.n8086 VSS.n8081 2.24011
R69049 VSS.n7052 VSS.n7051 2.24011
R69050 VSS.n7106 VSS.n7105 2.24011
R69051 VSS.n7121 VSS.n7120 2.24011
R69052 VSS.n7124 VSS.n7123 2.24011
R69053 VSS.n7113 VSS.n2593 2.24011
R69054 VSS.n8599 VSS.n1550 2.24011
R69055 VSS.n8601 VSS.n1550 2.24011
R69056 VSS.n7099 VSS.n7098 2.24011
R69057 VSS.n7099 VSS.n7097 2.24011
R69058 VSS.n2560 VSS.n2557 2.24011
R69059 VSS.n7160 VSS.n7159 2.24011
R69060 VSS.n7260 VSS.n2480 2.24011
R69061 VSS.n7243 VSS.n2503 2.24011
R69062 VSS.n8607 VSS.n1546 2.24011
R69063 VSS.n8607 VSS.n1545 2.24011
R69064 VSS.n8594 VSS.n8572 2.24011
R69065 VSS.n8587 VSS.n8574 2.24011
R69066 VSS.n8588 VSS.n8587 2.24011
R69067 VSS.n8581 VSS.n8576 2.24011
R69068 VSS.n8582 VSS.n8581 2.24011
R69069 VSS.n8084 VSS.n8079 2.24011
R69070 VSS.n7126 VSS.n2588 2.24011
R69071 VSS.n2591 VSS.n2505 2.24011
R69072 VSS.n7110 VSS.n7109 2.24011
R69073 VSS.n7102 VSS.n2602 2.24011
R69074 VSS.n7048 VSS.n2604 2.24011
R69075 VSS.n8600 VSS.n1549 2.24011
R69076 VSS.n7267 VSS.n2474 2.24011
R69077 VSS.n7071 VSS.n7070 2.24011
R69078 VSS.n6219 VSS.n6218 2.23714
R69079 VSS.n6221 VSS.n3884 2.23714
R69080 VSS.n6218 VSS.n3892 2.23714
R69081 VSS.n6221 VSS.n3883 2.23714
R69082 VSS.n6218 VSS.n3891 2.23714
R69083 VSS.n6221 VSS.n3882 2.23714
R69084 VSS.n6213 VSS.n3894 2.23714
R69085 VSS.n6215 VSS.n3900 2.23714
R69086 VSS.n6213 VSS.n3907 2.23714
R69087 VSS.n6215 VSS.n3899 2.23714
R69088 VSS.n6213 VSS.n3906 2.23714
R69089 VSS.n6059 VSS.n6058 2.23714
R69090 VSS.n6062 VSS.n6055 2.23714
R69091 VSS.n6060 VSS.n6059 2.23714
R69092 VSS.n6285 VSS.n6284 2.23714
R69093 VSS.n6288 VSS.n3819 2.23714
R69094 VSS.n6286 VSS.n6285 2.23714
R69095 VSS.n5731 VSS.n3830 2.18432
R69096 VSS.n5731 VSS.n3827 2.18432
R69097 VSS.n5896 VSS.n434 2.18432
R69098 VSS.n5896 VSS.n443 2.18432
R69099 VSS.n6056 VSS.n3821 1.5539
R69100 VSS.n6214 VSS.n3905 1.53005
R69101 VSS.n4571 VSS.n4570 1.52689
R69102 VSS.n9431 VSS.n709 1.5005
R69103 VSS.n9430 VSS.n9429 1.5005
R69104 VSS.n9428 VSS.n9427 1.5005
R69105 VSS.n9426 VSS.n9425 1.5005
R69106 VSS.n9424 VSS.n9423 1.5005
R69107 VSS.n9422 VSS.n9421 1.5005
R69108 VSS.n9420 VSS.n9419 1.5005
R69109 VSS.n9418 VSS.n9417 1.5005
R69110 VSS.n9416 VSS.n9415 1.5005
R69111 VSS.n9414 VSS.n9413 1.5005
R69112 VSS.n9412 VSS.n9411 1.5005
R69113 VSS.n9410 VSS.n9409 1.5005
R69114 VSS.n9408 VSS.n9407 1.5005
R69115 VSS.n9406 VSS.n9405 1.5005
R69116 VSS.n9404 VSS.n9403 1.5005
R69117 VSS.n9402 VSS.n9401 1.5005
R69118 VSS.n9400 VSS.n9399 1.5005
R69119 VSS.n9398 VSS.n9397 1.5005
R69120 VSS.n9396 VSS.n9395 1.5005
R69121 VSS.n9394 VSS.n9393 1.5005
R69122 VSS.n9392 VSS.n9391 1.5005
R69123 VSS.n9390 VSS.n9389 1.5005
R69124 VSS.n9388 VSS.n9387 1.5005
R69125 VSS.n9386 VSS.n9385 1.5005
R69126 VSS.n9384 VSS.n9383 1.5005
R69127 VSS.n9382 VSS.n9381 1.5005
R69128 VSS.n9380 VSS.n9379 1.5005
R69129 VSS.n759 VSS.n758 1.5005
R69130 VSS.n9456 VSS.n756 1.5005
R69131 VSS.n9458 VSS.n9457 1.5005
R69132 VSS.n757 VSS.n754 1.5005
R69133 VSS.n1170 VSS.n1169 1.5005
R69134 VSS.n1172 VSS.n1171 1.5005
R69135 VSS.n1174 VSS.n1173 1.5005
R69136 VSS.n1176 VSS.n1175 1.5005
R69137 VSS.n1178 VSS.n1177 1.5005
R69138 VSS.n1180 VSS.n1179 1.5005
R69139 VSS.n1182 VSS.n1181 1.5005
R69140 VSS.n1184 VSS.n1183 1.5005
R69141 VSS.n1186 VSS.n1185 1.5005
R69142 VSS.n1188 VSS.n1187 1.5005
R69143 VSS.n1190 VSS.n1189 1.5005
R69144 VSS.n1192 VSS.n1191 1.5005
R69145 VSS.n1194 VSS.n1193 1.5005
R69146 VSS.n1196 VSS.n1195 1.5005
R69147 VSS.n1198 VSS.n1197 1.5005
R69148 VSS.n1200 VSS.n1199 1.5005
R69149 VSS.n1202 VSS.n1201 1.5005
R69150 VSS.n1204 VSS.n1203 1.5005
R69151 VSS.n1206 VSS.n1205 1.5005
R69152 VSS.n1208 VSS.n1207 1.5005
R69153 VSS.n1210 VSS.n1209 1.5005
R69154 VSS.n1212 VSS.n1211 1.5005
R69155 VSS.n1214 VSS.n1213 1.5005
R69156 VSS.n1216 VSS.n1215 1.5005
R69157 VSS.n1218 VSS.n1217 1.5005
R69158 VSS.n2372 VSS.n1863 1.5005
R69159 VSS.n2374 VSS.n2373 1.5005
R69160 VSS.n2376 VSS.n2375 1.5005
R69161 VSS.n2378 VSS.n2377 1.5005
R69162 VSS.n2380 VSS.n2379 1.5005
R69163 VSS.n2382 VSS.n2381 1.5005
R69164 VSS.n2384 VSS.n2383 1.5005
R69165 VSS.n2386 VSS.n2385 1.5005
R69166 VSS.n2388 VSS.n2387 1.5005
R69167 VSS.n2390 VSS.n2389 1.5005
R69168 VSS.n2392 VSS.n2391 1.5005
R69169 VSS.n2394 VSS.n2393 1.5005
R69170 VSS.n2396 VSS.n2395 1.5005
R69171 VSS.n2398 VSS.n2397 1.5005
R69172 VSS.n2400 VSS.n2399 1.5005
R69173 VSS.n2402 VSS.n2401 1.5005
R69174 VSS.n2404 VSS.n2403 1.5005
R69175 VSS.n2406 VSS.n2405 1.5005
R69176 VSS.n2408 VSS.n2407 1.5005
R69177 VSS.n2410 VSS.n2409 1.5005
R69178 VSS.n2412 VSS.n2411 1.5005
R69179 VSS.n2414 VSS.n2413 1.5005
R69180 VSS.n2416 VSS.n2415 1.5005
R69181 VSS.n2418 VSS.n2417 1.5005
R69182 VSS.n2420 VSS.n2419 1.5005
R69183 VSS.n2422 VSS.n2421 1.5005
R69184 VSS.n2424 VSS.n2423 1.5005
R69185 VSS.n2426 VSS.n2425 1.5005
R69186 VSS.n7890 VSS.n2169 1.5005
R69187 VSS.n7892 VSS.n7891 1.5005
R69188 VSS.n2329 VSS.n2166 1.5005
R69189 VSS.n2328 VSS.n2327 1.5005
R69190 VSS.n2326 VSS.n2325 1.5005
R69191 VSS.n2324 VSS.n2323 1.5005
R69192 VSS.n2322 VSS.n2321 1.5005
R69193 VSS.n2320 VSS.n2319 1.5005
R69194 VSS.n2318 VSS.n2317 1.5005
R69195 VSS.n2316 VSS.n2315 1.5005
R69196 VSS.n2314 VSS.n2313 1.5005
R69197 VSS.n2312 VSS.n2311 1.5005
R69198 VSS.n2310 VSS.n2309 1.5005
R69199 VSS.n2308 VSS.n2307 1.5005
R69200 VSS.n2306 VSS.n2305 1.5005
R69201 VSS.n2304 VSS.n2303 1.5005
R69202 VSS.n2302 VSS.n2301 1.5005
R69203 VSS.n2300 VSS.n2299 1.5005
R69204 VSS.n2298 VSS.n2297 1.5005
R69205 VSS.n2296 VSS.n2295 1.5005
R69206 VSS.n2294 VSS.n2293 1.5005
R69207 VSS.n2292 VSS.n2291 1.5005
R69208 VSS.n2290 VSS.n2289 1.5005
R69209 VSS.n2288 VSS.n2287 1.5005
R69210 VSS.n2286 VSS.n2285 1.5005
R69211 VSS.n2284 VSS.n2283 1.5005
R69212 VSS.n2282 VSS.n2281 1.5005
R69213 VSS.n2280 VSS.n2279 1.5005
R69214 VSS.n7148 VSS.n7147 1.49571
R69215 VSS.n7205 VSS.n2496 1.35477
R69216 VSS.n2524 VSS.n2521 1.35477
R69217 VSS.n1614 VSS.n1553 1.35477
R69218 VSS.n1356 VSS.n1354 1.35477
R69219 VSS.n2787 VSS.n1687 1.3133
R69220 VSS.n2791 VSS.n1707 1.3133
R69221 VSS.n9573 VSS.n9570 1.3133
R69222 VSS.n7039 VSS.n1269 1.3133
R69223 VSS.n7048 VSS.n7047 1.17883
R69224 VSS.n7127 VSS.n7126 1.17883
R69225 VSS.n6217 VSS.n6216 0.8825
R69226 VSS.n7249 VSS.n7248 0.754554
R69227 VSS.n7088 VSS.n7057 0.754554
R69228 VSS.n2554 VSS.n2553 0.754554
R69229 VSS.n7253 VSS.n2493 0.754554
R69230 VSS.n7068 VSS.n2506 0.751716
R69231 VSS.n7078 VSS.n7058 0.751716
R69232 VSS.n7264 VSS.n7263 0.751716
R69233 VSS.n7161 VSS.n2563 0.751716
R69234 VSS.n8603 VSS.n8602 0.751716
R69235 VSS.n8592 VSS.n8591 0.751716
R69236 VSS.n7117 VSS.n7116 0.751716
R69237 VSS.n7108 VSS.n7107 0.751716
R69238 VSS.n8606 VSS.n1547 0.746446
R69239 VSS.n8586 VSS.n8585 0.746446
R69240 VSS.n7125 VSS.n7122 0.746446
R69241 VSS.n7054 VSS.n7053 0.746446
R69242 VSS.n7088 VSS.n2520 0.743357
R69243 VSS.n7227 VSS.n2520 0.743357
R69244 VSS.n7190 VSS.n2498 0.743357
R69245 VSS.n7251 VSS.n2498 0.743357
R69246 VSS.n7250 VSS.n7249 0.743357
R69247 VSS.n7251 VSS.n7250 0.743357
R69248 VSS.n7228 VSS.n2522 0.743357
R69249 VSS.n7228 VSS.n7227 0.743357
R69250 VSS.n2497 VSS.n2492 0.743357
R69251 VSS.n7251 VSS.n2497 0.743357
R69252 VSS.n2553 VSS.n2523 0.743357
R69253 VSS.n7227 VSS.n2523 0.743357
R69254 VSS.n7226 VSS.n7225 0.743357
R69255 VSS.n7227 VSS.n7226 0.743357
R69256 VSS.n7253 VSS.n7252 0.743357
R69257 VSS.n7252 VSS.n7251 0.743357
R69258 VSS.n9907 VSS.n9906 0.682336
R69259 VSS.n9905 VSS.n6 0.682336
R69260 VSS.n7302 VSS.n7 0.682078
R69261 VSS.n7879 VSS.n7878 0.682078
R69262 VSS.n536 DVSS 0.66425
R69263 VSS.n5780 DVSS 0.66425
R69264 VSS.n494 DVSS 0.66425
R69265 VSS.n6283 DVSS 0.66425
R69266 VSS.n437 DVSS 0.66425
R69267 VSS.n4092 DVSS 0.66425
R69268 VSS.n4158 DVSS 0.66425
R69269 VSS.n4756 DVSS 0.66425
R69270 VSS.n175 DVSS 0.66425
R69271 VSS.n2789 DVSS 0.66425
R69272 VSS.n3864 DVSS 0.66425
R69273 VSS.n5465 DVSS 0.66425
R69274 VSS.n6057 DVSS 0.66425
R69275 VSS.n428 DVSS 0.66425
R69276 VSS.n6582 DVSS 0.66425
R69277 VSS.n485 DVSS 0.66425
R69278 VSS.n6974 DVSS 0.66425
R69279 VSS.n527 DVSS 0.66425
R69280 VSS.n4730 VSS.n3859 0.623413
R69281 VSS.n6275 VSS.n6274 0.623413
R69282 VSS.n6580 VSS.n3229 0.623413
R69283 VSS.n9813 VSS.n174 0.623413
R69284 VSS.n9602 VSS.n9601 0.623413
R69285 VSS.n9589 VSS.n9588 0.623413
R69286 VSS.n6972 VSS.n2773 0.616858
R69287 VSS.n9576 VSS.n9575 0.616858
R69288 VSS.n5446 VSS.n219 0.612075
R69289 VSS.n5939 VSS.n3688 0.612075
R69290 VSS.n6640 VSS.n6639 0.612075
R69291 VSS.n5759 VSS.n3219 0.612075
R69292 VSS.n9688 VSS.n9687 0.612075
R69293 VSS.n5947 VSS.n3697 0.612075
R69294 VSS.n6758 VSS.n2966 0.612075
R69295 VSS.n4515 VSS.n4280 0.612075
R69296 VSS.n6041 VSS.n3801 0.612075
R69297 VSS.n5741 VSS.n3201 0.612075
R69298 VSS.n5253 VSS.n5252 0.612075
R69299 VSS.n6049 VSS.n3810 0.612075
R69300 VSS.n5750 VSS.n3210 0.612075
R69301 VSS.n5441 VSS.n205 0.612075
R69302 VSS.n5932 VSS.n3684 0.612075
R69303 VSS.n3659 VSS.n3109 0.612075
R69304 VSS.n2629 VSS.n2617 0.611189
R69305 VSS.n2783 VSS.n2763 0.611189
R69306 VSS.n2638 VSS.n2570 0.611189
R69307 VSS.n2745 VSS.n2576 0.611189
R69308 VSS.n2754 VSS.n2580 0.611189
R69309 VSS.n7032 VSS.n7031 0.611189
R69310 VSS.n6265 VSS.n6264 0.608354
R69311 VSS.n9607 VSS.n9606 0.608354
R69312 VSS.n9645 VSS.n359 0.602685
R69313 VSS.n9679 VSS.n325 0.602685
R69314 VSS.n6160 VSS.n3996 0.602685
R69315 VSS.n6196 VSS.n3952 0.602685
R69316 VSS.n9627 VSS.n397 0.602685
R69317 VSS.n4720 VSS.n4590 0.513801
R69318 VSS.n9825 VSS.n146 0.513519
R69319 VSS.n9828 VSS.n9824 0.5005
R69320 VSS.n4716 VSS.n4608 0.5005
R69321 VSS.n4715 VSS.n4609 0.5005
R69322 VSS.n4713 VSS.n4610 0.5005
R69323 VSS.n4613 VSS.n4611 0.5005
R69324 VSS.n4709 VSS.n4614 0.5005
R69325 VSS.n4708 VSS.n4615 0.5005
R69326 VSS.n4707 VSS.n4616 0.5005
R69327 VSS.n4681 VSS.n4617 0.5005
R69328 VSS.n4701 VSS.n4682 0.5005
R69329 VSS.n4700 VSS.n4683 0.5005
R69330 VSS.n4698 VSS.n4684 0.5005
R69331 VSS.n4687 VSS.n4685 0.5005
R69332 VSS.n4694 VSS.n4688 0.5005
R69333 VSS.n4693 VSS.n4689 0.5005
R69334 VSS.n4692 VSS.n4691 0.5005
R69335 VSS.n4690 VSS.n4358 0.5005
R69336 VSS.n5229 VSS.n4359 0.5005
R69337 VSS.n5228 VSS.n4360 0.5005
R69338 VSS.n5226 VSS.n4361 0.5005
R69339 VSS.n4364 VSS.n4362 0.5005
R69340 VSS.n5222 VSS.n4365 0.5005
R69341 VSS.n5221 VSS.n4366 0.5005
R69342 VSS.n5220 VSS.n4367 0.5005
R69343 VSS.n4370 VSS.n4368 0.5005
R69344 VSS.n5216 VSS.n4371 0.5005
R69345 VSS.n5215 VSS.n4372 0.5005
R69346 VSS.n5214 VSS.n4373 0.5005
R69347 VSS.n4376 VSS.n4374 0.5005
R69348 VSS.n5210 VSS.n4377 0.5005
R69349 VSS.n5209 VSS.n4378 0.5005
R69350 VSS.n5208 VSS.n4379 0.5005
R69351 VSS.n4401 VSS.n4380 0.5005
R69352 VSS.n5202 VSS.n4402 0.5005
R69353 VSS.n5201 VSS.n4403 0.5005
R69354 VSS.n5199 VSS.n4404 0.5005
R69355 VSS.n4407 VSS.n4405 0.5005
R69356 VSS.n5195 VSS.n4408 0.5005
R69357 VSS.n5194 VSS.n4409 0.5005
R69358 VSS.n5193 VSS.n4410 0.5005
R69359 VSS.n4413 VSS.n4411 0.5005
R69360 VSS.n5189 VSS.n4414 0.5005
R69361 VSS.n5188 VSS.n4415 0.5005
R69362 VSS.n5187 VSS.n4416 0.5005
R69363 VSS.n4419 VSS.n4417 0.5005
R69364 VSS.n5183 VSS.n4420 0.5005
R69365 VSS.n5182 VSS.n4421 0.5005
R69366 VSS.n5181 VSS.n4422 0.5005
R69367 VSS.n4442 VSS.n4423 0.5005
R69368 VSS.n4443 VSS.n4441 0.5005
R69369 VSS.n5175 VSS.n4444 0.5005
R69370 VSS.n5174 VSS.n4445 0.5005
R69371 VSS.n5173 VSS.n4446 0.5005
R69372 VSS.n5128 VSS.n4447 0.5005
R69373 VSS.n5165 VSS.n5129 0.5005
R69374 VSS.n5164 VSS.n5130 0.5005
R69375 VSS.n5163 VSS.n5131 0.5005
R69376 VSS.n5134 VSS.n5132 0.5005
R69377 VSS.n5159 VSS.n5135 0.5005
R69378 VSS.n5158 VSS.n5136 0.5005
R69379 VSS.n5157 VSS.n5137 0.5005
R69380 VSS.n5140 VSS.n5138 0.5005
R69381 VSS.n5153 VSS.n5141 0.5005
R69382 VSS.n5152 VSS.n5142 0.5005
R69383 VSS.n5151 VSS.n5143 0.5005
R69384 VSS.n5148 VSS.n5144 0.5005
R69385 VSS.n5147 VSS.n5146 0.5005
R69386 VSS.n5145 VSS.n46 0.5005
R69387 VSS.n9887 VSS.n47 0.5005
R69388 VSS.n9886 VSS.n48 0.5005
R69389 VSS.n9884 VSS.n49 0.5005
R69390 VSS.n52 VSS.n50 0.5005
R69391 VSS.n9880 VSS.n53 0.5005
R69392 VSS.n9879 VSS.n54 0.5005
R69393 VSS.n9878 VSS.n55 0.5005
R69394 VSS.n58 VSS.n56 0.5005
R69395 VSS.n9874 VSS.n59 0.5005
R69396 VSS.n9873 VSS.n60 0.5005
R69397 VSS.n9872 VSS.n61 0.5005
R69398 VSS.n64 VSS.n62 0.5005
R69399 VSS.n9868 VSS.n65 0.5005
R69400 VSS.n9867 VSS.n66 0.5005
R69401 VSS.n9866 VSS.n67 0.5005
R69402 VSS.n89 VSS.n68 0.5005
R69403 VSS.n9860 VSS.n90 0.5005
R69404 VSS.n9859 VSS.n91 0.5005
R69405 VSS.n9857 VSS.n92 0.5005
R69406 VSS.n95 VSS.n93 0.5005
R69407 VSS.n9853 VSS.n96 0.5005
R69408 VSS.n9852 VSS.n97 0.5005
R69409 VSS.n9851 VSS.n98 0.5005
R69410 VSS.n120 VSS.n99 0.5005
R69411 VSS.n9845 VSS.n121 0.5005
R69412 VSS.n9844 VSS.n122 0.5005
R69413 VSS.n9842 VSS.n123 0.5005
R69414 VSS.n126 VSS.n124 0.5005
R69415 VSS.n9838 VSS.n127 0.5005
R69416 VSS.n9837 VSS.n128 0.5005
R69417 VSS.n9836 VSS.n129 0.5005
R69418 VSS.n9823 VSS.n130 0.5005
R69419 VSS.n9827 VSS.n9826 0.5005
R69420 VSS.n9829 VSS.n9828 0.5005
R69421 VSS.n4607 VSS.n4595 0.5005
R69422 VSS.n4717 VSS.n4716 0.5005
R69423 VSS.n4715 VSS.n4714 0.5005
R69424 VSS.n4713 VSS.n4712 0.5005
R69425 VSS.n4711 VSS.n4611 0.5005
R69426 VSS.n4710 VSS.n4709 0.5005
R69427 VSS.n4708 VSS.n4612 0.5005
R69428 VSS.n4707 VSS.n4706 0.5005
R69429 VSS.n4623 VSS.n4617 0.5005
R69430 VSS.n4702 VSS.n4701 0.5005
R69431 VSS.n4700 VSS.n4699 0.5005
R69432 VSS.n4698 VSS.n4697 0.5005
R69433 VSS.n4696 VSS.n4685 0.5005
R69434 VSS.n4695 VSS.n4694 0.5005
R69435 VSS.n4693 VSS.n4686 0.5005
R69436 VSS.n4692 VSS.n4341 0.5005
R69437 VSS.n4358 VSS.n4346 0.5005
R69438 VSS.n5230 VSS.n5229 0.5005
R69439 VSS.n5228 VSS.n5227 0.5005
R69440 VSS.n5226 VSS.n5225 0.5005
R69441 VSS.n5224 VSS.n4362 0.5005
R69442 VSS.n5223 VSS.n5222 0.5005
R69443 VSS.n5221 VSS.n4363 0.5005
R69444 VSS.n5220 VSS.n5219 0.5005
R69445 VSS.n5218 VSS.n4368 0.5005
R69446 VSS.n5217 VSS.n5216 0.5005
R69447 VSS.n5215 VSS.n4369 0.5005
R69448 VSS.n5214 VSS.n5213 0.5005
R69449 VSS.n5212 VSS.n4374 0.5005
R69450 VSS.n5211 VSS.n5210 0.5005
R69451 VSS.n5209 VSS.n4375 0.5005
R69452 VSS.n5208 VSS.n5207 0.5005
R69453 VSS.n4386 VSS.n4380 0.5005
R69454 VSS.n5203 VSS.n5202 0.5005
R69455 VSS.n5201 VSS.n5200 0.5005
R69456 VSS.n5199 VSS.n5198 0.5005
R69457 VSS.n5197 VSS.n4405 0.5005
R69458 VSS.n5196 VSS.n5195 0.5005
R69459 VSS.n5194 VSS.n4406 0.5005
R69460 VSS.n5193 VSS.n5192 0.5005
R69461 VSS.n5191 VSS.n4411 0.5005
R69462 VSS.n5190 VSS.n5189 0.5005
R69463 VSS.n5188 VSS.n4412 0.5005
R69464 VSS.n5187 VSS.n5186 0.5005
R69465 VSS.n5185 VSS.n4417 0.5005
R69466 VSS.n5184 VSS.n5183 0.5005
R69467 VSS.n5182 VSS.n4418 0.5005
R69468 VSS.n5181 VSS.n5180 0.5005
R69469 VSS.n4429 VSS.n4423 0.5005
R69470 VSS.n4441 VSS.n4439 0.5005
R69471 VSS.n5176 VSS.n5175 0.5005
R69472 VSS.n5174 VSS.n4440 0.5005
R69473 VSS.n5173 VSS.n5172 0.5005
R69474 VSS.n4454 VSS.n4447 0.5005
R69475 VSS.n5166 VSS.n5165 0.5005
R69476 VSS.n5164 VSS.n5127 0.5005
R69477 VSS.n5163 VSS.n5162 0.5005
R69478 VSS.n5161 VSS.n5132 0.5005
R69479 VSS.n5160 VSS.n5159 0.5005
R69480 VSS.n5158 VSS.n5133 0.5005
R69481 VSS.n5157 VSS.n5156 0.5005
R69482 VSS.n5155 VSS.n5138 0.5005
R69483 VSS.n5154 VSS.n5153 0.5005
R69484 VSS.n5152 VSS.n5139 0.5005
R69485 VSS.n5151 VSS.n5150 0.5005
R69486 VSS.n5149 VSS.n5148 0.5005
R69487 VSS.n5147 VSS.n35 0.5005
R69488 VSS.n46 VSS.n41 0.5005
R69489 VSS.n9888 VSS.n9887 0.5005
R69490 VSS.n9886 VSS.n9885 0.5005
R69491 VSS.n9884 VSS.n9883 0.5005
R69492 VSS.n9882 VSS.n50 0.5005
R69493 VSS.n9881 VSS.n9880 0.5005
R69494 VSS.n9879 VSS.n51 0.5005
R69495 VSS.n9878 VSS.n9877 0.5005
R69496 VSS.n9876 VSS.n56 0.5005
R69497 VSS.n9875 VSS.n9874 0.5005
R69498 VSS.n9873 VSS.n57 0.5005
R69499 VSS.n9872 VSS.n9871 0.5005
R69500 VSS.n9870 VSS.n62 0.5005
R69501 VSS.n9869 VSS.n9868 0.5005
R69502 VSS.n9867 VSS.n63 0.5005
R69503 VSS.n9866 VSS.n9865 0.5005
R69504 VSS.n74 VSS.n68 0.5005
R69505 VSS.n9861 VSS.n9860 0.5005
R69506 VSS.n9859 VSS.n9858 0.5005
R69507 VSS.n9857 VSS.n9856 0.5005
R69508 VSS.n9855 VSS.n93 0.5005
R69509 VSS.n9854 VSS.n9853 0.5005
R69510 VSS.n9852 VSS.n94 0.5005
R69511 VSS.n9851 VSS.n9850 0.5005
R69512 VSS.n105 VSS.n99 0.5005
R69513 VSS.n9846 VSS.n9845 0.5005
R69514 VSS.n9844 VSS.n9843 0.5005
R69515 VSS.n9842 VSS.n9841 0.5005
R69516 VSS.n9840 VSS.n124 0.5005
R69517 VSS.n9839 VSS.n9838 0.5005
R69518 VSS.n9837 VSS.n125 0.5005
R69519 VSS.n9836 VSS.n9835 0.5005
R69520 VSS.n136 VSS.n130 0.5005
R69521 VSS.n4663 VSS.n4662 0.466338
R69522 VSS.n9898 VSS.n9897 0.466338
R69523 VSS.n4667 VSS.n4666 0.46307
R69524 VSS.n9895 VSS.n29 0.46307
R69525 VSS.n8298 VSS.n8281 0.462685
R69526 VSS.n6964 VSS.n2799 0.462685
R69527 VSS.n6263 VSS.n3836 0.462685
R69528 VSS.n6248 VSS.n3869 0.462685
R69529 VSS.n4762 VSS.n4731 0.462685
R69530 VSS.n8884 VSS.n540 0.462428
R69531 VSS.n6673 VSS.n502 0.462428
R69532 VSS.n425 VSS.n404 0.462428
R69533 VSS.n5482 VSS.n5428 0.462428
R69534 VSS.n9793 VSS.n178 0.462428
R69535 VSS.n7302 VSS.n7300 0.455549
R69536 VSS.n7414 VSS.n6 0.455549
R69537 VSS.n7878 VSS.n7272 0.455549
R69538 VSS.n9907 VSS.n3 0.455549
R69539 VSS.n7593 VSS.n7592 0.4505
R69540 VSS.n7591 VSS.n7291 0.4505
R69541 VSS.n7590 VSS.n7589 0.4505
R69542 VSS.n7325 VSS.n7324 0.4505
R69543 VSS.n7585 VSS.n7584 0.4505
R69544 VSS.n7583 VSS.n7327 0.4505
R69545 VSS.n7582 VSS.n7581 0.4505
R69546 VSS.n7329 VSS.n7328 0.4505
R69547 VSS.n7577 VSS.n7576 0.4505
R69548 VSS.n7575 VSS.n7331 0.4505
R69549 VSS.n7574 VSS.n7573 0.4505
R69550 VSS.n7333 VSS.n7332 0.4505
R69551 VSS.n7569 VSS.n7568 0.4505
R69552 VSS.n7567 VSS.n7335 0.4505
R69553 VSS.n7566 VSS.n7565 0.4505
R69554 VSS.n7337 VSS.n7336 0.4505
R69555 VSS.n7561 VSS.n7560 0.4505
R69556 VSS.n7559 VSS.n7339 0.4505
R69557 VSS.n7558 VSS.n7557 0.4505
R69558 VSS.n7341 VSS.n7340 0.4505
R69559 VSS.n7553 VSS.n7552 0.4505
R69560 VSS.n7551 VSS.n7343 0.4505
R69561 VSS.n7550 VSS.n7549 0.4505
R69562 VSS.n7345 VSS.n7344 0.4505
R69563 VSS.n7545 VSS.n7544 0.4505
R69564 VSS.n7543 VSS.n7347 0.4505
R69565 VSS.n7542 VSS.n7541 0.4505
R69566 VSS.n7349 VSS.n7348 0.4505
R69567 VSS.n7537 VSS.n7536 0.4505
R69568 VSS.n7535 VSS.n7351 0.4505
R69569 VSS.n7534 VSS.n7533 0.4505
R69570 VSS.n7353 VSS.n7352 0.4505
R69571 VSS.n7529 VSS.n7528 0.4505
R69572 VSS.n7527 VSS.n7355 0.4505
R69573 VSS.n7526 VSS.n7525 0.4505
R69574 VSS.n7357 VSS.n7356 0.4505
R69575 VSS.n7521 VSS.n7520 0.4505
R69576 VSS.n7519 VSS.n7359 0.4505
R69577 VSS.n7518 VSS.n7517 0.4505
R69578 VSS.n7361 VSS.n7360 0.4505
R69579 VSS.n7513 VSS.n7512 0.4505
R69580 VSS.n7511 VSS.n7363 0.4505
R69581 VSS.n7510 VSS.n7509 0.4505
R69582 VSS.n7365 VSS.n7364 0.4505
R69583 VSS.n7505 VSS.n7504 0.4505
R69584 VSS.n7503 VSS.n7367 0.4505
R69585 VSS.n7502 VSS.n7501 0.4505
R69586 VSS.n7369 VSS.n7368 0.4505
R69587 VSS.n7497 VSS.n7496 0.4505
R69588 VSS.n7495 VSS.n7371 0.4505
R69589 VSS.n7494 VSS.n7493 0.4505
R69590 VSS.n7373 VSS.n7372 0.4505
R69591 VSS.n7489 VSS.n7488 0.4505
R69592 VSS.n7487 VSS.n7375 0.4505
R69593 VSS.n7486 VSS.n7485 0.4505
R69594 VSS.n7377 VSS.n7376 0.4505
R69595 VSS.n7481 VSS.n7480 0.4505
R69596 VSS.n7479 VSS.n7379 0.4505
R69597 VSS.n7478 VSS.n7477 0.4505
R69598 VSS.n7381 VSS.n7380 0.4505
R69599 VSS.n7473 VSS.n7472 0.4505
R69600 VSS.n7471 VSS.n7383 0.4505
R69601 VSS.n7470 VSS.n7469 0.4505
R69602 VSS.n7385 VSS.n7384 0.4505
R69603 VSS.n7465 VSS.n7464 0.4505
R69604 VSS.n7463 VSS.n7387 0.4505
R69605 VSS.n7462 VSS.n7461 0.4505
R69606 VSS.n7389 VSS.n7388 0.4505
R69607 VSS.n7457 VSS.n7456 0.4505
R69608 VSS.n7455 VSS.n7391 0.4505
R69609 VSS.n7454 VSS.n7453 0.4505
R69610 VSS.n7393 VSS.n7392 0.4505
R69611 VSS.n7449 VSS.n7448 0.4505
R69612 VSS.n7447 VSS.n7395 0.4505
R69613 VSS.n7446 VSS.n7445 0.4505
R69614 VSS.n7397 VSS.n7396 0.4505
R69615 VSS.n7441 VSS.n7440 0.4505
R69616 VSS.n7439 VSS.n7399 0.4505
R69617 VSS.n7438 VSS.n7437 0.4505
R69618 VSS.n7401 VSS.n7400 0.4505
R69619 VSS.n7433 VSS.n7432 0.4505
R69620 VSS.n7431 VSS.n7403 0.4505
R69621 VSS.n7430 VSS.n7429 0.4505
R69622 VSS.n7405 VSS.n7404 0.4505
R69623 VSS.n7425 VSS.n7424 0.4505
R69624 VSS.n7423 VSS.n7407 0.4505
R69625 VSS.n7422 VSS.n7421 0.4505
R69626 VSS.n7418 VSS.n7408 0.4505
R69627 VSS.n7417 VSS.n7416 0.4505
R69628 VSS.n7415 VSS.n7410 0.4505
R69629 VSS.n7306 VSS.n7305 0.4505
R69630 VSS.n7307 VSS.n7299 0.4505
R69631 VSS.n7309 VSS.n7308 0.4505
R69632 VSS.n7297 VSS.n7296 0.4505
R69633 VSS.n7314 VSS.n7313 0.4505
R69634 VSS.n7315 VSS.n7295 0.4505
R69635 VSS.n7317 VSS.n7316 0.4505
R69636 VSS.n7293 VSS.n7292 0.4505
R69637 VSS.n7322 VSS.n7321 0.4505
R69638 VSS.n7323 VSS.n7290 0.4505
R69639 VSS.n9794 VSS.n187 0.4505
R69640 VSS.n4583 VSS.n4582 0.4505
R69641 VSS.n4767 VSS.n4766 0.4505
R69642 VSS.n4768 VSS.n4581 0.4505
R69643 VSS.n4770 VSS.n4769 0.4505
R69644 VSS.n4579 VSS.n4578 0.4505
R69645 VSS.n4775 VSS.n4774 0.4505
R69646 VSS.n4776 VSS.n4577 0.4505
R69647 VSS.n4778 VSS.n4777 0.4505
R69648 VSS.n4551 VSS.n4550 0.4505
R69649 VSS.n4789 VSS.n4788 0.4505
R69650 VSS.n4790 VSS.n4549 0.4505
R69651 VSS.n4792 VSS.n4791 0.4505
R69652 VSS.n4547 VSS.n4546 0.4505
R69653 VSS.n4797 VSS.n4796 0.4505
R69654 VSS.n4798 VSS.n4545 0.4505
R69655 VSS.n4800 VSS.n4799 0.4505
R69656 VSS.n4802 VSS.n4544 0.4505
R69657 VSS.n4805 VSS.n4804 0.4505
R69658 VSS.n4806 VSS.n4543 0.4505
R69659 VSS.n4808 VSS.n4807 0.4505
R69660 VSS.n4541 VSS.n4540 0.4505
R69661 VSS.n4813 VSS.n4812 0.4505
R69662 VSS.n4814 VSS.n4539 0.4505
R69663 VSS.n4816 VSS.n4815 0.4505
R69664 VSS.n4537 VSS.n4536 0.4505
R69665 VSS.n4821 VSS.n4820 0.4505
R69666 VSS.n4822 VSS.n4535 0.4505
R69667 VSS.n4824 VSS.n4823 0.4505
R69668 VSS.n4533 VSS.n4532 0.4505
R69669 VSS.n4829 VSS.n4828 0.4505
R69670 VSS.n4830 VSS.n4529 0.4505
R69671 VSS.n5059 VSS.n5058 0.4505
R69672 VSS.n5057 VSS.n4531 0.4505
R69673 VSS.n5056 VSS.n5055 0.4505
R69674 VSS.n5053 VSS.n4831 0.4505
R69675 VSS.n4835 VSS.n4832 0.4505
R69676 VSS.n5049 VSS.n5048 0.4505
R69677 VSS.n5047 VSS.n4834 0.4505
R69678 VSS.n5046 VSS.n5045 0.4505
R69679 VSS.n4837 VSS.n4836 0.4505
R69680 VSS.n5041 VSS.n5040 0.4505
R69681 VSS.n5039 VSS.n4839 0.4505
R69682 VSS.n5038 VSS.n5037 0.4505
R69683 VSS.n4841 VSS.n4840 0.4505
R69684 VSS.n5033 VSS.n5032 0.4505
R69685 VSS.n5031 VSS.n4843 0.4505
R69686 VSS.n5030 VSS.n5029 0.4505
R69687 VSS.n5028 VSS.n4844 0.4505
R69688 VSS.n5027 VSS.n5025 0.4505
R69689 VSS.n5024 VSS.n4845 0.4505
R69690 VSS.n5023 VSS.n5022 0.4505
R69691 VSS.n4847 VSS.n4846 0.4505
R69692 VSS.n4979 VSS.n4977 0.4505
R69693 VSS.n5016 VSS.n5015 0.4505
R69694 VSS.n5014 VSS.n4978 0.4505
R69695 VSS.n5013 VSS.n5012 0.4505
R69696 VSS.n4981 VSS.n4980 0.4505
R69697 VSS.n5008 VSS.n5007 0.4505
R69698 VSS.n5006 VSS.n4983 0.4505
R69699 VSS.n5005 VSS.n5004 0.4505
R69700 VSS.n4985 VSS.n4984 0.4505
R69701 VSS.n5000 VSS.n4999 0.4505
R69702 VSS.n4998 VSS.n4987 0.4505
R69703 VSS.n4997 VSS.n4996 0.4505
R69704 VSS.n4993 VSS.n4988 0.4505
R69705 VSS.n4992 VSS.n4991 0.4505
R69706 VSS.n4990 VSS.n4989 0.4505
R69707 VSS.n249 VSS.n248 0.4505
R69708 VSS.n9699 VSS.n9698 0.4505
R69709 VSS.n9700 VSS.n247 0.4505
R69710 VSS.n9702 VSS.n9701 0.4505
R69711 VSS.n245 VSS.n244 0.4505
R69712 VSS.n9707 VSS.n9706 0.4505
R69713 VSS.n9708 VSS.n243 0.4505
R69714 VSS.n9710 VSS.n9709 0.4505
R69715 VSS.n241 VSS.n240 0.4505
R69716 VSS.n9715 VSS.n9714 0.4505
R69717 VSS.n9716 VSS.n239 0.4505
R69718 VSS.n9718 VSS.n9717 0.4505
R69719 VSS.n237 VSS.n236 0.4505
R69720 VSS.n9723 VSS.n9722 0.4505
R69721 VSS.n9724 VSS.n233 0.4505
R69722 VSS.n9746 VSS.n9745 0.4505
R69723 VSS.n9744 VSS.n235 0.4505
R69724 VSS.n9743 VSS.n9742 0.4505
R69725 VSS.n9740 VSS.n9725 0.4505
R69726 VSS.n9729 VSS.n9726 0.4505
R69727 VSS.n9736 VSS.n9735 0.4505
R69728 VSS.n9734 VSS.n9728 0.4505
R69729 VSS.n9733 VSS.n9732 0.4505
R69730 VSS.n9731 VSS.n9730 0.4505
R69731 VSS.n193 VSS.n192 0.4505
R69732 VSS.n9781 VSS.n9780 0.4505
R69733 VSS.n9782 VSS.n191 0.4505
R69734 VSS.n9784 VSS.n9783 0.4505
R69735 VSS.n189 VSS.n188 0.4505
R69736 VSS.n9789 VSS.n9788 0.4505
R69737 VSS.n9790 VSS.n185 0.4505
R69738 VSS.n9796 VSS.n9795 0.4505
R69739 VSS.n8889 VSS.n8888 0.4505
R69740 VSS.n1705 VSS.n1704 0.4505
R69741 VSS.n8304 VSS.n8303 0.4505
R69742 VSS.n8305 VSS.n1703 0.4505
R69743 VSS.n8307 VSS.n8306 0.4505
R69744 VSS.n1701 VSS.n1700 0.4505
R69745 VSS.n8312 VSS.n8311 0.4505
R69746 VSS.n8313 VSS.n1699 0.4505
R69747 VSS.n8315 VSS.n8314 0.4505
R69748 VSS.n1685 VSS.n1684 0.4505
R69749 VSS.n8333 VSS.n8332 0.4505
R69750 VSS.n8334 VSS.n1683 0.4505
R69751 VSS.n8336 VSS.n8335 0.4505
R69752 VSS.n1681 VSS.n1680 0.4505
R69753 VSS.n8341 VSS.n8340 0.4505
R69754 VSS.n8342 VSS.n1679 0.4505
R69755 VSS.n8344 VSS.n8343 0.4505
R69756 VSS.n8346 VSS.n1678 0.4505
R69757 VSS.n8349 VSS.n8348 0.4505
R69758 VSS.n8350 VSS.n1677 0.4505
R69759 VSS.n8352 VSS.n8351 0.4505
R69760 VSS.n1675 VSS.n1674 0.4505
R69761 VSS.n8357 VSS.n8356 0.4505
R69762 VSS.n8358 VSS.n1673 0.4505
R69763 VSS.n8360 VSS.n8359 0.4505
R69764 VSS.n1671 VSS.n1670 0.4505
R69765 VSS.n8365 VSS.n8364 0.4505
R69766 VSS.n8366 VSS.n1669 0.4505
R69767 VSS.n8368 VSS.n8367 0.4505
R69768 VSS.n1667 VSS.n1666 0.4505
R69769 VSS.n8374 VSS.n8373 0.4505
R69770 VSS.n8375 VSS.n1665 0.4505
R69771 VSS.n8377 VSS.n8376 0.4505
R69772 VSS.n1654 VSS.n1653 0.4505
R69773 VSS.n8415 VSS.n8414 0.4505
R69774 VSS.n8416 VSS.n1652 0.4505
R69775 VSS.n8418 VSS.n8417 0.4505
R69776 VSS.n1650 VSS.n1649 0.4505
R69777 VSS.n8423 VSS.n8422 0.4505
R69778 VSS.n8424 VSS.n1648 0.4505
R69779 VSS.n8426 VSS.n8425 0.4505
R69780 VSS.n1646 VSS.n1645 0.4505
R69781 VSS.n8431 VSS.n8430 0.4505
R69782 VSS.n8432 VSS.n1644 0.4505
R69783 VSS.n8435 VSS.n8434 0.4505
R69784 VSS.n8433 VSS.n1641 0.4505
R69785 VSS.n8439 VSS.n1642 0.4505
R69786 VSS.n8440 VSS.n1640 0.4505
R69787 VSS.n8442 VSS.n8441 0.4505
R69788 VSS.n8443 VSS.n1638 0.4505
R69789 VSS.n8533 VSS.n8532 0.4505
R69790 VSS.n8531 VSS.n1639 0.4505
R69791 VSS.n8530 VSS.n8529 0.4505
R69792 VSS.n8528 VSS.n8444 0.4505
R69793 VSS.n8527 VSS.n8526 0.4505
R69794 VSS.n8525 VSS.n8445 0.4505
R69795 VSS.n8524 VSS.n8523 0.4505
R69796 VSS.n8447 VSS.n8446 0.4505
R69797 VSS.n8519 VSS.n8518 0.4505
R69798 VSS.n8517 VSS.n8450 0.4505
R69799 VSS.n8516 VSS.n8515 0.4505
R69800 VSS.n8452 VSS.n8451 0.4505
R69801 VSS.n8511 VSS.n8510 0.4505
R69802 VSS.n8509 VSS.n8454 0.4505
R69803 VSS.n8508 VSS.n8507 0.4505
R69804 VSS.n8504 VSS.n8455 0.4505
R69805 VSS.n8503 VSS.n8502 0.4505
R69806 VSS.n8501 VSS.n8456 0.4505
R69807 VSS.n8500 VSS.n8499 0.4505
R69808 VSS.n8497 VSS.n8457 0.4505
R69809 VSS.n8495 VSS.n8459 0.4505
R69810 VSS.n8462 VSS.n8458 0.4505
R69811 VSS.n8491 VSS.n8490 0.4505
R69812 VSS.n8489 VSS.n8461 0.4505
R69813 VSS.n8488 VSS.n8487 0.4505
R69814 VSS.n8464 VSS.n8463 0.4505
R69815 VSS.n8483 VSS.n8482 0.4505
R69816 VSS.n8481 VSS.n8466 0.4505
R69817 VSS.n8480 VSS.n8479 0.4505
R69818 VSS.n8468 VSS.n8467 0.4505
R69819 VSS.n8475 VSS.n8474 0.4505
R69820 VSS.n8473 VSS.n8470 0.4505
R69821 VSS.n8472 VSS.n8471 0.4505
R69822 VSS.n1287 VSS.n1286 0.4505
R69823 VSS.n8864 VSS.n8863 0.4505
R69824 VSS.n8865 VSS.n1285 0.4505
R69825 VSS.n8867 VSS.n8866 0.4505
R69826 VSS.n1283 VSS.n1282 0.4505
R69827 VSS.n8873 VSS.n8872 0.4505
R69828 VSS.n8874 VSS.n1281 0.4505
R69829 VSS.n8876 VSS.n8875 0.4505
R69830 VSS.n8877 VSS.n1280 0.4505
R69831 VSS.n8880 VSS.n8879 0.4505
R69832 VSS.n8881 VSS.n1278 0.4505
R69833 VSS.n8900 VSS.n8899 0.4505
R69834 VSS.n8898 VSS.n1279 0.4505
R69835 VSS.n8897 VSS.n8896 0.4505
R69836 VSS.n8893 VSS.n8882 0.4505
R69837 VSS.n8892 VSS.n8891 0.4505
R69838 VSS.n8890 VSS.n8883 0.4505
R69839 VSS.n8886 VSS.n8885 0.4505
R69840 VSS.n8888 VSS.n8887 0.4505
R69841 VSS.n8287 VSS.n8286 0.4505
R69842 VSS.n8293 VSS.n1705 0.4505
R69843 VSS.n8303 VSS.n8302 0.4505
R69844 VSS.n1703 VSS.n1702 0.4505
R69845 VSS.n8308 VSS.n8307 0.4505
R69846 VSS.n8309 VSS.n1701 0.4505
R69847 VSS.n8311 VSS.n8310 0.4505
R69848 VSS.n1699 VSS.n1694 0.4505
R69849 VSS.n8316 VSS.n8315 0.4505
R69850 VSS.n8322 VSS.n1685 0.4505
R69851 VSS.n8332 VSS.n8331 0.4505
R69852 VSS.n1683 VSS.n1682 0.4505
R69853 VSS.n8337 VSS.n8336 0.4505
R69854 VSS.n8338 VSS.n1681 0.4505
R69855 VSS.n8340 VSS.n8339 0.4505
R69856 VSS.n1679 VSS.n1571 0.4505
R69857 VSS.n8344 VSS.n1578 0.4505
R69858 VSS.n8346 VSS.n8345 0.4505
R69859 VSS.n8348 VSS.n8347 0.4505
R69860 VSS.n1677 VSS.n1676 0.4505
R69861 VSS.n8353 VSS.n8352 0.4505
R69862 VSS.n8354 VSS.n1675 0.4505
R69863 VSS.n8356 VSS.n8355 0.4505
R69864 VSS.n1673 VSS.n1672 0.4505
R69865 VSS.n8361 VSS.n8360 0.4505
R69866 VSS.n8362 VSS.n1671 0.4505
R69867 VSS.n8364 VSS.n8363 0.4505
R69868 VSS.n1669 VSS.n1668 0.4505
R69869 VSS.n8369 VSS.n8368 0.4505
R69870 VSS.n8370 VSS.n1667 0.4505
R69871 VSS.n8373 VSS.n8372 0.4505
R69872 VSS.n8371 VSS.n1665 0.4505
R69873 VSS.n8378 VSS.n8377 0.4505
R69874 VSS.n8384 VSS.n1654 0.4505
R69875 VSS.n8414 VSS.n8413 0.4505
R69876 VSS.n1652 VSS.n1651 0.4505
R69877 VSS.n8419 VSS.n8418 0.4505
R69878 VSS.n8420 VSS.n1650 0.4505
R69879 VSS.n8422 VSS.n8421 0.4505
R69880 VSS.n1648 VSS.n1647 0.4505
R69881 VSS.n8427 VSS.n8426 0.4505
R69882 VSS.n8428 VSS.n1646 0.4505
R69883 VSS.n8430 VSS.n8429 0.4505
R69884 VSS.n1644 VSS.n1643 0.4505
R69885 VSS.n8436 VSS.n8435 0.4505
R69886 VSS.n8437 VSS.n1641 0.4505
R69887 VSS.n8439 VSS.n8438 0.4505
R69888 VSS.n8440 VSS.n1619 0.4505
R69889 VSS.n8441 VSS.n1625 0.4505
R69890 VSS.n1638 VSS.n1634 0.4505
R69891 VSS.n8534 VSS.n8533 0.4505
R69892 VSS.n1639 VSS.n1637 0.4505
R69893 VSS.n8529 VSS.n1378 0.4505
R69894 VSS.n8528 VSS.n1369 0.4505
R69895 VSS.n8527 VSS.n1376 0.4505
R69896 VSS.n8448 VSS.n8445 0.4505
R69897 VSS.n8523 VSS.n8522 0.4505
R69898 VSS.n8521 VSS.n8447 0.4505
R69899 VSS.n8520 VSS.n8519 0.4505
R69900 VSS.n8450 VSS.n8449 0.4505
R69901 VSS.n8515 VSS.n8514 0.4505
R69902 VSS.n8513 VSS.n8452 0.4505
R69903 VSS.n8512 VSS.n8511 0.4505
R69904 VSS.n8454 VSS.n8453 0.4505
R69905 VSS.n8507 VSS.n8506 0.4505
R69906 VSS.n8505 VSS.n8504 0.4505
R69907 VSS.n8503 VSS.n1325 0.4505
R69908 VSS.n8456 VSS.n1331 0.4505
R69909 VSS.n8499 VSS.n8498 0.4505
R69910 VSS.n8497 VSS.n8496 0.4505
R69911 VSS.n8495 VSS.n8494 0.4505
R69912 VSS.n8493 VSS.n8458 0.4505
R69913 VSS.n8492 VSS.n8491 0.4505
R69914 VSS.n8461 VSS.n8460 0.4505
R69915 VSS.n8487 VSS.n8486 0.4505
R69916 VSS.n8485 VSS.n8464 0.4505
R69917 VSS.n8484 VSS.n8483 0.4505
R69918 VSS.n8466 VSS.n8465 0.4505
R69919 VSS.n8479 VSS.n8478 0.4505
R69920 VSS.n8477 VSS.n8468 0.4505
R69921 VSS.n8476 VSS.n8475 0.4505
R69922 VSS.n8470 VSS.n8469 0.4505
R69923 VSS.n8471 VSS.n1306 0.4505
R69924 VSS.n1309 VSS.n1287 0.4505
R69925 VSS.n8863 VSS.n8862 0.4505
R69926 VSS.n1294 VSS.n1285 0.4505
R69927 VSS.n8868 VSS.n8867 0.4505
R69928 VSS.n8869 VSS.n1283 0.4505
R69929 VSS.n8872 VSS.n8871 0.4505
R69930 VSS.n8870 VSS.n1281 0.4505
R69931 VSS.n8876 VSS.n1261 0.4505
R69932 VSS.n8877 VSS.n1267 0.4505
R69933 VSS.n8879 VSS.n8878 0.4505
R69934 VSS.n1278 VSS.n1276 0.4505
R69935 VSS.n8901 VSS.n8900 0.4505
R69936 VSS.n1279 VSS.n1277 0.4505
R69937 VSS.n8896 VSS.n8895 0.4505
R69938 VSS.n8894 VSS.n8893 0.4505
R69939 VSS.n8892 VSS.n542 0.4505
R69940 VSS.n8883 VSS.n548 0.4505
R69941 VSS.n6678 VSS.n6677 0.4505
R69942 VSS.n2821 VSS.n2820 0.4505
R69943 VSS.n2822 VSS.n2816 0.4505
R69944 VSS.n6955 VSS.n6954 0.4505
R69945 VSS.n6953 VSS.n2817 0.4505
R69946 VSS.n6952 VSS.n6951 0.4505
R69947 VSS.n2824 VSS.n2823 0.4505
R69948 VSS.n6947 VSS.n6946 0.4505
R69949 VSS.n6945 VSS.n2826 0.4505
R69950 VSS.n6944 VSS.n6943 0.4505
R69951 VSS.n2828 VSS.n2827 0.4505
R69952 VSS.n6932 VSS.n6931 0.4505
R69953 VSS.n6930 VSS.n2848 0.4505
R69954 VSS.n6929 VSS.n6928 0.4505
R69955 VSS.n2850 VSS.n2849 0.4505
R69956 VSS.n6924 VSS.n6923 0.4505
R69957 VSS.n6922 VSS.n2852 0.4505
R69958 VSS.n6921 VSS.n6920 0.4505
R69959 VSS.n2854 VSS.n2853 0.4505
R69960 VSS.n6909 VSS.n6908 0.4505
R69961 VSS.n6907 VSS.n2874 0.4505
R69962 VSS.n6906 VSS.n6905 0.4505
R69963 VSS.n2876 VSS.n2875 0.4505
R69964 VSS.n6901 VSS.n6900 0.4505
R69965 VSS.n6899 VSS.n2878 0.4505
R69966 VSS.n6898 VSS.n6897 0.4505
R69967 VSS.n2880 VSS.n2879 0.4505
R69968 VSS.n6893 VSS.n6892 0.4505
R69969 VSS.n6891 VSS.n2882 0.4505
R69970 VSS.n6890 VSS.n6889 0.4505
R69971 VSS.n2884 VSS.n2883 0.4505
R69972 VSS.n6885 VSS.n6884 0.4505
R69973 VSS.n6883 VSS.n2886 0.4505
R69974 VSS.n6882 VSS.n6881 0.4505
R69975 VSS.n2888 VSS.n2887 0.4505
R69976 VSS.n6870 VSS.n6869 0.4505
R69977 VSS.n6868 VSS.n2908 0.4505
R69978 VSS.n6867 VSS.n6866 0.4505
R69979 VSS.n2910 VSS.n2909 0.4505
R69980 VSS.n6862 VSS.n6861 0.4505
R69981 VSS.n6860 VSS.n2912 0.4505
R69982 VSS.n6859 VSS.n6858 0.4505
R69983 VSS.n2914 VSS.n2913 0.4505
R69984 VSS.n6854 VSS.n6853 0.4505
R69985 VSS.n6852 VSS.n2916 0.4505
R69986 VSS.n6851 VSS.n6850 0.4505
R69987 VSS.n2918 VSS.n2917 0.4505
R69988 VSS.n6846 VSS.n6845 0.4505
R69989 VSS.n6844 VSS.n2920 0.4505
R69990 VSS.n6843 VSS.n6842 0.4505
R69991 VSS.n2922 VSS.n2921 0.4505
R69992 VSS.n3012 VSS.n3011 0.4505
R69993 VSS.n3013 VSS.n3010 0.4505
R69994 VSS.n3016 VSS.n3015 0.4505
R69995 VSS.n3017 VSS.n3009 0.4505
R69996 VSS.n3019 VSS.n3018 0.4505
R69997 VSS.n3007 VSS.n3006 0.4505
R69998 VSS.n3024 VSS.n3023 0.4505
R69999 VSS.n3025 VSS.n3005 0.4505
R70000 VSS.n3027 VSS.n3026 0.4505
R70001 VSS.n3003 VSS.n3002 0.4505
R70002 VSS.n3032 VSS.n3031 0.4505
R70003 VSS.n3033 VSS.n3001 0.4505
R70004 VSS.n3036 VSS.n3035 0.4505
R70005 VSS.n3034 VSS.n2999 0.4505
R70006 VSS.n3040 VSS.n2998 0.4505
R70007 VSS.n3042 VSS.n3041 0.4505
R70008 VSS.n3043 VSS.n2995 0.4505
R70009 VSS.n6747 VSS.n6746 0.4505
R70010 VSS.n6745 VSS.n2997 0.4505
R70011 VSS.n6744 VSS.n6743 0.4505
R70012 VSS.n3045 VSS.n3044 0.4505
R70013 VSS.n6739 VSS.n6738 0.4505
R70014 VSS.n6737 VSS.n3047 0.4505
R70015 VSS.n6736 VSS.n6735 0.4505
R70016 VSS.n3049 VSS.n3048 0.4505
R70017 VSS.n6731 VSS.n6730 0.4505
R70018 VSS.n6729 VSS.n3051 0.4505
R70019 VSS.n6728 VSS.n6727 0.4505
R70020 VSS.n3053 VSS.n3052 0.4505
R70021 VSS.n6723 VSS.n6722 0.4505
R70022 VSS.n6721 VSS.n3055 0.4505
R70023 VSS.n6720 VSS.n6719 0.4505
R70024 VSS.n3057 VSS.n3056 0.4505
R70025 VSS.n3084 VSS.n3082 0.4505
R70026 VSS.n6713 VSS.n6712 0.4505
R70027 VSS.n6711 VSS.n3083 0.4505
R70028 VSS.n6710 VSS.n6709 0.4505
R70029 VSS.n3086 VSS.n3085 0.4505
R70030 VSS.n6705 VSS.n6704 0.4505
R70031 VSS.n6703 VSS.n3089 0.4505
R70032 VSS.n6702 VSS.n6701 0.4505
R70033 VSS.n3091 VSS.n3090 0.4505
R70034 VSS.n6670 VSS.n6668 0.4505
R70035 VSS.n6689 VSS.n6688 0.4505
R70036 VSS.n6687 VSS.n6669 0.4505
R70037 VSS.n6686 VSS.n6685 0.4505
R70038 VSS.n6682 VSS.n6671 0.4505
R70039 VSS.n6681 VSS.n6680 0.4505
R70040 VSS.n6679 VSS.n6672 0.4505
R70041 VSS.n6675 VSS.n6674 0.4505
R70042 VSS.n6677 VSS.n6676 0.4505
R70043 VSS.n2818 VSS.n2805 0.4505
R70044 VSS.n2820 VSS.n2819 0.4505
R70045 VSS.n2816 VSS.n2814 0.4505
R70046 VSS.n6956 VSS.n6955 0.4505
R70047 VSS.n2817 VSS.n2815 0.4505
R70048 VSS.n6951 VSS.n6950 0.4505
R70049 VSS.n6949 VSS.n2824 0.4505
R70050 VSS.n6948 VSS.n6947 0.4505
R70051 VSS.n2829 VSS.n2826 0.4505
R70052 VSS.n6943 VSS.n6942 0.4505
R70053 VSS.n2836 VSS.n2828 0.4505
R70054 VSS.n6933 VSS.n6932 0.4505
R70055 VSS.n2848 VSS.n2847 0.4505
R70056 VSS.n6928 VSS.n6927 0.4505
R70057 VSS.n6926 VSS.n2850 0.4505
R70058 VSS.n6925 VSS.n6924 0.4505
R70059 VSS.n2855 VSS.n2852 0.4505
R70060 VSS.n6920 VSS.n6919 0.4505
R70061 VSS.n2862 VSS.n2854 0.4505
R70062 VSS.n6910 VSS.n6909 0.4505
R70063 VSS.n2874 VSS.n2873 0.4505
R70064 VSS.n6905 VSS.n6904 0.4505
R70065 VSS.n6903 VSS.n2876 0.4505
R70066 VSS.n6902 VSS.n6901 0.4505
R70067 VSS.n2878 VSS.n2877 0.4505
R70068 VSS.n6897 VSS.n6896 0.4505
R70069 VSS.n6895 VSS.n2880 0.4505
R70070 VSS.n6894 VSS.n6893 0.4505
R70071 VSS.n2882 VSS.n2881 0.4505
R70072 VSS.n6889 VSS.n6888 0.4505
R70073 VSS.n6887 VSS.n2884 0.4505
R70074 VSS.n6886 VSS.n6885 0.4505
R70075 VSS.n2889 VSS.n2886 0.4505
R70076 VSS.n6881 VSS.n6880 0.4505
R70077 VSS.n2896 VSS.n2888 0.4505
R70078 VSS.n6871 VSS.n6870 0.4505
R70079 VSS.n2908 VSS.n2907 0.4505
R70080 VSS.n6866 VSS.n6865 0.4505
R70081 VSS.n6864 VSS.n2910 0.4505
R70082 VSS.n6863 VSS.n6862 0.4505
R70083 VSS.n2912 VSS.n2911 0.4505
R70084 VSS.n6858 VSS.n6857 0.4505
R70085 VSS.n6856 VSS.n2914 0.4505
R70086 VSS.n6855 VSS.n6854 0.4505
R70087 VSS.n2916 VSS.n2915 0.4505
R70088 VSS.n6850 VSS.n6849 0.4505
R70089 VSS.n6848 VSS.n2918 0.4505
R70090 VSS.n6847 VSS.n6846 0.4505
R70091 VSS.n2923 VSS.n2920 0.4505
R70092 VSS.n6842 VSS.n6841 0.4505
R70093 VSS.n2930 VSS.n2922 0.4505
R70094 VSS.n3012 VSS.n2942 0.4505
R70095 VSS.n3013 VSS.n2948 0.4505
R70096 VSS.n3015 VSS.n3014 0.4505
R70097 VSS.n3009 VSS.n3008 0.4505
R70098 VSS.n3020 VSS.n3019 0.4505
R70099 VSS.n3021 VSS.n3007 0.4505
R70100 VSS.n3023 VSS.n3022 0.4505
R70101 VSS.n3005 VSS.n3004 0.4505
R70102 VSS.n3028 VSS.n3027 0.4505
R70103 VSS.n3029 VSS.n3003 0.4505
R70104 VSS.n3031 VSS.n3030 0.4505
R70105 VSS.n3001 VSS.n3000 0.4505
R70106 VSS.n3037 VSS.n3036 0.4505
R70107 VSS.n3038 VSS.n2999 0.4505
R70108 VSS.n3040 VSS.n3039 0.4505
R70109 VSS.n3041 VSS.n2975 0.4505
R70110 VSS.n2995 VSS.n2981 0.4505
R70111 VSS.n6748 VSS.n6747 0.4505
R70112 VSS.n2997 VSS.n2996 0.4505
R70113 VSS.n6743 VSS.n6742 0.4505
R70114 VSS.n6741 VSS.n3045 0.4505
R70115 VSS.n6740 VSS.n6739 0.4505
R70116 VSS.n3047 VSS.n3046 0.4505
R70117 VSS.n6735 VSS.n6734 0.4505
R70118 VSS.n6733 VSS.n3049 0.4505
R70119 VSS.n6732 VSS.n6731 0.4505
R70120 VSS.n3051 VSS.n3050 0.4505
R70121 VSS.n6727 VSS.n6726 0.4505
R70122 VSS.n6725 VSS.n3053 0.4505
R70123 VSS.n6724 VSS.n6723 0.4505
R70124 VSS.n3055 VSS.n3054 0.4505
R70125 VSS.n6719 VSS.n6718 0.4505
R70126 VSS.n3063 VSS.n3057 0.4505
R70127 VSS.n3082 VSS.n3076 0.4505
R70128 VSS.n6714 VSS.n6713 0.4505
R70129 VSS.n3087 VSS.n3083 0.4505
R70130 VSS.n6709 VSS.n6708 0.4505
R70131 VSS.n6707 VSS.n3086 0.4505
R70132 VSS.n6706 VSS.n6705 0.4505
R70133 VSS.n3089 VSS.n3088 0.4505
R70134 VSS.n6701 VSS.n6700 0.4505
R70135 VSS.n3098 VSS.n3091 0.4505
R70136 VSS.n6668 VSS.n3105 0.4505
R70137 VSS.n6690 VSS.n6689 0.4505
R70138 VSS.n6669 VSS.n6667 0.4505
R70139 VSS.n6685 VSS.n6684 0.4505
R70140 VSS.n6683 VSS.n6682 0.4505
R70141 VSS.n6681 VSS.n504 0.4505
R70142 VSS.n6672 VSS.n510 0.4505
R70143 VSS.n9611 VSS.n9610 0.4505
R70144 VSS.n3918 VSS.n3915 0.4505
R70145 VSS.n3921 VSS.n3920 0.4505
R70146 VSS.n3922 VSS.n3914 0.4505
R70147 VSS.n3925 VSS.n3924 0.4505
R70148 VSS.n3923 VSS.n3912 0.4505
R70149 VSS.n3929 VSS.n3911 0.4505
R70150 VSS.n3931 VSS.n3930 0.4505
R70151 VSS.n3932 VSS.n3909 0.4505
R70152 VSS.n6211 VSS.n6210 0.4505
R70153 VSS.n6209 VSS.n3910 0.4505
R70154 VSS.n6208 VSS.n6207 0.4505
R70155 VSS.n3934 VSS.n3933 0.4505
R70156 VSS.n6203 VSS.n6202 0.4505
R70157 VSS.n6201 VSS.n3936 0.4505
R70158 VSS.n6200 VSS.n6199 0.4505
R70159 VSS.n3938 VSS.n3937 0.4505
R70160 VSS.n3963 VSS.n3962 0.4505
R70161 VSS.n3964 VSS.n3959 0.4505
R70162 VSS.n6191 VSS.n6190 0.4505
R70163 VSS.n6189 VSS.n3960 0.4505
R70164 VSS.n6188 VSS.n6187 0.4505
R70165 VSS.n3966 VSS.n3965 0.4505
R70166 VSS.n6183 VSS.n6182 0.4505
R70167 VSS.n6181 VSS.n3968 0.4505
R70168 VSS.n6180 VSS.n6179 0.4505
R70169 VSS.n3970 VSS.n3969 0.4505
R70170 VSS.n6175 VSS.n6174 0.4505
R70171 VSS.n6173 VSS.n3972 0.4505
R70172 VSS.n6172 VSS.n6171 0.4505
R70173 VSS.n3974 VSS.n3973 0.4505
R70174 VSS.n6167 VSS.n6166 0.4505
R70175 VSS.n6165 VSS.n3976 0.4505
R70176 VSS.n6164 VSS.n6163 0.4505
R70177 VSS.n3978 VSS.n3977 0.4505
R70178 VSS.n6155 VSS.n6154 0.4505
R70179 VSS.n6153 VSS.n3998 0.4505
R70180 VSS.n6152 VSS.n6151 0.4505
R70181 VSS.n4000 VSS.n3999 0.4505
R70182 VSS.n6147 VSS.n6146 0.4505
R70183 VSS.n6145 VSS.n4002 0.4505
R70184 VSS.n6144 VSS.n6143 0.4505
R70185 VSS.n4004 VSS.n4003 0.4505
R70186 VSS.n6139 VSS.n6138 0.4505
R70187 VSS.n6137 VSS.n4006 0.4505
R70188 VSS.n6136 VSS.n6135 0.4505
R70189 VSS.n4008 VSS.n4007 0.4505
R70190 VSS.n6131 VSS.n6130 0.4505
R70191 VSS.n6129 VSS.n4010 0.4505
R70192 VSS.n6128 VSS.n6127 0.4505
R70193 VSS.n4012 VSS.n4011 0.4505
R70194 VSS.n4181 VSS.n4179 0.4505
R70195 VSS.n4184 VSS.n4183 0.4505
R70196 VSS.n4185 VSS.n4177 0.4505
R70197 VSS.n4220 VSS.n4219 0.4505
R70198 VSS.n4218 VSS.n4178 0.4505
R70199 VSS.n4217 VSS.n4216 0.4505
R70200 VSS.n4187 VSS.n4186 0.4505
R70201 VSS.n4212 VSS.n4211 0.4505
R70202 VSS.n4210 VSS.n4189 0.4505
R70203 VSS.n4209 VSS.n4208 0.4505
R70204 VSS.n4191 VSS.n4190 0.4505
R70205 VSS.n4204 VSS.n4203 0.4505
R70206 VSS.n4202 VSS.n4193 0.4505
R70207 VSS.n4201 VSS.n4200 0.4505
R70208 VSS.n4197 VSS.n4194 0.4505
R70209 VSS.n4196 VSS.n4195 0.4505
R70210 VSS.n331 VSS.n328 0.4505
R70211 VSS.n9676 VSS.n9675 0.4505
R70212 VSS.n9674 VSS.n330 0.4505
R70213 VSS.n9673 VSS.n9672 0.4505
R70214 VSS.n333 VSS.n332 0.4505
R70215 VSS.n9668 VSS.n9667 0.4505
R70216 VSS.n9666 VSS.n335 0.4505
R70217 VSS.n9665 VSS.n9664 0.4505
R70218 VSS.n337 VSS.n336 0.4505
R70219 VSS.n9660 VSS.n9659 0.4505
R70220 VSS.n9658 VSS.n339 0.4505
R70221 VSS.n9657 VSS.n9656 0.4505
R70222 VSS.n341 VSS.n340 0.4505
R70223 VSS.n9652 VSS.n9651 0.4505
R70224 VSS.n9650 VSS.n343 0.4505
R70225 VSS.n9649 VSS.n9648 0.4505
R70226 VSS.n345 VSS.n344 0.4505
R70227 VSS.n372 VSS.n371 0.4505
R70228 VSS.n373 VSS.n368 0.4505
R70229 VSS.n9642 VSS.n9641 0.4505
R70230 VSS.n9640 VSS.n369 0.4505
R70231 VSS.n9639 VSS.n9638 0.4505
R70232 VSS.n375 VSS.n374 0.4505
R70233 VSS.n9634 VSS.n9633 0.4505
R70234 VSS.n9632 VSS.n377 0.4505
R70235 VSS.n9631 VSS.n9630 0.4505
R70236 VSS.n379 VSS.n378 0.4505
R70237 VSS.n9622 VSS.n9621 0.4505
R70238 VSS.n9620 VSS.n399 0.4505
R70239 VSS.n9619 VSS.n9618 0.4505
R70240 VSS.n401 VSS.n400 0.4505
R70241 VSS.n9614 VSS.n9613 0.4505
R70242 VSS.n9612 VSS.n403 0.4505
R70243 VSS.n413 VSS.n405 0.4505
R70244 VSS.n9610 VSS.n9609 0.4505
R70245 VSS.n3916 VSS.n3842 0.4505
R70246 VSS.n3918 VSS.n3917 0.4505
R70247 VSS.n3920 VSS.n3919 0.4505
R70248 VSS.n3914 VSS.n3913 0.4505
R70249 VSS.n3926 VSS.n3925 0.4505
R70250 VSS.n3927 VSS.n3912 0.4505
R70251 VSS.n3929 VSS.n3928 0.4505
R70252 VSS.n3930 VSS.n3895 0.4505
R70253 VSS.n3909 VSS.n3901 0.4505
R70254 VSS.n6212 VSS.n6211 0.4505
R70255 VSS.n3910 VSS.n3908 0.4505
R70256 VSS.n6207 VSS.n6206 0.4505
R70257 VSS.n6205 VSS.n3934 0.4505
R70258 VSS.n6204 VSS.n6203 0.4505
R70259 VSS.n3936 VSS.n3935 0.4505
R70260 VSS.n6199 VSS.n6198 0.4505
R70261 VSS.n3944 VSS.n3938 0.4505
R70262 VSS.n3962 VSS.n3961 0.4505
R70263 VSS.n3959 VSS.n3957 0.4505
R70264 VSS.n6192 VSS.n6191 0.4505
R70265 VSS.n3960 VSS.n3958 0.4505
R70266 VSS.n6187 VSS.n6186 0.4505
R70267 VSS.n6185 VSS.n3966 0.4505
R70268 VSS.n6184 VSS.n6183 0.4505
R70269 VSS.n3968 VSS.n3967 0.4505
R70270 VSS.n6179 VSS.n6178 0.4505
R70271 VSS.n6177 VSS.n3970 0.4505
R70272 VSS.n6176 VSS.n6175 0.4505
R70273 VSS.n3972 VSS.n3971 0.4505
R70274 VSS.n6171 VSS.n6170 0.4505
R70275 VSS.n6169 VSS.n3974 0.4505
R70276 VSS.n6168 VSS.n6167 0.4505
R70277 VSS.n3979 VSS.n3976 0.4505
R70278 VSS.n6163 VSS.n6162 0.4505
R70279 VSS.n3986 VSS.n3978 0.4505
R70280 VSS.n6156 VSS.n6155 0.4505
R70281 VSS.n3998 VSS.n3997 0.4505
R70282 VSS.n6151 VSS.n6150 0.4505
R70283 VSS.n6149 VSS.n4000 0.4505
R70284 VSS.n6148 VSS.n6147 0.4505
R70285 VSS.n4002 VSS.n4001 0.4505
R70286 VSS.n6143 VSS.n6142 0.4505
R70287 VSS.n6141 VSS.n4004 0.4505
R70288 VSS.n6140 VSS.n6139 0.4505
R70289 VSS.n4006 VSS.n4005 0.4505
R70290 VSS.n6135 VSS.n6134 0.4505
R70291 VSS.n6133 VSS.n4008 0.4505
R70292 VSS.n6132 VSS.n6131 0.4505
R70293 VSS.n4013 VSS.n4010 0.4505
R70294 VSS.n6127 VSS.n6126 0.4505
R70295 VSS.n4020 VSS.n4012 0.4505
R70296 VSS.n4181 VSS.n4180 0.4505
R70297 VSS.n4183 VSS.n4182 0.4505
R70298 VSS.n4177 VSS.n4172 0.4505
R70299 VSS.n4221 VSS.n4220 0.4505
R70300 VSS.n4178 VSS.n4176 0.4505
R70301 VSS.n4216 VSS.n4215 0.4505
R70302 VSS.n4214 VSS.n4187 0.4505
R70303 VSS.n4213 VSS.n4212 0.4505
R70304 VSS.n4189 VSS.n4188 0.4505
R70305 VSS.n4208 VSS.n4207 0.4505
R70306 VSS.n4206 VSS.n4191 0.4505
R70307 VSS.n4205 VSS.n4204 0.4505
R70308 VSS.n4193 VSS.n4192 0.4505
R70309 VSS.n4200 VSS.n4199 0.4505
R70310 VSS.n4198 VSS.n4197 0.4505
R70311 VSS.n4196 VSS.n311 0.4505
R70312 VSS.n328 VSS.n317 0.4505
R70313 VSS.n9677 VSS.n9676 0.4505
R70314 VSS.n330 VSS.n329 0.4505
R70315 VSS.n9672 VSS.n9671 0.4505
R70316 VSS.n9670 VSS.n333 0.4505
R70317 VSS.n9669 VSS.n9668 0.4505
R70318 VSS.n335 VSS.n334 0.4505
R70319 VSS.n9664 VSS.n9663 0.4505
R70320 VSS.n9662 VSS.n337 0.4505
R70321 VSS.n9661 VSS.n9660 0.4505
R70322 VSS.n339 VSS.n338 0.4505
R70323 VSS.n9656 VSS.n9655 0.4505
R70324 VSS.n9654 VSS.n341 0.4505
R70325 VSS.n9653 VSS.n9652 0.4505
R70326 VSS.n343 VSS.n342 0.4505
R70327 VSS.n9648 VSS.n9647 0.4505
R70328 VSS.n351 VSS.n345 0.4505
R70329 VSS.n371 VSS.n370 0.4505
R70330 VSS.n368 VSS.n363 0.4505
R70331 VSS.n9643 VSS.n9642 0.4505
R70332 VSS.n369 VSS.n367 0.4505
R70333 VSS.n9638 VSS.n9637 0.4505
R70334 VSS.n9636 VSS.n375 0.4505
R70335 VSS.n9635 VSS.n9634 0.4505
R70336 VSS.n380 VSS.n377 0.4505
R70337 VSS.n9630 VSS.n9629 0.4505
R70338 VSS.n387 VSS.n379 0.4505
R70339 VSS.n9623 VSS.n9622 0.4505
R70340 VSS.n399 VSS.n398 0.4505
R70341 VSS.n9618 VSS.n9617 0.4505
R70342 VSS.n9616 VSS.n401 0.4505
R70343 VSS.n9615 VSS.n9614 0.4505
R70344 VSS.n406 VSS.n403 0.4505
R70345 VSS.n5488 VSS.n5487 0.4505
R70346 VSS.n6236 VSS.n6234 0.4505
R70347 VSS.n6233 VSS.n3875 0.4505
R70348 VSS.n6232 VSS.n6231 0.4505
R70349 VSS.n3877 VSS.n3876 0.4505
R70350 VSS.n6227 VSS.n6226 0.4505
R70351 VSS.n6225 VSS.n3879 0.4505
R70352 VSS.n6224 VSS.n6223 0.4505
R70353 VSS.n3881 VSS.n3880 0.4505
R70354 VSS.n5278 VSS.n5277 0.4505
R70355 VSS.n5281 VSS.n5280 0.4505
R70356 VSS.n5282 VSS.n5276 0.4505
R70357 VSS.n5284 VSS.n5283 0.4505
R70358 VSS.n5274 VSS.n5273 0.4505
R70359 VSS.n5289 VSS.n5288 0.4505
R70360 VSS.n5290 VSS.n5272 0.4505
R70361 VSS.n5292 VSS.n5291 0.4505
R70362 VSS.n4312 VSS.n4311 0.4505
R70363 VSS.n5306 VSS.n5305 0.4505
R70364 VSS.n5307 VSS.n4310 0.4505
R70365 VSS.n5309 VSS.n5308 0.4505
R70366 VSS.n4308 VSS.n4307 0.4505
R70367 VSS.n5314 VSS.n5313 0.4505
R70368 VSS.n5315 VSS.n4306 0.4505
R70369 VSS.n5317 VSS.n5316 0.4505
R70370 VSS.n4304 VSS.n4303 0.4505
R70371 VSS.n5322 VSS.n5321 0.4505
R70372 VSS.n5323 VSS.n4302 0.4505
R70373 VSS.n5325 VSS.n5324 0.4505
R70374 VSS.n4300 VSS.n4299 0.4505
R70375 VSS.n5330 VSS.n5329 0.4505
R70376 VSS.n5331 VSS.n4296 0.4505
R70377 VSS.n5629 VSS.n5628 0.4505
R70378 VSS.n5627 VSS.n4298 0.4505
R70379 VSS.n5626 VSS.n5625 0.4505
R70380 VSS.n5623 VSS.n5332 0.4505
R70381 VSS.n5336 VSS.n5333 0.4505
R70382 VSS.n5619 VSS.n5618 0.4505
R70383 VSS.n5617 VSS.n5335 0.4505
R70384 VSS.n5616 VSS.n5615 0.4505
R70385 VSS.n5338 VSS.n5337 0.4505
R70386 VSS.n5611 VSS.n5610 0.4505
R70387 VSS.n5609 VSS.n5340 0.4505
R70388 VSS.n5608 VSS.n5607 0.4505
R70389 VSS.n5342 VSS.n5341 0.4505
R70390 VSS.n5603 VSS.n5602 0.4505
R70391 VSS.n5601 VSS.n5344 0.4505
R70392 VSS.n5600 VSS.n5599 0.4505
R70393 VSS.n5598 VSS.n5345 0.4505
R70394 VSS.n5597 VSS.n5595 0.4505
R70395 VSS.n5594 VSS.n5347 0.4505
R70396 VSS.n5593 VSS.n5592 0.4505
R70397 VSS.n5591 VSS.n5348 0.4505
R70398 VSS.n5590 VSS.n5588 0.4505
R70399 VSS.n5587 VSS.n5349 0.4505
R70400 VSS.n5586 VSS.n5585 0.4505
R70401 VSS.n5351 VSS.n5350 0.4505
R70402 VSS.n5581 VSS.n5580 0.4505
R70403 VSS.n5579 VSS.n5354 0.4505
R70404 VSS.n5578 VSS.n5577 0.4505
R70405 VSS.n5356 VSS.n5355 0.4505
R70406 VSS.n5573 VSS.n5572 0.4505
R70407 VSS.n5571 VSS.n5358 0.4505
R70408 VSS.n5570 VSS.n5569 0.4505
R70409 VSS.n5360 VSS.n5359 0.4505
R70410 VSS.n5565 VSS.n5564 0.4505
R70411 VSS.n5563 VSS.n5361 0.4505
R70412 VSS.n5562 VSS.n5561 0.4505
R70413 VSS.n5560 VSS.n5362 0.4505
R70414 VSS.n5558 VSS.n5556 0.4505
R70415 VSS.n5555 VSS.n5363 0.4505
R70416 VSS.n5554 VSS.n5553 0.4505
R70417 VSS.n5365 VSS.n5364 0.4505
R70418 VSS.n5549 VSS.n5548 0.4505
R70419 VSS.n5547 VSS.n5368 0.4505
R70420 VSS.n5546 VSS.n5545 0.4505
R70421 VSS.n5370 VSS.n5369 0.4505
R70422 VSS.n5541 VSS.n5540 0.4505
R70423 VSS.n5539 VSS.n5372 0.4505
R70424 VSS.n5538 VSS.n5537 0.4505
R70425 VSS.n5374 VSS.n5373 0.4505
R70426 VSS.n5533 VSS.n5532 0.4505
R70427 VSS.n5531 VSS.n5376 0.4505
R70428 VSS.n5530 VSS.n5529 0.4505
R70429 VSS.n5378 VSS.n5377 0.4505
R70430 VSS.n5399 VSS.n5397 0.4505
R70431 VSS.n5520 VSS.n5519 0.4505
R70432 VSS.n5518 VSS.n5398 0.4505
R70433 VSS.n5517 VSS.n5516 0.4505
R70434 VSS.n5401 VSS.n5400 0.4505
R70435 VSS.n5512 VSS.n5511 0.4505
R70436 VSS.n5510 VSS.n5403 0.4505
R70437 VSS.n5509 VSS.n5508 0.4505
R70438 VSS.n5405 VSS.n5404 0.4505
R70439 VSS.n5499 VSS.n5498 0.4505
R70440 VSS.n5497 VSS.n5423 0.4505
R70441 VSS.n5496 VSS.n5495 0.4505
R70442 VSS.n5425 VSS.n5424 0.4505
R70443 VSS.n5491 VSS.n5490 0.4505
R70444 VSS.n5489 VSS.n5427 0.4505
R70445 VSS.n5437 VSS.n5429 0.4505
R70446 VSS.n5487 VSS.n5486 0.4505
R70447 VSS.n6238 VSS.n6237 0.4505
R70448 VSS.n6236 VSS.n6235 0.4505
R70449 VSS.n3875 VSS.n3874 0.4505
R70450 VSS.n6231 VSS.n6230 0.4505
R70451 VSS.n6229 VSS.n3877 0.4505
R70452 VSS.n6228 VSS.n6227 0.4505
R70453 VSS.n3879 VSS.n3878 0.4505
R70454 VSS.n6223 VSS.n6222 0.4505
R70455 VSS.n3887 VSS.n3881 0.4505
R70456 VSS.n5278 VSS.n3893 0.4505
R70457 VSS.n5280 VSS.n5279 0.4505
R70458 VSS.n5276 VSS.n5275 0.4505
R70459 VSS.n5285 VSS.n5284 0.4505
R70460 VSS.n5286 VSS.n5274 0.4505
R70461 VSS.n5288 VSS.n5287 0.4505
R70462 VSS.n5272 VSS.n5269 0.4505
R70463 VSS.n5293 VSS.n5292 0.4505
R70464 VSS.n5295 VSS.n4312 0.4505
R70465 VSS.n5305 VSS.n5304 0.4505
R70466 VSS.n4310 VSS.n4309 0.4505
R70467 VSS.n5310 VSS.n5309 0.4505
R70468 VSS.n5311 VSS.n4308 0.4505
R70469 VSS.n5313 VSS.n5312 0.4505
R70470 VSS.n4306 VSS.n4305 0.4505
R70471 VSS.n5318 VSS.n5317 0.4505
R70472 VSS.n5319 VSS.n4304 0.4505
R70473 VSS.n5321 VSS.n5320 0.4505
R70474 VSS.n4302 VSS.n4301 0.4505
R70475 VSS.n5326 VSS.n5325 0.4505
R70476 VSS.n5327 VSS.n4300 0.4505
R70477 VSS.n5329 VSS.n5328 0.4505
R70478 VSS.n4296 VSS.n4292 0.4505
R70479 VSS.n5630 VSS.n5629 0.4505
R70480 VSS.n4298 VSS.n4297 0.4505
R70481 VSS.n5625 VSS.n5624 0.4505
R70482 VSS.n5623 VSS.n5622 0.4505
R70483 VSS.n5621 VSS.n5333 0.4505
R70484 VSS.n5620 VSS.n5619 0.4505
R70485 VSS.n5335 VSS.n5334 0.4505
R70486 VSS.n5615 VSS.n5614 0.4505
R70487 VSS.n5613 VSS.n5338 0.4505
R70488 VSS.n5612 VSS.n5611 0.4505
R70489 VSS.n5340 VSS.n5339 0.4505
R70490 VSS.n5607 VSS.n5606 0.4505
R70491 VSS.n5605 VSS.n5342 0.4505
R70492 VSS.n5604 VSS.n5603 0.4505
R70493 VSS.n5344 VSS.n5343 0.4505
R70494 VSS.n5599 VSS.n4265 0.4505
R70495 VSS.n5598 VSS.n4271 0.4505
R70496 VSS.n5597 VSS.n5596 0.4505
R70497 VSS.n5347 VSS.n5346 0.4505
R70498 VSS.n5592 VSS.n4247 0.4505
R70499 VSS.n5591 VSS.n4253 0.4505
R70500 VSS.n5590 VSS.n5589 0.4505
R70501 VSS.n5352 VSS.n5349 0.4505
R70502 VSS.n5585 VSS.n5584 0.4505
R70503 VSS.n5583 VSS.n5351 0.4505
R70504 VSS.n5582 VSS.n5581 0.4505
R70505 VSS.n5354 VSS.n5353 0.4505
R70506 VSS.n5577 VSS.n5576 0.4505
R70507 VSS.n5575 VSS.n5356 0.4505
R70508 VSS.n5574 VSS.n5573 0.4505
R70509 VSS.n5358 VSS.n5357 0.4505
R70510 VSS.n5569 VSS.n5568 0.4505
R70511 VSS.n5567 VSS.n5360 0.4505
R70512 VSS.n5566 VSS.n5565 0.4505
R70513 VSS.n5361 VSS.n290 0.4505
R70514 VSS.n5561 VSS.n295 0.4505
R70515 VSS.n5560 VSS.n5559 0.4505
R70516 VSS.n5558 VSS.n5557 0.4505
R70517 VSS.n5366 VSS.n5363 0.4505
R70518 VSS.n5553 VSS.n5552 0.4505
R70519 VSS.n5551 VSS.n5365 0.4505
R70520 VSS.n5550 VSS.n5549 0.4505
R70521 VSS.n5368 VSS.n5367 0.4505
R70522 VSS.n5545 VSS.n5544 0.4505
R70523 VSS.n5543 VSS.n5370 0.4505
R70524 VSS.n5542 VSS.n5541 0.4505
R70525 VSS.n5372 VSS.n5371 0.4505
R70526 VSS.n5537 VSS.n5536 0.4505
R70527 VSS.n5535 VSS.n5374 0.4505
R70528 VSS.n5534 VSS.n5533 0.4505
R70529 VSS.n5376 VSS.n5375 0.4505
R70530 VSS.n5529 VSS.n5528 0.4505
R70531 VSS.n5385 VSS.n5378 0.4505
R70532 VSS.n5397 VSS.n5392 0.4505
R70533 VSS.n5521 VSS.n5520 0.4505
R70534 VSS.n5398 VSS.n5396 0.4505
R70535 VSS.n5516 VSS.n5515 0.4505
R70536 VSS.n5514 VSS.n5401 0.4505
R70537 VSS.n5513 VSS.n5512 0.4505
R70538 VSS.n5406 VSS.n5403 0.4505
R70539 VSS.n5508 VSS.n5507 0.4505
R70540 VSS.n5413 VSS.n5405 0.4505
R70541 VSS.n5500 VSS.n5499 0.4505
R70542 VSS.n5423 VSS.n5422 0.4505
R70543 VSS.n5495 VSS.n5494 0.4505
R70544 VSS.n5493 VSS.n5425 0.4505
R70545 VSS.n5492 VSS.n5491 0.4505
R70546 VSS.n5430 VSS.n5427 0.4505
R70547 VSS.n9792 VSS.n9791 0.4505
R70548 VSS.n187 VSS.n186 0.4505
R70549 VSS.n4737 VSS.n4736 0.4505
R70550 VSS.n4728 VSS.n4583 0.4505
R70551 VSS.n4766 VSS.n4765 0.4505
R70552 VSS.n4581 VSS.n4580 0.4505
R70553 VSS.n4771 VSS.n4770 0.4505
R70554 VSS.n4772 VSS.n4579 0.4505
R70555 VSS.n4774 VSS.n4773 0.4505
R70556 VSS.n4577 VSS.n4572 0.4505
R70557 VSS.n4779 VSS.n4778 0.4505
R70558 VSS.n4562 VSS.n4551 0.4505
R70559 VSS.n4788 VSS.n4787 0.4505
R70560 VSS.n4549 VSS.n4548 0.4505
R70561 VSS.n4793 VSS.n4792 0.4505
R70562 VSS.n4794 VSS.n4547 0.4505
R70563 VSS.n4796 VSS.n4795 0.4505
R70564 VSS.n4545 VSS.n4333 0.4505
R70565 VSS.n4800 VSS.n4337 0.4505
R70566 VSS.n4802 VSS.n4801 0.4505
R70567 VSS.n4804 VSS.n4803 0.4505
R70568 VSS.n4543 VSS.n4542 0.4505
R70569 VSS.n4809 VSS.n4808 0.4505
R70570 VSS.n4810 VSS.n4541 0.4505
R70571 VSS.n4812 VSS.n4811 0.4505
R70572 VSS.n4539 VSS.n4538 0.4505
R70573 VSS.n4817 VSS.n4816 0.4505
R70574 VSS.n4818 VSS.n4537 0.4505
R70575 VSS.n4820 VSS.n4819 0.4505
R70576 VSS.n4535 VSS.n4534 0.4505
R70577 VSS.n4825 VSS.n4824 0.4505
R70578 VSS.n4826 VSS.n4533 0.4505
R70579 VSS.n4828 VSS.n4827 0.4505
R70580 VSS.n4529 VSS.n4525 0.4505
R70581 VSS.n5060 VSS.n5059 0.4505
R70582 VSS.n4531 VSS.n4530 0.4505
R70583 VSS.n5055 VSS.n5054 0.4505
R70584 VSS.n5053 VSS.n5052 0.4505
R70585 VSS.n5051 VSS.n4832 0.4505
R70586 VSS.n5050 VSS.n5049 0.4505
R70587 VSS.n4834 VSS.n4833 0.4505
R70588 VSS.n5045 VSS.n5044 0.4505
R70589 VSS.n5043 VSS.n4837 0.4505
R70590 VSS.n5042 VSS.n5041 0.4505
R70591 VSS.n4839 VSS.n4838 0.4505
R70592 VSS.n5037 VSS.n5036 0.4505
R70593 VSS.n5035 VSS.n4841 0.4505
R70594 VSS.n5034 VSS.n5033 0.4505
R70595 VSS.n4843 VSS.n4842 0.4505
R70596 VSS.n5029 VSS.n4494 0.4505
R70597 VSS.n5028 VSS.n4499 0.4505
R70598 VSS.n5027 VSS.n5026 0.4505
R70599 VSS.n4848 VSS.n4845 0.4505
R70600 VSS.n5022 VSS.n5021 0.4505
R70601 VSS.n4854 VSS.n4847 0.4505
R70602 VSS.n4977 VSS.n4975 0.4505
R70603 VSS.n5017 VSS.n5016 0.4505
R70604 VSS.n4978 VSS.n4976 0.4505
R70605 VSS.n5012 VSS.n5011 0.4505
R70606 VSS.n5010 VSS.n4981 0.4505
R70607 VSS.n5009 VSS.n5008 0.4505
R70608 VSS.n4983 VSS.n4982 0.4505
R70609 VSS.n5004 VSS.n5003 0.4505
R70610 VSS.n5002 VSS.n4985 0.4505
R70611 VSS.n5001 VSS.n5000 0.4505
R70612 VSS.n4987 VSS.n4986 0.4505
R70613 VSS.n4996 VSS.n4995 0.4505
R70614 VSS.n4994 VSS.n4993 0.4505
R70615 VSS.n4992 VSS.n259 0.4505
R70616 VSS.n4989 VSS.n263 0.4505
R70617 VSS.n268 VSS.n249 0.4505
R70618 VSS.n9698 VSS.n9697 0.4505
R70619 VSS.n247 VSS.n246 0.4505
R70620 VSS.n9703 VSS.n9702 0.4505
R70621 VSS.n9704 VSS.n245 0.4505
R70622 VSS.n9706 VSS.n9705 0.4505
R70623 VSS.n243 VSS.n242 0.4505
R70624 VSS.n9711 VSS.n9710 0.4505
R70625 VSS.n9712 VSS.n241 0.4505
R70626 VSS.n9714 VSS.n9713 0.4505
R70627 VSS.n239 VSS.n238 0.4505
R70628 VSS.n9719 VSS.n9718 0.4505
R70629 VSS.n9720 VSS.n237 0.4505
R70630 VSS.n9722 VSS.n9721 0.4505
R70631 VSS.n233 VSS.n229 0.4505
R70632 VSS.n9747 VSS.n9746 0.4505
R70633 VSS.n235 VSS.n234 0.4505
R70634 VSS.n9742 VSS.n9741 0.4505
R70635 VSS.n9740 VSS.n9739 0.4505
R70636 VSS.n9738 VSS.n9726 0.4505
R70637 VSS.n9737 VSS.n9736 0.4505
R70638 VSS.n9728 VSS.n9727 0.4505
R70639 VSS.n9732 VSS.n206 0.4505
R70640 VSS.n9731 VSS.n211 0.4505
R70641 VSS.n203 VSS.n193 0.4505
R70642 VSS.n9780 VSS.n9779 0.4505
R70643 VSS.n191 VSS.n190 0.4505
R70644 VSS.n9785 VSS.n9784 0.4505
R70645 VSS.n9786 VSS.n189 0.4505
R70646 VSS.n9788 VSS.n9787 0.4505
R70647 VSS.n185 VSS.n180 0.4505
R70648 VSS.n9797 VSS.n9796 0.4505
R70649 VSS.n7856 VSS.n7855 0.4505
R70650 VSS.n7285 VSS.n7284 0.4505
R70651 VSS.n7851 VSS.n7850 0.4505
R70652 VSS.n7849 VSS.n7600 0.4505
R70653 VSS.n7848 VSS.n7847 0.4505
R70654 VSS.n7602 VSS.n7601 0.4505
R70655 VSS.n7843 VSS.n7842 0.4505
R70656 VSS.n7841 VSS.n7604 0.4505
R70657 VSS.n7840 VSS.n7839 0.4505
R70658 VSS.n7606 VSS.n7605 0.4505
R70659 VSS.n7835 VSS.n7834 0.4505
R70660 VSS.n7833 VSS.n7608 0.4505
R70661 VSS.n7832 VSS.n7831 0.4505
R70662 VSS.n7610 VSS.n7609 0.4505
R70663 VSS.n7827 VSS.n7826 0.4505
R70664 VSS.n7825 VSS.n7612 0.4505
R70665 VSS.n7824 VSS.n7823 0.4505
R70666 VSS.n7614 VSS.n7613 0.4505
R70667 VSS.n7819 VSS.n7818 0.4505
R70668 VSS.n7817 VSS.n7616 0.4505
R70669 VSS.n7816 VSS.n7815 0.4505
R70670 VSS.n7618 VSS.n7617 0.4505
R70671 VSS.n7811 VSS.n7810 0.4505
R70672 VSS.n7809 VSS.n7620 0.4505
R70673 VSS.n7808 VSS.n7807 0.4505
R70674 VSS.n7622 VSS.n7621 0.4505
R70675 VSS.n7803 VSS.n7802 0.4505
R70676 VSS.n7801 VSS.n7624 0.4505
R70677 VSS.n7800 VSS.n7799 0.4505
R70678 VSS.n7626 VSS.n7625 0.4505
R70679 VSS.n7795 VSS.n7794 0.4505
R70680 VSS.n7793 VSS.n7628 0.4505
R70681 VSS.n7792 VSS.n7791 0.4505
R70682 VSS.n7630 VSS.n7629 0.4505
R70683 VSS.n7787 VSS.n7786 0.4505
R70684 VSS.n7785 VSS.n7632 0.4505
R70685 VSS.n7784 VSS.n7783 0.4505
R70686 VSS.n7634 VSS.n7633 0.4505
R70687 VSS.n7779 VSS.n7778 0.4505
R70688 VSS.n7777 VSS.n7636 0.4505
R70689 VSS.n7776 VSS.n7775 0.4505
R70690 VSS.n7638 VSS.n7637 0.4505
R70691 VSS.n7771 VSS.n7770 0.4505
R70692 VSS.n7769 VSS.n7640 0.4505
R70693 VSS.n7768 VSS.n7767 0.4505
R70694 VSS.n7642 VSS.n7641 0.4505
R70695 VSS.n7763 VSS.n7762 0.4505
R70696 VSS.n7761 VSS.n7644 0.4505
R70697 VSS.n7760 VSS.n7759 0.4505
R70698 VSS.n7646 VSS.n7645 0.4505
R70699 VSS.n7755 VSS.n7754 0.4505
R70700 VSS.n7753 VSS.n7648 0.4505
R70701 VSS.n7752 VSS.n7751 0.4505
R70702 VSS.n7650 VSS.n7649 0.4505
R70703 VSS.n7747 VSS.n7746 0.4505
R70704 VSS.n7745 VSS.n7652 0.4505
R70705 VSS.n7744 VSS.n7743 0.4505
R70706 VSS.n7654 VSS.n7653 0.4505
R70707 VSS.n7739 VSS.n7738 0.4505
R70708 VSS.n7737 VSS.n7656 0.4505
R70709 VSS.n7736 VSS.n7735 0.4505
R70710 VSS.n7658 VSS.n7657 0.4505
R70711 VSS.n7731 VSS.n7730 0.4505
R70712 VSS.n7729 VSS.n7660 0.4505
R70713 VSS.n7728 VSS.n7727 0.4505
R70714 VSS.n7662 VSS.n7661 0.4505
R70715 VSS.n7723 VSS.n7722 0.4505
R70716 VSS.n7721 VSS.n7664 0.4505
R70717 VSS.n7720 VSS.n7719 0.4505
R70718 VSS.n7666 VSS.n7665 0.4505
R70719 VSS.n7715 VSS.n7714 0.4505
R70720 VSS.n7713 VSS.n7668 0.4505
R70721 VSS.n7712 VSS.n7711 0.4505
R70722 VSS.n7670 VSS.n7669 0.4505
R70723 VSS.n7707 VSS.n7706 0.4505
R70724 VSS.n7705 VSS.n7672 0.4505
R70725 VSS.n7704 VSS.n7703 0.4505
R70726 VSS.n7674 VSS.n7673 0.4505
R70727 VSS.n7699 VSS.n7698 0.4505
R70728 VSS.n7697 VSS.n7676 0.4505
R70729 VSS.n7696 VSS.n7695 0.4505
R70730 VSS.n7678 VSS.n7677 0.4505
R70731 VSS.n7691 VSS.n7690 0.4505
R70732 VSS.n7689 VSS.n7680 0.4505
R70733 VSS.n7688 VSS.n7687 0.4505
R70734 VSS.n7684 VSS.n7681 0.4505
R70735 VSS.n7683 VSS.n7682 0.4505
R70736 VSS.n9914 VSS.n9913 0.4505
R70737 VSS.n9912 VSS.n2 0.4505
R70738 VSS.n9911 VSS.n9910 0.4505
R70739 VSS.n7875 VSS.n7874 0.4505
R70740 VSS.n7873 VSS.n7274 0.4505
R70741 VSS.n7872 VSS.n7871 0.4505
R70742 VSS.n7276 VSS.n7275 0.4505
R70743 VSS.n7867 VSS.n7866 0.4505
R70744 VSS.n7865 VSS.n7279 0.4505
R70745 VSS.n7864 VSS.n7863 0.4505
R70746 VSS.n7281 VSS.n7280 0.4505
R70747 VSS.n7859 VSS.n7858 0.4505
R70748 VSS.n7857 VSS.n7283 0.4505
R70749 VSS.n9908 VSS.n4 0.4505
R70750 VSS.n9910 VSS.n9909 0.4505
R70751 VSS.n2 VSS.n1 0.4505
R70752 VSS.n9915 VSS.n9914 0.4505
R70753 VSS.n7683 VSS.n0 0.4505
R70754 VSS.n7685 VSS.n7684 0.4505
R70755 VSS.n7687 VSS.n7686 0.4505
R70756 VSS.n7680 VSS.n7679 0.4505
R70757 VSS.n7692 VSS.n7691 0.4505
R70758 VSS.n7693 VSS.n7678 0.4505
R70759 VSS.n7695 VSS.n7694 0.4505
R70760 VSS.n7676 VSS.n7675 0.4505
R70761 VSS.n7700 VSS.n7699 0.4505
R70762 VSS.n7701 VSS.n7674 0.4505
R70763 VSS.n7703 VSS.n7702 0.4505
R70764 VSS.n7672 VSS.n7671 0.4505
R70765 VSS.n7708 VSS.n7707 0.4505
R70766 VSS.n7709 VSS.n7670 0.4505
R70767 VSS.n7711 VSS.n7710 0.4505
R70768 VSS.n7668 VSS.n7667 0.4505
R70769 VSS.n7716 VSS.n7715 0.4505
R70770 VSS.n7717 VSS.n7666 0.4505
R70771 VSS.n7719 VSS.n7718 0.4505
R70772 VSS.n7664 VSS.n7663 0.4505
R70773 VSS.n7724 VSS.n7723 0.4505
R70774 VSS.n7725 VSS.n7662 0.4505
R70775 VSS.n7727 VSS.n7726 0.4505
R70776 VSS.n7660 VSS.n7659 0.4505
R70777 VSS.n7732 VSS.n7731 0.4505
R70778 VSS.n7733 VSS.n7658 0.4505
R70779 VSS.n7735 VSS.n7734 0.4505
R70780 VSS.n7656 VSS.n7655 0.4505
R70781 VSS.n7740 VSS.n7739 0.4505
R70782 VSS.n7741 VSS.n7654 0.4505
R70783 VSS.n7743 VSS.n7742 0.4505
R70784 VSS.n7652 VSS.n7651 0.4505
R70785 VSS.n7748 VSS.n7747 0.4505
R70786 VSS.n7749 VSS.n7650 0.4505
R70787 VSS.n7751 VSS.n7750 0.4505
R70788 VSS.n7648 VSS.n7647 0.4505
R70789 VSS.n7756 VSS.n7755 0.4505
R70790 VSS.n7757 VSS.n7646 0.4505
R70791 VSS.n7759 VSS.n7758 0.4505
R70792 VSS.n7644 VSS.n7643 0.4505
R70793 VSS.n7764 VSS.n7763 0.4505
R70794 VSS.n7765 VSS.n7642 0.4505
R70795 VSS.n7767 VSS.n7766 0.4505
R70796 VSS.n7640 VSS.n7639 0.4505
R70797 VSS.n7772 VSS.n7771 0.4505
R70798 VSS.n7773 VSS.n7638 0.4505
R70799 VSS.n7775 VSS.n7774 0.4505
R70800 VSS.n7636 VSS.n7635 0.4505
R70801 VSS.n7780 VSS.n7779 0.4505
R70802 VSS.n7781 VSS.n7634 0.4505
R70803 VSS.n7783 VSS.n7782 0.4505
R70804 VSS.n7632 VSS.n7631 0.4505
R70805 VSS.n7788 VSS.n7787 0.4505
R70806 VSS.n7789 VSS.n7630 0.4505
R70807 VSS.n7791 VSS.n7790 0.4505
R70808 VSS.n7628 VSS.n7627 0.4505
R70809 VSS.n7796 VSS.n7795 0.4505
R70810 VSS.n7797 VSS.n7626 0.4505
R70811 VSS.n7799 VSS.n7798 0.4505
R70812 VSS.n7624 VSS.n7623 0.4505
R70813 VSS.n7804 VSS.n7803 0.4505
R70814 VSS.n7805 VSS.n7622 0.4505
R70815 VSS.n7807 VSS.n7806 0.4505
R70816 VSS.n7620 VSS.n7619 0.4505
R70817 VSS.n7812 VSS.n7811 0.4505
R70818 VSS.n7813 VSS.n7618 0.4505
R70819 VSS.n7815 VSS.n7814 0.4505
R70820 VSS.n7616 VSS.n7615 0.4505
R70821 VSS.n7820 VSS.n7819 0.4505
R70822 VSS.n7821 VSS.n7614 0.4505
R70823 VSS.n7823 VSS.n7822 0.4505
R70824 VSS.n7612 VSS.n7611 0.4505
R70825 VSS.n7828 VSS.n7827 0.4505
R70826 VSS.n7829 VSS.n7610 0.4505
R70827 VSS.n7831 VSS.n7830 0.4505
R70828 VSS.n7608 VSS.n7607 0.4505
R70829 VSS.n7836 VSS.n7835 0.4505
R70830 VSS.n7837 VSS.n7606 0.4505
R70831 VSS.n7839 VSS.n7838 0.4505
R70832 VSS.n7604 VSS.n7603 0.4505
R70833 VSS.n7844 VSS.n7843 0.4505
R70834 VSS.n7845 VSS.n7602 0.4505
R70835 VSS.n7847 VSS.n7846 0.4505
R70836 VSS.n7600 VSS.n7599 0.4505
R70837 VSS.n7852 VSS.n7851 0.4505
R70838 VSS.n7853 VSS.n7285 0.4505
R70839 VSS.n7855 VSS.n7854 0.4505
R70840 VSS.n7877 VSS.n7876 0.4505
R70841 VSS.n7875 VSS.n7273 0.4505
R70842 VSS.n7277 VSS.n7274 0.4505
R70843 VSS.n7871 VSS.n7870 0.4505
R70844 VSS.n7869 VSS.n7276 0.4505
R70845 VSS.n7868 VSS.n7867 0.4505
R70846 VSS.n7279 VSS.n7278 0.4505
R70847 VSS.n7863 VSS.n7862 0.4505
R70848 VSS.n7861 VSS.n7281 0.4505
R70849 VSS.n7860 VSS.n7859 0.4505
R70850 VSS.n7286 VSS.n7283 0.4505
R70851 VSS.n7413 VSS.n7412 0.4505
R70852 VSS.n7411 VSS.n7410 0.4505
R70853 VSS.n7417 VSS.n7409 0.4505
R70854 VSS.n7419 VSS.n7418 0.4505
R70855 VSS.n7421 VSS.n7420 0.4505
R70856 VSS.n7407 VSS.n7406 0.4505
R70857 VSS.n7426 VSS.n7425 0.4505
R70858 VSS.n7427 VSS.n7405 0.4505
R70859 VSS.n7429 VSS.n7428 0.4505
R70860 VSS.n7403 VSS.n7402 0.4505
R70861 VSS.n7434 VSS.n7433 0.4505
R70862 VSS.n7435 VSS.n7401 0.4505
R70863 VSS.n7437 VSS.n7436 0.4505
R70864 VSS.n7399 VSS.n7398 0.4505
R70865 VSS.n7442 VSS.n7441 0.4505
R70866 VSS.n7443 VSS.n7397 0.4505
R70867 VSS.n7445 VSS.n7444 0.4505
R70868 VSS.n7395 VSS.n7394 0.4505
R70869 VSS.n7450 VSS.n7449 0.4505
R70870 VSS.n7451 VSS.n7393 0.4505
R70871 VSS.n7453 VSS.n7452 0.4505
R70872 VSS.n7391 VSS.n7390 0.4505
R70873 VSS.n7458 VSS.n7457 0.4505
R70874 VSS.n7459 VSS.n7389 0.4505
R70875 VSS.n7461 VSS.n7460 0.4505
R70876 VSS.n7387 VSS.n7386 0.4505
R70877 VSS.n7466 VSS.n7465 0.4505
R70878 VSS.n7467 VSS.n7385 0.4505
R70879 VSS.n7469 VSS.n7468 0.4505
R70880 VSS.n7383 VSS.n7382 0.4505
R70881 VSS.n7474 VSS.n7473 0.4505
R70882 VSS.n7475 VSS.n7381 0.4505
R70883 VSS.n7477 VSS.n7476 0.4505
R70884 VSS.n7379 VSS.n7378 0.4505
R70885 VSS.n7482 VSS.n7481 0.4505
R70886 VSS.n7483 VSS.n7377 0.4505
R70887 VSS.n7485 VSS.n7484 0.4505
R70888 VSS.n7375 VSS.n7374 0.4505
R70889 VSS.n7490 VSS.n7489 0.4505
R70890 VSS.n7491 VSS.n7373 0.4505
R70891 VSS.n7493 VSS.n7492 0.4505
R70892 VSS.n7371 VSS.n7370 0.4505
R70893 VSS.n7498 VSS.n7497 0.4505
R70894 VSS.n7499 VSS.n7369 0.4505
R70895 VSS.n7501 VSS.n7500 0.4505
R70896 VSS.n7367 VSS.n7366 0.4505
R70897 VSS.n7506 VSS.n7505 0.4505
R70898 VSS.n7507 VSS.n7365 0.4505
R70899 VSS.n7509 VSS.n7508 0.4505
R70900 VSS.n7363 VSS.n7362 0.4505
R70901 VSS.n7514 VSS.n7513 0.4505
R70902 VSS.n7515 VSS.n7361 0.4505
R70903 VSS.n7517 VSS.n7516 0.4505
R70904 VSS.n7359 VSS.n7358 0.4505
R70905 VSS.n7522 VSS.n7521 0.4505
R70906 VSS.n7523 VSS.n7357 0.4505
R70907 VSS.n7525 VSS.n7524 0.4505
R70908 VSS.n7355 VSS.n7354 0.4505
R70909 VSS.n7530 VSS.n7529 0.4505
R70910 VSS.n7531 VSS.n7353 0.4505
R70911 VSS.n7533 VSS.n7532 0.4505
R70912 VSS.n7351 VSS.n7350 0.4505
R70913 VSS.n7538 VSS.n7537 0.4505
R70914 VSS.n7539 VSS.n7349 0.4505
R70915 VSS.n7541 VSS.n7540 0.4505
R70916 VSS.n7347 VSS.n7346 0.4505
R70917 VSS.n7546 VSS.n7545 0.4505
R70918 VSS.n7547 VSS.n7345 0.4505
R70919 VSS.n7549 VSS.n7548 0.4505
R70920 VSS.n7343 VSS.n7342 0.4505
R70921 VSS.n7554 VSS.n7553 0.4505
R70922 VSS.n7555 VSS.n7341 0.4505
R70923 VSS.n7557 VSS.n7556 0.4505
R70924 VSS.n7339 VSS.n7338 0.4505
R70925 VSS.n7562 VSS.n7561 0.4505
R70926 VSS.n7563 VSS.n7337 0.4505
R70927 VSS.n7565 VSS.n7564 0.4505
R70928 VSS.n7335 VSS.n7334 0.4505
R70929 VSS.n7570 VSS.n7569 0.4505
R70930 VSS.n7571 VSS.n7333 0.4505
R70931 VSS.n7573 VSS.n7572 0.4505
R70932 VSS.n7331 VSS.n7330 0.4505
R70933 VSS.n7578 VSS.n7577 0.4505
R70934 VSS.n7579 VSS.n7329 0.4505
R70935 VSS.n7581 VSS.n7580 0.4505
R70936 VSS.n7327 VSS.n7326 0.4505
R70937 VSS.n7586 VSS.n7585 0.4505
R70938 VSS.n7587 VSS.n7325 0.4505
R70939 VSS.n7589 VSS.n7588 0.4505
R70940 VSS.n7291 VSS.n7289 0.4505
R70941 VSS.n7594 VSS.n7593 0.4505
R70942 VSS.n7303 VSS.n7301 0.4505
R70943 VSS.n7305 VSS.n7304 0.4505
R70944 VSS.n7299 VSS.n7298 0.4505
R70945 VSS.n7310 VSS.n7309 0.4505
R70946 VSS.n7311 VSS.n7297 0.4505
R70947 VSS.n7313 VSS.n7312 0.4505
R70948 VSS.n7295 VSS.n7294 0.4505
R70949 VSS.n7318 VSS.n7317 0.4505
R70950 VSS.n7319 VSS.n7293 0.4505
R70951 VSS.n7321 VSS.n7320 0.4505
R70952 VSS.n7290 VSS.n7288 0.4505
R70953 VSS.n7199 VSS.n7198 0.444037
R70954 VSS.n7217 VSS.n7216 0.444037
R70955 VSS.n7241 VSS.n7235 0.444037
R70956 VSS.n7085 VSS.n7084 0.444037
R70957 VSS.n7258 VSS.n2487 0.444037
R70958 VSS.n7170 VSS.n7169 0.444037
R70959 VSS.n8546 VSS.n8545 0.444037
R70960 VSS.n8809 VSS.n8808 0.444037
R70961 VSS.n8066 VSS.n8065 0.444037
R70962 VSS.n8054 VSS.n8051 0.444037
R70963 VSS.n8403 VSS.n8402 0.444037
R70964 VSS.n8847 VSS.n1321 0.444037
R70965 VSS.n8551 VSS.n8550 0.440926
R70966 VSS.n8839 VSS.n8838 0.440926
R70967 VSS.n8071 VSS.n8070 0.440926
R70968 VSS.n8047 VSS.n8046 0.440926
R70969 VSS.n8391 VSS.n1565 0.440926
R70970 VSS.n8856 VSS.n8849 0.440926
R70971 VSS.n8579 VSS.n1360 0.433833
R70972 VSS.n8827 VSS.n1360 0.433833
R70973 VSS.n8005 VSS.n1555 0.433833
R70974 VSS.n8569 VSS.n1555 0.433833
R70975 VSS.n8570 VSS.n1552 0.433833
R70976 VSS.n8570 VSS.n8569 0.433833
R70977 VSS.n8829 VSS.n8828 0.433833
R70978 VSS.n8828 VSS.n8827 0.433833
R70979 VSS.n1558 VSS.n1554 0.433833
R70980 VSS.n8569 VSS.n1554 0.433833
R70981 VSS.n2607 VSS.n1359 0.433833
R70982 VSS.n8827 VSS.n1359 0.433833
R70983 VSS.n8826 VSS.n1353 0.433833
R70984 VSS.n8827 VSS.n8826 0.433833
R70985 VSS.n8568 VSS.n8567 0.433833
R70986 VSS.n8569 VSS.n8568 0.433833
R70987 VSS.n7596 VSS.n7287 0.412146
R70988 VSS.n7597 VSS.n7282 0.412128
R70989 VSS.n7596 VSS.n7595 0.412032
R70990 VSS.n7598 VSS.n7597 0.411993
R70991 VSS.n7109 VSS.n2599 0.400007
R70992 VSS.n7115 VSS.n2594 0.400007
R70993 VSS.n7192 VSS.n7191 0.384436
R70994 VSS.n7224 VSS.n7223 0.384436
R70995 VSS.n2508 VSS.n2502 0.384436
R70996 VSS.n7095 VSS.n7089 0.384436
R70997 VSS.n7255 VSS.n7254 0.384436
R70998 VSS.n7167 VSS.n2526 0.384436
R70999 VSS.n2612 DVSS 0.37265
R71000 VSS.n7131 DVSS 0.37265
R71001 VSS.n2359 VSS.n2356 0.369923
R71002 VSS.n9449 VSS.n9446 0.369923
R71003 VSS.n2440 VSS.n2439 0.369923
R71004 VSS.n2462 VSS.n2461 0.369923
R71005 VSS.n2364 VSS.n2361 0.365885
R71006 VSS.n9444 VSS.n9441 0.365885
R71007 VSS.n8095 VSS.n2084 0.365885
R71008 VSS.n2458 VSS.n1098 0.365885
R71009 VSS.n8080 VSS.n1552 0.356041
R71010 VSS.n8580 VSS.n8579 0.356041
R71011 VSS.n2608 VSS.n2607 0.356041
R71012 VSS.n8567 VSS.n1557 0.356041
R71013 VSS.n9749 VSS.n70 0.347921
R71014 VSS.n4619 VSS.n4558 0.347921
R71015 VSS.n9695 VSS.n38 0.347921
R71016 VSS.n5062 VSS.n4382 0.347921
R71017 VSS.n5236 VSS.n5234 0.347921
R71018 VSS.n4722 VSS.n4721 0.347921
R71019 VSS.n9799 VSS.n132 0.347921
R71020 VSS.n197 VSS.n101 0.347921
R71021 VSS.n5526 VSS.n352 0.347744
R71022 VSS.n9682 VSS.n9681 0.347744
R71023 VSS.n5640 VSS.n3988 0.347744
R71024 VSS.n5267 VSS.n3945 0.347744
R71025 VSS.n6247 VSS.n3844 0.347744
R71026 VSS.n5484 VSS.n415 0.347744
R71027 VSS.n5505 VSS.n389 0.347744
R71028 VSS.n2221 VSS.n1692 0.346681
R71029 VSS.n8279 VSS.n8278 0.346681
R71030 VSS.n9568 VSS.n9567 0.346681
R71031 VSS.n8911 VSS.n8910 0.346681
R71032 VSS.n7102 VSS.n7101 0.33552
R71033 VSS.n7247 VSS.n2505 0.33552
R71034 VSS.n5793 DVSS 0.332375
R71035 VSS.n2970 DVSS 0.332375
R71036 VSS.n6295 DVSS 0.332375
R71037 VSS.n6324 DVSS 0.332375
R71038 VSS.n4103 DVSS 0.332375
R71039 VSS.n4165 DVSS 0.332375
R71040 VSS.n4325 DVSS 0.332375
R71041 VSS.n276 DVSS 0.332375
R71042 VSS.n5255 DVSS 0.332375
R71043 VSS.n283 DVSS 0.332375
R71044 VSS.n6069 DVSS 0.332375
R71045 VSS.n5945 DVSS 0.332375
R71046 VSS.n6595 DVSS 0.332375
R71047 VSS.n6630 DVSS 0.332375
R71048 VSS.n6987 DVSS 0.332375
R71049 VSS.n7016 DVSS 0.332375
R71050 DVSS VSS.n7150 0.330584
R71051 VSS.n7140 DVSS 0.330584
R71052 VSS.n6966 VSS.n6965 0.288039
R71053 VSS.n9581 VSS.n9580 0.288039
R71054 VSS.n6716 VSS.n2626 0.28237
R71055 VSS.n6940 VSS.n2760 0.28237
R71056 VSS.n6750 VSS.n2635 0.28237
R71057 VSS.n6878 VSS.n2742 0.28237
R71058 VSS.n6917 VSS.n2751 0.28237
R71059 VSS.n6698 VSS.n2622 0.28237
R71060 VSS.n2557 VSS.n2470 0.27557
R71061 VSS.n7268 VSS.n7267 0.27557
R71062 VSS.n4608 VSS.n4590 0.256847
R71063 VSS.n9825 VSS.n9824 0.256847
R71064 VSS.n7306 VSS.n7300 0.231338
R71065 VSS.n7415 VSS.n7414 0.231338
R71066 VSS.n4731 VSS.n4582 0.231338
R71067 VSS.n9794 VSS.n9793 0.231338
R71068 VSS.n8281 VSS.n1704 0.231338
R71069 VSS.n8889 VSS.n8884 0.231338
R71070 VSS.n2821 VSS.n2799 0.231338
R71071 VSS.n6678 VSS.n6673 0.231338
R71072 VSS.n3915 VSS.n3836 0.231338
R71073 VSS.n9611 VSS.n404 0.231338
R71074 VSS.n6234 VSS.n3869 0.231338
R71075 VSS.n5488 VSS.n5428 0.231338
R71076 VSS.n7874 VSS.n7272 0.231338
R71077 VSS.n9911 VSS.n3 0.231338
R71078 VSS.n7159 VSS.n7156 0.231169
R71079 VSS.n7136 VSS.n2480 0.231169
R71080 VSS.n7131 VSS.n7130 0.225249
R71081 VSS.n7046 VSS.n2612 0.225249
R71082 VSS.n1612 VSS.n1452 0.224444
R71083 VSS.n8544 VSS.n1485 0.224444
R71084 VSS.n8271 VSS.n1793 0.220739
R71085 VSS.n8274 VSS.n1754 0.220739
R71086 VSS.n8277 VSS.n1715 0.220739
R71087 VSS.n6572 VSS.n3234 0.220739
R71088 VSS.n9542 VSS.n641 0.220619
R71089 VSS.n9470 VSS.n603 0.220619
R71090 VSS.n8923 VSS.n564 0.220619
R71091 VSS.n6371 VSS.n445 0.220619
R71092 VSS.n6386 VSS.n6370 0.214786
R71093 VSS.n6556 VSS.n3269 0.214786
R71094 VSS.n6555 VSS.n3270 0.214786
R71095 VSS.n6553 VSS.n3271 0.214786
R71096 VSS.n3274 VSS.n3272 0.214786
R71097 VSS.n6549 VSS.n3275 0.214786
R71098 VSS.n6548 VSS.n3276 0.214786
R71099 VSS.n6547 VSS.n3277 0.214786
R71100 VSS.n3330 VSS.n3278 0.214786
R71101 VSS.n3331 VSS.n3329 0.214786
R71102 VSS.n6541 VSS.n3332 0.214786
R71103 VSS.n6540 VSS.n3333 0.214786
R71104 VSS.n3336 VSS.n3334 0.214786
R71105 VSS.n6536 VSS.n3337 0.214786
R71106 VSS.n6535 VSS.n3338 0.214786
R71107 VSS.n6534 VSS.n3339 0.214786
R71108 VSS.n3392 VSS.n3340 0.214786
R71109 VSS.n3393 VSS.n3391 0.214786
R71110 VSS.n6528 VSS.n3394 0.214786
R71111 VSS.n6527 VSS.n3395 0.214786
R71112 VSS.n3398 VSS.n3396 0.214786
R71113 VSS.n6523 VSS.n3399 0.214786
R71114 VSS.n6522 VSS.n3400 0.214786
R71115 VSS.n6521 VSS.n3401 0.214786
R71116 VSS.n3404 VSS.n3402 0.214786
R71117 VSS.n6517 VSS.n3405 0.214786
R71118 VSS.n6516 VSS.n3406 0.214786
R71119 VSS.n6515 VSS.n3407 0.214786
R71120 VSS.n3410 VSS.n3408 0.214786
R71121 VSS.n6511 VSS.n3411 0.214786
R71122 VSS.n6510 VSS.n3412 0.214786
R71123 VSS.n6509 VSS.n3413 0.214786
R71124 VSS.n3466 VSS.n3414 0.214786
R71125 VSS.n3467 VSS.n3465 0.214786
R71126 VSS.n6503 VSS.n3468 0.214786
R71127 VSS.n6502 VSS.n3469 0.214786
R71128 VSS.n3472 VSS.n3470 0.214786
R71129 VSS.n6498 VSS.n3473 0.214786
R71130 VSS.n6497 VSS.n3474 0.214786
R71131 VSS.n6496 VSS.n3475 0.214786
R71132 VSS.n3478 VSS.n3476 0.214786
R71133 VSS.n6492 VSS.n3479 0.214786
R71134 VSS.n6491 VSS.n3480 0.214786
R71135 VSS.n6490 VSS.n3481 0.214786
R71136 VSS.n3484 VSS.n3482 0.214786
R71137 VSS.n6486 VSS.n3485 0.214786
R71138 VSS.n6485 VSS.n3486 0.214786
R71139 VSS.n6484 VSS.n3487 0.214786
R71140 VSS.n6483 VSS.n3488 0.214786
R71141 VSS.n6482 VSS.n3489 0.214786
R71142 VSS.n6479 VSS.n3490 0.214786
R71143 VSS.n6477 VSS.n3491 0.214786
R71144 VSS.n6476 VSS.n3492 0.214786
R71145 VSS.n6475 VSS.n3493 0.214786
R71146 VSS.n6473 VSS.n3494 0.214786
R71147 VSS.n3497 VSS.n3495 0.214786
R71148 VSS.n6469 VSS.n3498 0.214786
R71149 VSS.n6468 VSS.n3499 0.214786
R71150 VSS.n6467 VSS.n3500 0.214786
R71151 VSS.n3503 VSS.n3501 0.214786
R71152 VSS.n6463 VSS.n3504 0.214786
R71153 VSS.n6462 VSS.n3505 0.214786
R71154 VSS.n6461 VSS.n3506 0.214786
R71155 VSS.n3509 VSS.n3507 0.214786
R71156 VSS.n6457 VSS.n3510 0.214786
R71157 VSS.n6456 VSS.n3511 0.214786
R71158 VSS.n6455 VSS.n3512 0.214786
R71159 VSS.n3565 VSS.n3513 0.214786
R71160 VSS.n3566 VSS.n3564 0.214786
R71161 VSS.n6449 VSS.n3567 0.214786
R71162 VSS.n6448 VSS.n3568 0.214786
R71163 VSS.n3571 VSS.n3569 0.214786
R71164 VSS.n6444 VSS.n3572 0.214786
R71165 VSS.n6443 VSS.n3573 0.214786
R71166 VSS.n6442 VSS.n3574 0.214786
R71167 VSS.n3577 VSS.n3575 0.214786
R71168 VSS.n6438 VSS.n3578 0.214786
R71169 VSS.n6437 VSS.n3579 0.214786
R71170 VSS.n6436 VSS.n3580 0.214786
R71171 VSS.n3583 VSS.n3581 0.214786
R71172 VSS.n6432 VSS.n3584 0.214786
R71173 VSS.n6431 VSS.n3585 0.214786
R71174 VSS.n6430 VSS.n3586 0.214786
R71175 VSS.n3629 VSS.n3587 0.214786
R71176 VSS.n3631 VSS.n3630 0.214786
R71177 VSS.n3632 VSS.n3628 0.214786
R71178 VSS.n6412 VSS.n3633 0.214786
R71179 VSS.n6411 VSS.n3634 0.214786
R71180 VSS.n6410 VSS.n3635 0.214786
R71181 VSS.n3638 VSS.n3636 0.214786
R71182 VSS.n6406 VSS.n3639 0.214786
R71183 VSS.n6405 VSS.n3640 0.214786
R71184 VSS.n6362 VSS.n3641 0.214786
R71185 VSS.n6363 VSS.n6361 0.214786
R71186 VSS.n6394 VSS.n6364 0.214786
R71187 VSS.n6393 VSS.n6365 0.214786
R71188 VSS.n6392 VSS.n6366 0.214786
R71189 VSS.n6389 VSS.n6367 0.214786
R71190 VSS.n6388 VSS.n6368 0.214786
R71191 VSS.n6387 VSS.n6369 0.214786
R71192 VSS.n2244 VSS.n2231 0.214786
R71193 VSS.n2246 VSS.n2229 0.214786
R71194 VSS.n2249 VSS.n2248 0.214786
R71195 VSS.n2250 VSS.n2228 0.214786
R71196 VSS.n2253 VSS.n2252 0.214786
R71197 VSS.n2251 VSS.n2225 0.214786
R71198 VSS.n2257 VSS.n2226 0.214786
R71199 VSS.n2259 VSS.n2224 0.214786
R71200 VSS.n2262 VSS.n2261 0.214786
R71201 VSS.n2263 VSS.n2223 0.214786
R71202 VSS.n2267 VSS.n2264 0.214786
R71203 VSS.n2266 VSS.n2265 0.214786
R71204 VSS.n2133 VSS.n2132 0.214786
R71205 VSS.n7949 VSS.n7948 0.214786
R71206 VSS.n7953 VSS.n2130 0.214786
R71207 VSS.n7955 VSS.n2128 0.214786
R71208 VSS.n7958 VSS.n7957 0.214786
R71209 VSS.n7959 VSS.n2127 0.214786
R71210 VSS.n7998 VSS.n7960 0.214786
R71211 VSS.n7997 VSS.n7961 0.214786
R71212 VSS.n7996 VSS.n7962 0.214786
R71213 VSS.n7965 VSS.n7963 0.214786
R71214 VSS.n7992 VSS.n7966 0.214786
R71215 VSS.n7991 VSS.n7967 0.214786
R71216 VSS.n7990 VSS.n7968 0.214786
R71217 VSS.n7971 VSS.n7969 0.214786
R71218 VSS.n7986 VSS.n7972 0.214786
R71219 VSS.n7985 VSS.n7973 0.214786
R71220 VSS.n7984 VSS.n7974 0.214786
R71221 VSS.n7976 VSS.n7975 0.214786
R71222 VSS.n7980 VSS.n7977 0.214786
R71223 VSS.n7979 VSS.n7978 0.214786
R71224 VSS.n1522 VSS.n1521 0.214786
R71225 VSS.n8638 VSS.n8637 0.214786
R71226 VSS.n8639 VSS.n1520 0.214786
R71227 VSS.n8641 VSS.n8640 0.214786
R71228 VSS.n1517 VSS.n1516 0.214786
R71229 VSS.n8646 VSS.n8645 0.214786
R71230 VSS.n8648 VSS.n1515 0.214786
R71231 VSS.n8650 VSS.n8649 0.214786
R71232 VSS.n1513 VSS.n1512 0.214786
R71233 VSS.n8655 VSS.n8654 0.214786
R71234 VSS.n8656 VSS.n1511 0.214786
R71235 VSS.n8658 VSS.n8657 0.214786
R71236 VSS.n1509 VSS.n1508 0.214786
R71237 VSS.n8663 VSS.n8662 0.214786
R71238 VSS.n8664 VSS.n1507 0.214786
R71239 VSS.n8666 VSS.n8665 0.214786
R71240 VSS.n1476 VSS.n1475 0.214786
R71241 VSS.n8689 VSS.n8688 0.214786
R71242 VSS.n8690 VSS.n1474 0.214786
R71243 VSS.n8692 VSS.n8691 0.214786
R71244 VSS.n1443 VSS.n1442 0.214786
R71245 VSS.n8715 VSS.n8714 0.214786
R71246 VSS.n8716 VSS.n1441 0.214786
R71247 VSS.n8718 VSS.n8717 0.214786
R71248 VSS.n1439 VSS.n1438 0.214786
R71249 VSS.n8723 VSS.n8722 0.214786
R71250 VSS.n8724 VSS.n1437 0.214786
R71251 VSS.n8726 VSS.n8725 0.214786
R71252 VSS.n1435 VSS.n1434 0.214786
R71253 VSS.n8731 VSS.n8730 0.214786
R71254 VSS.n8735 VSS.n8734 0.214786
R71255 VSS.n8733 VSS.n1432 0.214786
R71256 VSS.n8739 VSS.n1431 0.214786
R71257 VSS.n8741 VSS.n8740 0.214786
R71258 VSS.n8742 VSS.n1430 0.214786
R71259 VSS.n8793 VSS.n8743 0.214786
R71260 VSS.n8792 VSS.n8744 0.214786
R71261 VSS.n8790 VSS.n8745 0.214786
R71262 VSS.n8748 VSS.n8746 0.214786
R71263 VSS.n8786 VSS.n8749 0.214786
R71264 VSS.n8785 VSS.n8750 0.214786
R71265 VSS.n8784 VSS.n8751 0.214786
R71266 VSS.n8754 VSS.n8752 0.214786
R71267 VSS.n8780 VSS.n8755 0.214786
R71268 VSS.n8779 VSS.n8756 0.214786
R71269 VSS.n8778 VSS.n8757 0.214786
R71270 VSS.n8760 VSS.n8758 0.214786
R71271 VSS.n8774 VSS.n8761 0.214786
R71272 VSS.n8773 VSS.n8762 0.214786
R71273 VSS.n8772 VSS.n8763 0.214786
R71274 VSS.n8770 VSS.n8764 0.214786
R71275 VSS.n8768 VSS.n8766 0.214786
R71276 VSS.n8765 VSS.n1140 0.214786
R71277 VSS.n8960 VSS.n1141 0.214786
R71278 VSS.n8958 VSS.n1142 0.214786
R71279 VSS.n1145 VSS.n1143 0.214786
R71280 VSS.n8954 VSS.n1146 0.214786
R71281 VSS.n8953 VSS.n1147 0.214786
R71282 VSS.n8952 VSS.n1148 0.214786
R71283 VSS.n8914 VSS.n1149 0.214786
R71284 VSS.n8915 VSS.n8913 0.214786
R71285 VSS.n8946 VSS.n8916 0.214786
R71286 VSS.n8945 VSS.n8917 0.214786
R71287 VSS.n8944 VSS.n8918 0.214786
R71288 VSS.n8941 VSS.n8919 0.214786
R71289 VSS.n8940 VSS.n8920 0.214786
R71290 VSS.n8939 VSS.n8921 0.214786
R71291 VSS.n8938 VSS.n8922 0.214786
R71292 VSS.n7913 VSS.n7899 0.214786
R71293 VSS.n7916 VSS.n7915 0.214786
R71294 VSS.n7917 VSS.n7898 0.214786
R71295 VSS.n7919 VSS.n7918 0.214786
R71296 VSS.n7896 VSS.n7895 0.214786
R71297 VSS.n7924 VSS.n7923 0.214786
R71298 VSS.n7925 VSS.n7894 0.214786
R71299 VSS.n7927 VSS.n7926 0.214786
R71300 VSS.n2141 VSS.n2140 0.214786
R71301 VSS.n7934 VSS.n7933 0.214786
R71302 VSS.n7935 VSS.n2139 0.214786
R71303 VSS.n7938 VSS.n7937 0.214786
R71304 VSS.n7936 VSS.n2137 0.214786
R71305 VSS.n7942 VSS.n2136 0.214786
R71306 VSS.n7945 VSS.n7944 0.214786
R71307 VSS.n2034 VSS.n2033 0.214786
R71308 VSS.n8106 VSS.n8105 0.214786
R71309 VSS.n8107 VSS.n2032 0.214786
R71310 VSS.n8109 VSS.n8108 0.214786
R71311 VSS.n2030 VSS.n2029 0.214786
R71312 VSS.n8114 VSS.n8113 0.214786
R71313 VSS.n8115 VSS.n2028 0.214786
R71314 VSS.n8117 VSS.n8116 0.214786
R71315 VSS.n2026 VSS.n2025 0.214786
R71316 VSS.n8122 VSS.n8121 0.214786
R71317 VSS.n8123 VSS.n2024 0.214786
R71318 VSS.n8125 VSS.n8124 0.214786
R71319 VSS.n2022 VSS.n2021 0.214786
R71320 VSS.n8131 VSS.n8130 0.214786
R71321 VSS.n8132 VSS.n2020 0.214786
R71322 VSS.n8134 VSS.n8133 0.214786
R71323 VSS.n8135 VSS.n2019 0.214786
R71324 VSS.n8138 VSS.n8137 0.214786
R71325 VSS.n8139 VSS.n2018 0.214786
R71326 VSS.n8148 VSS.n8140 0.214786
R71327 VSS.n8147 VSS.n8141 0.214786
R71328 VSS.n8146 VSS.n8142 0.214786
R71329 VSS.n8144 VSS.n8143 0.214786
R71330 VSS.n9170 VSS.n946 0.214786
R71331 VSS.n9169 VSS.n947 0.214786
R71332 VSS.n9168 VSS.n948 0.214786
R71333 VSS.n951 VSS.n949 0.214786
R71334 VSS.n9164 VSS.n952 0.214786
R71335 VSS.n9163 VSS.n953 0.214786
R71336 VSS.n9162 VSS.n954 0.214786
R71337 VSS.n957 VSS.n955 0.214786
R71338 VSS.n9158 VSS.n958 0.214786
R71339 VSS.n9157 VSS.n959 0.214786
R71340 VSS.n976 VSS.n960 0.214786
R71341 VSS.n9118 VSS.n977 0.214786
R71342 VSS.n9117 VSS.n978 0.214786
R71343 VSS.n9116 VSS.n979 0.214786
R71344 VSS.n997 VSS.n980 0.214786
R71345 VSS.n9077 VSS.n998 0.214786
R71346 VSS.n9076 VSS.n999 0.214786
R71347 VSS.n9075 VSS.n1000 0.214786
R71348 VSS.n1003 VSS.n1001 0.214786
R71349 VSS.n9071 VSS.n1004 0.214786
R71350 VSS.n9070 VSS.n1005 0.214786
R71351 VSS.n9069 VSS.n1006 0.214786
R71352 VSS.n1009 VSS.n1007 0.214786
R71353 VSS.n9065 VSS.n1010 0.214786
R71354 VSS.n9063 VSS.n1012 0.214786
R71355 VSS.n1015 VSS.n1013 0.214786
R71356 VSS.n9059 VSS.n1016 0.214786
R71357 VSS.n9058 VSS.n1017 0.214786
R71358 VSS.n9057 VSS.n1018 0.214786
R71359 VSS.n1057 VSS.n1019 0.214786
R71360 VSS.n1058 VSS.n1056 0.214786
R71361 VSS.n9037 VSS.n1059 0.214786
R71362 VSS.n9036 VSS.n1060 0.214786
R71363 VSS.n9035 VSS.n1061 0.214786
R71364 VSS.n1064 VSS.n1062 0.214786
R71365 VSS.n9031 VSS.n1065 0.214786
R71366 VSS.n9030 VSS.n1066 0.214786
R71367 VSS.n9029 VSS.n1067 0.214786
R71368 VSS.n1070 VSS.n1068 0.214786
R71369 VSS.n9025 VSS.n1071 0.214786
R71370 VSS.n9024 VSS.n1072 0.214786
R71371 VSS.n9023 VSS.n1073 0.214786
R71372 VSS.n1076 VSS.n1074 0.214786
R71373 VSS.n9019 VSS.n1077 0.214786
R71374 VSS.n9018 VSS.n1078 0.214786
R71375 VSS.n8996 VSS.n1079 0.214786
R71376 VSS.n8998 VSS.n8997 0.214786
R71377 VSS.n8999 VSS.n719 0.214786
R71378 VSS.n9508 VSS.n9507 0.214786
R71379 VSS.n722 VSS.n720 0.214786
R71380 VSS.n9503 VSS.n725 0.214786
R71381 VSS.n9502 VSS.n726 0.214786
R71382 VSS.n9501 VSS.n727 0.214786
R71383 VSS.n9459 VSS.n728 0.214786
R71384 VSS.n9495 VSS.n9460 0.214786
R71385 VSS.n9494 VSS.n9461 0.214786
R71386 VSS.n9464 VSS.n9462 0.214786
R71387 VSS.n9490 VSS.n9465 0.214786
R71388 VSS.n9489 VSS.n9466 0.214786
R71389 VSS.n9488 VSS.n9467 0.214786
R71390 VSS.n9486 VSS.n9468 0.214786
R71391 VSS.n9485 VSS.n9469 0.214786
R71392 VSS.n9545 VSS.n9541 0.214786
R71393 VSS.n8256 VSS.n1829 0.214786
R71394 VSS.n8255 VSS.n1830 0.214786
R71395 VSS.n8253 VSS.n1831 0.214786
R71396 VSS.n1834 VSS.n1832 0.214786
R71397 VSS.n8249 VSS.n1835 0.214786
R71398 VSS.n8248 VSS.n1836 0.214786
R71399 VSS.n8247 VSS.n1837 0.214786
R71400 VSS.n1870 VSS.n1838 0.214786
R71401 VSS.n1873 VSS.n1872 0.214786
R71402 VSS.n1874 VSS.n1869 0.214786
R71403 VSS.n8241 VSS.n1875 0.214786
R71404 VSS.n8240 VSS.n1876 0.214786
R71405 VSS.n8239 VSS.n1877 0.214786
R71406 VSS.n2134 VSS.n1878 0.214786
R71407 VSS.n8234 VSS.n1882 0.214786
R71408 VSS.n8233 VSS.n1883 0.214786
R71409 VSS.n1931 VSS.n1884 0.214786
R71410 VSS.n1932 VSS.n1930 0.214786
R71411 VSS.n8222 VSS.n1933 0.214786
R71412 VSS.n8221 VSS.n1934 0.214786
R71413 VSS.n8220 VSS.n1935 0.214786
R71414 VSS.n1938 VSS.n1936 0.214786
R71415 VSS.n8216 VSS.n1939 0.214786
R71416 VSS.n8215 VSS.n1940 0.214786
R71417 VSS.n8214 VSS.n1941 0.214786
R71418 VSS.n1944 VSS.n1942 0.214786
R71419 VSS.n8210 VSS.n1945 0.214786
R71420 VSS.n8209 VSS.n1946 0.214786
R71421 VSS.n8208 VSS.n1947 0.214786
R71422 VSS.n1950 VSS.n1948 0.214786
R71423 VSS.n8204 VSS.n1951 0.214786
R71424 VSS.n8203 VSS.n1952 0.214786
R71425 VSS.n8187 VSS.n1953 0.214786
R71426 VSS.n8188 VSS.n8186 0.214786
R71427 VSS.n8192 VSS.n8189 0.214786
R71428 VSS.n8191 VSS.n8190 0.214786
R71429 VSS.n939 VSS.n938 0.214786
R71430 VSS.n9176 VSS.n9175 0.214786
R71431 VSS.n9178 VSS.n936 0.214786
R71432 VSS.n9180 VSS.n9179 0.214786
R71433 VSS.n934 VSS.n933 0.214786
R71434 VSS.n9185 VSS.n9184 0.214786
R71435 VSS.n9186 VSS.n932 0.214786
R71436 VSS.n9188 VSS.n9187 0.214786
R71437 VSS.n930 VSS.n929 0.214786
R71438 VSS.n9193 VSS.n9192 0.214786
R71439 VSS.n9194 VSS.n928 0.214786
R71440 VSS.n9196 VSS.n9195 0.214786
R71441 VSS.n900 VSS.n899 0.214786
R71442 VSS.n9226 VSS.n9225 0.214786
R71443 VSS.n9227 VSS.n898 0.214786
R71444 VSS.n9229 VSS.n9228 0.214786
R71445 VSS.n872 VSS.n871 0.214786
R71446 VSS.n9259 VSS.n9258 0.214786
R71447 VSS.n9260 VSS.n870 0.214786
R71448 VSS.n9262 VSS.n9261 0.214786
R71449 VSS.n868 VSS.n867 0.214786
R71450 VSS.n9267 VSS.n9266 0.214786
R71451 VSS.n9268 VSS.n866 0.214786
R71452 VSS.n9270 VSS.n9269 0.214786
R71453 VSS.n864 VSS.n863 0.214786
R71454 VSS.n9275 VSS.n9274 0.214786
R71455 VSS.n9278 VSS.n9277 0.214786
R71456 VSS.n859 VSS.n858 0.214786
R71457 VSS.n9283 VSS.n9282 0.214786
R71458 VSS.n9284 VSS.n857 0.214786
R71459 VSS.n9286 VSS.n9285 0.214786
R71460 VSS.n830 VSS.n829 0.214786
R71461 VSS.n9317 VSS.n9316 0.214786
R71462 VSS.n9318 VSS.n828 0.214786
R71463 VSS.n9320 VSS.n9319 0.214786
R71464 VSS.n826 VSS.n825 0.214786
R71465 VSS.n9325 VSS.n9324 0.214786
R71466 VSS.n9326 VSS.n824 0.214786
R71467 VSS.n9328 VSS.n9327 0.214786
R71468 VSS.n822 VSS.n821 0.214786
R71469 VSS.n9333 VSS.n9332 0.214786
R71470 VSS.n9334 VSS.n820 0.214786
R71471 VSS.n9337 VSS.n9336 0.214786
R71472 VSS.n9335 VSS.n818 0.214786
R71473 VSS.n9341 VSS.n817 0.214786
R71474 VSS.n9343 VSS.n9342 0.214786
R71475 VSS.n9344 VSS.n816 0.214786
R71476 VSS.n9351 VSS.n9345 0.214786
R71477 VSS.n9350 VSS.n9346 0.214786
R71478 VSS.n9348 VSS.n717 0.214786
R71479 VSS.n9512 VSS.n9511 0.214786
R71480 VSS.n714 VSS.n713 0.214786
R71481 VSS.n9518 VSS.n9517 0.214786
R71482 VSS.n9519 VSS.n712 0.214786
R71483 VSS.n9521 VSS.n9520 0.214786
R71484 VSS.n684 VSS.n683 0.214786
R71485 VSS.n9529 VSS.n9528 0.214786
R71486 VSS.n9530 VSS.n682 0.214786
R71487 VSS.n9533 VSS.n9532 0.214786
R71488 VSS.n9531 VSS.n679 0.214786
R71489 VSS.n9537 VSS.n680 0.214786
R71490 VSS.n9539 VSS.n9538 0.214786
R71491 VSS.n9540 VSS.n678 0.214786
R71492 VSS.n9544 VSS.n9543 0.214786
R71493 VSS.n9546 VSS.n9545 0.214786
R71494 VSS.n1828 VSS.n1805 0.214786
R71495 VSS.n8257 VSS.n8256 0.214786
R71496 VSS.n8255 VSS.n8254 0.214786
R71497 VSS.n8253 VSS.n8252 0.214786
R71498 VSS.n8251 VSS.n1832 0.214786
R71499 VSS.n8250 VSS.n8249 0.214786
R71500 VSS.n8248 VSS.n1833 0.214786
R71501 VSS.n8247 VSS.n8246 0.214786
R71502 VSS.n1851 VSS.n1838 0.214786
R71503 VSS.n1872 VSS.n1871 0.214786
R71504 VSS.n1869 VSS.n1867 0.214786
R71505 VSS.n8242 VSS.n8241 0.214786
R71506 VSS.n8240 VSS.n1868 0.214786
R71507 VSS.n8239 VSS.n8238 0.214786
R71508 VSS.n8237 VSS.n1878 0.214786
R71509 VSS.n8235 VSS.n8234 0.214786
R71510 VSS.n8233 VSS.n8232 0.214786
R71511 VSS.n1885 VSS.n1884 0.214786
R71512 VSS.n1930 VSS.n1910 0.214786
R71513 VSS.n8223 VSS.n8222 0.214786
R71514 VSS.n8221 VSS.n1929 0.214786
R71515 VSS.n8220 VSS.n8219 0.214786
R71516 VSS.n8218 VSS.n1936 0.214786
R71517 VSS.n8217 VSS.n8216 0.214786
R71518 VSS.n8215 VSS.n1937 0.214786
R71519 VSS.n8214 VSS.n8213 0.214786
R71520 VSS.n8212 VSS.n1942 0.214786
R71521 VSS.n8211 VSS.n8210 0.214786
R71522 VSS.n8209 VSS.n1943 0.214786
R71523 VSS.n8208 VSS.n8207 0.214786
R71524 VSS.n8206 VSS.n1948 0.214786
R71525 VSS.n8205 VSS.n8204 0.214786
R71526 VSS.n8203 VSS.n8202 0.214786
R71527 VSS.n1954 VSS.n1953 0.214786
R71528 VSS.n8186 VSS.n8166 0.214786
R71529 VSS.n8193 VSS.n8192 0.214786
R71530 VSS.n8191 VSS.n8185 0.214786
R71531 VSS.n941 VSS.n939 0.214786
R71532 VSS.n9175 VSS.n9174 0.214786
R71533 VSS.n936 VSS.n935 0.214786
R71534 VSS.n9181 VSS.n9180 0.214786
R71535 VSS.n9182 VSS.n934 0.214786
R71536 VSS.n9184 VSS.n9183 0.214786
R71537 VSS.n932 VSS.n931 0.214786
R71538 VSS.n9189 VSS.n9188 0.214786
R71539 VSS.n9190 VSS.n930 0.214786
R71540 VSS.n9192 VSS.n9191 0.214786
R71541 VSS.n928 VSS.n916 0.214786
R71542 VSS.n9197 VSS.n9196 0.214786
R71543 VSS.n901 VSS.n900 0.214786
R71544 VSS.n9225 VSS.n9224 0.214786
R71545 VSS.n898 VSS.n887 0.214786
R71546 VSS.n9230 VSS.n9229 0.214786
R71547 VSS.n873 VSS.n872 0.214786
R71548 VSS.n9258 VSS.n9257 0.214786
R71549 VSS.n870 VSS.n869 0.214786
R71550 VSS.n9263 VSS.n9262 0.214786
R71551 VSS.n9264 VSS.n868 0.214786
R71552 VSS.n9266 VSS.n9265 0.214786
R71553 VSS.n866 VSS.n865 0.214786
R71554 VSS.n9271 VSS.n9270 0.214786
R71555 VSS.n9272 VSS.n864 0.214786
R71556 VSS.n9274 VSS.n9273 0.214786
R71557 VSS.n9279 VSS.n9278 0.214786
R71558 VSS.n9280 VSS.n859 0.214786
R71559 VSS.n9282 VSS.n9281 0.214786
R71560 VSS.n857 VSS.n845 0.214786
R71561 VSS.n9287 VSS.n9286 0.214786
R71562 VSS.n9298 VSS.n830 0.214786
R71563 VSS.n9316 VSS.n9315 0.214786
R71564 VSS.n828 VSS.n827 0.214786
R71565 VSS.n9321 VSS.n9320 0.214786
R71566 VSS.n9322 VSS.n826 0.214786
R71567 VSS.n9324 VSS.n9323 0.214786
R71568 VSS.n824 VSS.n823 0.214786
R71569 VSS.n9329 VSS.n9328 0.214786
R71570 VSS.n9330 VSS.n822 0.214786
R71571 VSS.n9332 VSS.n9331 0.214786
R71572 VSS.n820 VSS.n819 0.214786
R71573 VSS.n9338 VSS.n9337 0.214786
R71574 VSS.n9339 VSS.n818 0.214786
R71575 VSS.n9341 VSS.n9340 0.214786
R71576 VSS.n9342 VSS.n782 0.214786
R71577 VSS.n816 VSS.n795 0.214786
R71578 VSS.n9352 VSS.n9351 0.214786
R71579 VSS.n9350 VSS.n9349 0.214786
R71580 VSS.n9348 VSS.n9347 0.214786
R71581 VSS.n9513 VSS.n9512 0.214786
R71582 VSS.n9514 VSS.n714 0.214786
R71583 VSS.n9517 VSS.n9516 0.214786
R71584 VSS.n9515 VSS.n712 0.214786
R71585 VSS.n9522 VSS.n9521 0.214786
R71586 VSS.n9523 VSS.n684 0.214786
R71587 VSS.n9528 VSS.n9527 0.214786
R71588 VSS.n682 VSS.n681 0.214786
R71589 VSS.n9534 VSS.n9533 0.214786
R71590 VSS.n9535 VSS.n679 0.214786
R71591 VSS.n9537 VSS.n9536 0.214786
R71592 VSS.n9538 VSS.n643 0.214786
R71593 VSS.n678 VSS.n655 0.214786
R71594 VSS.n9472 VSS.n9471 0.214786
R71595 VSS.n9485 VSS.n9484 0.214786
R71596 VSS.n9486 VSS.n616 0.214786
R71597 VSS.n9488 VSS.n9487 0.214786
R71598 VSS.n9489 VSS.n9463 0.214786
R71599 VSS.n9491 VSS.n9490 0.214786
R71600 VSS.n9492 VSS.n9462 0.214786
R71601 VSS.n9494 VSS.n9493 0.214786
R71602 VSS.n9496 VSS.n9495 0.214786
R71603 VSS.n742 VSS.n728 0.214786
R71604 VSS.n9501 VSS.n9500 0.214786
R71605 VSS.n9502 VSS.n724 0.214786
R71606 VSS.n9504 VSS.n9503 0.214786
R71607 VSS.n9505 VSS.n722 0.214786
R71608 VSS.n9507 VSS.n9506 0.214786
R71609 VSS.n9000 VSS.n8999 0.214786
R71610 VSS.n8998 VSS.n8985 0.214786
R71611 VSS.n8972 VSS.n1079 0.214786
R71612 VSS.n9018 VSS.n9017 0.214786
R71613 VSS.n9020 VSS.n9019 0.214786
R71614 VSS.n9021 VSS.n1074 0.214786
R71615 VSS.n9023 VSS.n9022 0.214786
R71616 VSS.n9024 VSS.n1069 0.214786
R71617 VSS.n9026 VSS.n9025 0.214786
R71618 VSS.n9027 VSS.n1068 0.214786
R71619 VSS.n9029 VSS.n9028 0.214786
R71620 VSS.n9030 VSS.n1063 0.214786
R71621 VSS.n9032 VSS.n9031 0.214786
R71622 VSS.n9033 VSS.n1062 0.214786
R71623 VSS.n9035 VSS.n9034 0.214786
R71624 VSS.n9036 VSS.n1055 0.214786
R71625 VSS.n9038 VSS.n9037 0.214786
R71626 VSS.n1056 VSS.n1044 0.214786
R71627 VSS.n9054 VSS.n1019 0.214786
R71628 VSS.n9057 VSS.n9056 0.214786
R71629 VSS.n9058 VSS.n1014 0.214786
R71630 VSS.n9060 VSS.n9059 0.214786
R71631 VSS.n9061 VSS.n1013 0.214786
R71632 VSS.n9063 VSS.n9062 0.214786
R71633 VSS.n9066 VSS.n9065 0.214786
R71634 VSS.n9067 VSS.n1007 0.214786
R71635 VSS.n9069 VSS.n9068 0.214786
R71636 VSS.n9070 VSS.n1002 0.214786
R71637 VSS.n9072 VSS.n9071 0.214786
R71638 VSS.n9073 VSS.n1001 0.214786
R71639 VSS.n9075 VSS.n9074 0.214786
R71640 VSS.n9076 VSS.n996 0.214786
R71641 VSS.n9078 VSS.n9077 0.214786
R71642 VSS.n982 VSS.n980 0.214786
R71643 VSS.n9116 VSS.n9115 0.214786
R71644 VSS.n9117 VSS.n975 0.214786
R71645 VSS.n9119 VSS.n9118 0.214786
R71646 VSS.n961 VSS.n960 0.214786
R71647 VSS.n9157 VSS.n9156 0.214786
R71648 VSS.n9159 VSS.n9158 0.214786
R71649 VSS.n9160 VSS.n955 0.214786
R71650 VSS.n9162 VSS.n9161 0.214786
R71651 VSS.n9163 VSS.n950 0.214786
R71652 VSS.n9165 VSS.n9164 0.214786
R71653 VSS.n9166 VSS.n949 0.214786
R71654 VSS.n9168 VSS.n9167 0.214786
R71655 VSS.n9169 VSS.n944 0.214786
R71656 VSS.n9171 VSS.n9170 0.214786
R71657 VSS.n8144 VSS.n943 0.214786
R71658 VSS.n8146 VSS.n8145 0.214786
R71659 VSS.n8147 VSS.n2017 0.214786
R71660 VSS.n8149 VSS.n8148 0.214786
R71661 VSS.n2018 VSS.n2016 0.214786
R71662 VSS.n8137 VSS.n8136 0.214786
R71663 VSS.n8135 VSS.n1994 0.214786
R71664 VSS.n8134 VSS.n1981 0.214786
R71665 VSS.n8128 VSS.n2020 0.214786
R71666 VSS.n8130 VSS.n8129 0.214786
R71667 VSS.n8127 VSS.n2022 0.214786
R71668 VSS.n8126 VSS.n8125 0.214786
R71669 VSS.n2024 VSS.n2023 0.214786
R71670 VSS.n8121 VSS.n8120 0.214786
R71671 VSS.n8119 VSS.n2026 0.214786
R71672 VSS.n8118 VSS.n8117 0.214786
R71673 VSS.n2028 VSS.n2027 0.214786
R71674 VSS.n8113 VSS.n8112 0.214786
R71675 VSS.n8111 VSS.n2030 0.214786
R71676 VSS.n8110 VSS.n8109 0.214786
R71677 VSS.n2047 VSS.n2032 0.214786
R71678 VSS.n8105 VSS.n8104 0.214786
R71679 VSS.n8098 VSS.n2034 0.214786
R71680 VSS.n7944 VSS.n2080 0.214786
R71681 VSS.n7942 VSS.n7941 0.214786
R71682 VSS.n7940 VSS.n2137 0.214786
R71683 VSS.n7939 VSS.n7938 0.214786
R71684 VSS.n2139 VSS.n2138 0.214786
R71685 VSS.n7933 VSS.n7932 0.214786
R71686 VSS.n2167 VSS.n2141 0.214786
R71687 VSS.n7928 VSS.n7927 0.214786
R71688 VSS.n7894 VSS.n7893 0.214786
R71689 VSS.n7923 VSS.n7922 0.214786
R71690 VSS.n7921 VSS.n7896 0.214786
R71691 VSS.n7920 VSS.n7919 0.214786
R71692 VSS.n7898 VSS.n7897 0.214786
R71693 VSS.n7915 VSS.n7914 0.214786
R71694 VSS.n7913 VSS.n7912 0.214786
R71695 VSS.n7900 VSS.n1766 0.214786
R71696 VSS.n8925 VSS.n8924 0.214786
R71697 VSS.n8938 VSS.n8937 0.214786
R71698 VSS.n8939 VSS.n578 0.214786
R71699 VSS.n8940 VSS.n566 0.214786
R71700 VSS.n8942 VSS.n8941 0.214786
R71701 VSS.n8944 VSS.n8943 0.214786
R71702 VSS.n8945 VSS.n8912 0.214786
R71703 VSS.n8947 VSS.n8946 0.214786
R71704 VSS.n8913 VSS.n1225 0.214786
R71705 VSS.n1152 VSS.n1149 0.214786
R71706 VSS.n8952 VSS.n8951 0.214786
R71707 VSS.n8953 VSS.n1144 0.214786
R71708 VSS.n8955 VSS.n8954 0.214786
R71709 VSS.n8956 VSS.n1143 0.214786
R71710 VSS.n8958 VSS.n8957 0.214786
R71711 VSS.n8961 VSS.n8960 0.214786
R71712 VSS.n1140 VSS.n1102 0.214786
R71713 VSS.n8768 VSS.n8767 0.214786
R71714 VSS.n8770 VSS.n8769 0.214786
R71715 VSS.n8772 VSS.n8771 0.214786
R71716 VSS.n8773 VSS.n8759 0.214786
R71717 VSS.n8775 VSS.n8774 0.214786
R71718 VSS.n8776 VSS.n8758 0.214786
R71719 VSS.n8778 VSS.n8777 0.214786
R71720 VSS.n8779 VSS.n8753 0.214786
R71721 VSS.n8781 VSS.n8780 0.214786
R71722 VSS.n8782 VSS.n8752 0.214786
R71723 VSS.n8784 VSS.n8783 0.214786
R71724 VSS.n8785 VSS.n8747 0.214786
R71725 VSS.n8787 VSS.n8786 0.214786
R71726 VSS.n8788 VSS.n8746 0.214786
R71727 VSS.n8790 VSS.n8789 0.214786
R71728 VSS.n8792 VSS.n8791 0.214786
R71729 VSS.n8794 VSS.n8793 0.214786
R71730 VSS.n1430 VSS.n1407 0.214786
R71731 VSS.n8740 VSS.n1395 0.214786
R71732 VSS.n8739 VSS.n8738 0.214786
R71733 VSS.n8737 VSS.n1432 0.214786
R71734 VSS.n8736 VSS.n8735 0.214786
R71735 VSS.n8730 VSS.n8729 0.214786
R71736 VSS.n8728 VSS.n1435 0.214786
R71737 VSS.n8727 VSS.n8726 0.214786
R71738 VSS.n1437 VSS.n1436 0.214786
R71739 VSS.n8722 VSS.n8721 0.214786
R71740 VSS.n8720 VSS.n1439 0.214786
R71741 VSS.n8719 VSS.n8718 0.214786
R71742 VSS.n1441 VSS.n1440 0.214786
R71743 VSS.n8714 VSS.n8713 0.214786
R71744 VSS.n1444 VSS.n1443 0.214786
R71745 VSS.n8693 VSS.n8692 0.214786
R71746 VSS.n1474 VSS.n1464 0.214786
R71747 VSS.n8688 VSS.n8687 0.214786
R71748 VSS.n1477 VSS.n1476 0.214786
R71749 VSS.n8667 VSS.n8666 0.214786
R71750 VSS.n1507 VSS.n1497 0.214786
R71751 VSS.n8662 VSS.n8661 0.214786
R71752 VSS.n8660 VSS.n1509 0.214786
R71753 VSS.n8659 VSS.n8658 0.214786
R71754 VSS.n1511 VSS.n1510 0.214786
R71755 VSS.n8654 VSS.n8653 0.214786
R71756 VSS.n8652 VSS.n1513 0.214786
R71757 VSS.n8651 VSS.n8650 0.214786
R71758 VSS.n1515 VSS.n1514 0.214786
R71759 VSS.n8645 VSS.n8644 0.214786
R71760 VSS.n8643 VSS.n1517 0.214786
R71761 VSS.n8642 VSS.n8641 0.214786
R71762 VSS.n1520 VSS.n1519 0.214786
R71763 VSS.n8637 VSS.n8636 0.214786
R71764 VSS.n8609 VSS.n1522 0.214786
R71765 VSS.n7979 VSS.n1543 0.214786
R71766 VSS.n7981 VSS.n7980 0.214786
R71767 VSS.n7982 VSS.n7975 0.214786
R71768 VSS.n7984 VSS.n7983 0.214786
R71769 VSS.n7985 VSS.n7970 0.214786
R71770 VSS.n7987 VSS.n7986 0.214786
R71771 VSS.n7988 VSS.n7969 0.214786
R71772 VSS.n7990 VSS.n7989 0.214786
R71773 VSS.n7991 VSS.n7964 0.214786
R71774 VSS.n7993 VSS.n7992 0.214786
R71775 VSS.n7994 VSS.n7963 0.214786
R71776 VSS.n7996 VSS.n7995 0.214786
R71777 VSS.n7997 VSS.n2126 0.214786
R71778 VSS.n7999 VSS.n7998 0.214786
R71779 VSS.n2127 VSS.n2092 0.214786
R71780 VSS.n7957 VSS.n7956 0.214786
R71781 VSS.n7955 VSS.n7954 0.214786
R71782 VSS.n7953 VSS.n7952 0.214786
R71783 VSS.n7950 VSS.n7949 0.214786
R71784 VSS.n2132 VSS.n2131 0.214786
R71785 VSS.n2266 VSS.n2222 0.214786
R71786 VSS.n2268 VSS.n2267 0.214786
R71787 VSS.n2223 VSS.n2177 0.214786
R71788 VSS.n2261 VSS.n2260 0.214786
R71789 VSS.n2259 VSS.n2258 0.214786
R71790 VSS.n2257 VSS.n2256 0.214786
R71791 VSS.n2255 VSS.n2225 0.214786
R71792 VSS.n2254 VSS.n2253 0.214786
R71793 VSS.n2228 VSS.n2227 0.214786
R71794 VSS.n2248 VSS.n2247 0.214786
R71795 VSS.n2246 VSS.n2245 0.214786
R71796 VSS.n2244 VSS.n2243 0.214786
R71797 VSS.n2230 VSS.n1727 0.214786
R71798 VSS.n6373 VSS.n6372 0.214786
R71799 VSS.n6386 VSS.n6385 0.214786
R71800 VSS.n3268 VSS.n3247 0.214786
R71801 VSS.n6557 VSS.n6556 0.214786
R71802 VSS.n6555 VSS.n6554 0.214786
R71803 VSS.n6553 VSS.n6552 0.214786
R71804 VSS.n6551 VSS.n3272 0.214786
R71805 VSS.n6550 VSS.n6549 0.214786
R71806 VSS.n6548 VSS.n3273 0.214786
R71807 VSS.n6547 VSS.n6546 0.214786
R71808 VSS.n3291 VSS.n3278 0.214786
R71809 VSS.n3329 VSS.n3316 0.214786
R71810 VSS.n6542 VSS.n6541 0.214786
R71811 VSS.n6540 VSS.n6539 0.214786
R71812 VSS.n6538 VSS.n3334 0.214786
R71813 VSS.n6537 VSS.n6536 0.214786
R71814 VSS.n6535 VSS.n3335 0.214786
R71815 VSS.n6534 VSS.n6533 0.214786
R71816 VSS.n3353 VSS.n3340 0.214786
R71817 VSS.n3391 VSS.n3390 0.214786
R71818 VSS.n6529 VSS.n6528 0.214786
R71819 VSS.n6527 VSS.n6526 0.214786
R71820 VSS.n6525 VSS.n3396 0.214786
R71821 VSS.n6524 VSS.n6523 0.214786
R71822 VSS.n6522 VSS.n3397 0.214786
R71823 VSS.n6521 VSS.n6520 0.214786
R71824 VSS.n6519 VSS.n3402 0.214786
R71825 VSS.n6518 VSS.n6517 0.214786
R71826 VSS.n6516 VSS.n3403 0.214786
R71827 VSS.n6515 VSS.n6514 0.214786
R71828 VSS.n6513 VSS.n3408 0.214786
R71829 VSS.n6512 VSS.n6511 0.214786
R71830 VSS.n6510 VSS.n3409 0.214786
R71831 VSS.n6509 VSS.n6508 0.214786
R71832 VSS.n3427 VSS.n3414 0.214786
R71833 VSS.n3465 VSS.n3464 0.214786
R71834 VSS.n6504 VSS.n6503 0.214786
R71835 VSS.n6502 VSS.n6501 0.214786
R71836 VSS.n6500 VSS.n3470 0.214786
R71837 VSS.n6499 VSS.n6498 0.214786
R71838 VSS.n6497 VSS.n3471 0.214786
R71839 VSS.n6496 VSS.n6495 0.214786
R71840 VSS.n6494 VSS.n3476 0.214786
R71841 VSS.n6493 VSS.n6492 0.214786
R71842 VSS.n6491 VSS.n3477 0.214786
R71843 VSS.n6490 VSS.n6489 0.214786
R71844 VSS.n6488 VSS.n3482 0.214786
R71845 VSS.n6487 VSS.n6486 0.214786
R71846 VSS.n6485 VSS.n3483 0.214786
R71847 VSS.n6484 VSS.n3166 0.214786
R71848 VSS.n6483 VSS.n3179 0.214786
R71849 VSS.n6482 VSS.n6481 0.214786
R71850 VSS.n6479 VSS.n6478 0.214786
R71851 VSS.n6477 VSS.n3136 0.214786
R71852 VSS.n6476 VSS.n3149 0.214786
R71853 VSS.n6475 VSS.n6474 0.214786
R71854 VSS.n6473 VSS.n6472 0.214786
R71855 VSS.n6471 VSS.n3495 0.214786
R71856 VSS.n6470 VSS.n6469 0.214786
R71857 VSS.n6468 VSS.n3496 0.214786
R71858 VSS.n6467 VSS.n6466 0.214786
R71859 VSS.n6465 VSS.n3501 0.214786
R71860 VSS.n6464 VSS.n6463 0.214786
R71861 VSS.n6462 VSS.n3502 0.214786
R71862 VSS.n6461 VSS.n6460 0.214786
R71863 VSS.n6459 VSS.n3507 0.214786
R71864 VSS.n6458 VSS.n6457 0.214786
R71865 VSS.n6456 VSS.n3508 0.214786
R71866 VSS.n6455 VSS.n6454 0.214786
R71867 VSS.n3526 VSS.n3513 0.214786
R71868 VSS.n3564 VSS.n3563 0.214786
R71869 VSS.n6450 VSS.n6449 0.214786
R71870 VSS.n6448 VSS.n6447 0.214786
R71871 VSS.n6446 VSS.n3569 0.214786
R71872 VSS.n6445 VSS.n6444 0.214786
R71873 VSS.n6443 VSS.n3570 0.214786
R71874 VSS.n6442 VSS.n6441 0.214786
R71875 VSS.n6440 VSS.n3575 0.214786
R71876 VSS.n6439 VSS.n6438 0.214786
R71877 VSS.n6437 VSS.n3576 0.214786
R71878 VSS.n6436 VSS.n6435 0.214786
R71879 VSS.n6434 VSS.n3581 0.214786
R71880 VSS.n6433 VSS.n6432 0.214786
R71881 VSS.n6431 VSS.n3582 0.214786
R71882 VSS.n6430 VSS.n6429 0.214786
R71883 VSS.n3599 VSS.n3587 0.214786
R71884 VSS.n3630 VSS.n3623 0.214786
R71885 VSS.n3628 VSS.n3625 0.214786
R71886 VSS.n6413 VSS.n6412 0.214786
R71887 VSS.n6411 VSS.n3627 0.214786
R71888 VSS.n6410 VSS.n6409 0.214786
R71889 VSS.n6408 VSS.n3636 0.214786
R71890 VSS.n6407 VSS.n6406 0.214786
R71891 VSS.n6405 VSS.n6404 0.214786
R71892 VSS.n3642 VSS.n3641 0.214786
R71893 VSS.n6361 VSS.n6341 0.214786
R71894 VSS.n6395 VSS.n6394 0.214786
R71895 VSS.n6393 VSS.n6360 0.214786
R71896 VSS.n6392 VSS.n6391 0.214786
R71897 VSS.n6390 VSS.n6389 0.214786
R71898 VSS.n6388 VSS.n447 0.214786
R71899 VSS.n6387 VSS.n459 0.214786
R71900 VSS.n8566 VSS.n1558 0.208878
R71901 VSS.n1591 VSS.n1558 0.208878
R71902 VSS.n8006 VSS.n1552 0.208878
R71903 VSS.n8830 VSS.n8829 0.208878
R71904 VSS.n8829 VSS.n1355 0.208878
R71905 VSS.n8579 VSS.n1355 0.208878
R71906 VSS.n8005 VSS.n1591 0.208878
R71907 VSS.n8006 VSS.n8005 0.208878
R71908 VSS.n2607 VSS.n2606 0.208878
R71909 VSS.n2606 VSS.n1353 0.208878
R71910 VSS.n8830 VSS.n1353 0.208878
R71911 VSS.n8567 VSS.n8566 0.208878
R71912 VSS.n4674 VSS.n4639 0.188545
R71913 VSS.n9820 VSS.n166 0.188545
R71914 VSS.n8837 VSS.n1352 0.188295
R71915 VSS.n8807 VSS.n8806 0.188295
R71916 VSS.n8549 VSS.n1535 0.188295
R71917 VSS.n8554 VSS.n1595 0.188295
R71918 VSS.n5079 DVSS 0.188139
R71919 VSS.n4973 DVSS 0.188139
R71920 VSS.n5650 DVSS 0.188139
R71921 VSS.n4921 DVSS 0.188139
R71922 VSS.n4113 DVSS 0.188139
R71923 VSS.n5726 DVSS 0.188139
R71924 VSS.n6076 DVSS 0.188139
R71925 VSS.n5957 DVSS 0.188139
R71926 VSS.n6302 DVSS 0.188139
R71927 DVSS VSS.n6317 0.188139
R71928 VSS.n6602 DVSS 0.188139
R71929 DVSS VSS.n6623 0.188139
R71930 VSS.n5888 DVSS 0.188139
R71931 VSS.n6765 DVSS 0.188139
R71932 VSS.n6994 DVSS 0.188139
R71933 DVSS VSS.n7009 0.188139
R71934 VSS.n4671 VSS.n4670 0.177483
R71935 VSS.n163 VSS.n162 0.177483
R71936 VSS.n2789 VSS.n2788 0.169941
R71937 VSS.n7040 VSS.n536 0.169941
R71938 VSS.n7191 VSS.n2496 0.167502
R71939 VSS.n7224 VSS.n2524 0.167502
R71940 VSS.n5251 VSS.n4325 0.156611
R71941 VSS.n276 VSS.n223 0.156611
R71942 VSS.n5262 VSS.n5255 0.156611
R71943 VSS.n5451 VSS.n283 0.156611
R71944 VSS.n4103 VSS.n4102 0.156611
R71945 VSS.n4165 VSS.n4164 0.156611
R71946 VSS.n6069 VSS.n6068 0.156611
R71947 VSS.n5945 VSS.n5944 0.156611
R71948 VSS.n6295 VSS.n6294 0.156611
R71949 VSS.n6326 VSS.n6324 0.156611
R71950 VSS.n6595 VSS.n6594 0.156611
R71951 VSS.n6632 VSS.n6630 0.156611
R71952 VSS.n5793 VSS.n5792 0.156611
R71953 VSS.n6649 VSS.n2970 0.156611
R71954 VSS.n6987 VSS.n6986 0.156611
R71955 VSS.n7018 VSS.n7016 0.156611
R71956 VSS.n2369 VSS.n2366 0.148192
R71957 VSS.n9439 VSS.n9436 0.148192
R71958 VSS.n2275 VSS.n2088 0.148192
R71959 VSS.n8969 VSS.n1094 0.148192
R71960 VSS.n8811 VSS.n8810 0.143739
R71961 VSS.n8541 VSS.n8539 0.143739
R71962 VSS.n7213 VSS.n2536 0.139092
R71963 VSS.n7061 VSS.n2534 0.139092
R71964 VSS.n7182 VSS.n7181 0.139092
R71965 VSS.n7203 VSS.n2518 0.139092
R71966 VSS.n8815 VSS.n1377 0.138035
R71967 VSS.n7113 VSS.n1627 0.138035
R71968 VSS.n2612 VSS.n2566 0.137763
R71969 VSS.n7132 VSS.n7131 0.137763
R71970 VSS.n7151 DVSS 0.136254
R71971 DVSS VSS.n7139 0.136254
R71972 VSS.n2562 VSS.n2546 0.135923
R71973 VSS.n7083 VSS.n7079 0.135923
R71974 VSS.n7265 VSS.n2478 0.135923
R71975 VSS.n7071 VSS.n2513 0.135923
R71976 VSS.n2782 DVSS 0.129215
R71977 DVSS VSS.n7043 0.129215
R71978 VSS.n8860 VSS.n1305 0.120618
R71979 VSS.n8841 VSS.n8840 0.120618
R71980 VSS.n8547 VSS.n1602 0.120618
R71981 VSS.n8558 VSS.n8557 0.120618
R71982 VSS.n7168 VSS.n2528 0.11672
R71983 VSS.n7222 VSS.n2532 0.11672
R71984 VSS.n7257 VSS.n2491 0.11672
R71985 VSS.n7197 VSS.n2511 0.11672
R71986 VSS.n5778 VSS.n2807 0.116189
R71987 VSS.n9584 VSS.n9583 0.116189
R71988 VSS.n7052 VSS.n1296 0.115835
R71989 VSS.n7106 VSS.n1333 0.115835
R71990 VSS.n7121 VSS.n1659 0.115835
R71991 VSS.n7124 VSS.n1580 0.115835
R71992 VSS.n4569 DVSS 0.114389
R71993 DVSS VSS.n4095 0.114389
R71994 DVSS VSS.n6062 0.114389
R71995 DVSS VSS.n6288 0.114389
R71996 VSS.n7166 VSS.n7162 0.114063
R71997 VSS.n7099 VSS.n7096 0.114063
R71998 VSS.n7262 VSS.n7259 0.114063
R71999 VSS.n7243 VSS.n7242 0.114063
R72000 VSS.n3269 VSS.n3234 0.110634
R72001 VSS.n6371 VSS.n6370 0.110634
R72002 VSS.n1829 VSS.n1793 0.110634
R72003 VSS.n9542 VSS.n9541 0.110634
R72004 VSS.n7899 VSS.n1754 0.110634
R72005 VSS.n9470 VSS.n9469 0.110634
R72006 VSS.n2231 VSS.n1715 0.110634
R72007 VSS.n8923 VSS.n8922 0.110634
R72008 VSS.n6643 VSS.n3064 0.11052
R72009 VSS.n5762 VSS.n2838 0.11052
R72010 VSS.n6753 VSS.n6752 0.11052
R72011 VSS.n5744 VSS.n2898 0.11052
R72012 VSS.n5753 VSS.n2864 0.11052
R72013 VSS.n6663 VSS.n6662 0.11052
R72014 VSS.n1591 VSS.n1553 0.110159
R72015 VSS.n8830 VSS.n1354 0.110159
R72016 VSS.n4519 VSS.n4325 0.108278
R72017 VSS.n9691 VSS.n276 0.108278
R72018 VSS.n5255 VSS.n4286 0.108278
R72019 VSS.n9686 VSS.n283 0.108278
R72020 VSS.n4104 VSS.n4103 0.108278
R72021 VSS.n4166 VSS.n4165 0.108278
R72022 VSS.n6071 VSS.n6069 0.108278
R72023 VSS.n5949 VSS.n5945 0.108278
R72024 VSS.n6297 VSS.n6295 0.108278
R72025 VSS.n6324 VSS.n6323 0.108278
R72026 VSS.n6597 VSS.n6595 0.108278
R72027 VSS.n6630 VSS.n6629 0.108278
R72028 VSS.n5795 VSS.n5793 0.108278
R72029 VSS.n6757 VSS.n2970 0.108278
R72030 VSS.n6989 VSS.n6987 0.108278
R72031 VSS.n7016 VSS.n7015 0.108278
R72032 VSS.n7254 VSS.n2492 0.101041
R72033 VSS.n7191 VSS.n2492 0.101041
R72034 VSS.n7249 VSS.n2502 0.101041
R72035 VSS.n7224 VSS.n2522 0.101041
R72036 VSS.n7089 VSS.n2522 0.101041
R72037 VSS.n7089 VSS.n7088 0.101041
R72038 VSS.n7191 VSS.n7190 0.101041
R72039 VSS.n7190 VSS.n2502 0.101041
R72040 VSS.n2553 VSS.n2526 0.101041
R72041 VSS.n7225 VSS.n2526 0.101041
R72042 VSS.n7225 VSS.n7224 0.101041
R72043 VSS.n7254 VSS.n7253 0.101041
R72044 VSS.n4756 VSS.n4755 0.0982778
R72045 VSS.n9773 VSS.n175 0.0982778
R72046 VSS.n5465 VSS.n5464 0.0982778
R72047 VSS.n4159 VSS.n4158 0.0982778
R72048 VSS.n5934 VSS.n428 0.0982778
R72049 VSS.n6338 VSS.n437 0.0982778
R72050 VSS.n6584 VSS.n6582 0.0982778
R72051 VSS.n3667 VSS.n485 0.0982778
R72052 VSS.n5782 VSS.n5780 0.0982778
R72053 VSS.n6661 VSS.n494 0.0982778
R72054 VSS.n6976 VSS.n6974 0.0982778
R72055 VSS.n7030 VSS.n527 0.0982778
R72056 VSS.n6281 VSS.n3246 0.0967008
R72057 VSS.n9597 VSS.n9596 0.0967008
R72058 VSS.n4564 VSS.n3864 0.0941111
R72059 VSS.n4093 VSS.n4092 0.0941111
R72060 VSS.n6059 VSS.n6057 0.0941111
R72061 VSS.n6285 VSS.n6283 0.0941111
R72062 VSS.n3691 VSS.n3624 0.0910315
R72063 VSS.n3700 VSS.n3525 0.0910315
R72064 VSS.n3804 VSS.n3426 0.0910315
R72065 VSS.n3813 VSS.n3352 0.0910315
R72066 VSS.n6340 VSS.n6339 0.0910315
R72067 VSS.n8555 VSS.n1591 0.0873883
R72068 VSS.n8831 VSS.n8830 0.0873883
R72069 VSS.n8074 VSS.n8006 0.0873883
R72070 VSS.n8042 VSS.n1355 0.0873883
R72071 VSS.n8566 VSS.n8565 0.0873883
R72072 VSS.n2606 VSS.n1312 0.0873883
R72073 DVSS VSS.n5078 0.0796667
R72074 DVSS VSS.n271 0.0796667
R72075 DVSS VSS.n5648 0.0796667
R72076 DVSS VSS.n279 0.0796667
R72077 DVSS VSS.n4110 0.0796667
R72078 DVSS VSS.n4168 0.0796667
R72079 DVSS VSS.n6075 0.0796667
R72080 DVSS VSS.n5952 0.0796667
R72081 DVSS VSS.n6301 0.0796667
R72082 VSS.n6319 DVSS 0.0796667
R72083 DVSS VSS.n6601 0.0796667
R72084 VSS.n6625 DVSS 0.0796667
R72085 DVSS VSS.n5799 0.0796667
R72086 DVSS VSS.n6760 0.0796667
R72087 DVSS VSS.n6993 0.0796667
R72088 VSS.n7011 DVSS 0.0796667
R72089 VSS.n7270 VSS.n7269 0.0786237
R72090 VSS.n4753 DVSS 0.0757778
R72091 VSS.n9766 DVSS 0.0757778
R72092 VSS.n5458 DVSS 0.0757778
R72093 DVSS VSS.n4161 0.0757778
R72094 DVSS VSS.n5937 0.0757778
R72095 VSS.n6332 DVSS 0.0757778
R72096 DVSS VSS.n6588 0.0757778
R72097 VSS.n3663 DVSS 0.0757778
R72098 DVSS VSS.n5786 0.0757778
R72099 VSS.n6655 DVSS 0.0757778
R72100 DVSS VSS.n6980 0.0757778
R72101 VSS.n7024 DVSS 0.0757778
R72102 VSS.n994 VSS.n874 0.0740211
R72103 VSS.n973 VSS.n902 0.0740211
R72104 VSS.n2649 VSS.n2468 0.0702987
R72105 VSS.n5893 VSS.n5892 0.0702987
R72106 VSS.n5894 VSS.n3133 0.0702987
R72107 VSS.n5895 VSS.n3711 0.0702987
R72108 VSS.n5899 VSS.n5898 0.0702987
R72109 VSS.n5730 VSS.n5729 0.0702987
R72110 VSS.n4277 VSS.n4073 0.0702987
R72111 VSS.n4510 VSS.n10 0.0702987
R72112 VSS.n9902 VSS.n9901 0.0702987
R72113 VSS.n9015 VSS.n794 0.0621535
R72114 VSS.n9313 VSS.n843 0.0621535
R72115 VSS.n8165 VSS.n8164 0.0621535
R72116 VSS.n8102 VSS.n1909 0.0621535
R72117 VSS.n8276 VSS.n8275 0.0621535
R72118 VSS.n8273 VSS.n8272 0.0621535
R72119 VSS.n9565 VSS.n9564 0.0621535
R72120 VSS.n9562 VSS.n9561 0.0621535
R72121 VSS.n7144 VSS.n2573 0.059675
R72122 VSS.n4974 VSS.n4966 0.0571197
R72123 VSS.n4923 VSS.n4922 0.0571197
R72124 VSS.n5907 VSS.n5905 0.0571197
R72125 VSS.n5959 VSS.n5958 0.0571197
R72126 VSS.n6311 VSS.n6310 0.0571197
R72127 VSS.n3721 VSS.n3709 0.0571197
R72128 VSS.n5827 VSS.n3131 0.0571197
R72129 VSS.n5880 VSS.n5879 0.0571197
R72130 VSS.n6767 VSS.n6766 0.0571197
R72131 VSS.n7003 VSS.n7002 0.0571197
R72132 VSS.n2736 VSS.n2647 0.0571197
R72133 VSS.n5082 VSS.n4507 0.0571197
R72134 VSS.n4925 VSS.n4275 0.0571197
R72135 VSS.n6082 VSS.n6081 0.0571197
R72136 VSS.n6036 VSS.n6035 0.0571197
R72137 VSS.n6308 VSS.n6307 0.0571197
R72138 VSS.n3798 VSS.n3797 0.0571197
R72139 VSS.n5825 VSS.n3195 0.0571197
R72140 VSS.n5885 VSS.n5884 0.0571197
R72141 VSS.n5738 VSS.n2956 0.0571197
R72142 VSS.n7000 VSS.n6999 0.0571197
R72143 VSS.n2739 VSS.n2738 0.0571197
R72144 VSS.n6219 VSS.n3884 0.0569562
R72145 VSS.n3892 VSS.n3883 0.0569562
R72146 VSS.n3891 VSS.n3882 0.0569562
R72147 VSS.n3900 VSS.n3894 0.0569562
R72148 VSS.n3907 VSS.n3899 0.0569562
R72149 VSS.n6060 VSS.n6055 0.0569562
R72150 VSS.n6058 VSS.n6055 0.0569562
R72151 VSS.n6286 VSS.n3819 0.0569562
R72152 VSS.n6284 VSS.n3819 0.0569562
R72153 VSS.n3892 VSS.n3884 0.0569562
R72154 VSS.n3891 VSS.n3883 0.0569562
R72155 VSS.n3907 VSS.n3900 0.0569562
R72156 VSS.n3906 VSS.n3899 0.0569562
R72157 VSS.n6061 VSS.n3905 0.0563
R72158 VSS.n6287 VSS.n3821 0.0563
R72159 VSS.n7145 VSS.n2572 0.0560634
R72160 VSS.n7143 VSS.n2574 0.0560634
R72161 DVSS VSS.n2583 0.0487682
R72162 VSS.n7044 DVSS 0.0487682
R72163 VSS.n5724 VSS.n4029 0.0459225
R72164 VSS.n6124 VSS.n6123 0.0459225
R72165 VSS.n7246 VSS.n2503 0.0450718
R72166 VSS.n7098 VSS.n7056 0.0450718
R72167 VSS.n7097 VSS.n7056 0.0450718
R72168 VSS.n7260 VSS.n2482 0.0450718
R72169 VSS.n7160 VSS.n2555 0.0450718
R72170 VSS.n8084 VSS.n8082 0.0450718
R72171 VSS.n8605 VSS.n1546 0.0450718
R72172 VSS.n1548 VSS.n1546 0.0450718
R72173 VSS.n1548 VSS.n1545 0.0450718
R72174 VSS.n8601 VSS.n8600 0.0450718
R72175 VSS.n8600 VSS.n8599 0.0450718
R72176 VSS.n8595 VSS.n8594 0.0450718
R72177 VSS.n8594 VSS.n8593 0.0450718
R72178 VSS.n8589 VSS.n8574 0.0450718
R72179 VSS.n8589 VSS.n8588 0.0450718
R72180 VSS.n8588 VSS.n8575 0.0450718
R72181 VSS.n8583 VSS.n8576 0.0450718
R72182 VSS.n8583 VSS.n8582 0.0450718
R72183 VSS.n8582 VSS.n8577 0.0450718
R72184 VSS.n7123 VSS.n2588 0.0450718
R72185 VSS.n7120 VSS.n2591 0.0450718
R72186 VSS.n7105 VSS.n2602 0.0450718
R72187 VSS.n7051 VSS.n2604 0.0450718
R72188 VSS.n7245 VSS.n7244 0.0442838
R72189 VSS.n7244 VSS.n2506 0.0442838
R72190 VSS.n7069 VSS.n7066 0.0442838
R72191 VSS.n7072 VSS.n7066 0.0442838
R72192 VSS.n7077 VSS.n7076 0.0442838
R72193 VSS.n7078 VSS.n7077 0.0442838
R72194 VSS.n7058 VSS.n7055 0.0442838
R72195 VSS.n7261 VSS.n2479 0.0442838
R72196 VSS.n7263 VSS.n2479 0.0442838
R72197 VSS.n2477 VSS.n2475 0.0442838
R72198 VSS.n7266 VSS.n2475 0.0442838
R72199 VSS.n2559 VSS.n2556 0.0442838
R72200 VSS.n2563 VSS.n2556 0.0442838
R72201 VSS.n7158 VSS.n7157 0.0442838
R72202 VSS.n7157 VSS.n2554 0.0442838
R72203 VSS.n8085 VSS.n8083 0.0442838
R72204 VSS.n2590 VSS.n2589 0.0442838
R72205 VSS.n7125 VSS.n2590 0.0442838
R72206 VSS.n7119 VSS.n7118 0.0442838
R72207 VSS.n7118 VSS.n7117 0.0442838
R72208 VSS.n2597 VSS.n2596 0.0442838
R72209 VSS.n7114 VSS.n2597 0.0442838
R72210 VSS.n2601 VSS.n2598 0.0442838
R72211 VSS.n7108 VSS.n2601 0.0442838
R72212 VSS.n7104 VSS.n7103 0.0442838
R72213 VSS.n7103 VSS.n7054 0.0442838
R72214 VSS.n7050 VSS.n7049 0.0442838
R72215 VSS.n7049 VSS.n2608 0.0442838
R72216 VSS.n4865 VSS.n4510 0.0437
R72217 VSS.n4924 VSS.n4277 0.0437
R72218 VSS.n5729 VSS.n4075 0.0437
R72219 VSS.n5899 VSS.n4068 0.0437
R72220 VSS.n6309 VSS.n3711 0.0437
R72221 VSS.n6612 VSS.n3133 0.0437
R72222 VSS.n5892 VSS.n5733 0.0437
R72223 VSS.n7001 VSS.n2649 0.0437
R72224 VSS.n7073 VSS.n7072 0.0333378
R72225 VSS.n7074 VSS.n7073 0.0333378
R72226 VSS.n7266 VSS.n2476 0.0333378
R72227 VSS.n2561 VSS.n2476 0.0333378
R72228 VSS.n8598 VSS.n8597 0.0333378
R72229 VSS.n8597 VSS.n8596 0.0333378
R72230 VSS.n7114 VSS.n7112 0.0333378
R72231 VSS.n7112 VSS.n7111 0.0333378
R72232 VSS.n4088 VSS.n3898 0.03245
R72233 VSS.n4094 VSS.n3902 0.03245
R72234 VSS.n4091 VSS.n3897 0.03245
R72235 VSS.n4089 VSS.n3903 0.03245
R72236 VSS.n3904 VSS.n3896 0.03245
R72237 DVSS VSS.n4322 0.0313333
R72238 DVSS VSS.n9765 0.0313333
R72239 DVSS VSS.n4319 0.0313333
R72240 DVSS VSS.n5457 0.0313333
R72241 VSS.n4096 DVSS 0.0313333
R72242 VSS.n4162 DVSS 0.0313333
R72243 VSS.n6064 DVSS 0.0313333
R72244 VSS.n5941 DVSS 0.0313333
R72245 VSS.n6290 DVSS 0.0313333
R72246 DVSS VSS.n6330 0.0313333
R72247 VSS.n6590 DVSS 0.0313333
R72248 VSS.n6638 DVSS 0.0313333
R72249 VSS.n5788 DVSS 0.0313333
R72250 DVSS VSS.n6653 0.0313333
R72251 VSS.n6982 DVSS 0.0313333
R72252 DVSS VSS.n7022 0.0313333
R72253 VSS.n4568 VSS.n3888 0.03065
R72254 VSS.n4567 VSS.n3886 0.03065
R72255 VSS.n4565 VSS.n3889 0.03065
R72256 VSS.n3890 VSS.n3885 0.03065
R72257 VSS.n7073 VSS.n2501 0.0292293
R72258 VSS.n2501 VSS.n2499 0.0292293
R72259 VSS.n2499 VSS.n2494 0.0292293
R72260 VSS.n2494 VSS.n2476 0.0292293
R72261 VSS.n3906 VSS.n3898 0.0287281
R72262 VSS.n6058 VSS.n6056 0.0287281
R72263 VSS.n6284 VSS.n3820 0.0287281
R72264 VSS.n6220 VSS.n6219 0.0287281
R72265 VSS.n6217 VSS.n3882 0.0287281
R72266 VSS.n6216 VSS.n3894 0.0287281
R72267 VSS.n6061 VSS.n6060 0.0287281
R72268 VSS.n6287 VSS.n6286 0.0287281
R72269 VSS.n7889 VSS.n7888 0.0286081
R72270 VSS.n9455 VSS.n9454 0.0286081
R72271 VSS.n5897 VSS.n5731 0.0279406
R72272 VSS.n5897 VSS.n5896 0.0279406
R72273 VSS.n2567 VSS.n2566 0.0276508
R72274 VSS.n7137 VSS.n7134 0.0276508
R72275 VSS.n7137 VSS.n7135 0.0276508
R72276 VSS.n7140 VSS.n2472 0.0276508
R72277 VSS.n2786 VSS.n2781 0.0276508
R72278 VSS.n2786 VSS.n2785 0.0276508
R72279 VSS.n7128 VSS.n2585 0.0276508
R72280 VSS.n7128 VSS.n2586 0.0276508
R72281 VSS.n2613 VSS.n2611 0.0276508
R72282 VSS.n2615 VSS.n2611 0.0276508
R72283 VSS.n7040 VSS.n7036 0.0276508
R72284 VSS.n7195 VSS.n7194 0.0263511
R72285 VSS.n7198 VSS.n7186 0.0263511
R72286 VSS.n7204 VSS.n2537 0.0263511
R72287 VSS.n7220 VSS.n7219 0.0263511
R72288 VSS.n7223 VSS.n2527 0.0263511
R72289 VSS.n7239 VSS.n7238 0.0263511
R72290 VSS.n7241 VSS.n2510 0.0263511
R72291 VSS.n7232 VSS.n2517 0.0263511
R72292 VSS.n7084 VSS.n7060 0.0263511
R72293 VSS.n7093 VSS.n7092 0.0263511
R72294 VSS.n7095 VSS.n7087 0.0263511
R72295 VSS.n2489 VSS.n2485 0.0263511
R72296 VSS.n7258 VSS.n2486 0.0263511
R72297 VSS.n7180 VSS.n2540 0.0263511
R72298 VSS.n7170 VSS.n2545 0.0263511
R72299 VSS.n7165 VSS.n7164 0.0263511
R72300 VSS.n7167 VSS.n2551 0.0263511
R72301 VSS.n8555 VSS.n1592 0.0263511
R72302 VSS.n8548 VSS.n1600 0.0263511
R72303 VSS.n8548 VSS.n1601 0.0263511
R72304 VSS.n1608 VSS.n1607 0.0263511
R72305 VSS.n1610 VSS.n1609 0.0263511
R72306 VSS.n1390 VSS.n1345 0.0263511
R72307 VSS.n1346 VSS.n1345 0.0263511
R72308 VSS.n8836 VSS.n8833 0.0263511
R72309 VSS.n8836 VSS.n8835 0.0263511
R72310 VSS.n8009 VSS.n8004 0.0263511
R72311 VSS.n8068 VSS.n8016 0.0263511
R72312 VSS.n8021 VSS.n8020 0.0263511
R72313 VSS.n8025 VSS.n8024 0.0263511
R72314 VSS.n8049 VSS.n8031 0.0263511
R72315 VSS.n8044 VSS.n8039 0.0263511
R72316 VSS.n8563 VSS.n1566 0.0263511
R72317 VSS.n8390 VSS.n8389 0.0263511
R72318 VSS.n8402 VSS.n8395 0.0263511
R72319 VSS.n8822 VSS.n1364 0.0263511
R72320 VSS.n8845 VSS.n1320 0.0263511
R72321 VSS.n8852 VSS.n1313 0.0263511
R72322 VSS.n4570 VSS.n3888 0.02615
R72323 VSS.n4568 VSS.n3886 0.02615
R72324 VSS.n4567 VSS.n3889 0.02615
R72325 VSS.n4565 VSS.n3885 0.02615
R72326 VSS.n6220 VSS.n3890 0.02615
R72327 VSS.n8573 VSS.n1445 0.0256408
R72328 VSS.n1550 VSS.n1478 0.0256408
R72329 VSS.n2472 VSS.n2469 0.0248855
R72330 VSS.n5124 VSS.n5122 0.0248
R72331 VSS.n5122 VSS.n5120 0.0248
R72332 VSS.n5120 VSS.n5118 0.0248
R72333 VSS.n5118 VSS.n5116 0.0248
R72334 VSS.n5116 VSS.n4461 0.0248
R72335 VSS.n5112 VSS.n4461 0.0248
R72336 VSS.n5112 VSS.n5111 0.0248
R72337 VSS.n5111 VSS.n5110 0.0248
R72338 VSS.n5110 VSS.n4467 0.0248
R72339 VSS.n5106 VSS.n4467 0.0248
R72340 VSS.n5106 VSS.n5105 0.0248
R72341 VSS.n5105 VSS.n5104 0.0248
R72342 VSS.n5104 VSS.n4473 0.0248
R72343 VSS.n5100 VSS.n4473 0.0248
R72344 VSS.n5100 VSS.n5099 0.0248
R72345 VSS.n5098 VSS.n4479 0.0248
R72346 VSS.n5094 VSS.n4479 0.0248
R72347 VSS.n5094 VSS.n5093 0.0248
R72348 VSS.n5093 VSS.n5092 0.0248
R72349 VSS.n5092 VSS.n4485 0.0248
R72350 VSS.n5088 VSS.n4485 0.0248
R72351 VSS.n5088 VSS.n5087 0.0248
R72352 VSS.n5087 VSS.n4490 0.0248
R72353 VSS.n4861 VSS.n4490 0.0248
R72354 VSS.n4863 VSS.n4861 0.0248
R72355 VSS.n4865 VSS.n4863 0.0248
R72356 VSS.n4965 VSS.n4964 0.0248
R72357 VSS.n4964 VSS.n4875 0.0248
R72358 VSS.n4960 VSS.n4875 0.0248
R72359 VSS.n4960 VSS.n4959 0.0248
R72360 VSS.n4959 VSS.n4958 0.0248
R72361 VSS.n4958 VSS.n4881 0.0248
R72362 VSS.n4954 VSS.n4881 0.0248
R72363 VSS.n4954 VSS.n4953 0.0248
R72364 VSS.n4953 VSS.n4952 0.0248
R72365 VSS.n4952 VSS.n4887 0.0248
R72366 VSS.n4948 VSS.n4887 0.0248
R72367 VSS.n4948 VSS.n4947 0.0248
R72368 VSS.n4947 VSS.n4946 0.0248
R72369 VSS.n4946 VSS.n4893 0.0248
R72370 VSS.n4942 VSS.n4893 0.0248
R72371 VSS.n4941 VSS.n4940 0.0248
R72372 VSS.n4940 VSS.n4899 0.0248
R72373 VSS.n4936 VSS.n4899 0.0248
R72374 VSS.n4936 VSS.n4935 0.0248
R72375 VSS.n4935 VSS.n4934 0.0248
R72376 VSS.n4934 VSS.n4905 0.0248
R72377 VSS.n4930 VSS.n4905 0.0248
R72378 VSS.n4930 VSS.n4929 0.0248
R72379 VSS.n4929 VSS.n4928 0.0248
R72380 VSS.n4928 VSS.n4911 0.0248
R72381 VSS.n4924 VSS.n4911 0.0248
R72382 VSS.n5660 VSS.n5658 0.0248
R72383 VSS.n5660 VSS.n4260 0.0248
R72384 VSS.n5666 VSS.n4260 0.0248
R72385 VSS.n5666 VSS.n4243 0.0248
R72386 VSS.n5672 VSS.n4243 0.0248
R72387 VSS.n5672 VSS.n4241 0.0248
R72388 VSS.n5676 VSS.n4241 0.0248
R72389 VSS.n5676 VSS.n4239 0.0248
R72390 VSS.n5680 VSS.n4239 0.0248
R72391 VSS.n5680 VSS.n4237 0.0248
R72392 VSS.n5684 VSS.n4237 0.0248
R72393 VSS.n5684 VSS.n4235 0.0248
R72394 VSS.n5688 VSS.n4235 0.0248
R72395 VSS.n5688 VSS.n4233 0.0248
R72396 VSS.n5692 VSS.n4233 0.0248
R72397 VSS.n5696 VSS.n4231 0.0248
R72398 VSS.n5696 VSS.n4229 0.0248
R72399 VSS.n5700 VSS.n4229 0.0248
R72400 VSS.n5700 VSS.n4227 0.0248
R72401 VSS.n5705 VSS.n4227 0.0248
R72402 VSS.n5705 VSS.n4224 0.0248
R72403 VSS.n5709 VSS.n4224 0.0248
R72404 VSS.n5712 VSS.n5709 0.0248
R72405 VSS.n5714 VSS.n5712 0.0248
R72406 VSS.n5716 VSS.n5714 0.0248
R72407 VSS.n5716 VSS.n4075 0.0248
R72408 VSS.n6122 VSS.n6121 0.0248
R72409 VSS.n6121 VSS.n6120 0.0248
R72410 VSS.n6120 VSS.n4032 0.0248
R72411 VSS.n6116 VSS.n4032 0.0248
R72412 VSS.n6116 VSS.n6115 0.0248
R72413 VSS.n6115 VSS.n6114 0.0248
R72414 VSS.n6114 VSS.n4038 0.0248
R72415 VSS.n6110 VSS.n4038 0.0248
R72416 VSS.n6110 VSS.n6109 0.0248
R72417 VSS.n6109 VSS.n6108 0.0248
R72418 VSS.n6108 VSS.n4044 0.0248
R72419 VSS.n6104 VSS.n4044 0.0248
R72420 VSS.n6104 VSS.n6103 0.0248
R72421 VSS.n6103 VSS.n6102 0.0248
R72422 VSS.n6102 VSS.n4050 0.0248
R72423 VSS.n6098 VSS.n6097 0.0248
R72424 VSS.n6097 VSS.n6096 0.0248
R72425 VSS.n6096 VSS.n4056 0.0248
R72426 VSS.n6092 VSS.n4056 0.0248
R72427 VSS.n6092 VSS.n6091 0.0248
R72428 VSS.n6091 VSS.n6090 0.0248
R72429 VSS.n6090 VSS.n4062 0.0248
R72430 VSS.n6086 VSS.n4062 0.0248
R72431 VSS.n6086 VSS.n6085 0.0248
R72432 VSS.n6085 VSS.n6084 0.0248
R72433 VSS.n6084 VSS.n4068 0.0248
R72434 VSS.n6034 VSS.n6033 0.0248
R72435 VSS.n6033 VSS.n6032 0.0248
R72436 VSS.n6032 VSS.n5962 0.0248
R72437 VSS.n6028 VSS.n5962 0.0248
R72438 VSS.n6028 VSS.n6027 0.0248
R72439 VSS.n6027 VSS.n6026 0.0248
R72440 VSS.n6026 VSS.n5968 0.0248
R72441 VSS.n6022 VSS.n5968 0.0248
R72442 VSS.n6022 VSS.n6021 0.0248
R72443 VSS.n6021 VSS.n6020 0.0248
R72444 VSS.n6020 VSS.n5974 0.0248
R72445 VSS.n6016 VSS.n5974 0.0248
R72446 VSS.n6016 VSS.n6015 0.0248
R72447 VSS.n6015 VSS.n6014 0.0248
R72448 VSS.n6014 VSS.n5980 0.0248
R72449 VSS.n6010 VSS.n6009 0.0248
R72450 VSS.n6009 VSS.n6008 0.0248
R72451 VSS.n6008 VSS.n5986 0.0248
R72452 VSS.n6004 VSS.n5986 0.0248
R72453 VSS.n6004 VSS.n6003 0.0248
R72454 VSS.n6003 VSS.n6002 0.0248
R72455 VSS.n6002 VSS.n5992 0.0248
R72456 VSS.n5998 VSS.n5992 0.0248
R72457 VSS.n5998 VSS.n5997 0.0248
R72458 VSS.n5997 VSS.n3713 0.0248
R72459 VSS.n6309 VSS.n3713 0.0248
R72460 VSS.n3796 VSS.n3795 0.0248
R72461 VSS.n3795 VSS.n3794 0.0248
R72462 VSS.n3794 VSS.n3792 0.0248
R72463 VSS.n3792 VSS.n3790 0.0248
R72464 VSS.n3790 VSS.n3788 0.0248
R72465 VSS.n3788 VSS.n3786 0.0248
R72466 VSS.n3786 VSS.n3784 0.0248
R72467 VSS.n3784 VSS.n3782 0.0248
R72468 VSS.n3782 VSS.n3779 0.0248
R72469 VSS.n3779 VSS.n3778 0.0248
R72470 VSS.n3778 VSS.n3776 0.0248
R72471 VSS.n3776 VSS.n3774 0.0248
R72472 VSS.n3774 VSS.n3772 0.0248
R72473 VSS.n3772 VSS.n3770 0.0248
R72474 VSS.n3770 VSS.n3768 0.0248
R72475 VSS.n3765 VSS.n3764 0.0248
R72476 VSS.n3764 VSS.n3762 0.0248
R72477 VSS.n3762 VSS.n3760 0.0248
R72478 VSS.n3760 VSS.n3758 0.0248
R72479 VSS.n3758 VSS.n3756 0.0248
R72480 VSS.n3756 VSS.n3754 0.0248
R72481 VSS.n3754 VSS.n3752 0.0248
R72482 VSS.n3752 VSS.n3749 0.0248
R72483 VSS.n3749 VSS.n3748 0.0248
R72484 VSS.n3748 VSS.n3162 0.0248
R72485 VSS.n6612 VSS.n3162 0.0248
R72486 VSS.n5826 VSS.n5824 0.0248
R72487 VSS.n5830 VSS.n5824 0.0248
R72488 VSS.n5830 VSS.n5822 0.0248
R72489 VSS.n5834 VSS.n5822 0.0248
R72490 VSS.n5834 VSS.n5820 0.0248
R72491 VSS.n5838 VSS.n5820 0.0248
R72492 VSS.n5838 VSS.n5818 0.0248
R72493 VSS.n5842 VSS.n5818 0.0248
R72494 VSS.n5842 VSS.n5816 0.0248
R72495 VSS.n5846 VSS.n5816 0.0248
R72496 VSS.n5846 VSS.n5814 0.0248
R72497 VSS.n5851 VSS.n5814 0.0248
R72498 VSS.n5851 VSS.n5812 0.0248
R72499 VSS.n5855 VSS.n5812 0.0248
R72500 VSS.n5856 VSS.n5855 0.0248
R72501 VSS.n5859 VSS.n5809 0.0248
R72502 VSS.n5863 VSS.n5809 0.0248
R72503 VSS.n5863 VSS.n5807 0.0248
R72504 VSS.n5867 VSS.n5807 0.0248
R72505 VSS.n5867 VSS.n5805 0.0248
R72506 VSS.n5871 VSS.n5805 0.0248
R72507 VSS.n5871 VSS.n5803 0.0248
R72508 VSS.n5875 VSS.n5803 0.0248
R72509 VSS.n5875 VSS.n5801 0.0248
R72510 VSS.n5882 VSS.n5801 0.0248
R72511 VSS.n5882 VSS.n5733 0.0248
R72512 VSS.n6770 VSS.n2957 0.0248
R72513 VSS.n6770 VSS.n2954 0.0248
R72514 VSS.n6774 VSS.n2954 0.0248
R72515 VSS.n6777 VSS.n6774 0.0248
R72516 VSS.n6780 VSS.n6777 0.0248
R72517 VSS.n6783 VSS.n6780 0.0248
R72518 VSS.n6786 VSS.n6783 0.0248
R72519 VSS.n6787 VSS.n6786 0.0248
R72520 VSS.n6792 VSS.n6787 0.0248
R72521 VSS.n6795 VSS.n6792 0.0248
R72522 VSS.n6798 VSS.n6795 0.0248
R72523 VSS.n6800 VSS.n6798 0.0248
R72524 VSS.n6802 VSS.n6800 0.0248
R72525 VSS.n6802 VSS.n2938 0.0248
R72526 VSS.n6837 VSS.n2938 0.0248
R72527 VSS.n6836 VSS.n6835 0.0248
R72528 VSS.n6835 VSS.n6810 0.0248
R72529 VSS.n6831 VSS.n6810 0.0248
R72530 VSS.n6831 VSS.n6830 0.0248
R72531 VSS.n6830 VSS.n6829 0.0248
R72532 VSS.n6829 VSS.n6816 0.0248
R72533 VSS.n6825 VSS.n6816 0.0248
R72534 VSS.n6825 VSS.n6824 0.0248
R72535 VSS.n6824 VSS.n6823 0.0248
R72536 VSS.n6823 VSS.n2651 0.0248
R72537 VSS.n7001 VSS.n2651 0.0248
R72538 VSS.n2737 VSS.n2659 0.0248
R72539 VSS.n2733 VSS.n2659 0.0248
R72540 VSS.n2733 VSS.n2661 0.0248
R72541 VSS.n2729 VSS.n2661 0.0248
R72542 VSS.n2729 VSS.n2728 0.0248
R72543 VSS.n2728 VSS.n2727 0.0248
R72544 VSS.n2727 VSS.n2666 0.0248
R72545 VSS.n2723 VSS.n2666 0.0248
R72546 VSS.n2723 VSS.n2722 0.0248
R72547 VSS.n2722 VSS.n2721 0.0248
R72548 VSS.n2721 VSS.n2672 0.0248
R72549 VSS.n2717 VSS.n2672 0.0248
R72550 VSS.n2717 VSS.n2716 0.0248
R72551 VSS.n2716 VSS.n2715 0.0248
R72552 VSS.n2715 VSS.n2678 0.0248
R72553 VSS.n2711 VSS.n2710 0.0248
R72554 VSS.n2710 VSS.n2709 0.0248
R72555 VSS.n2709 VSS.n2684 0.0248
R72556 VSS.n2705 VSS.n2684 0.0248
R72557 VSS.n2705 VSS.n2704 0.0248
R72558 VSS.n2704 VSS.n2703 0.0248
R72559 VSS.n2703 VSS.n2690 0.0248
R72560 VSS.n2699 VSS.n2690 0.0248
R72561 VSS.n2699 VSS.n2698 0.0248
R72562 VSS.n2698 VSS.n2697 0.0248
R72563 VSS.n2697 VSS.n2573 0.0248
R72564 VSS.n7144 VSS.n2469 0.0248
R72565 VSS.n7269 VSS.n2469 0.0248
R72566 VSS.n4088 VSS.n3902 0.02435
R72567 VSS.n4094 VSS.n3897 0.02435
R72568 VSS.n4091 VSS.n3903 0.02435
R72569 VSS.n4089 VSS.n3896 0.02435
R72570 VSS.n6214 VSS.n3904 0.02435
R72571 VSS.n2339 VSS.n2338 0.0243462
R72572 VSS.n2364 VSS.n2339 0.0243462
R72573 VSS.n2346 VSS.n2345 0.0243462
R72574 VSS.n2359 VSS.n2346 0.0243462
R72575 VSS.n2356 VSS.n2350 0.0243462
R72576 VSS.n2350 VSS.n762 0.0243462
R72577 VSS.n9451 VSS.n764 0.0243462
R72578 VSS.n9449 VSS.n764 0.0243462
R72579 VSS.n774 VSS.n773 0.0243462
R72580 VSS.n9444 VSS.n774 0.0243462
R72581 VSS.n9371 VSS.n9370 0.0243462
R72582 VSS.n9439 VSS.n9371 0.0243462
R72583 VSS.n8597 VSS.n8571 0.0237143
R72584 VSS.n8571 VSS.n1358 0.0237143
R72585 VSS.n1556 VSS.n1358 0.0237143
R72586 VSS.n7112 VSS.n1556 0.0237143
R72587 VSS.n9452 VSS.n762 0.0233846
R72588 VSS.n9452 VSS.n9451 0.0233846
R72589 VSS.n2466 VSS.n2445 0.0233846
R72590 VSS.n2466 VSS.n2465 0.0233846
R72591 VSS.n4463 VSS.n4460 0.0233169
R72592 VSS.n4464 VSS.n4463 0.0233169
R72593 VSS.n4465 VSS.n4464 0.0233169
R72594 VSS.n4466 VSS.n4465 0.0233169
R72595 VSS.n4469 VSS.n4466 0.0233169
R72596 VSS.n4470 VSS.n4469 0.0233169
R72597 VSS.n4471 VSS.n4470 0.0233169
R72598 VSS.n4472 VSS.n4471 0.0233169
R72599 VSS.n4475 VSS.n4472 0.0233169
R72600 VSS.n4476 VSS.n4475 0.0233169
R72601 VSS.n4477 VSS.n4476 0.0233169
R72602 VSS.n4478 VSS.n4477 0.0233169
R72603 VSS.n4481 VSS.n4478 0.0233169
R72604 VSS.n4482 VSS.n4481 0.0233169
R72605 VSS.n4483 VSS.n4482 0.0233169
R72606 VSS.n4484 VSS.n4483 0.0233169
R72607 VSS.n4487 VSS.n4484 0.0233169
R72608 VSS.n4488 VSS.n4487 0.0233169
R72609 VSS.n4966 VSS.n4874 0.0233169
R72610 VSS.n4877 VSS.n4874 0.0233169
R72611 VSS.n4878 VSS.n4877 0.0233169
R72612 VSS.n4879 VSS.n4878 0.0233169
R72613 VSS.n4880 VSS.n4879 0.0233169
R72614 VSS.n4883 VSS.n4880 0.0233169
R72615 VSS.n4884 VSS.n4883 0.0233169
R72616 VSS.n4885 VSS.n4884 0.0233169
R72617 VSS.n4886 VSS.n4885 0.0233169
R72618 VSS.n4889 VSS.n4886 0.0233169
R72619 VSS.n4890 VSS.n4889 0.0233169
R72620 VSS.n4891 VSS.n4890 0.0233169
R72621 VSS.n4892 VSS.n4891 0.0233169
R72622 VSS.n4895 VSS.n4892 0.0233169
R72623 VSS.n4896 VSS.n4895 0.0233169
R72624 VSS.n4897 VSS.n4896 0.0233169
R72625 VSS.n4898 VSS.n4897 0.0233169
R72626 VSS.n4901 VSS.n4898 0.0233169
R72627 VSS.n4902 VSS.n4901 0.0233169
R72628 VSS.n4903 VSS.n4902 0.0233169
R72629 VSS.n4904 VSS.n4903 0.0233169
R72630 VSS.n4907 VSS.n4904 0.0233169
R72631 VSS.n4908 VSS.n4907 0.0233169
R72632 VSS.n4909 VSS.n4908 0.0233169
R72633 VSS.n4910 VSS.n4909 0.0233169
R72634 VSS.n4912 VSS.n4910 0.0233169
R72635 VSS.n4923 VSS.n4912 0.0233169
R72636 VSS.n5671 VSS.n4240 0.0233169
R72637 VSS.n5677 VSS.n4240 0.0233169
R72638 VSS.n5678 VSS.n5677 0.0233169
R72639 VSS.n5679 VSS.n5678 0.0233169
R72640 VSS.n5679 VSS.n4236 0.0233169
R72641 VSS.n5685 VSS.n4236 0.0233169
R72642 VSS.n5686 VSS.n5685 0.0233169
R72643 VSS.n5687 VSS.n5686 0.0233169
R72644 VSS.n5687 VSS.n4232 0.0233169
R72645 VSS.n5693 VSS.n4232 0.0233169
R72646 VSS.n5694 VSS.n5693 0.0233169
R72647 VSS.n5695 VSS.n5694 0.0233169
R72648 VSS.n5695 VSS.n4228 0.0233169
R72649 VSS.n5701 VSS.n4228 0.0233169
R72650 VSS.n5702 VSS.n5701 0.0233169
R72651 VSS.n5704 VSS.n5702 0.0233169
R72652 VSS.n5704 VSS.n5703 0.0233169
R72653 VSS.n5703 VSS.n4225 0.0233169
R72654 VSS.n4030 VSS.n4029 0.0233169
R72655 VSS.n4031 VSS.n4030 0.0233169
R72656 VSS.n4034 VSS.n4031 0.0233169
R72657 VSS.n4035 VSS.n4034 0.0233169
R72658 VSS.n4036 VSS.n4035 0.0233169
R72659 VSS.n4037 VSS.n4036 0.0233169
R72660 VSS.n4040 VSS.n4037 0.0233169
R72661 VSS.n4041 VSS.n4040 0.0233169
R72662 VSS.n4042 VSS.n4041 0.0233169
R72663 VSS.n4043 VSS.n4042 0.0233169
R72664 VSS.n4046 VSS.n4043 0.0233169
R72665 VSS.n4047 VSS.n4046 0.0233169
R72666 VSS.n4048 VSS.n4047 0.0233169
R72667 VSS.n4049 VSS.n4048 0.0233169
R72668 VSS.n4052 VSS.n4049 0.0233169
R72669 VSS.n4053 VSS.n4052 0.0233169
R72670 VSS.n4054 VSS.n4053 0.0233169
R72671 VSS.n4055 VSS.n4054 0.0233169
R72672 VSS.n4058 VSS.n4055 0.0233169
R72673 VSS.n4059 VSS.n4058 0.0233169
R72674 VSS.n4060 VSS.n4059 0.0233169
R72675 VSS.n4061 VSS.n4060 0.0233169
R72676 VSS.n4064 VSS.n4061 0.0233169
R72677 VSS.n4065 VSS.n4064 0.0233169
R72678 VSS.n4066 VSS.n4065 0.0233169
R72679 VSS.n4067 VSS.n4066 0.0233169
R72680 VSS.n5905 VSS.n4067 0.0233169
R72681 VSS.n5960 VSS.n5959 0.0233169
R72682 VSS.n5961 VSS.n5960 0.0233169
R72683 VSS.n5964 VSS.n5961 0.0233169
R72684 VSS.n5965 VSS.n5964 0.0233169
R72685 VSS.n5966 VSS.n5965 0.0233169
R72686 VSS.n5967 VSS.n5966 0.0233169
R72687 VSS.n5970 VSS.n5967 0.0233169
R72688 VSS.n5971 VSS.n5970 0.0233169
R72689 VSS.n5972 VSS.n5971 0.0233169
R72690 VSS.n5973 VSS.n5972 0.0233169
R72691 VSS.n5976 VSS.n5973 0.0233169
R72692 VSS.n5977 VSS.n5976 0.0233169
R72693 VSS.n5978 VSS.n5977 0.0233169
R72694 VSS.n5979 VSS.n5978 0.0233169
R72695 VSS.n5982 VSS.n5979 0.0233169
R72696 VSS.n5983 VSS.n5982 0.0233169
R72697 VSS.n5984 VSS.n5983 0.0233169
R72698 VSS.n5985 VSS.n5984 0.0233169
R72699 VSS.n5988 VSS.n5985 0.0233169
R72700 VSS.n5989 VSS.n5988 0.0233169
R72701 VSS.n5990 VSS.n5989 0.0233169
R72702 VSS.n5991 VSS.n5990 0.0233169
R72703 VSS.n5994 VSS.n5991 0.0233169
R72704 VSS.n5995 VSS.n5994 0.0233169
R72705 VSS.n5996 VSS.n5995 0.0233169
R72706 VSS.n5996 VSS.n3712 0.0233169
R72707 VSS.n6310 VSS.n3712 0.0233169
R72708 VSS.n3722 VSS.n3721 0.0233169
R72709 VSS.n3723 VSS.n3722 0.0233169
R72710 VSS.n3730 VSS.n3729 0.0233169
R72711 VSS.n3737 VSS.n3736 0.0233169
R72712 VSS.n3745 VSS.n3744 0.0233169
R72713 VSS.n5828 VSS.n5827 0.0233169
R72714 VSS.n5829 VSS.n5828 0.0233169
R72715 VSS.n5829 VSS.n5821 0.0233169
R72716 VSS.n5835 VSS.n5821 0.0233169
R72717 VSS.n5836 VSS.n5835 0.0233169
R72718 VSS.n5837 VSS.n5836 0.0233169
R72719 VSS.n5837 VSS.n5817 0.0233169
R72720 VSS.n5843 VSS.n5817 0.0233169
R72721 VSS.n5844 VSS.n5843 0.0233169
R72722 VSS.n5845 VSS.n5844 0.0233169
R72723 VSS.n5845 VSS.n5813 0.0233169
R72724 VSS.n5852 VSS.n5813 0.0233169
R72725 VSS.n5853 VSS.n5852 0.0233169
R72726 VSS.n5854 VSS.n5853 0.0233169
R72727 VSS.n5854 VSS.n5810 0.0233169
R72728 VSS.n5860 VSS.n5810 0.0233169
R72729 VSS.n5861 VSS.n5860 0.0233169
R72730 VSS.n5862 VSS.n5861 0.0233169
R72731 VSS.n5862 VSS.n5806 0.0233169
R72732 VSS.n5868 VSS.n5806 0.0233169
R72733 VSS.n5869 VSS.n5868 0.0233169
R72734 VSS.n5870 VSS.n5869 0.0233169
R72735 VSS.n5870 VSS.n5802 0.0233169
R72736 VSS.n5876 VSS.n5802 0.0233169
R72737 VSS.n5877 VSS.n5876 0.0233169
R72738 VSS.n5881 VSS.n5877 0.0233169
R72739 VSS.n5881 VSS.n5880 0.0233169
R72740 VSS.n6769 VSS.n6767 0.0233169
R72741 VSS.n6769 VSS.n6768 0.0233169
R72742 VSS.n6768 VSS.n2955 0.0233169
R72743 VSS.n6789 VSS.n6788 0.0233169
R72744 VSS.n6808 VSS.n6807 0.0233169
R72745 VSS.n6809 VSS.n6808 0.0233169
R72746 VSS.n6812 VSS.n6809 0.0233169
R72747 VSS.n6813 VSS.n6812 0.0233169
R72748 VSS.n6814 VSS.n6813 0.0233169
R72749 VSS.n6815 VSS.n6814 0.0233169
R72750 VSS.n6818 VSS.n6815 0.0233169
R72751 VSS.n6819 VSS.n6818 0.0233169
R72752 VSS.n6820 VSS.n6819 0.0233169
R72753 VSS.n6821 VSS.n6820 0.0233169
R72754 VSS.n6821 VSS.n2650 0.0233169
R72755 VSS.n7002 VSS.n2650 0.0233169
R72756 VSS.n2736 VSS.n2735 0.0233169
R72757 VSS.n2735 VSS.n2734 0.0233169
R72758 VSS.n2734 VSS.n2660 0.0233169
R72759 VSS.n2663 VSS.n2660 0.0233169
R72760 VSS.n2664 VSS.n2663 0.0233169
R72761 VSS.n2665 VSS.n2664 0.0233169
R72762 VSS.n2668 VSS.n2665 0.0233169
R72763 VSS.n2669 VSS.n2668 0.0233169
R72764 VSS.n2670 VSS.n2669 0.0233169
R72765 VSS.n2671 VSS.n2670 0.0233169
R72766 VSS.n2674 VSS.n2671 0.0233169
R72767 VSS.n2675 VSS.n2674 0.0233169
R72768 VSS.n2676 VSS.n2675 0.0233169
R72769 VSS.n2677 VSS.n2676 0.0233169
R72770 VSS.n2680 VSS.n2677 0.0233169
R72771 VSS.n2681 VSS.n2680 0.0233169
R72772 VSS.n2682 VSS.n2681 0.0233169
R72773 VSS.n2683 VSS.n2682 0.0233169
R72774 VSS.n2686 VSS.n2683 0.0233169
R72775 VSS.n2687 VSS.n2686 0.0233169
R72776 VSS.n2688 VSS.n2687 0.0233169
R72777 VSS.n2689 VSS.n2688 0.0233169
R72778 VSS.n2692 VSS.n2689 0.0233169
R72779 VSS.n2693 VSS.n2692 0.0233169
R72780 VSS.n2694 VSS.n2693 0.0233169
R72781 VSS.n2695 VSS.n2694 0.0233169
R72782 VSS.n2695 VSS.n2572 0.0233169
R72783 VSS.n7148 VSS.n7145 0.0233169
R72784 VSS.n5115 VSS.n5114 0.0233169
R72785 VSS.n5114 VSS.n5113 0.0233169
R72786 VSS.n5113 VSS.n4462 0.0233169
R72787 VSS.n5109 VSS.n4462 0.0233169
R72788 VSS.n5109 VSS.n5108 0.0233169
R72789 VSS.n5108 VSS.n5107 0.0233169
R72790 VSS.n5107 VSS.n4468 0.0233169
R72791 VSS.n5103 VSS.n4468 0.0233169
R72792 VSS.n5103 VSS.n5102 0.0233169
R72793 VSS.n5102 VSS.n5101 0.0233169
R72794 VSS.n5101 VSS.n4474 0.0233169
R72795 VSS.n5097 VSS.n4474 0.0233169
R72796 VSS.n5097 VSS.n5096 0.0233169
R72797 VSS.n5096 VSS.n5095 0.0233169
R72798 VSS.n5095 VSS.n4480 0.0233169
R72799 VSS.n5091 VSS.n4480 0.0233169
R72800 VSS.n5091 VSS.n5090 0.0233169
R72801 VSS.n5090 VSS.n5089 0.0233169
R72802 VSS.n4963 VSS.n4507 0.0233169
R72803 VSS.n4963 VSS.n4962 0.0233169
R72804 VSS.n4962 VSS.n4961 0.0233169
R72805 VSS.n4961 VSS.n4876 0.0233169
R72806 VSS.n4957 VSS.n4876 0.0233169
R72807 VSS.n4957 VSS.n4956 0.0233169
R72808 VSS.n4956 VSS.n4955 0.0233169
R72809 VSS.n4955 VSS.n4882 0.0233169
R72810 VSS.n4951 VSS.n4882 0.0233169
R72811 VSS.n4951 VSS.n4950 0.0233169
R72812 VSS.n4950 VSS.n4949 0.0233169
R72813 VSS.n4949 VSS.n4888 0.0233169
R72814 VSS.n4945 VSS.n4888 0.0233169
R72815 VSS.n4945 VSS.n4944 0.0233169
R72816 VSS.n4944 VSS.n4943 0.0233169
R72817 VSS.n4943 VSS.n4894 0.0233169
R72818 VSS.n4939 VSS.n4894 0.0233169
R72819 VSS.n4939 VSS.n4938 0.0233169
R72820 VSS.n4938 VSS.n4937 0.0233169
R72821 VSS.n4937 VSS.n4900 0.0233169
R72822 VSS.n4933 VSS.n4900 0.0233169
R72823 VSS.n4933 VSS.n4932 0.0233169
R72824 VSS.n4932 VSS.n4931 0.0233169
R72825 VSS.n4931 VSS.n4906 0.0233169
R72826 VSS.n4927 VSS.n4906 0.0233169
R72827 VSS.n4927 VSS.n4926 0.0233169
R72828 VSS.n4926 VSS.n4925 0.0233169
R72829 VSS.n5674 VSS.n5673 0.0233169
R72830 VSS.n5675 VSS.n5674 0.0233169
R72831 VSS.n5675 VSS.n4238 0.0233169
R72832 VSS.n5681 VSS.n4238 0.0233169
R72833 VSS.n5682 VSS.n5681 0.0233169
R72834 VSS.n5683 VSS.n5682 0.0233169
R72835 VSS.n5683 VSS.n4234 0.0233169
R72836 VSS.n5689 VSS.n4234 0.0233169
R72837 VSS.n5690 VSS.n5689 0.0233169
R72838 VSS.n5691 VSS.n5690 0.0233169
R72839 VSS.n5691 VSS.n4230 0.0233169
R72840 VSS.n5697 VSS.n4230 0.0233169
R72841 VSS.n5698 VSS.n5697 0.0233169
R72842 VSS.n5699 VSS.n5698 0.0233169
R72843 VSS.n5699 VSS.n4226 0.0233169
R72844 VSS.n5706 VSS.n4226 0.0233169
R72845 VSS.n5707 VSS.n5706 0.0233169
R72846 VSS.n5708 VSS.n5707 0.0233169
R72847 VSS.n6123 VSS.n4028 0.0233169
R72848 VSS.n6119 VSS.n4028 0.0233169
R72849 VSS.n6119 VSS.n6118 0.0233169
R72850 VSS.n6118 VSS.n6117 0.0233169
R72851 VSS.n6117 VSS.n4033 0.0233169
R72852 VSS.n6113 VSS.n4033 0.0233169
R72853 VSS.n6113 VSS.n6112 0.0233169
R72854 VSS.n6112 VSS.n6111 0.0233169
R72855 VSS.n6111 VSS.n4039 0.0233169
R72856 VSS.n6107 VSS.n4039 0.0233169
R72857 VSS.n6107 VSS.n6106 0.0233169
R72858 VSS.n6106 VSS.n6105 0.0233169
R72859 VSS.n6105 VSS.n4045 0.0233169
R72860 VSS.n6101 VSS.n4045 0.0233169
R72861 VSS.n6101 VSS.n6100 0.0233169
R72862 VSS.n6100 VSS.n6099 0.0233169
R72863 VSS.n6099 VSS.n4051 0.0233169
R72864 VSS.n6095 VSS.n4051 0.0233169
R72865 VSS.n6095 VSS.n6094 0.0233169
R72866 VSS.n6094 VSS.n6093 0.0233169
R72867 VSS.n6093 VSS.n4057 0.0233169
R72868 VSS.n6089 VSS.n4057 0.0233169
R72869 VSS.n6089 VSS.n6088 0.0233169
R72870 VSS.n6088 VSS.n6087 0.0233169
R72871 VSS.n6087 VSS.n4063 0.0233169
R72872 VSS.n6083 VSS.n4063 0.0233169
R72873 VSS.n6083 VSS.n6082 0.0233169
R72874 VSS.n6035 VSS.n5901 0.0233169
R72875 VSS.n6031 VSS.n5901 0.0233169
R72876 VSS.n6031 VSS.n6030 0.0233169
R72877 VSS.n6030 VSS.n6029 0.0233169
R72878 VSS.n6029 VSS.n5963 0.0233169
R72879 VSS.n6025 VSS.n5963 0.0233169
R72880 VSS.n6025 VSS.n6024 0.0233169
R72881 VSS.n6024 VSS.n6023 0.0233169
R72882 VSS.n6023 VSS.n5969 0.0233169
R72883 VSS.n6019 VSS.n5969 0.0233169
R72884 VSS.n6019 VSS.n6018 0.0233169
R72885 VSS.n6018 VSS.n6017 0.0233169
R72886 VSS.n6017 VSS.n5975 0.0233169
R72887 VSS.n6013 VSS.n5975 0.0233169
R72888 VSS.n6013 VSS.n6012 0.0233169
R72889 VSS.n6012 VSS.n6011 0.0233169
R72890 VSS.n6011 VSS.n5981 0.0233169
R72891 VSS.n6007 VSS.n5981 0.0233169
R72892 VSS.n6007 VSS.n6006 0.0233169
R72893 VSS.n6006 VSS.n6005 0.0233169
R72894 VSS.n6005 VSS.n5987 0.0233169
R72895 VSS.n6001 VSS.n5987 0.0233169
R72896 VSS.n6001 VSS.n6000 0.0233169
R72897 VSS.n6000 VSS.n5999 0.0233169
R72898 VSS.n5999 VSS.n5993 0.0233169
R72899 VSS.n5993 VSS.n3714 0.0233169
R72900 VSS.n6308 VSS.n3714 0.0233169
R72901 VSS.n3797 VSS.n3720 0.0233169
R72902 VSS.n3793 VSS.n3720 0.0233169
R72903 VSS.n3781 VSS.n3780 0.0233169
R72904 VSS.n3767 VSS.n3766 0.0233169
R72905 VSS.n3751 VSS.n3750 0.0233169
R72906 VSS.n5825 VSS.n5823 0.0233169
R72907 VSS.n5831 VSS.n5823 0.0233169
R72908 VSS.n5832 VSS.n5831 0.0233169
R72909 VSS.n5833 VSS.n5832 0.0233169
R72910 VSS.n5833 VSS.n5819 0.0233169
R72911 VSS.n5839 VSS.n5819 0.0233169
R72912 VSS.n5840 VSS.n5839 0.0233169
R72913 VSS.n5841 VSS.n5840 0.0233169
R72914 VSS.n5841 VSS.n5815 0.0233169
R72915 VSS.n5847 VSS.n5815 0.0233169
R72916 VSS.n5848 VSS.n5847 0.0233169
R72917 VSS.n5850 VSS.n5848 0.0233169
R72918 VSS.n5850 VSS.n5849 0.0233169
R72919 VSS.n5849 VSS.n5811 0.0233169
R72920 VSS.n5857 VSS.n5811 0.0233169
R72921 VSS.n5858 VSS.n5857 0.0233169
R72922 VSS.n5858 VSS.n5808 0.0233169
R72923 VSS.n5864 VSS.n5808 0.0233169
R72924 VSS.n5865 VSS.n5864 0.0233169
R72925 VSS.n5866 VSS.n5865 0.0233169
R72926 VSS.n5866 VSS.n5804 0.0233169
R72927 VSS.n5872 VSS.n5804 0.0233169
R72928 VSS.n5873 VSS.n5872 0.0233169
R72929 VSS.n5874 VSS.n5873 0.0233169
R72930 VSS.n5874 VSS.n5800 0.0233169
R72931 VSS.n5883 VSS.n5800 0.0233169
R72932 VSS.n5884 VSS.n5883 0.0233169
R72933 VSS.n6771 VSS.n2956 0.0233169
R72934 VSS.n6772 VSS.n6771 0.0233169
R72935 VSS.n6773 VSS.n6772 0.0233169
R72936 VSS.n6791 VSS.n6790 0.0233169
R72937 VSS.n6838 VSS.n2937 0.0233169
R72938 VSS.n6834 VSS.n2937 0.0233169
R72939 VSS.n6834 VSS.n6833 0.0233169
R72940 VSS.n6833 VSS.n6832 0.0233169
R72941 VSS.n6832 VSS.n6811 0.0233169
R72942 VSS.n6828 VSS.n6811 0.0233169
R72943 VSS.n6828 VSS.n6827 0.0233169
R72944 VSS.n6827 VSS.n6826 0.0233169
R72945 VSS.n6826 VSS.n6817 0.0233169
R72946 VSS.n6822 VSS.n6817 0.0233169
R72947 VSS.n6822 VSS.n2652 0.0233169
R72948 VSS.n7000 VSS.n2652 0.0233169
R72949 VSS.n2738 VSS.n2658 0.0233169
R72950 VSS.n2732 VSS.n2658 0.0233169
R72951 VSS.n2732 VSS.n2731 0.0233169
R72952 VSS.n2731 VSS.n2730 0.0233169
R72953 VSS.n2730 VSS.n2662 0.0233169
R72954 VSS.n2726 VSS.n2662 0.0233169
R72955 VSS.n2726 VSS.n2725 0.0233169
R72956 VSS.n2725 VSS.n2724 0.0233169
R72957 VSS.n2724 VSS.n2667 0.0233169
R72958 VSS.n2720 VSS.n2667 0.0233169
R72959 VSS.n2720 VSS.n2719 0.0233169
R72960 VSS.n2719 VSS.n2718 0.0233169
R72961 VSS.n2718 VSS.n2673 0.0233169
R72962 VSS.n2714 VSS.n2673 0.0233169
R72963 VSS.n2714 VSS.n2713 0.0233169
R72964 VSS.n2713 VSS.n2712 0.0233169
R72965 VSS.n2712 VSS.n2679 0.0233169
R72966 VSS.n2708 VSS.n2679 0.0233169
R72967 VSS.n2708 VSS.n2707 0.0233169
R72968 VSS.n2707 VSS.n2706 0.0233169
R72969 VSS.n2706 VSS.n2685 0.0233169
R72970 VSS.n2702 VSS.n2685 0.0233169
R72971 VSS.n2702 VSS.n2701 0.0233169
R72972 VSS.n2701 VSS.n2700 0.0233169
R72973 VSS.n2700 VSS.n2691 0.0233169
R72974 VSS.n2696 VSS.n2691 0.0233169
R72975 VSS.n2696 VSS.n2574 0.0233169
R72976 VSS.n3728 VSS.n3152 0.0231056
R72977 VSS.n6793 VSS.n2945 0.0231056
R72978 VSS.n3783 VSS.n3182 0.0231056
R72979 VSS.n6794 VSS.n2927 0.0231056
R72980 VSS.n1373 VSS.n1365 0.0228944
R72981 VSS.n8396 VSS.n1622 0.0228944
R72982 VSS.n7246 VSS.n7245 0.0227859
R72983 VSS.n7070 VSS.n7068 0.0227859
R72984 VSS.n7076 VSS.n7075 0.0227859
R72985 VSS.n7097 VSS.n7057 0.0227859
R72986 VSS.n7098 VSS.n7055 0.0227859
R72987 VSS.n7075 VSS.n7074 0.0227859
R72988 VSS.n7264 VSS.n2474 0.0227859
R72989 VSS.n2561 VSS.n2560 0.0227859
R72990 VSS.n7158 VSS.n2555 0.0227859
R72991 VSS.n2560 VSS.n2559 0.0227859
R72992 VSS.n7161 VSS.n7160 0.0227859
R72993 VSS.n7261 VSS.n7260 0.0227859
R72994 VSS.n2493 VSS.n2482 0.0227859
R72995 VSS.n7248 VSS.n2503 0.0227859
R72996 VSS.n8083 VSS.n8081 0.0227859
R72997 VSS.n8082 VSS.n1547 0.0227859
R72998 VSS.n8603 VSS.n1545 0.0227859
R72999 VSS.n8599 VSS.n8598 0.0227859
R73000 VSS.n8593 VSS.n8592 0.0227859
R73001 VSS.n8586 VSS.n8575 0.0227859
R73002 VSS.n8580 VSS.n8577 0.0227859
R73003 VSS.n8591 VSS.n8574 0.0227859
R73004 VSS.n8585 VSS.n8576 0.0227859
R73005 VSS.n8596 VSS.n8595 0.0227859
R73006 VSS.n8606 VSS.n8605 0.0227859
R73007 VSS.n8085 VSS.n8084 0.0227859
R73008 VSS.n8081 VSS.n8080 0.0227859
R73009 VSS.n7123 VSS.n2589 0.0227859
R73010 VSS.n7120 VSS.n7119 0.0227859
R73011 VSS.n2596 VSS.n2593 0.0227859
R73012 VSS.n7111 VSS.n7110 0.0227859
R73013 VSS.n7105 VSS.n7104 0.0227859
R73014 VSS.n7051 VSS.n7050 0.0227859
R73015 VSS.n2588 VSS.n1557 0.0227859
R73016 VSS.n7122 VSS.n2591 0.0227859
R73017 VSS.n7110 VSS.n2598 0.0227859
R73018 VSS.n7107 VSS.n2602 0.0227859
R73019 VSS.n7053 VSS.n2604 0.0227859
R73020 VSS.n7116 VSS.n2593 0.0227859
R73021 VSS.n8602 VSS.n8601 0.0227859
R73022 VSS.n2477 VSS.n2474 0.0227859
R73023 VSS.n7070 VSS.n7069 0.0227859
R73024 VSS.n3738 VSS.n3142 0.0226831
R73025 VSS.n3763 VSS.n3172 0.0226831
R73026 VSS.n4459 VSS.n4449 0.0224718
R73027 VSS.n5117 VSS.n4425 0.0224718
R73028 VSS.n8572 VSS.n1455 0.0222606
R73029 VSS.n1549 VSS.n1488 0.0222606
R73030 VSS.n6574 VSS.n6573 0.021937
R73031 VSS.n9594 VSS.n9593 0.021937
R73032 DVSS VSS.n5098 0.021875
R73033 DVSS VSS.n4941 0.021875
R73034 DVSS VSS.n4231 0.021875
R73035 VSS.n6098 DVSS 0.021875
R73036 VSS.n6010 DVSS 0.021875
R73037 VSS.n3765 DVSS 0.021875
R73038 VSS.n5859 DVSS 0.021875
R73039 DVSS VSS.n6836 0.021875
R73040 VSS.n2711 DVSS 0.021875
R73041 VSS.n5670 VSS.n4244 0.021838
R73042 VSS.n3746 VSS.n3159 0.021838
R73043 VSS.n4263 VSS.n4242 0.021838
R73044 VSS.n3747 VSS.n3189 0.021838
R73045 VSS.n8584 VSS.n1118 0.0215827
R73046 VSS.n8590 VSS.n1400 0.0215827
R73047 VSS.n8604 VSS.n1528 0.0215827
R73048 VSS.n8086 VSS.n2108 0.0215827
R73049 VSS.n5710 VSS.n4222 0.0214155
R73050 VSS.n3743 VSS.n3139 0.0214155
R73051 VSS.n5711 VSS.n4021 0.0214155
R73052 VSS.n3753 VSS.n3169 0.0214155
R73053 VSS.n1218 VSS.n1216 0.0212692
R73054 VSS.n1216 VSS.n1214 0.0212692
R73055 VSS.n1214 VSS.n1212 0.0212692
R73056 VSS.n1212 VSS.n1210 0.0212692
R73057 VSS.n1210 VSS.n1207 0.0212692
R73058 VSS.n1207 VSS.n1206 0.0212692
R73059 VSS.n1206 VSS.n1204 0.0212692
R73060 VSS.n1204 VSS.n1202 0.0212692
R73061 VSS.n1202 VSS.n1200 0.0212692
R73062 VSS.n1200 VSS.n1198 0.0212692
R73063 VSS.n1198 VSS.n1196 0.0212692
R73064 VSS.n1196 VSS.n1194 0.0212692
R73065 VSS.n1194 VSS.n1191 0.0212692
R73066 VSS.n1191 VSS.n1190 0.0212692
R73067 VSS.n1190 VSS.n1188 0.0212692
R73068 VSS.n1188 VSS.n1186 0.0212692
R73069 VSS.n1186 VSS.n1184 0.0212692
R73070 VSS.n1184 VSS.n1182 0.0212692
R73071 VSS.n1182 VSS.n1180 0.0212692
R73072 VSS.n1180 VSS.n1177 0.0212692
R73073 VSS.n1177 VSS.n1176 0.0212692
R73074 VSS.n1176 VSS.n1174 0.0212692
R73075 VSS.n1174 VSS.n1172 0.0212692
R73076 VSS.n1172 VSS.n1170 0.0212692
R73077 VSS.n1170 VSS.n757 0.0212692
R73078 VSS.n9457 VSS.n757 0.0212692
R73079 VSS.n9457 VSS.n9456 0.0212692
R73080 VSS.n9379 VSS.n759 0.0212692
R73081 VSS.n9382 VSS.n9379 0.0212692
R73082 VSS.n9384 VSS.n9382 0.0212692
R73083 VSS.n9386 VSS.n9384 0.0212692
R73084 VSS.n9388 VSS.n9386 0.0212692
R73085 VSS.n9390 VSS.n9388 0.0212692
R73086 VSS.n9392 VSS.n9390 0.0212692
R73087 VSS.n9393 VSS.n9392 0.0212692
R73088 VSS.n9396 VSS.n9393 0.0212692
R73089 VSS.n9398 VSS.n9396 0.0212692
R73090 VSS.n9400 VSS.n9398 0.0212692
R73091 VSS.n9402 VSS.n9400 0.0212692
R73092 VSS.n9404 VSS.n9402 0.0212692
R73093 VSS.n9406 VSS.n9404 0.0212692
R73094 VSS.n9408 VSS.n9406 0.0212692
R73095 VSS.n9409 VSS.n9408 0.0212692
R73096 VSS.n9412 VSS.n9409 0.0212692
R73097 VSS.n9414 VSS.n9412 0.0212692
R73098 VSS.n9416 VSS.n9414 0.0212692
R73099 VSS.n9418 VSS.n9416 0.0212692
R73100 VSS.n9420 VSS.n9418 0.0212692
R73101 VSS.n9422 VSS.n9420 0.0212692
R73102 VSS.n9424 VSS.n9422 0.0212692
R73103 VSS.n9425 VSS.n9424 0.0212692
R73104 VSS.n9428 VSS.n9425 0.0212692
R73105 VSS.n9430 VSS.n9428 0.0212692
R73106 VSS.n9431 VSS.n9430 0.0212692
R73107 VSS.n2370 VSS.n2369 0.0212692
R73108 VSS.n9436 VSS.n9375 0.0212692
R73109 VSS.n2282 VSS.n2280 0.0212692
R73110 VSS.n2284 VSS.n2282 0.0212692
R73111 VSS.n2286 VSS.n2284 0.0212692
R73112 VSS.n2287 VSS.n2286 0.0212692
R73113 VSS.n2290 VSS.n2287 0.0212692
R73114 VSS.n2292 VSS.n2290 0.0212692
R73115 VSS.n2294 VSS.n2292 0.0212692
R73116 VSS.n2296 VSS.n2294 0.0212692
R73117 VSS.n2298 VSS.n2296 0.0212692
R73118 VSS.n2300 VSS.n2298 0.0212692
R73119 VSS.n2302 VSS.n2300 0.0212692
R73120 VSS.n2303 VSS.n2302 0.0212692
R73121 VSS.n2306 VSS.n2303 0.0212692
R73122 VSS.n2308 VSS.n2306 0.0212692
R73123 VSS.n2310 VSS.n2308 0.0212692
R73124 VSS.n2312 VSS.n2310 0.0212692
R73125 VSS.n2314 VSS.n2312 0.0212692
R73126 VSS.n2316 VSS.n2314 0.0212692
R73127 VSS.n2317 VSS.n2316 0.0212692
R73128 VSS.n2320 VSS.n2317 0.0212692
R73129 VSS.n2322 VSS.n2320 0.0212692
R73130 VSS.n2324 VSS.n2322 0.0212692
R73131 VSS.n2326 VSS.n2324 0.0212692
R73132 VSS.n2328 VSS.n2326 0.0212692
R73133 VSS.n2329 VSS.n2328 0.0212692
R73134 VSS.n7891 VSS.n2329 0.0212692
R73135 VSS.n7891 VSS.n7890 0.0212692
R73136 VSS.n2426 VSS.n2424 0.0212692
R73137 VSS.n2424 VSS.n2421 0.0212692
R73138 VSS.n2421 VSS.n2420 0.0212692
R73139 VSS.n2420 VSS.n2418 0.0212692
R73140 VSS.n2418 VSS.n2416 0.0212692
R73141 VSS.n2416 VSS.n2414 0.0212692
R73142 VSS.n2414 VSS.n2412 0.0212692
R73143 VSS.n2412 VSS.n2410 0.0212692
R73144 VSS.n2410 VSS.n2407 0.0212692
R73145 VSS.n2407 VSS.n2406 0.0212692
R73146 VSS.n2406 VSS.n2404 0.0212692
R73147 VSS.n2404 VSS.n2402 0.0212692
R73148 VSS.n2402 VSS.n2400 0.0212692
R73149 VSS.n2400 VSS.n2398 0.0212692
R73150 VSS.n2398 VSS.n2396 0.0212692
R73151 VSS.n2396 VSS.n2394 0.0212692
R73152 VSS.n2394 VSS.n2391 0.0212692
R73153 VSS.n2391 VSS.n2390 0.0212692
R73154 VSS.n2390 VSS.n2388 0.0212692
R73155 VSS.n2388 VSS.n2386 0.0212692
R73156 VSS.n2386 VSS.n2384 0.0212692
R73157 VSS.n2384 VSS.n2382 0.0212692
R73158 VSS.n2382 VSS.n2380 0.0212692
R73159 VSS.n2380 VSS.n2378 0.0212692
R73160 VSS.n2378 VSS.n2375 0.0212692
R73161 VSS.n2375 VSS.n2374 0.0212692
R73162 VSS.n2374 VSS.n2372 0.0212692
R73163 VSS.n9901 VSS.n11 0.0208631
R73164 VSS.n9901 VSS.n9900 0.0208631
R73165 VSS.n8056 VSS.n1451 0.0207817
R73166 VSS.n8064 VSS.n1484 0.0207817
R73167 VSS.n4855 VSS.n4489 0.0205704
R73168 VSS.n3735 VSS.n3155 0.0205704
R73169 VSS.n5086 VSS.n4486 0.0205704
R73170 VSS.n3769 VSS.n3185 0.0205704
R73171 VSS.n7230 VSS.n2499 0.020197
R73172 VSS.n7231 VSS.n7230 0.020197
R73173 VSS.n7206 VSS.n2499 0.020197
R73174 VSS.n7207 VSS.n7206 0.020197
R73175 VSS.n7174 VSS.n2499 0.020197
R73176 VSS.n7175 VSS.n7174 0.020197
R73177 VSS.n4866 VSS.n4851 0.0201479
R73178 VSS.n3731 VSS.n3145 0.0201479
R73179 VSS.n6784 VSS.n2951 0.0201479
R73180 VSS.n4864 VSS.n4497 0.0201479
R73181 VSS.n3777 VSS.n3175 0.0201479
R73182 VSS.n6785 VSS.n2933 0.0201479
R73183 VSS.n7207 VSS.n7204 0.0198883
R73184 VSS.n7210 VSS.n7207 0.0198883
R73185 VSS.n7232 VSS.n7231 0.0198883
R73186 VSS.n7231 VSS.n2519 0.0198883
R73187 VSS.n7180 VSS.n7175 0.0198883
R73188 VSS.n7175 VSS.n7173 0.0198883
R73189 VSS.n8542 VSS.n1616 0.0198883
R73190 VSS.n1616 VSS.n1613 0.0198883
R73191 VSS.n8062 VSS.n8059 0.0198883
R73192 VSS.n8059 VSS.n8057 0.0198883
R73193 VSS.n8823 VSS.n1362 0.0198883
R73194 VSS.n8823 VSS.n8822 0.0198883
R73195 VSS.n2276 VSS.n2173 0.019811
R73196 VSS.n1164 VSS.n1151 0.019811
R73197 VSS.n3727 VSS.n3146 0.0197254
R73198 VSS.n6796 VSS.n2952 0.0197254
R73199 VSS.n3785 VSS.n3176 0.0197254
R73200 VSS.n6797 VSS.n2934 0.0197254
R73201 VSS.n2289 VSS.n2288 0.0196339
R73202 VSS.n2305 VSS.n2304 0.0196339
R73203 VSS.n2319 VSS.n2318 0.0196339
R73204 VSS.n7892 VSS.n2169 0.0196339
R73205 VSS.n2425 VSS.n2169 0.0196339
R73206 VSS.n2423 VSS.n2422 0.0196339
R73207 VSS.n2409 VSS.n2408 0.0196339
R73208 VSS.n2393 VSS.n2392 0.0196339
R73209 VSS.n2377 VSS.n2376 0.0196339
R73210 VSS.n2792 VSS.n2791 0.0196339
R73211 VSS.n9604 VSS.n431 0.0196339
R73212 VSS.n9604 VSS.n432 0.0196339
R73213 VSS.n9599 VSS.n440 0.0196339
R73214 VSS.n9599 VSS.n441 0.0196339
R73215 VSS.n9591 VSS.n488 0.0196339
R73216 VSS.n9591 VSS.n489 0.0196339
R73217 VSS.n9586 VSS.n497 0.0196339
R73218 VSS.n9586 VSS.n498 0.0196339
R73219 VSS.n9578 VSS.n530 0.0196339
R73220 VSS.n9578 VSS.n531 0.0196339
R73221 VSS.n9573 VSS.n538 0.0196339
R73222 VSS.n1209 VSS.n1208 0.0196339
R73223 VSS.n1193 VSS.n1192 0.0196339
R73224 VSS.n1179 VSS.n1178 0.0196339
R73225 VSS.n9458 VSS.n756 0.0196339
R73226 VSS.n758 VSS.n756 0.0196339
R73227 VSS.n9381 VSS.n9380 0.0196339
R73228 VSS.n9395 VSS.n9394 0.0196339
R73229 VSS.n9411 VSS.n9410 0.0196339
R73230 VSS.n9427 VSS.n9426 0.0196339
R73231 VSS.n2301 VSS.n2160 0.0194567
R73232 VSS.n2425 VSS.n1850 0.0194567
R73233 VSS.n1195 VSS.n748 0.0194567
R73234 VSS.n758 VSS.n697 0.0194567
R73235 VSS.n3739 VSS.n3156 0.0193028
R73236 VSS.n6617 VSS.n6616 0.0193028
R73237 VSS.n3761 VSS.n3186 0.0193028
R73238 VSS.n6608 VSS.n6607 0.0193028
R73239 VSS.n8854 VSS.n1291 0.0192795
R73240 VSS.n8843 VSS.n1315 0.0192795
R73241 VSS.n8404 VSS.n1658 0.0192795
R73242 VSS.n8561 VSS.n8560 0.0192795
R73243 VSS.n2790 VSS.n2789 0.0191034
R73244 VSS.n9574 VSS.n536 0.0191034
R73245 VSS.n2321 VSS.n2145 0.0191024
R73246 VSS.n2405 VSS.n1855 0.0191024
R73247 VSS.n1175 VSS.n732 0.0191024
R73248 VSS.n9397 VSS.n701 0.0191024
R73249 VSS.n4458 VSS.n4456 0.0190915
R73250 VSS.n5119 VSS.n4432 0.0190915
R73251 VSS.n5657 VSS.n4250 0.0188803
R73252 VSS.n5656 VSS.n4268 0.0188803
R73253 VSS.n8581 VSS.n1119 0.018748
R73254 VSS.n2285 VSS.n2152 0.018748
R73255 VSS.n2379 VSS.n1840 0.018748
R73256 VSS.n8587 VSS.n1419 0.018748
R73257 VSS.n8607 VSS.n1539 0.018748
R73258 VSS.n8087 VSS.n8079 0.018748
R73259 VSS.n6259 VSS.n3839 0.018748
R73260 VSS.n4156 VSS.n410 0.018748
R73261 VSS.n1211 VSS.n739 0.018748
R73262 VSS.n9423 VSS.n687 0.018748
R73263 VSS.n9899 VSS.n14 0.0184577
R73264 VSS.n5667 VSS.n4248 0.0184577
R73265 VSS.n3160 VSS.n3138 0.0184577
R73266 VSS.n4434 VSS.n4433 0.0184577
R73267 VSS.n5665 VSS.n5664 0.0184577
R73268 VSS.n3168 VSS.n3167 0.0184577
R73269 VSS.n2389 VSS.n1843 0.0183937
R73270 VSS.n9413 VSS.n690 0.0183937
R73271 VSS.n2467 VSS.n2466 0.0181271
R73272 VSS.n9453 VSS.n9452 0.0181271
R73273 VSS.n2395 VSS.n1858 0.0180394
R73274 VSS.n9407 VSS.n704 0.0180394
R73275 VSS.n4223 VSS.n4175 0.0180352
R73276 VSS.n3742 VSS.n3158 0.0180352
R73277 VSS.n5713 VSS.n4019 0.0180352
R73278 VSS.n3755 VSS.n3188 0.0180352
R73279 VSS.n7147 VSS.n7146 0.0178648
R73280 VSS.n6068 VSS.n6046 0.0177222
R73281 VSS.n6075 VSS.n6038 0.0177222
R73282 VSS.n6079 VSS.n4071 0.0177222
R73283 VSS.n5957 VSS.n5904 0.0177222
R73284 VSS.n5949 VSS.n5915 0.0177222
R73285 VSS.n5941 VSS.n5922 0.0177222
R73286 VSS.n5934 VSS.n5929 0.0177222
R73287 VSS.n6294 VSS.n3809 0.0177222
R73288 VSS.n6301 VSS.n3800 0.0177222
R73289 VSS.n6305 VSS.n3717 0.0177222
R73290 VSS.n6317 VSS.n3705 0.0177222
R73291 VSS.n6323 VSS.n3696 0.0177222
R73292 VSS.n6330 VSS.n3687 0.0177222
R73293 VSS.n6338 VSS.n3683 0.0177222
R73294 VSS.n6588 VSS.n3215 0.0177222
R73295 VSS.n6594 VSS.n3206 0.0177222
R73296 VSS.n6601 VSS.n3197 0.0177222
R73297 VSS.n6605 VSS.n3192 0.0177222
R73298 VSS.n6623 VSS.n3127 0.0177222
R73299 VSS.n6629 VSS.n3119 0.0177222
R73300 VSS.n6638 VSS.n3115 0.0177222
R73301 VSS.n3667 VSS.n3656 0.0177222
R73302 VSS.n5786 VSS.n5758 0.0177222
R73303 VSS.n5792 VSS.n5749 0.0177222
R73304 VSS.n5799 VSS.n5740 0.0177222
R73305 VSS.n5891 VSS.n5734 0.0177222
R73306 VSS.n6765 VSS.n2960 0.0177222
R73307 VSS.n6757 VSS.n2968 0.0177222
R73308 VSS.n6653 VSS.n3112 0.0177222
R73309 VSS.n6661 VSS.n3108 0.0177222
R73310 VSS.n6980 VSS.n2759 0.0177222
R73311 VSS.n6986 VSS.n2750 0.0177222
R73312 VSS.n6993 VSS.n2741 0.0177222
R73313 VSS.n6997 VSS.n2655 0.0177222
R73314 VSS.n7009 VSS.n2643 0.0177222
R73315 VSS.n7015 VSS.n2634 0.0177222
R73316 VSS.n7022 VSS.n2625 0.0177222
R73317 VSS.n7030 VSS.n2621 0.0177222
R73318 VSS.n2291 VSS.n2157 0.017685
R73319 VSS.n2373 VSS.n1862 0.017685
R73320 VSS.n1205 VSS.n745 0.017685
R73321 VSS.n9429 VSS.n708 0.017685
R73322 VSS.n3724 VSS.n3148 0.0176127
R73323 VSS.n6806 VSS.n2939 0.0176127
R73324 VSS.n3791 VSS.n3178 0.0176127
R73325 VSS.n6839 VSS.n2936 0.0176127
R73326 VSS.n8045 VSS.n1137 0.0175079
R73327 VSS.n8050 VSS.n1406 0.0175079
R73328 VSS.n8069 VSS.n1534 0.0175079
R73329 VSS.n8075 VSS.n2125 0.0175079
R73330 VSS.n2315 VSS.n2163 0.0173307
R73331 VSS.n2411 VSS.n1847 0.0173307
R73332 VSS.n1181 VSS.n751 0.0173307
R73333 VSS.n9391 VSS.n694 0.0173307
R73334 VSS.n4856 VSS.n4853 0.0171901
R73335 VSS.n3734 VSS.n3143 0.0171901
R73336 VSS.n6775 VSS.n2949 0.0171901
R73337 VSS.n5085 VSS.n4492 0.0171901
R73338 VSS.n3771 VSS.n3173 0.0171901
R73339 VSS.n6776 VSS.n2931 0.0171901
R73340 VSS.n9904 VSS.n9903 0.0171667
R73341 VSS.n7884 VSS.n7883 0.0171667
R73342 VSS.n7883 VSS.n761 0.0171667
R73343 VSS.n5081 VSS.n4510 0.0170278
R73344 VSS.n4971 VSS.n4510 0.0170278
R73345 VSS.n5652 VSS.n4277 0.0170278
R73346 VSS.n4914 VSS.n4277 0.0170278
R73347 VSS.n5729 VSS.n4115 0.0170278
R73348 VSS.n5729 VSS.n5728 0.0170278
R73349 VSS.n6079 VSS.n5899 0.0170278
R73350 VSS.n5903 VSS.n5899 0.0170278
R73351 VSS.n6305 VSS.n3711 0.0170278
R73352 VSS.n6314 VSS.n3711 0.0170278
R73353 VSS.n6605 VSS.n3133 0.0170278
R73354 VSS.n6620 VSS.n3133 0.0170278
R73355 VSS.n5892 VSS.n5891 0.0170278
R73356 VSS.n5892 VSS.n2959 0.0170278
R73357 VSS.n6997 VSS.n2649 0.0170278
R73358 VSS.n7006 VSS.n2649 0.0170278
R73359 VSS.n2272 VSS.n2270 0.0169764
R73360 VSS.n2307 VSS.n2148 0.0169764
R73361 VSS.n2419 VSS.n1852 0.0169764
R73362 VSS.n8949 VSS.n1224 0.0169764
R73363 VSS.n1189 VSS.n735 0.0169764
R73364 VSS.n9383 VSS.n698 0.0169764
R73365 VSS.n4867 VSS.n4858 0.0167676
R73366 VSS.n3732 VSS.n3153 0.0167676
R73367 VSS.n6781 VSS.n2946 0.0167676
R73368 VSS.n4862 VSS.n4501 0.0167676
R73369 VSS.n3775 VSS.n3183 0.0167676
R73370 VSS.n6782 VSS.n2928 0.0167676
R73371 VSS.n2299 VSS.n2149 0.016622
R73372 VSS.n1197 VSS.n736 0.016622
R73373 VSS.n3726 VSS.n3151 0.0163451
R73374 VSS.n2953 VSS.n2944 0.0163451
R73375 VSS.n1465 VSS.n1460 0.0163451
R73376 VSS.n8711 VSS.n1463 0.0163451
R73377 VSS.n3787 VSS.n3181 0.0163451
R73378 VSS.n6799 VSS.n2926 0.0163451
R73379 VSS.n1498 VSS.n1493 0.0163451
R73380 VSS.n8685 VSS.n1496 0.0163451
R73381 VSS.n6427 VSS.n3116 0.0162677
R73382 VSS.n6544 VSS.n3216 0.0162677
R73383 VSS.n2323 VSS.n2164 0.0162677
R73384 VSS.n2403 VSS.n1846 0.0162677
R73385 VSS.n6452 VSS.n3120 0.0162677
R73386 VSS.n6506 VSS.n3198 0.0162677
R73387 VSS.n6531 VSS.n3207 0.0162677
R73388 VSS.n4763 VSS.n4727 0.0162677
R73389 VSS.n6252 VSS.n3862 0.0162677
R73390 VSS.n9811 VSS.n172 0.0162677
R73391 VSS.n5475 VSS.n5473 0.0162677
R73392 VSS.n3669 VSS.n3668 0.0162677
R73393 VSS.n1173 VSS.n752 0.0162677
R73394 VSS.n9399 VSS.n693 0.0162677
R73395 VSS.n8058 VSS.n1358 0.0162576
R73396 VSS.n8059 VSS.n8058 0.0162576
R73397 VSS.n1615 VSS.n1358 0.0162576
R73398 VSS.n1616 VSS.n1615 0.0162576
R73399 VSS.n8824 VSS.n1358 0.0162576
R73400 VSS.n8824 VSS.n8823 0.0162576
R73401 VSS.n4967 VSS.n4850 0.0159225
R73402 VSS.n4972 VSS.n4869 0.0159225
R73403 VSS.n4969 VSS.n4849 0.0159225
R73404 VSS.n5019 VSS.n4870 0.0159225
R73405 VSS.n5721 VSS.n5719 0.0159225
R73406 VSS.n3740 VSS.n3141 0.0159225
R73407 VSS.n4508 VSS.n4496 0.0159225
R73408 VSS.n5080 VSS.n4504 0.0159225
R73409 VSS.n4511 VSS.n4495 0.0159225
R73410 VSS.n5083 VSS.n4505 0.0159225
R73411 VSS.n4074 VSS.n4024 0.0159225
R73412 VSS.n3759 VSS.n3171 0.0159225
R73413 VSS.n2283 VSS.n2156 0.0159134
R73414 VSS.n2381 VSS.n1861 0.0159134
R73415 VSS.n6257 VSS.n3851 0.0159134
R73416 VSS.n4153 VSS.n420 0.0159134
R73417 VSS.n1213 VSS.n744 0.0159134
R73418 VSS.n9421 VSS.n707 0.0159134
R73419 VSS.n4457 VSS.n4450 0.0157113
R73420 VSS.n5121 VSS.n4426 0.0157113
R73421 VSS.n79 VSS.n78 0.0155591
R73422 VSS.n2387 VSS.n1859 0.0155591
R73423 VSS.n4628 VSS.n4627 0.0155591
R73424 VSS.n9896 VSS.n22 0.0155591
R73425 VSS.n4391 VSS.n4390 0.0155591
R73426 VSS.n4354 VSS.n4353 0.0155591
R73427 VSS.n4603 VSS.n4602 0.0155591
R73428 VSS.n6264 VSS.n3832 0.0155591
R73429 VSS.n141 VSS.n140 0.0155591
R73430 VSS.n9607 VSS.n422 0.0155591
R73431 VSS.n110 VSS.n109 0.0155591
R73432 VSS.n9415 VSS.n705 0.0155591
R73433 VSS.n5167 VSS.n13 0.0155
R73434 VSS.n5659 VSS.n4258 0.0155
R73435 VSS.n4173 VSS.n4116 0.0155
R73436 VSS.n5727 VSS.n4120 0.0155
R73437 VSS.n4122 VSS.n4119 0.0155
R73438 VSS.n5722 VSS.n4117 0.0155
R73439 VSS.n5725 VSS.n4169 0.0155
R73440 VSS.n4661 VSS.n4430 0.0155
R73441 VSS.n5662 VSS.n5661 0.0155
R73442 VSS.n4076 VSS.n4017 0.0155
R73443 VSS.n4114 VSS.n4025 0.0155
R73444 VSS.n4078 VSS.n4016 0.0155
R73445 VSS.n4111 VSS.n4026 0.0155
R73446 VSS.n4027 VSS.n4015 0.0155
R73447 VSS.n6273 VSS.n6267 0.0155
R73448 VSS.n6280 VSS.n6278 0.0155
R73449 VSS.n6579 VSS.n6577 0.0155
R73450 VSS.n5777 VSS.n5775 0.0155
R73451 VSS.n6971 VSS.n6969 0.0155
R73452 VSS.n7930 VSS.n2166 0.0152047
R73453 VSS.n2397 VSS.n1844 0.0152047
R73454 VSS.n4761 VSS.n4760 0.0152047
R73455 VSS.n6239 VSS.n3857 0.0152047
R73456 VSS.n9807 VSS.n170 0.0152047
R73457 VSS.n5470 VSS.n5438 0.0152047
R73458 VSS.n9498 VSS.n754 0.0152047
R73459 VSS.n9405 VSS.n691 0.0152047
R73460 VSS.n4452 VSS.n16 0.0150775
R73461 VSS.n5668 VSS.n4259 0.0150775
R73462 VSS.n6614 VSS.n6613 0.0150775
R73463 VSS.n5178 VSS.n4438 0.0150775
R73464 VSS.n4266 VSS.n4261 0.0150775
R73465 VSS.n6611 VSS.n3163 0.0150775
R73466 VSS.n5126 VSS.n5125 0.0148662
R73467 VSS.n5123 VSS.n4427 0.0148662
R73468 VSS.n2293 VSS.n2151 0.0148504
R73469 VSS.n1863 VSS.n1839 0.0148504
R73470 VSS.n1203 VSS.n738 0.0148504
R73471 VSS.n709 VSS.n686 0.0148504
R73472 VSS.n4920 VSS.n4254 0.0146549
R73473 VSS.n4919 VSS.n4252 0.0146549
R73474 VSS.n4915 VSS.n4255 0.0146549
R73475 VSS.n4918 VSS.n4251 0.0146549
R73476 VSS.n5718 VSS.n5717 0.0146549
R73477 VSS.n3741 VSS.n3140 0.0146549
R73478 VSS.n5651 VSS.n4272 0.0146549
R73479 VSS.n4278 VSS.n4270 0.0146549
R73480 VSS.n5649 VSS.n4273 0.0146549
R73481 VSS.n5653 VSS.n4269 0.0146549
R73482 VSS.n5715 VSS.n4022 0.0146549
R73483 VSS.n3757 VSS.n3170 0.0146549
R73484 VSS.n7150 VSS.n2571 0.0145346
R73485 VSS.n2569 VSS.n2565 0.0145346
R73486 VSS.n7154 VSS.n2569 0.0145346
R73487 VSS.n2568 VSS.n2567 0.0145346
R73488 VSS.n7155 VSS.n7154 0.0145346
R73489 VSS.n7155 VSS.n2568 0.0145346
R73490 VSS.n7151 VSS.n2565 0.0145346
R73491 VSS.n7146 VSS.n2571 0.0145346
R73492 VSS.n7134 VSS.n7133 0.0145346
R73493 VSS.n7139 VSS.n2575 0.0145346
R73494 VSS.n7133 VSS.n7132 0.0145346
R73495 VSS.n7135 VSS.n2575 0.0145346
R73496 VSS.n2775 VSS.n2774 0.0145346
R73497 VSS.n2776 VSS.n2775 0.0145346
R73498 VSS.n2781 VSS.n2777 0.0145346
R73499 VSS.n2782 VSS.n2780 0.0145346
R73500 VSS.n2585 VSS.n2584 0.0145346
R73501 VSS.n7130 VSS.n2579 0.0145346
R73502 VSS.n2788 VSS.n2777 0.0145346
R73503 VSS.n2584 VSS.n2583 0.0145346
R73504 VSS.n2586 VSS.n2579 0.0145346
R73505 VSS.n2785 VSS.n2780 0.0145346
R73506 VSS.n2790 VSS.n2776 0.0145346
R73507 VSS.n2794 VSS.n2774 0.0145346
R73508 VSS.n4637 VSS.n4635 0.0145346
R73509 VSS.n4635 VSS.n4634 0.0145346
R73510 VSS.n4673 VSS.n4640 0.0145346
R73511 VSS.n4640 VSS.n4633 0.0145346
R73512 VSS.n4643 VSS.n4641 0.0145346
R73513 VSS.n4641 VSS.n4632 0.0145346
R73514 VSS.n4669 VSS.n4644 0.0145346
R73515 VSS.n4645 VSS.n4644 0.0145346
R73516 VSS.n4648 VSS.n4647 0.0145346
R73517 VSS.n4649 VSS.n4648 0.0145346
R73518 VSS.n4665 VSS.n4650 0.0145346
R73519 VSS.n4651 VSS.n4650 0.0145346
R73520 VSS.n4654 VSS.n4653 0.0145346
R73521 VSS.n4655 VSS.n4654 0.0145346
R73522 VSS.n4662 VSS.n4656 0.0145346
R73523 VSS.n4660 VSS.n4658 0.0145346
R73524 VSS.n4658 VSS.n4657 0.0145346
R73525 VSS.n9900 VSS.n12 0.0145346
R73526 VSS.n17 VSS.n15 0.0145346
R73527 VSS.n19 VSS.n15 0.0145346
R73528 VSS.n24 VSS.n21 0.0145346
R73529 VSS.n26 VSS.n24 0.0145346
R73530 VSS.n31 VSS.n23 0.0145346
R73531 VSS.n28 VSS.n23 0.0145346
R73532 VSS.n160 VSS.n159 0.0145346
R73533 VSS.n159 VSS.n158 0.0145346
R73534 VSS.n156 VSS.n155 0.0145346
R73535 VSS.n155 VSS.n154 0.0145346
R73536 VSS.n164 VSS.n153 0.0145346
R73537 VSS.n153 VSS.n152 0.0145346
R73538 VSS.n150 VSS.n149 0.0145346
R73539 VSS.n149 VSS.n148 0.0145346
R73540 VSS.n9819 VSS.n9818 0.0145346
R73541 VSS.n9818 VSS.n147 0.0145346
R73542 VSS.n4637 VSS.n4636 0.0145346
R73543 VSS.n4674 VSS.n4673 0.0145346
R73544 VSS.n4643 VSS.n4642 0.0145346
R73545 VSS.n4670 VSS.n4669 0.0145346
R73546 VSS.n4647 VSS.n4646 0.0145346
R73547 VSS.n4666 VSS.n4665 0.0145346
R73548 VSS.n4653 VSS.n4652 0.0145346
R73549 VSS.n4660 VSS.n4659 0.0145346
R73550 VSS.n18 VSS.n17 0.0145346
R73551 VSS.n9897 VSS.n21 0.0145346
R73552 VSS.n31 VSS.n27 0.0145346
R73553 VSS.n160 VSS.n29 0.0145346
R73554 VSS.n157 VSS.n156 0.0145346
R73555 VSS.n4639 VSS.n4634 0.0145346
R73556 VSS.n4642 VSS.n4633 0.0145346
R73557 VSS.n4671 VSS.n4632 0.0145346
R73558 VSS.n4646 VSS.n4645 0.0145346
R73559 VSS.n4667 VSS.n4649 0.0145346
R73560 VSS.n4652 VSS.n4651 0.0145346
R73561 VSS.n4663 VSS.n4655 0.0145346
R73562 VSS.n4659 VSS.n4656 0.0145346
R73563 VSS.n4657 VSS.n11 0.0145346
R73564 VSS.n18 VSS.n12 0.0145346
R73565 VSS.n9898 VSS.n19 0.0145346
R73566 VSS.n27 VSS.n26 0.0145346
R73567 VSS.n9895 VSS.n28 0.0145346
R73568 VSS.n158 VSS.n157 0.0145346
R73569 VSS.n162 VSS.n154 0.0145346
R73570 VSS.n9816 VSS.n147 0.0145346
R73571 VSS.n9820 VSS.n9819 0.0145346
R73572 VSS.n2614 VSS.n2613 0.0145346
R73573 VSS.n7044 VSS.n2610 0.0145346
R73574 VSS.n7034 VSS.n2618 0.0145346
R73575 VSS.n7035 VSS.n7034 0.0145346
R73576 VSS.n7037 VSS.n7036 0.0145346
R73577 VSS.n537 VSS.n534 0.0145346
R73578 VSS.n9572 VSS.n534 0.0145346
R73579 VSS.n9574 VSS.n537 0.0145346
R73580 VSS.n7046 VSS.n2614 0.0145346
R73581 VSS.n2615 VSS.n2610 0.0145346
R73582 VSS.n9572 VSS.n9571 0.0145346
R73583 VSS.n7038 VSS.n7035 0.0145346
R73584 VSS.n7038 VSS.n7037 0.0145346
R73585 VSS.n164 VSS.n163 0.0145346
R73586 VSS.n151 VSS.n150 0.0145346
R73587 VSS.n152 VSS.n151 0.0145346
R73588 VSS.n166 VSS.n148 0.0145346
R73589 VSS.n7043 VSS.n2618 0.0145346
R73590 VSS.n2313 VSS.n2146 0.0144961
R73591 VSS.n2413 VSS.n1854 0.0144961
R73592 VSS.n1183 VSS.n733 0.0144961
R73593 VSS.n9389 VSS.n700 0.0144961
R73594 VSS.n3725 VSS.n3150 0.0142324
R73595 VSS.n6803 VSS.n2943 0.0142324
R73596 VSS.n3789 VSS.n3180 0.0142324
R73597 VSS.n6801 VSS.n2925 0.0142324
R73598 VSS.n2309 VSS.n2161 0.0141417
R73599 VSS.n2417 VSS.n1849 0.0141417
R73600 VSS.n1187 VSS.n749 0.0141417
R73601 VSS.n9385 VSS.n696 0.0141417
R73602 VSS.n5170 VSS.n14 0.0140606
R73603 VSS.n5126 VSS.n4451 0.0140606
R73604 VSS.n4871 VSS.n4868 0.0140606
R73605 VSS.n4256 VSS.n4250 0.0140606
R73606 VSS.n5720 VSS.n4173 0.0140606
R73607 VSS.n5908 VSS.n5907 0.0140606
R73608 VSS.n5956 VSS.n5954 0.0140606
R73609 VSS.n5955 VSS.n5909 0.0140606
R73610 VSS.n5958 VSS.n5902 0.0140606
R73611 VSS.n6311 VSS.n3706 0.0140606
R73612 VSS.n6316 VSS.n3710 0.0140606
R73613 VSS.n6315 VSS.n3707 0.0140606
R73614 VSS.n3709 VSS.n3708 0.0140606
R73615 VSS.n6616 VSS.n3134 0.0140606
R73616 VSS.n6617 VSS.n3128 0.0140606
R73617 VSS.n6622 VSS.n3132 0.0140606
R73618 VSS.n6621 VSS.n3129 0.0140606
R73619 VSS.n3131 VSS.n3130 0.0140606
R73620 VSS.n5879 VSS.n2961 0.0140606
R73621 VSS.n6764 VSS.n6762 0.0140606
R73622 VSS.n6763 VSS.n2962 0.0140606
R73623 VSS.n6766 VSS.n2958 0.0140606
R73624 VSS.n7003 VSS.n2644 0.0140606
R73625 VSS.n7008 VSS.n2648 0.0140606
R73626 VSS.n7007 VSS.n2645 0.0140606
R73627 VSS.n2647 VSS.n2646 0.0140606
R73628 VSS.n8814 VSS.n8813 0.0140606
R73629 VSS.n8813 VSS.n1375 0.0140606
R73630 VSS.n1384 VSS.n1382 0.0140606
R73631 VSS.n1382 VSS.n1374 0.0140606
R73632 VSS.n1371 VSS.n1367 0.0140606
R73633 VSS.n1372 VSS.n1371 0.0140606
R73634 VSS.n1381 VSS.n1379 0.0140606
R73635 VSS.n1379 VSS.n1370 0.0140606
R73636 VSS.n1461 VSS.n1453 0.0140606
R73637 VSS.n1473 VSS.n1472 0.0140606
R73638 VSS.n1473 VSS.n1450 0.0140606
R73639 VSS.n8694 VSS.n1471 0.0140606
R73640 VSS.n1471 VSS.n1449 0.0140606
R73641 VSS.n8696 VSS.n1470 0.0140606
R73642 VSS.n1470 VSS.n1448 0.0140606
R73643 VSS.n8698 VSS.n1469 0.0140606
R73644 VSS.n1469 VSS.n1447 0.0140606
R73645 VSS.n8700 VSS.n1446 0.0140606
R73646 VSS.n8703 VSS.n8702 0.0140606
R73647 VSS.n8703 VSS.n1456 0.0140606
R73648 VSS.n8705 VSS.n8704 0.0140606
R73649 VSS.n8705 VSS.n1457 0.0140606
R73650 VSS.n8707 VSS.n8706 0.0140606
R73651 VSS.n8707 VSS.n1458 0.0140606
R73652 VSS.n8709 VSS.n8708 0.0140606
R73653 VSS.n8709 VSS.n1459 0.0140606
R73654 VSS.n2464 VSS.n2463 0.0140606
R73655 VSS.n2448 VSS.n2446 0.0140606
R73656 VSS.n9080 VSS.n983 0.0140606
R73657 VSS.n9081 VSS.n9080 0.0140606
R73658 VSS.n9083 VSS.n984 0.0140606
R73659 VSS.n9084 VSS.n9083 0.0140606
R73660 VSS.n9086 VSS.n985 0.0140606
R73661 VSS.n9087 VSS.n9086 0.0140606
R73662 VSS.n9089 VSS.n986 0.0140606
R73663 VSS.n9090 VSS.n9089 0.0140606
R73664 VSS.n9092 VSS.n987 0.0140606
R73665 VSS.n9093 VSS.n9092 0.0140606
R73666 VSS.n9095 VSS.n988 0.0140606
R73667 VSS.n9096 VSS.n9095 0.0140606
R73668 VSS.n9098 VSS.n989 0.0140606
R73669 VSS.n9099 VSS.n9098 0.0140606
R73670 VSS.n9101 VSS.n990 0.0140606
R73671 VSS.n9102 VSS.n9101 0.0140606
R73672 VSS.n9104 VSS.n991 0.0140606
R73673 VSS.n9105 VSS.n9104 0.0140606
R73674 VSS.n9107 VSS.n992 0.0140606
R73675 VSS.n9108 VSS.n9107 0.0140606
R73676 VSS.n9110 VSS.n993 0.0140606
R73677 VSS.n9111 VSS.n9110 0.0140606
R73678 VSS.n9113 VSS.n994 0.0140606
R73679 VSS.n9240 VSS.n9231 0.0140606
R73680 VSS.n9231 VSS.n875 0.0140606
R73681 VSS.n9241 VSS.n9232 0.0140606
R73682 VSS.n9232 VSS.n876 0.0140606
R73683 VSS.n9242 VSS.n9233 0.0140606
R73684 VSS.n9233 VSS.n877 0.0140606
R73685 VSS.n9243 VSS.n9234 0.0140606
R73686 VSS.n9234 VSS.n878 0.0140606
R73687 VSS.n9244 VSS.n9235 0.0140606
R73688 VSS.n9235 VSS.n879 0.0140606
R73689 VSS.n9245 VSS.n9236 0.0140606
R73690 VSS.n9236 VSS.n880 0.0140606
R73691 VSS.n9246 VSS.n9237 0.0140606
R73692 VSS.n9237 VSS.n881 0.0140606
R73693 VSS.n9247 VSS.n9238 0.0140606
R73694 VSS.n9238 VSS.n882 0.0140606
R73695 VSS.n9248 VSS.n9239 0.0140606
R73696 VSS.n9239 VSS.n883 0.0140606
R73697 VSS.n9252 VSS.n9251 0.0140606
R73698 VSS.n9252 VSS.n884 0.0140606
R73699 VSS.n9254 VSS.n886 0.0140606
R73700 VSS.n9255 VSS.n9254 0.0140606
R73701 VSS.n9249 VSS.n766 0.0140606
R73702 VSS.n768 VSS.n767 0.0140606
R73703 VSS.n9448 VSS.n765 0.0140606
R73704 VSS.n9447 VSS.n763 0.0140606
R73705 VSS.n4871 VSS.n4851 0.0140606
R73706 VSS.n4257 VSS.n4256 0.0140606
R73707 VSS.n5721 VSS.n5720 0.0140606
R73708 VSS.n3137 VSS.n3134 0.0140606
R73709 VSS.n8815 VSS.n8814 0.0140606
R73710 VSS.n1383 VSS.n1375 0.0140606
R73711 VSS.n1384 VSS.n1383 0.0140606
R73712 VSS.n1385 VSS.n1374 0.0140606
R73713 VSS.n8817 VSS.n1367 0.0140606
R73714 VSS.n1380 VSS.n1372 0.0140606
R73715 VSS.n1381 VSS.n1380 0.0140606
R73716 VSS.n8811 VSS.n1370 0.0140606
R73717 VSS.n1461 VSS.n1452 0.0140606
R73718 VSS.n1472 VSS.n1454 0.0140606
R73719 VSS.n8695 VSS.n1450 0.0140606
R73720 VSS.n8695 VSS.n8694 0.0140606
R73721 VSS.n8697 VSS.n1449 0.0140606
R73722 VSS.n8697 VSS.n8696 0.0140606
R73723 VSS.n8699 VSS.n1448 0.0140606
R73724 VSS.n8699 VSS.n8698 0.0140606
R73725 VSS.n8701 VSS.n1447 0.0140606
R73726 VSS.n8701 VSS.n8700 0.0140606
R73727 VSS.n8702 VSS.n1445 0.0140606
R73728 VSS.n1468 VSS.n1456 0.0140606
R73729 VSS.n8704 VSS.n1468 0.0140606
R73730 VSS.n1467 VSS.n1457 0.0140606
R73731 VSS.n8706 VSS.n1467 0.0140606
R73732 VSS.n1466 VSS.n1458 0.0140606
R73733 VSS.n8708 VSS.n1466 0.0140606
R73734 VSS.n1465 VSS.n1459 0.0140606
R73735 VSS.n995 VSS.n983 0.0140606
R73736 VSS.n9081 VSS.n9079 0.0140606
R73737 VSS.n9079 VSS.n984 0.0140606
R73738 VSS.n9084 VSS.n9082 0.0140606
R73739 VSS.n9082 VSS.n985 0.0140606
R73740 VSS.n9087 VSS.n9085 0.0140606
R73741 VSS.n9085 VSS.n986 0.0140606
R73742 VSS.n9090 VSS.n9088 0.0140606
R73743 VSS.n9088 VSS.n987 0.0140606
R73744 VSS.n9093 VSS.n9091 0.0140606
R73745 VSS.n9091 VSS.n988 0.0140606
R73746 VSS.n9096 VSS.n9094 0.0140606
R73747 VSS.n9094 VSS.n989 0.0140606
R73748 VSS.n9099 VSS.n9097 0.0140606
R73749 VSS.n9097 VSS.n990 0.0140606
R73750 VSS.n9102 VSS.n9100 0.0140606
R73751 VSS.n9100 VSS.n991 0.0140606
R73752 VSS.n9105 VSS.n9103 0.0140606
R73753 VSS.n9103 VSS.n992 0.0140606
R73754 VSS.n9108 VSS.n9106 0.0140606
R73755 VSS.n9106 VSS.n993 0.0140606
R73756 VSS.n9112 VSS.n9111 0.0140606
R73757 VSS.n9113 VSS.n9112 0.0140606
R73758 VSS.n9240 VSS.n874 0.0140606
R73759 VSS.n897 VSS.n875 0.0140606
R73760 VSS.n9241 VSS.n897 0.0140606
R73761 VSS.n896 VSS.n876 0.0140606
R73762 VSS.n9242 VSS.n896 0.0140606
R73763 VSS.n895 VSS.n877 0.0140606
R73764 VSS.n9243 VSS.n895 0.0140606
R73765 VSS.n894 VSS.n878 0.0140606
R73766 VSS.n9244 VSS.n894 0.0140606
R73767 VSS.n893 VSS.n879 0.0140606
R73768 VSS.n9245 VSS.n893 0.0140606
R73769 VSS.n892 VSS.n880 0.0140606
R73770 VSS.n9246 VSS.n892 0.0140606
R73771 VSS.n891 VSS.n881 0.0140606
R73772 VSS.n9247 VSS.n891 0.0140606
R73773 VSS.n890 VSS.n882 0.0140606
R73774 VSS.n9248 VSS.n890 0.0140606
R73775 VSS.n889 VSS.n883 0.0140606
R73776 VSS.n9251 VSS.n889 0.0140606
R73777 VSS.n888 VSS.n884 0.0140606
R73778 VSS.n888 VSS.n886 0.0140606
R73779 VSS.n9255 VSS.n885 0.0140606
R73780 VSS.n9249 VSS.n885 0.0140606
R73781 VSS.n4436 VSS.n4433 0.0140606
R73782 VSS.n4435 VSS.n4427 0.0140606
R73783 VSS.n4503 VSS.n4502 0.0140606
R73784 VSS.n5654 VSS.n4268 0.0140606
R73785 VSS.n4023 VSS.n4017 0.0140606
R73786 VSS.n6081 VSS.n6080 0.0140606
R73787 VSS.n6078 VSS.n6037 0.0140606
R73788 VSS.n6077 VSS.n4072 0.0140606
R73789 VSS.n6036 VSS.n5900 0.0140606
R73790 VSS.n6307 VSS.n6306 0.0140606
R73791 VSS.n6304 VSS.n3799 0.0140606
R73792 VSS.n6303 VSS.n3718 0.0140606
R73793 VSS.n3798 VSS.n3719 0.0140606
R73794 VSS.n6608 VSS.n3164 0.0140606
R73795 VSS.n6607 VSS.n6606 0.0140606
R73796 VSS.n6604 VSS.n3196 0.0140606
R73797 VSS.n6603 VSS.n3193 0.0140606
R73798 VSS.n3195 VSS.n3194 0.0140606
R73799 VSS.n5885 VSS.n5735 0.0140606
R73800 VSS.n5890 VSS.n5739 0.0140606
R73801 VSS.n5889 VSS.n5736 0.0140606
R73802 VSS.n5738 VSS.n5737 0.0140606
R73803 VSS.n6999 VSS.n6998 0.0140606
R73804 VSS.n6996 VSS.n2740 0.0140606
R73805 VSS.n6995 VSS.n2656 0.0140606
R73806 VSS.n2739 VSS.n2657 0.0140606
R73807 VSS.n1626 VSS.n1624 0.0140606
R73808 VSS.n1636 VSS.n1624 0.0140606
R73809 VSS.n1628 VSS.n1623 0.0140606
R73810 VSS.n1635 VSS.n1623 0.0140606
R73811 VSS.n1631 VSS.n1621 0.0140606
R73812 VSS.n8536 VSS.n1621 0.0140606
R73813 VSS.n1633 VSS.n1620 0.0140606
R73814 VSS.n1620 VSS.n1618 0.0140606
R73815 VSS.n1494 VSS.n1486 0.0140606
R73816 VSS.n1506 VSS.n1505 0.0140606
R73817 VSS.n1506 VSS.n1483 0.0140606
R73818 VSS.n8668 VSS.n1504 0.0140606
R73819 VSS.n1504 VSS.n1482 0.0140606
R73820 VSS.n8670 VSS.n1503 0.0140606
R73821 VSS.n1503 VSS.n1481 0.0140606
R73822 VSS.n8672 VSS.n1502 0.0140606
R73823 VSS.n1502 VSS.n1480 0.0140606
R73824 VSS.n8674 VSS.n1479 0.0140606
R73825 VSS.n8677 VSS.n8676 0.0140606
R73826 VSS.n8677 VSS.n1489 0.0140606
R73827 VSS.n8679 VSS.n8678 0.0140606
R73828 VSS.n8679 VSS.n1490 0.0140606
R73829 VSS.n8681 VSS.n8680 0.0140606
R73830 VSS.n8681 VSS.n1491 0.0140606
R73831 VSS.n8683 VSS.n8682 0.0140606
R73832 VSS.n8683 VSS.n1492 0.0140606
R73833 VSS.n2444 VSS.n2429 0.0140606
R73834 VSS.n2443 VSS.n2428 0.0140606
R73835 VSS.n9121 VSS.n962 0.0140606
R73836 VSS.n9122 VSS.n9121 0.0140606
R73837 VSS.n9124 VSS.n963 0.0140606
R73838 VSS.n9125 VSS.n9124 0.0140606
R73839 VSS.n9127 VSS.n964 0.0140606
R73840 VSS.n9128 VSS.n9127 0.0140606
R73841 VSS.n9130 VSS.n965 0.0140606
R73842 VSS.n9131 VSS.n9130 0.0140606
R73843 VSS.n9133 VSS.n966 0.0140606
R73844 VSS.n9134 VSS.n9133 0.0140606
R73845 VSS.n9136 VSS.n967 0.0140606
R73846 VSS.n9137 VSS.n9136 0.0140606
R73847 VSS.n9139 VSS.n968 0.0140606
R73848 VSS.n9140 VSS.n9139 0.0140606
R73849 VSS.n9142 VSS.n969 0.0140606
R73850 VSS.n9143 VSS.n9142 0.0140606
R73851 VSS.n9145 VSS.n970 0.0140606
R73852 VSS.n9146 VSS.n9145 0.0140606
R73853 VSS.n9148 VSS.n971 0.0140606
R73854 VSS.n9149 VSS.n9148 0.0140606
R73855 VSS.n9151 VSS.n972 0.0140606
R73856 VSS.n9152 VSS.n9151 0.0140606
R73857 VSS.n9154 VSS.n973 0.0140606
R73858 VSS.n9208 VSS.n9198 0.0140606
R73859 VSS.n9198 VSS.n903 0.0140606
R73860 VSS.n9209 VSS.n9199 0.0140606
R73861 VSS.n9199 VSS.n904 0.0140606
R73862 VSS.n9210 VSS.n9200 0.0140606
R73863 VSS.n9200 VSS.n905 0.0140606
R73864 VSS.n9211 VSS.n9201 0.0140606
R73865 VSS.n9201 VSS.n906 0.0140606
R73866 VSS.n9212 VSS.n9202 0.0140606
R73867 VSS.n9202 VSS.n907 0.0140606
R73868 VSS.n9213 VSS.n9203 0.0140606
R73869 VSS.n9203 VSS.n908 0.0140606
R73870 VSS.n9214 VSS.n9204 0.0140606
R73871 VSS.n9204 VSS.n909 0.0140606
R73872 VSS.n9215 VSS.n9205 0.0140606
R73873 VSS.n9205 VSS.n910 0.0140606
R73874 VSS.n9216 VSS.n9206 0.0140606
R73875 VSS.n9206 VSS.n911 0.0140606
R73876 VSS.n9217 VSS.n9207 0.0140606
R73877 VSS.n9207 VSS.n912 0.0140606
R73878 VSS.n9220 VSS.n9219 0.0140606
R73879 VSS.n9220 VSS.n913 0.0140606
R73880 VSS.n9222 VSS.n914 0.0140606
R73881 VSS.n2352 VSS.n2351 0.0140606
R73882 VSS.n2355 VSS.n2354 0.0140606
R73883 VSS.n2353 VSS.n2349 0.0140606
R73884 VSS.n4502 VSS.n4497 0.0140606
R73885 VSS.n5655 VSS.n5654 0.0140606
R73886 VSS.n4024 VSS.n4023 0.0140606
R73887 VSS.n6610 VSS.n3164 0.0140606
R73888 VSS.n1627 VSS.n1626 0.0140606
R73889 VSS.n1636 VSS.n1629 0.0140606
R73890 VSS.n1629 VSS.n1628 0.0140606
R73891 VSS.n1635 VSS.n1630 0.0140606
R73892 VSS.n1632 VSS.n1631 0.0140606
R73893 VSS.n8537 VSS.n8536 0.0140606
R73894 VSS.n8537 VSS.n1633 0.0140606
R73895 VSS.n8539 VSS.n1618 0.0140606
R73896 VSS.n1494 VSS.n1485 0.0140606
R73897 VSS.n1505 VSS.n1487 0.0140606
R73898 VSS.n8669 VSS.n1483 0.0140606
R73899 VSS.n8669 VSS.n8668 0.0140606
R73900 VSS.n8671 VSS.n1482 0.0140606
R73901 VSS.n8671 VSS.n8670 0.0140606
R73902 VSS.n8673 VSS.n1481 0.0140606
R73903 VSS.n8673 VSS.n8672 0.0140606
R73904 VSS.n8675 VSS.n1480 0.0140606
R73905 VSS.n8675 VSS.n8674 0.0140606
R73906 VSS.n8676 VSS.n1478 0.0140606
R73907 VSS.n1501 VSS.n1489 0.0140606
R73908 VSS.n8678 VSS.n1501 0.0140606
R73909 VSS.n1500 VSS.n1490 0.0140606
R73910 VSS.n8680 VSS.n1500 0.0140606
R73911 VSS.n1499 VSS.n1491 0.0140606
R73912 VSS.n8682 VSS.n1499 0.0140606
R73913 VSS.n1498 VSS.n1492 0.0140606
R73914 VSS.n974 VSS.n962 0.0140606
R73915 VSS.n9122 VSS.n9120 0.0140606
R73916 VSS.n9120 VSS.n963 0.0140606
R73917 VSS.n9125 VSS.n9123 0.0140606
R73918 VSS.n9123 VSS.n964 0.0140606
R73919 VSS.n9128 VSS.n9126 0.0140606
R73920 VSS.n9126 VSS.n965 0.0140606
R73921 VSS.n9131 VSS.n9129 0.0140606
R73922 VSS.n9129 VSS.n966 0.0140606
R73923 VSS.n9134 VSS.n9132 0.0140606
R73924 VSS.n9132 VSS.n967 0.0140606
R73925 VSS.n9137 VSS.n9135 0.0140606
R73926 VSS.n9135 VSS.n968 0.0140606
R73927 VSS.n9140 VSS.n9138 0.0140606
R73928 VSS.n9138 VSS.n969 0.0140606
R73929 VSS.n9143 VSS.n9141 0.0140606
R73930 VSS.n9141 VSS.n970 0.0140606
R73931 VSS.n9146 VSS.n9144 0.0140606
R73932 VSS.n9144 VSS.n971 0.0140606
R73933 VSS.n9149 VSS.n9147 0.0140606
R73934 VSS.n9147 VSS.n972 0.0140606
R73935 VSS.n9153 VSS.n9152 0.0140606
R73936 VSS.n9154 VSS.n9153 0.0140606
R73937 VSS.n9208 VSS.n902 0.0140606
R73938 VSS.n927 VSS.n903 0.0140606
R73939 VSS.n9209 VSS.n927 0.0140606
R73940 VSS.n926 VSS.n904 0.0140606
R73941 VSS.n9210 VSS.n926 0.0140606
R73942 VSS.n925 VSS.n905 0.0140606
R73943 VSS.n9211 VSS.n925 0.0140606
R73944 VSS.n924 VSS.n906 0.0140606
R73945 VSS.n9212 VSS.n924 0.0140606
R73946 VSS.n923 VSS.n907 0.0140606
R73947 VSS.n9213 VSS.n923 0.0140606
R73948 VSS.n922 VSS.n908 0.0140606
R73949 VSS.n9214 VSS.n922 0.0140606
R73950 VSS.n921 VSS.n909 0.0140606
R73951 VSS.n9215 VSS.n921 0.0140606
R73952 VSS.n920 VSS.n910 0.0140606
R73953 VSS.n9216 VSS.n920 0.0140606
R73954 VSS.n919 VSS.n911 0.0140606
R73955 VSS.n9217 VSS.n919 0.0140606
R73956 VSS.n918 VSS.n912 0.0140606
R73957 VSS.n9219 VSS.n918 0.0140606
R73958 VSS.n917 VSS.n913 0.0140606
R73959 VSS.n917 VSS.n914 0.0140606
R73960 VSS.n4435 VSS.n4430 0.0140606
R73961 VSS.n4436 VSS.n4424 0.0140606
R73962 VSS.n5167 VSS.n4451 0.0140606
R73963 VSS.n5170 VSS.n5169 0.0140606
R73964 VSS.n5900 VSS.n4072 0.0140606
R73965 VSS.n5909 VSS.n5902 0.0140606
R73966 VSS.n6078 VSS.n6077 0.0140606
R73967 VSS.n5956 VSS.n5955 0.0140606
R73968 VSS.n6037 VSS.n4070 0.0140606
R73969 VSS.n6080 VSS.n4070 0.0140606
R73970 VSS.n5954 VSS.n5953 0.0140606
R73971 VSS.n5953 VSS.n5908 0.0140606
R73972 VSS.n3719 VSS.n3718 0.0140606
R73973 VSS.n3708 VSS.n3707 0.0140606
R73974 VSS.n6304 VSS.n6303 0.0140606
R73975 VSS.n6316 VSS.n6315 0.0140606
R73976 VSS.n3799 VSS.n3716 0.0140606
R73977 VSS.n6306 VSS.n3716 0.0140606
R73978 VSS.n6313 VSS.n3710 0.0140606
R73979 VSS.n6313 VSS.n3706 0.0140606
R73980 VSS.n3194 VSS.n3193 0.0140606
R73981 VSS.n3130 VSS.n3129 0.0140606
R73982 VSS.n6604 VSS.n6603 0.0140606
R73983 VSS.n6622 VSS.n6621 0.0140606
R73984 VSS.n3196 VSS.n3191 0.0140606
R73985 VSS.n6606 VSS.n3191 0.0140606
R73986 VSS.n6619 VSS.n3132 0.0140606
R73987 VSS.n6619 VSS.n3128 0.0140606
R73988 VSS.n5737 VSS.n5736 0.0140606
R73989 VSS.n2962 VSS.n2958 0.0140606
R73990 VSS.n5890 VSS.n5889 0.0140606
R73991 VSS.n6764 VSS.n6763 0.0140606
R73992 VSS.n5887 VSS.n5739 0.0140606
R73993 VSS.n5887 VSS.n5735 0.0140606
R73994 VSS.n6762 VSS.n6761 0.0140606
R73995 VSS.n6761 VSS.n2961 0.0140606
R73996 VSS.n2657 VSS.n2656 0.0140606
R73997 VSS.n2646 VSS.n2645 0.0140606
R73998 VSS.n6996 VSS.n6995 0.0140606
R73999 VSS.n7008 VSS.n7007 0.0140606
R74000 VSS.n2740 VSS.n2654 0.0140606
R74001 VSS.n6998 VSS.n2654 0.0140606
R74002 VSS.n7005 VSS.n2648 0.0140606
R74003 VSS.n7005 VSS.n2644 0.0140606
R74004 VSS.n2354 VSS.n2353 0.0140606
R74005 VSS.n9448 VSS.n9447 0.0140606
R74006 VSS.n2355 VSS.n2352 0.0140606
R74007 VSS.n768 VSS.n765 0.0140606
R74008 VSS.n2351 VSS.n915 0.0140606
R74009 VSS.n9450 VSS.n767 0.0140606
R74010 VSS.n2444 VSS.n2443 0.0140606
R74011 VSS.n2463 VSS.n2448 0.0140606
R74012 VSS.n2429 VSS.n1496 0.0140606
R74013 VSS.n2464 VSS.n1463 0.0140606
R74014 VSS.n7194 VSS.n7193 0.0138885
R74015 VSS.n7200 VSS.n7199 0.0138885
R74016 VSS.n7212 VSS.n7210 0.0138885
R74017 VSS.n7214 VSS.n2535 0.0138885
R74018 VSS.n7219 VSS.n7218 0.0138885
R74019 VSS.n7211 VSS.n2535 0.0138885
R74020 VSS.n7212 VSS.n7211 0.0138885
R74021 VSS.n7218 VSS.n7217 0.0138885
R74022 VSS.n7238 VSS.n7237 0.0138885
R74023 VSS.n7235 VSS.n2512 0.0138885
R74024 VSS.n7080 VSS.n2519 0.0138885
R74025 VSS.n7092 VSS.n7091 0.0138885
R74026 VSS.n7081 VSS.n7080 0.0138885
R74027 VSS.n7091 VSS.n7085 0.0138885
R74028 VSS.n2489 VSS.n2484 0.0138885
R74029 VSS.n7177 VSS.n2487 0.0138885
R74030 VSS.n7173 VSS.n2541 0.0138885
R74031 VSS.n7164 VSS.n2547 0.0138885
R74032 VSS.n2543 VSS.n2541 0.0138885
R74033 VSS.n7169 VSS.n2547 0.0138885
R74034 VSS.n7237 VSS.n2508 0.0138885
R74035 VSS.n7193 VSS.n7192 0.0138885
R74036 VSS.n7255 VSS.n2484 0.0138885
R74037 VSS.n8553 VSS.n1589 0.0138885
R74038 VSS.n8552 VSS.n1594 0.0138885
R74039 VSS.n8551 VSS.n1588 0.0138885
R74040 VSS.n1600 VSS.n1597 0.0138885
R74041 VSS.n8545 VSS.n1605 0.0138885
R74042 VSS.n1613 VSS.n1387 0.0138885
R74043 VSS.n1390 VSS.n1344 0.0138885
R74044 VSS.n8833 VSS.n1350 0.0138885
R74045 VSS.n1592 VSS.n1589 0.0138885
R74046 VSS.n1594 VSS.n1588 0.0138885
R74047 VSS.n8550 VSS.n1597 0.0138885
R74048 VSS.n1610 VSS.n1387 0.0138885
R74049 VSS.n8808 VSS.n1344 0.0138885
R74050 VSS.n8838 VSS.n1350 0.0138885
R74051 VSS.n8553 VSS.n8552 0.0138885
R74052 VSS.n8073 VSS.n8002 0.0138885
R74053 VSS.n8007 VSS.n8002 0.0138885
R74054 VSS.n8013 VSS.n8012 0.0138885
R74055 VSS.n8015 VSS.n8013 0.0138885
R74056 VSS.n8065 VSS.n8019 0.0138885
R74057 VSS.n8057 VSS.n8023 0.0138885
R74058 VSS.n8028 VSS.n8027 0.0138885
R74059 VSS.n8030 VSS.n8028 0.0138885
R74060 VSS.n8035 VSS.n8034 0.0138885
R74061 VSS.n8038 VSS.n8035 0.0138885
R74062 VSS.n8074 VSS.n8073 0.0138885
R74063 VSS.n8070 VSS.n8012 0.0138885
R74064 VSS.n8024 VSS.n8023 0.0138885
R74065 VSS.n8051 VSS.n8027 0.0138885
R74066 VSS.n8046 VSS.n8034 0.0138885
R74067 VSS.n8044 VSS.n8038 0.0138885
R74068 VSS.n8049 VSS.n8030 0.0138885
R74069 VSS.n8068 VSS.n8015 0.0138885
R74070 VSS.n8007 VSS.n8004 0.0138885
R74071 VSS.n1566 VSS.n1560 0.0138885
R74072 VSS.n8562 VSS.n1562 0.0138885
R74073 VSS.n1564 VSS.n1562 0.0138885
R74074 VSS.n8389 VSS.n8386 0.0138885
R74075 VSS.n8387 VSS.n8385 0.0138885
R74076 VSS.n8393 VSS.n8387 0.0138885
R74077 VSS.n8400 VSS.n8398 0.0138885
R74078 VSS.n8399 VSS.n1362 0.0138885
R74079 VSS.n8820 VSS.n8818 0.0138885
R74080 VSS.n8819 VSS.n1321 0.0138885
R74081 VSS.n8846 VSS.n8845 0.0138885
R74082 VSS.n1319 VSS.n1317 0.0138885
R74083 VSS.n1317 VSS.n1314 0.0138885
R74084 VSS.n8855 VSS.n8852 0.0138885
R74085 VSS.n8853 VSS.n1311 0.0138885
R74086 VSS.n8850 VSS.n1311 0.0138885
R74087 VSS.n8565 VSS.n1560 0.0138885
R74088 VSS.n8563 VSS.n8562 0.0138885
R74089 VSS.n8391 VSS.n8386 0.0138885
R74090 VSS.n8390 VSS.n8385 0.0138885
R74091 VSS.n8818 VSS.n1364 0.0138885
R74092 VSS.n8847 VSS.n8846 0.0138885
R74093 VSS.n1320 VSS.n1319 0.0138885
R74094 VSS.n8856 VSS.n8855 0.0138885
R74095 VSS.n8853 VSS.n1313 0.0138885
R74096 VSS.n8850 VSS.n1312 0.0138885
R74097 VSS.n8849 VSS.n1314 0.0138885
R74098 VSS.n8820 VSS.n8819 0.0138885
R74099 VSS.n8403 VSS.n8393 0.0138885
R74100 VSS.n1565 VSS.n1564 0.0138885
R74101 VSS.n8398 VSS.n8395 0.0138885
R74102 VSS.n8400 VSS.n8399 0.0138885
R74103 VSS.n1607 VSS.n1605 0.0138885
R74104 VSS.n8020 VSS.n8019 0.0138885
R74105 VSS.n2515 VSS.n2512 0.0138885
R74106 VSS.n7201 VSS.n7200 0.0138885
R74107 VSS.n7178 VSS.n7177 0.0138885
R74108 VSS.n7196 VSS.n7195 0.0138885
R74109 VSS.n7202 VSS.n7201 0.0138885
R74110 VSS.n7215 VSS.n7214 0.0138885
R74111 VSS.n7221 VSS.n7220 0.0138885
R74112 VSS.n7216 VSS.n7215 0.0138885
R74113 VSS.n7221 VSS.n2527 0.0138885
R74114 VSS.n7239 VSS.n2509 0.0138885
R74115 VSS.n2516 VSS.n2515 0.0138885
R74116 VSS.n7082 VSS.n7081 0.0138885
R74117 VSS.n7093 VSS.n7086 0.0138885
R74118 VSS.n7082 VSS.n7060 0.0138885
R74119 VSS.n7087 VSS.n7086 0.0138885
R74120 VSS.n7256 VSS.n2485 0.0138885
R74121 VSS.n7178 VSS.n2539 0.0138885
R74122 VSS.n2544 VSS.n2543 0.0138885
R74123 VSS.n7165 VSS.n2550 0.0138885
R74124 VSS.n2545 VSS.n2544 0.0138885
R74125 VSS.n2551 VSS.n2550 0.0138885
R74126 VSS.n7256 VSS.n2486 0.0138885
R74127 VSS.n7196 VSS.n7186 0.0138885
R74128 VSS.n2510 VSS.n2509 0.0138885
R74129 VSS.n8546 VSS.n1599 0.0138885
R74130 VSS.n8543 VSS.n8542 0.0138885
R74131 VSS.n8809 VSS.n1388 0.0138885
R74132 VSS.n8839 VSS.n1347 0.0138885
R74133 VSS.n8832 VSS.n8831 0.0138885
R74134 VSS.n8835 VSS.n8832 0.0138885
R74135 VSS.n1347 VSS.n1346 0.0138885
R74136 VSS.n1609 VSS.n1388 0.0138885
R74137 VSS.n1601 VSS.n1599 0.0138885
R74138 VSS.n8071 VSS.n8003 0.0138885
R74139 VSS.n8066 VSS.n8014 0.0138885
R74140 VSS.n8063 VSS.n8062 0.0138885
R74141 VSS.n8055 VSS.n8054 0.0138885
R74142 VSS.n8047 VSS.n8029 0.0138885
R74143 VSS.n8042 VSS.n8037 0.0138885
R74144 VSS.n8039 VSS.n8037 0.0138885
R74145 VSS.n8031 VSS.n8029 0.0138885
R74146 VSS.n8055 VSS.n8025 0.0138885
R74147 VSS.n8016 VSS.n8014 0.0138885
R74148 VSS.n8009 VSS.n8003 0.0138885
R74149 VSS.n8543 VSS.n1608 0.0138885
R74150 VSS.n8063 VSS.n8021 0.0138885
R74151 VSS.n2540 VSS.n2539 0.0138885
R74152 VSS.n7202 VSS.n2537 0.0138885
R74153 VSS.n2517 VSS.n2516 0.0138885
R74154 VSS.n4859 VSS.n4857 0.0138099
R74155 VSS.n3733 VSS.n3154 0.0138099
R74156 VSS.n6778 VSS.n2947 0.0138099
R74157 VSS.n4860 VSS.n4500 0.0138099
R74158 VSS.n3773 VSS.n3184 0.0138099
R74159 VSS.n6779 VSS.n2929 0.0138099
R74160 VSS.n8964 VSS.n1096 0.0137874
R74161 VSS.n8963 VSS.n1093 0.0137874
R74162 VSS.n2297 VSS.n2159 0.0137874
R74163 VSS.n1428 VSS.n1396 0.0137874
R74164 VSS.n8804 VSS.n1429 0.0137874
R74165 VSS.n1544 VSS.n1540 0.0137874
R74166 VSS.n8634 VSS.n1542 0.0137874
R74167 VSS.n8090 VSS.n2086 0.0137874
R74168 VSS.n8089 VSS.n2083 0.0137874
R74169 VSS.n1199 VSS.n747 0.0137874
R74170 VSS.n221 VSS.n217 0.0134331
R74171 VSS.n9764 VSS.n224 0.0134331
R74172 VSS.n225 VSS.n220 0.0134331
R74173 VSS.n9760 VSS.n9759 0.0134331
R74174 VSS.n2325 VSS.n2144 0.0134331
R74175 VSS.n2401 VSS.n1856 0.0134331
R74176 VSS.n4746 VSS.n4554 0.0134331
R74177 VSS.n4754 VSS.n4560 0.0134331
R74178 VSS.n4748 VSS.n4553 0.0134331
R74179 VSS.n4785 VSS.n4561 0.0134331
R74180 VSS.n9692 VSS.n254 0.0134331
R74181 VSS.n9690 VSS.n253 0.0134331
R74182 VSS.n9689 VSS.n252 0.0134331
R74183 VSS.n274 VSS.n251 0.0134331
R74184 VSS.n4517 VSS.n4513 0.0134331
R74185 VSS.n5077 VSS.n4520 0.0134331
R74186 VSS.n4521 VSS.n4516 0.0134331
R74187 VSS.n5073 VSS.n5072 0.0134331
R74188 VSS.n4327 VSS.n4323 0.0134331
R74189 VSS.n5250 VSS.n4329 0.0134331
R74190 VSS.n5246 VSS.n4326 0.0134331
R74191 VSS.n5247 VSS.n4320 0.0134331
R74192 VSS.n4758 VSS.n4585 0.0134331
R74193 VSS.n3860 VSS.n3856 0.0134331
R74194 VSS.n9810 VSS.n171 0.0134331
R74195 VSS.n5467 VSS.n5435 0.0134331
R74196 VSS.n9774 VSS.n196 0.0134331
R74197 VSS.n9772 VSS.n201 0.0134331
R74198 VSS.n9771 VSS.n195 0.0134331
R74199 VSS.n9777 VSS.n202 0.0134331
R74200 VSS.n1171 VSS.n731 0.0134331
R74201 VSS.n9401 VSS.n702 0.0134331
R74202 VSS.n4859 VSS.n4852 0.0133873
R74203 VSS.n3733 VSS.n3144 0.0133873
R74204 VSS.n6778 VSS.n2950 0.0133873
R74205 VSS.n4860 VSS.n4498 0.0133873
R74206 VSS.n3773 VSS.n3174 0.0133873
R74207 VSS.n6779 VSS.n2932 0.0133873
R74208 VSS.n161 VSS.n75 0.0130787
R74209 VSS.n4132 VSS.n348 0.0130787
R74210 VSS.n4163 VSS.n355 0.0130787
R74211 VSS.n4134 VSS.n347 0.0130787
R74212 VSS.n4138 VSS.n356 0.0130787
R74213 VSS.n357 VSS.n346 0.0130787
R74214 VSS.n2281 VSS.n2153 0.0130787
R74215 VSS.n2383 VSS.n1841 0.0130787
R74216 VSS.n4672 VSS.n4624 0.0130787
R74217 VSS.n9894 VSS.n9893 0.0130787
R74218 VSS.n4124 VSS.n314 0.0130787
R74219 VSS.n4167 VSS.n322 0.0130787
R74220 VSS.n4126 VSS.n313 0.0130787
R74221 VSS.n4130 VSS.n323 0.0130787
R74222 VSS.n324 VSS.n312 0.0130787
R74223 VSS.n4664 VSS.n4387 0.0130787
R74224 VSS.n4080 VSS.n3983 0.0130787
R74225 VSS.n4109 VSS.n3993 0.0130787
R74226 VSS.n4082 VSS.n3982 0.0130787
R74227 VSS.n4105 VSS.n3994 0.0130787
R74228 VSS.n3995 VSS.n3981 0.0130787
R74229 VSS.n4668 VSS.n4347 0.0130787
R74230 VSS.n4084 VSS.n3941 0.0130787
R74231 VSS.n4101 VSS.n3948 0.0130787
R74232 VSS.n4086 VSS.n3940 0.0130787
R74233 VSS.n4097 VSS.n3949 0.0130787
R74234 VSS.n3950 VSS.n3939 0.0130787
R74235 VSS.n4638 VSS.n4596 0.0130787
R74236 VSS.n3852 VSS.n3838 0.0130787
R74237 VSS.n9817 VSS.n137 0.0130787
R74238 VSS.n4150 VSS.n409 0.0130787
R74239 VSS.n165 VSS.n106 0.0130787
R74240 VSS.n4140 VSS.n384 0.0130787
R74241 VSS.n4160 VSS.n394 0.0130787
R74242 VSS.n4142 VSS.n383 0.0130787
R74243 VSS.n4146 VSS.n395 0.0130787
R74244 VSS.n396 VSS.n382 0.0130787
R74245 VSS.n1215 VSS.n740 0.0130787
R74246 VSS.n9419 VSS.n688 0.0130787
R74247 VSS.n3725 VSS.n3147 0.0129648
R74248 VSS.n6804 VSS.n6803 0.0129648
R74249 VSS.n3789 VSS.n3177 0.0129648
R74250 VSS.n6801 VSS.n2935 0.0129648
R74251 VSS.n2366 VSS.n2335 0.0128916
R74252 VSS.n2361 VSS.n2342 0.0128916
R74253 VSS.n9446 VSS.n769 0.0128916
R74254 VSS.n9441 VSS.n777 0.0128916
R74255 VSS.n2338 VSS.n2335 0.0128916
R74256 VSS.n2345 VSS.n2342 0.0128916
R74257 VSS.n773 VSS.n769 0.0128916
R74258 VSS.n9370 VSS.n777 0.0128916
R74259 VSS.n2088 VSS.n2082 0.0128916
R74260 VSS.n8093 VSS.n8092 0.0128916
R74261 VSS.n8094 VSS.n8093 0.0128916
R74262 VSS.n2433 VSS.n2084 0.0128916
R74263 VSS.n2437 VSS.n2435 0.0128916
R74264 VSS.n2438 VSS.n2437 0.0128916
R74265 VSS.n2441 VSS.n2440 0.0128916
R74266 VSS.n2442 VSS.n2427 0.0128916
R74267 VSS.n2465 VSS.n2447 0.0128916
R74268 VSS.n2450 VSS.n2449 0.0128916
R74269 VSS.n2461 VSS.n2451 0.0128916
R74270 VSS.n2456 VSS.n2455 0.0128916
R74271 VSS.n2457 VSS.n2456 0.0128916
R74272 VSS.n1098 VSS.n1092 0.0128916
R74273 VSS.n8967 VSS.n8966 0.0128916
R74274 VSS.n8968 VSS.n8967 0.0128916
R74275 VSS.n8091 VSS.n2082 0.0128916
R74276 VSS.n2434 VSS.n2433 0.0128916
R74277 VSS.n2453 VSS.n2451 0.0128916
R74278 VSS.n8965 VSS.n1092 0.0128916
R74279 VSS.n8092 VSS.n8091 0.0128916
R74280 VSS.n2435 VSS.n2434 0.0128916
R74281 VSS.n2445 VSS.n2427 0.0128916
R74282 VSS.n2462 VSS.n2450 0.0128916
R74283 VSS.n2455 VSS.n2453 0.0128916
R74284 VSS.n8966 VSS.n8965 0.0128916
R74285 VSS.n8095 VSS.n8094 0.0128916
R74286 VSS.n2439 VSS.n2438 0.0128916
R74287 VSS.n2442 VSS.n2441 0.0128916
R74288 VSS.n2449 VSS.n2447 0.0128916
R74289 VSS.n2458 VSS.n2457 0.0128916
R74290 VSS.n8969 VSS.n8968 0.0128916
R74291 VSS.n9863 VSS.n83 0.0127244
R74292 VSS.n2279 VSS.n2154 0.0127244
R74293 VSS.n2385 VSS.n1842 0.0127244
R74294 VSS.n4704 VSS.n4675 0.0127244
R74295 VSS.n25 VSS.n20 0.0127244
R74296 VSS.n5205 VSS.n4395 0.0127244
R74297 VSS.n5232 VSS.n4355 0.0127244
R74298 VSS.n4719 VSS.n4604 0.0127244
R74299 VSS.n6261 VSS.n3837 0.0127244
R74300 VSS.n9833 VSS.n9821 0.0127244
R74301 VSS.n4149 VSS.n408 0.0127244
R74302 VSS.n9848 VSS.n114 0.0127244
R74303 VSS.n1217 VSS.n741 0.0127244
R74304 VSS.n9417 VSS.n689 0.0127244
R74305 VSS.n4922 VSS.n4254 0.0125423
R74306 VSS.n4920 VSS.n4252 0.0125423
R74307 VSS.n4919 VSS.n4255 0.0125423
R74308 VSS.n4915 VSS.n4251 0.0125423
R74309 VSS.n4918 VSS.n4257 0.0125423
R74310 VSS.n5717 VSS.n4174 0.0125423
R74311 VSS.n3741 VSS.n3157 0.0125423
R74312 VSS.n4275 VSS.n4272 0.0125423
R74313 VSS.n5651 VSS.n4270 0.0125423
R74314 VSS.n4278 VSS.n4273 0.0125423
R74315 VSS.n5649 VSS.n4269 0.0125423
R74316 VSS.n5655 VSS.n5653 0.0125423
R74317 VSS.n5715 VSS.n4018 0.0125423
R74318 VSS.n3757 VSS.n3187 0.0125423
R74319 VSS.n2371 VSS.n2330 0.0124231
R74320 VSS.n9433 VSS.n9432 0.0124231
R74321 VSS.n2278 VSS.n2170 0.0124231
R74322 VSS.n1223 VSS.n1219 0.0124231
R74323 VSS.n2562 VSS.n2558 0.0123796
R74324 VSS.n7171 VSS.n2542 0.0123796
R74325 VSS.n7172 VSS.n2536 0.0123796
R74326 VSS.n7208 VSS.n2533 0.0123796
R74327 VSS.n7209 VSS.n7208 0.0123796
R74328 VSS.n7063 VSS.n7062 0.0123796
R74329 VSS.n7083 VSS.n7064 0.0123796
R74330 VSS.n7065 VSS.n2599 0.0123796
R74331 VSS.n2600 VSS.n1377 0.0123796
R74332 VSS.n8821 VSS.n1366 0.0123796
R74333 VSS.n1389 VSS.n1386 0.0123796
R74334 VSS.n1612 VSS.n1611 0.0123796
R74335 VSS.n8052 VSS.n8022 0.0123796
R74336 VSS.n7079 VSS.n7065 0.0123796
R74337 VSS.n7213 VSS.n2533 0.0123796
R74338 VSS.n7209 VSS.n2534 0.0123796
R74339 VSS.n7064 VSS.n7063 0.0123796
R74340 VSS.n7062 VSS.n7061 0.0123796
R74341 VSS.n7172 VSS.n7171 0.0123796
R74342 VSS.n2546 VSS.n2542 0.0123796
R74343 VSS.n2558 VSS.n2557 0.0123796
R74344 VSS.n8810 VSS.n1386 0.0123796
R74345 VSS.n1611 VSS.n1389 0.0123796
R74346 VSS.n8053 VSS.n8052 0.0123796
R74347 VSS.n1366 VSS.n1363 0.0123796
R74348 VSS.n7109 VSS.n2600 0.0123796
R74349 VSS.n7142 VSS.n7141 0.0123796
R74350 VSS.n7268 VSS.n2471 0.0123796
R74351 VSS.n7265 VSS.n2473 0.0123796
R74352 VSS.n7179 VSS.n7176 0.0123796
R74353 VSS.n7181 VSS.n2538 0.0123796
R74354 VSS.n7184 VSS.n7183 0.0123796
R74355 VSS.n7203 VSS.n7185 0.0123796
R74356 VSS.n7233 VSS.n2514 0.0123796
R74357 VSS.n7234 VSS.n2513 0.0123796
R74358 VSS.n7067 VSS.n2594 0.0123796
R74359 VSS.n7113 VSS.n2595 0.0123796
R74360 VSS.n8401 VSS.n8397 0.0123796
R74361 VSS.n8540 VSS.n1604 0.0123796
R74362 VSS.n8544 VSS.n1606 0.0123796
R74363 VSS.n8060 VSS.n8018 0.0123796
R74364 VSS.n7115 VSS.n2595 0.0123796
R74365 VSS.n8397 VSS.n8394 0.0123796
R74366 VSS.n8541 VSS.n8540 0.0123796
R74367 VSS.n1606 VSS.n1604 0.0123796
R74368 VSS.n8061 VSS.n8060 0.0123796
R74369 VSS.n7267 VSS.n2473 0.0123796
R74370 VSS.n7071 VSS.n7067 0.0123796
R74371 VSS.n7234 VSS.n7233 0.0123796
R74372 VSS.n2518 VSS.n2514 0.0123796
R74373 VSS.n7185 VSS.n7184 0.0123796
R74374 VSS.n7183 VSS.n7182 0.0123796
R74375 VSS.n7179 VSS.n2538 0.0123796
R74376 VSS.n7176 VSS.n2478 0.0123796
R74377 VSS.n7141 VSS.n2471 0.0123796
R74378 VSS.n7143 VSS.n7142 0.0123796
R74379 VSS.n7149 VSS.n7148 0.0123796
R74380 VSS.n7149 VSS.n2470 0.0123796
R74381 VSS.n5456 VSS.n5386 0.0123701
R74382 VSS.n5449 VSS.n5384 0.0123701
R74383 VSS.n5452 VSS.n5387 0.0123701
R74384 VSS.n5448 VSS.n5383 0.0123701
R74385 VSS.n2327 VSS.n2143 0.0123701
R74386 VSS.n2399 VSS.n1857 0.0123701
R74387 VSS.n9685 VSS.n280 0.0123701
R74388 VSS.n9684 VSS.n286 0.0123701
R74389 VSS.n298 VSS.n297 0.0123701
R74390 VSS.n294 VSS.n285 0.0123701
R74391 VSS.n5647 VSS.n4284 0.0123701
R74392 VSS.n4287 VSS.n4283 0.0123701
R74393 VSS.n5643 VSS.n4288 0.0123701
R74394 VSS.n5642 VSS.n4282 0.0123701
R74395 VSS.n5261 VSS.n4316 0.0123701
R74396 VSS.n5256 VSS.n4315 0.0123701
R74397 VSS.n5258 VSS.n4317 0.0123701
R74398 VSS.n5263 VSS.n4314 0.0123701
R74399 VSS.n4744 VSS.n4586 0.0123701
R74400 VSS.n6250 VSS.n3865 0.0123701
R74401 VSS.n181 VSS.n169 0.0123701
R74402 VSS.n5471 VSS.n5436 0.0123701
R74403 VSS.n5463 VSS.n5414 0.0123701
R74404 VSS.n5444 VSS.n5412 0.0123701
R74405 VSS.n5459 VSS.n5415 0.0123701
R74406 VSS.n5443 VSS.n5411 0.0123701
R74407 VSS.n1169 VSS.n730 0.0123701
R74408 VSS.n9403 VSS.n703 0.0123701
R74409 VSS.n5125 VSS.n4455 0.012331
R74410 VSS.n5123 VSS.n4431 0.012331
R74411 VSS.n4453 VSS.n4452 0.0121197
R74412 VSS.n4259 VSS.n4249 0.0121197
R74413 VSS.n6613 VSS.n3137 0.0121197
R74414 VSS.n4438 VSS.n4428 0.0121197
R74415 VSS.n4267 VSS.n4266 0.0121197
R74416 VSS.n6611 VSS.n6610 0.0121197
R74417 VSS.n2295 VSS.n2158 0.0120157
R74418 VSS.n8244 VSS.n1866 0.0120157
R74419 VSS.n1201 VSS.n746 0.0120157
R74420 VSS.n9525 VSS.n711 0.0120157
R74421 VSS.n84 VSS.n78 0.0119575
R74422 VSS.n88 VSS.n72 0.0119575
R74423 VSS.n80 VSS.n76 0.0119575
R74424 VSS.n87 VSS.n71 0.0119575
R74425 VSS.n81 VSS.n77 0.0119575
R74426 VSS.n86 VSS.n70 0.0119575
R74427 VSS.n9748 VSS.n232 0.0119575
R74428 VSS.n9752 VSS.n9750 0.0119575
R74429 VSS.n9751 VSS.n231 0.0119575
R74430 VSS.n9755 VSS.n9753 0.0119575
R74431 VSS.n9754 VSS.n230 0.0119575
R74432 VSS.n9757 VSS.n9756 0.0119575
R74433 VSS.n5391 VSS.n5382 0.0119575
R74434 VSS.n5395 VSS.n5394 0.0119575
R74435 VSS.n5390 VSS.n5381 0.0119575
R74436 VSS.n5524 VSS.n5523 0.0119575
R74437 VSS.n5389 VSS.n5380 0.0119575
R74438 VSS.n5526 VSS.n5388 0.0119575
R74439 VSS.n366 VSS.n350 0.0119575
R74440 VSS.n360 VSS.n353 0.0119575
R74441 VSS.n365 VSS.n349 0.0119575
R74442 VSS.n361 VSS.n354 0.0119575
R74443 VSS.n364 VSS.n348 0.0119575
R74444 VSS.n5943 VSS.n5942 0.0119575
R74445 VSS.n5940 VSS.n5919 0.0119575
R74446 VSS.n5923 VSS.n5917 0.0119575
R74447 VSS.n5939 VSS.n5938 0.0119575
R74448 VSS.n6329 VSS.n3693 0.0119575
R74449 VSS.n3694 VSS.n3692 0.0119575
R74450 VSS.n6325 VSS.n3689 0.0119575
R74451 VSS.n3691 VSS.n3690 0.0119575
R74452 VSS.n6425 VSS.n3600 0.0119575
R74453 VSS.n3626 VSS.n3598 0.0119575
R74454 VSS.n6414 VSS.n3601 0.0119575
R74455 VSS.n3621 VSS.n3597 0.0119575
R74456 VSS.n6415 VSS.n3602 0.0119575
R74457 VSS.n3620 VSS.n3596 0.0119575
R74458 VSS.n6416 VSS.n3603 0.0119575
R74459 VSS.n3619 VSS.n3595 0.0119575
R74460 VSS.n6417 VSS.n3604 0.0119575
R74461 VSS.n3618 VSS.n3594 0.0119575
R74462 VSS.n6418 VSS.n3605 0.0119575
R74463 VSS.n3617 VSS.n3593 0.0119575
R74464 VSS.n6419 VSS.n3606 0.0119575
R74465 VSS.n3616 VSS.n3592 0.0119575
R74466 VSS.n6420 VSS.n3607 0.0119575
R74467 VSS.n3615 VSS.n3591 0.0119575
R74468 VSS.n6421 VSS.n3608 0.0119575
R74469 VSS.n3614 VSS.n3590 0.0119575
R74470 VSS.n6422 VSS.n3609 0.0119575
R74471 VSS.n3613 VSS.n3589 0.0119575
R74472 VSS.n6423 VSS.n3610 0.0119575
R74473 VSS.n3612 VSS.n3588 0.0119575
R74474 VSS.n6427 VSS.n3611 0.0119575
R74475 VSS.n6637 VSS.n6633 0.0119575
R74476 VSS.n6634 VSS.n3118 0.0119575
R74477 VSS.n6631 VSS.n3117 0.0119575
R74478 VSS.n6639 VSS.n3113 0.0119575
R74479 VSS.n6652 VSS.n6645 0.0119575
R74480 VSS.n6646 VSS.n6644 0.0119575
R74481 VSS.n6648 VSS.n6641 0.0119575
R74482 VSS.n6643 VSS.n6642 0.0119575
R74483 VSS.n3074 VSS.n3062 0.0119575
R74484 VSS.n3080 VSS.n3065 0.0119575
R74485 VSS.n3073 VSS.n3061 0.0119575
R74486 VSS.n3079 VSS.n3066 0.0119575
R74487 VSS.n3072 VSS.n3060 0.0119575
R74488 VSS.n3078 VSS.n3067 0.0119575
R74489 VSS.n3071 VSS.n3059 0.0119575
R74490 VSS.n3077 VSS.n3068 0.0119575
R74491 VSS.n3070 VSS.n3058 0.0119575
R74492 VSS.n6716 VSS.n3069 0.0119575
R74493 VSS.n7021 VSS.n2631 0.0119575
R74494 VSS.n2632 VSS.n2630 0.0119575
R74495 VSS.n7017 VSS.n2627 0.0119575
R74496 VSS.n2629 VSS.n2628 0.0119575
R74497 VSS.n1295 VSS.n1293 0.0119575
R74498 VSS.n1299 VSS.n1297 0.0119575
R74499 VSS.n1298 VSS.n1292 0.0119575
R74500 VSS.n1301 VSS.n1300 0.0119575
R74501 VSS.n1308 VSS.n1290 0.0119575
R74502 VSS.n1307 VSS.n1303 0.0119575
R74503 VSS.n1302 VSS.n1289 0.0119575
R74504 VSS.n8860 VSS.n1304 0.0119575
R74505 VSS.n8040 VSS.n1138 0.0119575
R74506 VSS.n1136 VSS.n1135 0.0119575
R74507 VSS.n1134 VSS.n1133 0.0119575
R74508 VSS.n1132 VSS.n1131 0.0119575
R74509 VSS.n1130 VSS.n1129 0.0119575
R74510 VSS.n1128 VSS.n1127 0.0119575
R74511 VSS.n1126 VSS.n1125 0.0119575
R74512 VSS.n1124 VSS.n1123 0.0119575
R74513 VSS.n1122 VSS.n1121 0.0119575
R74514 VSS.n8578 VSS.n1120 0.0119575
R74515 VSS.n1117 VSS.n1116 0.0119575
R74516 VSS.n1115 VSS.n1114 0.0119575
R74517 VSS.n1113 VSS.n1112 0.0119575
R74518 VSS.n1111 VSS.n1110 0.0119575
R74519 VSS.n1109 VSS.n1108 0.0119575
R74520 VSS.n1107 VSS.n1106 0.0119575
R74521 VSS.n1105 VSS.n1104 0.0119575
R74522 VSS.n1103 VSS.n1096 0.0119575
R74523 VSS.n1097 VSS.n1095 0.0119575
R74524 VSS.n8970 VSS.n1091 0.0119575
R74525 VSS.n9001 VSS.n8986 0.0119575
R74526 VSS.n8984 VSS.n1090 0.0119575
R74527 VSS.n9002 VSS.n8987 0.0119575
R74528 VSS.n8983 VSS.n1089 0.0119575
R74529 VSS.n9003 VSS.n8988 0.0119575
R74530 VSS.n8982 VSS.n1088 0.0119575
R74531 VSS.n9004 VSS.n8989 0.0119575
R74532 VSS.n8981 VSS.n1087 0.0119575
R74533 VSS.n9005 VSS.n8990 0.0119575
R74534 VSS.n8980 VSS.n1086 0.0119575
R74535 VSS.n9006 VSS.n8991 0.0119575
R74536 VSS.n8979 VSS.n1085 0.0119575
R74537 VSS.n9007 VSS.n8992 0.0119575
R74538 VSS.n8978 VSS.n1084 0.0119575
R74539 VSS.n9008 VSS.n8993 0.0119575
R74540 VSS.n8977 VSS.n1083 0.0119575
R74541 VSS.n9009 VSS.n8994 0.0119575
R74542 VSS.n8976 VSS.n1082 0.0119575
R74543 VSS.n9010 VSS.n8995 0.0119575
R74544 VSS.n8975 VSS.n1081 0.0119575
R74545 VSS.n9013 VSS.n9012 0.0119575
R74546 VSS.n8974 VSS.n1080 0.0119575
R74547 VSS.n9015 VSS.n8973 0.0119575
R74548 VSS.n9353 VSS.n797 0.0119575
R74549 VSS.n796 VSS.n793 0.0119575
R74550 VSS.n9354 VSS.n799 0.0119575
R74551 VSS.n798 VSS.n792 0.0119575
R74552 VSS.n9355 VSS.n801 0.0119575
R74553 VSS.n800 VSS.n791 0.0119575
R74554 VSS.n9356 VSS.n803 0.0119575
R74555 VSS.n802 VSS.n790 0.0119575
R74556 VSS.n9357 VSS.n805 0.0119575
R74557 VSS.n804 VSS.n789 0.0119575
R74558 VSS.n9358 VSS.n807 0.0119575
R74559 VSS.n806 VSS.n788 0.0119575
R74560 VSS.n9359 VSS.n809 0.0119575
R74561 VSS.n808 VSS.n787 0.0119575
R74562 VSS.n9360 VSS.n811 0.0119575
R74563 VSS.n810 VSS.n786 0.0119575
R74564 VSS.n9361 VSS.n813 0.0119575
R74565 VSS.n812 VSS.n785 0.0119575
R74566 VSS.n9362 VSS.n815 0.0119575
R74567 VSS.n814 VSS.n784 0.0119575
R74568 VSS.n9366 VSS.n9364 0.0119575
R74569 VSS.n9365 VSS.n783 0.0119575
R74570 VSS.n9368 VSS.n779 0.0119575
R74571 VSS.n9372 VSS.n9369 0.0119575
R74572 VSS.n9438 VSS.n778 0.0119575
R74573 VSS.n9437 VSS.n9373 0.0119575
R74574 VSS.n5393 VSS.n5382 0.0119575
R74575 VSS.n5395 VSS.n5391 0.0119575
R74576 VSS.n5394 VSS.n5381 0.0119575
R74577 VSS.n5523 VSS.n5390 0.0119575
R74578 VSS.n5524 VSS.n5380 0.0119575
R74579 VSS.n5389 VSS.n5388 0.0119575
R74580 VSS.n366 VSS.n352 0.0119575
R74581 VSS.n360 VSS.n350 0.0119575
R74582 VSS.n365 VSS.n353 0.0119575
R74583 VSS.n361 VSS.n349 0.0119575
R74584 VSS.n364 VSS.n354 0.0119575
R74585 VSS.n3074 VSS.n3064 0.0119575
R74586 VSS.n3080 VSS.n3062 0.0119575
R74587 VSS.n3073 VSS.n3065 0.0119575
R74588 VSS.n3079 VSS.n3061 0.0119575
R74589 VSS.n3072 VSS.n3066 0.0119575
R74590 VSS.n3078 VSS.n3060 0.0119575
R74591 VSS.n3071 VSS.n3067 0.0119575
R74592 VSS.n3077 VSS.n3059 0.0119575
R74593 VSS.n3070 VSS.n3068 0.0119575
R74594 VSS.n3069 VSS.n3058 0.0119575
R74595 VSS.n1296 VSS.n1295 0.0119575
R74596 VSS.n1297 VSS.n1293 0.0119575
R74597 VSS.n1299 VSS.n1298 0.0119575
R74598 VSS.n1300 VSS.n1292 0.0119575
R74599 VSS.n8858 VSS.n1290 0.0119575
R74600 VSS.n1308 VSS.n1307 0.0119575
R74601 VSS.n1303 VSS.n1302 0.0119575
R74602 VSS.n1304 VSS.n1289 0.0119575
R74603 VSS.n1352 VSS.n1138 0.0119575
R74604 VSS.n8036 VSS.n1136 0.0119575
R74605 VSS.n1135 VSS.n1134 0.0119575
R74606 VSS.n1133 VSS.n1132 0.0119575
R74607 VSS.n1131 VSS.n1130 0.0119575
R74608 VSS.n1129 VSS.n1128 0.0119575
R74609 VSS.n1127 VSS.n1126 0.0119575
R74610 VSS.n1125 VSS.n1124 0.0119575
R74611 VSS.n1123 VSS.n1122 0.0119575
R74612 VSS.n1121 VSS.n1120 0.0119575
R74613 VSS.n1118 VSS.n1117 0.0119575
R74614 VSS.n1116 VSS.n1115 0.0119575
R74615 VSS.n1114 VSS.n1113 0.0119575
R74616 VSS.n1112 VSS.n1111 0.0119575
R74617 VSS.n1110 VSS.n1109 0.0119575
R74618 VSS.n1108 VSS.n1107 0.0119575
R74619 VSS.n1106 VSS.n1105 0.0119575
R74620 VSS.n1104 VSS.n1103 0.0119575
R74621 VSS.n8986 VSS.n8971 0.0119575
R74622 VSS.n9001 VSS.n1090 0.0119575
R74623 VSS.n9002 VSS.n8984 0.0119575
R74624 VSS.n8987 VSS.n1089 0.0119575
R74625 VSS.n9003 VSS.n8983 0.0119575
R74626 VSS.n8988 VSS.n1088 0.0119575
R74627 VSS.n9004 VSS.n8982 0.0119575
R74628 VSS.n8989 VSS.n1087 0.0119575
R74629 VSS.n9005 VSS.n8981 0.0119575
R74630 VSS.n8990 VSS.n1086 0.0119575
R74631 VSS.n9006 VSS.n8980 0.0119575
R74632 VSS.n8991 VSS.n1085 0.0119575
R74633 VSS.n9007 VSS.n8979 0.0119575
R74634 VSS.n8992 VSS.n1084 0.0119575
R74635 VSS.n9008 VSS.n8978 0.0119575
R74636 VSS.n8993 VSS.n1083 0.0119575
R74637 VSS.n9009 VSS.n8977 0.0119575
R74638 VSS.n8994 VSS.n1082 0.0119575
R74639 VSS.n9010 VSS.n8976 0.0119575
R74640 VSS.n8995 VSS.n1081 0.0119575
R74641 VSS.n9012 VSS.n8975 0.0119575
R74642 VSS.n9013 VSS.n1080 0.0119575
R74643 VSS.n8974 VSS.n8973 0.0119575
R74644 VSS.n9353 VSS.n794 0.0119575
R74645 VSS.n797 VSS.n796 0.0119575
R74646 VSS.n9354 VSS.n793 0.0119575
R74647 VSS.n799 VSS.n798 0.0119575
R74648 VSS.n9355 VSS.n792 0.0119575
R74649 VSS.n801 VSS.n800 0.0119575
R74650 VSS.n9356 VSS.n791 0.0119575
R74651 VSS.n803 VSS.n802 0.0119575
R74652 VSS.n9357 VSS.n790 0.0119575
R74653 VSS.n805 VSS.n804 0.0119575
R74654 VSS.n9358 VSS.n789 0.0119575
R74655 VSS.n807 VSS.n806 0.0119575
R74656 VSS.n9359 VSS.n788 0.0119575
R74657 VSS.n809 VSS.n808 0.0119575
R74658 VSS.n9360 VSS.n787 0.0119575
R74659 VSS.n811 VSS.n810 0.0119575
R74660 VSS.n9361 VSS.n786 0.0119575
R74661 VSS.n813 VSS.n812 0.0119575
R74662 VSS.n9362 VSS.n785 0.0119575
R74663 VSS.n815 VSS.n814 0.0119575
R74664 VSS.n9364 VSS.n784 0.0119575
R74665 VSS.n9366 VSS.n9365 0.0119575
R74666 VSS.n783 VSS.n779 0.0119575
R74667 VSS.n3624 VSS.n3600 0.0119575
R74668 VSS.n6425 VSS.n3626 0.0119575
R74669 VSS.n6414 VSS.n3598 0.0119575
R74670 VSS.n3621 VSS.n3601 0.0119575
R74671 VSS.n6415 VSS.n3597 0.0119575
R74672 VSS.n3620 VSS.n3602 0.0119575
R74673 VSS.n6416 VSS.n3596 0.0119575
R74674 VSS.n3619 VSS.n3603 0.0119575
R74675 VSS.n6417 VSS.n3595 0.0119575
R74676 VSS.n3618 VSS.n3604 0.0119575
R74677 VSS.n6418 VSS.n3594 0.0119575
R74678 VSS.n3617 VSS.n3605 0.0119575
R74679 VSS.n6419 VSS.n3593 0.0119575
R74680 VSS.n3616 VSS.n3606 0.0119575
R74681 VSS.n6420 VSS.n3592 0.0119575
R74682 VSS.n3615 VSS.n3607 0.0119575
R74683 VSS.n6421 VSS.n3591 0.0119575
R74684 VSS.n3614 VSS.n3608 0.0119575
R74685 VSS.n6422 VSS.n3590 0.0119575
R74686 VSS.n3613 VSS.n3609 0.0119575
R74687 VSS.n6423 VSS.n3589 0.0119575
R74688 VSS.n3612 VSS.n3610 0.0119575
R74689 VSS.n3611 VSS.n3588 0.0119575
R74690 VSS.n3327 VSS.n3292 0.0119575
R74691 VSS.n3314 VSS.n3289 0.0119575
R74692 VSS.n3326 VSS.n3293 0.0119575
R74693 VSS.n3313 VSS.n3288 0.0119575
R74694 VSS.n3325 VSS.n3294 0.0119575
R74695 VSS.n3312 VSS.n3287 0.0119575
R74696 VSS.n3324 VSS.n3295 0.0119575
R74697 VSS.n3311 VSS.n3286 0.0119575
R74698 VSS.n3323 VSS.n3296 0.0119575
R74699 VSS.n3310 VSS.n3285 0.0119575
R74700 VSS.n3322 VSS.n3297 0.0119575
R74701 VSS.n3309 VSS.n3284 0.0119575
R74702 VSS.n3321 VSS.n3298 0.0119575
R74703 VSS.n3308 VSS.n3283 0.0119575
R74704 VSS.n3320 VSS.n3299 0.0119575
R74705 VSS.n3307 VSS.n3282 0.0119575
R74706 VSS.n3319 VSS.n3300 0.0119575
R74707 VSS.n3306 VSS.n3281 0.0119575
R74708 VSS.n3318 VSS.n3301 0.0119575
R74709 VSS.n3305 VSS.n3280 0.0119575
R74710 VSS.n3317 VSS.n3302 0.0119575
R74711 VSS.n3304 VSS.n3279 0.0119575
R74712 VSS.n6544 VSS.n3303 0.0119575
R74713 VSS.n6587 VSS.n3221 0.0119575
R74714 VSS.n3222 VSS.n3220 0.0119575
R74715 VSS.n6583 VSS.n3217 0.0119575
R74716 VSS.n3219 VSS.n3218 0.0119575
R74717 VSS.n5785 VSS.n5764 0.0119575
R74718 VSS.n5765 VSS.n5763 0.0119575
R74719 VSS.n5781 VSS.n5760 0.0119575
R74720 VSS.n5762 VSS.n5761 0.0119575
R74721 VSS.n2837 VSS.n2835 0.0119575
R74722 VSS.n6934 VSS.n2840 0.0119575
R74723 VSS.n2839 VSS.n2834 0.0119575
R74724 VSS.n6935 VSS.n2842 0.0119575
R74725 VSS.n2841 VSS.n2833 0.0119575
R74726 VSS.n6936 VSS.n2844 0.0119575
R74727 VSS.n2843 VSS.n2832 0.0119575
R74728 VSS.n6937 VSS.n2846 0.0119575
R74729 VSS.n2845 VSS.n2831 0.0119575
R74730 VSS.n6940 VSS.n6939 0.0119575
R74731 VSS.n6979 VSS.n2765 0.0119575
R74732 VSS.n2766 VSS.n2764 0.0119575
R74733 VSS.n6975 VSS.n2761 0.0119575
R74734 VSS.n2763 VSS.n2762 0.0119575
R74735 VSS.n8321 VSS.n1698 0.0119575
R74736 VSS.n8317 VSS.n1688 0.0119575
R74737 VSS.n8320 VSS.n1697 0.0119575
R74738 VSS.n8318 VSS.n1689 0.0119575
R74739 VSS.n8319 VSS.n1696 0.0119575
R74740 VSS.n8325 VSS.n1690 0.0119575
R74741 VSS.n8324 VSS.n1695 0.0119575
R74742 VSS.n8326 VSS.n1691 0.0119575
R74743 VSS.n8328 VSS.n1693 0.0119575
R74744 VSS.n8329 VSS.n1692 0.0119575
R74745 VSS.n2220 VSS.n2219 0.0119575
R74746 VSS.n2218 VSS.n2217 0.0119575
R74747 VSS.n2216 VSS.n2215 0.0119575
R74748 VSS.n2214 VSS.n2213 0.0119575
R74749 VSS.n2212 VSS.n2211 0.0119575
R74750 VSS.n2210 VSS.n2209 0.0119575
R74751 VSS.n2208 VSS.n2207 0.0119575
R74752 VSS.n2206 VSS.n2205 0.0119575
R74753 VSS.n2204 VSS.n2203 0.0119575
R74754 VSS.n2202 VSS.n2201 0.0119575
R74755 VSS.n2200 VSS.n2199 0.0119575
R74756 VSS.n2198 VSS.n2197 0.0119575
R74757 VSS.n2196 VSS.n2195 0.0119575
R74758 VSS.n2194 VSS.n2193 0.0119575
R74759 VSS.n2192 VSS.n2191 0.0119575
R74760 VSS.n2190 VSS.n2189 0.0119575
R74761 VSS.n2188 VSS.n2187 0.0119575
R74762 VSS.n2186 VSS.n2185 0.0119575
R74763 VSS.n2184 VSS.n2183 0.0119575
R74764 VSS.n2182 VSS.n2181 0.0119575
R74765 VSS.n2180 VSS.n2179 0.0119575
R74766 VSS.n2178 VSS.n2173 0.0119575
R74767 VSS.n3327 VSS.n3290 0.0119575
R74768 VSS.n3314 VSS.n3292 0.0119575
R74769 VSS.n3326 VSS.n3289 0.0119575
R74770 VSS.n3313 VSS.n3293 0.0119575
R74771 VSS.n3325 VSS.n3288 0.0119575
R74772 VSS.n3312 VSS.n3294 0.0119575
R74773 VSS.n3324 VSS.n3287 0.0119575
R74774 VSS.n3311 VSS.n3295 0.0119575
R74775 VSS.n3323 VSS.n3286 0.0119575
R74776 VSS.n3310 VSS.n3296 0.0119575
R74777 VSS.n3322 VSS.n3285 0.0119575
R74778 VSS.n3309 VSS.n3297 0.0119575
R74779 VSS.n3321 VSS.n3284 0.0119575
R74780 VSS.n3308 VSS.n3298 0.0119575
R74781 VSS.n3320 VSS.n3283 0.0119575
R74782 VSS.n3307 VSS.n3299 0.0119575
R74783 VSS.n3319 VSS.n3282 0.0119575
R74784 VSS.n3306 VSS.n3300 0.0119575
R74785 VSS.n3318 VSS.n3281 0.0119575
R74786 VSS.n3305 VSS.n3301 0.0119575
R74787 VSS.n3317 VSS.n3280 0.0119575
R74788 VSS.n3304 VSS.n3302 0.0119575
R74789 VSS.n3303 VSS.n3279 0.0119575
R74790 VSS.n2838 VSS.n2837 0.0119575
R74791 VSS.n6934 VSS.n2835 0.0119575
R74792 VSS.n2840 VSS.n2839 0.0119575
R74793 VSS.n6935 VSS.n2834 0.0119575
R74794 VSS.n2842 VSS.n2841 0.0119575
R74795 VSS.n6936 VSS.n2833 0.0119575
R74796 VSS.n2844 VSS.n2843 0.0119575
R74797 VSS.n6937 VSS.n2832 0.0119575
R74798 VSS.n2846 VSS.n2845 0.0119575
R74799 VSS.n6939 VSS.n2831 0.0119575
R74800 VSS.n8321 VSS.n1687 0.0119575
R74801 VSS.n1698 VSS.n1688 0.0119575
R74802 VSS.n8320 VSS.n8317 0.0119575
R74803 VSS.n1697 VSS.n1689 0.0119575
R74804 VSS.n8319 VSS.n8318 0.0119575
R74805 VSS.n1696 VSS.n1690 0.0119575
R74806 VSS.n8325 VSS.n8324 0.0119575
R74807 VSS.n1695 VSS.n1691 0.0119575
R74808 VSS.n8326 VSS.n1693 0.0119575
R74809 VSS.n8329 VSS.n8328 0.0119575
R74810 VSS.n2221 VSS.n2220 0.0119575
R74811 VSS.n2219 VSS.n2218 0.0119575
R74812 VSS.n2217 VSS.n2216 0.0119575
R74813 VSS.n2215 VSS.n2214 0.0119575
R74814 VSS.n2213 VSS.n2212 0.0119575
R74815 VSS.n2211 VSS.n2210 0.0119575
R74816 VSS.n2209 VSS.n2208 0.0119575
R74817 VSS.n2207 VSS.n2206 0.0119575
R74818 VSS.n2205 VSS.n2204 0.0119575
R74819 VSS.n2203 VSS.n2202 0.0119575
R74820 VSS.n2201 VSS.n2200 0.0119575
R74821 VSS.n2199 VSS.n2198 0.0119575
R74822 VSS.n2197 VSS.n2196 0.0119575
R74823 VSS.n2195 VSS.n2194 0.0119575
R74824 VSS.n2193 VSS.n2192 0.0119575
R74825 VSS.n2191 VSS.n2190 0.0119575
R74826 VSS.n2189 VSS.n2188 0.0119575
R74827 VSS.n2187 VSS.n2186 0.0119575
R74828 VSS.n2185 VSS.n2184 0.0119575
R74829 VSS.n2183 VSS.n2182 0.0119575
R74830 VSS.n2181 VSS.n2180 0.0119575
R74831 VSS.n2179 VSS.n2178 0.0119575
R74832 VSS.n4676 VSS.n4627 0.0119575
R74833 VSS.n4680 VSS.n4621 0.0119575
R74834 VSS.n4629 VSS.n4625 0.0119575
R74835 VSS.n4679 VSS.n4620 0.0119575
R74836 VSS.n4630 VSS.n4626 0.0119575
R74837 VSS.n4678 VSS.n4619 0.0119575
R74838 VSS.n4576 VSS.n4557 0.0119575
R74839 VSS.n4781 VSS.n4780 0.0119575
R74840 VSS.n4575 VSS.n4556 0.0119575
R74841 VSS.n4783 VSS.n4782 0.0119575
R74842 VSS.n4574 VSS.n4555 0.0119575
R74843 VSS.n4573 VSS.n4559 0.0119575
R74844 VSS.n4576 VSS.n4558 0.0119575
R74845 VSS.n4780 VSS.n4557 0.0119575
R74846 VSS.n4781 VSS.n4556 0.0119575
R74847 VSS.n4782 VSS.n4575 0.0119575
R74848 VSS.n4783 VSS.n4555 0.0119575
R74849 VSS.n4574 VSS.n4573 0.0119575
R74850 VSS.n9749 VSS.n9748 0.0119575
R74851 VSS.n9750 VSS.n232 0.0119575
R74852 VSS.n9752 VSS.n9751 0.0119575
R74853 VSS.n9753 VSS.n231 0.0119575
R74854 VSS.n9755 VSS.n9754 0.0119575
R74855 VSS.n9756 VSS.n230 0.0119575
R74856 VSS.n36 VSS.n22 0.0119575
R74857 VSS.n40 VSS.n32 0.0119575
R74858 VSS.n43 VSS.n42 0.0119575
R74859 VSS.n45 VSS.n39 0.0119575
R74860 VSS.n9891 VSS.n44 0.0119575
R74861 VSS.n9890 VSS.n38 0.0119575
R74862 VSS.n262 VSS.n258 0.0119575
R74863 VSS.n264 VSS.n257 0.0119575
R74864 VSS.n267 VSS.n261 0.0119575
R74865 VSS.n265 VSS.n256 0.0119575
R74866 VSS.n266 VSS.n260 0.0119575
R74867 VSS.n9693 VSS.n255 0.0119575
R74868 VSS.n299 VSS.n293 0.0119575
R74869 VSS.n303 VSS.n301 0.0119575
R74870 VSS.n302 VSS.n292 0.0119575
R74871 VSS.n306 VSS.n304 0.0119575
R74872 VSS.n305 VSS.n291 0.0119575
R74873 VSS.n9682 VSS.n307 0.0119575
R74874 VSS.n316 VSS.n308 0.0119575
R74875 VSS.n319 VSS.n318 0.0119575
R74876 VSS.n327 VSS.n315 0.0119575
R74877 VSS.n321 VSS.n320 0.0119575
R74878 VSS.n326 VSS.n314 0.0119575
R74879 VSS.n5951 VSS.n5950 0.0119575
R74880 VSS.n5948 VSS.n5912 0.0119575
R74881 VSS.n5916 VSS.n5910 0.0119575
R74882 VSS.n5947 VSS.n5946 0.0119575
R74883 VSS.n6322 VSS.n3702 0.0119575
R74884 VSS.n3703 VSS.n3701 0.0119575
R74885 VSS.n6318 VSS.n3698 0.0119575
R74886 VSS.n3700 VSS.n3699 0.0119575
R74887 VSS.n3551 VSS.n3527 0.0119575
R74888 VSS.n3549 VSS.n3524 0.0119575
R74889 VSS.n3552 VSS.n3528 0.0119575
R74890 VSS.n3548 VSS.n3523 0.0119575
R74891 VSS.n3553 VSS.n3529 0.0119575
R74892 VSS.n3547 VSS.n3522 0.0119575
R74893 VSS.n3554 VSS.n3530 0.0119575
R74894 VSS.n3546 VSS.n3521 0.0119575
R74895 VSS.n3555 VSS.n3531 0.0119575
R74896 VSS.n3545 VSS.n3520 0.0119575
R74897 VSS.n3556 VSS.n3532 0.0119575
R74898 VSS.n3544 VSS.n3519 0.0119575
R74899 VSS.n3557 VSS.n3533 0.0119575
R74900 VSS.n3543 VSS.n3518 0.0119575
R74901 VSS.n3558 VSS.n3534 0.0119575
R74902 VSS.n3542 VSS.n3517 0.0119575
R74903 VSS.n3559 VSS.n3535 0.0119575
R74904 VSS.n3541 VSS.n3516 0.0119575
R74905 VSS.n3560 VSS.n3536 0.0119575
R74906 VSS.n3540 VSS.n3515 0.0119575
R74907 VSS.n3561 VSS.n3537 0.0119575
R74908 VSS.n3539 VSS.n3514 0.0119575
R74909 VSS.n6452 VSS.n3538 0.0119575
R74910 VSS.n6628 VSS.n3124 0.0119575
R74911 VSS.n3125 VSS.n3123 0.0119575
R74912 VSS.n6624 VSS.n3122 0.0119575
R74913 VSS.n3121 VSS.n2966 0.0119575
R74914 VSS.n6759 VSS.n2965 0.0119575
R74915 VSS.n6756 VSS.n6754 0.0119575
R74916 VSS.n2969 VSS.n2963 0.0119575
R74917 VSS.n6753 VSS.n2971 0.0119575
R74918 VSS.n2980 VSS.n2972 0.0119575
R74919 VSS.n2983 VSS.n2982 0.0119575
R74920 VSS.n2994 VSS.n2979 0.0119575
R74921 VSS.n2985 VSS.n2984 0.0119575
R74922 VSS.n2993 VSS.n2978 0.0119575
R74923 VSS.n2987 VSS.n2986 0.0119575
R74924 VSS.n2992 VSS.n2977 0.0119575
R74925 VSS.n2989 VSS.n2988 0.0119575
R74926 VSS.n2991 VSS.n2976 0.0119575
R74927 VSS.n6750 VSS.n2990 0.0119575
R74928 VSS.n7014 VSS.n2640 0.0119575
R74929 VSS.n2641 VSS.n2639 0.0119575
R74930 VSS.n7010 VSS.n2636 0.0119575
R74931 VSS.n2638 VSS.n2637 0.0119575
R74932 VSS.n1332 VSS.n1330 0.0119575
R74933 VSS.n1336 VSS.n1334 0.0119575
R74934 VSS.n1335 VSS.n1329 0.0119575
R74935 VSS.n1338 VSS.n1337 0.0119575
R74936 VSS.n1328 VSS.n1327 0.0119575
R74937 VSS.n1341 VSS.n1339 0.0119575
R74938 VSS.n1340 VSS.n1326 0.0119575
R74939 VSS.n8841 VSS.n1342 0.0119575
R74940 VSS.n1408 VSS.n1392 0.0119575
R74941 VSS.n1409 VSS.n1405 0.0119575
R74942 VSS.n8795 VSS.n1412 0.0119575
R74943 VSS.n1411 VSS.n1404 0.0119575
R74944 VSS.n8796 VSS.n1414 0.0119575
R74945 VSS.n1413 VSS.n1403 0.0119575
R74946 VSS.n8797 VSS.n1416 0.0119575
R74947 VSS.n1415 VSS.n1402 0.0119575
R74948 VSS.n8798 VSS.n1418 0.0119575
R74949 VSS.n1417 VSS.n1401 0.0119575
R74950 VSS.n8799 VSS.n1421 0.0119575
R74951 VSS.n1420 VSS.n1399 0.0119575
R74952 VSS.n8800 VSS.n1423 0.0119575
R74953 VSS.n1422 VSS.n1398 0.0119575
R74954 VSS.n8801 VSS.n1425 0.0119575
R74955 VSS.n1424 VSS.n1397 0.0119575
R74956 VSS.n8802 VSS.n1427 0.0119575
R74957 VSS.n1426 VSS.n1396 0.0119575
R74958 VSS.n2460 VSS.n2459 0.0119575
R74959 VSS.n2454 VSS.n2452 0.0119575
R74960 VSS.n9039 VSS.n1045 0.0119575
R74961 VSS.n1043 VSS.n1031 0.0119575
R74962 VSS.n9040 VSS.n1046 0.0119575
R74963 VSS.n1042 VSS.n1030 0.0119575
R74964 VSS.n9041 VSS.n1047 0.0119575
R74965 VSS.n1041 VSS.n1029 0.0119575
R74966 VSS.n9042 VSS.n1048 0.0119575
R74967 VSS.n1040 VSS.n1028 0.0119575
R74968 VSS.n9043 VSS.n1049 0.0119575
R74969 VSS.n1039 VSS.n1027 0.0119575
R74970 VSS.n9044 VSS.n1050 0.0119575
R74971 VSS.n1038 VSS.n1026 0.0119575
R74972 VSS.n9045 VSS.n1051 0.0119575
R74973 VSS.n1037 VSS.n1025 0.0119575
R74974 VSS.n9046 VSS.n1052 0.0119575
R74975 VSS.n1036 VSS.n1024 0.0119575
R74976 VSS.n9047 VSS.n1053 0.0119575
R74977 VSS.n1035 VSS.n1023 0.0119575
R74978 VSS.n9048 VSS.n1054 0.0119575
R74979 VSS.n1034 VSS.n1022 0.0119575
R74980 VSS.n9052 VSS.n9051 0.0119575
R74981 VSS.n1033 VSS.n1021 0.0119575
R74982 VSS.n9049 VSS.n843 0.0119575
R74983 VSS.n9288 VSS.n844 0.0119575
R74984 VSS.n856 VSS.n842 0.0119575
R74985 VSS.n9299 VSS.n9289 0.0119575
R74986 VSS.n855 VSS.n841 0.0119575
R74987 VSS.n9300 VSS.n9290 0.0119575
R74988 VSS.n854 VSS.n840 0.0119575
R74989 VSS.n9301 VSS.n9291 0.0119575
R74990 VSS.n853 VSS.n839 0.0119575
R74991 VSS.n9302 VSS.n9292 0.0119575
R74992 VSS.n852 VSS.n838 0.0119575
R74993 VSS.n9303 VSS.n9293 0.0119575
R74994 VSS.n851 VSS.n837 0.0119575
R74995 VSS.n9304 VSS.n9294 0.0119575
R74996 VSS.n850 VSS.n836 0.0119575
R74997 VSS.n9305 VSS.n9295 0.0119575
R74998 VSS.n849 VSS.n835 0.0119575
R74999 VSS.n9306 VSS.n9296 0.0119575
R75000 VSS.n848 VSS.n834 0.0119575
R75001 VSS.n9307 VSS.n9297 0.0119575
R75002 VSS.n847 VSS.n833 0.0119575
R75003 VSS.n9311 VSS.n9310 0.0119575
R75004 VSS.n846 VSS.n832 0.0119575
R75005 VSS.n9308 VSS.n771 0.0119575
R75006 VSS.n775 VSS.n772 0.0119575
R75007 VSS.n9443 VSS.n770 0.0119575
R75008 VSS.n9442 VSS.n776 0.0119575
R75009 VSS.n9695 VSS.n258 0.0119575
R75010 VSS.n262 VSS.n257 0.0119575
R75011 VSS.n267 VSS.n264 0.0119575
R75012 VSS.n261 VSS.n256 0.0119575
R75013 VSS.n266 VSS.n265 0.0119575
R75014 VSS.n260 VSS.n255 0.0119575
R75015 VSS.n300 VSS.n299 0.0119575
R75016 VSS.n301 VSS.n293 0.0119575
R75017 VSS.n303 VSS.n302 0.0119575
R75018 VSS.n304 VSS.n292 0.0119575
R75019 VSS.n306 VSS.n305 0.0119575
R75020 VSS.n307 VSS.n291 0.0119575
R75021 VSS.n9681 VSS.n308 0.0119575
R75022 VSS.n318 VSS.n316 0.0119575
R75023 VSS.n327 VSS.n319 0.0119575
R75024 VSS.n320 VSS.n315 0.0119575
R75025 VSS.n326 VSS.n321 0.0119575
R75026 VSS.n3551 VSS.n3525 0.0119575
R75027 VSS.n3549 VSS.n3527 0.0119575
R75028 VSS.n3552 VSS.n3524 0.0119575
R75029 VSS.n3548 VSS.n3528 0.0119575
R75030 VSS.n3553 VSS.n3523 0.0119575
R75031 VSS.n3547 VSS.n3529 0.0119575
R75032 VSS.n3554 VSS.n3522 0.0119575
R75033 VSS.n3546 VSS.n3530 0.0119575
R75034 VSS.n3555 VSS.n3521 0.0119575
R75035 VSS.n3545 VSS.n3531 0.0119575
R75036 VSS.n3556 VSS.n3520 0.0119575
R75037 VSS.n3544 VSS.n3532 0.0119575
R75038 VSS.n3557 VSS.n3519 0.0119575
R75039 VSS.n3543 VSS.n3533 0.0119575
R75040 VSS.n3558 VSS.n3518 0.0119575
R75041 VSS.n3542 VSS.n3534 0.0119575
R75042 VSS.n3559 VSS.n3517 0.0119575
R75043 VSS.n3541 VSS.n3535 0.0119575
R75044 VSS.n3560 VSS.n3516 0.0119575
R75045 VSS.n3540 VSS.n3536 0.0119575
R75046 VSS.n3561 VSS.n3515 0.0119575
R75047 VSS.n3539 VSS.n3537 0.0119575
R75048 VSS.n3538 VSS.n3514 0.0119575
R75049 VSS.n6752 VSS.n2972 0.0119575
R75050 VSS.n2982 VSS.n2980 0.0119575
R75051 VSS.n2994 VSS.n2983 0.0119575
R75052 VSS.n2984 VSS.n2979 0.0119575
R75053 VSS.n2993 VSS.n2985 0.0119575
R75054 VSS.n2986 VSS.n2978 0.0119575
R75055 VSS.n2992 VSS.n2987 0.0119575
R75056 VSS.n2988 VSS.n2977 0.0119575
R75057 VSS.n2991 VSS.n2989 0.0119575
R75058 VSS.n2990 VSS.n2976 0.0119575
R75059 VSS.n1333 VSS.n1332 0.0119575
R75060 VSS.n1334 VSS.n1330 0.0119575
R75061 VSS.n1336 VSS.n1335 0.0119575
R75062 VSS.n1337 VSS.n1329 0.0119575
R75063 VSS.n1327 VSS.n1318 0.0119575
R75064 VSS.n1339 VSS.n1328 0.0119575
R75065 VSS.n1341 VSS.n1340 0.0119575
R75066 VSS.n1342 VSS.n1326 0.0119575
R75067 VSS.n8806 VSS.n1392 0.0119575
R75068 VSS.n1410 VSS.n1409 0.0119575
R75069 VSS.n8795 VSS.n1405 0.0119575
R75070 VSS.n1412 VSS.n1411 0.0119575
R75071 VSS.n8796 VSS.n1404 0.0119575
R75072 VSS.n1414 VSS.n1413 0.0119575
R75073 VSS.n8797 VSS.n1403 0.0119575
R75074 VSS.n1416 VSS.n1415 0.0119575
R75075 VSS.n8798 VSS.n1402 0.0119575
R75076 VSS.n1418 VSS.n1417 0.0119575
R75077 VSS.n8799 VSS.n1400 0.0119575
R75078 VSS.n1421 VSS.n1420 0.0119575
R75079 VSS.n8800 VSS.n1399 0.0119575
R75080 VSS.n1423 VSS.n1422 0.0119575
R75081 VSS.n8801 VSS.n1398 0.0119575
R75082 VSS.n1425 VSS.n1424 0.0119575
R75083 VSS.n8802 VSS.n1397 0.0119575
R75084 VSS.n1427 VSS.n1426 0.0119575
R75085 VSS.n1045 VSS.n1032 0.0119575
R75086 VSS.n9039 VSS.n1031 0.0119575
R75087 VSS.n9040 VSS.n1043 0.0119575
R75088 VSS.n1046 VSS.n1030 0.0119575
R75089 VSS.n9041 VSS.n1042 0.0119575
R75090 VSS.n1047 VSS.n1029 0.0119575
R75091 VSS.n9042 VSS.n1041 0.0119575
R75092 VSS.n1048 VSS.n1028 0.0119575
R75093 VSS.n9043 VSS.n1040 0.0119575
R75094 VSS.n1049 VSS.n1027 0.0119575
R75095 VSS.n9044 VSS.n1039 0.0119575
R75096 VSS.n1050 VSS.n1026 0.0119575
R75097 VSS.n9045 VSS.n1038 0.0119575
R75098 VSS.n1051 VSS.n1025 0.0119575
R75099 VSS.n9046 VSS.n1037 0.0119575
R75100 VSS.n1052 VSS.n1024 0.0119575
R75101 VSS.n9047 VSS.n1036 0.0119575
R75102 VSS.n1053 VSS.n1023 0.0119575
R75103 VSS.n9048 VSS.n1035 0.0119575
R75104 VSS.n1054 VSS.n1022 0.0119575
R75105 VSS.n9051 VSS.n1034 0.0119575
R75106 VSS.n9052 VSS.n1021 0.0119575
R75107 VSS.n9049 VSS.n1033 0.0119575
R75108 VSS.n9313 VSS.n844 0.0119575
R75109 VSS.n9288 VSS.n842 0.0119575
R75110 VSS.n9299 VSS.n856 0.0119575
R75111 VSS.n9289 VSS.n841 0.0119575
R75112 VSS.n9300 VSS.n855 0.0119575
R75113 VSS.n9290 VSS.n840 0.0119575
R75114 VSS.n9301 VSS.n854 0.0119575
R75115 VSS.n9291 VSS.n839 0.0119575
R75116 VSS.n9302 VSS.n853 0.0119575
R75117 VSS.n9292 VSS.n838 0.0119575
R75118 VSS.n9303 VSS.n852 0.0119575
R75119 VSS.n9293 VSS.n837 0.0119575
R75120 VSS.n9304 VSS.n851 0.0119575
R75121 VSS.n9294 VSS.n836 0.0119575
R75122 VSS.n9305 VSS.n850 0.0119575
R75123 VSS.n9295 VSS.n835 0.0119575
R75124 VSS.n9306 VSS.n849 0.0119575
R75125 VSS.n9296 VSS.n834 0.0119575
R75126 VSS.n9307 VSS.n848 0.0119575
R75127 VSS.n9297 VSS.n833 0.0119575
R75128 VSS.n9310 VSS.n847 0.0119575
R75129 VSS.n9311 VSS.n832 0.0119575
R75130 VSS.n9308 VSS.n846 0.0119575
R75131 VSS.n4396 VSS.n4390 0.0119575
R75132 VSS.n4400 VSS.n4384 0.0119575
R75133 VSS.n4392 VSS.n4388 0.0119575
R75134 VSS.n4399 VSS.n4383 0.0119575
R75135 VSS.n4393 VSS.n4389 0.0119575
R75136 VSS.n4398 VSS.n4382 0.0119575
R75137 VSS.n5061 VSS.n4528 0.0119575
R75138 VSS.n5065 VSS.n5063 0.0119575
R75139 VSS.n5064 VSS.n4527 0.0119575
R75140 VSS.n5068 VSS.n5066 0.0119575
R75141 VSS.n5067 VSS.n4526 0.0119575
R75142 VSS.n5070 VSS.n5069 0.0119575
R75143 VSS.n5631 VSS.n4295 0.0119575
R75144 VSS.n5635 VSS.n5633 0.0119575
R75145 VSS.n5634 VSS.n4294 0.0119575
R75146 VSS.n5638 VSS.n5636 0.0119575
R75147 VSS.n5637 VSS.n4293 0.0119575
R75148 VSS.n5640 VSS.n5639 0.0119575
R75149 VSS.n3987 VSS.n3985 0.0119575
R75150 VSS.n6157 VSS.n3990 0.0119575
R75151 VSS.n3989 VSS.n3984 0.0119575
R75152 VSS.n6158 VSS.n3992 0.0119575
R75153 VSS.n3991 VSS.n3983 0.0119575
R75154 VSS.n6074 VSS.n6043 0.0119575
R75155 VSS.n6044 VSS.n6042 0.0119575
R75156 VSS.n6070 VSS.n6039 0.0119575
R75157 VSS.n6041 VSS.n6040 0.0119575
R75158 VSS.n6300 VSS.n3806 0.0119575
R75159 VSS.n3807 VSS.n3805 0.0119575
R75160 VSS.n6296 VSS.n3802 0.0119575
R75161 VSS.n3804 VSS.n3803 0.0119575
R75162 VSS.n3452 VSS.n3428 0.0119575
R75163 VSS.n3450 VSS.n3425 0.0119575
R75164 VSS.n3453 VSS.n3429 0.0119575
R75165 VSS.n3449 VSS.n3424 0.0119575
R75166 VSS.n3454 VSS.n3430 0.0119575
R75167 VSS.n3448 VSS.n3423 0.0119575
R75168 VSS.n3455 VSS.n3431 0.0119575
R75169 VSS.n3447 VSS.n3422 0.0119575
R75170 VSS.n3456 VSS.n3432 0.0119575
R75171 VSS.n3446 VSS.n3421 0.0119575
R75172 VSS.n3457 VSS.n3433 0.0119575
R75173 VSS.n3445 VSS.n3420 0.0119575
R75174 VSS.n3458 VSS.n3434 0.0119575
R75175 VSS.n3444 VSS.n3419 0.0119575
R75176 VSS.n3459 VSS.n3435 0.0119575
R75177 VSS.n3443 VSS.n3418 0.0119575
R75178 VSS.n3460 VSS.n3436 0.0119575
R75179 VSS.n3442 VSS.n3417 0.0119575
R75180 VSS.n3461 VSS.n3437 0.0119575
R75181 VSS.n3441 VSS.n3416 0.0119575
R75182 VSS.n3462 VSS.n3438 0.0119575
R75183 VSS.n3440 VSS.n3415 0.0119575
R75184 VSS.n6506 VSS.n3439 0.0119575
R75185 VSS.n6600 VSS.n3203 0.0119575
R75186 VSS.n3204 VSS.n3202 0.0119575
R75187 VSS.n6596 VSS.n3199 0.0119575
R75188 VSS.n3201 VSS.n3200 0.0119575
R75189 VSS.n5798 VSS.n5746 0.0119575
R75190 VSS.n5747 VSS.n5745 0.0119575
R75191 VSS.n5794 VSS.n5742 0.0119575
R75192 VSS.n5744 VSS.n5743 0.0119575
R75193 VSS.n2897 VSS.n2895 0.0119575
R75194 VSS.n6872 VSS.n2900 0.0119575
R75195 VSS.n2899 VSS.n2894 0.0119575
R75196 VSS.n6873 VSS.n2902 0.0119575
R75197 VSS.n2901 VSS.n2893 0.0119575
R75198 VSS.n6874 VSS.n2904 0.0119575
R75199 VSS.n2903 VSS.n2892 0.0119575
R75200 VSS.n6875 VSS.n2906 0.0119575
R75201 VSS.n2905 VSS.n2891 0.0119575
R75202 VSS.n6878 VSS.n6877 0.0119575
R75203 VSS.n6992 VSS.n2747 0.0119575
R75204 VSS.n2748 VSS.n2746 0.0119575
R75205 VSS.n6988 VSS.n2743 0.0119575
R75206 VSS.n2745 VSS.n2744 0.0119575
R75207 VSS.n8383 VSS.n8382 0.0119575
R75208 VSS.n8380 VSS.n1660 0.0119575
R75209 VSS.n8381 VSS.n8379 0.0119575
R75210 VSS.n8405 VSS.n1661 0.0119575
R75211 VSS.n1663 VSS.n1657 0.0119575
R75212 VSS.n8407 VSS.n8406 0.0119575
R75213 VSS.n8408 VSS.n1656 0.0119575
R75214 VSS.n8409 VSS.n1602 0.0119575
R75215 VSS.n8610 VSS.n1536 0.0119575
R75216 VSS.n1537 VSS.n1533 0.0119575
R75217 VSS.n8612 VSS.n8611 0.0119575
R75218 VSS.n8614 VSS.n1532 0.0119575
R75219 VSS.n8615 VSS.n8613 0.0119575
R75220 VSS.n8617 VSS.n1531 0.0119575
R75221 VSS.n8618 VSS.n8616 0.0119575
R75222 VSS.n8620 VSS.n1530 0.0119575
R75223 VSS.n8621 VSS.n8619 0.0119575
R75224 VSS.n8608 VSS.n1529 0.0119575
R75225 VSS.n8623 VSS.n8622 0.0119575
R75226 VSS.n8625 VSS.n1527 0.0119575
R75227 VSS.n8626 VSS.n8624 0.0119575
R75228 VSS.n8628 VSS.n1526 0.0119575
R75229 VSS.n8629 VSS.n8627 0.0119575
R75230 VSS.n8631 VSS.n1525 0.0119575
R75231 VSS.n8632 VSS.n8630 0.0119575
R75232 VSS.n1544 VSS.n1524 0.0119575
R75233 VSS.n2432 VSS.n2431 0.0119575
R75234 VSS.n2436 VSS.n2430 0.0119575
R75235 VSS.n1997 VSS.n1995 0.0119575
R75236 VSS.n1996 VSS.n1992 0.0119575
R75237 VSS.n8150 VSS.n1999 0.0119575
R75238 VSS.n1998 VSS.n1991 0.0119575
R75239 VSS.n8151 VSS.n2001 0.0119575
R75240 VSS.n2000 VSS.n1990 0.0119575
R75241 VSS.n8152 VSS.n2003 0.0119575
R75242 VSS.n2002 VSS.n1989 0.0119575
R75243 VSS.n8153 VSS.n2005 0.0119575
R75244 VSS.n2004 VSS.n1988 0.0119575
R75245 VSS.n8154 VSS.n2007 0.0119575
R75246 VSS.n2006 VSS.n1987 0.0119575
R75247 VSS.n8155 VSS.n2009 0.0119575
R75248 VSS.n2008 VSS.n1986 0.0119575
R75249 VSS.n8156 VSS.n2011 0.0119575
R75250 VSS.n2010 VSS.n1985 0.0119575
R75251 VSS.n8157 VSS.n2013 0.0119575
R75252 VSS.n2012 VSS.n1984 0.0119575
R75253 VSS.n8158 VSS.n2015 0.0119575
R75254 VSS.n2014 VSS.n1983 0.0119575
R75255 VSS.n8162 VSS.n8160 0.0119575
R75256 VSS.n8161 VSS.n1982 0.0119575
R75257 VSS.n8164 VSS.n1978 0.0119575
R75258 VSS.n8167 VSS.n1955 0.0119575
R75259 VSS.n8184 VSS.n1977 0.0119575
R75260 VSS.n8168 VSS.n1956 0.0119575
R75261 VSS.n8183 VSS.n1976 0.0119575
R75262 VSS.n8169 VSS.n1957 0.0119575
R75263 VSS.n8182 VSS.n1975 0.0119575
R75264 VSS.n8170 VSS.n1958 0.0119575
R75265 VSS.n8181 VSS.n1974 0.0119575
R75266 VSS.n8171 VSS.n1959 0.0119575
R75267 VSS.n8180 VSS.n1973 0.0119575
R75268 VSS.n8172 VSS.n1960 0.0119575
R75269 VSS.n8179 VSS.n1972 0.0119575
R75270 VSS.n8173 VSS.n1961 0.0119575
R75271 VSS.n8178 VSS.n1971 0.0119575
R75272 VSS.n8174 VSS.n1962 0.0119575
R75273 VSS.n8177 VSS.n1970 0.0119575
R75274 VSS.n8175 VSS.n1963 0.0119575
R75275 VSS.n8176 VSS.n1969 0.0119575
R75276 VSS.n8196 VSS.n1964 0.0119575
R75277 VSS.n8195 VSS.n1968 0.0119575
R75278 VSS.n8197 VSS.n1965 0.0119575
R75279 VSS.n8199 VSS.n1967 0.0119575
R75280 VSS.n8200 VSS.n1966 0.0119575
R75281 VSS.n2347 VSS.n2344 0.0119575
R75282 VSS.n2358 VSS.n2343 0.0119575
R75283 VSS.n2357 VSS.n2348 0.0119575
R75284 VSS.n5062 VSS.n5061 0.0119575
R75285 VSS.n5063 VSS.n4528 0.0119575
R75286 VSS.n5065 VSS.n5064 0.0119575
R75287 VSS.n5066 VSS.n4527 0.0119575
R75288 VSS.n5068 VSS.n5067 0.0119575
R75289 VSS.n5069 VSS.n4526 0.0119575
R75290 VSS.n5632 VSS.n5631 0.0119575
R75291 VSS.n5633 VSS.n4295 0.0119575
R75292 VSS.n5635 VSS.n5634 0.0119575
R75293 VSS.n5636 VSS.n4294 0.0119575
R75294 VSS.n5638 VSS.n5637 0.0119575
R75295 VSS.n5639 VSS.n4293 0.0119575
R75296 VSS.n3988 VSS.n3987 0.0119575
R75297 VSS.n6157 VSS.n3985 0.0119575
R75298 VSS.n3990 VSS.n3989 0.0119575
R75299 VSS.n6158 VSS.n3984 0.0119575
R75300 VSS.n3992 VSS.n3991 0.0119575
R75301 VSS.n3452 VSS.n3426 0.0119575
R75302 VSS.n3450 VSS.n3428 0.0119575
R75303 VSS.n3453 VSS.n3425 0.0119575
R75304 VSS.n3449 VSS.n3429 0.0119575
R75305 VSS.n3454 VSS.n3424 0.0119575
R75306 VSS.n3448 VSS.n3430 0.0119575
R75307 VSS.n3455 VSS.n3423 0.0119575
R75308 VSS.n3447 VSS.n3431 0.0119575
R75309 VSS.n3456 VSS.n3422 0.0119575
R75310 VSS.n3446 VSS.n3432 0.0119575
R75311 VSS.n3457 VSS.n3421 0.0119575
R75312 VSS.n3445 VSS.n3433 0.0119575
R75313 VSS.n3458 VSS.n3420 0.0119575
R75314 VSS.n3444 VSS.n3434 0.0119575
R75315 VSS.n3459 VSS.n3419 0.0119575
R75316 VSS.n3443 VSS.n3435 0.0119575
R75317 VSS.n3460 VSS.n3418 0.0119575
R75318 VSS.n3442 VSS.n3436 0.0119575
R75319 VSS.n3461 VSS.n3417 0.0119575
R75320 VSS.n3441 VSS.n3437 0.0119575
R75321 VSS.n3462 VSS.n3416 0.0119575
R75322 VSS.n3440 VSS.n3438 0.0119575
R75323 VSS.n3439 VSS.n3415 0.0119575
R75324 VSS.n2898 VSS.n2897 0.0119575
R75325 VSS.n6872 VSS.n2895 0.0119575
R75326 VSS.n2900 VSS.n2899 0.0119575
R75327 VSS.n6873 VSS.n2894 0.0119575
R75328 VSS.n2902 VSS.n2901 0.0119575
R75329 VSS.n6874 VSS.n2893 0.0119575
R75330 VSS.n2904 VSS.n2903 0.0119575
R75331 VSS.n6875 VSS.n2892 0.0119575
R75332 VSS.n2906 VSS.n2905 0.0119575
R75333 VSS.n6877 VSS.n2891 0.0119575
R75334 VSS.n8383 VSS.n1659 0.0119575
R75335 VSS.n8382 VSS.n1660 0.0119575
R75336 VSS.n8381 VSS.n8380 0.0119575
R75337 VSS.n8379 VSS.n1661 0.0119575
R75338 VSS.n8411 VSS.n1663 0.0119575
R75339 VSS.n8407 VSS.n1657 0.0119575
R75340 VSS.n8406 VSS.n1656 0.0119575
R75341 VSS.n8409 VSS.n8408 0.0119575
R75342 VSS.n8610 VSS.n1535 0.0119575
R75343 VSS.n1538 VSS.n1537 0.0119575
R75344 VSS.n8612 VSS.n1533 0.0119575
R75345 VSS.n8611 VSS.n1532 0.0119575
R75346 VSS.n8615 VSS.n8614 0.0119575
R75347 VSS.n8613 VSS.n1531 0.0119575
R75348 VSS.n8618 VSS.n8617 0.0119575
R75349 VSS.n8616 VSS.n1530 0.0119575
R75350 VSS.n8621 VSS.n8620 0.0119575
R75351 VSS.n8619 VSS.n1529 0.0119575
R75352 VSS.n8623 VSS.n1528 0.0119575
R75353 VSS.n8622 VSS.n1527 0.0119575
R75354 VSS.n8626 VSS.n8625 0.0119575
R75355 VSS.n8624 VSS.n1526 0.0119575
R75356 VSS.n8629 VSS.n8628 0.0119575
R75357 VSS.n8627 VSS.n1525 0.0119575
R75358 VSS.n8632 VSS.n8631 0.0119575
R75359 VSS.n8630 VSS.n1524 0.0119575
R75360 VSS.n1995 VSS.n1993 0.0119575
R75361 VSS.n1997 VSS.n1996 0.0119575
R75362 VSS.n8150 VSS.n1992 0.0119575
R75363 VSS.n1999 VSS.n1998 0.0119575
R75364 VSS.n8151 VSS.n1991 0.0119575
R75365 VSS.n2001 VSS.n2000 0.0119575
R75366 VSS.n8152 VSS.n1990 0.0119575
R75367 VSS.n2003 VSS.n2002 0.0119575
R75368 VSS.n8153 VSS.n1989 0.0119575
R75369 VSS.n2005 VSS.n2004 0.0119575
R75370 VSS.n8154 VSS.n1988 0.0119575
R75371 VSS.n2007 VSS.n2006 0.0119575
R75372 VSS.n8155 VSS.n1987 0.0119575
R75373 VSS.n2009 VSS.n2008 0.0119575
R75374 VSS.n8156 VSS.n1986 0.0119575
R75375 VSS.n2011 VSS.n2010 0.0119575
R75376 VSS.n8157 VSS.n1985 0.0119575
R75377 VSS.n2013 VSS.n2012 0.0119575
R75378 VSS.n8158 VSS.n1984 0.0119575
R75379 VSS.n2015 VSS.n2014 0.0119575
R75380 VSS.n8160 VSS.n1983 0.0119575
R75381 VSS.n8162 VSS.n8161 0.0119575
R75382 VSS.n1982 VSS.n1978 0.0119575
R75383 VSS.n8165 VSS.n1955 0.0119575
R75384 VSS.n8184 VSS.n8167 0.0119575
R75385 VSS.n1977 VSS.n1956 0.0119575
R75386 VSS.n8183 VSS.n8168 0.0119575
R75387 VSS.n1976 VSS.n1957 0.0119575
R75388 VSS.n8182 VSS.n8169 0.0119575
R75389 VSS.n1975 VSS.n1958 0.0119575
R75390 VSS.n8181 VSS.n8170 0.0119575
R75391 VSS.n1974 VSS.n1959 0.0119575
R75392 VSS.n8180 VSS.n8171 0.0119575
R75393 VSS.n1973 VSS.n1960 0.0119575
R75394 VSS.n8179 VSS.n8172 0.0119575
R75395 VSS.n1972 VSS.n1961 0.0119575
R75396 VSS.n8178 VSS.n8173 0.0119575
R75397 VSS.n1971 VSS.n1962 0.0119575
R75398 VSS.n8177 VSS.n8174 0.0119575
R75399 VSS.n1970 VSS.n1963 0.0119575
R75400 VSS.n8176 VSS.n8175 0.0119575
R75401 VSS.n1969 VSS.n1964 0.0119575
R75402 VSS.n8196 VSS.n8195 0.0119575
R75403 VSS.n1968 VSS.n1965 0.0119575
R75404 VSS.n8197 VSS.n1967 0.0119575
R75405 VSS.n8200 VSS.n8199 0.0119575
R75406 VSS.n4353 VSS.n4352 0.0119575
R75407 VSS.n4357 VSS.n4344 0.0119575
R75408 VSS.n4349 VSS.n4348 0.0119575
R75409 VSS.n4356 VSS.n4343 0.0119575
R75410 VSS.n4351 VSS.n4350 0.0119575
R75411 VSS.n5234 VSS.n4338 0.0119575
R75412 VSS.n5235 VSS.n4336 0.0119575
R75413 VSS.n5239 VSS.n5237 0.0119575
R75414 VSS.n5238 VSS.n4335 0.0119575
R75415 VSS.n5242 VSS.n5240 0.0119575
R75416 VSS.n5241 VSS.n4334 0.0119575
R75417 VSS.n5244 VSS.n5243 0.0119575
R75418 VSS.n5294 VSS.n5271 0.0119575
R75419 VSS.n5298 VSS.n5265 0.0119575
R75420 VSS.n5297 VSS.n5270 0.0119575
R75421 VSS.n5299 VSS.n5266 0.0119575
R75422 VSS.n5301 VSS.n5268 0.0119575
R75423 VSS.n5302 VSS.n5267 0.0119575
R75424 VSS.n3955 VSS.n3943 0.0119575
R75425 VSS.n6193 VSS.n3946 0.0119575
R75426 VSS.n3954 VSS.n3942 0.0119575
R75427 VSS.n6194 VSS.n3947 0.0119575
R75428 VSS.n3953 VSS.n3941 0.0119575
R75429 VSS.n6067 VSS.n6051 0.0119575
R75430 VSS.n6052 VSS.n6050 0.0119575
R75431 VSS.n6063 VSS.n6047 0.0119575
R75432 VSS.n6049 VSS.n6048 0.0119575
R75433 VSS.n6293 VSS.n3815 0.0119575
R75434 VSS.n3816 VSS.n3814 0.0119575
R75435 VSS.n6289 VSS.n3811 0.0119575
R75436 VSS.n3813 VSS.n3812 0.0119575
R75437 VSS.n3378 VSS.n3354 0.0119575
R75438 VSS.n3376 VSS.n3351 0.0119575
R75439 VSS.n3379 VSS.n3355 0.0119575
R75440 VSS.n3375 VSS.n3350 0.0119575
R75441 VSS.n3380 VSS.n3356 0.0119575
R75442 VSS.n3374 VSS.n3349 0.0119575
R75443 VSS.n3381 VSS.n3357 0.0119575
R75444 VSS.n3373 VSS.n3348 0.0119575
R75445 VSS.n3382 VSS.n3358 0.0119575
R75446 VSS.n3372 VSS.n3347 0.0119575
R75447 VSS.n3383 VSS.n3359 0.0119575
R75448 VSS.n3371 VSS.n3346 0.0119575
R75449 VSS.n3384 VSS.n3360 0.0119575
R75450 VSS.n3370 VSS.n3345 0.0119575
R75451 VSS.n3385 VSS.n3361 0.0119575
R75452 VSS.n3369 VSS.n3344 0.0119575
R75453 VSS.n3386 VSS.n3362 0.0119575
R75454 VSS.n3368 VSS.n3343 0.0119575
R75455 VSS.n3387 VSS.n3363 0.0119575
R75456 VSS.n3367 VSS.n3342 0.0119575
R75457 VSS.n3388 VSS.n3364 0.0119575
R75458 VSS.n3366 VSS.n3341 0.0119575
R75459 VSS.n6531 VSS.n3365 0.0119575
R75460 VSS.n6593 VSS.n3212 0.0119575
R75461 VSS.n3213 VSS.n3211 0.0119575
R75462 VSS.n6589 VSS.n3208 0.0119575
R75463 VSS.n3210 VSS.n3209 0.0119575
R75464 VSS.n5791 VSS.n5755 0.0119575
R75465 VSS.n5756 VSS.n5754 0.0119575
R75466 VSS.n5787 VSS.n5751 0.0119575
R75467 VSS.n5753 VSS.n5752 0.0119575
R75468 VSS.n2863 VSS.n2861 0.0119575
R75469 VSS.n6911 VSS.n2866 0.0119575
R75470 VSS.n2865 VSS.n2860 0.0119575
R75471 VSS.n6912 VSS.n2868 0.0119575
R75472 VSS.n2867 VSS.n2859 0.0119575
R75473 VSS.n6913 VSS.n2870 0.0119575
R75474 VSS.n2869 VSS.n2858 0.0119575
R75475 VSS.n6914 VSS.n2872 0.0119575
R75476 VSS.n2871 VSS.n2857 0.0119575
R75477 VSS.n6917 VSS.n6916 0.0119575
R75478 VSS.n6985 VSS.n2756 0.0119575
R75479 VSS.n2757 VSS.n2755 0.0119575
R75480 VSS.n6981 VSS.n2752 0.0119575
R75481 VSS.n2754 VSS.n2753 0.0119575
R75482 VSS.n1579 VSS.n1577 0.0119575
R75483 VSS.n1583 VSS.n1581 0.0119575
R75484 VSS.n1582 VSS.n1576 0.0119575
R75485 VSS.n1575 VSS.n1567 0.0119575
R75486 VSS.n1574 VSS.n1573 0.0119575
R75487 VSS.n1586 VSS.n1584 0.0119575
R75488 VSS.n1585 VSS.n1572 0.0119575
R75489 VSS.n8558 VSS.n1587 0.0119575
R75490 VSS.n8001 VSS.n8000 0.0119575
R75491 VSS.n8076 VSS.n2124 0.0119575
R75492 VSS.n2123 VSS.n2122 0.0119575
R75493 VSS.n2121 VSS.n2120 0.0119575
R75494 VSS.n2119 VSS.n2118 0.0119575
R75495 VSS.n2117 VSS.n2116 0.0119575
R75496 VSS.n2115 VSS.n2114 0.0119575
R75497 VSS.n2113 VSS.n2112 0.0119575
R75498 VSS.n2111 VSS.n2110 0.0119575
R75499 VSS.n8078 VSS.n2109 0.0119575
R75500 VSS.n2107 VSS.n2106 0.0119575
R75501 VSS.n2105 VSS.n2104 0.0119575
R75502 VSS.n2103 VSS.n2102 0.0119575
R75503 VSS.n2101 VSS.n2100 0.0119575
R75504 VSS.n2099 VSS.n2098 0.0119575
R75505 VSS.n2097 VSS.n2096 0.0119575
R75506 VSS.n2095 VSS.n2094 0.0119575
R75507 VSS.n2093 VSS.n2086 0.0119575
R75508 VSS.n2087 VSS.n2085 0.0119575
R75509 VSS.n8096 VSS.n2081 0.0119575
R75510 VSS.n8100 VSS.n2048 0.0119575
R75511 VSS.n8099 VSS.n2046 0.0119575
R75512 VSS.n2051 VSS.n2049 0.0119575
R75513 VSS.n2050 VSS.n2045 0.0119575
R75514 VSS.n2054 VSS.n2052 0.0119575
R75515 VSS.n2053 VSS.n2044 0.0119575
R75516 VSS.n2057 VSS.n2055 0.0119575
R75517 VSS.n2056 VSS.n2043 0.0119575
R75518 VSS.n2060 VSS.n2058 0.0119575
R75519 VSS.n2059 VSS.n2042 0.0119575
R75520 VSS.n2063 VSS.n2061 0.0119575
R75521 VSS.n2062 VSS.n2041 0.0119575
R75522 VSS.n2066 VSS.n2064 0.0119575
R75523 VSS.n2065 VSS.n2040 0.0119575
R75524 VSS.n2069 VSS.n2067 0.0119575
R75525 VSS.n2068 VSS.n2039 0.0119575
R75526 VSS.n2072 VSS.n2070 0.0119575
R75527 VSS.n2071 VSS.n2038 0.0119575
R75528 VSS.n2075 VSS.n2073 0.0119575
R75529 VSS.n2074 VSS.n2037 0.0119575
R75530 VSS.n2078 VSS.n2076 0.0119575
R75531 VSS.n2077 VSS.n2036 0.0119575
R75532 VSS.n8102 VSS.n2079 0.0119575
R75533 VSS.n1911 VSS.n1886 0.0119575
R75534 VSS.n1928 VSS.n1908 0.0119575
R75535 VSS.n1912 VSS.n1887 0.0119575
R75536 VSS.n1927 VSS.n1907 0.0119575
R75537 VSS.n1913 VSS.n1888 0.0119575
R75538 VSS.n1926 VSS.n1906 0.0119575
R75539 VSS.n1914 VSS.n1889 0.0119575
R75540 VSS.n1925 VSS.n1905 0.0119575
R75541 VSS.n1915 VSS.n1890 0.0119575
R75542 VSS.n1924 VSS.n1904 0.0119575
R75543 VSS.n1916 VSS.n1891 0.0119575
R75544 VSS.n1923 VSS.n1903 0.0119575
R75545 VSS.n1917 VSS.n1892 0.0119575
R75546 VSS.n1922 VSS.n1902 0.0119575
R75547 VSS.n1918 VSS.n1893 0.0119575
R75548 VSS.n1921 VSS.n1901 0.0119575
R75549 VSS.n1919 VSS.n1894 0.0119575
R75550 VSS.n1920 VSS.n1900 0.0119575
R75551 VSS.n8226 VSS.n1895 0.0119575
R75552 VSS.n8225 VSS.n1899 0.0119575
R75553 VSS.n8227 VSS.n1896 0.0119575
R75554 VSS.n8229 VSS.n1898 0.0119575
R75555 VSS.n8230 VSS.n1897 0.0119575
R75556 VSS.n2340 VSS.n2337 0.0119575
R75557 VSS.n2363 VSS.n2336 0.0119575
R75558 VSS.n2362 VSS.n2341 0.0119575
R75559 VSS.n5236 VSS.n5235 0.0119575
R75560 VSS.n5237 VSS.n4336 0.0119575
R75561 VSS.n5239 VSS.n5238 0.0119575
R75562 VSS.n5240 VSS.n4335 0.0119575
R75563 VSS.n5242 VSS.n5241 0.0119575
R75564 VSS.n5243 VSS.n4334 0.0119575
R75565 VSS.n5294 VSS.n5264 0.0119575
R75566 VSS.n5271 VSS.n5265 0.0119575
R75567 VSS.n5298 VSS.n5297 0.0119575
R75568 VSS.n5270 VSS.n5266 0.0119575
R75569 VSS.n5299 VSS.n5268 0.0119575
R75570 VSS.n5302 VSS.n5301 0.0119575
R75571 VSS.n3955 VSS.n3945 0.0119575
R75572 VSS.n6193 VSS.n3943 0.0119575
R75573 VSS.n3954 VSS.n3946 0.0119575
R75574 VSS.n6194 VSS.n3942 0.0119575
R75575 VSS.n3953 VSS.n3947 0.0119575
R75576 VSS.n3378 VSS.n3352 0.0119575
R75577 VSS.n3376 VSS.n3354 0.0119575
R75578 VSS.n3379 VSS.n3351 0.0119575
R75579 VSS.n3375 VSS.n3355 0.0119575
R75580 VSS.n3380 VSS.n3350 0.0119575
R75581 VSS.n3374 VSS.n3356 0.0119575
R75582 VSS.n3381 VSS.n3349 0.0119575
R75583 VSS.n3373 VSS.n3357 0.0119575
R75584 VSS.n3382 VSS.n3348 0.0119575
R75585 VSS.n3372 VSS.n3358 0.0119575
R75586 VSS.n3383 VSS.n3347 0.0119575
R75587 VSS.n3371 VSS.n3359 0.0119575
R75588 VSS.n3384 VSS.n3346 0.0119575
R75589 VSS.n3370 VSS.n3360 0.0119575
R75590 VSS.n3385 VSS.n3345 0.0119575
R75591 VSS.n3369 VSS.n3361 0.0119575
R75592 VSS.n3386 VSS.n3344 0.0119575
R75593 VSS.n3368 VSS.n3362 0.0119575
R75594 VSS.n3387 VSS.n3343 0.0119575
R75595 VSS.n3367 VSS.n3363 0.0119575
R75596 VSS.n3388 VSS.n3342 0.0119575
R75597 VSS.n3366 VSS.n3364 0.0119575
R75598 VSS.n3365 VSS.n3341 0.0119575
R75599 VSS.n2864 VSS.n2863 0.0119575
R75600 VSS.n6911 VSS.n2861 0.0119575
R75601 VSS.n2866 VSS.n2865 0.0119575
R75602 VSS.n6912 VSS.n2860 0.0119575
R75603 VSS.n2868 VSS.n2867 0.0119575
R75604 VSS.n6913 VSS.n2859 0.0119575
R75605 VSS.n2870 VSS.n2869 0.0119575
R75606 VSS.n6914 VSS.n2858 0.0119575
R75607 VSS.n2872 VSS.n2871 0.0119575
R75608 VSS.n6916 VSS.n2857 0.0119575
R75609 VSS.n1580 VSS.n1579 0.0119575
R75610 VSS.n1581 VSS.n1577 0.0119575
R75611 VSS.n1583 VSS.n1582 0.0119575
R75612 VSS.n1576 VSS.n1575 0.0119575
R75613 VSS.n1573 VSS.n1563 0.0119575
R75614 VSS.n1584 VSS.n1574 0.0119575
R75615 VSS.n1586 VSS.n1585 0.0119575
R75616 VSS.n1587 VSS.n1572 0.0119575
R75617 VSS.n8000 VSS.n1595 0.0119575
R75618 VSS.n8077 VSS.n8076 0.0119575
R75619 VSS.n2124 VSS.n2123 0.0119575
R75620 VSS.n2122 VSS.n2121 0.0119575
R75621 VSS.n2120 VSS.n2119 0.0119575
R75622 VSS.n2118 VSS.n2117 0.0119575
R75623 VSS.n2116 VSS.n2115 0.0119575
R75624 VSS.n2114 VSS.n2113 0.0119575
R75625 VSS.n2112 VSS.n2111 0.0119575
R75626 VSS.n2110 VSS.n2109 0.0119575
R75627 VSS.n2108 VSS.n2107 0.0119575
R75628 VSS.n2106 VSS.n2105 0.0119575
R75629 VSS.n2104 VSS.n2103 0.0119575
R75630 VSS.n2102 VSS.n2101 0.0119575
R75631 VSS.n2100 VSS.n2099 0.0119575
R75632 VSS.n2098 VSS.n2097 0.0119575
R75633 VSS.n2096 VSS.n2095 0.0119575
R75634 VSS.n2094 VSS.n2093 0.0119575
R75635 VSS.n8097 VSS.n2048 0.0119575
R75636 VSS.n8100 VSS.n8099 0.0119575
R75637 VSS.n2049 VSS.n2046 0.0119575
R75638 VSS.n2051 VSS.n2050 0.0119575
R75639 VSS.n2052 VSS.n2045 0.0119575
R75640 VSS.n2054 VSS.n2053 0.0119575
R75641 VSS.n2055 VSS.n2044 0.0119575
R75642 VSS.n2057 VSS.n2056 0.0119575
R75643 VSS.n2058 VSS.n2043 0.0119575
R75644 VSS.n2060 VSS.n2059 0.0119575
R75645 VSS.n2061 VSS.n2042 0.0119575
R75646 VSS.n2063 VSS.n2062 0.0119575
R75647 VSS.n2064 VSS.n2041 0.0119575
R75648 VSS.n2066 VSS.n2065 0.0119575
R75649 VSS.n2067 VSS.n2040 0.0119575
R75650 VSS.n2069 VSS.n2068 0.0119575
R75651 VSS.n2070 VSS.n2039 0.0119575
R75652 VSS.n2072 VSS.n2071 0.0119575
R75653 VSS.n2073 VSS.n2038 0.0119575
R75654 VSS.n2075 VSS.n2074 0.0119575
R75655 VSS.n2076 VSS.n2037 0.0119575
R75656 VSS.n2078 VSS.n2077 0.0119575
R75657 VSS.n2079 VSS.n2036 0.0119575
R75658 VSS.n1909 VSS.n1886 0.0119575
R75659 VSS.n1928 VSS.n1911 0.0119575
R75660 VSS.n1908 VSS.n1887 0.0119575
R75661 VSS.n1927 VSS.n1912 0.0119575
R75662 VSS.n1907 VSS.n1888 0.0119575
R75663 VSS.n1926 VSS.n1913 0.0119575
R75664 VSS.n1906 VSS.n1889 0.0119575
R75665 VSS.n1925 VSS.n1914 0.0119575
R75666 VSS.n1905 VSS.n1890 0.0119575
R75667 VSS.n1924 VSS.n1915 0.0119575
R75668 VSS.n1904 VSS.n1891 0.0119575
R75669 VSS.n1923 VSS.n1916 0.0119575
R75670 VSS.n1903 VSS.n1892 0.0119575
R75671 VSS.n1922 VSS.n1917 0.0119575
R75672 VSS.n1902 VSS.n1893 0.0119575
R75673 VSS.n1921 VSS.n1918 0.0119575
R75674 VSS.n1901 VSS.n1894 0.0119575
R75675 VSS.n1920 VSS.n1919 0.0119575
R75676 VSS.n1900 VSS.n1895 0.0119575
R75677 VSS.n8226 VSS.n8225 0.0119575
R75678 VSS.n1899 VSS.n1896 0.0119575
R75679 VSS.n8227 VSS.n1898 0.0119575
R75680 VSS.n8230 VSS.n8229 0.0119575
R75681 VSS.n4602 VSS.n4601 0.0119575
R75682 VSS.n4606 VSS.n4593 0.0119575
R75683 VSS.n4598 VSS.n4597 0.0119575
R75684 VSS.n4605 VSS.n4592 0.0119575
R75685 VSS.n4600 VSS.n4599 0.0119575
R75686 VSS.n4721 VSS.n4587 0.0119575
R75687 VSS.n4735 VSS.n4734 0.0119575
R75688 VSS.n4739 VSS.n4723 0.0119575
R75689 VSS.n4738 VSS.n4733 0.0119575
R75690 VSS.n4741 VSS.n4724 0.0119575
R75691 VSS.n4740 VSS.n4732 0.0119575
R75692 VSS.n4761 VSS.n4725 0.0119575
R75693 VSS.n3873 VSS.n3872 0.0119575
R75694 VSS.n6242 VSS.n6240 0.0119575
R75695 VSS.n6241 VSS.n3871 0.0119575
R75696 VSS.n6245 VSS.n6243 0.0119575
R75697 VSS.n6244 VSS.n3870 0.0119575
R75698 VSS.n6247 VSS.n6246 0.0119575
R75699 VSS.n3843 VSS.n3841 0.0119575
R75700 VSS.n3847 VSS.n3845 0.0119575
R75701 VSS.n3846 VSS.n3840 0.0119575
R75702 VSS.n3850 VSS.n3848 0.0119575
R75703 VSS.n3849 VSS.n3839 0.0119575
R75704 VSS.n6558 VSS.n3249 0.0119575
R75705 VSS.n3248 VSS.n3245 0.0119575
R75706 VSS.n6559 VSS.n3251 0.0119575
R75707 VSS.n3250 VSS.n3244 0.0119575
R75708 VSS.n6560 VSS.n3253 0.0119575
R75709 VSS.n3252 VSS.n3243 0.0119575
R75710 VSS.n6561 VSS.n3255 0.0119575
R75711 VSS.n3254 VSS.n3242 0.0119575
R75712 VSS.n6562 VSS.n3257 0.0119575
R75713 VSS.n3256 VSS.n3241 0.0119575
R75714 VSS.n6563 VSS.n3259 0.0119575
R75715 VSS.n3258 VSS.n3240 0.0119575
R75716 VSS.n6564 VSS.n3261 0.0119575
R75717 VSS.n3260 VSS.n3239 0.0119575
R75718 VSS.n6565 VSS.n3263 0.0119575
R75719 VSS.n3262 VSS.n3238 0.0119575
R75720 VSS.n6566 VSS.n3265 0.0119575
R75721 VSS.n3264 VSS.n3237 0.0119575
R75722 VSS.n6567 VSS.n3267 0.0119575
R75723 VSS.n3266 VSS.n3236 0.0119575
R75724 VSS.n6571 VSS.n6569 0.0119575
R75725 VSS.n6570 VSS.n3235 0.0119575
R75726 VSS.n6573 VSS.n3231 0.0119575
R75727 VSS.n2806 VSS.n2804 0.0119575
R75728 VSS.n6957 VSS.n2809 0.0119575
R75729 VSS.n2808 VSS.n2803 0.0119575
R75730 VSS.n6958 VSS.n2811 0.0119575
R75731 VSS.n2810 VSS.n2802 0.0119575
R75732 VSS.n6959 VSS.n2813 0.0119575
R75733 VSS.n2812 VSS.n2801 0.0119575
R75734 VSS.n6963 VSS.n6961 0.0119575
R75735 VSS.n6962 VSS.n2800 0.0119575
R75736 VSS.n6965 VSS.n2796 0.0119575
R75737 VSS.n8292 VSS.n8285 0.0119575
R75738 VSS.n8288 VSS.n1708 0.0119575
R75739 VSS.n8291 VSS.n8284 0.0119575
R75740 VSS.n8289 VSS.n1709 0.0119575
R75741 VSS.n8290 VSS.n8283 0.0119575
R75742 VSS.n8296 VSS.n1710 0.0119575
R75743 VSS.n8295 VSS.n8282 0.0119575
R75744 VSS.n8297 VSS.n1711 0.0119575
R75745 VSS.n8299 VSS.n8280 0.0119575
R75746 VSS.n8300 VSS.n8279 0.0119575
R75747 VSS.n1729 VSS.n1712 0.0119575
R75748 VSS.n1728 VSS.n1726 0.0119575
R75749 VSS.n2232 VSS.n1731 0.0119575
R75750 VSS.n1730 VSS.n1725 0.0119575
R75751 VSS.n2233 VSS.n1733 0.0119575
R75752 VSS.n1732 VSS.n1724 0.0119575
R75753 VSS.n2234 VSS.n1735 0.0119575
R75754 VSS.n1734 VSS.n1723 0.0119575
R75755 VSS.n2235 VSS.n1737 0.0119575
R75756 VSS.n1736 VSS.n1722 0.0119575
R75757 VSS.n2236 VSS.n1739 0.0119575
R75758 VSS.n1738 VSS.n1721 0.0119575
R75759 VSS.n2237 VSS.n1741 0.0119575
R75760 VSS.n1740 VSS.n1720 0.0119575
R75761 VSS.n2238 VSS.n1743 0.0119575
R75762 VSS.n1742 VSS.n1719 0.0119575
R75763 VSS.n2239 VSS.n1745 0.0119575
R75764 VSS.n1744 VSS.n1718 0.0119575
R75765 VSS.n2240 VSS.n1747 0.0119575
R75766 VSS.n1746 VSS.n1717 0.0119575
R75767 VSS.n2241 VSS.n1749 0.0119575
R75768 VSS.n1748 VSS.n1716 0.0119575
R75769 VSS.n8276 VSS.n1750 0.0119575
R75770 VSS.n1768 VSS.n1751 0.0119575
R75771 VSS.n1767 VSS.n1765 0.0119575
R75772 VSS.n7901 VSS.n1770 0.0119575
R75773 VSS.n1769 VSS.n1764 0.0119575
R75774 VSS.n7902 VSS.n1772 0.0119575
R75775 VSS.n1771 VSS.n1763 0.0119575
R75776 VSS.n7903 VSS.n1774 0.0119575
R75777 VSS.n1773 VSS.n1762 0.0119575
R75778 VSS.n7904 VSS.n1776 0.0119575
R75779 VSS.n1775 VSS.n1761 0.0119575
R75780 VSS.n7905 VSS.n1778 0.0119575
R75781 VSS.n1777 VSS.n1760 0.0119575
R75782 VSS.n7906 VSS.n1780 0.0119575
R75783 VSS.n1779 VSS.n1759 0.0119575
R75784 VSS.n7907 VSS.n1782 0.0119575
R75785 VSS.n1781 VSS.n1758 0.0119575
R75786 VSS.n7908 VSS.n1784 0.0119575
R75787 VSS.n1783 VSS.n1757 0.0119575
R75788 VSS.n7909 VSS.n1786 0.0119575
R75789 VSS.n1785 VSS.n1756 0.0119575
R75790 VSS.n7910 VSS.n1788 0.0119575
R75791 VSS.n1787 VSS.n1755 0.0119575
R75792 VSS.n8273 VSS.n1789 0.0119575
R75793 VSS.n1807 VSS.n1790 0.0119575
R75794 VSS.n1806 VSS.n1804 0.0119575
R75795 VSS.n8258 VSS.n1809 0.0119575
R75796 VSS.n1808 VSS.n1803 0.0119575
R75797 VSS.n8259 VSS.n1811 0.0119575
R75798 VSS.n1810 VSS.n1802 0.0119575
R75799 VSS.n8260 VSS.n1813 0.0119575
R75800 VSS.n1812 VSS.n1801 0.0119575
R75801 VSS.n8261 VSS.n1815 0.0119575
R75802 VSS.n1814 VSS.n1800 0.0119575
R75803 VSS.n8262 VSS.n1817 0.0119575
R75804 VSS.n1816 VSS.n1799 0.0119575
R75805 VSS.n8263 VSS.n1819 0.0119575
R75806 VSS.n1818 VSS.n1798 0.0119575
R75807 VSS.n8264 VSS.n1821 0.0119575
R75808 VSS.n1820 VSS.n1797 0.0119575
R75809 VSS.n8265 VSS.n1823 0.0119575
R75810 VSS.n1822 VSS.n1796 0.0119575
R75811 VSS.n8266 VSS.n1825 0.0119575
R75812 VSS.n1824 VSS.n1795 0.0119575
R75813 VSS.n8267 VSS.n1827 0.0119575
R75814 VSS.n1826 VSS.n1794 0.0119575
R75815 VSS.n8270 VSS.n8269 0.0119575
R75816 VSS.n4734 VSS.n4722 0.0119575
R75817 VSS.n4735 VSS.n4723 0.0119575
R75818 VSS.n4739 VSS.n4738 0.0119575
R75819 VSS.n4733 VSS.n4724 0.0119575
R75820 VSS.n4741 VSS.n4740 0.0119575
R75821 VSS.n4732 VSS.n4725 0.0119575
R75822 VSS.n3872 VSS.n3862 0.0119575
R75823 VSS.n6240 VSS.n3873 0.0119575
R75824 VSS.n6242 VSS.n6241 0.0119575
R75825 VSS.n6243 VSS.n3871 0.0119575
R75826 VSS.n6245 VSS.n6244 0.0119575
R75827 VSS.n6246 VSS.n3870 0.0119575
R75828 VSS.n3844 VSS.n3843 0.0119575
R75829 VSS.n3845 VSS.n3841 0.0119575
R75830 VSS.n3847 VSS.n3846 0.0119575
R75831 VSS.n3848 VSS.n3840 0.0119575
R75832 VSS.n3850 VSS.n3849 0.0119575
R75833 VSS.n6558 VSS.n3246 0.0119575
R75834 VSS.n3249 VSS.n3248 0.0119575
R75835 VSS.n6559 VSS.n3245 0.0119575
R75836 VSS.n3251 VSS.n3250 0.0119575
R75837 VSS.n6560 VSS.n3244 0.0119575
R75838 VSS.n3253 VSS.n3252 0.0119575
R75839 VSS.n6561 VSS.n3243 0.0119575
R75840 VSS.n3255 VSS.n3254 0.0119575
R75841 VSS.n6562 VSS.n3242 0.0119575
R75842 VSS.n3257 VSS.n3256 0.0119575
R75843 VSS.n6563 VSS.n3241 0.0119575
R75844 VSS.n3259 VSS.n3258 0.0119575
R75845 VSS.n6564 VSS.n3240 0.0119575
R75846 VSS.n3261 VSS.n3260 0.0119575
R75847 VSS.n6565 VSS.n3239 0.0119575
R75848 VSS.n3263 VSS.n3262 0.0119575
R75849 VSS.n6566 VSS.n3238 0.0119575
R75850 VSS.n3265 VSS.n3264 0.0119575
R75851 VSS.n6567 VSS.n3237 0.0119575
R75852 VSS.n3267 VSS.n3266 0.0119575
R75853 VSS.n6569 VSS.n3236 0.0119575
R75854 VSS.n6571 VSS.n6570 0.0119575
R75855 VSS.n3235 VSS.n3231 0.0119575
R75856 VSS.n2807 VSS.n2806 0.0119575
R75857 VSS.n6957 VSS.n2804 0.0119575
R75858 VSS.n2809 VSS.n2808 0.0119575
R75859 VSS.n6958 VSS.n2803 0.0119575
R75860 VSS.n2811 VSS.n2810 0.0119575
R75861 VSS.n6959 VSS.n2802 0.0119575
R75862 VSS.n2813 VSS.n2812 0.0119575
R75863 VSS.n6961 VSS.n2801 0.0119575
R75864 VSS.n6963 VSS.n6962 0.0119575
R75865 VSS.n2800 VSS.n2796 0.0119575
R75866 VSS.n8292 VSS.n1707 0.0119575
R75867 VSS.n8285 VSS.n1708 0.0119575
R75868 VSS.n8291 VSS.n8288 0.0119575
R75869 VSS.n8284 VSS.n1709 0.0119575
R75870 VSS.n8290 VSS.n8289 0.0119575
R75871 VSS.n8283 VSS.n1710 0.0119575
R75872 VSS.n8296 VSS.n8295 0.0119575
R75873 VSS.n8282 VSS.n1711 0.0119575
R75874 VSS.n8297 VSS.n8280 0.0119575
R75875 VSS.n8300 VSS.n8299 0.0119575
R75876 VSS.n8278 VSS.n1712 0.0119575
R75877 VSS.n1729 VSS.n1728 0.0119575
R75878 VSS.n2232 VSS.n1726 0.0119575
R75879 VSS.n1731 VSS.n1730 0.0119575
R75880 VSS.n2233 VSS.n1725 0.0119575
R75881 VSS.n1733 VSS.n1732 0.0119575
R75882 VSS.n2234 VSS.n1724 0.0119575
R75883 VSS.n1735 VSS.n1734 0.0119575
R75884 VSS.n2235 VSS.n1723 0.0119575
R75885 VSS.n1737 VSS.n1736 0.0119575
R75886 VSS.n2236 VSS.n1722 0.0119575
R75887 VSS.n1739 VSS.n1738 0.0119575
R75888 VSS.n2237 VSS.n1721 0.0119575
R75889 VSS.n1741 VSS.n1740 0.0119575
R75890 VSS.n2238 VSS.n1720 0.0119575
R75891 VSS.n1743 VSS.n1742 0.0119575
R75892 VSS.n2239 VSS.n1719 0.0119575
R75893 VSS.n1745 VSS.n1744 0.0119575
R75894 VSS.n2240 VSS.n1718 0.0119575
R75895 VSS.n1747 VSS.n1746 0.0119575
R75896 VSS.n2241 VSS.n1717 0.0119575
R75897 VSS.n1749 VSS.n1748 0.0119575
R75898 VSS.n1750 VSS.n1716 0.0119575
R75899 VSS.n8275 VSS.n1751 0.0119575
R75900 VSS.n1768 VSS.n1767 0.0119575
R75901 VSS.n7901 VSS.n1765 0.0119575
R75902 VSS.n1770 VSS.n1769 0.0119575
R75903 VSS.n7902 VSS.n1764 0.0119575
R75904 VSS.n1772 VSS.n1771 0.0119575
R75905 VSS.n7903 VSS.n1763 0.0119575
R75906 VSS.n1774 VSS.n1773 0.0119575
R75907 VSS.n7904 VSS.n1762 0.0119575
R75908 VSS.n1776 VSS.n1775 0.0119575
R75909 VSS.n7905 VSS.n1761 0.0119575
R75910 VSS.n1778 VSS.n1777 0.0119575
R75911 VSS.n7906 VSS.n1760 0.0119575
R75912 VSS.n1780 VSS.n1779 0.0119575
R75913 VSS.n7907 VSS.n1759 0.0119575
R75914 VSS.n1782 VSS.n1781 0.0119575
R75915 VSS.n7908 VSS.n1758 0.0119575
R75916 VSS.n1784 VSS.n1783 0.0119575
R75917 VSS.n7909 VSS.n1757 0.0119575
R75918 VSS.n1786 VSS.n1785 0.0119575
R75919 VSS.n7910 VSS.n1756 0.0119575
R75920 VSS.n1788 VSS.n1787 0.0119575
R75921 VSS.n1789 VSS.n1755 0.0119575
R75922 VSS.n8272 VSS.n1790 0.0119575
R75923 VSS.n1807 VSS.n1806 0.0119575
R75924 VSS.n8258 VSS.n1804 0.0119575
R75925 VSS.n1809 VSS.n1808 0.0119575
R75926 VSS.n8259 VSS.n1803 0.0119575
R75927 VSS.n1811 VSS.n1810 0.0119575
R75928 VSS.n8260 VSS.n1802 0.0119575
R75929 VSS.n1813 VSS.n1812 0.0119575
R75930 VSS.n8261 VSS.n1801 0.0119575
R75931 VSS.n1815 VSS.n1814 0.0119575
R75932 VSS.n8262 VSS.n1800 0.0119575
R75933 VSS.n1817 VSS.n1816 0.0119575
R75934 VSS.n8263 VSS.n1799 0.0119575
R75935 VSS.n1819 VSS.n1818 0.0119575
R75936 VSS.n8264 VSS.n1798 0.0119575
R75937 VSS.n1821 VSS.n1820 0.0119575
R75938 VSS.n8265 VSS.n1797 0.0119575
R75939 VSS.n1823 VSS.n1822 0.0119575
R75940 VSS.n8266 VSS.n1796 0.0119575
R75941 VSS.n1825 VSS.n1824 0.0119575
R75942 VSS.n8267 VSS.n1795 0.0119575
R75943 VSS.n1827 VSS.n1826 0.0119575
R75944 VSS.n8269 VSS.n1794 0.0119575
R75945 VSS.n4606 VSS.n4596 0.0119575
R75946 VSS.n4597 VSS.n4593 0.0119575
R75947 VSS.n4605 VSS.n4598 0.0119575
R75948 VSS.n4599 VSS.n4592 0.0119575
R75949 VSS.n4600 VSS.n4587 0.0119575
R75950 VSS.n4601 VSS.n4591 0.0119575
R75951 VSS.n4680 VSS.n4624 0.0119575
R75952 VSS.n4629 VSS.n4621 0.0119575
R75953 VSS.n4679 VSS.n4625 0.0119575
R75954 VSS.n4630 VSS.n4620 0.0119575
R75955 VSS.n4678 VSS.n4626 0.0119575
R75956 VSS.n4676 VSS.n4618 0.0119575
R75957 VSS.n4357 VSS.n4347 0.0119575
R75958 VSS.n4348 VSS.n4344 0.0119575
R75959 VSS.n4356 VSS.n4349 0.0119575
R75960 VSS.n4350 VSS.n4343 0.0119575
R75961 VSS.n4351 VSS.n4338 0.0119575
R75962 VSS.n4352 VSS.n4342 0.0119575
R75963 VSS.n4400 VSS.n4387 0.0119575
R75964 VSS.n4392 VSS.n4384 0.0119575
R75965 VSS.n4399 VSS.n4388 0.0119575
R75966 VSS.n4393 VSS.n4383 0.0119575
R75967 VSS.n4398 VSS.n4389 0.0119575
R75968 VSS.n4396 VSS.n4381 0.0119575
R75969 VSS.n9893 VSS.n32 0.0119575
R75970 VSS.n42 VSS.n40 0.0119575
R75971 VSS.n45 VSS.n43 0.0119575
R75972 VSS.n44 VSS.n39 0.0119575
R75973 VSS.n9891 VSS.n9890 0.0119575
R75974 VSS.n37 VSS.n36 0.0119575
R75975 VSS.n88 VSS.n75 0.0119575
R75976 VSS.n80 VSS.n72 0.0119575
R75977 VSS.n87 VSS.n76 0.0119575
R75978 VSS.n81 VSS.n71 0.0119575
R75979 VSS.n86 VSS.n77 0.0119575
R75980 VSS.n84 VSS.n69 0.0119575
R75981 VSS.n142 VSS.n131 0.0119575
R75982 VSS.n145 VSS.n134 0.0119575
R75983 VSS.n9830 VSS.n138 0.0119575
R75984 VSS.n144 VSS.n133 0.0119575
R75985 VSS.n9831 VSS.n139 0.0119575
R75986 VSS.n143 VSS.n132 0.0119575
R75987 VSS.n9798 VSS.n184 0.0119575
R75988 VSS.n9802 VSS.n9800 0.0119575
R75989 VSS.n9801 VSS.n183 0.0119575
R75990 VSS.n9805 VSS.n9803 0.0119575
R75991 VSS.n9804 VSS.n182 0.0119575
R75992 VSS.n9807 VSS.n9806 0.0119575
R75993 VSS.n5474 VSS.n5434 0.0119575
R75994 VSS.n5480 VSS.n5477 0.0119575
R75995 VSS.n5476 VSS.n5433 0.0119575
R75996 VSS.n5481 VSS.n5479 0.0119575
R75997 VSS.n5478 VSS.n5432 0.0119575
R75998 VSS.n5484 VSS.n5483 0.0119575
R75999 VSS.n414 VSS.n412 0.0119575
R76000 VSS.n423 VSS.n417 0.0119575
R76001 VSS.n416 VSS.n411 0.0119575
R76002 VSS.n424 VSS.n419 0.0119575
R76003 VSS.n418 VSS.n410 0.0119575
R76004 VSS.n461 VSS.n444 0.0119575
R76005 VSS.n460 VSS.n458 0.0119575
R76006 VSS.n6374 VSS.n463 0.0119575
R76007 VSS.n462 VSS.n457 0.0119575
R76008 VSS.n6375 VSS.n465 0.0119575
R76009 VSS.n464 VSS.n456 0.0119575
R76010 VSS.n6376 VSS.n467 0.0119575
R76011 VSS.n466 VSS.n455 0.0119575
R76012 VSS.n6377 VSS.n469 0.0119575
R76013 VSS.n468 VSS.n454 0.0119575
R76014 VSS.n6378 VSS.n471 0.0119575
R76015 VSS.n470 VSS.n453 0.0119575
R76016 VSS.n6379 VSS.n473 0.0119575
R76017 VSS.n472 VSS.n452 0.0119575
R76018 VSS.n6380 VSS.n475 0.0119575
R76019 VSS.n474 VSS.n451 0.0119575
R76020 VSS.n6381 VSS.n477 0.0119575
R76021 VSS.n476 VSS.n450 0.0119575
R76022 VSS.n6382 VSS.n479 0.0119575
R76023 VSS.n478 VSS.n449 0.0119575
R76024 VSS.n6383 VSS.n481 0.0119575
R76025 VSS.n480 VSS.n448 0.0119575
R76026 VSS.n9594 VSS.n482 0.0119575
R76027 VSS.n509 VSS.n501 0.0119575
R76028 VSS.n512 VSS.n511 0.0119575
R76029 VSS.n523 VSS.n508 0.0119575
R76030 VSS.n514 VSS.n513 0.0119575
R76031 VSS.n522 VSS.n507 0.0119575
R76032 VSS.n516 VSS.n515 0.0119575
R76033 VSS.n521 VSS.n506 0.0119575
R76034 VSS.n518 VSS.n517 0.0119575
R76035 VSS.n520 VSS.n505 0.0119575
R76036 VSS.n9581 VSS.n519 0.0119575
R76037 VSS.n547 VSS.n539 0.0119575
R76038 VSS.n550 VSS.n549 0.0119575
R76039 VSS.n561 VSS.n546 0.0119575
R76040 VSS.n552 VSS.n551 0.0119575
R76041 VSS.n560 VSS.n545 0.0119575
R76042 VSS.n554 VSS.n553 0.0119575
R76043 VSS.n559 VSS.n544 0.0119575
R76044 VSS.n556 VSS.n555 0.0119575
R76045 VSS.n558 VSS.n543 0.0119575
R76046 VSS.n9568 VSS.n557 0.0119575
R76047 VSS.n580 VSS.n563 0.0119575
R76048 VSS.n579 VSS.n577 0.0119575
R76049 VSS.n8926 VSS.n582 0.0119575
R76050 VSS.n581 VSS.n576 0.0119575
R76051 VSS.n8927 VSS.n584 0.0119575
R76052 VSS.n583 VSS.n575 0.0119575
R76053 VSS.n8928 VSS.n586 0.0119575
R76054 VSS.n585 VSS.n574 0.0119575
R76055 VSS.n8929 VSS.n588 0.0119575
R76056 VSS.n587 VSS.n573 0.0119575
R76057 VSS.n8930 VSS.n590 0.0119575
R76058 VSS.n589 VSS.n572 0.0119575
R76059 VSS.n8931 VSS.n592 0.0119575
R76060 VSS.n591 VSS.n571 0.0119575
R76061 VSS.n8932 VSS.n594 0.0119575
R76062 VSS.n593 VSS.n570 0.0119575
R76063 VSS.n8933 VSS.n596 0.0119575
R76064 VSS.n595 VSS.n569 0.0119575
R76065 VSS.n8934 VSS.n598 0.0119575
R76066 VSS.n597 VSS.n568 0.0119575
R76067 VSS.n8935 VSS.n600 0.0119575
R76068 VSS.n599 VSS.n567 0.0119575
R76069 VSS.n9565 VSS.n601 0.0119575
R76070 VSS.n618 VSS.n602 0.0119575
R76071 VSS.n617 VSS.n615 0.0119575
R76072 VSS.n9473 VSS.n620 0.0119575
R76073 VSS.n619 VSS.n614 0.0119575
R76074 VSS.n9474 VSS.n622 0.0119575
R76075 VSS.n621 VSS.n613 0.0119575
R76076 VSS.n9475 VSS.n624 0.0119575
R76077 VSS.n623 VSS.n612 0.0119575
R76078 VSS.n9476 VSS.n626 0.0119575
R76079 VSS.n625 VSS.n611 0.0119575
R76080 VSS.n9477 VSS.n628 0.0119575
R76081 VSS.n627 VSS.n610 0.0119575
R76082 VSS.n9478 VSS.n630 0.0119575
R76083 VSS.n629 VSS.n609 0.0119575
R76084 VSS.n9479 VSS.n632 0.0119575
R76085 VSS.n631 VSS.n608 0.0119575
R76086 VSS.n9480 VSS.n634 0.0119575
R76087 VSS.n633 VSS.n607 0.0119575
R76088 VSS.n9481 VSS.n636 0.0119575
R76089 VSS.n635 VSS.n606 0.0119575
R76090 VSS.n9482 VSS.n638 0.0119575
R76091 VSS.n637 VSS.n605 0.0119575
R76092 VSS.n9562 VSS.n639 0.0119575
R76093 VSS.n657 VSS.n640 0.0119575
R76094 VSS.n656 VSS.n654 0.0119575
R76095 VSS.n9547 VSS.n659 0.0119575
R76096 VSS.n658 VSS.n653 0.0119575
R76097 VSS.n9548 VSS.n661 0.0119575
R76098 VSS.n660 VSS.n652 0.0119575
R76099 VSS.n9549 VSS.n663 0.0119575
R76100 VSS.n662 VSS.n651 0.0119575
R76101 VSS.n9550 VSS.n665 0.0119575
R76102 VSS.n664 VSS.n650 0.0119575
R76103 VSS.n9551 VSS.n667 0.0119575
R76104 VSS.n666 VSS.n649 0.0119575
R76105 VSS.n9552 VSS.n669 0.0119575
R76106 VSS.n668 VSS.n648 0.0119575
R76107 VSS.n9553 VSS.n671 0.0119575
R76108 VSS.n670 VSS.n647 0.0119575
R76109 VSS.n9554 VSS.n673 0.0119575
R76110 VSS.n672 VSS.n646 0.0119575
R76111 VSS.n9555 VSS.n675 0.0119575
R76112 VSS.n674 VSS.n645 0.0119575
R76113 VSS.n9556 VSS.n677 0.0119575
R76114 VSS.n676 VSS.n644 0.0119575
R76115 VSS.n9559 VSS.n9558 0.0119575
R76116 VSS.n145 VSS.n137 0.0119575
R76117 VSS.n9830 VSS.n134 0.0119575
R76118 VSS.n144 VSS.n138 0.0119575
R76119 VSS.n9831 VSS.n133 0.0119575
R76120 VSS.n143 VSS.n139 0.0119575
R76121 VSS.n9799 VSS.n9798 0.0119575
R76122 VSS.n9800 VSS.n184 0.0119575
R76123 VSS.n9802 VSS.n9801 0.0119575
R76124 VSS.n9803 VSS.n183 0.0119575
R76125 VSS.n9805 VSS.n9804 0.0119575
R76126 VSS.n9806 VSS.n182 0.0119575
R76127 VSS.n5475 VSS.n5474 0.0119575
R76128 VSS.n5480 VSS.n5434 0.0119575
R76129 VSS.n5477 VSS.n5476 0.0119575
R76130 VSS.n5481 VSS.n5433 0.0119575
R76131 VSS.n5479 VSS.n5478 0.0119575
R76132 VSS.n5483 VSS.n5432 0.0119575
R76133 VSS.n415 VSS.n414 0.0119575
R76134 VSS.n423 VSS.n412 0.0119575
R76135 VSS.n417 VSS.n416 0.0119575
R76136 VSS.n424 VSS.n411 0.0119575
R76137 VSS.n419 VSS.n418 0.0119575
R76138 VSS.n9596 VSS.n444 0.0119575
R76139 VSS.n461 VSS.n460 0.0119575
R76140 VSS.n6374 VSS.n458 0.0119575
R76141 VSS.n463 VSS.n462 0.0119575
R76142 VSS.n6375 VSS.n457 0.0119575
R76143 VSS.n465 VSS.n464 0.0119575
R76144 VSS.n6376 VSS.n456 0.0119575
R76145 VSS.n467 VSS.n466 0.0119575
R76146 VSS.n6377 VSS.n455 0.0119575
R76147 VSS.n469 VSS.n468 0.0119575
R76148 VSS.n6378 VSS.n454 0.0119575
R76149 VSS.n471 VSS.n470 0.0119575
R76150 VSS.n6379 VSS.n453 0.0119575
R76151 VSS.n473 VSS.n472 0.0119575
R76152 VSS.n6380 VSS.n452 0.0119575
R76153 VSS.n475 VSS.n474 0.0119575
R76154 VSS.n6381 VSS.n451 0.0119575
R76155 VSS.n477 VSS.n476 0.0119575
R76156 VSS.n6382 VSS.n450 0.0119575
R76157 VSS.n479 VSS.n478 0.0119575
R76158 VSS.n6383 VSS.n449 0.0119575
R76159 VSS.n481 VSS.n480 0.0119575
R76160 VSS.n482 VSS.n448 0.0119575
R76161 VSS.n9583 VSS.n501 0.0119575
R76162 VSS.n511 VSS.n509 0.0119575
R76163 VSS.n523 VSS.n512 0.0119575
R76164 VSS.n513 VSS.n508 0.0119575
R76165 VSS.n522 VSS.n514 0.0119575
R76166 VSS.n515 VSS.n507 0.0119575
R76167 VSS.n521 VSS.n516 0.0119575
R76168 VSS.n517 VSS.n506 0.0119575
R76169 VSS.n520 VSS.n518 0.0119575
R76170 VSS.n519 VSS.n505 0.0119575
R76171 VSS.n9570 VSS.n539 0.0119575
R76172 VSS.n549 VSS.n547 0.0119575
R76173 VSS.n561 VSS.n550 0.0119575
R76174 VSS.n551 VSS.n546 0.0119575
R76175 VSS.n560 VSS.n552 0.0119575
R76176 VSS.n553 VSS.n545 0.0119575
R76177 VSS.n559 VSS.n554 0.0119575
R76178 VSS.n555 VSS.n544 0.0119575
R76179 VSS.n558 VSS.n556 0.0119575
R76180 VSS.n557 VSS.n543 0.0119575
R76181 VSS.n9567 VSS.n563 0.0119575
R76182 VSS.n580 VSS.n579 0.0119575
R76183 VSS.n8926 VSS.n577 0.0119575
R76184 VSS.n582 VSS.n581 0.0119575
R76185 VSS.n8927 VSS.n576 0.0119575
R76186 VSS.n584 VSS.n583 0.0119575
R76187 VSS.n8928 VSS.n575 0.0119575
R76188 VSS.n586 VSS.n585 0.0119575
R76189 VSS.n8929 VSS.n574 0.0119575
R76190 VSS.n588 VSS.n587 0.0119575
R76191 VSS.n8930 VSS.n573 0.0119575
R76192 VSS.n590 VSS.n589 0.0119575
R76193 VSS.n8931 VSS.n572 0.0119575
R76194 VSS.n592 VSS.n591 0.0119575
R76195 VSS.n8932 VSS.n571 0.0119575
R76196 VSS.n594 VSS.n593 0.0119575
R76197 VSS.n8933 VSS.n570 0.0119575
R76198 VSS.n596 VSS.n595 0.0119575
R76199 VSS.n8934 VSS.n569 0.0119575
R76200 VSS.n598 VSS.n597 0.0119575
R76201 VSS.n8935 VSS.n568 0.0119575
R76202 VSS.n600 VSS.n599 0.0119575
R76203 VSS.n601 VSS.n567 0.0119575
R76204 VSS.n9564 VSS.n602 0.0119575
R76205 VSS.n618 VSS.n617 0.0119575
R76206 VSS.n9473 VSS.n615 0.0119575
R76207 VSS.n620 VSS.n619 0.0119575
R76208 VSS.n9474 VSS.n614 0.0119575
R76209 VSS.n622 VSS.n621 0.0119575
R76210 VSS.n9475 VSS.n613 0.0119575
R76211 VSS.n624 VSS.n623 0.0119575
R76212 VSS.n9476 VSS.n612 0.0119575
R76213 VSS.n626 VSS.n625 0.0119575
R76214 VSS.n9477 VSS.n611 0.0119575
R76215 VSS.n628 VSS.n627 0.0119575
R76216 VSS.n9478 VSS.n610 0.0119575
R76217 VSS.n630 VSS.n629 0.0119575
R76218 VSS.n9479 VSS.n609 0.0119575
R76219 VSS.n632 VSS.n631 0.0119575
R76220 VSS.n9480 VSS.n608 0.0119575
R76221 VSS.n634 VSS.n633 0.0119575
R76222 VSS.n9481 VSS.n607 0.0119575
R76223 VSS.n636 VSS.n635 0.0119575
R76224 VSS.n9482 VSS.n606 0.0119575
R76225 VSS.n638 VSS.n637 0.0119575
R76226 VSS.n639 VSS.n605 0.0119575
R76227 VSS.n9561 VSS.n640 0.0119575
R76228 VSS.n657 VSS.n656 0.0119575
R76229 VSS.n9547 VSS.n654 0.0119575
R76230 VSS.n659 VSS.n658 0.0119575
R76231 VSS.n9548 VSS.n653 0.0119575
R76232 VSS.n661 VSS.n660 0.0119575
R76233 VSS.n9549 VSS.n652 0.0119575
R76234 VSS.n663 VSS.n662 0.0119575
R76235 VSS.n9550 VSS.n651 0.0119575
R76236 VSS.n665 VSS.n664 0.0119575
R76237 VSS.n9551 VSS.n650 0.0119575
R76238 VSS.n667 VSS.n666 0.0119575
R76239 VSS.n9552 VSS.n649 0.0119575
R76240 VSS.n669 VSS.n668 0.0119575
R76241 VSS.n9553 VSS.n648 0.0119575
R76242 VSS.n671 VSS.n670 0.0119575
R76243 VSS.n9554 VSS.n647 0.0119575
R76244 VSS.n673 VSS.n672 0.0119575
R76245 VSS.n9555 VSS.n646 0.0119575
R76246 VSS.n675 VSS.n674 0.0119575
R76247 VSS.n9556 VSS.n645 0.0119575
R76248 VSS.n677 VSS.n676 0.0119575
R76249 VSS.n9558 VSS.n644 0.0119575
R76250 VSS.n142 VSS.n140 0.0119575
R76251 VSS.n6048 VSS.n6047 0.0119575
R76252 VSS.n6040 VSS.n6039 0.0119575
R76253 VSS.n5946 VSS.n5916 0.0119575
R76254 VSS.n5938 VSS.n5923 0.0119575
R76255 VSS.n6063 VSS.n6050 0.0119575
R76256 VSS.n6070 VSS.n6042 0.0119575
R76257 VSS.n5948 VSS.n5910 0.0119575
R76258 VSS.n5940 VSS.n5917 0.0119575
R76259 VSS.n6051 VSS.n3952 0.0119575
R76260 VSS.n6043 VSS.n3996 0.0119575
R76261 VSS.n5951 VSS.n325 0.0119575
R76262 VSS.n5943 VSS.n359 0.0119575
R76263 VSS.n6067 VSS.n6052 0.0119575
R76264 VSS.n6074 VSS.n6044 0.0119575
R76265 VSS.n5950 VSS.n5912 0.0119575
R76266 VSS.n5942 VSS.n5919 0.0119575
R76267 VSS.n3812 VSS.n3811 0.0119575
R76268 VSS.n3803 VSS.n3802 0.0119575
R76269 VSS.n3699 VSS.n3698 0.0119575
R76270 VSS.n3690 VSS.n3689 0.0119575
R76271 VSS.n6289 VSS.n3814 0.0119575
R76272 VSS.n6296 VSS.n3805 0.0119575
R76273 VSS.n6318 VSS.n3701 0.0119575
R76274 VSS.n6325 VSS.n3692 0.0119575
R76275 VSS.n3815 VSS.n3810 0.0119575
R76276 VSS.n3806 VSS.n3801 0.0119575
R76277 VSS.n3702 VSS.n3697 0.0119575
R76278 VSS.n3693 VSS.n3688 0.0119575
R76279 VSS.n6293 VSS.n3816 0.0119575
R76280 VSS.n6300 VSS.n3807 0.0119575
R76281 VSS.n6322 VSS.n3703 0.0119575
R76282 VSS.n6329 VSS.n3694 0.0119575
R76283 VSS.n3218 VSS.n3217 0.0119575
R76284 VSS.n3209 VSS.n3208 0.0119575
R76285 VSS.n3200 VSS.n3199 0.0119575
R76286 VSS.n3122 VSS.n3121 0.0119575
R76287 VSS.n3117 VSS.n3113 0.0119575
R76288 VSS.n6583 VSS.n3220 0.0119575
R76289 VSS.n6589 VSS.n3211 0.0119575
R76290 VSS.n6596 VSS.n3202 0.0119575
R76291 VSS.n6624 VSS.n3123 0.0119575
R76292 VSS.n6631 VSS.n3118 0.0119575
R76293 VSS.n3221 VSS.n3216 0.0119575
R76294 VSS.n3212 VSS.n3207 0.0119575
R76295 VSS.n3203 VSS.n3198 0.0119575
R76296 VSS.n3124 VSS.n3120 0.0119575
R76297 VSS.n6633 VSS.n3116 0.0119575
R76298 VSS.n6587 VSS.n3222 0.0119575
R76299 VSS.n6593 VSS.n3213 0.0119575
R76300 VSS.n6600 VSS.n3204 0.0119575
R76301 VSS.n6628 VSS.n3125 0.0119575
R76302 VSS.n6637 VSS.n6634 0.0119575
R76303 VSS.n5761 VSS.n5760 0.0119575
R76304 VSS.n5752 VSS.n5751 0.0119575
R76305 VSS.n5743 VSS.n5742 0.0119575
R76306 VSS.n2971 VSS.n2969 0.0119575
R76307 VSS.n6642 VSS.n6641 0.0119575
R76308 VSS.n5781 VSS.n5763 0.0119575
R76309 VSS.n5787 VSS.n5754 0.0119575
R76310 VSS.n5794 VSS.n5745 0.0119575
R76311 VSS.n6756 VSS.n2963 0.0119575
R76312 VSS.n6648 VSS.n6644 0.0119575
R76313 VSS.n5764 VSS.n5759 0.0119575
R76314 VSS.n5755 VSS.n5750 0.0119575
R76315 VSS.n5746 VSS.n5741 0.0119575
R76316 VSS.n6759 VSS.n6758 0.0119575
R76317 VSS.n6645 VSS.n6640 0.0119575
R76318 VSS.n5785 VSS.n5765 0.0119575
R76319 VSS.n5791 VSS.n5756 0.0119575
R76320 VSS.n5798 VSS.n5747 0.0119575
R76321 VSS.n6754 VSS.n2965 0.0119575
R76322 VSS.n6652 VSS.n6646 0.0119575
R76323 VSS.n2762 VSS.n2761 0.0119575
R76324 VSS.n2753 VSS.n2752 0.0119575
R76325 VSS.n2744 VSS.n2743 0.0119575
R76326 VSS.n2637 VSS.n2636 0.0119575
R76327 VSS.n2628 VSS.n2627 0.0119575
R76328 VSS.n6975 VSS.n2764 0.0119575
R76329 VSS.n6981 VSS.n2755 0.0119575
R76330 VSS.n6988 VSS.n2746 0.0119575
R76331 VSS.n7010 VSS.n2639 0.0119575
R76332 VSS.n7017 VSS.n2630 0.0119575
R76333 VSS.n2765 VSS.n2760 0.0119575
R76334 VSS.n2756 VSS.n2751 0.0119575
R76335 VSS.n2747 VSS.n2742 0.0119575
R76336 VSS.n2640 VSS.n2635 0.0119575
R76337 VSS.n2631 VSS.n2626 0.0119575
R76338 VSS.n6979 VSS.n2766 0.0119575
R76339 VSS.n6985 VSS.n2757 0.0119575
R76340 VSS.n6992 VSS.n2748 0.0119575
R76341 VSS.n7014 VSS.n2641 0.0119575
R76342 VSS.n7021 VSS.n2632 0.0119575
R76343 VSS.n115 VSS.n109 0.0119575
R76344 VSS.n119 VSS.n103 0.0119575
R76345 VSS.n111 VSS.n107 0.0119575
R76346 VSS.n118 VSS.n102 0.0119575
R76347 VSS.n112 VSS.n108 0.0119575
R76348 VSS.n117 VSS.n101 0.0119575
R76349 VSS.n210 VSS.n209 0.0119575
R76350 VSS.n213 VSS.n198 0.0119575
R76351 VSS.n212 VSS.n208 0.0119575
R76352 VSS.n215 VSS.n199 0.0119575
R76353 VSS.n214 VSS.n207 0.0119575
R76354 VSS.n9775 VSS.n200 0.0119575
R76355 VSS.n5416 VSS.n5410 0.0119575
R76356 VSS.n5501 VSS.n5419 0.0119575
R76357 VSS.n5418 VSS.n5409 0.0119575
R76358 VSS.n5502 VSS.n5421 0.0119575
R76359 VSS.n5420 VSS.n5408 0.0119575
R76360 VSS.n5505 VSS.n5504 0.0119575
R76361 VSS.n388 VSS.n386 0.0119575
R76362 VSS.n9624 VSS.n391 0.0119575
R76363 VSS.n390 VSS.n385 0.0119575
R76364 VSS.n9625 VSS.n393 0.0119575
R76365 VSS.n392 VSS.n384 0.0119575
R76366 VSS.n5936 VSS.n5935 0.0119575
R76367 VSS.n5933 VSS.n5926 0.0119575
R76368 VSS.n5930 VSS.n5924 0.0119575
R76369 VSS.n5932 VSS.n5931 0.0119575
R76370 VSS.n6337 VSS.n6333 0.0119575
R76371 VSS.n6334 VSS.n3686 0.0119575
R76372 VSS.n6331 VSS.n3685 0.0119575
R76373 VSS.n6339 VSS.n3681 0.0119575
R76374 VSS.n6342 VSS.n3643 0.0119575
R76375 VSS.n6359 VSS.n3680 0.0119575
R76376 VSS.n6343 VSS.n3644 0.0119575
R76377 VSS.n6358 VSS.n3679 0.0119575
R76378 VSS.n6344 VSS.n3645 0.0119575
R76379 VSS.n6357 VSS.n3678 0.0119575
R76380 VSS.n6345 VSS.n3646 0.0119575
R76381 VSS.n6356 VSS.n3677 0.0119575
R76382 VSS.n6346 VSS.n3647 0.0119575
R76383 VSS.n6355 VSS.n3676 0.0119575
R76384 VSS.n6347 VSS.n3648 0.0119575
R76385 VSS.n6354 VSS.n3675 0.0119575
R76386 VSS.n6348 VSS.n3649 0.0119575
R76387 VSS.n6353 VSS.n3674 0.0119575
R76388 VSS.n6349 VSS.n3650 0.0119575
R76389 VSS.n6352 VSS.n3673 0.0119575
R76390 VSS.n6350 VSS.n3651 0.0119575
R76391 VSS.n6351 VSS.n3672 0.0119575
R76392 VSS.n6398 VSS.n3652 0.0119575
R76393 VSS.n6397 VSS.n3671 0.0119575
R76394 VSS.n6399 VSS.n3653 0.0119575
R76395 VSS.n6401 VSS.n3670 0.0119575
R76396 VSS.n6402 VSS.n3669 0.0119575
R76397 VSS.n3666 VSS.n3655 0.0119575
R76398 VSS.n3661 VSS.n3660 0.0119575
R76399 VSS.n3662 VSS.n3657 0.0119575
R76400 VSS.n3659 VSS.n3658 0.0119575
R76401 VSS.n6660 VSS.n6656 0.0119575
R76402 VSS.n6657 VSS.n3111 0.0119575
R76403 VSS.n6654 VSS.n3110 0.0119575
R76404 VSS.n6662 VSS.n3106 0.0119575
R76405 VSS.n3104 VSS.n3097 0.0119575
R76406 VSS.n6691 VSS.n6664 0.0119575
R76407 VSS.n3103 VSS.n3096 0.0119575
R76408 VSS.n6692 VSS.n6665 0.0119575
R76409 VSS.n3102 VSS.n3095 0.0119575
R76410 VSS.n6693 VSS.n6666 0.0119575
R76411 VSS.n3101 VSS.n3094 0.0119575
R76412 VSS.n6696 VSS.n6695 0.0119575
R76413 VSS.n3100 VSS.n3093 0.0119575
R76414 VSS.n6698 VSS.n3099 0.0119575
R76415 VSS.n7029 VSS.n7025 0.0119575
R76416 VSS.n7026 VSS.n2624 0.0119575
R76417 VSS.n7023 VSS.n2623 0.0119575
R76418 VSS.n7031 VSS.n2619 0.0119575
R76419 VSS.n1268 VSS.n1266 0.0119575
R76420 VSS.n8902 VSS.n1271 0.0119575
R76421 VSS.n1270 VSS.n1265 0.0119575
R76422 VSS.n8903 VSS.n1273 0.0119575
R76423 VSS.n1272 VSS.n1264 0.0119575
R76424 VSS.n8904 VSS.n1275 0.0119575
R76425 VSS.n1274 VSS.n1263 0.0119575
R76426 VSS.n8908 VSS.n8906 0.0119575
R76427 VSS.n8907 VSS.n1262 0.0119575
R76428 VSS.n8910 VSS.n1258 0.0119575
R76429 VSS.n1256 VSS.n1153 0.0119575
R76430 VSS.n1257 VSS.n1255 0.0119575
R76431 VSS.n1253 VSS.n1154 0.0119575
R76432 VSS.n1254 VSS.n1252 0.0119575
R76433 VSS.n1250 VSS.n1155 0.0119575
R76434 VSS.n1251 VSS.n1249 0.0119575
R76435 VSS.n1247 VSS.n1156 0.0119575
R76436 VSS.n1248 VSS.n1246 0.0119575
R76437 VSS.n1244 VSS.n1157 0.0119575
R76438 VSS.n1245 VSS.n1243 0.0119575
R76439 VSS.n1241 VSS.n1158 0.0119575
R76440 VSS.n1242 VSS.n1240 0.0119575
R76441 VSS.n1238 VSS.n1159 0.0119575
R76442 VSS.n1239 VSS.n1237 0.0119575
R76443 VSS.n1235 VSS.n1160 0.0119575
R76444 VSS.n1236 VSS.n1234 0.0119575
R76445 VSS.n1232 VSS.n1161 0.0119575
R76446 VSS.n1233 VSS.n1231 0.0119575
R76447 VSS.n1229 VSS.n1162 0.0119575
R76448 VSS.n1230 VSS.n1228 0.0119575
R76449 VSS.n1226 VSS.n1163 0.0119575
R76450 VSS.n1227 VSS.n1151 0.0119575
R76451 VSS.n2623 VSS.n2619 0.0119575
R76452 VSS.n7023 VSS.n2624 0.0119575
R76453 VSS.n3110 VSS.n3106 0.0119575
R76454 VSS.n6654 VSS.n3111 0.0119575
R76455 VSS.n3658 VSS.n3657 0.0119575
R76456 VSS.n3662 VSS.n3660 0.0119575
R76457 VSS.n3685 VSS.n3681 0.0119575
R76458 VSS.n6331 VSS.n3686 0.0119575
R76459 VSS.n5931 VSS.n5930 0.0119575
R76460 VSS.n5933 VSS.n5924 0.0119575
R76461 VSS.n5936 VSS.n397 0.0119575
R76462 VSS.n5935 VSS.n5926 0.0119575
R76463 VSS.n6333 VSS.n3684 0.0119575
R76464 VSS.n6337 VSS.n6334 0.0119575
R76465 VSS.n3668 VSS.n3655 0.0119575
R76466 VSS.n3666 VSS.n3661 0.0119575
R76467 VSS.n6656 VSS.n3109 0.0119575
R76468 VSS.n6660 VSS.n6657 0.0119575
R76469 VSS.n7025 VSS.n2622 0.0119575
R76470 VSS.n7029 VSS.n7026 0.0119575
R76471 VSS.n119 VSS.n106 0.0119575
R76472 VSS.n111 VSS.n103 0.0119575
R76473 VSS.n118 VSS.n107 0.0119575
R76474 VSS.n112 VSS.n102 0.0119575
R76475 VSS.n117 VSS.n108 0.0119575
R76476 VSS.n209 VSS.n197 0.0119575
R76477 VSS.n210 VSS.n198 0.0119575
R76478 VSS.n213 VSS.n212 0.0119575
R76479 VSS.n208 VSS.n199 0.0119575
R76480 VSS.n215 VSS.n214 0.0119575
R76481 VSS.n207 VSS.n200 0.0119575
R76482 VSS.n5417 VSS.n5416 0.0119575
R76483 VSS.n5501 VSS.n5410 0.0119575
R76484 VSS.n5419 VSS.n5418 0.0119575
R76485 VSS.n5502 VSS.n5409 0.0119575
R76486 VSS.n5421 VSS.n5420 0.0119575
R76487 VSS.n5504 VSS.n5408 0.0119575
R76488 VSS.n389 VSS.n388 0.0119575
R76489 VSS.n9624 VSS.n386 0.0119575
R76490 VSS.n391 VSS.n390 0.0119575
R76491 VSS.n9625 VSS.n385 0.0119575
R76492 VSS.n393 VSS.n392 0.0119575
R76493 VSS.n6340 VSS.n3643 0.0119575
R76494 VSS.n6359 VSS.n6342 0.0119575
R76495 VSS.n3680 VSS.n3644 0.0119575
R76496 VSS.n6358 VSS.n6343 0.0119575
R76497 VSS.n3679 VSS.n3645 0.0119575
R76498 VSS.n6357 VSS.n6344 0.0119575
R76499 VSS.n3678 VSS.n3646 0.0119575
R76500 VSS.n6356 VSS.n6345 0.0119575
R76501 VSS.n3677 VSS.n3647 0.0119575
R76502 VSS.n6355 VSS.n6346 0.0119575
R76503 VSS.n3676 VSS.n3648 0.0119575
R76504 VSS.n6354 VSS.n6347 0.0119575
R76505 VSS.n3675 VSS.n3649 0.0119575
R76506 VSS.n6353 VSS.n6348 0.0119575
R76507 VSS.n3674 VSS.n3650 0.0119575
R76508 VSS.n6352 VSS.n6349 0.0119575
R76509 VSS.n3673 VSS.n3651 0.0119575
R76510 VSS.n6351 VSS.n6350 0.0119575
R76511 VSS.n3672 VSS.n3652 0.0119575
R76512 VSS.n6398 VSS.n6397 0.0119575
R76513 VSS.n3671 VSS.n3653 0.0119575
R76514 VSS.n6399 VSS.n3670 0.0119575
R76515 VSS.n6402 VSS.n6401 0.0119575
R76516 VSS.n6663 VSS.n3097 0.0119575
R76517 VSS.n6691 VSS.n3104 0.0119575
R76518 VSS.n6664 VSS.n3096 0.0119575
R76519 VSS.n6692 VSS.n3103 0.0119575
R76520 VSS.n6665 VSS.n3095 0.0119575
R76521 VSS.n6693 VSS.n3102 0.0119575
R76522 VSS.n6666 VSS.n3094 0.0119575
R76523 VSS.n6695 VSS.n3101 0.0119575
R76524 VSS.n6696 VSS.n3093 0.0119575
R76525 VSS.n3100 VSS.n3099 0.0119575
R76526 VSS.n1269 VSS.n1268 0.0119575
R76527 VSS.n8902 VSS.n1266 0.0119575
R76528 VSS.n1271 VSS.n1270 0.0119575
R76529 VSS.n8903 VSS.n1265 0.0119575
R76530 VSS.n1273 VSS.n1272 0.0119575
R76531 VSS.n8904 VSS.n1264 0.0119575
R76532 VSS.n1275 VSS.n1274 0.0119575
R76533 VSS.n8906 VSS.n1263 0.0119575
R76534 VSS.n8908 VSS.n8907 0.0119575
R76535 VSS.n1262 VSS.n1258 0.0119575
R76536 VSS.n8911 VSS.n1153 0.0119575
R76537 VSS.n1257 VSS.n1256 0.0119575
R76538 VSS.n1255 VSS.n1154 0.0119575
R76539 VSS.n1254 VSS.n1253 0.0119575
R76540 VSS.n1252 VSS.n1155 0.0119575
R76541 VSS.n1251 VSS.n1250 0.0119575
R76542 VSS.n1249 VSS.n1156 0.0119575
R76543 VSS.n1248 VSS.n1247 0.0119575
R76544 VSS.n1246 VSS.n1157 0.0119575
R76545 VSS.n1245 VSS.n1244 0.0119575
R76546 VSS.n1243 VSS.n1158 0.0119575
R76547 VSS.n1242 VSS.n1241 0.0119575
R76548 VSS.n1240 VSS.n1159 0.0119575
R76549 VSS.n1239 VSS.n1238 0.0119575
R76550 VSS.n1237 VSS.n1160 0.0119575
R76551 VSS.n1236 VSS.n1235 0.0119575
R76552 VSS.n1234 VSS.n1161 0.0119575
R76553 VSS.n1233 VSS.n1232 0.0119575
R76554 VSS.n1231 VSS.n1162 0.0119575
R76555 VSS.n1230 VSS.n1229 0.0119575
R76556 VSS.n1228 VSS.n1163 0.0119575
R76557 VSS.n1227 VSS.n1226 0.0119575
R76558 VSS.n115 VSS.n100 0.0119575
R76559 VSS.n2363 VSS.n2362 0.0119575
R76560 VSS.n2358 VSS.n2357 0.0119575
R76561 VSS.n9443 VSS.n9442 0.0119575
R76562 VSS.n9438 VSS.n9437 0.0119575
R76563 VSS.n2340 VSS.n2336 0.0119575
R76564 VSS.n2347 VSS.n2343 0.0119575
R76565 VSS.n775 VSS.n770 0.0119575
R76566 VSS.n9372 VSS.n778 0.0119575
R76567 VSS.n2365 VSS.n2337 0.0119575
R76568 VSS.n2360 VSS.n2344 0.0119575
R76569 VSS.n9445 VSS.n772 0.0119575
R76570 VSS.n9440 VSS.n9369 0.0119575
R76571 VSS.n2085 VSS.n2081 0.0119575
R76572 VSS.n2436 VSS.n2432 0.0119575
R76573 VSS.n2459 VSS.n2452 0.0119575
R76574 VSS.n1095 VSS.n1091 0.0119575
R76575 VSS.n2087 VSS.n2083 0.0119575
R76576 VSS.n2431 VSS.n1542 0.0119575
R76577 VSS.n2460 VSS.n1429 0.0119575
R76578 VSS.n1097 VSS.n1093 0.0119575
R76579 VSS.n4453 VSS.n13 0.0116972
R76580 VSS.n5659 VSS.n4249 0.0116972
R76581 VSS.n4120 VSS.n4116 0.0116972
R76582 VSS.n5727 VSS.n4122 0.0116972
R76583 VSS.n5722 VSS.n4119 0.0116972
R76584 VSS.n4169 VSS.n4117 0.0116972
R76585 VSS.n5725 VSS.n5724 0.0116972
R76586 VSS.n4661 VSS.n4428 0.0116972
R76587 VSS.n5661 VSS.n4267 0.0116972
R76588 VSS.n4076 VSS.n4025 0.0116972
R76589 VSS.n4114 VSS.n4016 0.0116972
R76590 VSS.n4078 VSS.n4026 0.0116972
R76591 VSS.n4111 VSS.n4015 0.0116972
R76592 VSS.n6124 VSS.n4027 0.0116972
R76593 VSS.n2311 VSS.n2162 0.0116614
R76594 VSS.n2415 VSS.n1848 0.0116614
R76595 VSS.n1185 VSS.n750 0.0116614
R76596 VSS.n9387 VSS.n695 0.0116614
R76597 VSS.n4457 VSS.n4455 0.0114859
R76598 VSS.n5121 VSS.n4431 0.0114859
R76599 VSS.n2277 VSS.n2172 0.0113607
R76600 VSS.n1166 VSS.n1094 0.0113607
R76601 VSS.n2275 VSS.n2172 0.0113607
R76602 VSS.n1167 VSS.n1166 0.0113607
R76603 VSS.n2311 VSS.n2147 0.0113071
R76604 VSS.n2415 VSS.n1853 0.0113071
R76605 VSS.n1185 VSS.n734 0.0113071
R76606 VSS.n9387 VSS.n699 0.0113071
R76607 VSS.n4967 VSS.n4868 0.0112746
R76608 VSS.n4972 VSS.n4850 0.0112746
R76609 VSS.n4969 VSS.n4869 0.0112746
R76610 VSS.n4870 VSS.n4849 0.0112746
R76611 VSS.n5019 VSS.n4974 0.0112746
R76612 VSS.n5719 VSS.n4174 0.0112746
R76613 VSS.n3740 VSS.n3157 0.0112746
R76614 VSS.n9450 VSS.n766 0.0112746
R76615 VSS.n4508 VSS.n4503 0.0112746
R76616 VSS.n5080 VSS.n4496 0.0112746
R76617 VSS.n4511 VSS.n4504 0.0112746
R76618 VSS.n4505 VSS.n4495 0.0112746
R76619 VSS.n5083 VSS.n5082 0.0112746
R76620 VSS.n4074 VSS.n4018 0.0112746
R76621 VSS.n3759 VSS.n3187 0.0112746
R76622 VSS.n9222 VSS.n915 0.0112746
R76623 VSS.n2295 VSS.n2150 0.0109528
R76624 VSS.n1201 VSS.n737 0.0109528
R76625 VSS.n9456 VSS.n9455 0.0108846
R76626 VSS.n9455 VSS.n759 0.0108846
R76627 VSS.n7890 VSS.n7889 0.0108846
R76628 VSS.n7889 VSS.n2426 0.0108846
R76629 VSS.n3726 VSS.n3147 0.0108521
R76630 VSS.n6804 VSS.n2953 0.0108521
R76631 VSS.n8711 VSS.n1460 0.0108521
R76632 VSS.n3787 VSS.n3177 0.0108521
R76633 VSS.n6799 VSS.n2935 0.0108521
R76634 VSS.n8685 VSS.n1493 0.0108521
R76635 VSS.n4759 VSS.n4756 0.0107778
R76636 VSS.n9812 VSS.n175 0.0107778
R76637 VSS.n6251 VSS.n3864 0.0107778
R76638 VSS.n5466 VSS.n5465 0.0107778
R76639 VSS.n4092 VSS.n3854 0.0107778
R76640 VSS.n4158 VSS.n4157 0.0107778
R76641 VSS.n6057 VSS.n3829 0.0107778
R76642 VSS.n9605 VSS.n428 0.0107778
R76643 VSS.n6283 VSS.n6282 0.0107778
R76644 VSS.n9600 VSS.n437 0.0107778
R76645 VSS.n6582 VSS.n6581 0.0107778
R76646 VSS.n9592 VSS.n485 0.0107778
R76647 VSS.n5780 VSS.n5779 0.0107778
R76648 VSS.n9587 VSS.n494 0.0107778
R76649 VSS.n6974 VSS.n6973 0.0107778
R76650 VSS.n9579 VSS.n527 0.0107778
R76651 VSS.n5446 VSS.n5386 0.0105984
R76652 VSS.n5456 VSS.n5384 0.0105984
R76653 VSS.n5449 VSS.n5387 0.0105984
R76654 VSS.n5452 VSS.n5383 0.0105984
R76655 VSS.n5448 VSS.n5393 0.0105984
R76656 VSS.n2327 VSS.n2165 0.0105984
R76657 VSS.n2399 VSS.n1845 0.0105984
R76658 VSS.n9687 VSS.n280 0.0105984
R76659 VSS.n9685 VSS.n9684 0.0105984
R76660 VSS.n298 VSS.n286 0.0105984
R76661 VSS.n297 VSS.n294 0.0105984
R76662 VSS.n300 VSS.n285 0.0105984
R76663 VSS.n4284 VSS.n4280 0.0105984
R76664 VSS.n5647 VSS.n4287 0.0105984
R76665 VSS.n4288 VSS.n4283 0.0105984
R76666 VSS.n5643 VSS.n5642 0.0105984
R76667 VSS.n5632 VSS.n4282 0.0105984
R76668 VSS.n5253 VSS.n4316 0.0105984
R76669 VSS.n5261 VSS.n4315 0.0105984
R76670 VSS.n5256 VSS.n4317 0.0105984
R76671 VSS.n5258 VSS.n4314 0.0105984
R76672 VSS.n5264 VSS.n5263 0.0105984
R76673 VSS.n4744 VSS.n4726 0.0105984
R76674 VSS.n6250 VSS.n6249 0.0105984
R76675 VSS.n9808 VSS.n169 0.0105984
R76676 VSS.n5471 VSS.n5439 0.0105984
R76677 VSS.n5441 VSS.n5414 0.0105984
R76678 VSS.n5463 VSS.n5412 0.0105984
R76679 VSS.n5444 VSS.n5415 0.0105984
R76680 VSS.n5459 VSS.n5411 0.0105984
R76681 VSS.n5443 VSS.n5417 0.0105984
R76682 VSS.n1169 VSS.n753 0.0105984
R76683 VSS.n9403 VSS.n692 0.0105984
R76684 VSS.n7045 VSS.n2616 0.0105466
R76685 VSS.n7047 VSS.n2609 0.0105466
R76686 VSS.n7052 VSS.n2605 0.0105466
R76687 VSS.n8857 VSS.n1310 0.0105466
R76688 VSS.n8834 VSS.n1349 0.0105466
R76689 VSS.n8837 VSS.n1351 0.0105466
R76690 VSS.n8041 VSS.n8033 0.0105466
R76691 VSS.n2784 VSS.n2778 0.0105466
R76692 VSS.n2787 VSS.n2779 0.0105466
R76693 VSS.n2274 VSS.n2273 0.0105466
R76694 VSS.n2271 VSS.n2171 0.0105466
R76695 VSS.n2333 VSS.n2331 0.0105466
R76696 VSS.n2368 VSS.n2367 0.0105466
R76697 VSS.n2334 VSS.n2332 0.0105466
R76698 VSS.n7152 VSS.n2570 0.0105466
R76699 VSS.n7156 VSS.n2564 0.0105466
R76700 VSS.n7162 VSS.n2552 0.0105466
R76701 VSS.n7163 VSS.n2548 0.0105466
R76702 VSS.n7168 VSS.n2549 0.0105466
R76703 VSS.n2530 VSS.n2529 0.0105466
R76704 VSS.n7222 VSS.n2531 0.0105466
R76705 VSS.n7094 VSS.n7090 0.0105466
R76706 VSS.n7096 VSS.n7059 0.0105466
R76707 VSS.n7100 VSS.n7099 0.0105466
R76708 VSS.n7106 VSS.n2603 0.0105466
R76709 VSS.n8848 VSS.n1316 0.0105466
R76710 VSS.n1348 VSS.n1343 0.0105466
R76711 VSS.n8807 VSS.n1391 0.0105466
R76712 VSS.n8032 VSS.n8026 0.0105466
R76713 VSS.n7153 VSS.n7152 0.0105466
R76714 VSS.n7153 VSS.n2564 0.0105466
R76715 VSS.n7101 VSS.n7100 0.0105466
R76716 VSS.n2531 VSS.n2530 0.0105466
R76717 VSS.n2529 VSS.n2528 0.0105466
R76718 VSS.n7094 VSS.n7059 0.0105466
R76719 VSS.n7090 VSS.n2532 0.0105466
R76720 VSS.n2549 VSS.n2548 0.0105466
R76721 VSS.n7166 VSS.n7163 0.0105466
R76722 VSS.n7159 VSS.n2552 0.0105466
R76723 VSS.n7138 VSS.n2577 0.0105466
R76724 VSS.n7136 VSS.n2578 0.0105466
R76725 VSS.n7262 VSS.n2481 0.0105466
R76726 VSS.n2488 VSS.n2483 0.0105466
R76727 VSS.n7257 VSS.n2490 0.0105466
R76728 VSS.n7188 VSS.n7187 0.0105466
R76729 VSS.n7197 VSS.n7189 0.0105466
R76730 VSS.n7240 VSS.n7236 0.0105466
R76731 VSS.n7242 VSS.n2507 0.0105466
R76732 VSS.n7247 VSS.n2504 0.0105466
R76733 VSS.n7121 VSS.n2592 0.0105466
R76734 VSS.n8388 VSS.n1662 0.0105466
R76735 VSS.n1603 VSS.n1596 0.0105466
R76736 VSS.n8549 VSS.n1598 0.0105466
R76737 VSS.n8017 VSS.n8011 0.0105466
R76738 VSS.n2481 VSS.n2480 0.0105466
R76739 VSS.n7243 VSS.n2504 0.0105466
R76740 VSS.n7240 VSS.n2507 0.0105466
R76741 VSS.n7236 VSS.n2511 0.0105466
R76742 VSS.n7189 VSS.n7188 0.0105466
R76743 VSS.n7187 VSS.n2491 0.0105466
R76744 VSS.n2490 VSS.n2488 0.0105466
R76745 VSS.n7259 VSS.n2483 0.0105466
R76746 VSS.n7129 VSS.n2581 0.0105466
R76747 VSS.n7127 VSS.n2582 0.0105466
R76748 VSS.n7124 VSS.n2587 0.0105466
R76749 VSS.n8564 VSS.n1561 0.0105466
R76750 VSS.n8557 VSS.n8556 0.0105466
R76751 VSS.n8554 VSS.n1593 0.0105466
R76752 VSS.n8010 VSS.n8008 0.0105466
R76753 VSS.n8547 VSS.n1603 0.0105466
R76754 VSS.n8840 VSS.n1343 0.0105466
R76755 VSS.n8834 VSS.n1305 0.0105466
R76756 VSS.n1351 VSS.n1349 0.0105466
R76757 VSS.n1391 VSS.n1348 0.0105466
R76758 VSS.n1598 VSS.n1596 0.0105466
R76759 VSS.n1593 VSS.n1590 0.0105466
R76760 VSS.n8556 VSS.n1590 0.0105466
R76761 VSS.n8072 VSS.n8010 0.0105466
R76762 VSS.n8067 VSS.n8017 0.0105466
R76763 VSS.n8048 VSS.n8032 0.0105466
R76764 VSS.n8043 VSS.n8041 0.0105466
R76765 VSS.n8851 VSS.n1310 0.0105466
R76766 VSS.n8844 VSS.n1316 0.0105466
R76767 VSS.n8392 VSS.n8388 0.0105466
R76768 VSS.n1561 VSS.n1559 0.0105466
R76769 VSS.n7126 VSS.n2587 0.0105466
R76770 VSS.n2592 VSS.n2505 0.0105466
R76771 VSS.n7102 VSS.n2603 0.0105466
R76772 VSS.n7048 VSS.n2605 0.0105466
R76773 VSS.n7138 VSS.n2578 0.0105466
R76774 VSS.n2577 VSS.n2576 0.0105466
R76775 VSS.n2779 VSS.n2778 0.0105466
R76776 VSS.n7129 VSS.n2582 0.0105466
R76777 VSS.n2784 VSS.n2783 0.0105466
R76778 VSS.n2581 VSS.n2580 0.0105466
R76779 VSS.n6269 VSS.n3831 0.0105466
R76780 VSS.n6271 VSS.n6270 0.0105466
R76781 VSS.n6272 VSS.n6271 0.0105466
R76782 VSS.n6274 VSS.n3828 0.0105466
R76783 VSS.n6276 VSS.n3823 0.0105466
R76784 VSS.n6277 VSS.n3824 0.0105466
R76785 VSS.n6279 VSS.n3824 0.0105466
R76786 VSS.n6281 VSS.n3826 0.0105466
R76787 VSS.n6575 VSS.n3225 0.0105466
R76788 VSS.n6576 VSS.n3226 0.0105466
R76789 VSS.n6578 VSS.n3226 0.0105466
R76790 VSS.n6580 VSS.n3228 0.0105466
R76791 VSS.n5773 VSS.n5768 0.0105466
R76792 VSS.n5774 VSS.n5769 0.0105466
R76793 VSS.n5776 VSS.n5769 0.0105466
R76794 VSS.n5778 VSS.n5771 0.0105466
R76795 VSS.n6967 VSS.n2769 0.0105466
R76796 VSS.n6968 VSS.n2770 0.0105466
R76797 VSS.n6970 VSS.n2770 0.0105466
R76798 VSS.n6972 VSS.n2772 0.0105466
R76799 VSS.n2793 VSS.n2773 0.0105466
R76800 VSS.n2793 VSS.n2792 0.0105466
R76801 VSS.n9606 VSS.n427 0.0105466
R76802 VSS.n432 VSS.n430 0.0105466
R76803 VSS.n9601 VSS.n436 0.0105466
R76804 VSS.n441 VSS.n439 0.0105466
R76805 VSS.n9593 VSS.n484 0.0105466
R76806 VSS.n489 VSS.n487 0.0105466
R76807 VSS.n9588 VSS.n493 0.0105466
R76808 VSS.n498 VSS.n496 0.0105466
R76809 VSS.n9580 VSS.n526 0.0105466
R76810 VSS.n531 VSS.n529 0.0105466
R76811 VSS.n9575 VSS.n535 0.0105466
R76812 VSS.n9602 VSS.n430 0.0105466
R76813 VSS.n6270 VSS.n6269 0.0105466
R76814 VSS.n6265 VSS.n3831 0.0105466
R76815 VSS.n431 VSS.n427 0.0105466
R76816 VSS.n6268 VSS.n3828 0.0105466
R76817 VSS.n6272 VSS.n6268 0.0105466
R76818 VSS.n9597 VSS.n439 0.0105466
R76819 VSS.n6277 VSS.n3823 0.0105466
R76820 VSS.n6276 VSS.n6275 0.0105466
R76821 VSS.n440 VSS.n436 0.0105466
R76822 VSS.n3826 VSS.n3822 0.0105466
R76823 VSS.n6279 VSS.n3822 0.0105466
R76824 VSS.n9589 VSS.n487 0.0105466
R76825 VSS.n6576 VSS.n3225 0.0105466
R76826 VSS.n6575 VSS.n6574 0.0105466
R76827 VSS.n488 VSS.n484 0.0105466
R76828 VSS.n3228 VSS.n3224 0.0105466
R76829 VSS.n6578 VSS.n3224 0.0105466
R76830 VSS.n9584 VSS.n496 0.0105466
R76831 VSS.n5774 VSS.n5768 0.0105466
R76832 VSS.n5773 VSS.n3229 0.0105466
R76833 VSS.n497 VSS.n493 0.0105466
R76834 VSS.n5771 VSS.n5767 0.0105466
R76835 VSS.n5776 VSS.n5767 0.0105466
R76836 VSS.n9576 VSS.n529 0.0105466
R76837 VSS.n6968 VSS.n2769 0.0105466
R76838 VSS.n6967 VSS.n6966 0.0105466
R76839 VSS.n530 VSS.n526 0.0105466
R76840 VSS.n2772 VSS.n2768 0.0105466
R76841 VSS.n6970 VSS.n2768 0.0105466
R76842 VSS.n7045 VSS.n2609 0.0105466
R76843 VSS.n2617 VSS.n2616 0.0105466
R76844 VSS.n538 VSS.n535 0.0105466
R76845 VSS.n7042 VSS.n7032 0.0105466
R76846 VSS.n7039 VSS.n7033 0.0105466
R76847 VSS.n1222 VSS.n1168 0.0105466
R76848 VSS.n1221 VSS.n1220 0.0105466
R76849 VSS.n9377 VSS.n9376 0.0105466
R76850 VSS.n9435 VSS.n9434 0.0105466
R76851 VSS.n9378 VSS.n9374 0.0105466
R76852 VSS.n7042 VSS.n7041 0.0105466
R76853 VSS.n7041 VSS.n7033 0.0105466
R76854 VSS.n2368 VSS.n2332 0.0105466
R76855 VSS.n2367 VSS.n2333 0.0105466
R76856 VSS.n2331 VSS.n1866 0.0105466
R76857 VSS.n9434 VSS.n9378 0.0105466
R76858 VSS.n9435 VSS.n9377 0.0105466
R76859 VSS.n9376 VSS.n711 0.0105466
R76860 VSS.n2274 VSS.n2171 0.0105466
R76861 VSS.n2273 VSS.n2272 0.0105466
R76862 VSS.n1222 VSS.n1221 0.0105466
R76863 VSS.n1224 VSS.n1168 0.0105466
R76864 VSS.n4716 VSS.n4607 0.0105
R76865 VSS.n4716 VSS.n4715 0.0105
R76866 VSS.n4715 VSS.n4713 0.0105
R76867 VSS.n4713 VSS.n4611 0.0105
R76868 VSS.n4709 VSS.n4611 0.0105
R76869 VSS.n4709 VSS.n4708 0.0105
R76870 VSS.n4708 VSS.n4707 0.0105
R76871 VSS.n4707 VSS.n4617 0.0105
R76872 VSS.n4701 VSS.n4617 0.0105
R76873 VSS.n4701 VSS.n4700 0.0105
R76874 VSS.n4700 VSS.n4698 0.0105
R76875 VSS.n4698 VSS.n4685 0.0105
R76876 VSS.n4694 VSS.n4685 0.0105
R76877 VSS.n4694 VSS.n4693 0.0105
R76878 VSS.n4693 VSS.n4692 0.0105
R76879 VSS.n4692 VSS.n4358 0.0105
R76880 VSS.n5229 VSS.n4358 0.0105
R76881 VSS.n5229 VSS.n5228 0.0105
R76882 VSS.n5228 VSS.n5226 0.0105
R76883 VSS.n5226 VSS.n4362 0.0105
R76884 VSS.n5222 VSS.n4362 0.0105
R76885 VSS.n5222 VSS.n5221 0.0105
R76886 VSS.n5221 VSS.n5220 0.0105
R76887 VSS.n5220 VSS.n4368 0.0105
R76888 VSS.n5216 VSS.n4368 0.0105
R76889 VSS.n5216 VSS.n5215 0.0105
R76890 VSS.n5215 VSS.n5214 0.0105
R76891 VSS.n5214 VSS.n4374 0.0105
R76892 VSS.n5210 VSS.n4374 0.0105
R76893 VSS.n5210 VSS.n5209 0.0105
R76894 VSS.n5209 VSS.n5208 0.0105
R76895 VSS.n5208 VSS.n4380 0.0105
R76896 VSS.n5202 VSS.n4380 0.0105
R76897 VSS.n5202 VSS.n5201 0.0105
R76898 VSS.n5201 VSS.n5199 0.0105
R76899 VSS.n5199 VSS.n4405 0.0105
R76900 VSS.n5195 VSS.n4405 0.0105
R76901 VSS.n5195 VSS.n5194 0.0105
R76902 VSS.n5194 VSS.n5193 0.0105
R76903 VSS.n5193 VSS.n4411 0.0105
R76904 VSS.n5189 VSS.n4411 0.0105
R76905 VSS.n5189 VSS.n5188 0.0105
R76906 VSS.n5188 VSS.n5187 0.0105
R76907 VSS.n5187 VSS.n4417 0.0105
R76908 VSS.n5183 VSS.n4417 0.0105
R76909 VSS.n5183 VSS.n5182 0.0105
R76910 VSS.n5182 VSS.n5181 0.0105
R76911 VSS.n5181 VSS.n4423 0.0105
R76912 VSS.n4441 VSS.n4423 0.0105
R76913 VSS.n5175 VSS.n4441 0.0105
R76914 VSS.n5175 VSS.n5174 0.0105
R76915 VSS.n5174 VSS.n5173 0.0105
R76916 VSS.n5173 VSS.n4447 0.0105
R76917 VSS.n5165 VSS.n4447 0.0105
R76918 VSS.n5165 VSS.n5164 0.0105
R76919 VSS.n5164 VSS.n5163 0.0105
R76920 VSS.n5163 VSS.n5132 0.0105
R76921 VSS.n5159 VSS.n5132 0.0105
R76922 VSS.n5159 VSS.n5158 0.0105
R76923 VSS.n5158 VSS.n5157 0.0105
R76924 VSS.n5157 VSS.n5138 0.0105
R76925 VSS.n5153 VSS.n5138 0.0105
R76926 VSS.n5153 VSS.n5152 0.0105
R76927 VSS.n5152 VSS.n5151 0.0105
R76928 VSS.n5151 VSS.n5148 0.0105
R76929 VSS.n5148 VSS.n5147 0.0105
R76930 VSS.n5147 VSS.n46 0.0105
R76931 VSS.n9887 VSS.n46 0.0105
R76932 VSS.n9887 VSS.n9886 0.0105
R76933 VSS.n9886 VSS.n9884 0.0105
R76934 VSS.n9884 VSS.n50 0.0105
R76935 VSS.n9880 VSS.n50 0.0105
R76936 VSS.n9880 VSS.n9879 0.0105
R76937 VSS.n9879 VSS.n9878 0.0105
R76938 VSS.n9878 VSS.n56 0.0105
R76939 VSS.n9874 VSS.n56 0.0105
R76940 VSS.n9874 VSS.n9873 0.0105
R76941 VSS.n9873 VSS.n9872 0.0105
R76942 VSS.n9872 VSS.n62 0.0105
R76943 VSS.n9868 VSS.n62 0.0105
R76944 VSS.n9868 VSS.n9867 0.0105
R76945 VSS.n9867 VSS.n9866 0.0105
R76946 VSS.n9866 VSS.n68 0.0105
R76947 VSS.n9860 VSS.n68 0.0105
R76948 VSS.n9860 VSS.n9859 0.0105
R76949 VSS.n9859 VSS.n9857 0.0105
R76950 VSS.n9857 VSS.n93 0.0105
R76951 VSS.n9853 VSS.n93 0.0105
R76952 VSS.n9853 VSS.n9852 0.0105
R76953 VSS.n9852 VSS.n9851 0.0105
R76954 VSS.n9851 VSS.n99 0.0105
R76955 VSS.n9845 VSS.n99 0.0105
R76956 VSS.n9845 VSS.n9844 0.0105
R76957 VSS.n9844 VSS.n9842 0.0105
R76958 VSS.n9842 VSS.n124 0.0105
R76959 VSS.n9838 VSS.n124 0.0105
R76960 VSS.n9838 VSS.n9837 0.0105
R76961 VSS.n9836 VSS.n130 0.0105
R76962 VSS.n9828 VSS.n130 0.0105
R76963 VSS.n9828 VSS.n9827 0.0105
R76964 VSS.n4712 VSS.n4711 0.0105
R76965 VSS.n4711 VSS.n4710 0.0105
R76966 VSS.n4710 VSS.n4612 0.0105
R76967 VSS.n4706 VSS.n4612 0.0105
R76968 VSS.n4697 VSS.n4696 0.0105
R76969 VSS.n4696 VSS.n4695 0.0105
R76970 VSS.n4695 VSS.n4686 0.0105
R76971 VSS.n4686 VSS.n4341 0.0105
R76972 VSS.n5225 VSS.n5224 0.0105
R76973 VSS.n5224 VSS.n5223 0.0105
R76974 VSS.n5223 VSS.n4363 0.0105
R76975 VSS.n5219 VSS.n4363 0.0105
R76976 VSS.n5219 VSS.n5218 0.0105
R76977 VSS.n5218 VSS.n5217 0.0105
R76978 VSS.n5217 VSS.n4369 0.0105
R76979 VSS.n5213 VSS.n4369 0.0105
R76980 VSS.n5213 VSS.n5212 0.0105
R76981 VSS.n5212 VSS.n5211 0.0105
R76982 VSS.n5211 VSS.n4375 0.0105
R76983 VSS.n5207 VSS.n4375 0.0105
R76984 VSS.n5198 VSS.n5197 0.0105
R76985 VSS.n5197 VSS.n5196 0.0105
R76986 VSS.n5196 VSS.n4406 0.0105
R76987 VSS.n5192 VSS.n4406 0.0105
R76988 VSS.n5192 VSS.n5191 0.0105
R76989 VSS.n5191 VSS.n5190 0.0105
R76990 VSS.n5190 VSS.n4412 0.0105
R76991 VSS.n5186 VSS.n4412 0.0105
R76992 VSS.n5186 VSS.n5185 0.0105
R76993 VSS.n5185 VSS.n5184 0.0105
R76994 VSS.n5184 VSS.n4418 0.0105
R76995 VSS.n5180 VSS.n4418 0.0105
R76996 VSS.n5176 VSS.n4440 0.0105
R76997 VSS.n5166 VSS.n5127 0.0105
R76998 VSS.n5162 VSS.n5127 0.0105
R76999 VSS.n5162 VSS.n5161 0.0105
R77000 VSS.n5161 VSS.n5160 0.0105
R77001 VSS.n5160 VSS.n5133 0.0105
R77002 VSS.n5156 VSS.n5133 0.0105
R77003 VSS.n5156 VSS.n5155 0.0105
R77004 VSS.n5155 VSS.n5154 0.0105
R77005 VSS.n5154 VSS.n5139 0.0105
R77006 VSS.n5150 VSS.n5139 0.0105
R77007 VSS.n5150 VSS.n5149 0.0105
R77008 VSS.n5149 VSS.n35 0.0105
R77009 VSS.n9883 VSS.n9882 0.0105
R77010 VSS.n9882 VSS.n9881 0.0105
R77011 VSS.n9881 VSS.n51 0.0105
R77012 VSS.n9877 VSS.n51 0.0105
R77013 VSS.n9877 VSS.n9876 0.0105
R77014 VSS.n9876 VSS.n9875 0.0105
R77015 VSS.n9875 VSS.n57 0.0105
R77016 VSS.n9871 VSS.n57 0.0105
R77017 VSS.n9871 VSS.n9870 0.0105
R77018 VSS.n9870 VSS.n9869 0.0105
R77019 VSS.n9869 VSS.n63 0.0105
R77020 VSS.n9865 VSS.n63 0.0105
R77021 VSS.n9856 VSS.n9855 0.0105
R77022 VSS.n9855 VSS.n9854 0.0105
R77023 VSS.n9854 VSS.n94 0.0105
R77024 VSS.n9850 VSS.n94 0.0105
R77025 VSS.n9841 VSS.n9840 0.0105
R77026 VSS.n9840 VSS.n9839 0.0105
R77027 VSS.n9839 VSS.n125 0.0105
R77028 VSS.n4858 VSS.n4852 0.0104296
R77029 VSS.n3732 VSS.n3144 0.0104296
R77030 VSS.n6781 VSS.n2950 0.0104296
R77031 VSS.n4862 VSS.n4498 0.0104296
R77032 VSS.n3775 VSS.n3174 0.0104296
R77033 VSS.n6782 VSS.n2932 0.0104296
R77034 VSS.n83 VSS.n73 0.0102441
R77035 VSS.n2279 VSS.n2155 0.0102441
R77036 VSS.n2385 VSS.n1860 0.0102441
R77037 VSS.n4675 VSS.n4622 0.0102441
R77038 VSS.n30 VSS.n20 0.0102441
R77039 VSS.n4395 VSS.n4385 0.0102441
R77040 VSS.n4355 VSS.n4345 0.0102441
R77041 VSS.n4604 VSS.n4594 0.0102441
R77042 VSS.n6262 VSS.n6261 0.0102441
R77043 VSS.n9821 VSS.n135 0.0102441
R77044 VSS.n4149 VSS.n421 0.0102441
R77045 VSS.n114 VSS.n104 0.0102441
R77046 VSS.n1217 VSS.n743 0.0102441
R77047 VSS.n9417 VSS.n706 0.0102441
R77048 VSS.n4857 VSS.n4856 0.010007
R77049 VSS.n3734 VSS.n3154 0.010007
R77050 VSS.n6775 VSS.n2947 0.010007
R77051 VSS.n4500 VSS.n4492 0.010007
R77052 VSS.n3771 VSS.n3184 0.010007
R77053 VSS.n6776 VSS.n2929 0.010007
R77054 VSS.n161 VSS.n73 0.00988976
R77055 VSS.n4132 VSS.n355 0.00988976
R77056 VSS.n4163 VSS.n347 0.00988976
R77057 VSS.n4134 VSS.n356 0.00988976
R77058 VSS.n4138 VSS.n346 0.00988976
R77059 VSS.n9645 VSS.n357 0.00988976
R77060 VSS.n2281 VSS.n2155 0.00988976
R77061 VSS.n2383 VSS.n1860 0.00988976
R77062 VSS.n4672 VSS.n4622 0.00988976
R77063 VSS.n9894 VSS.n30 0.00988976
R77064 VSS.n4124 VSS.n322 0.00988976
R77065 VSS.n4167 VSS.n313 0.00988976
R77066 VSS.n4126 VSS.n323 0.00988976
R77067 VSS.n4130 VSS.n312 0.00988976
R77068 VSS.n9679 VSS.n324 0.00988976
R77069 VSS.n4664 VSS.n4385 0.00988976
R77070 VSS.n4080 VSS.n3993 0.00988976
R77071 VSS.n4109 VSS.n3982 0.00988976
R77072 VSS.n4082 VSS.n3994 0.00988976
R77073 VSS.n4105 VSS.n3981 0.00988976
R77074 VSS.n6160 VSS.n3995 0.00988976
R77075 VSS.n4668 VSS.n4345 0.00988976
R77076 VSS.n4084 VSS.n3948 0.00988976
R77077 VSS.n4101 VSS.n3940 0.00988976
R77078 VSS.n4086 VSS.n3949 0.00988976
R77079 VSS.n4097 VSS.n3939 0.00988976
R77080 VSS.n6196 VSS.n3950 0.00988976
R77081 VSS.n4638 VSS.n4594 0.00988976
R77082 VSS.n6262 VSS.n3852 0.00988976
R77083 VSS.n9817 VSS.n135 0.00988976
R77084 VSS.n4150 VSS.n421 0.00988976
R77085 VSS.n165 VSS.n104 0.00988976
R77086 VSS.n4140 VSS.n394 0.00988976
R77087 VSS.n4160 VSS.n383 0.00988976
R77088 VSS.n4142 VSS.n395 0.00988976
R77089 VSS.n4146 VSS.n382 0.00988976
R77090 VSS.n9627 VSS.n396 0.00988976
R77091 VSS.n1215 VSS.n743 0.00988976
R77092 VSS.n9419 VSS.n706 0.00988976
R77093 VSS.n5180 VSS.n5179 0.00979577
R77094 VSS.n7305 VSS.n7301 0.00962857
R77095 VSS.n7305 VSS.n7299 0.00962857
R77096 VSS.n7309 VSS.n7299 0.00962857
R77097 VSS.n7309 VSS.n7297 0.00962857
R77098 VSS.n7313 VSS.n7297 0.00962857
R77099 VSS.n7313 VSS.n7295 0.00962857
R77100 VSS.n7317 VSS.n7295 0.00962857
R77101 VSS.n7317 VSS.n7293 0.00962857
R77102 VSS.n7321 VSS.n7293 0.00962857
R77103 VSS.n7321 VSS.n7290 0.00962857
R77104 VSS.n7593 VSS.n7290 0.00962857
R77105 VSS.n7593 VSS.n7291 0.00962857
R77106 VSS.n7589 VSS.n7291 0.00962857
R77107 VSS.n7589 VSS.n7325 0.00962857
R77108 VSS.n7585 VSS.n7325 0.00962857
R77109 VSS.n7585 VSS.n7327 0.00962857
R77110 VSS.n7581 VSS.n7327 0.00962857
R77111 VSS.n7581 VSS.n7329 0.00962857
R77112 VSS.n7577 VSS.n7329 0.00962857
R77113 VSS.n7577 VSS.n7331 0.00962857
R77114 VSS.n7573 VSS.n7331 0.00962857
R77115 VSS.n7573 VSS.n7333 0.00962857
R77116 VSS.n7569 VSS.n7333 0.00962857
R77117 VSS.n7569 VSS.n7335 0.00962857
R77118 VSS.n7565 VSS.n7335 0.00962857
R77119 VSS.n7565 VSS.n7337 0.00962857
R77120 VSS.n7561 VSS.n7337 0.00962857
R77121 VSS.n7561 VSS.n7339 0.00962857
R77122 VSS.n7557 VSS.n7339 0.00962857
R77123 VSS.n7557 VSS.n7341 0.00962857
R77124 VSS.n7553 VSS.n7341 0.00962857
R77125 VSS.n7553 VSS.n7343 0.00962857
R77126 VSS.n7549 VSS.n7343 0.00962857
R77127 VSS.n7549 VSS.n7345 0.00962857
R77128 VSS.n7545 VSS.n7345 0.00962857
R77129 VSS.n7545 VSS.n7347 0.00962857
R77130 VSS.n7541 VSS.n7347 0.00962857
R77131 VSS.n7541 VSS.n7349 0.00962857
R77132 VSS.n7537 VSS.n7349 0.00962857
R77133 VSS.n7537 VSS.n7351 0.00962857
R77134 VSS.n7533 VSS.n7351 0.00962857
R77135 VSS.n7533 VSS.n7353 0.00962857
R77136 VSS.n7529 VSS.n7353 0.00962857
R77137 VSS.n7529 VSS.n7355 0.00962857
R77138 VSS.n7525 VSS.n7355 0.00962857
R77139 VSS.n7525 VSS.n7357 0.00962857
R77140 VSS.n7521 VSS.n7357 0.00962857
R77141 VSS.n7521 VSS.n7359 0.00962857
R77142 VSS.n7517 VSS.n7359 0.00962857
R77143 VSS.n7517 VSS.n7361 0.00962857
R77144 VSS.n7513 VSS.n7361 0.00962857
R77145 VSS.n7513 VSS.n7363 0.00962857
R77146 VSS.n7509 VSS.n7363 0.00962857
R77147 VSS.n7509 VSS.n7365 0.00962857
R77148 VSS.n7505 VSS.n7365 0.00962857
R77149 VSS.n7505 VSS.n7367 0.00962857
R77150 VSS.n7501 VSS.n7367 0.00962857
R77151 VSS.n7501 VSS.n7369 0.00962857
R77152 VSS.n7497 VSS.n7369 0.00962857
R77153 VSS.n7497 VSS.n7371 0.00962857
R77154 VSS.n7493 VSS.n7371 0.00962857
R77155 VSS.n7493 VSS.n7373 0.00962857
R77156 VSS.n7489 VSS.n7373 0.00962857
R77157 VSS.n7489 VSS.n7375 0.00962857
R77158 VSS.n7485 VSS.n7375 0.00962857
R77159 VSS.n7485 VSS.n7377 0.00962857
R77160 VSS.n7481 VSS.n7377 0.00962857
R77161 VSS.n7481 VSS.n7379 0.00962857
R77162 VSS.n7477 VSS.n7379 0.00962857
R77163 VSS.n7477 VSS.n7381 0.00962857
R77164 VSS.n7473 VSS.n7381 0.00962857
R77165 VSS.n7473 VSS.n7383 0.00962857
R77166 VSS.n7469 VSS.n7383 0.00962857
R77167 VSS.n7469 VSS.n7385 0.00962857
R77168 VSS.n7465 VSS.n7385 0.00962857
R77169 VSS.n7465 VSS.n7387 0.00962857
R77170 VSS.n7461 VSS.n7387 0.00962857
R77171 VSS.n7461 VSS.n7389 0.00962857
R77172 VSS.n7457 VSS.n7389 0.00962857
R77173 VSS.n7457 VSS.n7391 0.00962857
R77174 VSS.n7453 VSS.n7391 0.00962857
R77175 VSS.n7453 VSS.n7393 0.00962857
R77176 VSS.n7449 VSS.n7393 0.00962857
R77177 VSS.n7449 VSS.n7395 0.00962857
R77178 VSS.n7445 VSS.n7395 0.00962857
R77179 VSS.n7445 VSS.n7397 0.00962857
R77180 VSS.n7441 VSS.n7397 0.00962857
R77181 VSS.n7441 VSS.n7399 0.00962857
R77182 VSS.n7437 VSS.n7399 0.00962857
R77183 VSS.n7437 VSS.n7401 0.00962857
R77184 VSS.n7433 VSS.n7401 0.00962857
R77185 VSS.n7433 VSS.n7403 0.00962857
R77186 VSS.n7429 VSS.n7403 0.00962857
R77187 VSS.n7429 VSS.n7405 0.00962857
R77188 VSS.n7425 VSS.n7405 0.00962857
R77189 VSS.n7425 VSS.n7407 0.00962857
R77190 VSS.n7421 VSS.n7407 0.00962857
R77191 VSS.n7418 VSS.n7417 0.00962857
R77192 VSS.n7417 VSS.n7410 0.00962857
R77193 VSS.n7413 VSS.n7410 0.00962857
R77194 VSS.n4736 VSS.n4583 0.00962857
R77195 VSS.n4766 VSS.n4583 0.00962857
R77196 VSS.n4766 VSS.n4581 0.00962857
R77197 VSS.n4770 VSS.n4581 0.00962857
R77198 VSS.n4770 VSS.n4579 0.00962857
R77199 VSS.n4774 VSS.n4579 0.00962857
R77200 VSS.n4774 VSS.n4577 0.00962857
R77201 VSS.n4778 VSS.n4577 0.00962857
R77202 VSS.n4778 VSS.n4551 0.00962857
R77203 VSS.n4788 VSS.n4551 0.00962857
R77204 VSS.n4788 VSS.n4549 0.00962857
R77205 VSS.n4792 VSS.n4549 0.00962857
R77206 VSS.n4792 VSS.n4547 0.00962857
R77207 VSS.n4796 VSS.n4547 0.00962857
R77208 VSS.n4796 VSS.n4545 0.00962857
R77209 VSS.n4800 VSS.n4545 0.00962857
R77210 VSS.n4802 VSS.n4800 0.00962857
R77211 VSS.n4804 VSS.n4802 0.00962857
R77212 VSS.n4804 VSS.n4543 0.00962857
R77213 VSS.n4808 VSS.n4543 0.00962857
R77214 VSS.n4808 VSS.n4541 0.00962857
R77215 VSS.n4812 VSS.n4541 0.00962857
R77216 VSS.n4812 VSS.n4539 0.00962857
R77217 VSS.n4816 VSS.n4539 0.00962857
R77218 VSS.n4816 VSS.n4537 0.00962857
R77219 VSS.n4820 VSS.n4537 0.00962857
R77220 VSS.n4820 VSS.n4535 0.00962857
R77221 VSS.n4824 VSS.n4535 0.00962857
R77222 VSS.n4824 VSS.n4533 0.00962857
R77223 VSS.n4828 VSS.n4533 0.00962857
R77224 VSS.n4828 VSS.n4529 0.00962857
R77225 VSS.n5059 VSS.n4529 0.00962857
R77226 VSS.n5059 VSS.n4531 0.00962857
R77227 VSS.n5055 VSS.n4531 0.00962857
R77228 VSS.n5055 VSS.n5053 0.00962857
R77229 VSS.n5053 VSS.n4832 0.00962857
R77230 VSS.n5049 VSS.n4832 0.00962857
R77231 VSS.n5049 VSS.n4834 0.00962857
R77232 VSS.n5045 VSS.n4834 0.00962857
R77233 VSS.n5045 VSS.n4837 0.00962857
R77234 VSS.n5041 VSS.n4837 0.00962857
R77235 VSS.n5041 VSS.n4839 0.00962857
R77236 VSS.n5037 VSS.n4839 0.00962857
R77237 VSS.n5037 VSS.n4841 0.00962857
R77238 VSS.n5033 VSS.n4841 0.00962857
R77239 VSS.n5033 VSS.n4843 0.00962857
R77240 VSS.n5029 VSS.n4843 0.00962857
R77241 VSS.n5029 VSS.n5028 0.00962857
R77242 VSS.n5028 VSS.n5027 0.00962857
R77243 VSS.n5027 VSS.n4845 0.00962857
R77244 VSS.n5022 VSS.n4845 0.00962857
R77245 VSS.n5022 VSS.n4847 0.00962857
R77246 VSS.n4977 VSS.n4847 0.00962857
R77247 VSS.n5016 VSS.n4977 0.00962857
R77248 VSS.n5016 VSS.n4978 0.00962857
R77249 VSS.n5012 VSS.n4978 0.00962857
R77250 VSS.n5012 VSS.n4981 0.00962857
R77251 VSS.n5008 VSS.n4981 0.00962857
R77252 VSS.n5008 VSS.n4983 0.00962857
R77253 VSS.n5004 VSS.n4983 0.00962857
R77254 VSS.n5004 VSS.n4985 0.00962857
R77255 VSS.n5000 VSS.n4985 0.00962857
R77256 VSS.n5000 VSS.n4987 0.00962857
R77257 VSS.n4996 VSS.n4987 0.00962857
R77258 VSS.n4996 VSS.n4993 0.00962857
R77259 VSS.n4993 VSS.n4992 0.00962857
R77260 VSS.n4992 VSS.n4989 0.00962857
R77261 VSS.n4989 VSS.n249 0.00962857
R77262 VSS.n9698 VSS.n249 0.00962857
R77263 VSS.n9698 VSS.n247 0.00962857
R77264 VSS.n9702 VSS.n247 0.00962857
R77265 VSS.n9702 VSS.n245 0.00962857
R77266 VSS.n9706 VSS.n245 0.00962857
R77267 VSS.n9706 VSS.n243 0.00962857
R77268 VSS.n9710 VSS.n243 0.00962857
R77269 VSS.n9710 VSS.n241 0.00962857
R77270 VSS.n9714 VSS.n241 0.00962857
R77271 VSS.n9714 VSS.n239 0.00962857
R77272 VSS.n9718 VSS.n239 0.00962857
R77273 VSS.n9718 VSS.n237 0.00962857
R77274 VSS.n9722 VSS.n237 0.00962857
R77275 VSS.n9722 VSS.n233 0.00962857
R77276 VSS.n9746 VSS.n233 0.00962857
R77277 VSS.n9746 VSS.n235 0.00962857
R77278 VSS.n9742 VSS.n235 0.00962857
R77279 VSS.n9742 VSS.n9740 0.00962857
R77280 VSS.n9740 VSS.n9726 0.00962857
R77281 VSS.n9736 VSS.n9726 0.00962857
R77282 VSS.n9736 VSS.n9728 0.00962857
R77283 VSS.n9732 VSS.n9728 0.00962857
R77284 VSS.n9732 VSS.n9731 0.00962857
R77285 VSS.n9731 VSS.n193 0.00962857
R77286 VSS.n9780 VSS.n193 0.00962857
R77287 VSS.n9780 VSS.n191 0.00962857
R77288 VSS.n9784 VSS.n191 0.00962857
R77289 VSS.n9784 VSS.n189 0.00962857
R77290 VSS.n9788 VSS.n189 0.00962857
R77291 VSS.n9796 VSS.n185 0.00962857
R77292 VSS.n9796 VSS.n187 0.00962857
R77293 VSS.n9792 VSS.n187 0.00962857
R77294 VSS.n8286 VSS.n1705 0.00962857
R77295 VSS.n8303 VSS.n1705 0.00962857
R77296 VSS.n8303 VSS.n1703 0.00962857
R77297 VSS.n8307 VSS.n1703 0.00962857
R77298 VSS.n8307 VSS.n1701 0.00962857
R77299 VSS.n8311 VSS.n1701 0.00962857
R77300 VSS.n8311 VSS.n1699 0.00962857
R77301 VSS.n8315 VSS.n1699 0.00962857
R77302 VSS.n8315 VSS.n1685 0.00962857
R77303 VSS.n8332 VSS.n1685 0.00962857
R77304 VSS.n8332 VSS.n1683 0.00962857
R77305 VSS.n8336 VSS.n1683 0.00962857
R77306 VSS.n8336 VSS.n1681 0.00962857
R77307 VSS.n8340 VSS.n1681 0.00962857
R77308 VSS.n8340 VSS.n1679 0.00962857
R77309 VSS.n8344 VSS.n1679 0.00962857
R77310 VSS.n8346 VSS.n8344 0.00962857
R77311 VSS.n8348 VSS.n8346 0.00962857
R77312 VSS.n8348 VSS.n1677 0.00962857
R77313 VSS.n8352 VSS.n1677 0.00962857
R77314 VSS.n8352 VSS.n1675 0.00962857
R77315 VSS.n8356 VSS.n1675 0.00962857
R77316 VSS.n8356 VSS.n1673 0.00962857
R77317 VSS.n8360 VSS.n1673 0.00962857
R77318 VSS.n8360 VSS.n1671 0.00962857
R77319 VSS.n8364 VSS.n1671 0.00962857
R77320 VSS.n8364 VSS.n1669 0.00962857
R77321 VSS.n8368 VSS.n1669 0.00962857
R77322 VSS.n8368 VSS.n1667 0.00962857
R77323 VSS.n8373 VSS.n1667 0.00962857
R77324 VSS.n8373 VSS.n1665 0.00962857
R77325 VSS.n8377 VSS.n1665 0.00962857
R77326 VSS.n8377 VSS.n1654 0.00962857
R77327 VSS.n8414 VSS.n1654 0.00962857
R77328 VSS.n8414 VSS.n1652 0.00962857
R77329 VSS.n8418 VSS.n1652 0.00962857
R77330 VSS.n8418 VSS.n1650 0.00962857
R77331 VSS.n8422 VSS.n1650 0.00962857
R77332 VSS.n8422 VSS.n1648 0.00962857
R77333 VSS.n8426 VSS.n1648 0.00962857
R77334 VSS.n8426 VSS.n1646 0.00962857
R77335 VSS.n8430 VSS.n1646 0.00962857
R77336 VSS.n8430 VSS.n1644 0.00962857
R77337 VSS.n8435 VSS.n1644 0.00962857
R77338 VSS.n8435 VSS.n1641 0.00962857
R77339 VSS.n8439 VSS.n1641 0.00962857
R77340 VSS.n8440 VSS.n8439 0.00962857
R77341 VSS.n8441 VSS.n8440 0.00962857
R77342 VSS.n8441 VSS.n1638 0.00962857
R77343 VSS.n8533 VSS.n1638 0.00962857
R77344 VSS.n8533 VSS.n1639 0.00962857
R77345 VSS.n8529 VSS.n1639 0.00962857
R77346 VSS.n8529 VSS.n8528 0.00962857
R77347 VSS.n8528 VSS.n8527 0.00962857
R77348 VSS.n8527 VSS.n8445 0.00962857
R77349 VSS.n8523 VSS.n8445 0.00962857
R77350 VSS.n8523 VSS.n8447 0.00962857
R77351 VSS.n8519 VSS.n8447 0.00962857
R77352 VSS.n8519 VSS.n8450 0.00962857
R77353 VSS.n8515 VSS.n8450 0.00962857
R77354 VSS.n8515 VSS.n8452 0.00962857
R77355 VSS.n8511 VSS.n8452 0.00962857
R77356 VSS.n8511 VSS.n8454 0.00962857
R77357 VSS.n8507 VSS.n8454 0.00962857
R77358 VSS.n8507 VSS.n8504 0.00962857
R77359 VSS.n8504 VSS.n8503 0.00962857
R77360 VSS.n8503 VSS.n8456 0.00962857
R77361 VSS.n8499 VSS.n8456 0.00962857
R77362 VSS.n8499 VSS.n8497 0.00962857
R77363 VSS.n8497 VSS.n8495 0.00962857
R77364 VSS.n8495 VSS.n8458 0.00962857
R77365 VSS.n8491 VSS.n8458 0.00962857
R77366 VSS.n8491 VSS.n8461 0.00962857
R77367 VSS.n8487 VSS.n8461 0.00962857
R77368 VSS.n8487 VSS.n8464 0.00962857
R77369 VSS.n8483 VSS.n8464 0.00962857
R77370 VSS.n8483 VSS.n8466 0.00962857
R77371 VSS.n8479 VSS.n8466 0.00962857
R77372 VSS.n8479 VSS.n8468 0.00962857
R77373 VSS.n8475 VSS.n8468 0.00962857
R77374 VSS.n8475 VSS.n8470 0.00962857
R77375 VSS.n8471 VSS.n8470 0.00962857
R77376 VSS.n8471 VSS.n1287 0.00962857
R77377 VSS.n8863 VSS.n1287 0.00962857
R77378 VSS.n8863 VSS.n1285 0.00962857
R77379 VSS.n8867 VSS.n1285 0.00962857
R77380 VSS.n8867 VSS.n1283 0.00962857
R77381 VSS.n8872 VSS.n1283 0.00962857
R77382 VSS.n8872 VSS.n1281 0.00962857
R77383 VSS.n8876 VSS.n1281 0.00962857
R77384 VSS.n8877 VSS.n8876 0.00962857
R77385 VSS.n8879 VSS.n8877 0.00962857
R77386 VSS.n8879 VSS.n1278 0.00962857
R77387 VSS.n8900 VSS.n1278 0.00962857
R77388 VSS.n8900 VSS.n1279 0.00962857
R77389 VSS.n8896 VSS.n1279 0.00962857
R77390 VSS.n8896 VSS.n8893 0.00962857
R77391 VSS.n8892 VSS.n8883 0.00962857
R77392 VSS.n8888 VSS.n8883 0.00962857
R77393 VSS.n8888 VSS.n8886 0.00962857
R77394 VSS.n8308 VSS.n1702 0.00962857
R77395 VSS.n8309 VSS.n8308 0.00962857
R77396 VSS.n8310 VSS.n8309 0.00962857
R77397 VSS.n8310 VSS.n1694 0.00962857
R77398 VSS.n8337 VSS.n1682 0.00962857
R77399 VSS.n8338 VSS.n8337 0.00962857
R77400 VSS.n8339 VSS.n8338 0.00962857
R77401 VSS.n8339 VSS.n1571 0.00962857
R77402 VSS.n8353 VSS.n1676 0.00962857
R77403 VSS.n8354 VSS.n8353 0.00962857
R77404 VSS.n8355 VSS.n8354 0.00962857
R77405 VSS.n8355 VSS.n1672 0.00962857
R77406 VSS.n8361 VSS.n1672 0.00962857
R77407 VSS.n8362 VSS.n8361 0.00962857
R77408 VSS.n8363 VSS.n8362 0.00962857
R77409 VSS.n8363 VSS.n1668 0.00962857
R77410 VSS.n8369 VSS.n1668 0.00962857
R77411 VSS.n8370 VSS.n8369 0.00962857
R77412 VSS.n8372 VSS.n8370 0.00962857
R77413 VSS.n8372 VSS.n8371 0.00962857
R77414 VSS.n8419 VSS.n1651 0.00962857
R77415 VSS.n8420 VSS.n8419 0.00962857
R77416 VSS.n8421 VSS.n8420 0.00962857
R77417 VSS.n8421 VSS.n1647 0.00962857
R77418 VSS.n8427 VSS.n1647 0.00962857
R77419 VSS.n8428 VSS.n8427 0.00962857
R77420 VSS.n8429 VSS.n8428 0.00962857
R77421 VSS.n8429 VSS.n1643 0.00962857
R77422 VSS.n8436 VSS.n1643 0.00962857
R77423 VSS.n8437 VSS.n8436 0.00962857
R77424 VSS.n8438 VSS.n8437 0.00962857
R77425 VSS.n8438 VSS.n1619 0.00962857
R77426 VSS.n8534 VSS.n1637 0.00962857
R77427 VSS.n8448 VSS.n1376 0.00962857
R77428 VSS.n8522 VSS.n8448 0.00962857
R77429 VSS.n8522 VSS.n8521 0.00962857
R77430 VSS.n8521 VSS.n8520 0.00962857
R77431 VSS.n8520 VSS.n8449 0.00962857
R77432 VSS.n8514 VSS.n8449 0.00962857
R77433 VSS.n8514 VSS.n8513 0.00962857
R77434 VSS.n8513 VSS.n8512 0.00962857
R77435 VSS.n8512 VSS.n8453 0.00962857
R77436 VSS.n8506 VSS.n8453 0.00962857
R77437 VSS.n8506 VSS.n8505 0.00962857
R77438 VSS.n8505 VSS.n1325 0.00962857
R77439 VSS.n8494 VSS.n8493 0.00962857
R77440 VSS.n8493 VSS.n8492 0.00962857
R77441 VSS.n8492 VSS.n8460 0.00962857
R77442 VSS.n8486 VSS.n8460 0.00962857
R77443 VSS.n8486 VSS.n8485 0.00962857
R77444 VSS.n8485 VSS.n8484 0.00962857
R77445 VSS.n8484 VSS.n8465 0.00962857
R77446 VSS.n8478 VSS.n8465 0.00962857
R77447 VSS.n8478 VSS.n8477 0.00962857
R77448 VSS.n8477 VSS.n8476 0.00962857
R77449 VSS.n8476 VSS.n8469 0.00962857
R77450 VSS.n8469 VSS.n1306 0.00962857
R77451 VSS.n8869 VSS.n8868 0.00962857
R77452 VSS.n8871 VSS.n8869 0.00962857
R77453 VSS.n8871 VSS.n8870 0.00962857
R77454 VSS.n8870 VSS.n1261 0.00962857
R77455 VSS.n8901 VSS.n1277 0.00962857
R77456 VSS.n8895 VSS.n1277 0.00962857
R77457 VSS.n8895 VSS.n8894 0.00962857
R77458 VSS.n2820 VSS.n2818 0.00962857
R77459 VSS.n2820 VSS.n2816 0.00962857
R77460 VSS.n6955 VSS.n2816 0.00962857
R77461 VSS.n6955 VSS.n2817 0.00962857
R77462 VSS.n6951 VSS.n2817 0.00962857
R77463 VSS.n6951 VSS.n2824 0.00962857
R77464 VSS.n6947 VSS.n2824 0.00962857
R77465 VSS.n6947 VSS.n2826 0.00962857
R77466 VSS.n6943 VSS.n2826 0.00962857
R77467 VSS.n6943 VSS.n2828 0.00962857
R77468 VSS.n6932 VSS.n2828 0.00962857
R77469 VSS.n6932 VSS.n2848 0.00962857
R77470 VSS.n6928 VSS.n2848 0.00962857
R77471 VSS.n6928 VSS.n2850 0.00962857
R77472 VSS.n6924 VSS.n2850 0.00962857
R77473 VSS.n6924 VSS.n2852 0.00962857
R77474 VSS.n6920 VSS.n2852 0.00962857
R77475 VSS.n6920 VSS.n2854 0.00962857
R77476 VSS.n6909 VSS.n2854 0.00962857
R77477 VSS.n6909 VSS.n2874 0.00962857
R77478 VSS.n6905 VSS.n2874 0.00962857
R77479 VSS.n6905 VSS.n2876 0.00962857
R77480 VSS.n6901 VSS.n2876 0.00962857
R77481 VSS.n6901 VSS.n2878 0.00962857
R77482 VSS.n6897 VSS.n2878 0.00962857
R77483 VSS.n6897 VSS.n2880 0.00962857
R77484 VSS.n6893 VSS.n2880 0.00962857
R77485 VSS.n6893 VSS.n2882 0.00962857
R77486 VSS.n6889 VSS.n2882 0.00962857
R77487 VSS.n6889 VSS.n2884 0.00962857
R77488 VSS.n6885 VSS.n2884 0.00962857
R77489 VSS.n6885 VSS.n2886 0.00962857
R77490 VSS.n6881 VSS.n2886 0.00962857
R77491 VSS.n6881 VSS.n2888 0.00962857
R77492 VSS.n6870 VSS.n2888 0.00962857
R77493 VSS.n6870 VSS.n2908 0.00962857
R77494 VSS.n6866 VSS.n2908 0.00962857
R77495 VSS.n6866 VSS.n2910 0.00962857
R77496 VSS.n6862 VSS.n2910 0.00962857
R77497 VSS.n6862 VSS.n2912 0.00962857
R77498 VSS.n6858 VSS.n2912 0.00962857
R77499 VSS.n6858 VSS.n2914 0.00962857
R77500 VSS.n6854 VSS.n2914 0.00962857
R77501 VSS.n6854 VSS.n2916 0.00962857
R77502 VSS.n6850 VSS.n2916 0.00962857
R77503 VSS.n6850 VSS.n2918 0.00962857
R77504 VSS.n6846 VSS.n2918 0.00962857
R77505 VSS.n6846 VSS.n2920 0.00962857
R77506 VSS.n6842 VSS.n2920 0.00962857
R77507 VSS.n6842 VSS.n2922 0.00962857
R77508 VSS.n3012 VSS.n2922 0.00962857
R77509 VSS.n3013 VSS.n3012 0.00962857
R77510 VSS.n3015 VSS.n3013 0.00962857
R77511 VSS.n3015 VSS.n3009 0.00962857
R77512 VSS.n3019 VSS.n3009 0.00962857
R77513 VSS.n3019 VSS.n3007 0.00962857
R77514 VSS.n3023 VSS.n3007 0.00962857
R77515 VSS.n3023 VSS.n3005 0.00962857
R77516 VSS.n3027 VSS.n3005 0.00962857
R77517 VSS.n3027 VSS.n3003 0.00962857
R77518 VSS.n3031 VSS.n3003 0.00962857
R77519 VSS.n3031 VSS.n3001 0.00962857
R77520 VSS.n3036 VSS.n3001 0.00962857
R77521 VSS.n3036 VSS.n2999 0.00962857
R77522 VSS.n3040 VSS.n2999 0.00962857
R77523 VSS.n3041 VSS.n3040 0.00962857
R77524 VSS.n3041 VSS.n2995 0.00962857
R77525 VSS.n6747 VSS.n2995 0.00962857
R77526 VSS.n6747 VSS.n2997 0.00962857
R77527 VSS.n6743 VSS.n2997 0.00962857
R77528 VSS.n6743 VSS.n3045 0.00962857
R77529 VSS.n6739 VSS.n3045 0.00962857
R77530 VSS.n6739 VSS.n3047 0.00962857
R77531 VSS.n6735 VSS.n3047 0.00962857
R77532 VSS.n6735 VSS.n3049 0.00962857
R77533 VSS.n6731 VSS.n3049 0.00962857
R77534 VSS.n6731 VSS.n3051 0.00962857
R77535 VSS.n6727 VSS.n3051 0.00962857
R77536 VSS.n6727 VSS.n3053 0.00962857
R77537 VSS.n6723 VSS.n3053 0.00962857
R77538 VSS.n6723 VSS.n3055 0.00962857
R77539 VSS.n6719 VSS.n3055 0.00962857
R77540 VSS.n6719 VSS.n3057 0.00962857
R77541 VSS.n3082 VSS.n3057 0.00962857
R77542 VSS.n6713 VSS.n3082 0.00962857
R77543 VSS.n6713 VSS.n3083 0.00962857
R77544 VSS.n6709 VSS.n3083 0.00962857
R77545 VSS.n6709 VSS.n3086 0.00962857
R77546 VSS.n6705 VSS.n3086 0.00962857
R77547 VSS.n6705 VSS.n3089 0.00962857
R77548 VSS.n6701 VSS.n3089 0.00962857
R77549 VSS.n6701 VSS.n3091 0.00962857
R77550 VSS.n6668 VSS.n3091 0.00962857
R77551 VSS.n6689 VSS.n6668 0.00962857
R77552 VSS.n6689 VSS.n6669 0.00962857
R77553 VSS.n6685 VSS.n6669 0.00962857
R77554 VSS.n6685 VSS.n6682 0.00962857
R77555 VSS.n6681 VSS.n6672 0.00962857
R77556 VSS.n6677 VSS.n6672 0.00962857
R77557 VSS.n6677 VSS.n6675 0.00962857
R77558 VSS.n6956 VSS.n2815 0.00962857
R77559 VSS.n6950 VSS.n2815 0.00962857
R77560 VSS.n6950 VSS.n6949 0.00962857
R77561 VSS.n6949 VSS.n6948 0.00962857
R77562 VSS.n6933 VSS.n2847 0.00962857
R77563 VSS.n6927 VSS.n2847 0.00962857
R77564 VSS.n6927 VSS.n6926 0.00962857
R77565 VSS.n6926 VSS.n6925 0.00962857
R77566 VSS.n6910 VSS.n2873 0.00962857
R77567 VSS.n6904 VSS.n2873 0.00962857
R77568 VSS.n6904 VSS.n6903 0.00962857
R77569 VSS.n6903 VSS.n6902 0.00962857
R77570 VSS.n6902 VSS.n2877 0.00962857
R77571 VSS.n6896 VSS.n2877 0.00962857
R77572 VSS.n6896 VSS.n6895 0.00962857
R77573 VSS.n6895 VSS.n6894 0.00962857
R77574 VSS.n6894 VSS.n2881 0.00962857
R77575 VSS.n6888 VSS.n2881 0.00962857
R77576 VSS.n6888 VSS.n6887 0.00962857
R77577 VSS.n6887 VSS.n6886 0.00962857
R77578 VSS.n6871 VSS.n2907 0.00962857
R77579 VSS.n6865 VSS.n2907 0.00962857
R77580 VSS.n6865 VSS.n6864 0.00962857
R77581 VSS.n6864 VSS.n6863 0.00962857
R77582 VSS.n6863 VSS.n2911 0.00962857
R77583 VSS.n6857 VSS.n2911 0.00962857
R77584 VSS.n6857 VSS.n6856 0.00962857
R77585 VSS.n6856 VSS.n6855 0.00962857
R77586 VSS.n6855 VSS.n2915 0.00962857
R77587 VSS.n6849 VSS.n2915 0.00962857
R77588 VSS.n6849 VSS.n6848 0.00962857
R77589 VSS.n6848 VSS.n6847 0.00962857
R77590 VSS.n2942 VSS.n2930 0.00962857
R77591 VSS.n3020 VSS.n3008 0.00962857
R77592 VSS.n3021 VSS.n3020 0.00962857
R77593 VSS.n3022 VSS.n3021 0.00962857
R77594 VSS.n3022 VSS.n3004 0.00962857
R77595 VSS.n3028 VSS.n3004 0.00962857
R77596 VSS.n3029 VSS.n3028 0.00962857
R77597 VSS.n3030 VSS.n3029 0.00962857
R77598 VSS.n3030 VSS.n3000 0.00962857
R77599 VSS.n3037 VSS.n3000 0.00962857
R77600 VSS.n3038 VSS.n3037 0.00962857
R77601 VSS.n3039 VSS.n3038 0.00962857
R77602 VSS.n3039 VSS.n2975 0.00962857
R77603 VSS.n6742 VSS.n6741 0.00962857
R77604 VSS.n6741 VSS.n6740 0.00962857
R77605 VSS.n6740 VSS.n3046 0.00962857
R77606 VSS.n6734 VSS.n3046 0.00962857
R77607 VSS.n6734 VSS.n6733 0.00962857
R77608 VSS.n6733 VSS.n6732 0.00962857
R77609 VSS.n6732 VSS.n3050 0.00962857
R77610 VSS.n6726 VSS.n3050 0.00962857
R77611 VSS.n6726 VSS.n6725 0.00962857
R77612 VSS.n6725 VSS.n6724 0.00962857
R77613 VSS.n6724 VSS.n3054 0.00962857
R77614 VSS.n6718 VSS.n3054 0.00962857
R77615 VSS.n6708 VSS.n3087 0.00962857
R77616 VSS.n6708 VSS.n6707 0.00962857
R77617 VSS.n6707 VSS.n6706 0.00962857
R77618 VSS.n6706 VSS.n3088 0.00962857
R77619 VSS.n6690 VSS.n6667 0.00962857
R77620 VSS.n6684 VSS.n6667 0.00962857
R77621 VSS.n6684 VSS.n6683 0.00962857
R77622 VSS.n3918 VSS.n3916 0.00962857
R77623 VSS.n3920 VSS.n3918 0.00962857
R77624 VSS.n3920 VSS.n3914 0.00962857
R77625 VSS.n3925 VSS.n3914 0.00962857
R77626 VSS.n3925 VSS.n3912 0.00962857
R77627 VSS.n3929 VSS.n3912 0.00962857
R77628 VSS.n3930 VSS.n3929 0.00962857
R77629 VSS.n3930 VSS.n3909 0.00962857
R77630 VSS.n6211 VSS.n3909 0.00962857
R77631 VSS.n6211 VSS.n3910 0.00962857
R77632 VSS.n6207 VSS.n3910 0.00962857
R77633 VSS.n6207 VSS.n3934 0.00962857
R77634 VSS.n6203 VSS.n3934 0.00962857
R77635 VSS.n6203 VSS.n3936 0.00962857
R77636 VSS.n6199 VSS.n3936 0.00962857
R77637 VSS.n6199 VSS.n3938 0.00962857
R77638 VSS.n3962 VSS.n3938 0.00962857
R77639 VSS.n3962 VSS.n3959 0.00962857
R77640 VSS.n6191 VSS.n3959 0.00962857
R77641 VSS.n6191 VSS.n3960 0.00962857
R77642 VSS.n6187 VSS.n3960 0.00962857
R77643 VSS.n6187 VSS.n3966 0.00962857
R77644 VSS.n6183 VSS.n3966 0.00962857
R77645 VSS.n6183 VSS.n3968 0.00962857
R77646 VSS.n6179 VSS.n3968 0.00962857
R77647 VSS.n6179 VSS.n3970 0.00962857
R77648 VSS.n6175 VSS.n3970 0.00962857
R77649 VSS.n6175 VSS.n3972 0.00962857
R77650 VSS.n6171 VSS.n3972 0.00962857
R77651 VSS.n6171 VSS.n3974 0.00962857
R77652 VSS.n6167 VSS.n3974 0.00962857
R77653 VSS.n6167 VSS.n3976 0.00962857
R77654 VSS.n6163 VSS.n3976 0.00962857
R77655 VSS.n6163 VSS.n3978 0.00962857
R77656 VSS.n6155 VSS.n3978 0.00962857
R77657 VSS.n6155 VSS.n3998 0.00962857
R77658 VSS.n6151 VSS.n3998 0.00962857
R77659 VSS.n6151 VSS.n4000 0.00962857
R77660 VSS.n6147 VSS.n4000 0.00962857
R77661 VSS.n6147 VSS.n4002 0.00962857
R77662 VSS.n6143 VSS.n4002 0.00962857
R77663 VSS.n6143 VSS.n4004 0.00962857
R77664 VSS.n6139 VSS.n4004 0.00962857
R77665 VSS.n6139 VSS.n4006 0.00962857
R77666 VSS.n6135 VSS.n4006 0.00962857
R77667 VSS.n6135 VSS.n4008 0.00962857
R77668 VSS.n6131 VSS.n4008 0.00962857
R77669 VSS.n6131 VSS.n4010 0.00962857
R77670 VSS.n6127 VSS.n4010 0.00962857
R77671 VSS.n6127 VSS.n4012 0.00962857
R77672 VSS.n4181 VSS.n4012 0.00962857
R77673 VSS.n4183 VSS.n4181 0.00962857
R77674 VSS.n4183 VSS.n4177 0.00962857
R77675 VSS.n4220 VSS.n4177 0.00962857
R77676 VSS.n4220 VSS.n4178 0.00962857
R77677 VSS.n4216 VSS.n4178 0.00962857
R77678 VSS.n4216 VSS.n4187 0.00962857
R77679 VSS.n4212 VSS.n4187 0.00962857
R77680 VSS.n4212 VSS.n4189 0.00962857
R77681 VSS.n4208 VSS.n4189 0.00962857
R77682 VSS.n4208 VSS.n4191 0.00962857
R77683 VSS.n4204 VSS.n4191 0.00962857
R77684 VSS.n4204 VSS.n4193 0.00962857
R77685 VSS.n4200 VSS.n4193 0.00962857
R77686 VSS.n4200 VSS.n4197 0.00962857
R77687 VSS.n4197 VSS.n4196 0.00962857
R77688 VSS.n4196 VSS.n328 0.00962857
R77689 VSS.n9676 VSS.n328 0.00962857
R77690 VSS.n9676 VSS.n330 0.00962857
R77691 VSS.n9672 VSS.n330 0.00962857
R77692 VSS.n9672 VSS.n333 0.00962857
R77693 VSS.n9668 VSS.n333 0.00962857
R77694 VSS.n9668 VSS.n335 0.00962857
R77695 VSS.n9664 VSS.n335 0.00962857
R77696 VSS.n9664 VSS.n337 0.00962857
R77697 VSS.n9660 VSS.n337 0.00962857
R77698 VSS.n9660 VSS.n339 0.00962857
R77699 VSS.n9656 VSS.n339 0.00962857
R77700 VSS.n9656 VSS.n341 0.00962857
R77701 VSS.n9652 VSS.n341 0.00962857
R77702 VSS.n9652 VSS.n343 0.00962857
R77703 VSS.n9648 VSS.n343 0.00962857
R77704 VSS.n9648 VSS.n345 0.00962857
R77705 VSS.n371 VSS.n345 0.00962857
R77706 VSS.n371 VSS.n368 0.00962857
R77707 VSS.n9642 VSS.n368 0.00962857
R77708 VSS.n9642 VSS.n369 0.00962857
R77709 VSS.n9638 VSS.n369 0.00962857
R77710 VSS.n9638 VSS.n375 0.00962857
R77711 VSS.n9634 VSS.n375 0.00962857
R77712 VSS.n9634 VSS.n377 0.00962857
R77713 VSS.n9630 VSS.n377 0.00962857
R77714 VSS.n9630 VSS.n379 0.00962857
R77715 VSS.n9622 VSS.n379 0.00962857
R77716 VSS.n9622 VSS.n399 0.00962857
R77717 VSS.n9618 VSS.n399 0.00962857
R77718 VSS.n9618 VSS.n401 0.00962857
R77719 VSS.n9614 VSS.n403 0.00962857
R77720 VSS.n9610 VSS.n403 0.00962857
R77721 VSS.n9610 VSS.n405 0.00962857
R77722 VSS.n3926 VSS.n3913 0.00962857
R77723 VSS.n3927 VSS.n3926 0.00962857
R77724 VSS.n3928 VSS.n3927 0.00962857
R77725 VSS.n3928 VSS.n3895 0.00962857
R77726 VSS.n6212 VSS.n3908 0.00962857
R77727 VSS.n6206 VSS.n3908 0.00962857
R77728 VSS.n6206 VSS.n6205 0.00962857
R77729 VSS.n6205 VSS.n6204 0.00962857
R77730 VSS.n6204 VSS.n3935 0.00962857
R77731 VSS.n6198 VSS.n3935 0.00962857
R77732 VSS.n6192 VSS.n3958 0.00962857
R77733 VSS.n6186 VSS.n3958 0.00962857
R77734 VSS.n6186 VSS.n6185 0.00962857
R77735 VSS.n6185 VSS.n6184 0.00962857
R77736 VSS.n6184 VSS.n3967 0.00962857
R77737 VSS.n6178 VSS.n3967 0.00962857
R77738 VSS.n6178 VSS.n6177 0.00962857
R77739 VSS.n6177 VSS.n6176 0.00962857
R77740 VSS.n6176 VSS.n3971 0.00962857
R77741 VSS.n6170 VSS.n3971 0.00962857
R77742 VSS.n6170 VSS.n6169 0.00962857
R77743 VSS.n6169 VSS.n6168 0.00962857
R77744 VSS.n6156 VSS.n3997 0.00962857
R77745 VSS.n6150 VSS.n3997 0.00962857
R77746 VSS.n6150 VSS.n6149 0.00962857
R77747 VSS.n6149 VSS.n6148 0.00962857
R77748 VSS.n6148 VSS.n4001 0.00962857
R77749 VSS.n6142 VSS.n4001 0.00962857
R77750 VSS.n6142 VSS.n6141 0.00962857
R77751 VSS.n6141 VSS.n6140 0.00962857
R77752 VSS.n6140 VSS.n4005 0.00962857
R77753 VSS.n6134 VSS.n4005 0.00962857
R77754 VSS.n6134 VSS.n6133 0.00962857
R77755 VSS.n6133 VSS.n6132 0.00962857
R77756 VSS.n4180 VSS.n4020 0.00962857
R77757 VSS.n4221 VSS.n4176 0.00962857
R77758 VSS.n4215 VSS.n4176 0.00962857
R77759 VSS.n4215 VSS.n4214 0.00962857
R77760 VSS.n4214 VSS.n4213 0.00962857
R77761 VSS.n4213 VSS.n4188 0.00962857
R77762 VSS.n4207 VSS.n4188 0.00962857
R77763 VSS.n4207 VSS.n4206 0.00962857
R77764 VSS.n4206 VSS.n4205 0.00962857
R77765 VSS.n4205 VSS.n4192 0.00962857
R77766 VSS.n4199 VSS.n4192 0.00962857
R77767 VSS.n4199 VSS.n4198 0.00962857
R77768 VSS.n4198 VSS.n311 0.00962857
R77769 VSS.n9671 VSS.n9670 0.00962857
R77770 VSS.n9670 VSS.n9669 0.00962857
R77771 VSS.n9669 VSS.n334 0.00962857
R77772 VSS.n9663 VSS.n334 0.00962857
R77773 VSS.n9663 VSS.n9662 0.00962857
R77774 VSS.n9662 VSS.n9661 0.00962857
R77775 VSS.n9661 VSS.n338 0.00962857
R77776 VSS.n9655 VSS.n338 0.00962857
R77777 VSS.n9655 VSS.n9654 0.00962857
R77778 VSS.n9654 VSS.n9653 0.00962857
R77779 VSS.n9653 VSS.n342 0.00962857
R77780 VSS.n9647 VSS.n342 0.00962857
R77781 VSS.n9643 VSS.n367 0.00962857
R77782 VSS.n9637 VSS.n367 0.00962857
R77783 VSS.n9637 VSS.n9636 0.00962857
R77784 VSS.n9636 VSS.n9635 0.00962857
R77785 VSS.n9623 VSS.n398 0.00962857
R77786 VSS.n9617 VSS.n398 0.00962857
R77787 VSS.n9617 VSS.n9616 0.00962857
R77788 VSS.n6237 VSS.n6236 0.00962857
R77789 VSS.n6236 VSS.n3875 0.00962857
R77790 VSS.n6231 VSS.n3875 0.00962857
R77791 VSS.n6231 VSS.n3877 0.00962857
R77792 VSS.n6227 VSS.n3877 0.00962857
R77793 VSS.n6227 VSS.n3879 0.00962857
R77794 VSS.n6223 VSS.n3879 0.00962857
R77795 VSS.n6223 VSS.n3881 0.00962857
R77796 VSS.n5278 VSS.n3881 0.00962857
R77797 VSS.n5280 VSS.n5278 0.00962857
R77798 VSS.n5280 VSS.n5276 0.00962857
R77799 VSS.n5284 VSS.n5276 0.00962857
R77800 VSS.n5284 VSS.n5274 0.00962857
R77801 VSS.n5288 VSS.n5274 0.00962857
R77802 VSS.n5288 VSS.n5272 0.00962857
R77803 VSS.n5292 VSS.n5272 0.00962857
R77804 VSS.n5292 VSS.n4312 0.00962857
R77805 VSS.n5305 VSS.n4312 0.00962857
R77806 VSS.n5305 VSS.n4310 0.00962857
R77807 VSS.n5309 VSS.n4310 0.00962857
R77808 VSS.n5309 VSS.n4308 0.00962857
R77809 VSS.n5313 VSS.n4308 0.00962857
R77810 VSS.n5313 VSS.n4306 0.00962857
R77811 VSS.n5317 VSS.n4306 0.00962857
R77812 VSS.n5317 VSS.n4304 0.00962857
R77813 VSS.n5321 VSS.n4304 0.00962857
R77814 VSS.n5321 VSS.n4302 0.00962857
R77815 VSS.n5325 VSS.n4302 0.00962857
R77816 VSS.n5325 VSS.n4300 0.00962857
R77817 VSS.n5329 VSS.n4300 0.00962857
R77818 VSS.n5329 VSS.n4296 0.00962857
R77819 VSS.n5629 VSS.n4296 0.00962857
R77820 VSS.n5629 VSS.n4298 0.00962857
R77821 VSS.n5625 VSS.n4298 0.00962857
R77822 VSS.n5625 VSS.n5623 0.00962857
R77823 VSS.n5623 VSS.n5333 0.00962857
R77824 VSS.n5619 VSS.n5333 0.00962857
R77825 VSS.n5619 VSS.n5335 0.00962857
R77826 VSS.n5615 VSS.n5335 0.00962857
R77827 VSS.n5615 VSS.n5338 0.00962857
R77828 VSS.n5611 VSS.n5338 0.00962857
R77829 VSS.n5611 VSS.n5340 0.00962857
R77830 VSS.n5607 VSS.n5340 0.00962857
R77831 VSS.n5607 VSS.n5342 0.00962857
R77832 VSS.n5603 VSS.n5342 0.00962857
R77833 VSS.n5603 VSS.n5344 0.00962857
R77834 VSS.n5599 VSS.n5344 0.00962857
R77835 VSS.n5599 VSS.n5598 0.00962857
R77836 VSS.n5598 VSS.n5597 0.00962857
R77837 VSS.n5597 VSS.n5347 0.00962857
R77838 VSS.n5592 VSS.n5347 0.00962857
R77839 VSS.n5592 VSS.n5591 0.00962857
R77840 VSS.n5591 VSS.n5590 0.00962857
R77841 VSS.n5590 VSS.n5349 0.00962857
R77842 VSS.n5585 VSS.n5349 0.00962857
R77843 VSS.n5585 VSS.n5351 0.00962857
R77844 VSS.n5581 VSS.n5351 0.00962857
R77845 VSS.n5581 VSS.n5354 0.00962857
R77846 VSS.n5577 VSS.n5354 0.00962857
R77847 VSS.n5577 VSS.n5356 0.00962857
R77848 VSS.n5573 VSS.n5356 0.00962857
R77849 VSS.n5573 VSS.n5358 0.00962857
R77850 VSS.n5569 VSS.n5358 0.00962857
R77851 VSS.n5569 VSS.n5360 0.00962857
R77852 VSS.n5565 VSS.n5360 0.00962857
R77853 VSS.n5565 VSS.n5361 0.00962857
R77854 VSS.n5561 VSS.n5361 0.00962857
R77855 VSS.n5561 VSS.n5560 0.00962857
R77856 VSS.n5560 VSS.n5558 0.00962857
R77857 VSS.n5558 VSS.n5363 0.00962857
R77858 VSS.n5553 VSS.n5363 0.00962857
R77859 VSS.n5553 VSS.n5365 0.00962857
R77860 VSS.n5549 VSS.n5365 0.00962857
R77861 VSS.n5549 VSS.n5368 0.00962857
R77862 VSS.n5545 VSS.n5368 0.00962857
R77863 VSS.n5545 VSS.n5370 0.00962857
R77864 VSS.n5541 VSS.n5370 0.00962857
R77865 VSS.n5541 VSS.n5372 0.00962857
R77866 VSS.n5537 VSS.n5372 0.00962857
R77867 VSS.n5537 VSS.n5374 0.00962857
R77868 VSS.n5533 VSS.n5374 0.00962857
R77869 VSS.n5533 VSS.n5376 0.00962857
R77870 VSS.n5529 VSS.n5376 0.00962857
R77871 VSS.n5529 VSS.n5378 0.00962857
R77872 VSS.n5397 VSS.n5378 0.00962857
R77873 VSS.n5520 VSS.n5397 0.00962857
R77874 VSS.n5520 VSS.n5398 0.00962857
R77875 VSS.n5516 VSS.n5398 0.00962857
R77876 VSS.n5516 VSS.n5401 0.00962857
R77877 VSS.n5512 VSS.n5401 0.00962857
R77878 VSS.n5512 VSS.n5403 0.00962857
R77879 VSS.n5508 VSS.n5403 0.00962857
R77880 VSS.n5508 VSS.n5405 0.00962857
R77881 VSS.n5499 VSS.n5405 0.00962857
R77882 VSS.n5499 VSS.n5423 0.00962857
R77883 VSS.n5495 VSS.n5423 0.00962857
R77884 VSS.n5495 VSS.n5425 0.00962857
R77885 VSS.n5491 VSS.n5427 0.00962857
R77886 VSS.n5487 VSS.n5427 0.00962857
R77887 VSS.n5487 VSS.n5429 0.00962857
R77888 VSS.n6230 VSS.n6229 0.00962857
R77889 VSS.n6229 VSS.n6228 0.00962857
R77890 VSS.n6228 VSS.n3878 0.00962857
R77891 VSS.n6222 VSS.n3878 0.00962857
R77892 VSS.n5279 VSS.n3893 0.00962857
R77893 VSS.n5279 VSS.n5275 0.00962857
R77894 VSS.n5285 VSS.n5275 0.00962857
R77895 VSS.n5286 VSS.n5285 0.00962857
R77896 VSS.n5287 VSS.n5286 0.00962857
R77897 VSS.n5287 VSS.n5269 0.00962857
R77898 VSS.n5310 VSS.n4309 0.00962857
R77899 VSS.n5311 VSS.n5310 0.00962857
R77900 VSS.n5312 VSS.n5311 0.00962857
R77901 VSS.n5312 VSS.n4305 0.00962857
R77902 VSS.n5318 VSS.n4305 0.00962857
R77903 VSS.n5319 VSS.n5318 0.00962857
R77904 VSS.n5320 VSS.n5319 0.00962857
R77905 VSS.n5320 VSS.n4301 0.00962857
R77906 VSS.n5326 VSS.n4301 0.00962857
R77907 VSS.n5327 VSS.n5326 0.00962857
R77908 VSS.n5328 VSS.n5327 0.00962857
R77909 VSS.n5328 VSS.n4292 0.00962857
R77910 VSS.n5622 VSS.n5621 0.00962857
R77911 VSS.n5621 VSS.n5620 0.00962857
R77912 VSS.n5620 VSS.n5334 0.00962857
R77913 VSS.n5614 VSS.n5334 0.00962857
R77914 VSS.n5614 VSS.n5613 0.00962857
R77915 VSS.n5613 VSS.n5612 0.00962857
R77916 VSS.n5612 VSS.n5339 0.00962857
R77917 VSS.n5606 VSS.n5339 0.00962857
R77918 VSS.n5606 VSS.n5605 0.00962857
R77919 VSS.n5605 VSS.n5604 0.00962857
R77920 VSS.n5604 VSS.n5343 0.00962857
R77921 VSS.n5343 VSS.n4265 0.00962857
R77922 VSS.n5346 VSS.n4247 0.00962857
R77923 VSS.n5584 VSS.n5352 0.00962857
R77924 VSS.n5584 VSS.n5583 0.00962857
R77925 VSS.n5583 VSS.n5582 0.00962857
R77926 VSS.n5582 VSS.n5353 0.00962857
R77927 VSS.n5576 VSS.n5353 0.00962857
R77928 VSS.n5576 VSS.n5575 0.00962857
R77929 VSS.n5575 VSS.n5574 0.00962857
R77930 VSS.n5574 VSS.n5357 0.00962857
R77931 VSS.n5568 VSS.n5357 0.00962857
R77932 VSS.n5568 VSS.n5567 0.00962857
R77933 VSS.n5567 VSS.n5566 0.00962857
R77934 VSS.n5566 VSS.n290 0.00962857
R77935 VSS.n5552 VSS.n5366 0.00962857
R77936 VSS.n5552 VSS.n5551 0.00962857
R77937 VSS.n5551 VSS.n5550 0.00962857
R77938 VSS.n5550 VSS.n5367 0.00962857
R77939 VSS.n5544 VSS.n5367 0.00962857
R77940 VSS.n5544 VSS.n5543 0.00962857
R77941 VSS.n5543 VSS.n5542 0.00962857
R77942 VSS.n5542 VSS.n5371 0.00962857
R77943 VSS.n5536 VSS.n5371 0.00962857
R77944 VSS.n5536 VSS.n5535 0.00962857
R77945 VSS.n5535 VSS.n5534 0.00962857
R77946 VSS.n5534 VSS.n5375 0.00962857
R77947 VSS.n5521 VSS.n5396 0.00962857
R77948 VSS.n5515 VSS.n5396 0.00962857
R77949 VSS.n5515 VSS.n5514 0.00962857
R77950 VSS.n5514 VSS.n5513 0.00962857
R77951 VSS.n5500 VSS.n5422 0.00962857
R77952 VSS.n5494 VSS.n5422 0.00962857
R77953 VSS.n5494 VSS.n5493 0.00962857
R77954 VSS.n4771 VSS.n4580 0.00962857
R77955 VSS.n4772 VSS.n4771 0.00962857
R77956 VSS.n4773 VSS.n4772 0.00962857
R77957 VSS.n4773 VSS.n4572 0.00962857
R77958 VSS.n4793 VSS.n4548 0.00962857
R77959 VSS.n4794 VSS.n4793 0.00962857
R77960 VSS.n4795 VSS.n4794 0.00962857
R77961 VSS.n4795 VSS.n4333 0.00962857
R77962 VSS.n4809 VSS.n4542 0.00962857
R77963 VSS.n4810 VSS.n4809 0.00962857
R77964 VSS.n4811 VSS.n4810 0.00962857
R77965 VSS.n4811 VSS.n4538 0.00962857
R77966 VSS.n4817 VSS.n4538 0.00962857
R77967 VSS.n4818 VSS.n4817 0.00962857
R77968 VSS.n4819 VSS.n4818 0.00962857
R77969 VSS.n4819 VSS.n4534 0.00962857
R77970 VSS.n4825 VSS.n4534 0.00962857
R77971 VSS.n4826 VSS.n4825 0.00962857
R77972 VSS.n4827 VSS.n4826 0.00962857
R77973 VSS.n4827 VSS.n4525 0.00962857
R77974 VSS.n5052 VSS.n5051 0.00962857
R77975 VSS.n5051 VSS.n5050 0.00962857
R77976 VSS.n5050 VSS.n4833 0.00962857
R77977 VSS.n5044 VSS.n4833 0.00962857
R77978 VSS.n5044 VSS.n5043 0.00962857
R77979 VSS.n5043 VSS.n5042 0.00962857
R77980 VSS.n5042 VSS.n4838 0.00962857
R77981 VSS.n5036 VSS.n4838 0.00962857
R77982 VSS.n5036 VSS.n5035 0.00962857
R77983 VSS.n5035 VSS.n5034 0.00962857
R77984 VSS.n5034 VSS.n4842 0.00962857
R77985 VSS.n4842 VSS.n4494 0.00962857
R77986 VSS.n5021 VSS.n4848 0.00962857
R77987 VSS.n5017 VSS.n4976 0.00962857
R77988 VSS.n5011 VSS.n4976 0.00962857
R77989 VSS.n5011 VSS.n5010 0.00962857
R77990 VSS.n5010 VSS.n5009 0.00962857
R77991 VSS.n5009 VSS.n4982 0.00962857
R77992 VSS.n5003 VSS.n4982 0.00962857
R77993 VSS.n5003 VSS.n5002 0.00962857
R77994 VSS.n5002 VSS.n5001 0.00962857
R77995 VSS.n5001 VSS.n4986 0.00962857
R77996 VSS.n4995 VSS.n4986 0.00962857
R77997 VSS.n4995 VSS.n4994 0.00962857
R77998 VSS.n4994 VSS.n259 0.00962857
R77999 VSS.n9703 VSS.n246 0.00962857
R78000 VSS.n9704 VSS.n9703 0.00962857
R78001 VSS.n9705 VSS.n9704 0.00962857
R78002 VSS.n9705 VSS.n242 0.00962857
R78003 VSS.n9711 VSS.n242 0.00962857
R78004 VSS.n9712 VSS.n9711 0.00962857
R78005 VSS.n9713 VSS.n9712 0.00962857
R78006 VSS.n9713 VSS.n238 0.00962857
R78007 VSS.n9719 VSS.n238 0.00962857
R78008 VSS.n9720 VSS.n9719 0.00962857
R78009 VSS.n9721 VSS.n9720 0.00962857
R78010 VSS.n9721 VSS.n229 0.00962857
R78011 VSS.n9739 VSS.n9738 0.00962857
R78012 VSS.n9738 VSS.n9737 0.00962857
R78013 VSS.n9737 VSS.n9727 0.00962857
R78014 VSS.n9727 VSS.n206 0.00962857
R78015 VSS.n9785 VSS.n190 0.00962857
R78016 VSS.n9786 VSS.n9785 0.00962857
R78017 VSS.n9787 VSS.n9786 0.00962857
R78018 VSS.n7876 VSS.n7875 0.00962857
R78019 VSS.n7875 VSS.n7274 0.00962857
R78020 VSS.n7871 VSS.n7274 0.00962857
R78021 VSS.n7871 VSS.n7276 0.00962857
R78022 VSS.n7867 VSS.n7276 0.00962857
R78023 VSS.n7867 VSS.n7279 0.00962857
R78024 VSS.n7863 VSS.n7279 0.00962857
R78025 VSS.n7863 VSS.n7281 0.00962857
R78026 VSS.n7859 VSS.n7281 0.00962857
R78027 VSS.n7859 VSS.n7283 0.00962857
R78028 VSS.n7855 VSS.n7283 0.00962857
R78029 VSS.n7855 VSS.n7285 0.00962857
R78030 VSS.n7851 VSS.n7285 0.00962857
R78031 VSS.n7851 VSS.n7600 0.00962857
R78032 VSS.n7847 VSS.n7600 0.00962857
R78033 VSS.n7847 VSS.n7602 0.00962857
R78034 VSS.n7843 VSS.n7602 0.00962857
R78035 VSS.n7843 VSS.n7604 0.00962857
R78036 VSS.n7839 VSS.n7604 0.00962857
R78037 VSS.n7839 VSS.n7606 0.00962857
R78038 VSS.n7835 VSS.n7606 0.00962857
R78039 VSS.n7835 VSS.n7608 0.00962857
R78040 VSS.n7831 VSS.n7608 0.00962857
R78041 VSS.n7831 VSS.n7610 0.00962857
R78042 VSS.n7827 VSS.n7610 0.00962857
R78043 VSS.n7827 VSS.n7612 0.00962857
R78044 VSS.n7823 VSS.n7612 0.00962857
R78045 VSS.n7823 VSS.n7614 0.00962857
R78046 VSS.n7819 VSS.n7614 0.00962857
R78047 VSS.n7819 VSS.n7616 0.00962857
R78048 VSS.n7815 VSS.n7616 0.00962857
R78049 VSS.n7815 VSS.n7618 0.00962857
R78050 VSS.n7811 VSS.n7618 0.00962857
R78051 VSS.n7811 VSS.n7620 0.00962857
R78052 VSS.n7807 VSS.n7620 0.00962857
R78053 VSS.n7807 VSS.n7622 0.00962857
R78054 VSS.n7803 VSS.n7622 0.00962857
R78055 VSS.n7803 VSS.n7624 0.00962857
R78056 VSS.n7799 VSS.n7624 0.00962857
R78057 VSS.n7799 VSS.n7626 0.00962857
R78058 VSS.n7795 VSS.n7626 0.00962857
R78059 VSS.n7795 VSS.n7628 0.00962857
R78060 VSS.n7791 VSS.n7628 0.00962857
R78061 VSS.n7791 VSS.n7630 0.00962857
R78062 VSS.n7787 VSS.n7630 0.00962857
R78063 VSS.n7787 VSS.n7632 0.00962857
R78064 VSS.n7783 VSS.n7632 0.00962857
R78065 VSS.n7783 VSS.n7634 0.00962857
R78066 VSS.n7779 VSS.n7634 0.00962857
R78067 VSS.n7779 VSS.n7636 0.00962857
R78068 VSS.n7775 VSS.n7636 0.00962857
R78069 VSS.n7775 VSS.n7638 0.00962857
R78070 VSS.n7771 VSS.n7638 0.00962857
R78071 VSS.n7771 VSS.n7640 0.00962857
R78072 VSS.n7767 VSS.n7640 0.00962857
R78073 VSS.n7767 VSS.n7642 0.00962857
R78074 VSS.n7763 VSS.n7642 0.00962857
R78075 VSS.n7763 VSS.n7644 0.00962857
R78076 VSS.n7759 VSS.n7644 0.00962857
R78077 VSS.n7759 VSS.n7646 0.00962857
R78078 VSS.n7755 VSS.n7646 0.00962857
R78079 VSS.n7755 VSS.n7648 0.00962857
R78080 VSS.n7751 VSS.n7648 0.00962857
R78081 VSS.n7751 VSS.n7650 0.00962857
R78082 VSS.n7747 VSS.n7650 0.00962857
R78083 VSS.n7747 VSS.n7652 0.00962857
R78084 VSS.n7743 VSS.n7652 0.00962857
R78085 VSS.n7743 VSS.n7654 0.00962857
R78086 VSS.n7739 VSS.n7654 0.00962857
R78087 VSS.n7739 VSS.n7656 0.00962857
R78088 VSS.n7735 VSS.n7656 0.00962857
R78089 VSS.n7735 VSS.n7658 0.00962857
R78090 VSS.n7731 VSS.n7658 0.00962857
R78091 VSS.n7731 VSS.n7660 0.00962857
R78092 VSS.n7727 VSS.n7660 0.00962857
R78093 VSS.n7727 VSS.n7662 0.00962857
R78094 VSS.n7723 VSS.n7662 0.00962857
R78095 VSS.n7723 VSS.n7664 0.00962857
R78096 VSS.n7719 VSS.n7664 0.00962857
R78097 VSS.n7719 VSS.n7666 0.00962857
R78098 VSS.n7715 VSS.n7666 0.00962857
R78099 VSS.n7715 VSS.n7668 0.00962857
R78100 VSS.n7711 VSS.n7668 0.00962857
R78101 VSS.n7711 VSS.n7670 0.00962857
R78102 VSS.n7707 VSS.n7670 0.00962857
R78103 VSS.n7707 VSS.n7672 0.00962857
R78104 VSS.n7703 VSS.n7672 0.00962857
R78105 VSS.n7703 VSS.n7674 0.00962857
R78106 VSS.n7699 VSS.n7674 0.00962857
R78107 VSS.n7699 VSS.n7676 0.00962857
R78108 VSS.n7695 VSS.n7676 0.00962857
R78109 VSS.n7695 VSS.n7678 0.00962857
R78110 VSS.n7691 VSS.n7678 0.00962857
R78111 VSS.n7691 VSS.n7680 0.00962857
R78112 VSS.n7687 VSS.n7680 0.00962857
R78113 VSS.n7687 VSS.n7684 0.00962857
R78114 VSS.n7684 VSS.n7683 0.00962857
R78115 VSS.n9914 VSS.n2 0.00962857
R78116 VSS.n9910 VSS.n2 0.00962857
R78117 VSS.n9910 VSS.n4 0.00962857
R78118 VSS.n7878 VSS.n7877 0.00962857
R78119 VSS.n7877 VSS.n7273 0.00962857
R78120 VSS.n7277 VSS.n7273 0.00962857
R78121 VSS.n7870 VSS.n7277 0.00962857
R78122 VSS.n7870 VSS.n7869 0.00962857
R78123 VSS.n7869 VSS.n7868 0.00962857
R78124 VSS.n7868 VSS.n7278 0.00962857
R78125 VSS.n7862 VSS.n7278 0.00962857
R78126 VSS.n7862 VSS.n7861 0.00962857
R78127 VSS.n7861 VSS.n7860 0.00962857
R78128 VSS.n7854 VSS.n7853 0.00962857
R78129 VSS.n7853 VSS.n7852 0.00962857
R78130 VSS.n7852 VSS.n7599 0.00962857
R78131 VSS.n7846 VSS.n7599 0.00962857
R78132 VSS.n7846 VSS.n7845 0.00962857
R78133 VSS.n7845 VSS.n7844 0.00962857
R78134 VSS.n7844 VSS.n7603 0.00962857
R78135 VSS.n7838 VSS.n7603 0.00962857
R78136 VSS.n7838 VSS.n7837 0.00962857
R78137 VSS.n7837 VSS.n7836 0.00962857
R78138 VSS.n7836 VSS.n7607 0.00962857
R78139 VSS.n7830 VSS.n7607 0.00962857
R78140 VSS.n7830 VSS.n7829 0.00962857
R78141 VSS.n7829 VSS.n7828 0.00962857
R78142 VSS.n7828 VSS.n7611 0.00962857
R78143 VSS.n7822 VSS.n7611 0.00962857
R78144 VSS.n7822 VSS.n7821 0.00962857
R78145 VSS.n7821 VSS.n7820 0.00962857
R78146 VSS.n7820 VSS.n7615 0.00962857
R78147 VSS.n7814 VSS.n7615 0.00962857
R78148 VSS.n7814 VSS.n7813 0.00962857
R78149 VSS.n7813 VSS.n7812 0.00962857
R78150 VSS.n7812 VSS.n7619 0.00962857
R78151 VSS.n7806 VSS.n7619 0.00962857
R78152 VSS.n7806 VSS.n7805 0.00962857
R78153 VSS.n7805 VSS.n7804 0.00962857
R78154 VSS.n7804 VSS.n7623 0.00962857
R78155 VSS.n7798 VSS.n7623 0.00962857
R78156 VSS.n7798 VSS.n7797 0.00962857
R78157 VSS.n7797 VSS.n7796 0.00962857
R78158 VSS.n7796 VSS.n7627 0.00962857
R78159 VSS.n7790 VSS.n7627 0.00962857
R78160 VSS.n7790 VSS.n7789 0.00962857
R78161 VSS.n7789 VSS.n7788 0.00962857
R78162 VSS.n7788 VSS.n7631 0.00962857
R78163 VSS.n7782 VSS.n7631 0.00962857
R78164 VSS.n7782 VSS.n7781 0.00962857
R78165 VSS.n7781 VSS.n7780 0.00962857
R78166 VSS.n7780 VSS.n7635 0.00962857
R78167 VSS.n7774 VSS.n7635 0.00962857
R78168 VSS.n7774 VSS.n7773 0.00962857
R78169 VSS.n7773 VSS.n7772 0.00962857
R78170 VSS.n7772 VSS.n7639 0.00962857
R78171 VSS.n7766 VSS.n7639 0.00962857
R78172 VSS.n7766 VSS.n7765 0.00962857
R78173 VSS.n7765 VSS.n7764 0.00962857
R78174 VSS.n7764 VSS.n7643 0.00962857
R78175 VSS.n7758 VSS.n7643 0.00962857
R78176 VSS.n7758 VSS.n7757 0.00962857
R78177 VSS.n7757 VSS.n7756 0.00962857
R78178 VSS.n7756 VSS.n7647 0.00962857
R78179 VSS.n7750 VSS.n7647 0.00962857
R78180 VSS.n7750 VSS.n7749 0.00962857
R78181 VSS.n7749 VSS.n7748 0.00962857
R78182 VSS.n7748 VSS.n7651 0.00962857
R78183 VSS.n7742 VSS.n7651 0.00962857
R78184 VSS.n7742 VSS.n7741 0.00962857
R78185 VSS.n7741 VSS.n7740 0.00962857
R78186 VSS.n7740 VSS.n7655 0.00962857
R78187 VSS.n7734 VSS.n7655 0.00962857
R78188 VSS.n7734 VSS.n7733 0.00962857
R78189 VSS.n7733 VSS.n7732 0.00962857
R78190 VSS.n7732 VSS.n7659 0.00962857
R78191 VSS.n7726 VSS.n7659 0.00962857
R78192 VSS.n7726 VSS.n7725 0.00962857
R78193 VSS.n7725 VSS.n7724 0.00962857
R78194 VSS.n7724 VSS.n7663 0.00962857
R78195 VSS.n7718 VSS.n7663 0.00962857
R78196 VSS.n7718 VSS.n7717 0.00962857
R78197 VSS.n7717 VSS.n7716 0.00962857
R78198 VSS.n7716 VSS.n7667 0.00962857
R78199 VSS.n7710 VSS.n7667 0.00962857
R78200 VSS.n7710 VSS.n7709 0.00962857
R78201 VSS.n7709 VSS.n7708 0.00962857
R78202 VSS.n7708 VSS.n7671 0.00962857
R78203 VSS.n7702 VSS.n7671 0.00962857
R78204 VSS.n7702 VSS.n7701 0.00962857
R78205 VSS.n7701 VSS.n7700 0.00962857
R78206 VSS.n7700 VSS.n7675 0.00962857
R78207 VSS.n7694 VSS.n7675 0.00962857
R78208 VSS.n7694 VSS.n7693 0.00962857
R78209 VSS.n7693 VSS.n7692 0.00962857
R78210 VSS.n7692 VSS.n7679 0.00962857
R78211 VSS.n7686 VSS.n7679 0.00962857
R78212 VSS.n7686 VSS.n7685 0.00962857
R78213 VSS.n7685 VSS.n0 0.00962857
R78214 VSS.n9915 VSS.n1 0.00962857
R78215 VSS.n9909 VSS.n1 0.00962857
R78216 VSS.n9909 VSS.n9908 0.00962857
R78217 VSS.n9908 VSS.n9907 0.00962857
R78218 VSS.n7303 VSS.n7302 0.00962857
R78219 VSS.n7304 VSS.n7303 0.00962857
R78220 VSS.n7304 VSS.n7298 0.00962857
R78221 VSS.n7310 VSS.n7298 0.00962857
R78222 VSS.n7311 VSS.n7310 0.00962857
R78223 VSS.n7312 VSS.n7311 0.00962857
R78224 VSS.n7312 VSS.n7294 0.00962857
R78225 VSS.n7318 VSS.n7294 0.00962857
R78226 VSS.n7319 VSS.n7318 0.00962857
R78227 VSS.n7320 VSS.n7319 0.00962857
R78228 VSS.n7594 VSS.n7289 0.00962857
R78229 VSS.n7588 VSS.n7289 0.00962857
R78230 VSS.n7588 VSS.n7587 0.00962857
R78231 VSS.n7587 VSS.n7586 0.00962857
R78232 VSS.n7586 VSS.n7326 0.00962857
R78233 VSS.n7580 VSS.n7326 0.00962857
R78234 VSS.n7580 VSS.n7579 0.00962857
R78235 VSS.n7579 VSS.n7578 0.00962857
R78236 VSS.n7578 VSS.n7330 0.00962857
R78237 VSS.n7572 VSS.n7330 0.00962857
R78238 VSS.n7572 VSS.n7571 0.00962857
R78239 VSS.n7571 VSS.n7570 0.00962857
R78240 VSS.n7570 VSS.n7334 0.00962857
R78241 VSS.n7564 VSS.n7334 0.00962857
R78242 VSS.n7564 VSS.n7563 0.00962857
R78243 VSS.n7563 VSS.n7562 0.00962857
R78244 VSS.n7562 VSS.n7338 0.00962857
R78245 VSS.n7556 VSS.n7338 0.00962857
R78246 VSS.n7556 VSS.n7555 0.00962857
R78247 VSS.n7555 VSS.n7554 0.00962857
R78248 VSS.n7554 VSS.n7342 0.00962857
R78249 VSS.n7548 VSS.n7342 0.00962857
R78250 VSS.n7548 VSS.n7547 0.00962857
R78251 VSS.n7547 VSS.n7546 0.00962857
R78252 VSS.n7546 VSS.n7346 0.00962857
R78253 VSS.n7540 VSS.n7346 0.00962857
R78254 VSS.n7540 VSS.n7539 0.00962857
R78255 VSS.n7539 VSS.n7538 0.00962857
R78256 VSS.n7538 VSS.n7350 0.00962857
R78257 VSS.n7532 VSS.n7350 0.00962857
R78258 VSS.n7532 VSS.n7531 0.00962857
R78259 VSS.n7531 VSS.n7530 0.00962857
R78260 VSS.n7530 VSS.n7354 0.00962857
R78261 VSS.n7524 VSS.n7354 0.00962857
R78262 VSS.n7524 VSS.n7523 0.00962857
R78263 VSS.n7523 VSS.n7522 0.00962857
R78264 VSS.n7522 VSS.n7358 0.00962857
R78265 VSS.n7516 VSS.n7358 0.00962857
R78266 VSS.n7516 VSS.n7515 0.00962857
R78267 VSS.n7515 VSS.n7514 0.00962857
R78268 VSS.n7514 VSS.n7362 0.00962857
R78269 VSS.n7508 VSS.n7362 0.00962857
R78270 VSS.n7508 VSS.n7507 0.00962857
R78271 VSS.n7507 VSS.n7506 0.00962857
R78272 VSS.n7506 VSS.n7366 0.00962857
R78273 VSS.n7500 VSS.n7366 0.00962857
R78274 VSS.n7500 VSS.n7499 0.00962857
R78275 VSS.n7499 VSS.n7498 0.00962857
R78276 VSS.n7498 VSS.n7370 0.00962857
R78277 VSS.n7492 VSS.n7370 0.00962857
R78278 VSS.n7492 VSS.n7491 0.00962857
R78279 VSS.n7491 VSS.n7490 0.00962857
R78280 VSS.n7490 VSS.n7374 0.00962857
R78281 VSS.n7484 VSS.n7374 0.00962857
R78282 VSS.n7484 VSS.n7483 0.00962857
R78283 VSS.n7483 VSS.n7482 0.00962857
R78284 VSS.n7482 VSS.n7378 0.00962857
R78285 VSS.n7476 VSS.n7378 0.00962857
R78286 VSS.n7476 VSS.n7475 0.00962857
R78287 VSS.n7475 VSS.n7474 0.00962857
R78288 VSS.n7474 VSS.n7382 0.00962857
R78289 VSS.n7468 VSS.n7382 0.00962857
R78290 VSS.n7468 VSS.n7467 0.00962857
R78291 VSS.n7467 VSS.n7466 0.00962857
R78292 VSS.n7466 VSS.n7386 0.00962857
R78293 VSS.n7460 VSS.n7386 0.00962857
R78294 VSS.n7460 VSS.n7459 0.00962857
R78295 VSS.n7459 VSS.n7458 0.00962857
R78296 VSS.n7458 VSS.n7390 0.00962857
R78297 VSS.n7452 VSS.n7390 0.00962857
R78298 VSS.n7452 VSS.n7451 0.00962857
R78299 VSS.n7451 VSS.n7450 0.00962857
R78300 VSS.n7450 VSS.n7394 0.00962857
R78301 VSS.n7444 VSS.n7394 0.00962857
R78302 VSS.n7444 VSS.n7443 0.00962857
R78303 VSS.n7443 VSS.n7442 0.00962857
R78304 VSS.n7442 VSS.n7398 0.00962857
R78305 VSS.n7436 VSS.n7398 0.00962857
R78306 VSS.n7436 VSS.n7435 0.00962857
R78307 VSS.n7435 VSS.n7434 0.00962857
R78308 VSS.n7434 VSS.n7402 0.00962857
R78309 VSS.n7428 VSS.n7402 0.00962857
R78310 VSS.n7428 VSS.n7427 0.00962857
R78311 VSS.n7427 VSS.n7426 0.00962857
R78312 VSS.n7426 VSS.n7406 0.00962857
R78313 VSS.n7420 VSS.n7406 0.00962857
R78314 VSS.n7419 VSS.n7409 0.00962857
R78315 VSS.n7411 VSS.n7409 0.00962857
R78316 VSS.n7412 VSS.n7411 0.00962857
R78317 VSS.n7412 VSS.n6 0.00962857
R78318 VSS.n4755 VSS.n4747 0.00959466
R78319 VSS.n4750 VSS.n4749 0.00959466
R78320 VSS.n4752 VSS.n4749 0.00959466
R78321 VSS.n5248 VSS.n4322 0.00959466
R78322 VSS.n4328 VSS.n4321 0.00959466
R78323 VSS.n4328 VSS.n4324 0.00959466
R78324 VSS.n5074 VSS.n4519 0.00959466
R78325 VSS.n5075 VSS.n4518 0.00959466
R78326 VSS.n4518 VSS.n4514 0.00959466
R78327 VSS.n4512 VSS.n4506 0.00959466
R78328 VSS.n4512 VSS.n4509 0.00959466
R78329 VSS.n4970 VSS.n4873 0.00959466
R78330 VSS.n4970 VSS.n4968 0.00959466
R78331 VSS.n273 VSS.n271 0.00959466
R78332 VSS.n277 VSS.n270 0.00959466
R78333 VSS.n275 VSS.n270 0.00959466
R78334 VSS.n9761 VSS.n223 0.00959466
R78335 VSS.n9762 VSS.n222 0.00959466
R78336 VSS.n222 VSS.n218 0.00959466
R78337 VSS.n9767 VSS.n9766 0.00959466
R78338 VSS.n9768 VSS.n216 0.00959466
R78339 VSS.n9770 VSS.n216 0.00959466
R78340 VSS.n4751 VSS.n4750 0.00959466
R78341 VSS.n5249 VSS.n4321 0.00959466
R78342 VSS.n5076 VSS.n5075 0.00959466
R78343 VSS.n5079 VSS.n4506 0.00959466
R78344 VSS.n4971 VSS.n4873 0.00959466
R78345 VSS.n277 VSS.n272 0.00959466
R78346 VSS.n9763 VSS.n9762 0.00959466
R78347 VSS.n4751 VSS.n4747 0.00959466
R78348 VSS.n4753 VSS.n4752 0.00959466
R78349 VSS.n5249 VSS.n5248 0.00959466
R78350 VSS.n5251 VSS.n4324 0.00959466
R78351 VSS.n5076 VSS.n5074 0.00959466
R78352 VSS.n5078 VSS.n4514 0.00959466
R78353 VSS.n5081 VSS.n4509 0.00959466
R78354 VSS.n4973 VSS.n4968 0.00959466
R78355 VSS.n273 VSS.n272 0.00959466
R78356 VSS.n9691 VSS.n275 0.00959466
R78357 VSS.n9763 VSS.n9761 0.00959466
R78358 VSS.n9765 VSS.n218 0.00959466
R78359 VSS.n4566 VSS.n4564 0.00959466
R78360 VSS.n5259 VSS.n4319 0.00959466
R78361 VSS.n5257 VSS.n4318 0.00959466
R78362 VSS.n5257 VSS.n5254 0.00959466
R78363 VSS.n5644 VSS.n4286 0.00959466
R78364 VSS.n5645 VSS.n4285 0.00959466
R78365 VSS.n4285 VSS.n4281 0.00959466
R78366 VSS.n4279 VSS.n4274 0.00959466
R78367 VSS.n4279 VSS.n4276 0.00959466
R78368 VSS.n4917 VSS.n4913 0.00959466
R78369 VSS.n4916 VSS.n4913 0.00959466
R78370 VSS.n296 VSS.n279 0.00959466
R78371 VSS.n284 VSS.n278 0.00959466
R78372 VSS.n282 VSS.n278 0.00959466
R78373 VSS.n5453 VSS.n5451 0.00959466
R78374 VSS.n5454 VSS.n5450 0.00959466
R78375 VSS.n5450 VSS.n5447 0.00959466
R78376 VSS.n5460 VSS.n5458 0.00959466
R78377 VSS.n5461 VSS.n5445 0.00959466
R78378 VSS.n5445 VSS.n5442 0.00959466
R78379 VSS.n4569 VSS.n4566 0.00959466
R78380 VSS.n5260 VSS.n4318 0.00959466
R78381 VSS.n5646 VSS.n5645 0.00959466
R78382 VSS.n5650 VSS.n4274 0.00959466
R78383 VSS.n4917 VSS.n4914 0.00959466
R78384 VSS.n284 VSS.n281 0.00959466
R78385 VSS.n5455 VSS.n5454 0.00959466
R78386 VSS.n5260 VSS.n5259 0.00959466
R78387 VSS.n5262 VSS.n5254 0.00959466
R78388 VSS.n5646 VSS.n5644 0.00959466
R78389 VSS.n5648 VSS.n4281 0.00959466
R78390 VSS.n5652 VSS.n4276 0.00959466
R78391 VSS.n4921 VSS.n4916 0.00959466
R78392 VSS.n296 VSS.n281 0.00959466
R78393 VSS.n9686 VSS.n282 0.00959466
R78394 VSS.n5455 VSS.n5453 0.00959466
R78395 VSS.n5457 VSS.n5447 0.00959466
R78396 VSS.n4093 VSS.n4090 0.00959466
R78397 VSS.n4098 VSS.n4096 0.00959466
R78398 VSS.n4099 VSS.n4087 0.00959466
R78399 VSS.n4087 VSS.n4085 0.00959466
R78400 VSS.n4106 VSS.n4104 0.00959466
R78401 VSS.n4107 VSS.n4083 0.00959466
R78402 VSS.n4083 VSS.n4081 0.00959466
R78403 VSS.n4112 VSS.n4079 0.00959466
R78404 VSS.n4079 VSS.n4077 0.00959466
R78405 VSS.n4121 VSS.n4118 0.00959466
R78406 VSS.n4123 VSS.n4121 0.00959466
R78407 VSS.n4168 VSS.n4125 0.00959466
R78408 VSS.n4128 VSS.n4127 0.00959466
R78409 VSS.n4131 VSS.n4127 0.00959466
R78410 VSS.n4164 VSS.n4133 0.00959466
R78411 VSS.n4136 VSS.n4135 0.00959466
R78412 VSS.n4139 VSS.n4135 0.00959466
R78413 VSS.n4161 VSS.n4141 0.00959466
R78414 VSS.n4144 VSS.n4143 0.00959466
R78415 VSS.n4147 VSS.n4143 0.00959466
R78416 VSS.n4095 VSS.n4090 0.00959466
R78417 VSS.n4100 VSS.n4099 0.00959466
R78418 VSS.n4108 VSS.n4107 0.00959466
R78419 VSS.n4113 VSS.n4112 0.00959466
R78420 VSS.n5728 VSS.n4118 0.00959466
R78421 VSS.n4129 VSS.n4128 0.00959466
R78422 VSS.n4137 VSS.n4136 0.00959466
R78423 VSS.n4100 VSS.n4098 0.00959466
R78424 VSS.n4102 VSS.n4085 0.00959466
R78425 VSS.n4108 VSS.n4106 0.00959466
R78426 VSS.n4110 VSS.n4081 0.00959466
R78427 VSS.n4115 VSS.n4077 0.00959466
R78428 VSS.n5726 VSS.n4123 0.00959466
R78429 VSS.n4129 VSS.n4125 0.00959466
R78430 VSS.n4166 VSS.n4131 0.00959466
R78431 VSS.n4137 VSS.n4133 0.00959466
R78432 VSS.n4162 VSS.n4139 0.00959466
R78433 VSS.n6059 VSS.n6054 0.00959466
R78434 VSS.n6065 VSS.n6064 0.00959466
R78435 VSS.n6053 VSS.n6046 0.00959466
R78436 VSS.n6072 VSS.n6071 0.00959466
R78437 VSS.n6045 VSS.n6038 0.00959466
R78438 VSS.n4071 VSS.n4069 0.00959466
R78439 VSS.n5906 VSS.n5904 0.00959466
R78440 VSS.n5952 VSS.n5911 0.00959466
R78441 VSS.n5915 VSS.n5914 0.00959466
R78442 VSS.n5944 VSS.n5918 0.00959466
R78443 VSS.n5922 VSS.n5921 0.00959466
R78444 VSS.n5937 VSS.n5925 0.00959466
R78445 VSS.n5929 VSS.n5928 0.00959466
R78446 VSS.n6066 VSS.n6065 0.00959466
R78447 VSS.n6073 VSS.n6072 0.00959466
R78448 VSS.n5913 VSS.n5911 0.00959466
R78449 VSS.n5920 VSS.n5918 0.00959466
R78450 VSS.n6062 VSS.n6054 0.00959466
R78451 VSS.n6066 VSS.n6053 0.00959466
R78452 VSS.n6073 VSS.n6045 0.00959466
R78453 VSS.n6076 VSS.n4069 0.00959466
R78454 VSS.n5906 VSS.n5903 0.00959466
R78455 VSS.n5914 VSS.n5913 0.00959466
R78456 VSS.n5921 VSS.n5920 0.00959466
R78457 VSS.n6285 VSS.n3818 0.00959466
R78458 VSS.n6291 VSS.n6290 0.00959466
R78459 VSS.n3817 VSS.n3809 0.00959466
R78460 VSS.n6298 VSS.n6297 0.00959466
R78461 VSS.n3808 VSS.n3800 0.00959466
R78462 VSS.n3717 VSS.n3715 0.00959466
R78463 VSS.n6312 VSS.n3705 0.00959466
R78464 VSS.n6320 VSS.n6319 0.00959466
R78465 VSS.n3704 VSS.n3696 0.00959466
R78466 VSS.n6327 VSS.n6326 0.00959466
R78467 VSS.n3695 VSS.n3687 0.00959466
R78468 VSS.n6332 VSS.n3682 0.00959466
R78469 VSS.n6335 VSS.n3683 0.00959466
R78470 VSS.n6292 VSS.n6291 0.00959466
R78471 VSS.n6299 VSS.n6298 0.00959466
R78472 VSS.n6321 VSS.n6320 0.00959466
R78473 VSS.n6328 VSS.n6327 0.00959466
R78474 VSS.n6288 VSS.n3818 0.00959466
R78475 VSS.n6292 VSS.n3817 0.00959466
R78476 VSS.n6299 VSS.n3808 0.00959466
R78477 VSS.n6302 VSS.n3715 0.00959466
R78478 VSS.n6314 VSS.n6312 0.00959466
R78479 VSS.n6321 VSS.n3704 0.00959466
R78480 VSS.n6328 VSS.n3695 0.00959466
R78481 VSS.n6585 VSS.n6584 0.00959466
R78482 VSS.n3223 VSS.n3215 0.00959466
R78483 VSS.n6591 VSS.n6590 0.00959466
R78484 VSS.n3214 VSS.n3206 0.00959466
R78485 VSS.n6598 VSS.n6597 0.00959466
R78486 VSS.n3205 VSS.n3197 0.00959466
R78487 VSS.n3192 VSS.n3190 0.00959466
R78488 VSS.n6618 VSS.n3127 0.00959466
R78489 VSS.n6626 VSS.n6625 0.00959466
R78490 VSS.n3126 VSS.n3119 0.00959466
R78491 VSS.n6632 VSS.n3114 0.00959466
R78492 VSS.n6635 VSS.n3115 0.00959466
R78493 VSS.n3664 VSS.n3663 0.00959466
R78494 VSS.n3656 VSS.n3654 0.00959466
R78495 VSS.n6586 VSS.n6585 0.00959466
R78496 VSS.n6592 VSS.n6591 0.00959466
R78497 VSS.n6599 VSS.n6598 0.00959466
R78498 VSS.n6627 VSS.n6626 0.00959466
R78499 VSS.n6636 VSS.n3114 0.00959466
R78500 VSS.n6586 VSS.n3223 0.00959466
R78501 VSS.n6592 VSS.n3214 0.00959466
R78502 VSS.n6599 VSS.n3205 0.00959466
R78503 VSS.n6602 VSS.n3190 0.00959466
R78504 VSS.n6620 VSS.n6618 0.00959466
R78505 VSS.n6627 VSS.n3126 0.00959466
R78506 VSS.n6636 VSS.n6635 0.00959466
R78507 VSS.n5783 VSS.n5782 0.00959466
R78508 VSS.n5766 VSS.n5758 0.00959466
R78509 VSS.n5789 VSS.n5788 0.00959466
R78510 VSS.n5757 VSS.n5749 0.00959466
R78511 VSS.n5796 VSS.n5795 0.00959466
R78512 VSS.n5748 VSS.n5740 0.00959466
R78513 VSS.n5886 VSS.n5734 0.00959466
R78514 VSS.n5878 VSS.n2960 0.00959466
R78515 VSS.n6760 VSS.n2964 0.00959466
R78516 VSS.n2968 VSS.n2967 0.00959466
R78517 VSS.n6650 VSS.n6649 0.00959466
R78518 VSS.n6647 VSS.n3112 0.00959466
R78519 VSS.n6655 VSS.n3107 0.00959466
R78520 VSS.n6658 VSS.n3108 0.00959466
R78521 VSS.n5784 VSS.n5783 0.00959466
R78522 VSS.n5790 VSS.n5789 0.00959466
R78523 VSS.n5797 VSS.n5796 0.00959466
R78524 VSS.n6755 VSS.n2964 0.00959466
R78525 VSS.n6651 VSS.n6650 0.00959466
R78526 VSS.n5784 VSS.n5766 0.00959466
R78527 VSS.n5790 VSS.n5757 0.00959466
R78528 VSS.n5797 VSS.n5748 0.00959466
R78529 VSS.n5888 VSS.n5886 0.00959466
R78530 VSS.n5878 VSS.n2959 0.00959466
R78531 VSS.n6755 VSS.n2967 0.00959466
R78532 VSS.n6651 VSS.n6647 0.00959466
R78533 VSS.n6977 VSS.n6976 0.00959466
R78534 VSS.n2767 VSS.n2759 0.00959466
R78535 VSS.n6983 VSS.n6982 0.00959466
R78536 VSS.n2758 VSS.n2750 0.00959466
R78537 VSS.n6990 VSS.n6989 0.00959466
R78538 VSS.n2749 VSS.n2741 0.00959466
R78539 VSS.n2655 VSS.n2653 0.00959466
R78540 VSS.n7004 VSS.n2643 0.00959466
R78541 VSS.n7012 VSS.n7011 0.00959466
R78542 VSS.n2642 VSS.n2634 0.00959466
R78543 VSS.n7019 VSS.n7018 0.00959466
R78544 VSS.n2633 VSS.n2625 0.00959466
R78545 VSS.n7024 VSS.n2620 0.00959466
R78546 VSS.n7027 VSS.n2621 0.00959466
R78547 VSS.n6978 VSS.n6977 0.00959466
R78548 VSS.n6984 VSS.n6983 0.00959466
R78549 VSS.n6991 VSS.n6990 0.00959466
R78550 VSS.n7013 VSS.n7012 0.00959466
R78551 VSS.n7020 VSS.n7019 0.00959466
R78552 VSS.n6978 VSS.n2767 0.00959466
R78553 VSS.n6984 VSS.n2758 0.00959466
R78554 VSS.n6991 VSS.n2749 0.00959466
R78555 VSS.n6994 VSS.n2653 0.00959466
R78556 VSS.n7006 VSS.n7004 0.00959466
R78557 VSS.n7013 VSS.n2642 0.00959466
R78558 VSS.n7020 VSS.n2633 0.00959466
R78559 VSS.n7028 VSS.n2620 0.00959466
R78560 VSS.n6659 VSS.n3107 0.00959466
R78561 VSS.n3665 VSS.n3664 0.00959466
R78562 VSS.n6336 VSS.n3682 0.00959466
R78563 VSS.n5927 VSS.n5925 0.00959466
R78564 VSS.n4145 VSS.n4144 0.00959466
R78565 VSS.n4145 VSS.n4141 0.00959466
R78566 VSS.n4159 VSS.n4147 0.00959466
R78567 VSS.n5462 VSS.n5461 0.00959466
R78568 VSS.n5462 VSS.n5460 0.00959466
R78569 VSS.n5464 VSS.n5442 0.00959466
R78570 VSS.n9769 VSS.n9768 0.00959466
R78571 VSS.n9769 VSS.n9767 0.00959466
R78572 VSS.n9773 VSS.n9770 0.00959466
R78573 VSS.n5928 VSS.n5927 0.00959466
R78574 VSS.n6336 VSS.n6335 0.00959466
R78575 VSS.n3665 VSS.n3654 0.00959466
R78576 VSS.n6659 VSS.n6658 0.00959466
R78577 VSS.n7028 VSS.n7027 0.00959466
R78578 VSS.n3724 VSS.n3150 0.00958451
R78579 VSS.n2943 VSS.n2939 0.00958451
R78580 VSS.n3791 VSS.n3180 0.00958451
R78581 VSS.n2936 VSS.n2925 0.00958451
R78582 VSS.n9757 VSS.n217 0.00953543
R78583 VSS.n9764 VSS.n221 0.00953543
R78584 VSS.n224 VSS.n220 0.00953543
R78585 VSS.n9760 VSS.n225 0.00953543
R78586 VSS.n9759 VSS.n219 0.00953543
R78587 VSS.n9440 VSS.n9368 0.00953543
R78588 VSS.n2325 VSS.n2165 0.00953543
R78589 VSS.n2401 VSS.n1845 0.00953543
R78590 VSS.n4746 VSS.n4559 0.00953543
R78591 VSS.n4754 VSS.n4554 0.00953543
R78592 VSS.n4748 VSS.n4560 0.00953543
R78593 VSS.n4561 VSS.n4553 0.00953543
R78594 VSS.n4785 VSS.n4571 0.00953543
R78595 VSS.n9693 VSS.n9692 0.00953543
R78596 VSS.n9690 VSS.n254 0.00953543
R78597 VSS.n9689 VSS.n253 0.00953543
R78598 VSS.n274 VSS.n252 0.00953543
R78599 VSS.n9688 VSS.n251 0.00953543
R78600 VSS.n9445 VSS.n771 0.00953543
R78601 VSS.n5070 VSS.n4513 0.00953543
R78602 VSS.n5077 VSS.n4517 0.00953543
R78603 VSS.n4520 VSS.n4516 0.00953543
R78604 VSS.n5073 VSS.n4521 0.00953543
R78605 VSS.n5072 VSS.n4515 0.00953543
R78606 VSS.n2360 VSS.n1966 0.00953543
R78607 VSS.n5244 VSS.n4323 0.00953543
R78608 VSS.n5250 VSS.n4327 0.00953543
R78609 VSS.n4329 VSS.n4326 0.00953543
R78610 VSS.n5247 VSS.n5246 0.00953543
R78611 VSS.n5252 VSS.n4320 0.00953543
R78612 VSS.n2365 VSS.n1897 0.00953543
R78613 VSS.n4758 VSS.n4726 0.00953543
R78614 VSS.n6249 VSS.n3856 0.00953543
R78615 VSS.n9808 VSS.n171 0.00953543
R78616 VSS.n5467 VSS.n5439 0.00953543
R78617 VSS.n9775 VSS.n9774 0.00953543
R78618 VSS.n9772 VSS.n196 0.00953543
R78619 VSS.n9771 VSS.n201 0.00953543
R78620 VSS.n202 VSS.n195 0.00953543
R78621 VSS.n9777 VSS.n205 0.00953543
R78622 VSS.n1171 VSS.n753 0.00953543
R78623 VSS.n9401 VSS.n692 0.00953543
R78624 VSS.n5168 VSS.n5166 0.00951408
R78625 VSS.n7147 VSS.n2469 0.00943102
R78626 VSS.n1219 VSS.n1218 0.00934615
R78627 VSS.n9432 VSS.n9431 0.00934615
R78628 VSS.n2371 VSS.n2370 0.00934615
R78629 VSS.n9432 VSS.n9375 0.00934615
R78630 VSS.n2280 VSS.n2278 0.00934615
R78631 VSS.n2372 VSS.n2371 0.00934615
R78632 VSS.n2278 VSS.n2277 0.00934615
R78633 VSS.n1219 VSS.n1167 0.00934615
R78634 VSS.n8964 VSS.n8963 0.0091811
R78635 VSS.n2297 VSS.n2150 0.0091811
R78636 VSS.n8804 VSS.n1428 0.0091811
R78637 VSS.n8634 VSS.n1540 0.0091811
R78638 VSS.n8090 VSS.n8089 0.0091811
R78639 VSS.n1199 VSS.n737 0.0091811
R78640 VSS.n5718 VSS.n4223 0.00916197
R78641 VSS.n3742 VSS.n3140 0.00916197
R78642 VSS.n5713 VSS.n4022 0.00916197
R78643 VSS.n3755 VSS.n3170 0.00916197
R78644 VSS.n9 VSS.n5 0.00910927
R78645 VSS.n5732 VSS.n9 0.00910927
R78646 VSS.n7880 VSS.n8 0.00910927
R78647 VSS.n5732 VSS.n8 0.00910927
R78648 VSS.n8538 VSS.n1619 0.00898571
R78649 VSS.n6847 VSS.n2919 0.00898571
R78650 VSS.n6132 VSS.n4009 0.00898571
R78651 VSS.n5663 VSS.n4265 0.00898571
R78652 VSS.n5084 VSS.n4494 0.00898571
R78653 VSS.n2309 VSS.n2147 0.00882677
R78654 VSS.n2417 VSS.n1853 0.00882677
R78655 VSS.n1187 VSS.n734 0.00882677
R78656 VSS.n9385 VSS.n699 0.00882677
R78657 VSS.n9899 VSS.n16 0.00873944
R78658 VSS.n5668 VSS.n5667 0.00873944
R78659 VSS.n6614 VSS.n3160 0.00873944
R78660 VSS.n5178 VSS.n4434 0.00873944
R78661 VSS.n5665 VSS.n4261 0.00873944
R78662 VSS.n3167 VSS.n3163 0.00873944
R78663 VSS.n8816 VSS.n1376 0.00872857
R78664 VSS.n3008 VSS.n2941 0.00872857
R78665 VSS.n5723 VSS.n4221 0.00872857
R78666 VSS.n5352 VSS.n4246 0.00872857
R78667 VSS.n5018 VSS.n5017 0.00872857
R78668 VSS.n9837 DVSS 0.00852817
R78669 VSS.n4437 VSS.n4429 0.00852817
R78670 DVSS VSS.n125 0.00852817
R78671 VSS.n4757 VSS.n4742 0.00848752
R78672 VSS.n4745 VSS.n4742 0.00848752
R78673 VSS.n176 VSS.n173 0.00848752
R78674 VSS.n9814 VSS.n168 0.00848752
R78675 VSS.n173 VSS.n168 0.00848752
R78676 VSS.n4757 VSS.n4743 0.00848752
R78677 VSS.n4759 VSS.n4745 0.00848752
R78678 VSS.n9812 VSS.n176 0.00848752
R78679 VSS.n3861 VSS.n3858 0.00848752
R78680 VSS.n3863 VSS.n3861 0.00848752
R78681 VSS.n5469 VSS.n5440 0.00848752
R78682 VSS.n5472 VSS.n5468 0.00848752
R78683 VSS.n5468 VSS.n5440 0.00848752
R78684 VSS.n6253 VSS.n3858 0.00848752
R78685 VSS.n6251 VSS.n3863 0.00848752
R78686 VSS.n5469 VSS.n5466 0.00848752
R78687 VSS.n6258 VSS.n3853 0.00848752
R78688 VSS.n6256 VSS.n3853 0.00848752
R78689 VSS.n4151 VSS.n4148 0.00848752
R78690 VSS.n4155 VSS.n4152 0.00848752
R78691 VSS.n4152 VSS.n4151 0.00848752
R78692 VSS.n6260 VSS.n6258 0.00848752
R78693 VSS.n6256 VSS.n3854 0.00848752
R78694 VSS.n4157 VSS.n4148 0.00848752
R78695 VSS.n6267 VSS.n6266 0.00848752
R78696 VSS.n429 VSS.n426 0.00848752
R78697 VSS.n9603 VSS.n433 0.00848752
R78698 VSS.n433 VSS.n426 0.00848752
R78699 VSS.n9605 VSS.n429 0.00848752
R78700 VSS.n6266 VSS.n3829 0.00848752
R78701 VSS.n6278 VSS.n3825 0.00848752
R78702 VSS.n438 VSS.n435 0.00848752
R78703 VSS.n9598 VSS.n442 0.00848752
R78704 VSS.n442 VSS.n435 0.00848752
R78705 VSS.n9600 VSS.n438 0.00848752
R78706 VSS.n6282 VSS.n3825 0.00848752
R78707 VSS.n6577 VSS.n3227 0.00848752
R78708 VSS.n486 VSS.n483 0.00848752
R78709 VSS.n9590 VSS.n490 0.00848752
R78710 VSS.n490 VSS.n483 0.00848752
R78711 VSS.n9592 VSS.n486 0.00848752
R78712 VSS.n6581 VSS.n3227 0.00848752
R78713 VSS.n5775 VSS.n5770 0.00848752
R78714 VSS.n495 VSS.n492 0.00848752
R78715 VSS.n9585 VSS.n499 0.00848752
R78716 VSS.n499 VSS.n492 0.00848752
R78717 VSS.n9587 VSS.n495 0.00848752
R78718 VSS.n5779 VSS.n5770 0.00848752
R78719 VSS.n6969 VSS.n2771 0.00848752
R78720 VSS.n528 VSS.n525 0.00848752
R78721 VSS.n9577 VSS.n532 0.00848752
R78722 VSS.n532 VSS.n525 0.00848752
R78723 VSS.n9579 VSS.n528 0.00848752
R78724 VSS.n6973 VSS.n2771 0.00848752
R78725 VSS.n2313 VSS.n2162 0.00847244
R78726 VSS.n2413 VSS.n1848 0.00847244
R78727 VSS.n1183 VSS.n750 0.00847244
R78728 VSS.n9389 VSS.n695 0.00847244
R78729 VSS.n5657 VSS.n4258 0.0083169
R78730 VSS.n5662 VSS.n5656 0.0083169
R78731 VSS.n4706 VSS.n4705 0.0083169
R78732 VSS.n5233 VSS.n4341 0.0083169
R78733 VSS.n5207 VSS.n5206 0.0083169
R78734 VSS.n5171 VSS.n4454 0.00824648
R78735 VSS.n2293 VSS.n2158 0.00811811
R78736 VSS.n8244 VSS.n1863 0.00811811
R78737 VSS.n1203 VSS.n746 0.00811811
R78738 VSS.n9525 VSS.n709 0.00811811
R78739 VSS.n4458 VSS.n4450 0.00810563
R78740 VSS.n5119 VSS.n4426 0.00810563
R78741 VSS.n9883 VSS.n33 0.00803521
R78742 VSS.n9856 VSS.n82 0.00803521
R78743 VSS.n9841 VSS.n113 0.00803521
R78744 VSS.n3739 VSS.n3141 0.00789437
R78745 VSS.n3761 VSS.n3171 0.00789437
R78746 VSS.n7421 VSS 0.00782857
R78747 VSS.n9788 DVSS 0.00782857
R78748 VSS.n8893 DVSS 0.00782857
R78749 VSS.n1625 VSS.n1617 0.00782857
R78750 VSS.n8894 DVSS 0.00782857
R78751 VSS.n6682 DVSS 0.00782857
R78752 VSS.n2924 VSS.n2923 0.00782857
R78753 VSS.n6683 DVSS 0.00782857
R78754 DVSS VSS.n401 0.00782857
R78755 VSS.n4014 VSS.n4013 0.00782857
R78756 VSS.n9616 DVSS 0.00782857
R78757 DVSS VSS.n5425 0.00782857
R78758 VSS.n4271 VSS.n4262 0.00782857
R78759 VSS.n5493 DVSS 0.00782857
R78760 VSS.n4499 VSS.n4491 0.00782857
R78761 VSS.n9787 DVSS 0.00782857
R78762 VSS.n7683 VSS 0.00782857
R78763 VSS VSS.n0 0.00782857
R78764 VSS.n7420 VSS 0.00782857
R78765 VSS.n2166 VSS.n2143 0.00776378
R78766 VSS.n2397 VSS.n1857 0.00776378
R78767 VSS.n4760 VSS.n4586 0.00776378
R78768 VSS.n3865 VSS.n3857 0.00776378
R78769 VSS.n181 VSS.n170 0.00776378
R78770 VSS.n5470 VSS.n5436 0.00776378
R78771 VSS.n754 VSS.n730 0.00776378
R78772 VSS.n9405 VSS.n703 0.00776378
R78773 VSS.n8327 VSS.n1694 0.00763571
R78774 VSS.n8559 VSS.n1571 0.00763571
R78775 VSS.n8371 VSS.n1664 0.00763571
R78776 VSS.n6948 VSS.n2825 0.00763571
R78777 VSS.n6925 VSS.n2851 0.00763571
R78778 VSS.n6886 VSS.n2885 0.00763571
R78779 VSS.n6198 VSS.n6197 0.00763571
R78780 VSS.n6168 VSS.n3975 0.00763571
R78781 VSS.n5300 VSS.n5269 0.00763571
R78782 VSS.n5641 VSS.n4292 0.00763571
R78783 VSS.n4784 VSS.n4572 0.00763571
R78784 VSS.n5245 VSS.n4333 0.00763571
R78785 VSS.n5071 VSS.n4525 0.00763571
R78786 VSS.n8812 VSS.n1369 0.00757143
R78787 VSS.n3014 VSS.n2940 0.00757143
R78788 VSS.n4172 VSS.n4170 0.00757143
R78789 VSS.n5589 VSS.n4245 0.00757143
R78790 VSS.n4975 VSS.n4872 0.00757143
R78791 VSS.n3727 VSS.n3151 0.00747183
R78792 VSS.n6796 VSS.n2944 0.00747183
R78793 VSS.n3785 VSS.n3181 0.00747183
R78794 VSS.n6797 VSS.n2926 0.00747183
R78795 VSS.n9863 VSS.n79 0.00740945
R78796 VSS.n2271 VSS.n2154 0.00740945
R78797 VSS.n2387 VSS.n1842 0.00740945
R78798 VSS.n4704 VSS.n4628 0.00740945
R78799 VSS.n9896 VSS.n25 0.00740945
R78800 VSS.n5205 VSS.n4391 0.00740945
R78801 VSS.n5232 VSS.n4354 0.00740945
R78802 VSS.n4719 VSS.n4603 0.00740945
R78803 VSS.n3837 VSS.n3832 0.00740945
R78804 VSS.n9833 VSS.n141 0.00740945
R78805 VSS.n422 VSS.n408 0.00740945
R78806 VSS.n9848 VSS.n110 0.00740945
R78807 VSS.n1220 VSS.n741 0.00740945
R78808 VSS.n9415 VSS.n689 0.00740945
R78809 VSS.n8494 VSS.n1323 0.00737857
R78810 VSS.n8868 VSS.n1284 0.00737857
R78811 VSS.n8905 VSS.n8901 0.00737857
R78812 VSS.n6742 VSS.n2973 0.00737857
R78813 VSS.n3087 VSS.n3081 0.00737857
R78814 VSS.n6694 VSS.n6690 0.00737857
R78815 VSS.n9671 VSS.n309 0.00737857
R78816 VSS.n9644 VSS.n9643 0.00737857
R78817 VSS.n9626 VSS.n9623 0.00737857
R78818 VSS.n5366 VSS.n288 0.00737857
R78819 VSS.n5522 VSS.n5521 0.00737857
R78820 VSS.n5503 VSS.n5500 0.00737857
R78821 VSS.n9696 VSS.n246 0.00737857
R78822 VSS.n9739 VSS.n227 0.00737857
R78823 VSS.n9778 VSS.n190 0.00737857
R78824 VSS.n5177 VSS.n4439 0.00726056
R78825 VSS.n7860 VSS.n7282 0.00725
R78826 VSS.n7320 VSS.n7287 0.00725
R78827 VSS.n4609 VSS.n4608 0.00716667
R78828 VSS.n4610 VSS.n4609 0.00716667
R78829 VSS.n4613 VSS.n4610 0.00716667
R78830 VSS.n4614 VSS.n4613 0.00716667
R78831 VSS.n4615 VSS.n4614 0.00716667
R78832 VSS.n4616 VSS.n4615 0.00716667
R78833 VSS.n4681 VSS.n4616 0.00716667
R78834 VSS.n4682 VSS.n4681 0.00716667
R78835 VSS.n4683 VSS.n4682 0.00716667
R78836 VSS.n4684 VSS.n4683 0.00716667
R78837 VSS.n4687 VSS.n4684 0.00716667
R78838 VSS.n4688 VSS.n4687 0.00716667
R78839 VSS.n4689 VSS.n4688 0.00716667
R78840 VSS.n4691 VSS.n4689 0.00716667
R78841 VSS.n4691 VSS.n4690 0.00716667
R78842 VSS.n4690 VSS.n4359 0.00716667
R78843 VSS.n4360 VSS.n4359 0.00716667
R78844 VSS.n4361 VSS.n4360 0.00716667
R78845 VSS.n4364 VSS.n4361 0.00716667
R78846 VSS.n4365 VSS.n4364 0.00716667
R78847 VSS.n4366 VSS.n4365 0.00716667
R78848 VSS.n4367 VSS.n4366 0.00716667
R78849 VSS.n4370 VSS.n4367 0.00716667
R78850 VSS.n4371 VSS.n4370 0.00716667
R78851 VSS.n4372 VSS.n4371 0.00716667
R78852 VSS.n4373 VSS.n4372 0.00716667
R78853 VSS.n4376 VSS.n4373 0.00716667
R78854 VSS.n4377 VSS.n4376 0.00716667
R78855 VSS.n4378 VSS.n4377 0.00716667
R78856 VSS.n4379 VSS.n4378 0.00716667
R78857 VSS.n4401 VSS.n4379 0.00716667
R78858 VSS.n4402 VSS.n4401 0.00716667
R78859 VSS.n4403 VSS.n4402 0.00716667
R78860 VSS.n4404 VSS.n4403 0.00716667
R78861 VSS.n4407 VSS.n4404 0.00716667
R78862 VSS.n4408 VSS.n4407 0.00716667
R78863 VSS.n4409 VSS.n4408 0.00716667
R78864 VSS.n4410 VSS.n4409 0.00716667
R78865 VSS.n4413 VSS.n4410 0.00716667
R78866 VSS.n4414 VSS.n4413 0.00716667
R78867 VSS.n4415 VSS.n4414 0.00716667
R78868 VSS.n4416 VSS.n4415 0.00716667
R78869 VSS.n4419 VSS.n4416 0.00716667
R78870 VSS.n4420 VSS.n4419 0.00716667
R78871 VSS.n4421 VSS.n4420 0.00716667
R78872 VSS.n4422 VSS.n4421 0.00716667
R78873 VSS.n4442 VSS.n4422 0.00716667
R78874 VSS.n4443 VSS.n4442 0.00716667
R78875 VSS.n4444 VSS.n4443 0.00716667
R78876 VSS.n4445 VSS.n4444 0.00716667
R78877 VSS.n4446 VSS.n4445 0.00716667
R78878 VSS.n5128 VSS.n4446 0.00716667
R78879 VSS.n5129 VSS.n5128 0.00716667
R78880 VSS.n5130 VSS.n5129 0.00716667
R78881 VSS.n5131 VSS.n5130 0.00716667
R78882 VSS.n5134 VSS.n5131 0.00716667
R78883 VSS.n5135 VSS.n5134 0.00716667
R78884 VSS.n5136 VSS.n5135 0.00716667
R78885 VSS.n5137 VSS.n5136 0.00716667
R78886 VSS.n5140 VSS.n5137 0.00716667
R78887 VSS.n5141 VSS.n5140 0.00716667
R78888 VSS.n5142 VSS.n5141 0.00716667
R78889 VSS.n5143 VSS.n5142 0.00716667
R78890 VSS.n5144 VSS.n5143 0.00716667
R78891 VSS.n5146 VSS.n5144 0.00716667
R78892 VSS.n5146 VSS.n5145 0.00716667
R78893 VSS.n5145 VSS.n47 0.00716667
R78894 VSS.n48 VSS.n47 0.00716667
R78895 VSS.n49 VSS.n48 0.00716667
R78896 VSS.n52 VSS.n49 0.00716667
R78897 VSS.n53 VSS.n52 0.00716667
R78898 VSS.n54 VSS.n53 0.00716667
R78899 VSS.n55 VSS.n54 0.00716667
R78900 VSS.n58 VSS.n55 0.00716667
R78901 VSS.n59 VSS.n58 0.00716667
R78902 VSS.n60 VSS.n59 0.00716667
R78903 VSS.n61 VSS.n60 0.00716667
R78904 VSS.n64 VSS.n61 0.00716667
R78905 VSS.n65 VSS.n64 0.00716667
R78906 VSS.n66 VSS.n65 0.00716667
R78907 VSS.n67 VSS.n66 0.00716667
R78908 VSS.n89 VSS.n67 0.00716667
R78909 VSS.n90 VSS.n89 0.00716667
R78910 VSS.n91 VSS.n90 0.00716667
R78911 VSS.n92 VSS.n91 0.00716667
R78912 VSS.n95 VSS.n92 0.00716667
R78913 VSS.n96 VSS.n95 0.00716667
R78914 VSS.n97 VSS.n96 0.00716667
R78915 VSS.n98 VSS.n97 0.00716667
R78916 VSS.n120 VSS.n98 0.00716667
R78917 VSS.n121 VSS.n120 0.00716667
R78918 VSS.n122 VSS.n121 0.00716667
R78919 VSS.n123 VSS.n122 0.00716667
R78920 VSS.n126 VSS.n123 0.00716667
R78921 VSS.n127 VSS.n126 0.00716667
R78922 VSS.n128 VSS.n127 0.00716667
R78923 VSS.n129 VSS.n128 0.00716667
R78924 VSS.n9824 VSS.n9823 0.00716667
R78925 VSS.n4743 VSS.n3855 0.00716667
R78926 VSS.n9815 VSS.n9814 0.00716667
R78927 VSS.n6254 VSS.n6253 0.00716667
R78928 VSS.n5472 VSS.n167 0.00716667
R78929 VSS.n6260 VSS.n6255 0.00716667
R78930 VSS.n4155 VSS.n4154 0.00716667
R78931 VSS.n6273 VSS.n3830 0.00716667
R78932 VSS.n9603 VSS.n434 0.00716667
R78933 VSS.n6280 VSS.n3827 0.00716667
R78934 VSS.n9598 VSS.n443 0.00716667
R78935 VSS.n6579 VSS.n3230 0.00716667
R78936 VSS.n9590 VSS.n491 0.00716667
R78937 VSS.n5777 VSS.n5772 0.00716667
R78938 VSS.n9585 VSS.n500 0.00716667
R78939 VSS.n6971 VSS.n2795 0.00716667
R78940 VSS.n9577 VSS.n533 0.00716667
R78941 VSS.n2283 VSS.n2153 0.00705512
R78942 VSS.n2381 VSS.n1841 0.00705512
R78943 VSS.n6257 VSS.n3838 0.00705512
R78944 VSS.n4153 VSS.n409 0.00705512
R78945 VSS.n1213 VSS.n740 0.00705512
R78946 VSS.n9421 VSS.n688 0.00705512
R78947 VSS.n4867 VSS.n4866 0.0070493
R78948 VSS.n3731 VSS.n3153 0.0070493
R78949 VSS.n6784 VSS.n2946 0.0070493
R78950 VSS.n4864 VSS.n4501 0.0070493
R78951 VSS.n3777 VSS.n3183 0.0070493
R78952 VSS.n6785 VSS.n2928 0.0070493
R78953 VSS.n4718 VSS.n4595 0.0070493
R78954 VSS.n4703 VSS.n4623 0.0070493
R78955 VSS.n5231 VSS.n4346 0.0070493
R78956 VSS.n5204 VSS.n4386 0.0070493
R78957 VSS.n9823 DVSS 0.00697887
R78958 VSS.n5172 VSS.n4448 0.00697887
R78959 VSS.n7882 VSS.n7881 0.00678019
R78960 VSS.n7886 VSS.n7885 0.00678019
R78961 VSS.n9892 VSS.n35 0.00676761
R78962 VSS.n9885 VSS.n34 0.00676761
R78963 VSS.n9865 VSS.n9864 0.00676761
R78964 VSS.n9858 VSS.n85 0.00676761
R78965 VSS.n9850 VSS.n9849 0.00676761
R78966 VSS.n9843 VSS.n116 0.00676761
R78967 VSS.n9835 VSS.n9834 0.00676761
R78968 VSS.n9826 VSS.n9822 0.00676761
R78969 VSS.n2323 VSS.n2144 0.00670079
R78970 VSS.n2403 VSS.n1856 0.00670079
R78971 VSS.n4727 VSS.n4585 0.00670079
R78972 VSS.n6252 VSS.n3860 0.00670079
R78973 VSS.n9811 VSS.n9810 0.00670079
R78974 VSS.n5473 VSS.n5435 0.00670079
R78975 VSS.n1173 VSS.n731 0.00670079
R78976 VSS.n9399 VSS.n702 0.00670079
R78977 VSS.n8535 VSS.n1634 0.00667143
R78978 VSS.n6841 VSS.n6840 0.00667143
R78979 VSS.n6126 VSS.n6125 0.00667143
R78980 VSS.n5596 VSS.n4264 0.00667143
R78981 VSS.n5026 VSS.n4493 0.00667143
R78982 VSS.n4853 VSS.n4489 0.00662676
R78983 VSS.n3735 VSS.n3143 0.00662676
R78984 VSS.n2955 VSS.n2949 0.00662676
R78985 VSS.n5086 VSS.n5085 0.00662676
R78986 VSS.n3769 VSS.n3173 0.00662676
R78987 VSS.n6773 VSS.n2931 0.00662676
R78988 VSS.n7307 VSS.n7306 0.00658571
R78989 VSS.n7308 VSS.n7307 0.00658571
R78990 VSS.n7308 VSS.n7296 0.00658571
R78991 VSS.n7314 VSS.n7296 0.00658571
R78992 VSS.n7315 VSS.n7314 0.00658571
R78993 VSS.n7316 VSS.n7315 0.00658571
R78994 VSS.n7316 VSS.n7292 0.00658571
R78995 VSS.n7322 VSS.n7292 0.00658571
R78996 VSS.n7323 VSS.n7322 0.00658571
R78997 VSS.n7592 VSS.n7323 0.00658571
R78998 VSS.n7592 VSS.n7591 0.00658571
R78999 VSS.n7591 VSS.n7590 0.00658571
R79000 VSS.n7590 VSS.n7324 0.00658571
R79001 VSS.n7584 VSS.n7324 0.00658571
R79002 VSS.n7584 VSS.n7583 0.00658571
R79003 VSS.n7583 VSS.n7582 0.00658571
R79004 VSS.n7582 VSS.n7328 0.00658571
R79005 VSS.n7576 VSS.n7328 0.00658571
R79006 VSS.n7576 VSS.n7575 0.00658571
R79007 VSS.n7575 VSS.n7574 0.00658571
R79008 VSS.n7574 VSS.n7332 0.00658571
R79009 VSS.n7568 VSS.n7332 0.00658571
R79010 VSS.n7568 VSS.n7567 0.00658571
R79011 VSS.n7567 VSS.n7566 0.00658571
R79012 VSS.n7566 VSS.n7336 0.00658571
R79013 VSS.n7560 VSS.n7336 0.00658571
R79014 VSS.n7560 VSS.n7559 0.00658571
R79015 VSS.n7559 VSS.n7558 0.00658571
R79016 VSS.n7558 VSS.n7340 0.00658571
R79017 VSS.n7552 VSS.n7340 0.00658571
R79018 VSS.n7552 VSS.n7551 0.00658571
R79019 VSS.n7551 VSS.n7550 0.00658571
R79020 VSS.n7550 VSS.n7344 0.00658571
R79021 VSS.n7544 VSS.n7344 0.00658571
R79022 VSS.n7544 VSS.n7543 0.00658571
R79023 VSS.n7543 VSS.n7542 0.00658571
R79024 VSS.n7542 VSS.n7348 0.00658571
R79025 VSS.n7536 VSS.n7348 0.00658571
R79026 VSS.n7536 VSS.n7535 0.00658571
R79027 VSS.n7535 VSS.n7534 0.00658571
R79028 VSS.n7534 VSS.n7352 0.00658571
R79029 VSS.n7528 VSS.n7352 0.00658571
R79030 VSS.n7528 VSS.n7527 0.00658571
R79031 VSS.n7527 VSS.n7526 0.00658571
R79032 VSS.n7526 VSS.n7356 0.00658571
R79033 VSS.n7520 VSS.n7356 0.00658571
R79034 VSS.n7520 VSS.n7519 0.00658571
R79035 VSS.n7519 VSS.n7518 0.00658571
R79036 VSS.n7518 VSS.n7360 0.00658571
R79037 VSS.n7512 VSS.n7360 0.00658571
R79038 VSS.n7512 VSS.n7511 0.00658571
R79039 VSS.n7511 VSS.n7510 0.00658571
R79040 VSS.n7510 VSS.n7364 0.00658571
R79041 VSS.n7504 VSS.n7364 0.00658571
R79042 VSS.n7504 VSS.n7503 0.00658571
R79043 VSS.n7503 VSS.n7502 0.00658571
R79044 VSS.n7502 VSS.n7368 0.00658571
R79045 VSS.n7496 VSS.n7368 0.00658571
R79046 VSS.n7496 VSS.n7495 0.00658571
R79047 VSS.n7495 VSS.n7494 0.00658571
R79048 VSS.n7494 VSS.n7372 0.00658571
R79049 VSS.n7488 VSS.n7372 0.00658571
R79050 VSS.n7488 VSS.n7487 0.00658571
R79051 VSS.n7487 VSS.n7486 0.00658571
R79052 VSS.n7486 VSS.n7376 0.00658571
R79053 VSS.n7480 VSS.n7376 0.00658571
R79054 VSS.n7480 VSS.n7479 0.00658571
R79055 VSS.n7479 VSS.n7478 0.00658571
R79056 VSS.n7478 VSS.n7380 0.00658571
R79057 VSS.n7472 VSS.n7380 0.00658571
R79058 VSS.n7472 VSS.n7471 0.00658571
R79059 VSS.n7471 VSS.n7470 0.00658571
R79060 VSS.n7470 VSS.n7384 0.00658571
R79061 VSS.n7464 VSS.n7384 0.00658571
R79062 VSS.n7464 VSS.n7463 0.00658571
R79063 VSS.n7463 VSS.n7462 0.00658571
R79064 VSS.n7462 VSS.n7388 0.00658571
R79065 VSS.n7456 VSS.n7388 0.00658571
R79066 VSS.n7456 VSS.n7455 0.00658571
R79067 VSS.n7455 VSS.n7454 0.00658571
R79068 VSS.n7454 VSS.n7392 0.00658571
R79069 VSS.n7448 VSS.n7392 0.00658571
R79070 VSS.n7448 VSS.n7447 0.00658571
R79071 VSS.n7447 VSS.n7446 0.00658571
R79072 VSS.n7446 VSS.n7396 0.00658571
R79073 VSS.n7440 VSS.n7396 0.00658571
R79074 VSS.n7440 VSS.n7439 0.00658571
R79075 VSS.n7439 VSS.n7438 0.00658571
R79076 VSS.n7438 VSS.n7400 0.00658571
R79077 VSS.n7432 VSS.n7400 0.00658571
R79078 VSS.n7432 VSS.n7431 0.00658571
R79079 VSS.n7431 VSS.n7430 0.00658571
R79080 VSS.n7430 VSS.n7404 0.00658571
R79081 VSS.n7424 VSS.n7404 0.00658571
R79082 VSS.n7424 VSS.n7423 0.00658571
R79083 VSS.n7423 VSS.n7422 0.00658571
R79084 VSS.n7422 VSS.n7408 0.00658571
R79085 VSS.n7416 VSS.n7415 0.00658571
R79086 VSS.n4767 VSS.n4582 0.00658571
R79087 VSS.n4768 VSS.n4767 0.00658571
R79088 VSS.n4769 VSS.n4768 0.00658571
R79089 VSS.n4769 VSS.n4578 0.00658571
R79090 VSS.n4775 VSS.n4578 0.00658571
R79091 VSS.n4776 VSS.n4775 0.00658571
R79092 VSS.n4777 VSS.n4776 0.00658571
R79093 VSS.n4777 VSS.n4550 0.00658571
R79094 VSS.n4789 VSS.n4550 0.00658571
R79095 VSS.n4790 VSS.n4789 0.00658571
R79096 VSS.n4791 VSS.n4790 0.00658571
R79097 VSS.n4791 VSS.n4546 0.00658571
R79098 VSS.n4797 VSS.n4546 0.00658571
R79099 VSS.n4798 VSS.n4797 0.00658571
R79100 VSS.n4799 VSS.n4798 0.00658571
R79101 VSS.n4799 VSS.n4544 0.00658571
R79102 VSS.n4805 VSS.n4544 0.00658571
R79103 VSS.n4806 VSS.n4805 0.00658571
R79104 VSS.n4807 VSS.n4806 0.00658571
R79105 VSS.n4807 VSS.n4540 0.00658571
R79106 VSS.n4813 VSS.n4540 0.00658571
R79107 VSS.n4814 VSS.n4813 0.00658571
R79108 VSS.n4815 VSS.n4814 0.00658571
R79109 VSS.n4815 VSS.n4536 0.00658571
R79110 VSS.n4821 VSS.n4536 0.00658571
R79111 VSS.n4822 VSS.n4821 0.00658571
R79112 VSS.n4823 VSS.n4822 0.00658571
R79113 VSS.n4823 VSS.n4532 0.00658571
R79114 VSS.n4829 VSS.n4532 0.00658571
R79115 VSS.n4830 VSS.n4829 0.00658571
R79116 VSS.n5058 VSS.n4830 0.00658571
R79117 VSS.n5058 VSS.n5057 0.00658571
R79118 VSS.n5057 VSS.n5056 0.00658571
R79119 VSS.n5056 VSS.n4831 0.00658571
R79120 VSS.n4835 VSS.n4831 0.00658571
R79121 VSS.n5048 VSS.n4835 0.00658571
R79122 VSS.n5048 VSS.n5047 0.00658571
R79123 VSS.n5047 VSS.n5046 0.00658571
R79124 VSS.n5046 VSS.n4836 0.00658571
R79125 VSS.n5040 VSS.n4836 0.00658571
R79126 VSS.n5040 VSS.n5039 0.00658571
R79127 VSS.n5039 VSS.n5038 0.00658571
R79128 VSS.n5038 VSS.n4840 0.00658571
R79129 VSS.n5032 VSS.n4840 0.00658571
R79130 VSS.n5032 VSS.n5031 0.00658571
R79131 VSS.n5031 VSS.n5030 0.00658571
R79132 VSS.n5030 VSS.n4844 0.00658571
R79133 VSS.n5025 VSS.n4844 0.00658571
R79134 VSS.n5025 VSS.n5024 0.00658571
R79135 VSS.n5024 VSS.n5023 0.00658571
R79136 VSS.n5023 VSS.n4846 0.00658571
R79137 VSS.n4979 VSS.n4846 0.00658571
R79138 VSS.n5015 VSS.n4979 0.00658571
R79139 VSS.n5015 VSS.n5014 0.00658571
R79140 VSS.n5014 VSS.n5013 0.00658571
R79141 VSS.n5013 VSS.n4980 0.00658571
R79142 VSS.n5007 VSS.n4980 0.00658571
R79143 VSS.n5007 VSS.n5006 0.00658571
R79144 VSS.n5006 VSS.n5005 0.00658571
R79145 VSS.n5005 VSS.n4984 0.00658571
R79146 VSS.n4999 VSS.n4984 0.00658571
R79147 VSS.n4999 VSS.n4998 0.00658571
R79148 VSS.n4998 VSS.n4997 0.00658571
R79149 VSS.n4997 VSS.n4988 0.00658571
R79150 VSS.n4991 VSS.n4988 0.00658571
R79151 VSS.n4991 VSS.n4990 0.00658571
R79152 VSS.n4990 VSS.n248 0.00658571
R79153 VSS.n9699 VSS.n248 0.00658571
R79154 VSS.n9700 VSS.n9699 0.00658571
R79155 VSS.n9701 VSS.n9700 0.00658571
R79156 VSS.n9701 VSS.n244 0.00658571
R79157 VSS.n9707 VSS.n244 0.00658571
R79158 VSS.n9708 VSS.n9707 0.00658571
R79159 VSS.n9709 VSS.n9708 0.00658571
R79160 VSS.n9709 VSS.n240 0.00658571
R79161 VSS.n9715 VSS.n240 0.00658571
R79162 VSS.n9716 VSS.n9715 0.00658571
R79163 VSS.n9717 VSS.n9716 0.00658571
R79164 VSS.n9717 VSS.n236 0.00658571
R79165 VSS.n9723 VSS.n236 0.00658571
R79166 VSS.n9724 VSS.n9723 0.00658571
R79167 VSS.n9745 VSS.n9724 0.00658571
R79168 VSS.n9745 VSS.n9744 0.00658571
R79169 VSS.n9744 VSS.n9743 0.00658571
R79170 VSS.n9743 VSS.n9725 0.00658571
R79171 VSS.n9729 VSS.n9725 0.00658571
R79172 VSS.n9735 VSS.n9729 0.00658571
R79173 VSS.n9735 VSS.n9734 0.00658571
R79174 VSS.n9734 VSS.n9733 0.00658571
R79175 VSS.n9733 VSS.n9730 0.00658571
R79176 VSS.n9730 VSS.n192 0.00658571
R79177 VSS.n9781 VSS.n192 0.00658571
R79178 VSS.n9782 VSS.n9781 0.00658571
R79179 VSS.n9783 VSS.n9782 0.00658571
R79180 VSS.n9783 VSS.n188 0.00658571
R79181 VSS.n9789 VSS.n188 0.00658571
R79182 VSS.n9790 VSS.n9789 0.00658571
R79183 VSS.n9795 VSS.n9794 0.00658571
R79184 VSS.n8304 VSS.n1704 0.00658571
R79185 VSS.n8305 VSS.n8304 0.00658571
R79186 VSS.n8306 VSS.n8305 0.00658571
R79187 VSS.n8306 VSS.n1700 0.00658571
R79188 VSS.n8312 VSS.n1700 0.00658571
R79189 VSS.n8313 VSS.n8312 0.00658571
R79190 VSS.n8314 VSS.n8313 0.00658571
R79191 VSS.n8314 VSS.n1684 0.00658571
R79192 VSS.n8333 VSS.n1684 0.00658571
R79193 VSS.n8334 VSS.n8333 0.00658571
R79194 VSS.n8335 VSS.n8334 0.00658571
R79195 VSS.n8335 VSS.n1680 0.00658571
R79196 VSS.n8341 VSS.n1680 0.00658571
R79197 VSS.n8342 VSS.n8341 0.00658571
R79198 VSS.n8343 VSS.n8342 0.00658571
R79199 VSS.n8343 VSS.n1678 0.00658571
R79200 VSS.n8349 VSS.n1678 0.00658571
R79201 VSS.n8350 VSS.n8349 0.00658571
R79202 VSS.n8351 VSS.n8350 0.00658571
R79203 VSS.n8351 VSS.n1674 0.00658571
R79204 VSS.n8357 VSS.n1674 0.00658571
R79205 VSS.n8358 VSS.n8357 0.00658571
R79206 VSS.n8359 VSS.n8358 0.00658571
R79207 VSS.n8359 VSS.n1670 0.00658571
R79208 VSS.n8365 VSS.n1670 0.00658571
R79209 VSS.n8366 VSS.n8365 0.00658571
R79210 VSS.n8367 VSS.n8366 0.00658571
R79211 VSS.n8367 VSS.n1666 0.00658571
R79212 VSS.n8374 VSS.n1666 0.00658571
R79213 VSS.n8375 VSS.n8374 0.00658571
R79214 VSS.n8376 VSS.n8375 0.00658571
R79215 VSS.n8376 VSS.n1653 0.00658571
R79216 VSS.n8415 VSS.n1653 0.00658571
R79217 VSS.n8416 VSS.n8415 0.00658571
R79218 VSS.n8417 VSS.n8416 0.00658571
R79219 VSS.n8417 VSS.n1649 0.00658571
R79220 VSS.n8423 VSS.n1649 0.00658571
R79221 VSS.n8424 VSS.n8423 0.00658571
R79222 VSS.n8425 VSS.n8424 0.00658571
R79223 VSS.n8425 VSS.n1645 0.00658571
R79224 VSS.n8431 VSS.n1645 0.00658571
R79225 VSS.n8432 VSS.n8431 0.00658571
R79226 VSS.n8434 VSS.n8432 0.00658571
R79227 VSS.n8434 VSS.n8433 0.00658571
R79228 VSS.n8433 VSS.n1642 0.00658571
R79229 VSS.n1642 VSS.n1640 0.00658571
R79230 VSS.n8442 VSS.n1640 0.00658571
R79231 VSS.n8443 VSS.n8442 0.00658571
R79232 VSS.n8532 VSS.n8443 0.00658571
R79233 VSS.n8532 VSS.n8531 0.00658571
R79234 VSS.n8531 VSS.n8530 0.00658571
R79235 VSS.n8530 VSS.n8444 0.00658571
R79236 VSS.n8526 VSS.n8444 0.00658571
R79237 VSS.n8526 VSS.n8525 0.00658571
R79238 VSS.n8525 VSS.n8524 0.00658571
R79239 VSS.n8524 VSS.n8446 0.00658571
R79240 VSS.n8518 VSS.n8446 0.00658571
R79241 VSS.n8518 VSS.n8517 0.00658571
R79242 VSS.n8517 VSS.n8516 0.00658571
R79243 VSS.n8516 VSS.n8451 0.00658571
R79244 VSS.n8510 VSS.n8451 0.00658571
R79245 VSS.n8510 VSS.n8509 0.00658571
R79246 VSS.n8509 VSS.n8508 0.00658571
R79247 VSS.n8508 VSS.n8455 0.00658571
R79248 VSS.n8502 VSS.n8455 0.00658571
R79249 VSS.n8502 VSS.n8501 0.00658571
R79250 VSS.n8501 VSS.n8500 0.00658571
R79251 VSS.n8500 VSS.n8457 0.00658571
R79252 VSS.n8459 VSS.n8457 0.00658571
R79253 VSS.n8462 VSS.n8459 0.00658571
R79254 VSS.n8490 VSS.n8462 0.00658571
R79255 VSS.n8490 VSS.n8489 0.00658571
R79256 VSS.n8489 VSS.n8488 0.00658571
R79257 VSS.n8488 VSS.n8463 0.00658571
R79258 VSS.n8482 VSS.n8463 0.00658571
R79259 VSS.n8482 VSS.n8481 0.00658571
R79260 VSS.n8481 VSS.n8480 0.00658571
R79261 VSS.n8480 VSS.n8467 0.00658571
R79262 VSS.n8474 VSS.n8467 0.00658571
R79263 VSS.n8474 VSS.n8473 0.00658571
R79264 VSS.n8473 VSS.n8472 0.00658571
R79265 VSS.n8472 VSS.n1286 0.00658571
R79266 VSS.n8864 VSS.n1286 0.00658571
R79267 VSS.n8865 VSS.n8864 0.00658571
R79268 VSS.n8866 VSS.n8865 0.00658571
R79269 VSS.n8866 VSS.n1282 0.00658571
R79270 VSS.n8873 VSS.n1282 0.00658571
R79271 VSS.n8874 VSS.n8873 0.00658571
R79272 VSS.n8875 VSS.n8874 0.00658571
R79273 VSS.n8875 VSS.n1280 0.00658571
R79274 VSS.n8880 VSS.n1280 0.00658571
R79275 VSS.n8881 VSS.n8880 0.00658571
R79276 VSS.n8899 VSS.n8881 0.00658571
R79277 VSS.n8899 VSS.n8898 0.00658571
R79278 VSS.n8898 VSS.n8897 0.00658571
R79279 VSS.n8897 VSS.n8882 0.00658571
R79280 VSS.n8891 VSS.n8882 0.00658571
R79281 VSS.n8890 VSS.n8889 0.00658571
R79282 VSS.n2822 VSS.n2821 0.00658571
R79283 VSS.n6954 VSS.n2822 0.00658571
R79284 VSS.n6954 VSS.n6953 0.00658571
R79285 VSS.n6953 VSS.n6952 0.00658571
R79286 VSS.n6952 VSS.n2823 0.00658571
R79287 VSS.n6946 VSS.n2823 0.00658571
R79288 VSS.n6946 VSS.n6945 0.00658571
R79289 VSS.n6945 VSS.n6944 0.00658571
R79290 VSS.n6944 VSS.n2827 0.00658571
R79291 VSS.n6931 VSS.n2827 0.00658571
R79292 VSS.n6931 VSS.n6930 0.00658571
R79293 VSS.n6930 VSS.n6929 0.00658571
R79294 VSS.n6929 VSS.n2849 0.00658571
R79295 VSS.n6923 VSS.n2849 0.00658571
R79296 VSS.n6923 VSS.n6922 0.00658571
R79297 VSS.n6922 VSS.n6921 0.00658571
R79298 VSS.n6921 VSS.n2853 0.00658571
R79299 VSS.n6908 VSS.n2853 0.00658571
R79300 VSS.n6908 VSS.n6907 0.00658571
R79301 VSS.n6907 VSS.n6906 0.00658571
R79302 VSS.n6906 VSS.n2875 0.00658571
R79303 VSS.n6900 VSS.n2875 0.00658571
R79304 VSS.n6900 VSS.n6899 0.00658571
R79305 VSS.n6899 VSS.n6898 0.00658571
R79306 VSS.n6898 VSS.n2879 0.00658571
R79307 VSS.n6892 VSS.n2879 0.00658571
R79308 VSS.n6892 VSS.n6891 0.00658571
R79309 VSS.n6891 VSS.n6890 0.00658571
R79310 VSS.n6890 VSS.n2883 0.00658571
R79311 VSS.n6884 VSS.n2883 0.00658571
R79312 VSS.n6884 VSS.n6883 0.00658571
R79313 VSS.n6883 VSS.n6882 0.00658571
R79314 VSS.n6882 VSS.n2887 0.00658571
R79315 VSS.n6869 VSS.n2887 0.00658571
R79316 VSS.n6869 VSS.n6868 0.00658571
R79317 VSS.n6868 VSS.n6867 0.00658571
R79318 VSS.n6867 VSS.n2909 0.00658571
R79319 VSS.n6861 VSS.n2909 0.00658571
R79320 VSS.n6861 VSS.n6860 0.00658571
R79321 VSS.n6860 VSS.n6859 0.00658571
R79322 VSS.n6859 VSS.n2913 0.00658571
R79323 VSS.n6853 VSS.n2913 0.00658571
R79324 VSS.n6853 VSS.n6852 0.00658571
R79325 VSS.n6852 VSS.n6851 0.00658571
R79326 VSS.n6851 VSS.n2917 0.00658571
R79327 VSS.n6845 VSS.n2917 0.00658571
R79328 VSS.n6845 VSS.n6844 0.00658571
R79329 VSS.n6844 VSS.n6843 0.00658571
R79330 VSS.n6843 VSS.n2921 0.00658571
R79331 VSS.n3011 VSS.n2921 0.00658571
R79332 VSS.n3011 VSS.n3010 0.00658571
R79333 VSS.n3016 VSS.n3010 0.00658571
R79334 VSS.n3017 VSS.n3016 0.00658571
R79335 VSS.n3018 VSS.n3017 0.00658571
R79336 VSS.n3018 VSS.n3006 0.00658571
R79337 VSS.n3024 VSS.n3006 0.00658571
R79338 VSS.n3025 VSS.n3024 0.00658571
R79339 VSS.n3026 VSS.n3025 0.00658571
R79340 VSS.n3026 VSS.n3002 0.00658571
R79341 VSS.n3032 VSS.n3002 0.00658571
R79342 VSS.n3033 VSS.n3032 0.00658571
R79343 VSS.n3035 VSS.n3033 0.00658571
R79344 VSS.n3035 VSS.n3034 0.00658571
R79345 VSS.n3034 VSS.n2998 0.00658571
R79346 VSS.n3042 VSS.n2998 0.00658571
R79347 VSS.n3043 VSS.n3042 0.00658571
R79348 VSS.n6746 VSS.n3043 0.00658571
R79349 VSS.n6746 VSS.n6745 0.00658571
R79350 VSS.n6745 VSS.n6744 0.00658571
R79351 VSS.n6744 VSS.n3044 0.00658571
R79352 VSS.n6738 VSS.n3044 0.00658571
R79353 VSS.n6738 VSS.n6737 0.00658571
R79354 VSS.n6737 VSS.n6736 0.00658571
R79355 VSS.n6736 VSS.n3048 0.00658571
R79356 VSS.n6730 VSS.n3048 0.00658571
R79357 VSS.n6730 VSS.n6729 0.00658571
R79358 VSS.n6729 VSS.n6728 0.00658571
R79359 VSS.n6728 VSS.n3052 0.00658571
R79360 VSS.n6722 VSS.n3052 0.00658571
R79361 VSS.n6722 VSS.n6721 0.00658571
R79362 VSS.n6721 VSS.n6720 0.00658571
R79363 VSS.n6720 VSS.n3056 0.00658571
R79364 VSS.n3084 VSS.n3056 0.00658571
R79365 VSS.n6712 VSS.n3084 0.00658571
R79366 VSS.n6712 VSS.n6711 0.00658571
R79367 VSS.n6711 VSS.n6710 0.00658571
R79368 VSS.n6710 VSS.n3085 0.00658571
R79369 VSS.n6704 VSS.n3085 0.00658571
R79370 VSS.n6704 VSS.n6703 0.00658571
R79371 VSS.n6703 VSS.n6702 0.00658571
R79372 VSS.n6702 VSS.n3090 0.00658571
R79373 VSS.n6670 VSS.n3090 0.00658571
R79374 VSS.n6688 VSS.n6670 0.00658571
R79375 VSS.n6688 VSS.n6687 0.00658571
R79376 VSS.n6687 VSS.n6686 0.00658571
R79377 VSS.n6686 VSS.n6671 0.00658571
R79378 VSS.n6680 VSS.n6671 0.00658571
R79379 VSS.n6679 VSS.n6678 0.00658571
R79380 VSS.n3921 VSS.n3915 0.00658571
R79381 VSS.n3922 VSS.n3921 0.00658571
R79382 VSS.n3924 VSS.n3922 0.00658571
R79383 VSS.n3924 VSS.n3923 0.00658571
R79384 VSS.n3923 VSS.n3911 0.00658571
R79385 VSS.n3931 VSS.n3911 0.00658571
R79386 VSS.n3932 VSS.n3931 0.00658571
R79387 VSS.n6210 VSS.n3932 0.00658571
R79388 VSS.n6210 VSS.n6209 0.00658571
R79389 VSS.n6209 VSS.n6208 0.00658571
R79390 VSS.n6208 VSS.n3933 0.00658571
R79391 VSS.n6202 VSS.n3933 0.00658571
R79392 VSS.n6202 VSS.n6201 0.00658571
R79393 VSS.n6201 VSS.n6200 0.00658571
R79394 VSS.n6200 VSS.n3937 0.00658571
R79395 VSS.n3963 VSS.n3937 0.00658571
R79396 VSS.n3964 VSS.n3963 0.00658571
R79397 VSS.n6190 VSS.n3964 0.00658571
R79398 VSS.n6190 VSS.n6189 0.00658571
R79399 VSS.n6189 VSS.n6188 0.00658571
R79400 VSS.n6188 VSS.n3965 0.00658571
R79401 VSS.n6182 VSS.n3965 0.00658571
R79402 VSS.n6182 VSS.n6181 0.00658571
R79403 VSS.n6181 VSS.n6180 0.00658571
R79404 VSS.n6180 VSS.n3969 0.00658571
R79405 VSS.n6174 VSS.n3969 0.00658571
R79406 VSS.n6174 VSS.n6173 0.00658571
R79407 VSS.n6173 VSS.n6172 0.00658571
R79408 VSS.n6172 VSS.n3973 0.00658571
R79409 VSS.n6166 VSS.n3973 0.00658571
R79410 VSS.n6166 VSS.n6165 0.00658571
R79411 VSS.n6165 VSS.n6164 0.00658571
R79412 VSS.n6164 VSS.n3977 0.00658571
R79413 VSS.n6154 VSS.n3977 0.00658571
R79414 VSS.n6154 VSS.n6153 0.00658571
R79415 VSS.n6153 VSS.n6152 0.00658571
R79416 VSS.n6152 VSS.n3999 0.00658571
R79417 VSS.n6146 VSS.n3999 0.00658571
R79418 VSS.n6146 VSS.n6145 0.00658571
R79419 VSS.n6145 VSS.n6144 0.00658571
R79420 VSS.n6144 VSS.n4003 0.00658571
R79421 VSS.n6138 VSS.n4003 0.00658571
R79422 VSS.n6138 VSS.n6137 0.00658571
R79423 VSS.n6137 VSS.n6136 0.00658571
R79424 VSS.n6136 VSS.n4007 0.00658571
R79425 VSS.n6130 VSS.n4007 0.00658571
R79426 VSS.n6130 VSS.n6129 0.00658571
R79427 VSS.n6129 VSS.n6128 0.00658571
R79428 VSS.n6128 VSS.n4011 0.00658571
R79429 VSS.n4179 VSS.n4011 0.00658571
R79430 VSS.n4184 VSS.n4179 0.00658571
R79431 VSS.n4185 VSS.n4184 0.00658571
R79432 VSS.n4219 VSS.n4185 0.00658571
R79433 VSS.n4219 VSS.n4218 0.00658571
R79434 VSS.n4218 VSS.n4217 0.00658571
R79435 VSS.n4217 VSS.n4186 0.00658571
R79436 VSS.n4211 VSS.n4186 0.00658571
R79437 VSS.n4211 VSS.n4210 0.00658571
R79438 VSS.n4210 VSS.n4209 0.00658571
R79439 VSS.n4209 VSS.n4190 0.00658571
R79440 VSS.n4203 VSS.n4190 0.00658571
R79441 VSS.n4203 VSS.n4202 0.00658571
R79442 VSS.n4202 VSS.n4201 0.00658571
R79443 VSS.n4201 VSS.n4194 0.00658571
R79444 VSS.n4195 VSS.n4194 0.00658571
R79445 VSS.n4195 VSS.n331 0.00658571
R79446 VSS.n9675 VSS.n331 0.00658571
R79447 VSS.n9675 VSS.n9674 0.00658571
R79448 VSS.n9674 VSS.n9673 0.00658571
R79449 VSS.n9673 VSS.n332 0.00658571
R79450 VSS.n9667 VSS.n332 0.00658571
R79451 VSS.n9667 VSS.n9666 0.00658571
R79452 VSS.n9666 VSS.n9665 0.00658571
R79453 VSS.n9665 VSS.n336 0.00658571
R79454 VSS.n9659 VSS.n336 0.00658571
R79455 VSS.n9659 VSS.n9658 0.00658571
R79456 VSS.n9658 VSS.n9657 0.00658571
R79457 VSS.n9657 VSS.n340 0.00658571
R79458 VSS.n9651 VSS.n340 0.00658571
R79459 VSS.n9651 VSS.n9650 0.00658571
R79460 VSS.n9650 VSS.n9649 0.00658571
R79461 VSS.n9649 VSS.n344 0.00658571
R79462 VSS.n372 VSS.n344 0.00658571
R79463 VSS.n373 VSS.n372 0.00658571
R79464 VSS.n9641 VSS.n373 0.00658571
R79465 VSS.n9641 VSS.n9640 0.00658571
R79466 VSS.n9640 VSS.n9639 0.00658571
R79467 VSS.n9639 VSS.n374 0.00658571
R79468 VSS.n9633 VSS.n374 0.00658571
R79469 VSS.n9633 VSS.n9632 0.00658571
R79470 VSS.n9632 VSS.n9631 0.00658571
R79471 VSS.n9631 VSS.n378 0.00658571
R79472 VSS.n9621 VSS.n378 0.00658571
R79473 VSS.n9621 VSS.n9620 0.00658571
R79474 VSS.n9620 VSS.n9619 0.00658571
R79475 VSS.n9619 VSS.n400 0.00658571
R79476 VSS.n9613 VSS.n400 0.00658571
R79477 VSS.n9612 VSS.n9611 0.00658571
R79478 VSS.n6234 VSS.n6233 0.00658571
R79479 VSS.n6233 VSS.n6232 0.00658571
R79480 VSS.n6232 VSS.n3876 0.00658571
R79481 VSS.n6226 VSS.n3876 0.00658571
R79482 VSS.n6226 VSS.n6225 0.00658571
R79483 VSS.n6225 VSS.n6224 0.00658571
R79484 VSS.n6224 VSS.n3880 0.00658571
R79485 VSS.n5277 VSS.n3880 0.00658571
R79486 VSS.n5281 VSS.n5277 0.00658571
R79487 VSS.n5282 VSS.n5281 0.00658571
R79488 VSS.n5283 VSS.n5282 0.00658571
R79489 VSS.n5283 VSS.n5273 0.00658571
R79490 VSS.n5289 VSS.n5273 0.00658571
R79491 VSS.n5290 VSS.n5289 0.00658571
R79492 VSS.n5291 VSS.n5290 0.00658571
R79493 VSS.n5291 VSS.n4311 0.00658571
R79494 VSS.n5306 VSS.n4311 0.00658571
R79495 VSS.n5307 VSS.n5306 0.00658571
R79496 VSS.n5308 VSS.n5307 0.00658571
R79497 VSS.n5308 VSS.n4307 0.00658571
R79498 VSS.n5314 VSS.n4307 0.00658571
R79499 VSS.n5315 VSS.n5314 0.00658571
R79500 VSS.n5316 VSS.n5315 0.00658571
R79501 VSS.n5316 VSS.n4303 0.00658571
R79502 VSS.n5322 VSS.n4303 0.00658571
R79503 VSS.n5323 VSS.n5322 0.00658571
R79504 VSS.n5324 VSS.n5323 0.00658571
R79505 VSS.n5324 VSS.n4299 0.00658571
R79506 VSS.n5330 VSS.n4299 0.00658571
R79507 VSS.n5331 VSS.n5330 0.00658571
R79508 VSS.n5628 VSS.n5331 0.00658571
R79509 VSS.n5628 VSS.n5627 0.00658571
R79510 VSS.n5627 VSS.n5626 0.00658571
R79511 VSS.n5626 VSS.n5332 0.00658571
R79512 VSS.n5336 VSS.n5332 0.00658571
R79513 VSS.n5618 VSS.n5336 0.00658571
R79514 VSS.n5618 VSS.n5617 0.00658571
R79515 VSS.n5617 VSS.n5616 0.00658571
R79516 VSS.n5616 VSS.n5337 0.00658571
R79517 VSS.n5610 VSS.n5337 0.00658571
R79518 VSS.n5610 VSS.n5609 0.00658571
R79519 VSS.n5609 VSS.n5608 0.00658571
R79520 VSS.n5608 VSS.n5341 0.00658571
R79521 VSS.n5602 VSS.n5341 0.00658571
R79522 VSS.n5602 VSS.n5601 0.00658571
R79523 VSS.n5601 VSS.n5600 0.00658571
R79524 VSS.n5600 VSS.n5345 0.00658571
R79525 VSS.n5595 VSS.n5345 0.00658571
R79526 VSS.n5595 VSS.n5594 0.00658571
R79527 VSS.n5594 VSS.n5593 0.00658571
R79528 VSS.n5593 VSS.n5348 0.00658571
R79529 VSS.n5588 VSS.n5348 0.00658571
R79530 VSS.n5588 VSS.n5587 0.00658571
R79531 VSS.n5587 VSS.n5586 0.00658571
R79532 VSS.n5586 VSS.n5350 0.00658571
R79533 VSS.n5580 VSS.n5350 0.00658571
R79534 VSS.n5580 VSS.n5579 0.00658571
R79535 VSS.n5579 VSS.n5578 0.00658571
R79536 VSS.n5578 VSS.n5355 0.00658571
R79537 VSS.n5572 VSS.n5355 0.00658571
R79538 VSS.n5572 VSS.n5571 0.00658571
R79539 VSS.n5571 VSS.n5570 0.00658571
R79540 VSS.n5570 VSS.n5359 0.00658571
R79541 VSS.n5564 VSS.n5359 0.00658571
R79542 VSS.n5564 VSS.n5563 0.00658571
R79543 VSS.n5563 VSS.n5562 0.00658571
R79544 VSS.n5562 VSS.n5362 0.00658571
R79545 VSS.n5556 VSS.n5362 0.00658571
R79546 VSS.n5556 VSS.n5555 0.00658571
R79547 VSS.n5555 VSS.n5554 0.00658571
R79548 VSS.n5554 VSS.n5364 0.00658571
R79549 VSS.n5548 VSS.n5364 0.00658571
R79550 VSS.n5548 VSS.n5547 0.00658571
R79551 VSS.n5547 VSS.n5546 0.00658571
R79552 VSS.n5546 VSS.n5369 0.00658571
R79553 VSS.n5540 VSS.n5369 0.00658571
R79554 VSS.n5540 VSS.n5539 0.00658571
R79555 VSS.n5539 VSS.n5538 0.00658571
R79556 VSS.n5538 VSS.n5373 0.00658571
R79557 VSS.n5532 VSS.n5373 0.00658571
R79558 VSS.n5532 VSS.n5531 0.00658571
R79559 VSS.n5531 VSS.n5530 0.00658571
R79560 VSS.n5530 VSS.n5377 0.00658571
R79561 VSS.n5399 VSS.n5377 0.00658571
R79562 VSS.n5519 VSS.n5399 0.00658571
R79563 VSS.n5519 VSS.n5518 0.00658571
R79564 VSS.n5518 VSS.n5517 0.00658571
R79565 VSS.n5517 VSS.n5400 0.00658571
R79566 VSS.n5511 VSS.n5400 0.00658571
R79567 VSS.n5511 VSS.n5510 0.00658571
R79568 VSS.n5510 VSS.n5509 0.00658571
R79569 VSS.n5509 VSS.n5404 0.00658571
R79570 VSS.n5498 VSS.n5404 0.00658571
R79571 VSS.n5498 VSS.n5497 0.00658571
R79572 VSS.n5497 VSS.n5496 0.00658571
R79573 VSS.n5496 VSS.n5424 0.00658571
R79574 VSS.n5490 VSS.n5424 0.00658571
R79575 VSS.n5489 VSS.n5488 0.00658571
R79576 VSS.n7874 VSS.n7873 0.00658571
R79577 VSS.n7873 VSS.n7872 0.00658571
R79578 VSS.n7872 VSS.n7275 0.00658571
R79579 VSS.n7866 VSS.n7275 0.00658571
R79580 VSS.n7866 VSS.n7865 0.00658571
R79581 VSS.n7865 VSS.n7864 0.00658571
R79582 VSS.n7864 VSS.n7280 0.00658571
R79583 VSS.n7858 VSS.n7280 0.00658571
R79584 VSS.n7858 VSS.n7857 0.00658571
R79585 VSS.n7857 VSS.n7856 0.00658571
R79586 VSS.n7856 VSS.n7284 0.00658571
R79587 VSS.n7850 VSS.n7284 0.00658571
R79588 VSS.n7850 VSS.n7849 0.00658571
R79589 VSS.n7849 VSS.n7848 0.00658571
R79590 VSS.n7848 VSS.n7601 0.00658571
R79591 VSS.n7842 VSS.n7601 0.00658571
R79592 VSS.n7842 VSS.n7841 0.00658571
R79593 VSS.n7841 VSS.n7840 0.00658571
R79594 VSS.n7840 VSS.n7605 0.00658571
R79595 VSS.n7834 VSS.n7605 0.00658571
R79596 VSS.n7834 VSS.n7833 0.00658571
R79597 VSS.n7833 VSS.n7832 0.00658571
R79598 VSS.n7832 VSS.n7609 0.00658571
R79599 VSS.n7826 VSS.n7609 0.00658571
R79600 VSS.n7826 VSS.n7825 0.00658571
R79601 VSS.n7825 VSS.n7824 0.00658571
R79602 VSS.n7824 VSS.n7613 0.00658571
R79603 VSS.n7818 VSS.n7613 0.00658571
R79604 VSS.n7818 VSS.n7817 0.00658571
R79605 VSS.n7817 VSS.n7816 0.00658571
R79606 VSS.n7816 VSS.n7617 0.00658571
R79607 VSS.n7810 VSS.n7617 0.00658571
R79608 VSS.n7810 VSS.n7809 0.00658571
R79609 VSS.n7809 VSS.n7808 0.00658571
R79610 VSS.n7808 VSS.n7621 0.00658571
R79611 VSS.n7802 VSS.n7621 0.00658571
R79612 VSS.n7802 VSS.n7801 0.00658571
R79613 VSS.n7801 VSS.n7800 0.00658571
R79614 VSS.n7800 VSS.n7625 0.00658571
R79615 VSS.n7794 VSS.n7625 0.00658571
R79616 VSS.n7794 VSS.n7793 0.00658571
R79617 VSS.n7793 VSS.n7792 0.00658571
R79618 VSS.n7792 VSS.n7629 0.00658571
R79619 VSS.n7786 VSS.n7629 0.00658571
R79620 VSS.n7786 VSS.n7785 0.00658571
R79621 VSS.n7785 VSS.n7784 0.00658571
R79622 VSS.n7784 VSS.n7633 0.00658571
R79623 VSS.n7778 VSS.n7633 0.00658571
R79624 VSS.n7778 VSS.n7777 0.00658571
R79625 VSS.n7777 VSS.n7776 0.00658571
R79626 VSS.n7776 VSS.n7637 0.00658571
R79627 VSS.n7770 VSS.n7637 0.00658571
R79628 VSS.n7770 VSS.n7769 0.00658571
R79629 VSS.n7769 VSS.n7768 0.00658571
R79630 VSS.n7768 VSS.n7641 0.00658571
R79631 VSS.n7762 VSS.n7641 0.00658571
R79632 VSS.n7762 VSS.n7761 0.00658571
R79633 VSS.n7761 VSS.n7760 0.00658571
R79634 VSS.n7760 VSS.n7645 0.00658571
R79635 VSS.n7754 VSS.n7645 0.00658571
R79636 VSS.n7754 VSS.n7753 0.00658571
R79637 VSS.n7753 VSS.n7752 0.00658571
R79638 VSS.n7752 VSS.n7649 0.00658571
R79639 VSS.n7746 VSS.n7649 0.00658571
R79640 VSS.n7746 VSS.n7745 0.00658571
R79641 VSS.n7745 VSS.n7744 0.00658571
R79642 VSS.n7744 VSS.n7653 0.00658571
R79643 VSS.n7738 VSS.n7653 0.00658571
R79644 VSS.n7738 VSS.n7737 0.00658571
R79645 VSS.n7737 VSS.n7736 0.00658571
R79646 VSS.n7736 VSS.n7657 0.00658571
R79647 VSS.n7730 VSS.n7657 0.00658571
R79648 VSS.n7730 VSS.n7729 0.00658571
R79649 VSS.n7729 VSS.n7728 0.00658571
R79650 VSS.n7728 VSS.n7661 0.00658571
R79651 VSS.n7722 VSS.n7661 0.00658571
R79652 VSS.n7722 VSS.n7721 0.00658571
R79653 VSS.n7721 VSS.n7720 0.00658571
R79654 VSS.n7720 VSS.n7665 0.00658571
R79655 VSS.n7714 VSS.n7665 0.00658571
R79656 VSS.n7714 VSS.n7713 0.00658571
R79657 VSS.n7713 VSS.n7712 0.00658571
R79658 VSS.n7712 VSS.n7669 0.00658571
R79659 VSS.n7706 VSS.n7669 0.00658571
R79660 VSS.n7706 VSS.n7705 0.00658571
R79661 VSS.n7705 VSS.n7704 0.00658571
R79662 VSS.n7704 VSS.n7673 0.00658571
R79663 VSS.n7698 VSS.n7673 0.00658571
R79664 VSS.n7698 VSS.n7697 0.00658571
R79665 VSS.n7697 VSS.n7696 0.00658571
R79666 VSS.n7696 VSS.n7677 0.00658571
R79667 VSS.n7690 VSS.n7677 0.00658571
R79668 VSS.n7690 VSS.n7689 0.00658571
R79669 VSS.n7689 VSS.n7688 0.00658571
R79670 VSS.n7688 VSS.n7681 0.00658571
R79671 VSS.n7682 VSS.n7681 0.00658571
R79672 VSS.n9912 VSS.n9911 0.00658571
R79673 VSS.n9172 VSS.n942 0.0065
R79674 VSS.n1433 VSS.n1008 0.0065
R79675 VSS.n7943 VSS.n1881 0.0065
R79676 VSS.n945 VSS.n940 0.0065
R79677 VSS.n8959 VSS.n721 0.0065
R79678 VSS.n1518 VSS.n945 0.0065
R79679 VSS.n7943 VSS.n2129 0.0065
R79680 VSS.n9064 VSS.n1011 0.0065
R79681 VSS.n9064 VSS.n861 0.0065
R79682 VSS.n721 VSS.n716 0.0065
R79683 VSS.n8236 VSS.n1879 0.0065
R79684 VSS.n9173 VSS.n9172 0.0065
R79685 VSS.n1008 VSS.n860 0.0065
R79686 VSS.n1139 VSS.n723 0.0065
R79687 VSS.n723 VSS.n715 0.0065
R79688 VSS.n7951 VSS.n1879 0.0065
R79689 VSS.n4712 VSS.n4588 0.00648592
R79690 VSS.n4697 VSS.n4631 0.00648592
R79691 VSS.n5225 VSS.n4339 0.00648592
R79692 VSS.n5198 VSS.n4394 0.00648592
R79693 VSS.n8294 VSS.n8287 0.00647857
R79694 VSS.n8323 VSS.n8316 0.00647857
R79695 VSS.n1578 VSS.n1568 0.00647857
R79696 VSS.n8410 VSS.n8378 0.00647857
R79697 VSS.n2805 VSS.n2797 0.00647857
R79698 VSS.n2830 VSS.n2829 0.00647857
R79699 VSS.n2856 VSS.n2855 0.00647857
R79700 VSS.n2890 VSS.n2889 0.00647857
R79701 VSS.n3842 VSS.n3833 0.00647857
R79702 VSS.n3956 VSS.n3944 0.00647857
R79703 VSS.n3980 VSS.n3979 0.00647857
R79704 VSS.n6238 VSS.n3866 0.00647857
R79705 VSS.n5296 VSS.n5293 0.00647857
R79706 VSS.n5630 VSS.n4289 0.00647857
R79707 VSS.n4737 VSS.n4729 0.00647857
R79708 VSS.n4779 VSS.n4563 0.00647857
R79709 VSS.n4337 VSS.n4330 0.00647857
R79710 VSS.n5060 VSS.n4522 0.00647857
R79711 VSS.n8056 VSS.n1454 0.00641549
R79712 VSS.n8064 VSS.n1487 0.00641549
R79713 VSS.n7416 VSS 0.00641429
R79714 VSS.n9795 DVSS 0.00641429
R79715 DVSS VSS.n8890 0.00641429
R79716 VSS.n1378 VSS.n1368 0.00641429
R79717 DVSS VSS.n6679 0.00641429
R79718 VSS.n6805 VSS.n2948 0.00641429
R79719 DVSS VSS.n9612 0.00641429
R79720 VSS.n4182 VSS.n4171 0.00641429
R79721 DVSS VSS.n5489 0.00641429
R79722 VSS.n5669 VSS.n4253 0.00641429
R79723 VSS.n5020 VSS.n4854 0.00641429
R79724 VSS VSS.n9912 0.00641429
R79725 VSS.n2299 VSS.n2159 0.00634646
R79726 VSS.n1197 VSS.n747 0.00634646
R79727 VSS.n8842 VSS.n1325 0.00622143
R79728 VSS.n8496 VSS.n1324 0.00622143
R79729 VSS.n8859 VSS.n1306 0.00622143
R79730 VSS.n8861 VSS.n1294 0.00622143
R79731 VSS.n8909 VSS.n1261 0.00622143
R79732 VSS.n1276 VSS.n1260 0.00622143
R79733 VSS.n9569 VSS.n542 0.00622143
R79734 VSS.n8885 VSS.n541 0.00622143
R79735 VSS.n6751 VSS.n2975 0.00622143
R79736 VSS.n2996 VSS.n2974 0.00622143
R79737 VSS.n6718 VSS.n6717 0.00622143
R79738 VSS.n6715 VSS.n6714 0.00622143
R79739 VSS.n3092 VSS.n3088 0.00622143
R79740 VSS.n6697 VSS.n3105 0.00622143
R79741 VSS.n9582 VSS.n504 0.00622143
R79742 VSS.n6674 VSS.n503 0.00622143
R79743 VSS.n9680 VSS.n311 0.00622143
R79744 VSS.n329 VSS.n310 0.00622143
R79745 VSS.n9647 VSS.n9646 0.00622143
R79746 VSS.n363 VSS.n358 0.00622143
R79747 VSS.n9635 VSS.n376 0.00622143
R79748 VSS.n9628 VSS.n387 0.00622143
R79749 VSS.n9615 VSS.n402 0.00622143
R79750 VSS.n9608 VSS.n413 0.00622143
R79751 VSS.n9683 VSS.n290 0.00622143
R79752 VSS.n5557 VSS.n289 0.00622143
R79753 VSS.n5379 VSS.n5375 0.00622143
R79754 VSS.n5525 VSS.n5392 0.00622143
R79755 VSS.n5513 VSS.n5402 0.00622143
R79756 VSS.n5506 VSS.n5413 0.00622143
R79757 VSS.n5492 VSS.n5426 0.00622143
R79758 VSS.n5485 VSS.n5437 0.00622143
R79759 VSS.n9694 VSS.n259 0.00622143
R79760 VSS.n9697 VSS.n250 0.00622143
R79761 VSS.n9758 VSS.n229 0.00622143
R79762 VSS.n9741 VSS.n228 0.00622143
R79763 VSS.n9776 VSS.n206 0.00622143
R79764 VSS.n9779 VSS.n194 0.00622143
R79765 VSS.n9809 VSS.n180 0.00622143
R79766 VSS.n9791 VSS.n179 0.00622143
R79767 VSS.n3723 VSS.n3148 0.00620423
R79768 VSS.n6807 VSS.n6806 0.00620423
R79769 VSS.n3793 VSS.n3178 0.00620423
R79770 VSS.n6839 VSS.n6838 0.00620423
R79771 VSS.n7598 VSS.n7286 0.00609286
R79772 VSS.n7595 VSS.n7288 0.00609286
R79773 VSS.n2307 VSS.n2161 0.00599213
R79774 VSS.n2419 VSS.n1849 0.00599213
R79775 VSS.n1189 VSS.n749 0.00599213
R79776 VSS.n9383 VSS.n696 0.00599213
R79777 VSS.n8301 VSS.n1702 0.00596429
R79778 VSS.n8330 VSS.n1682 0.00596429
R79779 VSS.n1676 VSS.n1569 0.00596429
R79780 VSS.n8412 VSS.n1651 0.00596429
R79781 VSS.n6960 VSS.n6956 0.00596429
R79782 VSS.n6938 VSS.n6933 0.00596429
R79783 VSS.n6915 VSS.n6910 0.00596429
R79784 VSS.n6876 VSS.n6871 0.00596429
R79785 VSS.n3913 VSS.n3834 0.00596429
R79786 VSS.n6195 VSS.n6192 0.00596429
R79787 VSS.n6159 VSS.n6156 0.00596429
R79788 VSS.n6230 VSS.n3867 0.00596429
R79789 VSS.n5303 VSS.n4309 0.00596429
R79790 VSS.n5622 VSS.n4290 0.00596429
R79791 VSS.n4764 VSS.n4580 0.00596429
R79792 VSS.n4786 VSS.n4548 0.00596429
R79793 VSS.n4542 VSS.n4331 0.00596429
R79794 VSS.n5052 VSS.n4523 0.00596429
R79795 VSS.n9827 VSS.n9825 0.00591803
R79796 VSS.n4607 VSS.n4590 0.00591803
R79797 VSS.n5710 VSS.n4175 0.00578169
R79798 VSS.n3743 VSS.n3158 0.00578169
R79799 VSS.n2446 VSS.n995 0.00578169
R79800 VSS.n5711 VSS.n4019 0.00578169
R79801 VSS.n3753 VSS.n3188 0.00578169
R79802 VSS.n2428 VSS.n974 0.00578169
R79803 VSS.n4717 VSS.n4589 0.00578169
R79804 VSS.n4702 VSS.n4677 0.00578169
R79805 VSS.n5230 VSS.n4340 0.00578169
R79806 VSS.n5203 VSS.n4397 0.00578169
R79807 VSS.n6215 VSS.n3895 0.00570714
R79808 VSS.n6222 VSS.n6221 0.00570714
R79809 VSS.n2315 VSS.n2146 0.0056378
R79810 VSS.n2411 VSS.n1854 0.0056378
R79811 VSS.n1181 VSS.n733 0.0056378
R79812 VSS.n9391 VSS.n700 0.0056378
R79813 VSS.n6213 VSS.n6212 0.00557857
R79814 VSS.n6218 VSS.n3893 0.00557857
R79815 VSS.n9889 VSS.n41 0.0055
R79816 VSS.n9889 VSS.n9888 0.0055
R79817 VSS.n9862 VSS.n74 0.0055
R79818 VSS.n9862 VSS.n9861 0.0055
R79819 VSS.n9847 VSS.n105 0.0055
R79820 VSS.n9847 VSS.n9846 0.0055
R79821 VSS.n9832 VSS.n136 0.0055
R79822 VSS.n9832 VSS.n9829 0.0055
R79823 VSS.n7414 VSS.n7413 0.00548841
R79824 VSS.n7301 VSS.n7300 0.00548841
R79825 VSS.n9793 VSS.n9792 0.00548841
R79826 VSS.n4736 VSS.n4731 0.00548841
R79827 VSS.n8886 VSS.n8884 0.00548841
R79828 VSS.n8286 VSS.n8281 0.00548841
R79829 VSS.n6675 VSS.n6673 0.00548841
R79830 VSS.n2818 VSS.n2799 0.00548841
R79831 VSS.n405 VSS.n404 0.00548841
R79832 VSS.n3916 VSS.n3836 0.00548841
R79833 VSS.n5429 VSS.n5428 0.00548841
R79834 VSS.n6237 VSS.n3869 0.00548841
R79835 VSS.n4 VSS.n3 0.00548841
R79836 VSS.n7876 VSS.n7272 0.00548841
R79837 VSS.n8045 VSS.n8036 0.00546063
R79838 VSS.n8050 VSS.n1410 0.00546063
R79839 VSS.n8069 VSS.n1538 0.00546063
R79840 VSS.n8077 VSS.n8075 0.00546063
R79841 VSS.n7682 VSS 0.00538571
R79842 VSS.n4248 VSS.n4244 0.00535915
R79843 VSS.n3746 VSS.n3138 0.00535915
R79844 VSS.n5664 VSS.n4263 0.00535915
R79845 VSS.n3747 VSS.n3168 0.00535915
R79846 VSS.n8293 VSS.n1706 0.00532143
R79847 VSS.n8322 VSS.n1686 0.00532143
R79848 VSS.n8345 VSS.n1570 0.00532143
R79849 VSS.n8384 VSS.n1655 0.00532143
R79850 VSS.n2819 VSS.n2798 0.00532143
R79851 VSS.n6942 VSS.n6941 0.00532143
R79852 VSS.n6919 VSS.n6918 0.00532143
R79853 VSS.n6880 VSS.n6879 0.00532143
R79854 VSS.n3917 VSS.n3835 0.00532143
R79855 VSS.n3961 VSS.n3951 0.00532143
R79856 VSS.n6162 VSS.n6161 0.00532143
R79857 VSS.n6235 VSS.n3868 0.00532143
R79858 VSS.n5295 VSS.n4313 0.00532143
R79859 VSS.n4297 VSS.n4291 0.00532143
R79860 VSS.n4728 VSS.n4584 0.00532143
R79861 VSS.n4562 VSS.n4552 0.00532143
R79862 VSS.n4801 VSS.n4332 0.00532143
R79863 VSS.n4530 VSS.n4524 0.00532143
R79864 VSS.n2291 VSS.n2151 0.00528346
R79865 VSS.n2373 VSS.n1839 0.00528346
R79866 VSS.n1205 VSS.n738 0.00528346
R79867 VSS.n9429 VSS.n686 0.00528346
R79868 VSS.n4714 VSS.n4589 0.00521831
R79869 VSS.n4699 VSS.n4677 0.00521831
R79870 VSS.n5227 VSS.n4340 0.00521831
R79871 VSS.n5200 VSS.n4397 0.00521831
R79872 VSS.n1331 VSS.n1322 0.00506429
R79873 VSS.n8498 VSS.n1322 0.00506429
R79874 VSS.n1309 VSS.n1288 0.00506429
R79875 VSS.n8862 VSS.n1288 0.00506429
R79876 VSS.n1267 VSS.n1259 0.00506429
R79877 VSS.n8878 VSS.n1259 0.00506429
R79878 VSS.n562 VSS.n548 0.00506429
R79879 VSS.n8887 VSS.n562 0.00506429
R79880 VSS.n6749 VSS.n2981 0.00506429
R79881 VSS.n6749 VSS.n6748 0.00506429
R79882 VSS.n3075 VSS.n3063 0.00506429
R79883 VSS.n3076 VSS.n3075 0.00506429
R79884 VSS.n6700 VSS.n6699 0.00506429
R79885 VSS.n6699 VSS.n3098 0.00506429
R79886 VSS.n524 VSS.n510 0.00506429
R79887 VSS.n6676 VSS.n524 0.00506429
R79888 VSS.n9678 VSS.n317 0.00506429
R79889 VSS.n9678 VSS.n9677 0.00506429
R79890 VSS.n362 VSS.n351 0.00506429
R79891 VSS.n370 VSS.n362 0.00506429
R79892 VSS.n381 VSS.n380 0.00506429
R79893 VSS.n9629 VSS.n381 0.00506429
R79894 VSS.n407 VSS.n406 0.00506429
R79895 VSS.n9609 VSS.n407 0.00506429
R79896 VSS.n295 VSS.n287 0.00506429
R79897 VSS.n5559 VSS.n287 0.00506429
R79898 VSS.n5528 VSS.n5527 0.00506429
R79899 VSS.n5527 VSS.n5385 0.00506429
R79900 VSS.n5407 VSS.n5406 0.00506429
R79901 VSS.n5507 VSS.n5407 0.00506429
R79902 VSS.n5431 VSS.n5430 0.00506429
R79903 VSS.n5486 VSS.n5431 0.00506429
R79904 VSS.n269 VSS.n263 0.00506429
R79905 VSS.n269 VSS.n268 0.00506429
R79906 VSS.n9747 VSS.n226 0.00506429
R79907 VSS.n234 VSS.n226 0.00506429
R79908 VSS.n211 VSS.n204 0.00506429
R79909 VSS.n204 VSS.n203 0.00506429
R79910 VSS.n9797 VSS.n177 0.00506429
R79911 VSS.n186 VSS.n177 0.00506429
R79912 VSS.n8572 VSS.n1446 0.00493662
R79913 VSS.n1549 VSS.n1479 0.00493662
R79914 VSS.n8971 VSS.n8970 0.00492913
R79915 VSS.n7930 VSS.n7892 0.00492913
R79916 VSS.n2395 VSS.n1844 0.00492913
R79917 VSS.n2454 VSS.n1032 0.00492913
R79918 VSS.n2430 VSS.n1993 0.00492913
R79919 VSS.n8097 VSS.n8096 0.00492913
R79920 VSS.n6239 VSS.n3859 0.00492913
R79921 VSS.n5438 VSS.n174 0.00492913
R79922 VSS.n9498 VSS.n9458 0.00492913
R79923 VSS.n9407 VSS.n691 0.00492913
R79924 VSS.n8302 VSS.n1706 0.00480714
R79925 VSS.n8331 VSS.n1686 0.00480714
R79926 VSS.n8347 VSS.n1570 0.00480714
R79927 VSS.n8413 VSS.n1655 0.00480714
R79928 VSS.n2814 VSS.n2798 0.00480714
R79929 VSS.n6941 VSS.n2836 0.00480714
R79930 VSS.n6918 VSS.n2862 0.00480714
R79931 VSS.n6879 VSS.n2896 0.00480714
R79932 VSS.n3919 VSS.n3835 0.00480714
R79933 VSS.n3957 VSS.n3951 0.00480714
R79934 VSS.n6161 VSS.n3986 0.00480714
R79935 VSS.n3874 VSS.n3868 0.00480714
R79936 VSS.n5304 VSS.n4313 0.00480714
R79937 VSS.n5624 VSS.n4291 0.00480714
R79938 VSS.n4765 VSS.n4584 0.00480714
R79939 VSS.n4787 VSS.n4552 0.00480714
R79940 VSS.n4803 VSS.n4332 0.00480714
R79941 VSS.n5054 VSS.n4524 0.00480714
R79942 VSS.n6556 VSS.n3268 0.00476
R79943 VSS.n6556 VSS.n6555 0.00476
R79944 VSS.n6555 VSS.n6553 0.00476
R79945 VSS.n6553 VSS.n3272 0.00476
R79946 VSS.n6549 VSS.n3272 0.00476
R79947 VSS.n6549 VSS.n6548 0.00476
R79948 VSS.n6548 VSS.n6547 0.00476
R79949 VSS.n6547 VSS.n3278 0.00476
R79950 VSS.n3329 VSS.n3278 0.00476
R79951 VSS.n6541 VSS.n3329 0.00476
R79952 VSS.n6541 VSS.n6540 0.00476
R79953 VSS.n6540 VSS.n3334 0.00476
R79954 VSS.n6536 VSS.n3334 0.00476
R79955 VSS.n6536 VSS.n6535 0.00476
R79956 VSS.n6535 VSS.n6534 0.00476
R79957 VSS.n6534 VSS.n3340 0.00476
R79958 VSS.n3391 VSS.n3340 0.00476
R79959 VSS.n6528 VSS.n3391 0.00476
R79960 VSS.n6528 VSS.n6527 0.00476
R79961 VSS.n6527 VSS.n3396 0.00476
R79962 VSS.n6523 VSS.n3396 0.00476
R79963 VSS.n6523 VSS.n6522 0.00476
R79964 VSS.n6522 VSS.n6521 0.00476
R79965 VSS.n6521 VSS.n3402 0.00476
R79966 VSS.n6517 VSS.n3402 0.00476
R79967 VSS.n6517 VSS.n6516 0.00476
R79968 VSS.n6516 VSS.n6515 0.00476
R79969 VSS.n6515 VSS.n3408 0.00476
R79970 VSS.n6511 VSS.n3408 0.00476
R79971 VSS.n6511 VSS.n6510 0.00476
R79972 VSS.n6510 VSS.n6509 0.00476
R79973 VSS.n6509 VSS.n3414 0.00476
R79974 VSS.n3465 VSS.n3414 0.00476
R79975 VSS.n6503 VSS.n3465 0.00476
R79976 VSS.n6503 VSS.n6502 0.00476
R79977 VSS.n6502 VSS.n3470 0.00476
R79978 VSS.n6498 VSS.n3470 0.00476
R79979 VSS.n6498 VSS.n6497 0.00476
R79980 VSS.n6497 VSS.n6496 0.00476
R79981 VSS.n6496 VSS.n3476 0.00476
R79982 VSS.n6492 VSS.n3476 0.00476
R79983 VSS.n6492 VSS.n6491 0.00476
R79984 VSS.n6491 VSS.n6490 0.00476
R79985 VSS.n6490 VSS.n3482 0.00476
R79986 VSS.n6486 VSS.n3482 0.00476
R79987 VSS.n6486 VSS.n6485 0.00476
R79988 VSS.n6485 VSS.n6484 0.00476
R79989 VSS.n6484 VSS.n6483 0.00476
R79990 VSS.n6483 VSS.n6482 0.00476
R79991 VSS.n6482 VSS.n6479 0.00476
R79992 VSS.n6479 VSS.n6477 0.00476
R79993 VSS.n6477 VSS.n6476 0.00476
R79994 VSS.n6476 VSS.n6475 0.00476
R79995 VSS.n6475 VSS.n6473 0.00476
R79996 VSS.n6473 VSS.n3495 0.00476
R79997 VSS.n6469 VSS.n3495 0.00476
R79998 VSS.n6469 VSS.n6468 0.00476
R79999 VSS.n6468 VSS.n6467 0.00476
R80000 VSS.n6467 VSS.n3501 0.00476
R80001 VSS.n6463 VSS.n3501 0.00476
R80002 VSS.n6463 VSS.n6462 0.00476
R80003 VSS.n6462 VSS.n6461 0.00476
R80004 VSS.n6461 VSS.n3507 0.00476
R80005 VSS.n6457 VSS.n3507 0.00476
R80006 VSS.n6457 VSS.n6456 0.00476
R80007 VSS.n6456 VSS.n6455 0.00476
R80008 VSS.n6455 VSS.n3513 0.00476
R80009 VSS.n3564 VSS.n3513 0.00476
R80010 VSS.n6449 VSS.n3564 0.00476
R80011 VSS.n6449 VSS.n6448 0.00476
R80012 VSS.n6448 VSS.n3569 0.00476
R80013 VSS.n6444 VSS.n3569 0.00476
R80014 VSS.n6444 VSS.n6443 0.00476
R80015 VSS.n6443 VSS.n6442 0.00476
R80016 VSS.n6442 VSS.n3575 0.00476
R80017 VSS.n6438 VSS.n3575 0.00476
R80018 VSS.n6438 VSS.n6437 0.00476
R80019 VSS.n6437 VSS.n6436 0.00476
R80020 VSS.n6436 VSS.n3581 0.00476
R80021 VSS.n6432 VSS.n3581 0.00476
R80022 VSS.n6432 VSS.n6431 0.00476
R80023 VSS.n6431 VSS.n6430 0.00476
R80024 VSS.n6430 VSS.n3587 0.00476
R80025 VSS.n3630 VSS.n3587 0.00476
R80026 VSS.n3630 VSS.n3628 0.00476
R80027 VSS.n6412 VSS.n3628 0.00476
R80028 VSS.n6412 VSS.n6411 0.00476
R80029 VSS.n6411 VSS.n6410 0.00476
R80030 VSS.n6410 VSS.n3636 0.00476
R80031 VSS.n6406 VSS.n3636 0.00476
R80032 VSS.n6406 VSS.n6405 0.00476
R80033 VSS.n6405 VSS.n3641 0.00476
R80034 VSS.n6361 VSS.n3641 0.00476
R80035 VSS.n6394 VSS.n6361 0.00476
R80036 VSS.n6394 VSS.n6393 0.00476
R80037 VSS.n6393 VSS.n6392 0.00476
R80038 VSS.n6392 VSS.n6389 0.00476
R80039 VSS.n6388 VSS.n6387 0.00476
R80040 VSS.n6387 VSS.n6386 0.00476
R80041 VSS.n6386 VSS.n6373 0.00476
R80042 VSS.n2244 VSS.n2230 0.00476
R80043 VSS.n2246 VSS.n2244 0.00476
R80044 VSS.n2248 VSS.n2246 0.00476
R80045 VSS.n2248 VSS.n2228 0.00476
R80046 VSS.n2253 VSS.n2228 0.00476
R80047 VSS.n2253 VSS.n2225 0.00476
R80048 VSS.n2257 VSS.n2225 0.00476
R80049 VSS.n2259 VSS.n2257 0.00476
R80050 VSS.n2261 VSS.n2259 0.00476
R80051 VSS.n2261 VSS.n2223 0.00476
R80052 VSS.n2267 VSS.n2223 0.00476
R80053 VSS.n2267 VSS.n2266 0.00476
R80054 VSS.n2266 VSS.n2132 0.00476
R80055 VSS.n7949 VSS.n2132 0.00476
R80056 VSS.n7955 VSS.n7953 0.00476
R80057 VSS.n7957 VSS.n7955 0.00476
R80058 VSS.n7957 VSS.n2127 0.00476
R80059 VSS.n7998 VSS.n2127 0.00476
R80060 VSS.n7998 VSS.n7997 0.00476
R80061 VSS.n7997 VSS.n7996 0.00476
R80062 VSS.n7996 VSS.n7963 0.00476
R80063 VSS.n7992 VSS.n7963 0.00476
R80064 VSS.n7992 VSS.n7991 0.00476
R80065 VSS.n7991 VSS.n7990 0.00476
R80066 VSS.n7990 VSS.n7969 0.00476
R80067 VSS.n7986 VSS.n7969 0.00476
R80068 VSS.n7986 VSS.n7985 0.00476
R80069 VSS.n7985 VSS.n7984 0.00476
R80070 VSS.n7984 VSS.n7975 0.00476
R80071 VSS.n7980 VSS.n7975 0.00476
R80072 VSS.n7980 VSS.n7979 0.00476
R80073 VSS.n7979 VSS.n1522 0.00476
R80074 VSS.n8637 VSS.n1522 0.00476
R80075 VSS.n8637 VSS.n1520 0.00476
R80076 VSS.n8641 VSS.n1520 0.00476
R80077 VSS.n8641 VSS.n1517 0.00476
R80078 VSS.n8645 VSS.n1517 0.00476
R80079 VSS.n8650 VSS.n1515 0.00476
R80080 VSS.n8650 VSS.n1513 0.00476
R80081 VSS.n8654 VSS.n1513 0.00476
R80082 VSS.n8654 VSS.n1511 0.00476
R80083 VSS.n8658 VSS.n1511 0.00476
R80084 VSS.n8658 VSS.n1509 0.00476
R80085 VSS.n8662 VSS.n1509 0.00476
R80086 VSS.n8662 VSS.n1507 0.00476
R80087 VSS.n8666 VSS.n1507 0.00476
R80088 VSS.n8666 VSS.n1476 0.00476
R80089 VSS.n8688 VSS.n1476 0.00476
R80090 VSS.n8688 VSS.n1474 0.00476
R80091 VSS.n8692 VSS.n1474 0.00476
R80092 VSS.n8692 VSS.n1443 0.00476
R80093 VSS.n8714 VSS.n1443 0.00476
R80094 VSS.n8714 VSS.n1441 0.00476
R80095 VSS.n8718 VSS.n1441 0.00476
R80096 VSS.n8718 VSS.n1439 0.00476
R80097 VSS.n8722 VSS.n1439 0.00476
R80098 VSS.n8722 VSS.n1437 0.00476
R80099 VSS.n8726 VSS.n1437 0.00476
R80100 VSS.n8726 VSS.n1435 0.00476
R80101 VSS.n8730 VSS.n1435 0.00476
R80102 VSS.n8735 VSS.n1432 0.00476
R80103 VSS.n8739 VSS.n1432 0.00476
R80104 VSS.n8740 VSS.n8739 0.00476
R80105 VSS.n8740 VSS.n1430 0.00476
R80106 VSS.n8793 VSS.n1430 0.00476
R80107 VSS.n8793 VSS.n8792 0.00476
R80108 VSS.n8792 VSS.n8790 0.00476
R80109 VSS.n8790 VSS.n8746 0.00476
R80110 VSS.n8786 VSS.n8746 0.00476
R80111 VSS.n8786 VSS.n8785 0.00476
R80112 VSS.n8785 VSS.n8784 0.00476
R80113 VSS.n8784 VSS.n8752 0.00476
R80114 VSS.n8780 VSS.n8752 0.00476
R80115 VSS.n8780 VSS.n8779 0.00476
R80116 VSS.n8779 VSS.n8778 0.00476
R80117 VSS.n8778 VSS.n8758 0.00476
R80118 VSS.n8774 VSS.n8758 0.00476
R80119 VSS.n8774 VSS.n8773 0.00476
R80120 VSS.n8773 VSS.n8772 0.00476
R80121 VSS.n8772 VSS.n8770 0.00476
R80122 VSS.n8770 VSS.n8768 0.00476
R80123 VSS.n8768 VSS.n1140 0.00476
R80124 VSS.n8960 VSS.n1140 0.00476
R80125 VSS.n8958 VSS.n1143 0.00476
R80126 VSS.n8954 VSS.n1143 0.00476
R80127 VSS.n8954 VSS.n8953 0.00476
R80128 VSS.n8953 VSS.n8952 0.00476
R80129 VSS.n8952 VSS.n1149 0.00476
R80130 VSS.n8913 VSS.n1149 0.00476
R80131 VSS.n8946 VSS.n8913 0.00476
R80132 VSS.n8946 VSS.n8945 0.00476
R80133 VSS.n8945 VSS.n8944 0.00476
R80134 VSS.n8944 VSS.n8941 0.00476
R80135 VSS.n8940 VSS.n8939 0.00476
R80136 VSS.n8939 VSS.n8938 0.00476
R80137 VSS.n8938 VSS.n8925 0.00476
R80138 VSS.n7913 VSS.n7900 0.00476
R80139 VSS.n7915 VSS.n7913 0.00476
R80140 VSS.n7915 VSS.n7898 0.00476
R80141 VSS.n7919 VSS.n7898 0.00476
R80142 VSS.n7919 VSS.n7896 0.00476
R80143 VSS.n7923 VSS.n7896 0.00476
R80144 VSS.n7923 VSS.n7894 0.00476
R80145 VSS.n7927 VSS.n7894 0.00476
R80146 VSS.n7927 VSS.n2141 0.00476
R80147 VSS.n7933 VSS.n2141 0.00476
R80148 VSS.n7933 VSS.n2139 0.00476
R80149 VSS.n7938 VSS.n2139 0.00476
R80150 VSS.n7938 VSS.n2137 0.00476
R80151 VSS.n7942 VSS.n2137 0.00476
R80152 VSS.n7944 VSS.n2034 0.00476
R80153 VSS.n8105 VSS.n2034 0.00476
R80154 VSS.n8105 VSS.n2032 0.00476
R80155 VSS.n8109 VSS.n2032 0.00476
R80156 VSS.n8109 VSS.n2030 0.00476
R80157 VSS.n8113 VSS.n2030 0.00476
R80158 VSS.n8113 VSS.n2028 0.00476
R80159 VSS.n8117 VSS.n2028 0.00476
R80160 VSS.n8117 VSS.n2026 0.00476
R80161 VSS.n8121 VSS.n2026 0.00476
R80162 VSS.n8121 VSS.n2024 0.00476
R80163 VSS.n8125 VSS.n2024 0.00476
R80164 VSS.n8125 VSS.n2022 0.00476
R80165 VSS.n8130 VSS.n2022 0.00476
R80166 VSS.n8130 VSS.n2020 0.00476
R80167 VSS.n8134 VSS.n2020 0.00476
R80168 VSS.n8135 VSS.n8134 0.00476
R80169 VSS.n8137 VSS.n8135 0.00476
R80170 VSS.n8137 VSS.n2018 0.00476
R80171 VSS.n8148 VSS.n2018 0.00476
R80172 VSS.n8148 VSS.n8147 0.00476
R80173 VSS.n8147 VSS.n8146 0.00476
R80174 VSS.n8146 VSS.n8144 0.00476
R80175 VSS.n9170 VSS.n9169 0.00476
R80176 VSS.n9169 VSS.n9168 0.00476
R80177 VSS.n9168 VSS.n949 0.00476
R80178 VSS.n9164 VSS.n949 0.00476
R80179 VSS.n9164 VSS.n9163 0.00476
R80180 VSS.n9163 VSS.n9162 0.00476
R80181 VSS.n9162 VSS.n955 0.00476
R80182 VSS.n9158 VSS.n955 0.00476
R80183 VSS.n9158 VSS.n9157 0.00476
R80184 VSS.n9157 VSS.n960 0.00476
R80185 VSS.n9118 VSS.n960 0.00476
R80186 VSS.n9118 VSS.n9117 0.00476
R80187 VSS.n9117 VSS.n9116 0.00476
R80188 VSS.n9116 VSS.n980 0.00476
R80189 VSS.n9077 VSS.n980 0.00476
R80190 VSS.n9077 VSS.n9076 0.00476
R80191 VSS.n9076 VSS.n9075 0.00476
R80192 VSS.n9075 VSS.n1001 0.00476
R80193 VSS.n9071 VSS.n1001 0.00476
R80194 VSS.n9071 VSS.n9070 0.00476
R80195 VSS.n9070 VSS.n9069 0.00476
R80196 VSS.n9069 VSS.n1007 0.00476
R80197 VSS.n9065 VSS.n1007 0.00476
R80198 VSS.n9063 VSS.n1013 0.00476
R80199 VSS.n9059 VSS.n1013 0.00476
R80200 VSS.n9059 VSS.n9058 0.00476
R80201 VSS.n9058 VSS.n9057 0.00476
R80202 VSS.n9057 VSS.n1019 0.00476
R80203 VSS.n1056 VSS.n1019 0.00476
R80204 VSS.n9037 VSS.n1056 0.00476
R80205 VSS.n9037 VSS.n9036 0.00476
R80206 VSS.n9036 VSS.n9035 0.00476
R80207 VSS.n9035 VSS.n1062 0.00476
R80208 VSS.n9031 VSS.n1062 0.00476
R80209 VSS.n9031 VSS.n9030 0.00476
R80210 VSS.n9030 VSS.n9029 0.00476
R80211 VSS.n9029 VSS.n1068 0.00476
R80212 VSS.n9025 VSS.n1068 0.00476
R80213 VSS.n9025 VSS.n9024 0.00476
R80214 VSS.n9024 VSS.n9023 0.00476
R80215 VSS.n9023 VSS.n1074 0.00476
R80216 VSS.n9019 VSS.n1074 0.00476
R80217 VSS.n9019 VSS.n9018 0.00476
R80218 VSS.n9018 VSS.n1079 0.00476
R80219 VSS.n8998 VSS.n1079 0.00476
R80220 VSS.n8999 VSS.n8998 0.00476
R80221 VSS.n9507 VSS.n722 0.00476
R80222 VSS.n9503 VSS.n722 0.00476
R80223 VSS.n9503 VSS.n9502 0.00476
R80224 VSS.n9502 VSS.n9501 0.00476
R80225 VSS.n9501 VSS.n728 0.00476
R80226 VSS.n9495 VSS.n728 0.00476
R80227 VSS.n9495 VSS.n9494 0.00476
R80228 VSS.n9494 VSS.n9462 0.00476
R80229 VSS.n9490 VSS.n9462 0.00476
R80230 VSS.n9490 VSS.n9489 0.00476
R80231 VSS.n9489 VSS.n9488 0.00476
R80232 VSS.n9486 VSS.n9485 0.00476
R80233 VSS.n9485 VSS.n9472 0.00476
R80234 VSS.n8256 VSS.n1828 0.00476
R80235 VSS.n8256 VSS.n8255 0.00476
R80236 VSS.n8255 VSS.n8253 0.00476
R80237 VSS.n8253 VSS.n1832 0.00476
R80238 VSS.n8249 VSS.n1832 0.00476
R80239 VSS.n8249 VSS.n8248 0.00476
R80240 VSS.n8248 VSS.n8247 0.00476
R80241 VSS.n8247 VSS.n1838 0.00476
R80242 VSS.n1872 VSS.n1838 0.00476
R80243 VSS.n1872 VSS.n1869 0.00476
R80244 VSS.n8241 VSS.n1869 0.00476
R80245 VSS.n8241 VSS.n8240 0.00476
R80246 VSS.n8240 VSS.n8239 0.00476
R80247 VSS.n8239 VSS.n1878 0.00476
R80248 VSS.n8234 VSS.n8233 0.00476
R80249 VSS.n8233 VSS.n1884 0.00476
R80250 VSS.n1930 VSS.n1884 0.00476
R80251 VSS.n8222 VSS.n1930 0.00476
R80252 VSS.n8222 VSS.n8221 0.00476
R80253 VSS.n8221 VSS.n8220 0.00476
R80254 VSS.n8220 VSS.n1936 0.00476
R80255 VSS.n8216 VSS.n1936 0.00476
R80256 VSS.n8216 VSS.n8215 0.00476
R80257 VSS.n8215 VSS.n8214 0.00476
R80258 VSS.n8214 VSS.n1942 0.00476
R80259 VSS.n8210 VSS.n1942 0.00476
R80260 VSS.n8210 VSS.n8209 0.00476
R80261 VSS.n8209 VSS.n8208 0.00476
R80262 VSS.n8208 VSS.n1948 0.00476
R80263 VSS.n8204 VSS.n1948 0.00476
R80264 VSS.n8204 VSS.n8203 0.00476
R80265 VSS.n8203 VSS.n1953 0.00476
R80266 VSS.n8186 VSS.n1953 0.00476
R80267 VSS.n8192 VSS.n8186 0.00476
R80268 VSS.n8192 VSS.n8191 0.00476
R80269 VSS.n8191 VSS.n939 0.00476
R80270 VSS.n9175 VSS.n939 0.00476
R80271 VSS.n9180 VSS.n936 0.00476
R80272 VSS.n9180 VSS.n934 0.00476
R80273 VSS.n9184 VSS.n934 0.00476
R80274 VSS.n9184 VSS.n932 0.00476
R80275 VSS.n9188 VSS.n932 0.00476
R80276 VSS.n9188 VSS.n930 0.00476
R80277 VSS.n9192 VSS.n930 0.00476
R80278 VSS.n9192 VSS.n928 0.00476
R80279 VSS.n9196 VSS.n928 0.00476
R80280 VSS.n9196 VSS.n900 0.00476
R80281 VSS.n9225 VSS.n900 0.00476
R80282 VSS.n9225 VSS.n898 0.00476
R80283 VSS.n9229 VSS.n898 0.00476
R80284 VSS.n9229 VSS.n872 0.00476
R80285 VSS.n9258 VSS.n872 0.00476
R80286 VSS.n9258 VSS.n870 0.00476
R80287 VSS.n9262 VSS.n870 0.00476
R80288 VSS.n9262 VSS.n868 0.00476
R80289 VSS.n9266 VSS.n868 0.00476
R80290 VSS.n9266 VSS.n866 0.00476
R80291 VSS.n9270 VSS.n866 0.00476
R80292 VSS.n9270 VSS.n864 0.00476
R80293 VSS.n9274 VSS.n864 0.00476
R80294 VSS.n9278 VSS.n859 0.00476
R80295 VSS.n9282 VSS.n859 0.00476
R80296 VSS.n9282 VSS.n857 0.00476
R80297 VSS.n9286 VSS.n857 0.00476
R80298 VSS.n9286 VSS.n830 0.00476
R80299 VSS.n9316 VSS.n830 0.00476
R80300 VSS.n9316 VSS.n828 0.00476
R80301 VSS.n9320 VSS.n828 0.00476
R80302 VSS.n9320 VSS.n826 0.00476
R80303 VSS.n9324 VSS.n826 0.00476
R80304 VSS.n9324 VSS.n824 0.00476
R80305 VSS.n9328 VSS.n824 0.00476
R80306 VSS.n9328 VSS.n822 0.00476
R80307 VSS.n9332 VSS.n822 0.00476
R80308 VSS.n9332 VSS.n820 0.00476
R80309 VSS.n9337 VSS.n820 0.00476
R80310 VSS.n9337 VSS.n818 0.00476
R80311 VSS.n9341 VSS.n818 0.00476
R80312 VSS.n9342 VSS.n9341 0.00476
R80313 VSS.n9342 VSS.n816 0.00476
R80314 VSS.n9351 VSS.n816 0.00476
R80315 VSS.n9351 VSS.n9350 0.00476
R80316 VSS.n9350 VSS.n9348 0.00476
R80317 VSS.n9512 VSS.n714 0.00476
R80318 VSS.n9517 VSS.n714 0.00476
R80319 VSS.n9517 VSS.n712 0.00476
R80320 VSS.n9521 VSS.n712 0.00476
R80321 VSS.n9521 VSS.n684 0.00476
R80322 VSS.n9528 VSS.n684 0.00476
R80323 VSS.n9528 VSS.n682 0.00476
R80324 VSS.n9533 VSS.n682 0.00476
R80325 VSS.n9533 VSS.n679 0.00476
R80326 VSS.n9537 VSS.n679 0.00476
R80327 VSS.n9538 VSS.n678 0.00476
R80328 VSS.n9545 VSS.n678 0.00476
R80329 VSS.n9545 VSS.n9544 0.00476
R80330 VSS.n8252 VSS.n8251 0.00476
R80331 VSS.n8251 VSS.n8250 0.00476
R80332 VSS.n8250 VSS.n1833 0.00476
R80333 VSS.n8246 VSS.n1833 0.00476
R80334 VSS.n8242 VSS.n1868 0.00476
R80335 VSS.n8238 VSS.n1868 0.00476
R80336 VSS.n8238 VSS.n8237 0.00476
R80337 VSS.n8223 VSS.n1929 0.00476
R80338 VSS.n8219 VSS.n1929 0.00476
R80339 VSS.n8219 VSS.n8218 0.00476
R80340 VSS.n8218 VSS.n8217 0.00476
R80341 VSS.n8217 VSS.n1937 0.00476
R80342 VSS.n8213 VSS.n1937 0.00476
R80343 VSS.n8213 VSS.n8212 0.00476
R80344 VSS.n8212 VSS.n8211 0.00476
R80345 VSS.n8211 VSS.n1943 0.00476
R80346 VSS.n8207 VSS.n1943 0.00476
R80347 VSS.n8207 VSS.n8206 0.00476
R80348 VSS.n8206 VSS.n8205 0.00476
R80349 VSS.n8193 VSS.n8185 0.00476
R80350 VSS.n8185 VSS.n941 0.00476
R80351 VSS.n9174 VSS.n941 0.00476
R80352 VSS.n9181 VSS.n935 0.00476
R80353 VSS.n9182 VSS.n9181 0.00476
R80354 VSS.n9183 VSS.n9182 0.00476
R80355 VSS.n9183 VSS.n931 0.00476
R80356 VSS.n9189 VSS.n931 0.00476
R80357 VSS.n9190 VSS.n9189 0.00476
R80358 VSS.n9191 VSS.n9190 0.00476
R80359 VSS.n9191 VSS.n916 0.00476
R80360 VSS.n9224 VSS.n887 0.00476
R80361 VSS.n9257 VSS.n869 0.00476
R80362 VSS.n9263 VSS.n869 0.00476
R80363 VSS.n9264 VSS.n9263 0.00476
R80364 VSS.n9265 VSS.n9264 0.00476
R80365 VSS.n9265 VSS.n865 0.00476
R80366 VSS.n9271 VSS.n865 0.00476
R80367 VSS.n9272 VSS.n9271 0.00476
R80368 VSS.n9273 VSS.n9272 0.00476
R80369 VSS.n9280 VSS.n9279 0.00476
R80370 VSS.n9281 VSS.n9280 0.00476
R80371 VSS.n9281 VSS.n845 0.00476
R80372 VSS.n9321 VSS.n827 0.00476
R80373 VSS.n9322 VSS.n9321 0.00476
R80374 VSS.n9323 VSS.n9322 0.00476
R80375 VSS.n9323 VSS.n823 0.00476
R80376 VSS.n9329 VSS.n823 0.00476
R80377 VSS.n9330 VSS.n9329 0.00476
R80378 VSS.n9331 VSS.n9330 0.00476
R80379 VSS.n9331 VSS.n819 0.00476
R80380 VSS.n9338 VSS.n819 0.00476
R80381 VSS.n9339 VSS.n9338 0.00476
R80382 VSS.n9340 VSS.n9339 0.00476
R80383 VSS.n9340 VSS.n782 0.00476
R80384 VSS.n9514 VSS.n9513 0.00476
R80385 VSS.n9516 VSS.n9514 0.00476
R80386 VSS.n9516 VSS.n9515 0.00476
R80387 VSS.n9534 VSS.n681 0.00476
R80388 VSS.n9535 VSS.n9534 0.00476
R80389 VSS.n9536 VSS.n9535 0.00476
R80390 VSS.n7920 VSS.n7897 0.00476
R80391 VSS.n7921 VSS.n7920 0.00476
R80392 VSS.n7922 VSS.n7921 0.00476
R80393 VSS.n7922 VSS.n7893 0.00476
R80394 VSS.n7939 VSS.n2138 0.00476
R80395 VSS.n7940 VSS.n7939 0.00476
R80396 VSS.n7941 VSS.n7940 0.00476
R80397 VSS.n8111 VSS.n8110 0.00476
R80398 VSS.n8112 VSS.n8111 0.00476
R80399 VSS.n8112 VSS.n2027 0.00476
R80400 VSS.n8118 VSS.n2027 0.00476
R80401 VSS.n8119 VSS.n8118 0.00476
R80402 VSS.n8120 VSS.n8119 0.00476
R80403 VSS.n8120 VSS.n2023 0.00476
R80404 VSS.n8126 VSS.n2023 0.00476
R80405 VSS.n8127 VSS.n8126 0.00476
R80406 VSS.n8129 VSS.n8127 0.00476
R80407 VSS.n8129 VSS.n8128 0.00476
R80408 VSS.n8128 VSS.n1981 0.00476
R80409 VSS.n8149 VSS.n2017 0.00476
R80410 VSS.n8145 VSS.n2017 0.00476
R80411 VSS.n8145 VSS.n943 0.00476
R80412 VSS.n9171 VSS.n944 0.00476
R80413 VSS.n9167 VSS.n944 0.00476
R80414 VSS.n9167 VSS.n9166 0.00476
R80415 VSS.n9166 VSS.n9165 0.00476
R80416 VSS.n9165 VSS.n950 0.00476
R80417 VSS.n9161 VSS.n950 0.00476
R80418 VSS.n9161 VSS.n9160 0.00476
R80419 VSS.n9160 VSS.n9159 0.00476
R80420 VSS.n9119 VSS.n975 0.00476
R80421 VSS.n9078 VSS.n996 0.00476
R80422 VSS.n9074 VSS.n996 0.00476
R80423 VSS.n9074 VSS.n9073 0.00476
R80424 VSS.n9073 VSS.n9072 0.00476
R80425 VSS.n9072 VSS.n1002 0.00476
R80426 VSS.n9068 VSS.n1002 0.00476
R80427 VSS.n9068 VSS.n9067 0.00476
R80428 VSS.n9067 VSS.n9066 0.00476
R80429 VSS.n9062 VSS.n9061 0.00476
R80430 VSS.n9061 VSS.n9060 0.00476
R80431 VSS.n9060 VSS.n1014 0.00476
R80432 VSS.n9038 VSS.n1055 0.00476
R80433 VSS.n9034 VSS.n1055 0.00476
R80434 VSS.n9034 VSS.n9033 0.00476
R80435 VSS.n9033 VSS.n9032 0.00476
R80436 VSS.n9032 VSS.n1063 0.00476
R80437 VSS.n9028 VSS.n1063 0.00476
R80438 VSS.n9028 VSS.n9027 0.00476
R80439 VSS.n9027 VSS.n9026 0.00476
R80440 VSS.n9026 VSS.n1069 0.00476
R80441 VSS.n9022 VSS.n1069 0.00476
R80442 VSS.n9022 VSS.n9021 0.00476
R80443 VSS.n9021 VSS.n9020 0.00476
R80444 VSS.n9506 VSS.n9505 0.00476
R80445 VSS.n9505 VSS.n9504 0.00476
R80446 VSS.n9504 VSS.n724 0.00476
R80447 VSS.n9493 VSS.n9492 0.00476
R80448 VSS.n9492 VSS.n9491 0.00476
R80449 VSS.n9491 VSS.n9463 0.00476
R80450 VSS.n9487 VSS.n9463 0.00476
R80451 VSS.n2247 VSS.n2227 0.00476
R80452 VSS.n2254 VSS.n2227 0.00476
R80453 VSS.n2255 VSS.n2254 0.00476
R80454 VSS.n2256 VSS.n2255 0.00476
R80455 VSS.n2268 VSS.n2222 0.00476
R80456 VSS.n2222 VSS.n2131 0.00476
R80457 VSS.n7950 VSS.n2131 0.00476
R80458 VSS.n7999 VSS.n2126 0.00476
R80459 VSS.n7995 VSS.n2126 0.00476
R80460 VSS.n7995 VSS.n7994 0.00476
R80461 VSS.n7994 VSS.n7993 0.00476
R80462 VSS.n7993 VSS.n7964 0.00476
R80463 VSS.n7989 VSS.n7964 0.00476
R80464 VSS.n7989 VSS.n7988 0.00476
R80465 VSS.n7988 VSS.n7987 0.00476
R80466 VSS.n7987 VSS.n7970 0.00476
R80467 VSS.n7983 VSS.n7970 0.00476
R80468 VSS.n7983 VSS.n7982 0.00476
R80469 VSS.n7982 VSS.n7981 0.00476
R80470 VSS.n8642 VSS.n1519 0.00476
R80471 VSS.n8643 VSS.n8642 0.00476
R80472 VSS.n8644 VSS.n8643 0.00476
R80473 VSS.n8651 VSS.n1514 0.00476
R80474 VSS.n8652 VSS.n8651 0.00476
R80475 VSS.n8653 VSS.n8652 0.00476
R80476 VSS.n8653 VSS.n1510 0.00476
R80477 VSS.n8659 VSS.n1510 0.00476
R80478 VSS.n8660 VSS.n8659 0.00476
R80479 VSS.n8661 VSS.n8660 0.00476
R80480 VSS.n8661 VSS.n1497 0.00476
R80481 VSS.n8687 VSS.n1464 0.00476
R80482 VSS.n8713 VSS.n1440 0.00476
R80483 VSS.n8719 VSS.n1440 0.00476
R80484 VSS.n8720 VSS.n8719 0.00476
R80485 VSS.n8721 VSS.n8720 0.00476
R80486 VSS.n8721 VSS.n1436 0.00476
R80487 VSS.n8727 VSS.n1436 0.00476
R80488 VSS.n8728 VSS.n8727 0.00476
R80489 VSS.n8729 VSS.n8728 0.00476
R80490 VSS.n8737 VSS.n8736 0.00476
R80491 VSS.n8738 VSS.n8737 0.00476
R80492 VSS.n8738 VSS.n1395 0.00476
R80493 VSS.n8789 VSS.n8788 0.00476
R80494 VSS.n8788 VSS.n8787 0.00476
R80495 VSS.n8787 VSS.n8747 0.00476
R80496 VSS.n8783 VSS.n8747 0.00476
R80497 VSS.n8783 VSS.n8782 0.00476
R80498 VSS.n8782 VSS.n8781 0.00476
R80499 VSS.n8781 VSS.n8753 0.00476
R80500 VSS.n8777 VSS.n8753 0.00476
R80501 VSS.n8777 VSS.n8776 0.00476
R80502 VSS.n8776 VSS.n8775 0.00476
R80503 VSS.n8775 VSS.n8759 0.00476
R80504 VSS.n8771 VSS.n8759 0.00476
R80505 VSS.n8957 VSS.n8956 0.00476
R80506 VSS.n8956 VSS.n8955 0.00476
R80507 VSS.n8955 VSS.n1144 0.00476
R80508 VSS.n8947 VSS.n8912 0.00476
R80509 VSS.n8943 VSS.n8912 0.00476
R80510 VSS.n8943 VSS.n8942 0.00476
R80511 VSS.n6552 VSS.n6551 0.00476
R80512 VSS.n6551 VSS.n6550 0.00476
R80513 VSS.n6550 VSS.n3273 0.00476
R80514 VSS.n6546 VSS.n3273 0.00476
R80515 VSS.n6539 VSS.n6538 0.00476
R80516 VSS.n6538 VSS.n6537 0.00476
R80517 VSS.n6537 VSS.n3335 0.00476
R80518 VSS.n6533 VSS.n3335 0.00476
R80519 VSS.n6526 VSS.n6525 0.00476
R80520 VSS.n6525 VSS.n6524 0.00476
R80521 VSS.n6524 VSS.n3397 0.00476
R80522 VSS.n6520 VSS.n3397 0.00476
R80523 VSS.n6520 VSS.n6519 0.00476
R80524 VSS.n6519 VSS.n6518 0.00476
R80525 VSS.n6518 VSS.n3403 0.00476
R80526 VSS.n6514 VSS.n3403 0.00476
R80527 VSS.n6514 VSS.n6513 0.00476
R80528 VSS.n6513 VSS.n6512 0.00476
R80529 VSS.n6512 VSS.n3409 0.00476
R80530 VSS.n6508 VSS.n3409 0.00476
R80531 VSS.n6501 VSS.n6500 0.00476
R80532 VSS.n6500 VSS.n6499 0.00476
R80533 VSS.n6499 VSS.n3471 0.00476
R80534 VSS.n6495 VSS.n3471 0.00476
R80535 VSS.n6495 VSS.n6494 0.00476
R80536 VSS.n6494 VSS.n6493 0.00476
R80537 VSS.n6493 VSS.n3477 0.00476
R80538 VSS.n6489 VSS.n3477 0.00476
R80539 VSS.n6489 VSS.n6488 0.00476
R80540 VSS.n6488 VSS.n6487 0.00476
R80541 VSS.n6487 VSS.n3483 0.00476
R80542 VSS.n3483 VSS.n3166 0.00476
R80543 VSS.n6478 VSS.n3136 0.00476
R80544 VSS.n6472 VSS.n6471 0.00476
R80545 VSS.n6471 VSS.n6470 0.00476
R80546 VSS.n6470 VSS.n3496 0.00476
R80547 VSS.n6466 VSS.n3496 0.00476
R80548 VSS.n6466 VSS.n6465 0.00476
R80549 VSS.n6465 VSS.n6464 0.00476
R80550 VSS.n6464 VSS.n3502 0.00476
R80551 VSS.n6460 VSS.n3502 0.00476
R80552 VSS.n6460 VSS.n6459 0.00476
R80553 VSS.n6459 VSS.n6458 0.00476
R80554 VSS.n6458 VSS.n3508 0.00476
R80555 VSS.n6454 VSS.n3508 0.00476
R80556 VSS.n6447 VSS.n6446 0.00476
R80557 VSS.n6446 VSS.n6445 0.00476
R80558 VSS.n6445 VSS.n3570 0.00476
R80559 VSS.n6441 VSS.n3570 0.00476
R80560 VSS.n6441 VSS.n6440 0.00476
R80561 VSS.n6440 VSS.n6439 0.00476
R80562 VSS.n6439 VSS.n3576 0.00476
R80563 VSS.n6435 VSS.n3576 0.00476
R80564 VSS.n6435 VSS.n6434 0.00476
R80565 VSS.n6434 VSS.n6433 0.00476
R80566 VSS.n6433 VSS.n3582 0.00476
R80567 VSS.n6429 VSS.n3582 0.00476
R80568 VSS.n6413 VSS.n3627 0.00476
R80569 VSS.n6409 VSS.n3627 0.00476
R80570 VSS.n6409 VSS.n6408 0.00476
R80571 VSS.n6408 VSS.n6407 0.00476
R80572 VSS.n6395 VSS.n6360 0.00476
R80573 VSS.n6391 VSS.n6360 0.00476
R80574 VSS.n6391 VSS.n6390 0.00476
R80575 VSS.n4459 VSS.n4456 0.00472535
R80576 VSS.n5117 VSS.n4432 0.00472535
R80577 DVSS VSS.n9537 0.00458
R80578 VSS.n9536 DVSS 0.00458
R80579 VSS.n2389 VSS.n1859 0.0045748
R80580 VSS.n9413 VSS.n705 0.0045748
R80581 VSS.n6213 VSS.n3901 0.00455
R80582 VSS.n6218 VSS.n3887 0.00455
R80583 VSS.n3738 VSS.n3156 0.00451408
R80584 VSS.n3763 VSS.n3186 0.00451408
R80585 VSS.n4714 VSS.n4588 0.00451408
R80586 VSS.n4699 VSS.n4631 0.00451408
R80587 VSS.n5227 VSS.n4339 0.00451408
R80588 VSS.n5200 VSS.n4394 0.00451408
R80589 VSS.n8647 VSS.n937 0.0045
R80590 VSS.n8732 VSS.n862 0.0045
R80591 VSS.n7946 VSS.n2135 0.0045
R80592 VSS.n9177 VSS.n937 0.0045
R80593 VSS.n9276 VSS.n862 0.0045
R80594 VSS.n9509 VSS.n718 0.0045
R80595 VSS.n9510 VSS.n9509 0.0045
R80596 VSS.n7947 VSS.n7946 0.0045
R80597 VSS.n9221 VSS.n916 0.00446
R80598 VSS.n9159 VSS.n956 0.00446
R80599 VSS.n8684 VSS.n1497 0.00446
R80600 VSS.n6609 VSS.n3166 0.00446
R80601 VSS.n6215 VSS.n3901 0.00442143
R80602 VSS.n6221 VSS.n3887 0.00442143
R80603 VSS.n9257 VSS.n9256 0.00434
R80604 VSS.n9109 VSS.n9078 0.00434
R80605 VSS.n8713 VSS.n8712 0.00434
R80606 VSS.n6472 VSS.n3135 0.00434
R80607 VSS.n1385 VSS.n1365 0.00430282
R80608 VSS.n8396 VSS.n1630 0.00430282
R80609 VSS.n9892 VSS.n41 0.00423239
R80610 VSS.n9888 VSS.n34 0.00423239
R80611 VSS.n9864 VSS.n74 0.00423239
R80612 VSS.n9861 VSS.n85 0.00423239
R80613 VSS.n9849 VSS.n105 0.00423239
R80614 VSS.n9846 VSS.n116 0.00423239
R80615 VSS.n9834 VSS.n136 0.00423239
R80616 VSS.n9829 VSS.n9822 0.00423239
R80617 VSS.n8581 VSS.n8578 0.00422047
R80618 VSS.n2285 VSS.n2156 0.00422047
R80619 VSS.n2379 VSS.n1861 0.00422047
R80620 VSS.n8587 VSS.n1401 0.00422047
R80621 VSS.n8608 VSS.n8607 0.00422047
R80622 VSS.n8079 VSS.n8078 0.00422047
R80623 VSS.n6259 VSS.n3851 0.00422047
R80624 VSS.n4156 VSS.n420 0.00422047
R80625 VSS.n1211 VSS.n744 0.00422047
R80626 VSS.n9423 VSS.n707 0.00422047
R80627 VSS.n8302 VSS.n8301 0.00416429
R80628 VSS.n8331 VSS.n8330 0.00416429
R80629 VSS.n8347 VSS.n1569 0.00416429
R80630 VSS.n8413 VSS.n8412 0.00416429
R80631 VSS.n6960 VSS.n2814 0.00416429
R80632 VSS.n6938 VSS.n2836 0.00416429
R80633 VSS.n6915 VSS.n2862 0.00416429
R80634 VSS.n6876 VSS.n2896 0.00416429
R80635 VSS.n3919 VSS.n3834 0.00416429
R80636 VSS.n6195 VSS.n3957 0.00416429
R80637 VSS.n6159 VSS.n3986 0.00416429
R80638 VSS.n3874 VSS.n3867 0.00416429
R80639 VSS.n5304 VSS.n5303 0.00416429
R80640 VSS.n5624 VSS.n4290 0.00416429
R80641 VSS.n4765 VSS.n4764 0.00416429
R80642 VSS.n4787 VSS.n4786 0.00416429
R80643 VSS.n4803 VSS.n4331 0.00416429
R80644 VSS.n5054 VSS.n4523 0.00416429
R80645 VSS.n3728 VSS.n3146 0.00409155
R80646 VSS.n6793 VSS.n2952 0.00409155
R80647 VSS.n3783 VSS.n3176 0.00409155
R80648 VSS.n6794 VSS.n2934 0.00409155
R80649 VSS.n8959 VSS.n8958 0.00404
R80650 VSS.n9507 VSS.n721 0.00404
R80651 VSS.n9512 VSS.n716 0.00404
R80652 VSS.n9513 VSS.n715 0.00404
R80653 VSS.n9506 VSS.n723 0.00404
R80654 VSS.n8957 VSS.n1139 0.00404
R80655 VSS.n7854 VSS.n7598 0.00403571
R80656 VSS.n7595 VSS.n7594 0.00403571
R80657 VSS.n4448 VSS.n4440 0.00402113
R80658 VSS.n4718 VSS.n4717 0.0039507
R80659 VSS.n4703 VSS.n4702 0.0039507
R80660 VSS.n5231 VSS.n5230 0.0039507
R80661 VSS.n5204 VSS.n5203 0.0039507
R80662 VSS.n6389 DVSS 0.00392
R80663 VSS.n8941 DVSS 0.00392
R80664 VSS.n9218 VSS.n9197 0.00392
R80665 VSS.n9156 VSS.n9155 0.00392
R80666 VSS.n8667 VSS.n1495 0.00392
R80667 VSS.n8942 DVSS 0.00392
R80668 VSS.n6480 VSS.n3179 0.00392
R80669 VSS.n6390 DVSS 0.00392
R80670 VSS.n8842 VSS.n1331 0.00390714
R80671 VSS.n8498 VSS.n1324 0.00390714
R80672 VSS.n8859 VSS.n1309 0.00390714
R80673 VSS.n8862 VSS.n8861 0.00390714
R80674 VSS.n8909 VSS.n1267 0.00390714
R80675 VSS.n8878 VSS.n1260 0.00390714
R80676 VSS.n9569 VSS.n548 0.00390714
R80677 VSS.n8887 VSS.n541 0.00390714
R80678 VSS.n6751 VSS.n2981 0.00390714
R80679 VSS.n6748 VSS.n2974 0.00390714
R80680 VSS.n6717 VSS.n3063 0.00390714
R80681 VSS.n6715 VSS.n3076 0.00390714
R80682 VSS.n6700 VSS.n3092 0.00390714
R80683 VSS.n6697 VSS.n3098 0.00390714
R80684 VSS.n9582 VSS.n510 0.00390714
R80685 VSS.n6676 VSS.n503 0.00390714
R80686 VSS.n9680 VSS.n317 0.00390714
R80687 VSS.n9677 VSS.n310 0.00390714
R80688 VSS.n9646 VSS.n351 0.00390714
R80689 VSS.n370 VSS.n358 0.00390714
R80690 VSS.n380 VSS.n376 0.00390714
R80691 VSS.n9629 VSS.n9628 0.00390714
R80692 VSS.n406 VSS.n402 0.00390714
R80693 VSS.n9609 VSS.n9608 0.00390714
R80694 VSS.n9683 VSS.n295 0.00390714
R80695 VSS.n5559 VSS.n289 0.00390714
R80696 VSS.n5528 VSS.n5379 0.00390714
R80697 VSS.n5525 VSS.n5385 0.00390714
R80698 VSS.n5406 VSS.n5402 0.00390714
R80699 VSS.n5507 VSS.n5506 0.00390714
R80700 VSS.n5430 VSS.n5426 0.00390714
R80701 VSS.n5486 VSS.n5485 0.00390714
R80702 VSS.n9694 VSS.n263 0.00390714
R80703 VSS.n268 VSS.n250 0.00390714
R80704 VSS.n9758 VSS.n9747 0.00390714
R80705 VSS.n234 VSS.n228 0.00390714
R80706 VSS.n9776 VSS.n211 0.00390714
R80707 VSS.n203 VSS.n194 0.00390714
R80708 VSS.n9809 VSS.n9797 0.00390714
R80709 VSS.n186 VSS.n179 0.00390714
R80710 VSS.n2321 VSS.n2164 0.00386614
R80711 VSS.n2405 VSS.n1846 0.00386614
R80712 VSS.n4763 VSS.n4730 0.00386614
R80713 VSS.n9813 VSS.n172 0.00386614
R80714 VSS.n1175 VSS.n752 0.00386614
R80715 VSS.n9397 VSS.n693 0.00386614
R80716 VSS.n8246 VSS.n8245 0.00383
R80717 VSS.n8235 VSS.n1880 0.00383
R80718 VSS.n8205 VSS.n1949 0.00383
R80719 VSS.n7929 VSS.n7893 0.00383
R80720 VSS.n8101 VSS.n2080 0.00383
R80721 VSS.n8163 VSS.n1981 0.00383
R80722 VSS.n2256 VSS.n2176 0.00383
R80723 VSS.n7952 VSS.n2090 0.00383
R80724 VSS.n7981 VSS.n1541 0.00383
R80725 VSS.n6546 VSS.n6545 0.00383
R80726 VSS.n6533 VSS.n6532 0.00383
R80727 VSS.n6508 VSS.n6507 0.00383
R80728 VSS.n8735 VSS.n1011 0.0038
R80729 VSS.n9064 VSS.n9063 0.0038
R80730 VSS.n9278 VSS.n861 0.0038
R80731 VSS.n9250 VSS.n873 0.0038
R80732 VSS.n9279 VSS.n860 0.0038
R80733 VSS.n9114 VSS.n982 0.0038
R80734 VSS.n9062 VSS.n1008 0.0038
R80735 VSS.n1462 VSS.n1444 0.0038
R80736 VSS.n8736 VSS.n1433 0.0038
R80737 VSS.n6474 VSS.n3161 0.0038
R80738 VSS.n5177 VSS.n5176 0.00373944
R80739 VSS.n1637 VSS.n1368 0.00371429
R80740 VSS.n6805 VSS.n2942 0.00371429
R80741 VSS.n4180 VSS.n4171 0.00371429
R80742 VSS.n5669 VSS.n4247 0.00371429
R80743 VSS.n5021 VSS.n5020 0.00371429
R80744 VSS.n9314 VSS.n827 0.00371
R80745 VSS.n9347 VSS.n780 0.00371
R80746 VSS.n9526 VSS.n681 0.00371
R80747 VSS.n9050 VSS.n9038 0.00371
R80748 VSS.n9011 VSS.n9000 0.00371
R80749 VSS.n9493 VSS.n755 0.00371
R80750 VSS.n8789 VSS.n1393 0.00371
R80751 VSS.n8962 VSS.n8961 0.00371
R80752 VSS.n8948 VSS.n8947 0.00371
R80753 VSS.n6447 VSS.n3550 0.00371
R80754 VSS.n6424 VSS.n6413 0.00371
R80755 VSS.n6396 VSS.n6395 0.00371
R80756 VSS.n8854 VSS.n1301 0.00368898
R80757 VSS.n1338 VSS.n1315 0.00368898
R80758 VSS.n8405 VSS.n8404 0.00368898
R80759 VSS.n8561 VSS.n1567 0.00368898
R80760 VSS.n3730 VSS.n3145 0.00366901
R80761 VSS.n6788 VSS.n2951 0.00366901
R80762 VSS.n3780 VSS.n3175 0.00366901
R80763 VSS.n6790 VSS.n2933 0.00366901
R80764 VSS.n8294 VSS.n8293 0.00365
R80765 VSS.n8323 VSS.n8322 0.00365
R80766 VSS.n8345 VSS.n1568 0.00365
R80767 VSS.n8410 VSS.n8384 0.00365
R80768 VSS.n2819 VSS.n2797 0.00365
R80769 VSS.n6942 VSS.n2830 0.00365
R80770 VSS.n6919 VSS.n2856 0.00365
R80771 VSS.n6880 VSS.n2890 0.00365
R80772 VSS.n3917 VSS.n3833 0.00365
R80773 VSS.n3961 VSS.n3956 0.00365
R80774 VSS.n6162 VSS.n3980 0.00365
R80775 VSS.n6235 VSS.n3866 0.00365
R80776 VSS.n5296 VSS.n5295 0.00365
R80777 VSS.n4297 VSS.n4289 0.00365
R80778 VSS.n4729 VSS.n4728 0.00365
R80779 VSS.n4563 VSS.n4562 0.00365
R80780 VSS.n4801 VSS.n4330 0.00365
R80781 VSS.n4530 VSS.n4522 0.00365
R80782 VSS.n1518 VSS.n1515 0.00356
R80783 VSS.n9170 VSS.n945 0.00356
R80784 VSS.n940 VSS.n936 0.00356
R80785 VSS.n9173 VSS.n935 0.00356
R80786 VSS.n9172 VSS.n9171 0.00356
R80787 VSS.n1514 VSS.n942 0.00356
R80788 DVSS VSS.n9486 0.00353
R80789 VSS.n2301 VSS.n2149 0.00351181
R80790 VSS.n1195 VSS.n736 0.00351181
R80791 VSS.n8821 VSS.n8817 0.00345775
R80792 VSS.n8401 VSS.n1632 0.00345775
R80793 VSS.n8535 VSS.n8534 0.00345714
R80794 VSS.n6840 VSS.n2930 0.00345714
R80795 VSS.n6125 VSS.n4020 0.00345714
R80796 VSS.n5346 VSS.n4264 0.00345714
R80797 VSS.n4848 VSS.n4493 0.00345714
R80798 VSS.n5099 DVSS 0.003425
R80799 VSS.n4942 DVSS 0.003425
R80800 VSS.n5692 DVSS 0.003425
R80801 DVSS VSS.n4050 0.003425
R80802 DVSS VSS.n5980 0.003425
R80803 VSS.n3768 DVSS 0.003425
R80804 VSS.n5856 DVSS 0.003425
R80805 VSS.n6837 DVSS 0.003425
R80806 DVSS VSS.n2678 0.003425
R80807 VSS.n9223 VSS.n901 0.00338
R80808 VSS.n9150 VSS.n961 0.00338
R80809 VSS.n8686 VSS.n1477 0.00338
R80810 VSS.n6481 VSS.n3165 0.00338
R80811 VSS.n3270 VSS.n3269 0.00334
R80812 VSS.n3271 VSS.n3270 0.00334
R80813 VSS.n3274 VSS.n3271 0.00334
R80814 VSS.n3275 VSS.n3274 0.00334
R80815 VSS.n3276 VSS.n3275 0.00334
R80816 VSS.n3277 VSS.n3276 0.00334
R80817 VSS.n3330 VSS.n3277 0.00334
R80818 VSS.n3331 VSS.n3330 0.00334
R80819 VSS.n3332 VSS.n3331 0.00334
R80820 VSS.n3333 VSS.n3332 0.00334
R80821 VSS.n3336 VSS.n3333 0.00334
R80822 VSS.n3337 VSS.n3336 0.00334
R80823 VSS.n3338 VSS.n3337 0.00334
R80824 VSS.n3339 VSS.n3338 0.00334
R80825 VSS.n3392 VSS.n3339 0.00334
R80826 VSS.n3393 VSS.n3392 0.00334
R80827 VSS.n3394 VSS.n3393 0.00334
R80828 VSS.n3395 VSS.n3394 0.00334
R80829 VSS.n3398 VSS.n3395 0.00334
R80830 VSS.n3399 VSS.n3398 0.00334
R80831 VSS.n3400 VSS.n3399 0.00334
R80832 VSS.n3401 VSS.n3400 0.00334
R80833 VSS.n3404 VSS.n3401 0.00334
R80834 VSS.n3405 VSS.n3404 0.00334
R80835 VSS.n3406 VSS.n3405 0.00334
R80836 VSS.n3407 VSS.n3406 0.00334
R80837 VSS.n3410 VSS.n3407 0.00334
R80838 VSS.n3411 VSS.n3410 0.00334
R80839 VSS.n3412 VSS.n3411 0.00334
R80840 VSS.n3413 VSS.n3412 0.00334
R80841 VSS.n3466 VSS.n3413 0.00334
R80842 VSS.n3467 VSS.n3466 0.00334
R80843 VSS.n3468 VSS.n3467 0.00334
R80844 VSS.n3469 VSS.n3468 0.00334
R80845 VSS.n3472 VSS.n3469 0.00334
R80846 VSS.n3473 VSS.n3472 0.00334
R80847 VSS.n3474 VSS.n3473 0.00334
R80848 VSS.n3475 VSS.n3474 0.00334
R80849 VSS.n3478 VSS.n3475 0.00334
R80850 VSS.n3479 VSS.n3478 0.00334
R80851 VSS.n3480 VSS.n3479 0.00334
R80852 VSS.n3481 VSS.n3480 0.00334
R80853 VSS.n3484 VSS.n3481 0.00334
R80854 VSS.n3485 VSS.n3484 0.00334
R80855 VSS.n3486 VSS.n3485 0.00334
R80856 VSS.n3487 VSS.n3486 0.00334
R80857 VSS.n3488 VSS.n3487 0.00334
R80858 VSS.n3489 VSS.n3488 0.00334
R80859 VSS.n3490 VSS.n3489 0.00334
R80860 VSS.n3491 VSS.n3490 0.00334
R80861 VSS.n3492 VSS.n3491 0.00334
R80862 VSS.n3493 VSS.n3492 0.00334
R80863 VSS.n3494 VSS.n3493 0.00334
R80864 VSS.n3497 VSS.n3494 0.00334
R80865 VSS.n3498 VSS.n3497 0.00334
R80866 VSS.n3499 VSS.n3498 0.00334
R80867 VSS.n3500 VSS.n3499 0.00334
R80868 VSS.n3503 VSS.n3500 0.00334
R80869 VSS.n3504 VSS.n3503 0.00334
R80870 VSS.n3505 VSS.n3504 0.00334
R80871 VSS.n3506 VSS.n3505 0.00334
R80872 VSS.n3509 VSS.n3506 0.00334
R80873 VSS.n3510 VSS.n3509 0.00334
R80874 VSS.n3511 VSS.n3510 0.00334
R80875 VSS.n3512 VSS.n3511 0.00334
R80876 VSS.n3565 VSS.n3512 0.00334
R80877 VSS.n3566 VSS.n3565 0.00334
R80878 VSS.n3567 VSS.n3566 0.00334
R80879 VSS.n3568 VSS.n3567 0.00334
R80880 VSS.n3571 VSS.n3568 0.00334
R80881 VSS.n3572 VSS.n3571 0.00334
R80882 VSS.n3573 VSS.n3572 0.00334
R80883 VSS.n3574 VSS.n3573 0.00334
R80884 VSS.n3577 VSS.n3574 0.00334
R80885 VSS.n3578 VSS.n3577 0.00334
R80886 VSS.n3579 VSS.n3578 0.00334
R80887 VSS.n3580 VSS.n3579 0.00334
R80888 VSS.n3583 VSS.n3580 0.00334
R80889 VSS.n3584 VSS.n3583 0.00334
R80890 VSS.n3585 VSS.n3584 0.00334
R80891 VSS.n3586 VSS.n3585 0.00334
R80892 VSS.n3629 VSS.n3586 0.00334
R80893 VSS.n3631 VSS.n3629 0.00334
R80894 VSS.n3632 VSS.n3631 0.00334
R80895 VSS.n3633 VSS.n3632 0.00334
R80896 VSS.n3634 VSS.n3633 0.00334
R80897 VSS.n3635 VSS.n3634 0.00334
R80898 VSS.n3638 VSS.n3635 0.00334
R80899 VSS.n3639 VSS.n3638 0.00334
R80900 VSS.n3640 VSS.n3639 0.00334
R80901 VSS.n6362 VSS.n3640 0.00334
R80902 VSS.n6363 VSS.n6362 0.00334
R80903 VSS.n6364 VSS.n6363 0.00334
R80904 VSS.n6365 VSS.n6364 0.00334
R80905 VSS.n6366 VSS.n6365 0.00334
R80906 VSS.n6367 VSS.n6366 0.00334
R80907 VSS.n6370 VSS.n6369 0.00334
R80908 VSS.n1830 VSS.n1829 0.00334
R80909 VSS.n1831 VSS.n1830 0.00334
R80910 VSS.n1834 VSS.n1831 0.00334
R80911 VSS.n1835 VSS.n1834 0.00334
R80912 VSS.n1836 VSS.n1835 0.00334
R80913 VSS.n1837 VSS.n1836 0.00334
R80914 VSS.n1870 VSS.n1837 0.00334
R80915 VSS.n1873 VSS.n1870 0.00334
R80916 VSS.n1874 VSS.n1873 0.00334
R80917 VSS.n1875 VSS.n1874 0.00334
R80918 VSS.n1876 VSS.n1875 0.00334
R80919 VSS.n1877 VSS.n1876 0.00334
R80920 VSS.n2134 VSS.n1877 0.00334
R80921 VSS.n1883 VSS.n1882 0.00334
R80922 VSS.n1931 VSS.n1883 0.00334
R80923 VSS.n1932 VSS.n1931 0.00334
R80924 VSS.n1933 VSS.n1932 0.00334
R80925 VSS.n1934 VSS.n1933 0.00334
R80926 VSS.n1935 VSS.n1934 0.00334
R80927 VSS.n1938 VSS.n1935 0.00334
R80928 VSS.n1939 VSS.n1938 0.00334
R80929 VSS.n1940 VSS.n1939 0.00334
R80930 VSS.n1941 VSS.n1940 0.00334
R80931 VSS.n1944 VSS.n1941 0.00334
R80932 VSS.n1945 VSS.n1944 0.00334
R80933 VSS.n1946 VSS.n1945 0.00334
R80934 VSS.n1947 VSS.n1946 0.00334
R80935 VSS.n1950 VSS.n1947 0.00334
R80936 VSS.n1951 VSS.n1950 0.00334
R80937 VSS.n1952 VSS.n1951 0.00334
R80938 VSS.n8187 VSS.n1952 0.00334
R80939 VSS.n8188 VSS.n8187 0.00334
R80940 VSS.n8189 VSS.n8188 0.00334
R80941 VSS.n8190 VSS.n8189 0.00334
R80942 VSS.n8190 VSS.n938 0.00334
R80943 VSS.n9176 VSS.n938 0.00334
R80944 VSS.n9179 VSS.n9178 0.00334
R80945 VSS.n9179 VSS.n933 0.00334
R80946 VSS.n9185 VSS.n933 0.00334
R80947 VSS.n9186 VSS.n9185 0.00334
R80948 VSS.n9187 VSS.n9186 0.00334
R80949 VSS.n9187 VSS.n929 0.00334
R80950 VSS.n9193 VSS.n929 0.00334
R80951 VSS.n9194 VSS.n9193 0.00334
R80952 VSS.n9195 VSS.n9194 0.00334
R80953 VSS.n9195 VSS.n899 0.00334
R80954 VSS.n9226 VSS.n899 0.00334
R80955 VSS.n9227 VSS.n9226 0.00334
R80956 VSS.n9228 VSS.n9227 0.00334
R80957 VSS.n9228 VSS.n871 0.00334
R80958 VSS.n9259 VSS.n871 0.00334
R80959 VSS.n9260 VSS.n9259 0.00334
R80960 VSS.n9261 VSS.n9260 0.00334
R80961 VSS.n9261 VSS.n867 0.00334
R80962 VSS.n9267 VSS.n867 0.00334
R80963 VSS.n9268 VSS.n9267 0.00334
R80964 VSS.n9269 VSS.n9268 0.00334
R80965 VSS.n9269 VSS.n863 0.00334
R80966 VSS.n9275 VSS.n863 0.00334
R80967 VSS.n9277 VSS.n858 0.00334
R80968 VSS.n9283 VSS.n858 0.00334
R80969 VSS.n9284 VSS.n9283 0.00334
R80970 VSS.n9285 VSS.n9284 0.00334
R80971 VSS.n9285 VSS.n829 0.00334
R80972 VSS.n9317 VSS.n829 0.00334
R80973 VSS.n9318 VSS.n9317 0.00334
R80974 VSS.n9319 VSS.n9318 0.00334
R80975 VSS.n9319 VSS.n825 0.00334
R80976 VSS.n9325 VSS.n825 0.00334
R80977 VSS.n9326 VSS.n9325 0.00334
R80978 VSS.n9327 VSS.n9326 0.00334
R80979 VSS.n9327 VSS.n821 0.00334
R80980 VSS.n9333 VSS.n821 0.00334
R80981 VSS.n9334 VSS.n9333 0.00334
R80982 VSS.n9336 VSS.n9334 0.00334
R80983 VSS.n9336 VSS.n9335 0.00334
R80984 VSS.n9335 VSS.n817 0.00334
R80985 VSS.n9343 VSS.n817 0.00334
R80986 VSS.n9344 VSS.n9343 0.00334
R80987 VSS.n9345 VSS.n9344 0.00334
R80988 VSS.n9346 VSS.n9345 0.00334
R80989 VSS.n9346 VSS.n717 0.00334
R80990 VSS.n9511 VSS.n713 0.00334
R80991 VSS.n9518 VSS.n713 0.00334
R80992 VSS.n9519 VSS.n9518 0.00334
R80993 VSS.n9520 VSS.n9519 0.00334
R80994 VSS.n9520 VSS.n683 0.00334
R80995 VSS.n9529 VSS.n683 0.00334
R80996 VSS.n9530 VSS.n9529 0.00334
R80997 VSS.n9532 VSS.n9530 0.00334
R80998 VSS.n9532 VSS.n9531 0.00334
R80999 VSS.n9531 VSS.n680 0.00334
R81000 VSS.n9541 VSS.n9540 0.00334
R81001 VSS.n7916 VSS.n7899 0.00334
R81002 VSS.n7917 VSS.n7916 0.00334
R81003 VSS.n7918 VSS.n7917 0.00334
R81004 VSS.n7918 VSS.n7895 0.00334
R81005 VSS.n7924 VSS.n7895 0.00334
R81006 VSS.n7925 VSS.n7924 0.00334
R81007 VSS.n7926 VSS.n7925 0.00334
R81008 VSS.n7926 VSS.n2140 0.00334
R81009 VSS.n7934 VSS.n2140 0.00334
R81010 VSS.n7935 VSS.n7934 0.00334
R81011 VSS.n7937 VSS.n7935 0.00334
R81012 VSS.n7937 VSS.n7936 0.00334
R81013 VSS.n7936 VSS.n2136 0.00334
R81014 VSS.n7945 VSS.n2033 0.00334
R81015 VSS.n8106 VSS.n2033 0.00334
R81016 VSS.n8107 VSS.n8106 0.00334
R81017 VSS.n8108 VSS.n8107 0.00334
R81018 VSS.n8108 VSS.n2029 0.00334
R81019 VSS.n8114 VSS.n2029 0.00334
R81020 VSS.n8115 VSS.n8114 0.00334
R81021 VSS.n8116 VSS.n8115 0.00334
R81022 VSS.n8116 VSS.n2025 0.00334
R81023 VSS.n8122 VSS.n2025 0.00334
R81024 VSS.n8123 VSS.n8122 0.00334
R81025 VSS.n8124 VSS.n8123 0.00334
R81026 VSS.n8124 VSS.n2021 0.00334
R81027 VSS.n8131 VSS.n2021 0.00334
R81028 VSS.n8132 VSS.n8131 0.00334
R81029 VSS.n8133 VSS.n8132 0.00334
R81030 VSS.n8133 VSS.n2019 0.00334
R81031 VSS.n8138 VSS.n2019 0.00334
R81032 VSS.n8139 VSS.n8138 0.00334
R81033 VSS.n8140 VSS.n8139 0.00334
R81034 VSS.n8141 VSS.n8140 0.00334
R81035 VSS.n8142 VSS.n8141 0.00334
R81036 VSS.n8143 VSS.n8142 0.00334
R81037 VSS.n947 VSS.n946 0.00334
R81038 VSS.n948 VSS.n947 0.00334
R81039 VSS.n951 VSS.n948 0.00334
R81040 VSS.n952 VSS.n951 0.00334
R81041 VSS.n953 VSS.n952 0.00334
R81042 VSS.n954 VSS.n953 0.00334
R81043 VSS.n957 VSS.n954 0.00334
R81044 VSS.n958 VSS.n957 0.00334
R81045 VSS.n959 VSS.n958 0.00334
R81046 VSS.n976 VSS.n959 0.00334
R81047 VSS.n977 VSS.n976 0.00334
R81048 VSS.n978 VSS.n977 0.00334
R81049 VSS.n979 VSS.n978 0.00334
R81050 VSS.n997 VSS.n979 0.00334
R81051 VSS.n998 VSS.n997 0.00334
R81052 VSS.n999 VSS.n998 0.00334
R81053 VSS.n1000 VSS.n999 0.00334
R81054 VSS.n1003 VSS.n1000 0.00334
R81055 VSS.n1004 VSS.n1003 0.00334
R81056 VSS.n1005 VSS.n1004 0.00334
R81057 VSS.n1006 VSS.n1005 0.00334
R81058 VSS.n1009 VSS.n1006 0.00334
R81059 VSS.n1010 VSS.n1009 0.00334
R81060 VSS.n1015 VSS.n1012 0.00334
R81061 VSS.n1016 VSS.n1015 0.00334
R81062 VSS.n1017 VSS.n1016 0.00334
R81063 VSS.n1018 VSS.n1017 0.00334
R81064 VSS.n1057 VSS.n1018 0.00334
R81065 VSS.n1058 VSS.n1057 0.00334
R81066 VSS.n1059 VSS.n1058 0.00334
R81067 VSS.n1060 VSS.n1059 0.00334
R81068 VSS.n1061 VSS.n1060 0.00334
R81069 VSS.n1064 VSS.n1061 0.00334
R81070 VSS.n1065 VSS.n1064 0.00334
R81071 VSS.n1066 VSS.n1065 0.00334
R81072 VSS.n1067 VSS.n1066 0.00334
R81073 VSS.n1070 VSS.n1067 0.00334
R81074 VSS.n1071 VSS.n1070 0.00334
R81075 VSS.n1072 VSS.n1071 0.00334
R81076 VSS.n1073 VSS.n1072 0.00334
R81077 VSS.n1076 VSS.n1073 0.00334
R81078 VSS.n1077 VSS.n1076 0.00334
R81079 VSS.n1078 VSS.n1077 0.00334
R81080 VSS.n8996 VSS.n1078 0.00334
R81081 VSS.n8997 VSS.n8996 0.00334
R81082 VSS.n8997 VSS.n719 0.00334
R81083 VSS.n9508 VSS.n720 0.00334
R81084 VSS.n725 VSS.n720 0.00334
R81085 VSS.n726 VSS.n725 0.00334
R81086 VSS.n727 VSS.n726 0.00334
R81087 VSS.n9459 VSS.n727 0.00334
R81088 VSS.n9460 VSS.n9459 0.00334
R81089 VSS.n9461 VSS.n9460 0.00334
R81090 VSS.n9464 VSS.n9461 0.00334
R81091 VSS.n9465 VSS.n9464 0.00334
R81092 VSS.n9466 VSS.n9465 0.00334
R81093 VSS.n9467 VSS.n9466 0.00334
R81094 VSS.n9469 VSS.n9468 0.00334
R81095 VSS.n2231 VSS.n2229 0.00334
R81096 VSS.n2249 VSS.n2229 0.00334
R81097 VSS.n2250 VSS.n2249 0.00334
R81098 VSS.n2252 VSS.n2250 0.00334
R81099 VSS.n2252 VSS.n2251 0.00334
R81100 VSS.n2251 VSS.n2226 0.00334
R81101 VSS.n2226 VSS.n2224 0.00334
R81102 VSS.n2262 VSS.n2224 0.00334
R81103 VSS.n2263 VSS.n2262 0.00334
R81104 VSS.n2264 VSS.n2263 0.00334
R81105 VSS.n2265 VSS.n2264 0.00334
R81106 VSS.n2265 VSS.n2133 0.00334
R81107 VSS.n7948 VSS.n2133 0.00334
R81108 VSS.n2130 VSS.n2128 0.00334
R81109 VSS.n7958 VSS.n2128 0.00334
R81110 VSS.n7959 VSS.n7958 0.00334
R81111 VSS.n7960 VSS.n7959 0.00334
R81112 VSS.n7961 VSS.n7960 0.00334
R81113 VSS.n7962 VSS.n7961 0.00334
R81114 VSS.n7965 VSS.n7962 0.00334
R81115 VSS.n7966 VSS.n7965 0.00334
R81116 VSS.n7967 VSS.n7966 0.00334
R81117 VSS.n7968 VSS.n7967 0.00334
R81118 VSS.n7971 VSS.n7968 0.00334
R81119 VSS.n7972 VSS.n7971 0.00334
R81120 VSS.n7973 VSS.n7972 0.00334
R81121 VSS.n7974 VSS.n7973 0.00334
R81122 VSS.n7976 VSS.n7974 0.00334
R81123 VSS.n7977 VSS.n7976 0.00334
R81124 VSS.n7978 VSS.n7977 0.00334
R81125 VSS.n7978 VSS.n1521 0.00334
R81126 VSS.n8638 VSS.n1521 0.00334
R81127 VSS.n8639 VSS.n8638 0.00334
R81128 VSS.n8640 VSS.n8639 0.00334
R81129 VSS.n8640 VSS.n1516 0.00334
R81130 VSS.n8646 VSS.n1516 0.00334
R81131 VSS.n8649 VSS.n8648 0.00334
R81132 VSS.n8649 VSS.n1512 0.00334
R81133 VSS.n8655 VSS.n1512 0.00334
R81134 VSS.n8656 VSS.n8655 0.00334
R81135 VSS.n8657 VSS.n8656 0.00334
R81136 VSS.n8657 VSS.n1508 0.00334
R81137 VSS.n8663 VSS.n1508 0.00334
R81138 VSS.n8664 VSS.n8663 0.00334
R81139 VSS.n8665 VSS.n8664 0.00334
R81140 VSS.n8665 VSS.n1475 0.00334
R81141 VSS.n8689 VSS.n1475 0.00334
R81142 VSS.n8690 VSS.n8689 0.00334
R81143 VSS.n8691 VSS.n8690 0.00334
R81144 VSS.n8691 VSS.n1442 0.00334
R81145 VSS.n8715 VSS.n1442 0.00334
R81146 VSS.n8716 VSS.n8715 0.00334
R81147 VSS.n8717 VSS.n8716 0.00334
R81148 VSS.n8717 VSS.n1438 0.00334
R81149 VSS.n8723 VSS.n1438 0.00334
R81150 VSS.n8724 VSS.n8723 0.00334
R81151 VSS.n8725 VSS.n8724 0.00334
R81152 VSS.n8725 VSS.n1434 0.00334
R81153 VSS.n8731 VSS.n1434 0.00334
R81154 VSS.n8734 VSS.n8733 0.00334
R81155 VSS.n8733 VSS.n1431 0.00334
R81156 VSS.n8741 VSS.n1431 0.00334
R81157 VSS.n8742 VSS.n8741 0.00334
R81158 VSS.n8743 VSS.n8742 0.00334
R81159 VSS.n8744 VSS.n8743 0.00334
R81160 VSS.n8745 VSS.n8744 0.00334
R81161 VSS.n8748 VSS.n8745 0.00334
R81162 VSS.n8749 VSS.n8748 0.00334
R81163 VSS.n8750 VSS.n8749 0.00334
R81164 VSS.n8751 VSS.n8750 0.00334
R81165 VSS.n8754 VSS.n8751 0.00334
R81166 VSS.n8755 VSS.n8754 0.00334
R81167 VSS.n8756 VSS.n8755 0.00334
R81168 VSS.n8757 VSS.n8756 0.00334
R81169 VSS.n8760 VSS.n8757 0.00334
R81170 VSS.n8761 VSS.n8760 0.00334
R81171 VSS.n8762 VSS.n8761 0.00334
R81172 VSS.n8763 VSS.n8762 0.00334
R81173 VSS.n8764 VSS.n8763 0.00334
R81174 VSS.n8766 VSS.n8764 0.00334
R81175 VSS.n8766 VSS.n8765 0.00334
R81176 VSS.n8765 VSS.n1141 0.00334
R81177 VSS.n1145 VSS.n1142 0.00334
R81178 VSS.n1146 VSS.n1145 0.00334
R81179 VSS.n1147 VSS.n1146 0.00334
R81180 VSS.n1148 VSS.n1147 0.00334
R81181 VSS.n8914 VSS.n1148 0.00334
R81182 VSS.n8915 VSS.n8914 0.00334
R81183 VSS.n8916 VSS.n8915 0.00334
R81184 VSS.n8917 VSS.n8916 0.00334
R81185 VSS.n8918 VSS.n8917 0.00334
R81186 VSS.n8919 VSS.n8918 0.00334
R81187 VSS.n8920 VSS.n8919 0.00334
R81188 VSS.n8922 VSS.n8921 0.00334
R81189 VSS.n7953 VSS.n2129 0.00332
R81190 VSS.n7944 VSS.n7943 0.00332
R81191 VSS.n8234 VSS.n1881 0.00332
R81192 VSS.n8236 VSS.n8235 0.00332
R81193 VSS.n2080 VSS.n1879 0.00332
R81194 VSS.n7952 VSS.n7951 0.00332
R81195 VSS.n8268 VSS.n1805 0.00329
R81196 VSS.n1865 VSS.n1851 0.00329
R81197 VSS.n8232 VSS.n8231 0.00329
R81198 VSS.n8202 VSS.n8201 0.00329
R81199 VSS.n7911 VSS.n1766 0.00329
R81200 VSS.n7928 VSS.n2168 0.00329
R81201 VSS.n8098 VSS.n2035 0.00329
R81202 VSS.n1994 VSS.n1979 0.00329
R81203 VSS.n2242 VSS.n1727 0.00329
R81204 VSS.n2258 VSS.n2175 0.00329
R81205 VSS.n7954 VSS.n2091 0.00329
R81206 VSS.n8633 VSS.n1543 0.00329
R81207 VSS.n6568 VSS.n3247 0.00329
R81208 VSS.n3315 VSS.n3291 0.00329
R81209 VSS.n3389 VSS.n3353 0.00329
R81210 VSS.n3463 VSS.n3427 0.00329
R81211 VSS.n6369 DVSS 0.00326
R81212 VSS.n8921 DVSS 0.00326
R81213 VSS.n9253 VSS.n9230 0.00326
R81214 VSS.n9115 VSS.n981 0.00326
R81215 VSS.n8710 VSS.n8693 0.00326
R81216 VSS.n6615 VSS.n3149 0.00326
R81217 VSS.n4855 VSS.n4488 0.00324648
R81218 VSS.n3736 VSS.n3155 0.00324648
R81219 VSS.n5089 VSS.n4486 0.00324648
R81220 VSS.n3767 VSS.n3185 0.00324648
R81221 VSS.n680 DVSS 0.00322
R81222 VSS.n9312 VSS.n845 0.00317
R81223 VSS.n9315 VSS.n831 0.00317
R81224 VSS.n9367 VSS.n782 0.00317
R81225 VSS.n9349 VSS.n781 0.00317
R81226 VSS.n9515 VSS.n710 0.00317
R81227 VSS.n9527 VSS.n685 0.00317
R81228 VSS.n9560 VSS.n643 0.00317
R81229 VSS.n9543 VSS.n642 0.00317
R81230 VSS.n1020 VSS.n1014 0.00317
R81231 VSS.n9053 VSS.n1044 0.00317
R81232 VSS.n9020 VSS.n1075 0.00317
R81233 VSS.n9014 VSS.n8985 0.00317
R81234 VSS.n729 VSS.n724 0.00317
R81235 VSS.n9497 VSS.n9496 0.00317
R81236 VSS.n9471 VSS.n604 0.00317
R81237 VSS.n8805 VSS.n1395 0.00317
R81238 VSS.n8791 VSS.n1394 0.00317
R81239 VSS.n8771 VSS.n1100 0.00317
R81240 VSS.n1102 VSS.n1099 0.00317
R81241 VSS.n1150 VSS.n1144 0.00317
R81242 VSS.n1225 VSS.n1165 0.00317
R81243 VSS.n9566 VSS.n566 0.00317
R81244 VSS.n8924 VSS.n565 0.00317
R81245 VSS.n6454 VSS.n6453 0.00317
R81246 VSS.n6451 VSS.n6450 0.00317
R81247 VSS.n6429 VSS.n6428 0.00317
R81248 VSS.n6426 VSS.n3625 0.00317
R81249 VSS.n6407 VSS.n3637 0.00317
R81250 VSS.n6400 VSS.n6341 0.00317
R81251 VSS.n9595 VSS.n447 0.00317
R81252 VSS.n6372 VSS.n446 0.00317
R81253 VSS.n2276 VSS.n2270 0.00315748
R81254 VSS.n2305 VSS.n2148 0.00315748
R81255 VSS.n2422 VSS.n1852 0.00315748
R81256 VSS.n8949 VSS.n1164 0.00315748
R81257 VSS.n1192 VSS.n735 0.00315748
R81258 VSS.n9381 VSS.n698 0.00315748
R81259 VSS.n6373 VSS.n6371 0.00309529
R81260 VSS.n3268 VSS.n3234 0.00309529
R81261 VSS.n2230 VSS.n1715 0.00309529
R81262 VSS.n8925 VSS.n8923 0.00309529
R81263 VSS.n7900 VSS.n1754 0.00309529
R81264 VSS.n9472 VSS.n9470 0.00309529
R81265 VSS.n9544 VSS.n9542 0.00309529
R81266 VSS.n1828 VSS.n1793 0.00309529
R81267 VSS.n8252 VSS.n1791 0.00305
R81268 VSS.n8243 VSS.n8242 0.00305
R81269 VSS.n8224 VSS.n8223 0.00305
R81270 VSS.n8194 VSS.n8193 0.00305
R81271 VSS.n7897 VSS.n1752 0.00305
R81272 VSS.n7931 VSS.n2138 0.00305
R81273 VSS.n8110 VSS.n2031 0.00305
R81274 VSS.n8159 VSS.n8149 0.00305
R81275 VSS.n2247 VSS.n1713 0.00305
R81276 VSS.n2269 VSS.n2268 0.00305
R81277 VSS.n8088 VSS.n7999 0.00305
R81278 VSS.n8635 VSS.n1519 0.00305
R81279 VSS.n6552 VSS.n3232 0.00305
R81280 VSS.n6539 VSS.n3328 0.00305
R81281 VSS.n6526 VSS.n3377 0.00305
R81282 VSS.n6501 VSS.n3451 0.00305
R81283 VSS.n8022 VSS.n1451 0.00303521
R81284 VSS.n8018 VSS.n1484 0.00303521
R81285 VSS.n8858 VSS.n8857 0.00298032
R81286 VSS.n8848 VSS.n1318 0.00298032
R81287 VSS.n8411 VSS.n1662 0.00298032
R81288 VSS.n8564 VSS.n1563 0.00298032
R81289 VSS.n9885 VSS.n33 0.00296479
R81290 VSS.n9858 VSS.n82 0.00296479
R81291 VSS.n9843 VSS.n113 0.00296479
R81292 VSS.n9826 VSS.n146 0.00296479
R81293 VSS.n7286 VSS.n7282 0.00287857
R81294 VSS.n7288 VSS.n7287 0.00287857
R81295 VSS.n9511 VSS.n9510 0.00286
R81296 VSS.n9509 VSS.n9508 0.00286
R81297 VSS.n1142 VSS.n718 0.00286
R81298 VSS.n9540 DVSS 0.00282
R81299 VSS.n2318 VSS.n2163 0.00280315
R81300 VSS.n2409 VSS.n1847 0.00280315
R81301 VSS.n1179 VSS.n751 0.00280315
R81302 VSS.n9394 VSS.n694 0.00280315
R81303 DVSS VSS.n6367 0.00278
R81304 VSS.n5172 VSS.n5171 0.00275352
R81305 VSS.n8257 VSS.n1792 0.00275
R81306 VSS.n1871 VSS.n1864 0.00275
R81307 VSS.n8228 VSS.n1885 0.00275
R81308 VSS.n8198 VSS.n1954 0.00275
R81309 VSS.n7912 VSS.n1753 0.00275
R81310 VSS.n2167 VSS.n2142 0.00275
R81311 VSS.n8104 VSS.n8103 0.00275
R81312 VSS.n8136 VSS.n1980 0.00275
R81313 VSS.n2243 VSS.n1714 0.00275
R81314 VSS.n2260 VSS.n2174 0.00275
R81315 VSS.n7956 VSS.n2089 0.00275
R81316 VSS.n8609 VSS.n1523 0.00275
R81317 VSS.n8496 VSS.n1323 0.00275
R81318 VSS.n1294 VSS.n1284 0.00275
R81319 VSS.n8905 VSS.n1276 0.00275
R81320 VSS.n8885 VSS.n540 0.00275
R81321 VSS.n2996 VSS.n2973 0.00275
R81322 VSS.n6714 VSS.n3081 0.00275
R81323 VSS.n6694 VSS.n3105 0.00275
R81324 VSS.n6674 VSS.n502 0.00275
R81325 VSS.n329 VSS.n309 0.00275
R81326 VSS.n9644 VSS.n363 0.00275
R81327 VSS.n9626 VSS.n387 0.00275
R81328 VSS.n425 VSS.n413 0.00275
R81329 VSS.n5557 VSS.n288 0.00275
R81330 VSS.n5522 VSS.n5392 0.00275
R81331 VSS.n5503 VSS.n5413 0.00275
R81332 VSS.n5482 VSS.n5437 0.00275
R81333 VSS.n6557 VSS.n3233 0.00275
R81334 VSS.n6543 VSS.n3316 0.00275
R81335 VSS.n6530 VSS.n3390 0.00275
R81336 VSS.n6505 VSS.n3464 0.00275
R81337 VSS.n9697 VSS.n9696 0.00275
R81338 VSS.n9741 VSS.n227 0.00275
R81339 VSS.n9779 VSS.n9778 0.00275
R81340 VSS.n9791 VSS.n178 0.00275
R81341 VSS.n9277 VSS.n9276 0.0027
R81342 VSS.n1012 VSS.n862 0.0027
R81343 VSS.n8734 VSS.n8732 0.0027
R81344 VSS.n4720 VSS.n4595 0.0026831
R81345 VSS.n4705 VSS.n4623 0.0026831
R81346 VSS.n5233 VSS.n4346 0.0026831
R81347 VSS.n5206 VSS.n4386 0.0026831
R81348 VSS.n9309 VSS.n9287 0.00263
R81349 VSS.n9309 VSS.n9298 0.00263
R81350 VSS.n9363 VSS.n795 0.00263
R81351 VSS.n9363 VSS.n9352 0.00263
R81352 VSS.n9524 VSS.n9522 0.00263
R81353 VSS.n9524 VSS.n9523 0.00263
R81354 VSS.n9557 VSS.n655 0.00263
R81355 VSS.n9557 VSS.n9546 0.00263
R81356 VSS.n9056 VSS.n9055 0.00263
R81357 VSS.n9055 VSS.n9054 0.00263
R81358 VSS.n9017 VSS.n9016 0.00263
R81359 VSS.n9016 VSS.n8972 0.00263
R81360 VSS.n9500 VSS.n9499 0.00263
R81361 VSS.n9499 VSS.n742 0.00263
R81362 VSS.n9483 VSS.n616 0.00263
R81363 VSS.n9484 VSS.n9483 0.00263
R81364 VSS.n8803 VSS.n1407 0.00263
R81365 VSS.n8803 VSS.n8794 0.00263
R81366 VSS.n8769 VSS.n1101 0.00263
R81367 VSS.n8767 VSS.n1101 0.00263
R81368 VSS.n8951 VSS.n8950 0.00263
R81369 VSS.n8950 VSS.n1152 0.00263
R81370 VSS.n8936 VSS.n578 0.00263
R81371 VSS.n8937 VSS.n8936 0.00263
R81372 VSS.n3562 VSS.n3526 0.00263
R81373 VSS.n3563 VSS.n3562 0.00263
R81374 VSS.n3622 VSS.n3599 0.00263
R81375 VSS.n3623 VSS.n3622 0.00263
R81376 VSS.n6404 VSS.n6403 0.00263
R81377 VSS.n6403 VSS.n3642 0.00263
R81378 VSS.n6384 VSS.n459 0.00263
R81379 VSS.n6385 VSS.n6384 0.00263
R81380 VSS.n8033 VSS.n1137 0.00262598
R81381 VSS.n8026 VSS.n1406 0.00262598
R81382 VSS.n8011 VSS.n1534 0.00262598
R81383 VSS.n8008 VSS.n2125 0.00262598
R81384 VSS.n8812 VSS.n1378 0.00255714
R81385 VSS.n2948 VSS.n2940 0.00255714
R81386 VSS.n4182 VSS.n4170 0.00255714
R81387 VSS.n4253 VSS.n4245 0.00255714
R81388 VSS.n4872 VSS.n4854 0.00255714
R81389 VSS.n9178 VSS.n9177 0.00254
R81390 VSS.n946 VSS.n937 0.00254
R81391 VSS.n8648 VSS.n8647 0.00254
R81392 VSS.n8254 VSS.n1792 0.00251
R81393 VSS.n1867 VSS.n1864 0.00251
R81394 VSS.n8228 VSS.n1910 0.00251
R81395 VSS.n8198 VSS.n8166 0.00251
R81396 VSS.n7914 VSS.n1753 0.00251
R81397 VSS.n7932 VSS.n2142 0.00251
R81398 VSS.n8103 VSS.n2047 0.00251
R81399 VSS.n2016 VSS.n1980 0.00251
R81400 VSS.n2245 VSS.n1714 0.00251
R81401 VSS.n2177 VSS.n2174 0.00251
R81402 VSS.n2092 VSS.n2089 0.00251
R81403 VSS.n8636 VSS.n1523 0.00251
R81404 VSS.n6554 VSS.n3233 0.00251
R81405 VSS.n6543 VSS.n6542 0.00251
R81406 VSS.n6530 VSS.n6529 0.00251
R81407 VSS.n6505 VSS.n6504 0.00251
R81408 VSS.n8298 VSS.n8287 0.00249286
R81409 VSS.n8327 VSS.n8316 0.00249286
R81410 VSS.n8559 VSS.n1578 0.00249286
R81411 VSS.n8378 VSS.n1664 0.00249286
R81412 VSS.n6964 VSS.n2805 0.00249286
R81413 VSS.n2829 VSS.n2825 0.00249286
R81414 VSS.n2855 VSS.n2851 0.00249286
R81415 VSS.n2889 VSS.n2885 0.00249286
R81416 VSS.n6263 VSS.n3842 0.00249286
R81417 VSS.n6197 VSS.n3944 0.00249286
R81418 VSS.n3979 VSS.n3975 0.00249286
R81419 VSS.n6248 VSS.n6238 0.00249286
R81420 VSS.n5300 VSS.n5293 0.00249286
R81421 VSS.n5641 VSS.n5630 0.00249286
R81422 VSS.n4762 VSS.n4737 0.00249286
R81423 VSS.n4784 VSS.n4779 0.00249286
R81424 VSS.n5245 VSS.n4337 0.00249286
R81425 VSS.n5071 VSS.n5060 0.00249286
R81426 DVSS VSS.n9836 0.00247183
R81427 VSS.n4439 VSS.n4437 0.00247183
R81428 VSS.n9835 DVSS 0.00247183
R81429 VSS.n2289 VSS.n2157 0.00244882
R81430 VSS.n2376 VSS.n1862 0.00244882
R81431 VSS.n1208 VSS.n745 0.00244882
R81432 VSS.n9427 VSS.n708 0.00244882
R81433 VSS.n4225 VSS.n4222 0.00240141
R81434 VSS.n3744 VSS.n3139 0.00240141
R81435 VSS.n5708 VSS.n4021 0.00240141
R81436 VSS.n3751 VSS.n3169 0.00240141
R81437 VSS.n2135 VSS.n1882 0.00238
R81438 VSS.n7946 VSS.n7945 0.00238
R81439 VSS.n7947 VSS.n2130 0.00238
R81440 VSS.n7418 VSS 0.0023
R81441 DVSS VSS.n185 0.0023
R81442 DVSS VSS.n8892 0.0023
R81443 VSS.n1634 VSS.n1617 0.0023
R81444 DVSS VSS.n542 0.0023
R81445 DVSS VSS.n6681 0.0023
R81446 VSS.n6841 VSS.n2924 0.0023
R81447 DVSS VSS.n504 0.0023
R81448 VSS.n9614 DVSS 0.0023
R81449 VSS.n6126 VSS.n4014 0.0023
R81450 DVSS VSS.n9615 0.0023
R81451 VSS.n5491 DVSS 0.0023
R81452 VSS.n5596 VSS.n4262 0.0023
R81453 DVSS VSS.n5492 0.0023
R81454 VSS.n5026 VSS.n4491 0.0023
R81455 DVSS VSS.n180 0.0023
R81456 VSS.n9914 VSS 0.0023
R81457 VSS VSS.n9915 0.0023
R81458 VSS VSS.n7419 0.0023
R81459 VSS.n8254 VSS.n1791 0.00221
R81460 VSS.n8243 VSS.n1867 0.00221
R81461 VSS.n8224 VSS.n1910 0.00221
R81462 VSS.n8194 VSS.n8166 0.00221
R81463 VSS.n7914 VSS.n1752 0.00221
R81464 VSS.n7932 VSS.n7931 0.00221
R81465 VSS.n2047 VSS.n2031 0.00221
R81466 VSS.n8159 VSS.n2016 0.00221
R81467 VSS.n2245 VSS.n1713 0.00221
R81468 VSS.n2269 VSS.n2177 0.00221
R81469 VSS.n8088 VSS.n2092 0.00221
R81470 VSS.n8636 VSS.n8635 0.00221
R81471 VSS.n6554 VSS.n3232 0.00221
R81472 VSS.n6542 VSS.n3328 0.00221
R81473 VSS.n6529 VSS.n3377 0.00221
R81474 VSS.n6504 VSS.n3451 0.00221
R81475 VSS.n2393 VSS.n1858 0.00209449
R81476 VSS.n9410 VSS.n704 0.00209449
R81477 VSS.n9312 VSS.n9287 0.00209
R81478 VSS.n9298 VSS.n831 0.00209
R81479 VSS.n9367 VSS.n795 0.00209
R81480 VSS.n9352 VSS.n781 0.00209
R81481 VSS.n9522 VSS.n710 0.00209
R81482 VSS.n9523 VSS.n685 0.00209
R81483 VSS.n9560 VSS.n655 0.00209
R81484 VSS.n9546 VSS.n642 0.00209
R81485 VSS.n9056 VSS.n1020 0.00209
R81486 VSS.n9054 VSS.n9053 0.00209
R81487 VSS.n9017 VSS.n1075 0.00209
R81488 VSS.n9014 VSS.n8972 0.00209
R81489 VSS.n9500 VSS.n729 0.00209
R81490 VSS.n9497 VSS.n742 0.00209
R81491 VSS.n9563 VSS.n616 0.00209
R81492 VSS.n9484 VSS.n604 0.00209
R81493 VSS.n8805 VSS.n1407 0.00209
R81494 VSS.n8794 VSS.n1394 0.00209
R81495 VSS.n8769 VSS.n1100 0.00209
R81496 VSS.n8767 VSS.n1099 0.00209
R81497 VSS.n8951 VSS.n1150 0.00209
R81498 VSS.n1165 VSS.n1152 0.00209
R81499 VSS.n9566 VSS.n578 0.00209
R81500 VSS.n8937 VSS.n565 0.00209
R81501 VSS.n6453 VSS.n3526 0.00209
R81502 VSS.n6451 VSS.n3563 0.00209
R81503 VSS.n6428 VSS.n3599 0.00209
R81504 VSS.n6426 VSS.n3623 0.00209
R81505 VSS.n6404 VSS.n3637 0.00209
R81506 VSS.n6400 VSS.n3642 0.00209
R81507 VSS.n9595 VSS.n459 0.00209
R81508 VSS.n6385 VSS.n446 0.00209
R81509 VSS.n9253 VSS.n887 0.002
R81510 VSS.n981 VSS.n975 0.002
R81511 VSS.n8710 VSS.n1464 0.002
R81512 VSS.n6615 VSS.n3136 0.002
R81513 VSS.n5671 VSS.n5670 0.00197887
R81514 VSS.n3745 VSS.n3159 0.00197887
R81515 VSS.n5673 VSS.n4242 0.00197887
R81516 VSS.n3750 VSS.n3189 0.00197887
R81517 VSS.n8268 VSS.n8257 0.00197
R81518 VSS.n1871 VSS.n1865 0.00197
R81519 VSS.n8231 VSS.n1885 0.00197
R81520 VSS.n8201 VSS.n1954 0.00197
R81521 VSS.n7912 VSS.n7911 0.00197
R81522 VSS.n2168 VSS.n2167 0.00197
R81523 VSS.n8104 VSS.n2035 0.00197
R81524 VSS.n8136 VSS.n1979 0.00197
R81525 VSS.n2243 VSS.n2242 0.00197
R81526 VSS.n2260 VSS.n2175 0.00197
R81527 VSS.n7956 VSS.n2091 0.00197
R81528 VSS.n8633 VSS.n8609 0.00197
R81529 VSS.n6568 VSS.n6557 0.00197
R81530 VSS.n3316 VSS.n3315 0.00197
R81531 VSS.n3390 VSS.n3389 0.00197
R81532 VSS.n3464 VSS.n3463 0.00197
R81533 DVSS VSS.n9467 0.00196
R81534 VSS.n7949 VSS.n2129 0.00194
R81535 VSS.n7943 VSS.n7942 0.00194
R81536 VSS.n1881 VSS.n1878 0.00194
R81537 VSS.n8237 VSS.n8236 0.00194
R81538 VSS.n7941 VSS.n1879 0.00194
R81539 VSS.n9563 DVSS 0.00194
R81540 VSS.n7951 VSS.n7950 0.00194
R81541 VSS.n9468 DVSS 0.00188
R81542 VSS.n9224 VSS.n9223 0.00188
R81543 VSS.n9150 VSS.n9119 0.00188
R81544 VSS.n8687 VSS.n8686 0.00188
R81545 VSS.n6478 VSS.n3165 0.00188
R81546 VSS.n2392 VSS.n1843 0.00174016
R81547 VSS.n9411 VSS.n690 0.00174016
R81548 VSS.n9488 DVSS 0.00173
R81549 VSS.n9487 DVSS 0.00173
R81550 VSS.n8645 VSS.n1518 0.0017
R81551 VSS.n8144 VSS.n945 0.0017
R81552 VSS.n9175 VSS.n940 0.0017
R81553 VSS.n9174 VSS.n9173 0.0017
R81554 VSS.n9172 VSS.n943 0.0017
R81555 VSS.n8644 VSS.n942 0.0017
R81556 VSS.n9913 VSS 0.0017
R81557 VSS.n8573 VSS.n1455 0.00155634
R81558 VSS.n1550 VSS.n1488 0.00155634
R81559 VSS.n9315 VSS.n9314 0.00155
R81560 VSS.n9349 VSS.n780 0.00155
R81561 VSS.n9527 VSS.n9526 0.00155
R81562 VSS.n9543 VSS.n641 0.00155
R81563 VSS.n9050 VSS.n1044 0.00155
R81564 VSS.n9011 VSS.n8985 0.00155
R81565 VSS.n9496 VSS.n755 0.00155
R81566 VSS.n9471 VSS.n603 0.00155
R81567 VSS.n8791 VSS.n1393 0.00155
R81568 VSS.n8962 VSS.n1102 0.00155
R81569 VSS.n8948 VSS.n1225 0.00155
R81570 VSS.n8924 VSS.n564 0.00155
R81571 VSS.n6450 VSS.n3550 0.00155
R81572 VSS.n6424 VSS.n3625 0.00155
R81573 VSS.n6396 VSS.n6341 0.00155
R81574 VSS.n6372 VSS.n445 0.00155
R81575 VSS.n5168 VSS.n4454 0.00148592
R81576 VSS.n2135 VSS.n2134 0.00146
R81577 VSS.n7946 VSS.n2136 0.00146
R81578 VSS.n7948 VSS.n7947 0.00146
R81579 VSS.n8730 VSS.n1011 0.00146
R81580 VSS.n9065 VSS.n9064 0.00146
R81581 VSS.n9274 VSS.n861 0.00146
R81582 VSS.n9250 VSS.n9230 0.00146
R81583 VSS.n9273 VSS.n860 0.00146
R81584 VSS.n9115 VSS.n9114 0.00146
R81585 VSS.n9066 VSS.n1008 0.00146
R81586 VSS.n8693 VSS.n1462 0.00146
R81587 VSS.n8729 VSS.n1433 0.00146
R81588 VSS.n3161 VSS.n3149 0.00146
R81589 VSS.n8271 VSS.n1805 0.00143
R81590 VSS.n8245 VSS.n1851 0.00143
R81591 VSS.n8232 VSS.n1880 0.00143
R81592 VSS.n8202 VSS.n1949 0.00143
R81593 VSS.n8274 VSS.n1766 0.00143
R81594 VSS.n7929 VSS.n7928 0.00143
R81595 VSS.n8101 VSS.n8098 0.00143
R81596 VSS.n8163 VSS.n1994 0.00143
R81597 VSS.n8277 VSS.n1727 0.00143
R81598 VSS.n2258 VSS.n2176 0.00143
R81599 VSS.n7954 VSS.n2090 0.00143
R81600 VSS.n1543 VSS.n1541 0.00143
R81601 VSS.n6572 VSS.n3247 0.00143
R81602 VSS.n6545 VSS.n3291 0.00143
R81603 VSS.n6532 VSS.n3353 0.00143
R81604 VSS.n6507 VSS.n3427 0.00143
R81605 VSS.n8816 VSS.n1369 0.0014
R81606 VSS.n3014 VSS.n2941 0.0014
R81607 VSS.n5723 VSS.n4172 0.0014
R81608 VSS.n5589 VSS.n4246 0.0014
R81609 VSS.n5018 VSS.n4975 0.0014
R81610 VSS.n8584 VSS.n1119 0.00138583
R81611 VSS.n2288 VSS.n2152 0.00138583
R81612 VSS.n2377 VSS.n1840 0.00138583
R81613 VSS.n8590 VSS.n1419 0.00138583
R81614 VSS.n8604 VSS.n1539 0.00138583
R81615 VSS.n8087 VSS.n8086 0.00138583
R81616 VSS.n1209 VSS.n739 0.00138583
R81617 VSS.n9426 VSS.n687 0.00138583
R81618 VSS.n4460 VSS.n4449 0.00134507
R81619 VSS.n8053 VSS.n1453 0.00134507
R81620 VSS.n5115 VSS.n4425 0.00134507
R81621 VSS.n8061 VSS.n1486 0.00134507
R81622 DVSS VSS.n6388 0.00134
R81623 DVSS VSS.n8940 0.00134
R81624 VSS.n9218 VSS.n901 0.00134
R81625 VSS.n9155 VSS.n961 0.00134
R81626 VSS.n1495 VSS.n1477 0.00134
R81627 DVSS VSS.n566 0.00134
R81628 VSS.n6481 VSS.n6480 0.00134
R81629 DVSS VSS.n447 0.00134
R81630 VSS.n9177 VSS.n9176 0.0013
R81631 VSS.n8143 VSS.n937 0.0013
R81632 VSS.n8647 VSS.n8646 0.0013
R81633 VSS.n8960 VSS.n8959 0.00122
R81634 VSS.n8999 VSS.n721 0.00122
R81635 VSS.n9348 VSS.n716 0.00122
R81636 VSS.n9347 VSS.n715 0.00122
R81637 VSS.n9000 VSS.n723 0.00122
R81638 VSS.n8961 VSS.n1139 0.00122
R81639 VSS.n8043 VSS.n8040 0.00120866
R81640 VSS.n8048 VSS.n1408 0.00120866
R81641 VSS.n8067 VSS.n1536 0.00120866
R81642 VSS.n8072 VSS.n8001 0.00120866
R81643 VSS.n5179 VSS.n4429 0.00120422
R81644 VSS.n8538 VSS.n1625 0.00114286
R81645 VSS.n2923 VSS.n2919 0.00114286
R81646 VSS.n4013 VSS.n4009 0.00114286
R81647 VSS.n5663 VSS.n4271 0.00114286
R81648 VSS.n5084 VSS.n4499 0.00114286
R81649 VSS.n9276 VSS.n9275 0.00114
R81650 VSS.n1010 VSS.n862 0.00114
R81651 VSS.n8732 VSS.n8731 0.00114
R81652 VSS.n3737 VSS.n3142 0.0011338
R81653 VSS.n3766 VSS.n3172 0.0011338
R81654 VSS.n6368 DVSS 0.00106
R81655 VSS.n2319 VSS.n2145 0.0010315
R81656 VSS.n2408 VSS.n1855 0.0010315
R81657 VSS.n1178 VSS.n732 0.0010315
R81658 VSS.n9395 VSS.n701 0.0010315
R81659 DVSS VSS.n9539 0.00102
R81660 VSS.n9510 VSS.n717 0.00098
R81661 VSS.n9509 VSS.n719 0.00098
R81662 VSS.n1141 VSS.n718 0.00098
R81663 VSS.n1373 VSS.n1363 0.000922535
R81664 VSS.n8394 VSS.n1622 0.000922535
R81665 VSS.n9256 VSS.n873 0.00092
R81666 VSS.n9109 VSS.n982 0.00092
R81667 VSS.n8712 VSS.n1444 0.00092
R81668 VSS.n6474 VSS.n3135 0.00092
R81669 VSS.n8851 VSS.n1291 0.000854331
R81670 VSS.n8844 VSS.n8843 0.000854331
R81671 VSS.n8392 VSS.n1658 0.000854331
R81672 VSS.n8560 VSS.n1559 0.000854331
R81673 VSS.n9221 VSS.n9197 0.0008
R81674 VSS.n9156 VSS.n956 0.0008
R81675 VSS.n8684 VSS.n8667 0.0008
R81676 VSS.n6609 VSS.n3179 0.0008
R81677 VSS.n3729 VSS.n3152 0.000711268
R81678 VSS.n6789 VSS.n2945 0.000711268
R81679 VSS.n3781 VSS.n3182 0.000711268
R81680 VSS.n6791 VSS.n2927 0.000711268
R81681 DVSS VSS.n129 0.000687793
R81682 VSS.n9538 DVSS 0.00068
R81683 DVSS VSS.n643 0.00068
R81684 VSS.n2304 VSS.n2160 0.000677165
R81685 VSS.n2423 VSS.n1850 0.000677165
R81686 VSS.n1193 VSS.n748 0.000677165
R81687 VSS.n9380 VSS.n697 0.000677165
R81688 VSS VSS.n7408 0.000671429
R81689 DVSS VSS.n9790 0.000671429
R81690 VSS.n8891 DVSS 0.000671429
R81691 VSS.n6680 DVSS 0.000671429
R81692 VSS.n9613 DVSS 0.000671429
R81693 VSS.n5490 DVSS 0.000671429
R81694 VSS.n9913 VSS 0.000671429
R81695 VSS.n9539 DVSS 0.00062
R81696 DVSS VSS.n6368 0.00058
R81697 DVSS VSS.n8920 0.00058
C0 DVSS VDD 50.9753f
C1 DVDD VDD 48.1675f
C2 DVSS ASIG5V 0.485981p
C3 DVDD ASIG5V 0.626156p
C4 ASIG5V VDD 21.911001f
C5 DVSS DVDD 1.55543p
C6 VDD VSS 56.043198f
C7 ASIG5V VSS 0.258722p
C8 DVDD VSS 0.754874p
C9 DVSS VSS 0.389892p
C10 VDD.n0 VSS 0.618992f
C11 VDD.n1 VSS 0.902595f
C12 VDD.n2 VSS 12.7524f
C13 VDD.n3 VSS 0.081789f
C14 VDD.n4 VSS 0.618992f
C15 VDD.n5 VSS 26.8072f
C16 VDD.n6 VSS 0.021107f
C17 VDD.n7 VSS 0.246589f
C18 VDD.n8 VSS 0.902595f
C19 VDD.n9 VSS 0.101025f
C20 VDD.n10 VSS 1.13549f
C21 VDD.n11 VSS 1.13549f
C22 VDD.n12 VSS 0.101122f
C23 VDD.n13 VSS 0.081789f
C24 VDD.n14 VSS 12.752299f
C25 VDD.n15 VSS 27.137402f
C26 VDD.n16 VSS 15.5483f
C27 VDD.n17 VSS 0.246589f
C28 ASIG5V.n0 VSS 0.701152f
C29 ASIG5V.n1 VSS 0.470002f
C30 ASIG5V.n2 VSS 0.045974f
C31 ASIG5V.n3 VSS 0.076709f
C32 ASIG5V.n4 VSS 0.045974f
C33 ASIG5V.n5 VSS 0.076709f
C34 ASIG5V.n6 VSS 0.052746f
C35 ASIG5V.n7 VSS 0.052746f
C36 ASIG5V.n8 VSS 0.045974f
C37 ASIG5V.n9 VSS 0.045974f
C38 ASIG5V.n10 VSS 1.0941f
C39 ASIG5V.n52 VSS 0.970825f
C40 ASIG5V.n53 VSS 0.056945f
C41 ASIG5V.n54 VSS 0.0621f
C42 ASIG5V.n55 VSS 0.036092f
C43 ASIG5V.n56 VSS 0.123278f
C44 ASIG5V.n98 VSS 0.970825f
C45 ASIG5V.n99 VSS 0.056945f
C46 ASIG5V.n100 VSS 0.056945f
C47 ASIG5V.n101 VSS 0.056945f
C48 ASIG5V.n102 VSS 0.056945f
C49 ASIG5V.n103 VSS 0.056945f
C50 ASIG5V.n104 VSS 0.056945f
C51 ASIG5V.n105 VSS 0.056945f
C52 ASIG5V.n106 VSS 0.056945f
C53 ASIG5V.n107 VSS 0.056945f
C54 ASIG5V.n108 VSS 0.056945f
C55 ASIG5V.n109 VSS 0.056945f
C56 ASIG5V.n110 VSS 0.056945f
C57 ASIG5V.n111 VSS 0.056945f
C58 ASIG5V.n112 VSS 0.056945f
C59 ASIG5V.n113 VSS 0.056945f
C60 ASIG5V.n114 VSS 0.056945f
C61 ASIG5V.n115 VSS 0.056945f
C62 ASIG5V.n116 VSS 0.056945f
C63 ASIG5V.n117 VSS 0.056945f
C64 ASIG5V.n118 VSS 0.056945f
C65 ASIG5V.n119 VSS 0.056945f
C66 ASIG5V.n120 VSS 0.056945f
C67 ASIG5V.n121 VSS 0.056945f
C68 ASIG5V.n122 VSS 0.056945f
C69 ASIG5V.n123 VSS 0.056945f
C70 ASIG5V.n124 VSS 0.056945f
C71 ASIG5V.n125 VSS 0.056945f
C72 ASIG5V.n126 VSS 0.056945f
C73 ASIG5V.n127 VSS 0.056945f
C74 ASIG5V.n128 VSS 0.056945f
C75 ASIG5V.n129 VSS 0.056945f
C76 ASIG5V.n130 VSS 0.056945f
C77 ASIG5V.n131 VSS 0.056945f
C78 ASIG5V.n132 VSS 0.056945f
C79 ASIG5V.n133 VSS 0.056945f
C80 ASIG5V.n134 VSS 0.056945f
C81 ASIG5V.n135 VSS 0.056945f
C82 ASIG5V.n136 VSS 0.056945f
C83 ASIG5V.n137 VSS 0.056945f
C84 ASIG5V.n138 VSS 0.056945f
C85 ASIG5V.n139 VSS 0.056945f
C86 ASIG5V.n140 VSS 0.056945f
C87 ASIG5V.n141 VSS 0.056945f
C88 ASIG5V.n142 VSS 0.056945f
C89 ASIG5V.n143 VSS 0.056945f
C90 ASIG5V.n144 VSS 0.056945f
C91 ASIG5V.n145 VSS 0.056945f
C92 ASIG5V.n146 VSS 0.056945f
C93 ASIG5V.n147 VSS 0.056945f
C94 ASIG5V.n148 VSS 0.056945f
C95 ASIG5V.n149 VSS 0.056945f
C96 ASIG5V.n150 VSS 0.056945f
C97 ASIG5V.n151 VSS 0.056945f
C98 ASIG5V.n152 VSS 0.056945f
C99 ASIG5V.n153 VSS 0.056945f
C100 ASIG5V.n154 VSS 0.056945f
C101 ASIG5V.n155 VSS 0.056945f
C102 ASIG5V.n156 VSS 0.056945f
C103 ASIG5V.n157 VSS 0.056945f
C104 ASIG5V.n158 VSS 0.056945f
C105 ASIG5V.n159 VSS 0.056945f
C106 ASIG5V.n160 VSS 0.056945f
C107 ASIG5V.n161 VSS 0.072161f
C108 ASIG5V.n162 VSS 0.09726f
C109 ASIG5V.n163 VSS 0.0621f
C110 ASIG5V.n164 VSS 0.108961f
C111 ASIG5V.n165 VSS 0.0621f
C112 ASIG5V.n166 VSS 0.99394f
C113 ASIG5V.n167 VSS 0.0621f
C114 ASIG5V.n168 VSS 0.052133f
C115 ASIG5V.n169 VSS 0.536863f
C116 ASIG5V.n170 VSS 0.09726f
C117 ASIG5V.n171 VSS 0.108961f
C118 ASIG5V.n172 VSS 0.108961f
C119 ASIG5V.n173 VSS 0.832135f
C120 ASIG5V.n215 VSS 0.036092f
C121 ASIG5V.n216 VSS 0.693446f
C122 ASIG5V.n217 VSS 0.045974f
C123 ASIG5V.n218 VSS 0.036092f
C124 ASIG5V.n219 VSS 0.223443f
C125 ASIG5V.n220 VSS 0.056945f
C126 ASIG5V.n221 VSS 0.056945f
C127 ASIG5V.n222 VSS 0.056945f
C128 ASIG5V.n223 VSS 0.056945f
C129 ASIG5V.n224 VSS 0.056945f
C130 ASIG5V.n225 VSS 0.056945f
C131 ASIG5V.n226 VSS 0.056945f
C132 ASIG5V.n227 VSS 0.056945f
C133 ASIG5V.n228 VSS 0.056945f
C134 ASIG5V.n229 VSS 0.056945f
C135 ASIG5V.n230 VSS 0.056945f
C136 ASIG5V.n231 VSS 0.056945f
C137 ASIG5V.n232 VSS 0.056945f
C138 ASIG5V.n233 VSS 0.056945f
C139 ASIG5V.n234 VSS 0.056945f
C140 ASIG5V.n235 VSS 0.056945f
C141 ASIG5V.n236 VSS 0.056945f
C142 ASIG5V.n237 VSS 0.056945f
C143 ASIG5V.n238 VSS 0.056945f
C144 ASIG5V.n239 VSS 0.056945f
C145 ASIG5V.n240 VSS 0.056945f
C146 ASIG5V.n241 VSS 0.056945f
C147 ASIG5V.n242 VSS 0.056945f
C148 ASIG5V.n243 VSS 0.056945f
C149 ASIG5V.n244 VSS 0.056945f
C150 ASIG5V.n245 VSS 0.056945f
C151 ASIG5V.n246 VSS 0.056945f
C152 ASIG5V.n247 VSS 0.056945f
C153 ASIG5V.n248 VSS 0.056945f
C154 ASIG5V.n249 VSS 0.056945f
C155 ASIG5V.n250 VSS 0.056945f
C156 ASIG5V.n251 VSS 0.056945f
C157 ASIG5V.n252 VSS 0.056945f
C158 ASIG5V.n253 VSS 0.056945f
C159 ASIG5V.n254 VSS 0.056945f
C160 ASIG5V.n255 VSS 0.056945f
C161 ASIG5V.n256 VSS 0.056945f
C162 ASIG5V.n257 VSS 0.056945f
C163 ASIG5V.n258 VSS 0.056945f
C164 ASIG5V.n259 VSS 0.056945f
C165 ASIG5V.n260 VSS 0.036092f
C166 ASIG5V.n262 VSS 0.056945f
C167 ASIG5V.n263 VSS 0.056945f
C168 ASIG5V.n264 VSS 0.056945f
C169 ASIG5V.n265 VSS 0.056945f
C170 ASIG5V.n266 VSS 0.056945f
C171 ASIG5V.n267 VSS 0.056945f
C172 ASIG5V.n269 VSS 0.056945f
C173 ASIG5V.n270 VSS 0.056945f
C174 ASIG5V.n271 VSS 0.056945f
C175 ASIG5V.n273 VSS 0.056945f
C176 ASIG5V.n274 VSS 0.056945f
C177 ASIG5V.n275 VSS 0.056945f
C178 ASIG5V.n276 VSS 0.056945f
C179 ASIG5V.n277 VSS 0.056945f
C180 ASIG5V.n278 VSS 0.056945f
C181 ASIG5V.n279 VSS 0.056945f
C182 ASIG5V.n281 VSS 0.056945f
C183 ASIG5V.n282 VSS 0.056945f
C184 ASIG5V.n283 VSS 0.056945f
C185 ASIG5V.n285 VSS 0.056945f
C186 ASIG5V.n286 VSS 0.056945f
C187 ASIG5V.n287 VSS 0.056945f
C188 ASIG5V.n288 VSS 0.056945f
C189 ASIG5V.n289 VSS 0.056945f
C190 ASIG5V.n290 VSS 0.056945f
C191 ASIG5V.n291 VSS 0.056945f
C192 ASIG5V.n293 VSS 0.056945f
C193 ASIG5V.n294 VSS 0.056945f
C194 ASIG5V.n295 VSS 0.056945f
C195 ASIG5V.n297 VSS 0.056945f
C196 ASIG5V.n298 VSS 0.056945f
C197 ASIG5V.n299 VSS 0.056945f
C198 ASIG5V.n300 VSS 0.056945f
C199 ASIG5V.n301 VSS 0.056945f
C200 ASIG5V.n302 VSS 0.056945f
C201 ASIG5V.n303 VSS 0.056945f
C202 ASIG5V.n305 VSS 0.056945f
C203 ASIG5V.n306 VSS 0.056945f
C204 ASIG5V.n307 VSS 0.056945f
C205 ASIG5V.n309 VSS 0.056945f
C206 ASIG5V.n310 VSS 0.056945f
C207 ASIG5V.n311 VSS 0.056945f
C208 ASIG5V.n312 VSS 0.056945f
C209 ASIG5V.n313 VSS 0.056945f
C210 ASIG5V.n314 VSS 0.056945f
C211 ASIG5V.n315 VSS 0.056945f
C212 ASIG5V.n317 VSS 0.056945f
C213 ASIG5V.n318 VSS 0.056945f
C214 ASIG5V.n319 VSS 0.056945f
C215 ASIG5V.n321 VSS 0.056945f
C216 ASIG5V.n322 VSS 0.056945f
C217 ASIG5V.n323 VSS 0.056945f
C218 ASIG5V.n324 VSS 0.056945f
C219 ASIG5V.n325 VSS 0.056945f
C220 ASIG5V.n326 VSS 0.056945f
C221 ASIG5V.n327 VSS 0.056945f
C222 ASIG5V.n329 VSS 0.056945f
C223 ASIG5V.n330 VSS 0.056945f
C224 ASIG5V.n331 VSS 0.056945f
C225 ASIG5V.n333 VSS 0.056945f
C226 ASIG5V.n334 VSS 0.056945f
C227 ASIG5V.n335 VSS 0.056945f
C228 ASIG5V.n336 VSS 0.056945f
C229 ASIG5V.n337 VSS 0.056945f
C230 ASIG5V.n338 VSS 0.056945f
C231 ASIG5V.n339 VSS 0.056945f
C232 ASIG5V.n341 VSS 0.056945f
C233 ASIG5V.n342 VSS 0.056945f
C234 ASIG5V.n343 VSS 0.056945f
C235 ASIG5V.n345 VSS 0.056945f
C236 ASIG5V.n346 VSS 0.056945f
C237 ASIG5V.n347 VSS 0.056945f
C238 ASIG5V.n348 VSS 0.056945f
C239 ASIG5V.n349 VSS 0.056945f
C240 ASIG5V.n350 VSS 0.056945f
C241 ASIG5V.n351 VSS 0.056945f
C242 ASIG5V.n353 VSS 0.056945f
C243 ASIG5V.n354 VSS 0.056945f
C244 ASIG5V.n355 VSS 0.056945f
C245 ASIG5V.n357 VSS 0.056945f
C246 ASIG5V.n358 VSS 0.056945f
C247 ASIG5V.n359 VSS 0.056945f
C248 ASIG5V.n360 VSS 0.056945f
C249 ASIG5V.n361 VSS 0.056945f
C250 ASIG5V.n362 VSS 0.056945f
C251 ASIG5V.n363 VSS 0.056945f
C252 ASIG5V.n365 VSS 0.056945f
C253 ASIG5V.n366 VSS 0.056945f
C254 ASIG5V.n367 VSS 0.056945f
C255 ASIG5V.n369 VSS 0.056945f
C256 ASIG5V.n370 VSS 0.056945f
C257 ASIG5V.n371 VSS 0.056945f
C258 ASIG5V.n372 VSS 0.056945f
C259 ASIG5V.n373 VSS 0.056945f
C260 ASIG5V.n374 VSS 0.056945f
C261 ASIG5V.n375 VSS 0.056945f
C262 ASIG5V.n377 VSS 0.056945f
C263 ASIG5V.n378 VSS 0.056945f
C264 ASIG5V.n379 VSS 0.056945f
C265 ASIG5V.n381 VSS 0.056945f
C266 ASIG5V.n382 VSS 0.056945f
C267 ASIG5V.n383 VSS 0.056945f
C268 ASIG5V.n384 VSS 0.056945f
C269 ASIG5V.n385 VSS 0.056945f
C270 ASIG5V.n386 VSS 0.056945f
C271 ASIG5V.n387 VSS 0.056945f
C272 ASIG5V.n389 VSS 0.056945f
C273 ASIG5V.n390 VSS 0.056945f
C274 ASIG5V.n391 VSS 0.056945f
C275 ASIG5V.n393 VSS 0.056945f
C276 ASIG5V.n394 VSS 0.056945f
C277 ASIG5V.n395 VSS 0.056945f
C278 ASIG5V.n396 VSS 0.056945f
C279 ASIG5V.n397 VSS 0.056945f
C280 ASIG5V.n398 VSS 0.056945f
C281 ASIG5V.n399 VSS 0.056945f
C282 ASIG5V.n401 VSS 0.056945f
C283 ASIG5V.n402 VSS 0.056945f
C284 ASIG5V.n403 VSS 0.056945f
C285 ASIG5V.n405 VSS 0.056945f
C286 ASIG5V.n406 VSS 0.056945f
C287 ASIG5V.n407 VSS 0.056945f
C288 ASIG5V.n408 VSS 0.056945f
C289 ASIG5V.n409 VSS 0.056945f
C290 ASIG5V.n410 VSS 0.056945f
C291 ASIG5V.n411 VSS 0.056945f
C292 ASIG5V.n413 VSS 0.056945f
C293 ASIG5V.n414 VSS 0.056945f
C294 ASIG5V.n415 VSS 0.056945f
C295 ASIG5V.n417 VSS 0.056945f
C296 ASIG5V.n418 VSS 0.056945f
C297 ASIG5V.n419 VSS 0.056945f
C298 ASIG5V.n420 VSS 0.056945f
C299 ASIG5V.n421 VSS 0.056945f
C300 ASIG5V.n422 VSS 0.056945f
C301 ASIG5V.n423 VSS 0.056945f
C302 ASIG5V.n425 VSS 0.056945f
C303 ASIG5V.n426 VSS 0.056945f
C304 ASIG5V.n427 VSS 0.056945f
C305 ASIG5V.n429 VSS 0.056945f
C306 ASIG5V.n430 VSS 0.056945f
C307 ASIG5V.n431 VSS 0.056945f
C308 ASIG5V.n432 VSS 0.056945f
C309 ASIG5V.n433 VSS 0.056945f
C310 ASIG5V.n434 VSS 0.056945f
C311 ASIG5V.n435 VSS 0.056945f
C312 ASIG5V.n437 VSS 0.056945f
C313 ASIG5V.n438 VSS 0.056945f
C314 ASIG5V.n439 VSS 0.056945f
C315 ASIG5V.n441 VSS 0.056945f
C316 ASIG5V.n442 VSS 0.056945f
C317 ASIG5V.n443 VSS 0.056945f
C318 ASIG5V.n444 VSS 0.056945f
C319 ASIG5V.n445 VSS 0.056945f
C320 ASIG5V.n446 VSS 0.056945f
C321 ASIG5V.n447 VSS 0.056945f
C322 ASIG5V.n449 VSS 0.056945f
C323 ASIG5V.n450 VSS 0.056945f
C324 ASIG5V.n451 VSS 0.056945f
C325 ASIG5V.n453 VSS 0.056945f
C326 ASIG5V.n454 VSS 0.056945f
C327 ASIG5V.n455 VSS 0.056945f
C328 ASIG5V.n456 VSS 0.056945f
C329 ASIG5V.n457 VSS 0.056945f
C330 ASIG5V.n458 VSS 0.056945f
C331 ASIG5V.n459 VSS 0.056945f
C332 ASIG5V.n461 VSS 0.056945f
C333 ASIG5V.n462 VSS 0.056945f
C334 ASIG5V.n463 VSS 0.056945f
C335 ASIG5V.n465 VSS 0.056945f
C336 ASIG5V.n466 VSS 0.056945f
C337 ASIG5V.n467 VSS 0.056945f
C338 ASIG5V.n468 VSS 0.056945f
C339 ASIG5V.n469 VSS 0.056945f
C340 ASIG5V.n470 VSS 0.056945f
C341 ASIG5V.n471 VSS 0.056945f
C342 ASIG5V.n473 VSS 0.056945f
C343 ASIG5V.n474 VSS 0.056945f
C344 ASIG5V.n475 VSS 0.056945f
C345 ASIG5V.n477 VSS 0.056945f
C346 ASIG5V.n478 VSS 0.056945f
C347 ASIG5V.n479 VSS 0.056945f
C348 ASIG5V.n480 VSS 0.056945f
C349 ASIG5V.n481 VSS 0.056945f
C350 ASIG5V.n482 VSS 0.056945f
C351 ASIG5V.n483 VSS 0.056945f
C352 ASIG5V.n485 VSS 0.056945f
C353 ASIG5V.n486 VSS 0.056945f
C354 ASIG5V.n487 VSS 0.056945f
C355 ASIG5V.n489 VSS 0.056945f
C356 ASIG5V.n490 VSS 0.056945f
C357 ASIG5V.n491 VSS 0.056945f
C358 ASIG5V.n492 VSS 0.056945f
C359 ASIG5V.n493 VSS 0.056945f
C360 ASIG5V.n494 VSS 0.056945f
C361 ASIG5V.n495 VSS 0.056945f
C362 ASIG5V.n497 VSS 0.056945f
C363 ASIG5V.n498 VSS 0.056945f
C364 ASIG5V.n499 VSS 0.056945f
C365 ASIG5V.n501 VSS 0.056945f
C366 ASIG5V.n502 VSS 0.056945f
C367 ASIG5V.n503 VSS 0.056945f
C368 ASIG5V.n504 VSS 0.056945f
C369 ASIG5V.n505 VSS 0.047415f
C370 ASIG5V.n506 VSS 0.066995f
C371 ASIG5V.n507 VSS 0.076709f
C372 ASIG5V.n508 VSS 0.955415f
C373 ASIG5V.n509 VSS 0.066995f
C374 ASIG5V.n510 VSS 0.046943f
C375 ASIG5V.n511 VSS 0.05375f
C376 ASIG5V.n512 VSS 0.05375f
C377 ASIG5V.n513 VSS 0.955415f
C378 ASIG5V.n514 VSS 0.076709f
C379 ASIG5V.n515 VSS 0.05429f
C380 ASIG5V.n516 VSS 0.05429f
C381 ASIG5V.n517 VSS 0.045974f
C382 ASIG5V.n518 VSS 0.076709f
C383 ASIG5V.n519 VSS 0.047268f
C384 ASIG5V.n520 VSS 1.0941f
C385 ASIG5V.n521 VSS 0.639512f
C386 ASIG5V.n522 VSS 0.0621f
C387 ASIG5V.n523 VSS 0.0621f
C388 ASIG5V.n524 VSS 0.052133f
C389 ASIG5V.n525 VSS 0.09726f
C390 ASIG5V.n526 VSS 0.108961f
C391 ASIG5V.n527 VSS 0.108961f
C392 ASIG5V.n528 VSS 0.639512f
C393 ASIG5V.n570 VSS 0.036092f
C394 ASIG5V.n571 VSS 0.500822f
C395 ASIG5V.n572 VSS 0.045974f
C396 ASIG5V.n573 VSS 0.036092f
C397 ASIG5V.n574 VSS 0.056945f
C398 ASIG5V.n575 VSS 0.056945f
C399 ASIG5V.n576 VSS 0.056945f
C400 ASIG5V.n577 VSS 0.056945f
C401 ASIG5V.n578 VSS 0.056945f
C402 ASIG5V.n579 VSS 0.056945f
C403 ASIG5V.n580 VSS 0.056945f
C404 ASIG5V.n581 VSS 0.056945f
C405 ASIG5V.n582 VSS 0.056945f
C406 ASIG5V.n583 VSS 0.056945f
C407 ASIG5V.n584 VSS 0.056945f
C408 ASIG5V.n585 VSS 0.056945f
C409 ASIG5V.n586 VSS 0.056945f
C410 ASIG5V.n587 VSS 0.056945f
C411 ASIG5V.n588 VSS 0.056945f
C412 ASIG5V.n589 VSS 0.056945f
C413 ASIG5V.n590 VSS 0.056945f
C414 ASIG5V.n591 VSS 0.056945f
C415 ASIG5V.n592 VSS 0.056945f
C416 ASIG5V.n593 VSS 0.056945f
C417 ASIG5V.n594 VSS 0.056945f
C418 ASIG5V.n595 VSS 0.056945f
C419 ASIG5V.n596 VSS 0.056945f
C420 ASIG5V.n597 VSS 0.056945f
C421 ASIG5V.n598 VSS 0.056945f
C422 ASIG5V.n599 VSS 0.056945f
C423 ASIG5V.n600 VSS 0.056945f
C424 ASIG5V.n601 VSS 0.056945f
C425 ASIG5V.n602 VSS 0.056945f
C426 ASIG5V.n603 VSS 0.056945f
C427 ASIG5V.n604 VSS 0.056945f
C428 ASIG5V.n605 VSS 0.056945f
C429 ASIG5V.n606 VSS 0.056945f
C430 ASIG5V.n607 VSS 0.056945f
C431 ASIG5V.n608 VSS 0.056945f
C432 ASIG5V.n609 VSS 0.056945f
C433 ASIG5V.n610 VSS 0.056945f
C434 ASIG5V.n611 VSS 0.056945f
C435 ASIG5V.n612 VSS 0.056945f
C436 ASIG5V.n613 VSS 0.056945f
C437 ASIG5V.n614 VSS 0.036092f
C438 ASIG5V.n616 VSS 0.056945f
C439 ASIG5V.n617 VSS 0.056945f
C440 ASIG5V.n618 VSS 0.056945f
C441 ASIG5V.n619 VSS 0.056945f
C442 ASIG5V.n620 VSS 0.056945f
C443 ASIG5V.n621 VSS 0.056945f
C444 ASIG5V.n623 VSS 0.056945f
C445 ASIG5V.n624 VSS 0.056945f
C446 ASIG5V.n625 VSS 0.056945f
C447 ASIG5V.n627 VSS 0.056945f
C448 ASIG5V.n628 VSS 0.056945f
C449 ASIG5V.n629 VSS 0.056945f
C450 ASIG5V.n630 VSS 0.056945f
C451 ASIG5V.n631 VSS 0.056945f
C452 ASIG5V.n632 VSS 0.056945f
C453 ASIG5V.n633 VSS 0.056945f
C454 ASIG5V.n635 VSS 0.056945f
C455 ASIG5V.n636 VSS 0.056945f
C456 ASIG5V.n637 VSS 0.056945f
C457 ASIG5V.n639 VSS 0.056945f
C458 ASIG5V.n640 VSS 0.056945f
C459 ASIG5V.n641 VSS 0.056945f
C460 ASIG5V.n642 VSS 0.056945f
C461 ASIG5V.n643 VSS 0.056945f
C462 ASIG5V.n644 VSS 0.056945f
C463 ASIG5V.n645 VSS 0.056945f
C464 ASIG5V.n647 VSS 0.056945f
C465 ASIG5V.n648 VSS 0.056945f
C466 ASIG5V.n649 VSS 0.056945f
C467 ASIG5V.n651 VSS 0.056945f
C468 ASIG5V.n652 VSS 0.056945f
C469 ASIG5V.n653 VSS 0.056945f
C470 ASIG5V.n654 VSS 0.056945f
C471 ASIG5V.n655 VSS 0.056945f
C472 ASIG5V.n656 VSS 0.056945f
C473 ASIG5V.n657 VSS 0.056945f
C474 ASIG5V.n659 VSS 0.056945f
C475 ASIG5V.n660 VSS 0.056945f
C476 ASIG5V.n661 VSS 0.056945f
C477 ASIG5V.n663 VSS 0.056945f
C478 ASIG5V.n664 VSS 0.056945f
C479 ASIG5V.n665 VSS 0.056945f
C480 ASIG5V.n666 VSS 0.056945f
C481 ASIG5V.n667 VSS 0.056945f
C482 ASIG5V.n668 VSS 0.056945f
C483 ASIG5V.n669 VSS 0.056945f
C484 ASIG5V.n671 VSS 0.056945f
C485 ASIG5V.n672 VSS 0.056945f
C486 ASIG5V.n673 VSS 0.056945f
C487 ASIG5V.n675 VSS 0.056945f
C488 ASIG5V.n676 VSS 0.056945f
C489 ASIG5V.n677 VSS 0.056945f
C490 ASIG5V.n678 VSS 0.056945f
C491 ASIG5V.n679 VSS 0.056945f
C492 ASIG5V.n680 VSS 0.056945f
C493 ASIG5V.n681 VSS 0.056945f
C494 ASIG5V.n683 VSS 0.056945f
C495 ASIG5V.n684 VSS 0.056945f
C496 ASIG5V.n685 VSS 0.056945f
C497 ASIG5V.n687 VSS 0.056945f
C498 ASIG5V.n688 VSS 0.056945f
C499 ASIG5V.n689 VSS 0.056945f
C500 ASIG5V.n690 VSS 0.056945f
C501 ASIG5V.n691 VSS 0.056945f
C502 ASIG5V.n692 VSS 0.056945f
C503 ASIG5V.n693 VSS 0.056945f
C504 ASIG5V.n695 VSS 0.056945f
C505 ASIG5V.n696 VSS 0.056945f
C506 ASIG5V.n697 VSS 0.056945f
C507 ASIG5V.n699 VSS 0.056945f
C508 ASIG5V.n700 VSS 0.056945f
C509 ASIG5V.n701 VSS 0.056945f
C510 ASIG5V.n702 VSS 0.056945f
C511 ASIG5V.n703 VSS 0.056945f
C512 ASIG5V.n704 VSS 0.056945f
C513 ASIG5V.n705 VSS 0.056945f
C514 ASIG5V.n707 VSS 0.056945f
C515 ASIG5V.n708 VSS 0.056945f
C516 ASIG5V.n709 VSS 0.056945f
C517 ASIG5V.n711 VSS 0.056945f
C518 ASIG5V.n712 VSS 0.056945f
C519 ASIG5V.n713 VSS 0.056945f
C520 ASIG5V.n714 VSS 0.056945f
C521 ASIG5V.n715 VSS 0.056945f
C522 ASIG5V.n716 VSS 0.056945f
C523 ASIG5V.n717 VSS 0.056945f
C524 ASIG5V.n719 VSS 0.056945f
C525 ASIG5V.n720 VSS 0.056945f
C526 ASIG5V.n721 VSS 0.056945f
C527 ASIG5V.n723 VSS 0.056945f
C528 ASIG5V.n724 VSS 0.056945f
C529 ASIG5V.n725 VSS 0.056945f
C530 ASIG5V.n726 VSS 0.056945f
C531 ASIG5V.n727 VSS 0.056945f
C532 ASIG5V.n728 VSS 0.056945f
C533 ASIG5V.n729 VSS 0.056945f
C534 ASIG5V.n731 VSS 0.056945f
C535 ASIG5V.n732 VSS 0.056945f
C536 ASIG5V.n733 VSS 0.056945f
C537 ASIG5V.n735 VSS 0.056945f
C538 ASIG5V.n736 VSS 0.056945f
C539 ASIG5V.n737 VSS 0.056945f
C540 ASIG5V.n738 VSS 0.056945f
C541 ASIG5V.n739 VSS 0.056945f
C542 ASIG5V.n740 VSS 0.056945f
C543 ASIG5V.n741 VSS 0.056945f
C544 ASIG5V.n743 VSS 0.056945f
C545 ASIG5V.n744 VSS 0.056945f
C546 ASIG5V.n745 VSS 0.056945f
C547 ASIG5V.n747 VSS 0.056945f
C548 ASIG5V.n748 VSS 0.056945f
C549 ASIG5V.n749 VSS 0.056945f
C550 ASIG5V.n750 VSS 0.056945f
C551 ASIG5V.n751 VSS 0.056945f
C552 ASIG5V.n752 VSS 0.056945f
C553 ASIG5V.n753 VSS 0.056945f
C554 ASIG5V.n755 VSS 0.056945f
C555 ASIG5V.n756 VSS 0.056945f
C556 ASIG5V.n757 VSS 0.056945f
C557 ASIG5V.n759 VSS 0.056945f
C558 ASIG5V.n760 VSS 0.056945f
C559 ASIG5V.n761 VSS 0.056945f
C560 ASIG5V.n762 VSS 0.056945f
C561 ASIG5V.n763 VSS 0.056945f
C562 ASIG5V.n764 VSS 0.056945f
C563 ASIG5V.n765 VSS 0.056945f
C564 ASIG5V.n767 VSS 0.056945f
C565 ASIG5V.n768 VSS 0.056945f
C566 ASIG5V.n769 VSS 0.056945f
C567 ASIG5V.n771 VSS 0.056945f
C568 ASIG5V.n772 VSS 0.056945f
C569 ASIG5V.n773 VSS 0.056945f
C570 ASIG5V.n774 VSS 0.056945f
C571 ASIG5V.n775 VSS 0.056945f
C572 ASIG5V.n776 VSS 0.056945f
C573 ASIG5V.n777 VSS 0.056945f
C574 ASIG5V.n779 VSS 0.056945f
C575 ASIG5V.n780 VSS 0.056945f
C576 ASIG5V.n781 VSS 0.056945f
C577 ASIG5V.n783 VSS 0.056945f
C578 ASIG5V.n784 VSS 0.056945f
C579 ASIG5V.n785 VSS 0.056945f
C580 ASIG5V.n786 VSS 0.056945f
C581 ASIG5V.n787 VSS 0.056945f
C582 ASIG5V.n788 VSS 0.056945f
C583 ASIG5V.n789 VSS 0.056945f
C584 ASIG5V.n791 VSS 0.056945f
C585 ASIG5V.n792 VSS 0.056945f
C586 ASIG5V.n793 VSS 0.056945f
C587 ASIG5V.n795 VSS 0.056945f
C588 ASIG5V.n796 VSS 0.056945f
C589 ASIG5V.n797 VSS 0.056945f
C590 ASIG5V.n798 VSS 0.056945f
C591 ASIG5V.n799 VSS 0.056945f
C592 ASIG5V.n800 VSS 0.056945f
C593 ASIG5V.n801 VSS 0.056945f
C594 ASIG5V.n803 VSS 0.056945f
C595 ASIG5V.n804 VSS 0.056945f
C596 ASIG5V.n805 VSS 0.056945f
C597 ASIG5V.n807 VSS 0.056945f
C598 ASIG5V.n808 VSS 0.056945f
C599 ASIG5V.n809 VSS 0.056945f
C600 ASIG5V.n810 VSS 0.056945f
C601 ASIG5V.n811 VSS 0.056945f
C602 ASIG5V.n812 VSS 0.056945f
C603 ASIG5V.n813 VSS 0.056945f
C604 ASIG5V.n815 VSS 0.056945f
C605 ASIG5V.n816 VSS 0.056945f
C606 ASIG5V.n817 VSS 0.056945f
C607 ASIG5V.n819 VSS 0.056945f
C608 ASIG5V.n820 VSS 0.056945f
C609 ASIG5V.n821 VSS 0.056945f
C610 ASIG5V.n822 VSS 0.056945f
C611 ASIG5V.n823 VSS 0.056945f
C612 ASIG5V.n824 VSS 0.056945f
C613 ASIG5V.n825 VSS 0.056945f
C614 ASIG5V.n827 VSS 0.056945f
C615 ASIG5V.n828 VSS 0.056945f
C616 ASIG5V.n829 VSS 0.056945f
C617 ASIG5V.n831 VSS 0.056945f
C618 ASIG5V.n832 VSS 0.056945f
C619 ASIG5V.n833 VSS 0.056945f
C620 ASIG5V.n834 VSS 0.056945f
C621 ASIG5V.n835 VSS 0.056945f
C622 ASIG5V.n836 VSS 0.056945f
C623 ASIG5V.n837 VSS 0.056945f
C624 ASIG5V.n839 VSS 0.056945f
C625 ASIG5V.n840 VSS 0.056945f
C626 ASIG5V.n841 VSS 0.056945f
C627 ASIG5V.n843 VSS 0.056945f
C628 ASIG5V.n844 VSS 0.056945f
C629 ASIG5V.n845 VSS 0.056945f
C630 ASIG5V.n846 VSS 0.056945f
C631 ASIG5V.n847 VSS 0.056945f
C632 ASIG5V.n848 VSS 0.056945f
C633 ASIG5V.n849 VSS 0.056945f
C634 ASIG5V.n851 VSS 0.056945f
C635 ASIG5V.n852 VSS 0.056945f
C636 ASIG5V.n853 VSS 0.056945f
C637 ASIG5V.n855 VSS 0.056945f
C638 ASIG5V.n856 VSS 0.056945f
C639 ASIG5V.n857 VSS 0.056945f
C640 ASIG5V.n858 VSS 0.056945f
C641 ASIG5V.n859 VSS 0.041282f
C642 ASIG5V.n860 VSS 0.066995f
C643 ASIG5V.n861 VSS 0.047268f
C644 ASIG5V.n862 VSS 0.045974f
C645 ASIG5V.n863 VSS 0.076709f
C646 ASIG5V.n864 VSS 0.040245f
C647 ASIG5V.n865 VSS 1.0941f
C648 ASIG5V.n866 VSS 0.955416f
C649 ASIG5V.n867 VSS 0.063267f
C650 ASIG5V.n868 VSS 0.063267f
C651 ASIG5V.n869 VSS 0.052133f
C652 ASIG5V.n870 VSS 0.094123f
C653 ASIG5V.n871 VSS 0.0621f
C654 ASIG5V.n872 VSS 0.108961f
C655 ASIG5V.n873 VSS 0.0621f
C656 ASIG5V.n874 VSS 0.108961f
C657 ASIG5V.n875 VSS 0.485412f
C658 ASIG5V.n876 VSS 0.708856f
C659 ASIG5V.n877 VSS 0.855251f
C660 ASIG5V.n878 VSS 1.0941f
C661 ASIG5V.n879 VSS 0.045974f
C662 ASIG5V.n880 VSS 0.071577f
C663 ASIG5V.n881 VSS 0.045974f
C664 ASIG5V.n882 VSS 0.071577f
C665 ASIG5V.n883 VSS 0.056945f
C666 ASIG5V.n884 VSS 0.056945f
C667 ASIG5V.n885 VSS 0.056945f
C668 ASIG5V.n887 VSS 0.056945f
C669 ASIG5V.n888 VSS 0.056945f
C670 ASIG5V.n889 VSS 0.056945f
C671 ASIG5V.n891 VSS 0.056945f
C672 ASIG5V.n892 VSS 0.056945f
C673 ASIG5V.n893 VSS 0.056945f
C674 ASIG5V.n895 VSS 0.056945f
C675 ASIG5V.n896 VSS 0.056945f
C676 ASIG5V.n897 VSS 0.056945f
C677 ASIG5V.n899 VSS 0.056945f
C678 ASIG5V.n900 VSS 0.056945f
C679 ASIG5V.n901 VSS 0.056945f
C680 ASIG5V.n903 VSS 0.056945f
C681 ASIG5V.n904 VSS 0.056945f
C682 ASIG5V.n905 VSS 0.056945f
C683 ASIG5V.n907 VSS 0.056945f
C684 ASIG5V.n908 VSS 0.056945f
C685 ASIG5V.n909 VSS 0.056945f
C686 ASIG5V.n911 VSS 0.056945f
C687 ASIG5V.n912 VSS 0.056945f
C688 ASIG5V.n913 VSS 0.056945f
C689 ASIG5V.n915 VSS 0.056945f
C690 ASIG5V.n916 VSS 0.056945f
C691 ASIG5V.n917 VSS 0.056945f
C692 ASIG5V.n919 VSS 0.056945f
C693 ASIG5V.n920 VSS 0.056945f
C694 ASIG5V.n921 VSS 0.056945f
C695 ASIG5V.n923 VSS 0.056945f
C696 ASIG5V.n924 VSS 0.056945f
C697 ASIG5V.n925 VSS 0.056945f
C698 ASIG5V.n927 VSS 0.056945f
C699 ASIG5V.n928 VSS 0.056945f
C700 ASIG5V.n929 VSS 0.056945f
C701 ASIG5V.n931 VSS 0.056945f
C702 ASIG5V.n932 VSS 0.056945f
C703 ASIG5V.n933 VSS 0.056945f
C704 ASIG5V.n935 VSS 0.056945f
C705 ASIG5V.n936 VSS 0.056945f
C706 ASIG5V.n937 VSS 0.056945f
C707 ASIG5V.n939 VSS 0.056945f
C708 ASIG5V.n940 VSS 0.056945f
C709 ASIG5V.n941 VSS 0.056945f
C710 ASIG5V.n943 VSS 0.056945f
C711 ASIG5V.n944 VSS 0.056945f
C712 ASIG5V.n945 VSS 0.056945f
C713 ASIG5V.n947 VSS 0.056945f
C714 ASIG5V.n948 VSS 0.056945f
C715 ASIG5V.n949 VSS 0.056945f
C716 ASIG5V.n951 VSS 0.056945f
C717 ASIG5V.n952 VSS 0.056945f
C718 ASIG5V.n953 VSS 0.056945f
C719 ASIG5V.n955 VSS 0.056945f
C720 ASIG5V.n956 VSS 0.056945f
C721 ASIG5V.n957 VSS 0.056945f
C722 ASIG5V.n959 VSS 0.056945f
C723 ASIG5V.n960 VSS 0.056945f
C724 ASIG5V.n961 VSS 0.056945f
C725 ASIG5V.n963 VSS 0.056945f
C726 ASIG5V.n964 VSS 0.056945f
C727 ASIG5V.n965 VSS 0.056945f
C728 ASIG5V.n966 VSS 0.036092f
C729 ASIG5V.n967 VSS 0.036092f
C730 ASIG5V.n969 VSS 0.056945f
C731 ASIG5V.n971 VSS 0.056945f
C732 ASIG5V.n973 VSS 0.056945f
C733 ASIG5V.n974 VSS 0.056945f
C734 ASIG5V.n975 VSS 0.056945f
C735 ASIG5V.n976 VSS 0.056945f
C736 ASIG5V.n977 VSS 0.056945f
C737 ASIG5V.n978 VSS 0.056945f
C738 ASIG5V.n979 VSS 0.056945f
C739 ASIG5V.n981 VSS 0.056945f
C740 ASIG5V.n983 VSS 0.056945f
C741 ASIG5V.n985 VSS 0.056945f
C742 ASIG5V.n986 VSS 0.056945f
C743 ASIG5V.n987 VSS 0.056945f
C744 ASIG5V.n988 VSS 0.056945f
C745 ASIG5V.n989 VSS 0.056945f
C746 ASIG5V.n990 VSS 0.056945f
C747 ASIG5V.n991 VSS 0.056945f
C748 ASIG5V.n993 VSS 0.056945f
C749 ASIG5V.n995 VSS 0.056945f
C750 ASIG5V.n997 VSS 0.056945f
C751 ASIG5V.n998 VSS 0.056945f
C752 ASIG5V.n999 VSS 0.056945f
C753 ASIG5V.n1000 VSS 0.056945f
C754 ASIG5V.n1001 VSS 0.056945f
C755 ASIG5V.n1002 VSS 0.056945f
C756 ASIG5V.n1003 VSS 0.056945f
C757 ASIG5V.n1005 VSS 0.056945f
C758 ASIG5V.n1007 VSS 0.056945f
C759 ASIG5V.n1009 VSS 0.056945f
C760 ASIG5V.n1010 VSS 0.056945f
C761 ASIG5V.n1011 VSS 0.056945f
C762 ASIG5V.n1012 VSS 0.056945f
C763 ASIG5V.n1013 VSS 0.056945f
C764 ASIG5V.n1014 VSS 0.056945f
C765 ASIG5V.n1015 VSS 0.056945f
C766 ASIG5V.n1017 VSS 0.056945f
C767 ASIG5V.n1019 VSS 0.056945f
C768 ASIG5V.n1021 VSS 0.056945f
C769 ASIG5V.n1022 VSS 0.056945f
C770 ASIG5V.n1023 VSS 0.056945f
C771 ASIG5V.n1024 VSS 0.056945f
C772 ASIG5V.n1025 VSS 0.056945f
C773 ASIG5V.n1026 VSS 0.056945f
C774 ASIG5V.n1027 VSS 0.056945f
C775 ASIG5V.n1029 VSS 0.056945f
C776 ASIG5V.n1031 VSS 0.056945f
C777 ASIG5V.n1033 VSS 0.056945f
C778 ASIG5V.n1034 VSS 0.056945f
C779 ASIG5V.n1035 VSS 0.056945f
C780 ASIG5V.n1036 VSS 0.056945f
C781 ASIG5V.n1037 VSS 0.056945f
C782 ASIG5V.n1038 VSS 0.056945f
C783 ASIG5V.n1039 VSS 0.056945f
C784 ASIG5V.n1041 VSS 0.056945f
C785 ASIG5V.n1043 VSS 0.056945f
C786 ASIG5V.n1045 VSS 0.056945f
C787 ASIG5V.n1046 VSS 0.056945f
C788 ASIG5V.n1047 VSS 0.056945f
C789 ASIG5V.n1048 VSS 0.056945f
C790 ASIG5V.n1049 VSS 0.056945f
C791 ASIG5V.n1050 VSS 0.056945f
C792 ASIG5V.n1051 VSS 0.056945f
C793 ASIG5V.n1053 VSS 0.056945f
C794 ASIG5V.n1055 VSS 0.056945f
C795 ASIG5V.n1057 VSS 0.056945f
C796 ASIG5V.n1058 VSS 0.056945f
C797 ASIG5V.n1059 VSS 0.056945f
C798 ASIG5V.n1060 VSS 0.056945f
C799 ASIG5V.n1061 VSS 0.056945f
C800 ASIG5V.n1062 VSS 0.056945f
C801 ASIG5V.n1063 VSS 0.056945f
C802 ASIG5V.n1065 VSS 0.056945f
C803 ASIG5V.n1067 VSS 0.056945f
C804 ASIG5V.n1069 VSS 0.056945f
C805 ASIG5V.n1070 VSS 0.056945f
C806 ASIG5V.n1071 VSS 0.056945f
C807 ASIG5V.n1072 VSS 0.056945f
C808 ASIG5V.n1073 VSS 0.056945f
C809 ASIG5V.n1074 VSS 0.056945f
C810 ASIG5V.n1075 VSS 0.056945f
C811 ASIG5V.n1077 VSS 0.056945f
C812 ASIG5V.n1079 VSS 0.056945f
C813 ASIG5V.n1081 VSS 0.056945f
C814 ASIG5V.n1082 VSS 0.056945f
C815 ASIG5V.n1083 VSS 0.056945f
C816 ASIG5V.n1084 VSS 0.056945f
C817 ASIG5V.n1085 VSS 0.056945f
C818 ASIG5V.n1086 VSS 0.056945f
C819 ASIG5V.n1087 VSS 0.056945f
C820 ASIG5V.n1089 VSS 0.056945f
C821 ASIG5V.n1091 VSS 0.056945f
C822 ASIG5V.n1093 VSS 0.056945f
C823 ASIG5V.n1094 VSS 0.056945f
C824 ASIG5V.n1095 VSS 0.056945f
C825 ASIG5V.n1096 VSS 0.056945f
C826 ASIG5V.n1097 VSS 0.056945f
C827 ASIG5V.n1098 VSS 0.056945f
C828 ASIG5V.n1099 VSS 0.056945f
C829 ASIG5V.n1101 VSS 0.056945f
C830 ASIG5V.n1103 VSS 0.056945f
C831 ASIG5V.n1105 VSS 0.056945f
C832 ASIG5V.n1106 VSS 0.056945f
C833 ASIG5V.n1107 VSS 0.056945f
C834 ASIG5V.n1108 VSS 0.056945f
C835 ASIG5V.n1109 VSS 0.056945f
C836 ASIG5V.n1110 VSS 0.056945f
C837 ASIG5V.n1111 VSS 0.056945f
C838 ASIG5V.n1113 VSS 0.056945f
C839 ASIG5V.n1115 VSS 0.056945f
C840 ASIG5V.n1117 VSS 0.056945f
C841 ASIG5V.n1118 VSS 0.056945f
C842 ASIG5V.n1119 VSS 0.056945f
C843 ASIG5V.n1120 VSS 0.056945f
C844 ASIG5V.n1121 VSS 0.056945f
C845 ASIG5V.n1122 VSS 0.056945f
C846 ASIG5V.n1123 VSS 0.056945f
C847 ASIG5V.n1125 VSS 0.056945f
C848 ASIG5V.n1127 VSS 0.056945f
C849 ASIG5V.n1129 VSS 0.056945f
C850 ASIG5V.n1130 VSS 0.056945f
C851 ASIG5V.n1131 VSS 0.056945f
C852 ASIG5V.n1132 VSS 0.056945f
C853 ASIG5V.n1133 VSS 0.056945f
C854 ASIG5V.n1134 VSS 0.056945f
C855 ASIG5V.n1135 VSS 0.056945f
C856 ASIG5V.n1137 VSS 0.056945f
C857 ASIG5V.n1139 VSS 0.056945f
C858 ASIG5V.n1141 VSS 0.056945f
C859 ASIG5V.n1142 VSS 0.056945f
C860 ASIG5V.n1143 VSS 0.056945f
C861 ASIG5V.n1144 VSS 0.056945f
C862 ASIG5V.n1145 VSS 0.056945f
C863 ASIG5V.n1146 VSS 0.056945f
C864 ASIG5V.n1147 VSS 0.056945f
C865 ASIG5V.n1149 VSS 0.056945f
C866 ASIG5V.n1151 VSS 0.056945f
C867 ASIG5V.n1153 VSS 0.056945f
C868 ASIG5V.n1154 VSS 0.056945f
C869 ASIG5V.n1155 VSS 0.056945f
C870 ASIG5V.n1156 VSS 0.056945f
C871 ASIG5V.n1157 VSS 0.056945f
C872 ASIG5V.n1158 VSS 0.056945f
C873 ASIG5V.n1159 VSS 0.056945f
C874 ASIG5V.n1161 VSS 0.056945f
C875 ASIG5V.n1163 VSS 0.056945f
C876 ASIG5V.n1165 VSS 0.056945f
C877 ASIG5V.n1166 VSS 0.056945f
C878 ASIG5V.n1167 VSS 0.056945f
C879 ASIG5V.n1168 VSS 0.056945f
C880 ASIG5V.n1169 VSS 0.056945f
C881 ASIG5V.n1170 VSS 0.056945f
C882 ASIG5V.n1171 VSS 0.056945f
C883 ASIG5V.n1173 VSS 0.056945f
C884 ASIG5V.n1175 VSS 0.056945f
C885 ASIG5V.n1177 VSS 0.056945f
C886 ASIG5V.n1178 VSS 0.056945f
C887 ASIG5V.n1179 VSS 0.056945f
C888 ASIG5V.n1180 VSS 0.056945f
C889 ASIG5V.n1181 VSS 0.056945f
C890 ASIG5V.n1182 VSS 0.056945f
C891 ASIG5V.n1183 VSS 0.056945f
C892 ASIG5V.n1185 VSS 0.056945f
C893 ASIG5V.n1187 VSS 0.056945f
C894 ASIG5V.n1189 VSS 0.056945f
C895 ASIG5V.n1190 VSS 0.056945f
C896 ASIG5V.n1191 VSS 0.056945f
C897 ASIG5V.n1192 VSS 0.056945f
C898 ASIG5V.n1193 VSS 0.056945f
C899 ASIG5V.n1194 VSS 0.056945f
C900 ASIG5V.n1195 VSS 0.056945f
C901 ASIG5V.n1197 VSS 0.056945f
C902 ASIG5V.n1199 VSS 0.056945f
C903 ASIG5V.n1201 VSS 0.056945f
C904 ASIG5V.n1202 VSS 0.056945f
C905 ASIG5V.n1203 VSS 0.056945f
C906 ASIG5V.n1204 VSS 0.056945f
C907 ASIG5V.n1205 VSS 0.056945f
C908 ASIG5V.n1206 VSS 0.056945f
C909 ASIG5V.n1207 VSS 0.056945f
C910 ASIG5V.n1208 VSS 0.056945f
C911 ASIG5V.n1210 VSS 0.056945f
C912 ASIG5V.n1212 VSS 0.056945f
C913 ASIG5V.n1214 VSS 0.036092f
C914 ASIG5V.n1215 VSS 0.036092f
C915 ASIG5V.n1216 VSS 0.047722f
C916 ASIG5V.n1217 VSS 0.040245f
C917 ASIG5V.n1218 VSS 0.035149f
C918 ASIG5V.n1219 VSS 0.052746f
C919 ASIG5V.n1220 VSS 0.047722f
C920 ASIG5V.n1221 VSS 0.066995f
C921 ASIG5V.n1222 VSS 0.045974f
C922 ASIG5V.n1223 VSS 0.076709f
C923 ASIG5V.n1224 VSS 0.045974f
C924 ASIG5V.n1225 VSS 0.076709f
C925 ASIG5V.n1226 VSS 0.685742f
C926 ASIG5V.n1268 VSS 0.036092f
C927 ASIG5V.n1269 VSS 0.685742f
C928 ASIG5V.n1270 VSS 0.036092f
C929 ASIG5V.n1271 VSS 0.785906f
C930 ASIG5V.n1272 VSS 0.577872f
C931 ASIG5V.n1273 VSS 0.056945f
C932 ASIG5V.n1274 VSS 0.056945f
C933 ASIG5V.n1275 VSS 0.056945f
C934 ASIG5V.n1276 VSS 0.056945f
C935 ASIG5V.n1277 VSS 0.056945f
C936 ASIG5V.n1278 VSS 0.056945f
C937 ASIG5V.n1279 VSS 0.056945f
C938 ASIG5V.n1280 VSS 0.056945f
C939 ASIG5V.n1281 VSS 0.056945f
C940 ASIG5V.n1282 VSS 0.056945f
C941 ASIG5V.n1283 VSS 0.056945f
C942 ASIG5V.n1284 VSS 0.056945f
C943 ASIG5V.n1285 VSS 0.056945f
C944 ASIG5V.n1286 VSS 0.056945f
C945 ASIG5V.n1287 VSS 0.056945f
C946 ASIG5V.n1288 VSS 0.056945f
C947 ASIG5V.n1289 VSS 0.056945f
C948 ASIG5V.n1290 VSS 0.056945f
C949 ASIG5V.n1291 VSS 0.056945f
C950 ASIG5V.n1292 VSS 0.056945f
C951 ASIG5V.n1293 VSS 0.056945f
C952 ASIG5V.n1294 VSS 0.056945f
C953 ASIG5V.n1295 VSS 0.056945f
C954 ASIG5V.n1296 VSS 0.056945f
C955 ASIG5V.n1297 VSS 0.056945f
C956 ASIG5V.n1298 VSS 0.056945f
C957 ASIG5V.n1299 VSS 0.056945f
C958 ASIG5V.n1300 VSS 0.056945f
C959 ASIG5V.n1301 VSS 0.056945f
C960 ASIG5V.n1302 VSS 0.056945f
C961 ASIG5V.n1303 VSS 0.056945f
C962 ASIG5V.n1304 VSS 0.056945f
C963 ASIG5V.n1305 VSS 0.056945f
C964 ASIG5V.n1306 VSS 0.056945f
C965 ASIG5V.n1307 VSS 0.056945f
C966 ASIG5V.n1308 VSS 0.056945f
C967 ASIG5V.n1309 VSS 0.056945f
C968 ASIG5V.n1310 VSS 0.056945f
C969 ASIG5V.n1311 VSS 0.056945f
C970 ASIG5V.n1312 VSS 0.056945f
C971 ASIG5V.n1314 VSS 0.056945f
C972 ASIG5V.n1315 VSS 0.056945f
C973 ASIG5V.n1316 VSS 0.07229f
C974 ASIG5V.n1317 VSS 0.075569f
C975 ASIG5V.n1318 VSS 0.108961f
C976 ASIG5V.n1319 VSS 0.075569f
C977 ASIG5V.n1320 VSS 0.0621f
C978 ASIG5V.n1321 VSS 0.087871f
C979 ASIG5V.n1322 VSS 0.07229f
C980 ASIG5V.n1323 VSS 0.0621f
C981 ASIG5V.n1324 VSS 0.108961f
C982 ASIG5V.n1325 VSS 0.0621f
C983 ASIG5V.n1326 VSS 0.955415f
C984 ASIG5V.n1327 VSS 1.0941f
C985 ASIG5V.n1328 VSS 0.955415f
C986 ASIG5V.n1370 VSS 0.870661f
C987 ASIG5V.n1371 VSS 0.056945f
C988 ASIG5V.n1372 VSS 0.036092f
C989 ASIG5V.n1373 VSS 0.246558f
C990 ASIG5V.n1415 VSS 0.847545f
C991 ASIG5V.n1416 VSS 0.045974f
C992 ASIG5V.n1417 VSS 0.056945f
C993 ASIG5V.n1418 VSS 0.056945f
C994 ASIG5V.n1419 VSS 0.056945f
C995 ASIG5V.n1420 VSS 0.056945f
C996 ASIG5V.n1421 VSS 0.056945f
C997 ASIG5V.n1422 VSS 0.056945f
C998 ASIG5V.n1423 VSS 0.056945f
C999 ASIG5V.n1424 VSS 0.056945f
C1000 ASIG5V.n1425 VSS 0.056945f
C1001 ASIG5V.n1426 VSS 0.056945f
C1002 ASIG5V.n1427 VSS 0.056945f
C1003 ASIG5V.n1428 VSS 0.056945f
C1004 ASIG5V.n1429 VSS 0.056945f
C1005 ASIG5V.n1430 VSS 0.056945f
C1006 ASIG5V.n1431 VSS 0.056945f
C1007 ASIG5V.n1432 VSS 0.056945f
C1008 ASIG5V.n1433 VSS 0.056945f
C1009 ASIG5V.n1434 VSS 0.056945f
C1010 ASIG5V.n1435 VSS 0.056945f
C1011 ASIG5V.n1436 VSS 0.056945f
C1012 ASIG5V.n1437 VSS 0.056945f
C1013 ASIG5V.n1438 VSS 0.056945f
C1014 ASIG5V.n1439 VSS 0.056945f
C1015 ASIG5V.n1440 VSS 0.056945f
C1016 ASIG5V.n1441 VSS 0.056945f
C1017 ASIG5V.n1442 VSS 0.056945f
C1018 ASIG5V.n1443 VSS 0.056945f
C1019 ASIG5V.n1444 VSS 0.056945f
C1020 ASIG5V.n1445 VSS 0.056945f
C1021 ASIG5V.n1446 VSS 0.056945f
C1022 ASIG5V.n1447 VSS 0.056945f
C1023 ASIG5V.n1448 VSS 0.056945f
C1024 ASIG5V.n1449 VSS 0.056945f
C1025 ASIG5V.n1450 VSS 0.056945f
C1026 ASIG5V.n1451 VSS 0.056945f
C1027 ASIG5V.n1452 VSS 0.056945f
C1028 ASIG5V.n1453 VSS 0.056945f
C1029 ASIG5V.n1454 VSS 0.056945f
C1030 ASIG5V.n1455 VSS 0.056945f
C1031 ASIG5V.n1456 VSS 0.056945f
C1032 ASIG5V.n1457 VSS 0.056945f
C1033 ASIG5V.n1458 VSS 0.056945f
C1034 ASIG5V.n1459 VSS 0.056945f
C1035 ASIG5V.n1460 VSS 0.056945f
C1036 ASIG5V.n1461 VSS 0.056945f
C1037 ASIG5V.n1462 VSS 0.056945f
C1038 ASIG5V.n1463 VSS 0.056945f
C1039 ASIG5V.n1464 VSS 0.056945f
C1040 ASIG5V.n1465 VSS 0.056945f
C1041 ASIG5V.n1466 VSS 0.056945f
C1042 ASIG5V.n1467 VSS 0.056945f
C1043 ASIG5V.n1468 VSS 0.056945f
C1044 ASIG5V.n1469 VSS 0.056945f
C1045 ASIG5V.n1470 VSS 0.056945f
C1046 ASIG5V.n1471 VSS 0.056945f
C1047 ASIG5V.n1472 VSS 0.056945f
C1048 ASIG5V.n1473 VSS 0.056945f
C1049 ASIG5V.n1474 VSS 0.056945f
C1050 ASIG5V.n1475 VSS 0.056945f
C1051 ASIG5V.n1476 VSS 0.056945f
C1052 ASIG5V.n1477 VSS 0.056945f
C1053 ASIG5V.n1478 VSS 0.056945f
C1054 ASIG5V.n1479 VSS 0.052133f
C1055 ASIG5V.n1480 VSS 0.056945f
C1056 ASIG5V.n1481 VSS 0.056945f
C1057 ASIG5V.n1482 VSS 0.056945f
C1058 ASIG5V.n1483 VSS 0.056945f
C1059 ASIG5V.n1484 VSS 0.056945f
C1060 ASIG5V.n1485 VSS 0.056945f
C1061 ASIG5V.n1486 VSS 0.056945f
C1062 ASIG5V.n1487 VSS 0.056945f
C1063 ASIG5V.n1488 VSS 0.056945f
C1064 ASIG5V.n1489 VSS 0.056945f
C1065 ASIG5V.n1490 VSS 0.056945f
C1066 ASIG5V.n1491 VSS 0.056945f
C1067 ASIG5V.n1492 VSS 0.056945f
C1068 ASIG5V.n1493 VSS 0.056945f
C1069 ASIG5V.n1494 VSS 0.056945f
C1070 ASIG5V.n1495 VSS 0.056945f
C1071 ASIG5V.n1496 VSS 0.056945f
C1072 ASIG5V.n1497 VSS 0.056945f
C1073 ASIG5V.n1498 VSS 0.056945f
C1074 ASIG5V.n1499 VSS 0.056945f
C1075 ASIG5V.n1500 VSS 0.056945f
C1076 ASIG5V.n1501 VSS 0.056945f
C1077 ASIG5V.n1502 VSS 0.056945f
C1078 ASIG5V.n1503 VSS 0.056945f
C1079 ASIG5V.n1504 VSS 0.056945f
C1080 ASIG5V.n1505 VSS 0.056945f
C1081 ASIG5V.n1506 VSS 0.056945f
C1082 ASIG5V.n1507 VSS 0.056945f
C1083 ASIG5V.n1508 VSS 0.056945f
C1084 ASIG5V.n1509 VSS 0.056945f
C1085 ASIG5V.n1510 VSS 0.056945f
C1086 ASIG5V.n1511 VSS 0.056945f
C1087 ASIG5V.n1512 VSS 0.056945f
C1088 ASIG5V.n1513 VSS 0.056945f
C1089 ASIG5V.n1514 VSS 0.056945f
C1090 ASIG5V.n1515 VSS 0.056945f
C1091 ASIG5V.n1516 VSS 0.056945f
C1092 ASIG5V.n1517 VSS 0.056945f
C1093 ASIG5V.n1518 VSS 0.056945f
C1094 ASIG5V.n1519 VSS 0.056945f
C1095 ASIG5V.n1520 VSS 0.056945f
C1096 ASIG5V.n1521 VSS 0.056945f
C1097 ASIG5V.n1522 VSS 0.056945f
C1098 ASIG5V.n1523 VSS 0.056945f
C1099 ASIG5V.n1524 VSS 0.056945f
C1100 ASIG5V.n1525 VSS 0.056945f
C1101 ASIG5V.n1526 VSS 0.056945f
C1102 ASIG5V.n1527 VSS 0.056945f
C1103 ASIG5V.n1528 VSS 0.056945f
C1104 ASIG5V.n1529 VSS 0.056945f
C1105 ASIG5V.n1530 VSS 0.056945f
C1106 ASIG5V.n1531 VSS 0.056945f
C1107 ASIG5V.n1532 VSS 0.056945f
C1108 ASIG5V.n1533 VSS 0.056945f
C1109 ASIG5V.n1534 VSS 0.056945f
C1110 ASIG5V.n1535 VSS 0.056945f
C1111 ASIG5V.n1536 VSS 0.056945f
C1112 ASIG5V.n1537 VSS 0.056945f
C1113 ASIG5V.n1538 VSS 0.056945f
C1114 ASIG5V.n1539 VSS 0.056945f
C1115 ASIG5V.n1540 VSS 0.056945f
C1116 ASIG5V.n1541 VSS 0.056945f
C1117 ASIG5V.n1542 VSS 0.056945f
C1118 ASIG5V.n1543 VSS 0.056945f
C1119 ASIG5V.n1544 VSS 0.056945f
C1120 ASIG5V.n1545 VSS 0.056945f
C1121 ASIG5V.n1546 VSS 0.056945f
C1122 ASIG5V.n1547 VSS 0.056945f
C1123 ASIG5V.n1548 VSS 0.056945f
C1124 ASIG5V.n1549 VSS 0.056945f
C1125 ASIG5V.n1550 VSS 0.056945f
C1126 ASIG5V.n1551 VSS 0.056945f
C1127 ASIG5V.n1552 VSS 0.056945f
C1128 ASIG5V.n1553 VSS 0.056945f
C1129 ASIG5V.n1554 VSS 0.056945f
C1130 ASIG5V.n1555 VSS 0.056945f
C1131 ASIG5V.n1556 VSS 0.056945f
C1132 ASIG5V.n1557 VSS 0.056945f
C1133 ASIG5V.n1558 VSS 0.056945f
C1134 ASIG5V.n1559 VSS 0.056945f
C1135 ASIG5V.n1560 VSS 0.056945f
C1136 ASIG5V.n1561 VSS 0.056945f
C1137 ASIG5V.n1562 VSS 0.056945f
C1138 ASIG5V.n1563 VSS 0.056945f
C1139 ASIG5V.n1564 VSS 0.056945f
C1140 ASIG5V.n1565 VSS 0.056945f
C1141 ASIG5V.n1566 VSS 0.056945f
C1142 ASIG5V.n1567 VSS 0.056945f
C1143 ASIG5V.n1568 VSS 0.056945f
C1144 ASIG5V.n1569 VSS 0.056945f
C1145 ASIG5V.n1570 VSS 0.056945f
C1146 ASIG5V.n1571 VSS 0.056945f
C1147 ASIG5V.n1572 VSS 0.056945f
C1148 ASIG5V.n1573 VSS 0.056945f
C1149 ASIG5V.n1574 VSS 0.056945f
C1150 ASIG5V.n1575 VSS 0.056945f
C1151 ASIG5V.n1576 VSS 0.056945f
C1152 ASIG5V.n1577 VSS 0.056945f
C1153 ASIG5V.n1578 VSS 0.056945f
C1154 ASIG5V.n1579 VSS 0.056945f
C1155 ASIG5V.n1580 VSS 0.056945f
C1156 ASIG5V.n1581 VSS 0.056945f
C1157 ASIG5V.n1582 VSS 0.056945f
C1158 ASIG5V.n1583 VSS 0.056945f
C1159 ASIG5V.n1584 VSS 0.056945f
C1160 ASIG5V.n1585 VSS 0.056945f
C1161 ASIG5V.n1586 VSS 0.056945f
C1162 ASIG5V.n1587 VSS 0.056945f
C1163 ASIG5V.n1588 VSS 0.056945f
C1164 ASIG5V.n1589 VSS 0.056945f
C1165 ASIG5V.n1590 VSS 0.056945f
C1166 ASIG5V.n1591 VSS 0.056945f
C1167 ASIG5V.n1592 VSS 0.056945f
C1168 ASIG5V.n1593 VSS 0.056945f
C1169 ASIG5V.n1594 VSS 0.056945f
C1170 ASIG5V.n1595 VSS 0.056945f
C1171 ASIG5V.n1596 VSS 0.056945f
C1172 ASIG5V.n1597 VSS 0.056945f
C1173 ASIG5V.n1598 VSS 0.056945f
C1174 ASIG5V.n1599 VSS 0.056945f
C1175 ASIG5V.n1600 VSS 0.056945f
C1176 ASIG5V.n1601 VSS 0.056945f
C1177 ASIG5V.n1602 VSS 0.056945f
C1178 ASIG5V.n1603 VSS 0.056945f
C1179 ASIG5V.n1604 VSS 0.056945f
C1180 ASIG5V.n1605 VSS 0.056945f
C1181 ASIG5V.n1606 VSS 0.056945f
C1182 ASIG5V.n1607 VSS 0.056945f
C1183 ASIG5V.n1608 VSS 0.056945f
C1184 ASIG5V.n1609 VSS 0.056945f
C1185 ASIG5V.n1610 VSS 0.056945f
C1186 ASIG5V.n1611 VSS 0.056945f
C1187 ASIG5V.n1612 VSS 0.056945f
C1188 ASIG5V.n1613 VSS 0.056945f
C1189 ASIG5V.n1614 VSS 0.056945f
C1190 ASIG5V.n1615 VSS 0.056945f
C1191 ASIG5V.n1616 VSS 0.056945f
C1192 ASIG5V.n1617 VSS 0.056945f
C1193 ASIG5V.n1618 VSS 0.056945f
C1194 ASIG5V.n1619 VSS 0.056945f
C1195 ASIG5V.n1620 VSS 0.056945f
C1196 ASIG5V.n1621 VSS 0.056945f
C1197 ASIG5V.n1622 VSS 0.056945f
C1198 ASIG5V.n1623 VSS 0.056945f
C1199 ASIG5V.n1624 VSS 0.056945f
C1200 ASIG5V.n1625 VSS 0.056945f
C1201 ASIG5V.n1626 VSS 0.056945f
C1202 ASIG5V.n1627 VSS 0.056945f
C1203 ASIG5V.n1628 VSS 0.056945f
C1204 ASIG5V.n1629 VSS 0.056945f
C1205 ASIG5V.n1630 VSS 0.056945f
C1206 ASIG5V.n1631 VSS 0.056945f
C1207 ASIG5V.n1632 VSS 0.056945f
C1208 ASIG5V.n1633 VSS 0.056945f
C1209 ASIG5V.n1634 VSS 0.056945f
C1210 ASIG5V.n1635 VSS 0.056945f
C1211 ASIG5V.n1636 VSS 0.056945f
C1212 ASIG5V.n1637 VSS 0.056945f
C1213 ASIG5V.n1638 VSS 0.056945f
C1214 ASIG5V.n1639 VSS 0.056945f
C1215 ASIG5V.n1640 VSS 0.056945f
C1216 ASIG5V.n1641 VSS 0.056945f
C1217 ASIG5V.n1642 VSS 0.056945f
C1218 ASIG5V.n1643 VSS 0.056945f
C1219 ASIG5V.n1644 VSS 0.056945f
C1220 ASIG5V.n1645 VSS 0.056945f
C1221 ASIG5V.n1646 VSS 0.056945f
C1222 ASIG5V.n1647 VSS 0.056945f
C1223 ASIG5V.n1648 VSS 0.056945f
C1224 ASIG5V.n1649 VSS 0.056945f
C1225 ASIG5V.n1650 VSS 0.056945f
C1226 ASIG5V.n1651 VSS 0.056945f
C1227 ASIG5V.n1652 VSS 0.056945f
C1228 ASIG5V.n1653 VSS 0.056945f
C1229 ASIG5V.n1654 VSS 0.056945f
C1230 ASIG5V.n1655 VSS 0.056945f
C1231 ASIG5V.n1656 VSS 0.056945f
C1232 ASIG5V.n1657 VSS 0.056945f
C1233 ASIG5V.n1658 VSS 0.056945f
C1234 ASIG5V.n1659 VSS 0.056945f
C1235 ASIG5V.n1660 VSS 0.056945f
C1236 ASIG5V.n1661 VSS 0.056945f
C1237 ASIG5V.n1662 VSS 0.056945f
C1238 ASIG5V.n1663 VSS 0.047722f
C1239 ASIG5V.n1664 VSS 0.064554f
C1240 ASIG5V.n1665 VSS 0.064554f
C1241 ASIG5V.n1666 VSS 0.076709f
C1242 ASIG5V.n1667 VSS 0.050509f
C1243 ASIG5V.n1668 VSS 0.056379f
C1244 ASIG5V.n1669 VSS 0.052746f
C1245 ASIG5V.n1670 VSS 0.052746f
C1246 ASIG5V.n1671 VSS 0.045974f
C1247 ASIG5V.n1672 VSS 0.076709f
C1248 ASIG5V.n1673 VSS 0.045974f
C1249 ASIG5V.n1674 VSS 0.955415f
C1250 ASIG5V.n1675 VSS 1.0941f
C1251 ASIG5V.n1717 VSS 1.07099f
C1252 ASIG5V.n1718 VSS 0.056945f
C1253 ASIG5V.n1719 VSS 0.0621f
C1254 ASIG5V.n1720 VSS 0.036092f
C1255 ASIG5V.n1721 VSS 0.416067f
C1256 ASIG5V.n1763 VSS 1.07099f
C1257 ASIG5V.n1764 VSS 0.056945f
C1258 ASIG5V.n1765 VSS 0.056945f
C1259 ASIG5V.n1766 VSS 0.056945f
C1260 ASIG5V.n1767 VSS 0.056945f
C1261 ASIG5V.n1768 VSS 0.056945f
C1262 ASIG5V.n1769 VSS 0.056945f
C1263 ASIG5V.n1770 VSS 0.056945f
C1264 ASIG5V.n1771 VSS 0.056945f
C1265 ASIG5V.n1772 VSS 0.056945f
C1266 ASIG5V.n1773 VSS 0.056945f
C1267 ASIG5V.n1774 VSS 0.056945f
C1268 ASIG5V.n1775 VSS 0.056945f
C1269 ASIG5V.n1776 VSS 0.056945f
C1270 ASIG5V.n1777 VSS 0.056945f
C1271 ASIG5V.n1778 VSS 0.056945f
C1272 ASIG5V.n1779 VSS 0.056945f
C1273 ASIG5V.n1780 VSS 0.056945f
C1274 ASIG5V.n1781 VSS 0.056945f
C1275 ASIG5V.n1782 VSS 0.056945f
C1276 ASIG5V.n1783 VSS 0.056945f
C1277 ASIG5V.n1784 VSS 0.056945f
C1278 ASIG5V.n1785 VSS 0.056945f
C1279 ASIG5V.n1786 VSS 0.056945f
C1280 ASIG5V.n1787 VSS 0.056945f
C1281 ASIG5V.n1788 VSS 0.056945f
C1282 ASIG5V.n1789 VSS 0.056945f
C1283 ASIG5V.n1790 VSS 0.056945f
C1284 ASIG5V.n1791 VSS 0.056945f
C1285 ASIG5V.n1792 VSS 0.056945f
C1286 ASIG5V.n1793 VSS 0.056945f
C1287 ASIG5V.n1794 VSS 0.056945f
C1288 ASIG5V.n1795 VSS 0.056945f
C1289 ASIG5V.n1796 VSS 0.056945f
C1290 ASIG5V.n1797 VSS 0.056945f
C1291 ASIG5V.n1798 VSS 0.056945f
C1292 ASIG5V.n1799 VSS 0.056945f
C1293 ASIG5V.n1800 VSS 0.056945f
C1294 ASIG5V.n1801 VSS 0.056945f
C1295 ASIG5V.n1802 VSS 0.056945f
C1296 ASIG5V.n1803 VSS 0.056945f
C1297 ASIG5V.n1804 VSS 0.056945f
C1298 ASIG5V.n1805 VSS 0.056945f
C1299 ASIG5V.n1806 VSS 0.056945f
C1300 ASIG5V.n1807 VSS 0.056945f
C1301 ASIG5V.n1808 VSS 0.056945f
C1302 ASIG5V.n1809 VSS 0.056945f
C1303 ASIG5V.n1810 VSS 0.056945f
C1304 ASIG5V.n1811 VSS 0.056945f
C1305 ASIG5V.n1812 VSS 0.056945f
C1306 ASIG5V.n1813 VSS 0.056945f
C1307 ASIG5V.n1814 VSS 0.056945f
C1308 ASIG5V.n1815 VSS 0.056945f
C1309 ASIG5V.n1816 VSS 0.056945f
C1310 ASIG5V.n1817 VSS 0.056945f
C1311 ASIG5V.n1818 VSS 0.056945f
C1312 ASIG5V.n1819 VSS 0.056945f
C1313 ASIG5V.n1820 VSS 0.056945f
C1314 ASIG5V.n1821 VSS 0.056945f
C1315 ASIG5V.n1822 VSS 0.056945f
C1316 ASIG5V.n1823 VSS 0.056945f
C1317 ASIG5V.n1824 VSS 0.056945f
C1318 ASIG5V.n1825 VSS 0.056945f
C1319 ASIG5V.n1826 VSS 0.089417f
C1320 ASIG5V.n1827 VSS 0.09726f
C1321 ASIG5V.n1828 VSS 0.108961f
C1322 ASIG5V.n1829 VSS 0.09726f
C1323 ASIG5V.n1830 VSS 0.067455f
C1324 ASIG5V.n1831 VSS 0.075569f
C1325 ASIG5V.n1832 VSS 0.075569f
C1326 ASIG5V.n1833 VSS 0.108961f
C1327 ASIG5V.n1834 VSS 0.100173f
C1328 ASIG5V.n1835 VSS 0.100173f
C1329 ASIG5V.n1836 VSS 0.0621f
C1330 ASIG5V.n1837 VSS 0.108961f
C1331 ASIG5V.n1838 VSS 0.057995f
C1332 ASIG5V.n1839 VSS 0.916891f
C1333 ASIG5V.n1840 VSS 0.057995f
C1334 ASIG5V.n1841 VSS 0.536863f
C1335 ASIG5V.n1842 VSS 0.052133f
C1336 ASIG5V.n1843 VSS 0.09726f
C1337 ASIG5V.n1844 VSS 0.0621f
C1338 ASIG5V.n1845 VSS 0.108961f
C1339 ASIG5V.n1846 VSS 0.0621f
C1340 ASIG5V.n1847 VSS 0.108961f
C1341 ASIG5V.n1848 VSS 0.323607f
C1342 ASIG5V.n1849 VSS 0.685742f
C1343 ASIG5V.n1850 VSS 0.064554f
C1344 ASIG5V.n1851 VSS 0.043486f
C1345 ASIG5V.n1852 VSS 0.064554f
C1346 ASIG5V.n1853 VSS 0.043486f
C1347 ASIG5V.n1854 VSS 0.047722f
C1348 ASIG5V.n1855 VSS 0.066995f
C1349 ASIG5V.n1856 VSS 0.076709f
C1350 ASIG5V.n1857 VSS 0.045974f
C1351 ASIG5V.n1858 VSS 0.050246f
C1352 ASIG5V.n1859 VSS 0.057532f
C1353 ASIG5V.n1860 VSS 0.057532f
C1354 ASIG5V.n1861 VSS 0.955415f
C1355 ASIG5V.n1862 VSS 0.076709f
C1356 ASIG5V.n1863 VSS 0.045974f
C1357 ASIG5V.n1864 VSS 0.670332f
C1358 ASIG5V.n1906 VSS 0.036092f
C1359 ASIG5V.n1907 VSS 0.036092f
C1360 ASIG5V.n1908 VSS 0.056945f
C1361 ASIG5V.n1909 VSS 0.056945f
C1362 ASIG5V.n1910 VSS 0.056945f
C1363 ASIG5V.n1911 VSS 0.056945f
C1364 ASIG5V.n1912 VSS 0.056945f
C1365 ASIG5V.n1913 VSS 0.056945f
C1366 ASIG5V.n1914 VSS 0.056945f
C1367 ASIG5V.n1915 VSS 0.056945f
C1368 ASIG5V.n1916 VSS 0.056945f
C1369 ASIG5V.n1917 VSS 0.056945f
C1370 ASIG5V.n1918 VSS 0.056945f
C1371 ASIG5V.n1919 VSS 0.056945f
C1372 ASIG5V.n1920 VSS 0.056945f
C1373 ASIG5V.n1921 VSS 0.056945f
C1374 ASIG5V.n1922 VSS 0.056945f
C1375 ASIG5V.n1923 VSS 0.056945f
C1376 ASIG5V.n1924 VSS 0.056945f
C1377 ASIG5V.n1925 VSS 0.056945f
C1378 ASIG5V.n1926 VSS 0.056945f
C1379 ASIG5V.n1927 VSS 0.056945f
C1380 ASIG5V.n1928 VSS 0.056945f
C1381 ASIG5V.n1929 VSS 0.056945f
C1382 ASIG5V.n1930 VSS 0.056945f
C1383 ASIG5V.n1931 VSS 0.056945f
C1384 ASIG5V.n1932 VSS 0.056945f
C1385 ASIG5V.n1933 VSS 0.056945f
C1386 ASIG5V.n1934 VSS 0.056945f
C1387 ASIG5V.n1935 VSS 0.056945f
C1388 ASIG5V.n1936 VSS 0.056945f
C1389 ASIG5V.n1937 VSS 0.056945f
C1390 ASIG5V.n1938 VSS 0.056945f
C1391 ASIG5V.n1939 VSS 0.056945f
C1392 ASIG5V.n1940 VSS 0.056945f
C1393 ASIG5V.n1941 VSS 0.056945f
C1394 ASIG5V.n1942 VSS 0.056945f
C1395 ASIG5V.n1943 VSS 0.056945f
C1396 ASIG5V.n1944 VSS 0.056945f
C1397 ASIG5V.n1945 VSS 0.056945f
C1398 ASIG5V.n1946 VSS 0.056945f
C1399 ASIG5V.n1947 VSS 0.056945f
C1400 ASIG5V.n1948 VSS 0.036092f
C1401 ASIG5V.n1950 VSS 0.056945f
C1402 ASIG5V.n1951 VSS 0.056945f
C1403 ASIG5V.n1952 VSS 0.056945f
C1404 ASIG5V.n1953 VSS 0.056945f
C1405 ASIG5V.n1954 VSS 0.056945f
C1406 ASIG5V.n1955 VSS 0.056945f
C1407 ASIG5V.n1957 VSS 0.056945f
C1408 ASIG5V.n1958 VSS 0.056945f
C1409 ASIG5V.n1959 VSS 0.056945f
C1410 ASIG5V.n1961 VSS 0.056945f
C1411 ASIG5V.n1962 VSS 0.056945f
C1412 ASIG5V.n1963 VSS 0.056945f
C1413 ASIG5V.n1964 VSS 0.056945f
C1414 ASIG5V.n1965 VSS 0.056945f
C1415 ASIG5V.n1966 VSS 0.056945f
C1416 ASIG5V.n1967 VSS 0.056945f
C1417 ASIG5V.n1969 VSS 0.056945f
C1418 ASIG5V.n1970 VSS 0.056945f
C1419 ASIG5V.n1971 VSS 0.056945f
C1420 ASIG5V.n1973 VSS 0.056945f
C1421 ASIG5V.n1974 VSS 0.056945f
C1422 ASIG5V.n1975 VSS 0.056945f
C1423 ASIG5V.n1976 VSS 0.056945f
C1424 ASIG5V.n1977 VSS 0.056945f
C1425 ASIG5V.n1978 VSS 0.056945f
C1426 ASIG5V.n1979 VSS 0.056945f
C1427 ASIG5V.n1981 VSS 0.056945f
C1428 ASIG5V.n1982 VSS 0.056945f
C1429 ASIG5V.n1983 VSS 0.056945f
C1430 ASIG5V.n1985 VSS 0.056945f
C1431 ASIG5V.n1986 VSS 0.056945f
C1432 ASIG5V.n1987 VSS 0.056945f
C1433 ASIG5V.n1988 VSS 0.056945f
C1434 ASIG5V.n1989 VSS 0.056945f
C1435 ASIG5V.n1990 VSS 0.056945f
C1436 ASIG5V.n1991 VSS 0.056945f
C1437 ASIG5V.n1993 VSS 0.056945f
C1438 ASIG5V.n1994 VSS 0.056945f
C1439 ASIG5V.n1995 VSS 0.056945f
C1440 ASIG5V.n1997 VSS 0.056945f
C1441 ASIG5V.n1998 VSS 0.056945f
C1442 ASIG5V.n1999 VSS 0.056945f
C1443 ASIG5V.n2000 VSS 0.056945f
C1444 ASIG5V.n2001 VSS 0.056945f
C1445 ASIG5V.n2002 VSS 0.056945f
C1446 ASIG5V.n2003 VSS 0.056945f
C1447 ASIG5V.n2005 VSS 0.056945f
C1448 ASIG5V.n2006 VSS 0.056945f
C1449 ASIG5V.n2007 VSS 0.056945f
C1450 ASIG5V.n2009 VSS 0.056945f
C1451 ASIG5V.n2010 VSS 0.056945f
C1452 ASIG5V.n2011 VSS 0.056945f
C1453 ASIG5V.n2012 VSS 0.056945f
C1454 ASIG5V.n2013 VSS 0.056945f
C1455 ASIG5V.n2014 VSS 0.056945f
C1456 ASIG5V.n2015 VSS 0.056945f
C1457 ASIG5V.n2017 VSS 0.056945f
C1458 ASIG5V.n2018 VSS 0.056945f
C1459 ASIG5V.n2019 VSS 0.056945f
C1460 ASIG5V.n2021 VSS 0.056945f
C1461 ASIG5V.n2022 VSS 0.056945f
C1462 ASIG5V.n2023 VSS 0.056945f
C1463 ASIG5V.n2024 VSS 0.056945f
C1464 ASIG5V.n2025 VSS 0.056945f
C1465 ASIG5V.n2026 VSS 0.056945f
C1466 ASIG5V.n2027 VSS 0.056945f
C1467 ASIG5V.n2029 VSS 0.056945f
C1468 ASIG5V.n2030 VSS 0.056945f
C1469 ASIG5V.n2031 VSS 0.056945f
C1470 ASIG5V.n2033 VSS 0.056945f
C1471 ASIG5V.n2034 VSS 0.056945f
C1472 ASIG5V.n2035 VSS 0.056945f
C1473 ASIG5V.n2036 VSS 0.056945f
C1474 ASIG5V.n2037 VSS 0.056945f
C1475 ASIG5V.n2038 VSS 0.056945f
C1476 ASIG5V.n2039 VSS 0.056945f
C1477 ASIG5V.n2041 VSS 0.056945f
C1478 ASIG5V.n2042 VSS 0.056945f
C1479 ASIG5V.n2043 VSS 0.056945f
C1480 ASIG5V.n2045 VSS 0.056945f
C1481 ASIG5V.n2046 VSS 0.056945f
C1482 ASIG5V.n2047 VSS 0.056945f
C1483 ASIG5V.n2048 VSS 0.056945f
C1484 ASIG5V.n2049 VSS 0.056945f
C1485 ASIG5V.n2050 VSS 0.056945f
C1486 ASIG5V.n2051 VSS 0.056945f
C1487 ASIG5V.n2053 VSS 0.056945f
C1488 ASIG5V.n2054 VSS 0.056945f
C1489 ASIG5V.n2055 VSS 0.056945f
C1490 ASIG5V.n2057 VSS 0.056945f
C1491 ASIG5V.n2058 VSS 0.056945f
C1492 ASIG5V.n2059 VSS 0.056945f
C1493 ASIG5V.n2060 VSS 0.056945f
C1494 ASIG5V.n2061 VSS 0.056945f
C1495 ASIG5V.n2062 VSS 0.056945f
C1496 ASIG5V.n2063 VSS 0.056945f
C1497 ASIG5V.n2065 VSS 0.056945f
C1498 ASIG5V.n2066 VSS 0.056945f
C1499 ASIG5V.n2067 VSS 0.056945f
C1500 ASIG5V.n2069 VSS 0.056945f
C1501 ASIG5V.n2070 VSS 0.056945f
C1502 ASIG5V.n2071 VSS 0.056945f
C1503 ASIG5V.n2072 VSS 0.056945f
C1504 ASIG5V.n2073 VSS 0.056945f
C1505 ASIG5V.n2074 VSS 0.056945f
C1506 ASIG5V.n2075 VSS 0.056945f
C1507 ASIG5V.n2077 VSS 0.056945f
C1508 ASIG5V.n2078 VSS 0.056945f
C1509 ASIG5V.n2079 VSS 0.056945f
C1510 ASIG5V.n2081 VSS 0.056945f
C1511 ASIG5V.n2082 VSS 0.056945f
C1512 ASIG5V.n2083 VSS 0.056945f
C1513 ASIG5V.n2084 VSS 0.056945f
C1514 ASIG5V.n2085 VSS 0.056945f
C1515 ASIG5V.n2086 VSS 0.056945f
C1516 ASIG5V.n2087 VSS 0.056945f
C1517 ASIG5V.n2089 VSS 0.056945f
C1518 ASIG5V.n2090 VSS 0.056945f
C1519 ASIG5V.n2091 VSS 0.056945f
C1520 ASIG5V.n2093 VSS 0.056945f
C1521 ASIG5V.n2094 VSS 0.056945f
C1522 ASIG5V.n2095 VSS 0.056945f
C1523 ASIG5V.n2096 VSS 0.056945f
C1524 ASIG5V.n2097 VSS 0.056945f
C1525 ASIG5V.n2098 VSS 0.056945f
C1526 ASIG5V.n2099 VSS 0.056945f
C1527 ASIG5V.n2101 VSS 0.056945f
C1528 ASIG5V.n2102 VSS 0.056945f
C1529 ASIG5V.n2103 VSS 0.056945f
C1530 ASIG5V.n2105 VSS 0.056945f
C1531 ASIG5V.n2106 VSS 0.056945f
C1532 ASIG5V.n2107 VSS 0.056945f
C1533 ASIG5V.n2108 VSS 0.056945f
C1534 ASIG5V.n2109 VSS 0.056945f
C1535 ASIG5V.n2110 VSS 0.056945f
C1536 ASIG5V.n2111 VSS 0.056945f
C1537 ASIG5V.n2113 VSS 0.056945f
C1538 ASIG5V.n2114 VSS 0.056945f
C1539 ASIG5V.n2115 VSS 0.056945f
C1540 ASIG5V.n2117 VSS 0.056945f
C1541 ASIG5V.n2118 VSS 0.056945f
C1542 ASIG5V.n2119 VSS 0.056945f
C1543 ASIG5V.n2120 VSS 0.056945f
C1544 ASIG5V.n2121 VSS 0.056945f
C1545 ASIG5V.n2122 VSS 0.056945f
C1546 ASIG5V.n2123 VSS 0.056945f
C1547 ASIG5V.n2125 VSS 0.056945f
C1548 ASIG5V.n2126 VSS 0.056945f
C1549 ASIG5V.n2127 VSS 0.056945f
C1550 ASIG5V.n2129 VSS 0.056945f
C1551 ASIG5V.n2130 VSS 0.056945f
C1552 ASIG5V.n2131 VSS 0.056945f
C1553 ASIG5V.n2132 VSS 0.056945f
C1554 ASIG5V.n2133 VSS 0.056945f
C1555 ASIG5V.n2134 VSS 0.056945f
C1556 ASIG5V.n2135 VSS 0.056945f
C1557 ASIG5V.n2137 VSS 0.056945f
C1558 ASIG5V.n2138 VSS 0.056945f
C1559 ASIG5V.n2139 VSS 0.056945f
C1560 ASIG5V.n2141 VSS 0.056945f
C1561 ASIG5V.n2142 VSS 0.056945f
C1562 ASIG5V.n2143 VSS 0.056945f
C1563 ASIG5V.n2144 VSS 0.056945f
C1564 ASIG5V.n2145 VSS 0.056945f
C1565 ASIG5V.n2146 VSS 0.056945f
C1566 ASIG5V.n2147 VSS 0.056945f
C1567 ASIG5V.n2149 VSS 0.056945f
C1568 ASIG5V.n2150 VSS 0.056945f
C1569 ASIG5V.n2151 VSS 0.056945f
C1570 ASIG5V.n2153 VSS 0.056945f
C1571 ASIG5V.n2154 VSS 0.056945f
C1572 ASIG5V.n2155 VSS 0.056945f
C1573 ASIG5V.n2156 VSS 0.056945f
C1574 ASIG5V.n2157 VSS 0.056945f
C1575 ASIG5V.n2158 VSS 0.056945f
C1576 ASIG5V.n2159 VSS 0.056945f
C1577 ASIG5V.n2161 VSS 0.056945f
C1578 ASIG5V.n2162 VSS 0.056945f
C1579 ASIG5V.n2163 VSS 0.056945f
C1580 ASIG5V.n2165 VSS 0.056945f
C1581 ASIG5V.n2166 VSS 0.056945f
C1582 ASIG5V.n2167 VSS 0.056945f
C1583 ASIG5V.n2168 VSS 0.056945f
C1584 ASIG5V.n2169 VSS 0.056945f
C1585 ASIG5V.n2170 VSS 0.056945f
C1586 ASIG5V.n2171 VSS 0.056945f
C1587 ASIG5V.n2173 VSS 0.056945f
C1588 ASIG5V.n2174 VSS 0.056945f
C1589 ASIG5V.n2175 VSS 0.056945f
C1590 ASIG5V.n2177 VSS 0.056945f
C1591 ASIG5V.n2178 VSS 0.056945f
C1592 ASIG5V.n2179 VSS 0.056945f
C1593 ASIG5V.n2180 VSS 0.056945f
C1594 ASIG5V.n2181 VSS 0.056945f
C1595 ASIG5V.n2182 VSS 0.056945f
C1596 ASIG5V.n2183 VSS 0.056945f
C1597 ASIG5V.n2185 VSS 0.056945f
C1598 ASIG5V.n2186 VSS 0.056945f
C1599 ASIG5V.n2187 VSS 0.056945f
C1600 ASIG5V.n2189 VSS 0.056945f
C1601 ASIG5V.n2190 VSS 0.056945f
C1602 ASIG5V.n2191 VSS 0.056945f
C1603 ASIG5V.n2192 VSS 0.056945f
C1604 ASIG5V.n2193 VSS 0.056945f
C1605 ASIG5V.n2194 VSS 0.056945f
C1606 ASIG5V.n2195 VSS 0.056945f
C1607 ASIG5V.n2197 VSS 0.036092f
C1608 ASIG5V.n2198 VSS 0.809021f
C1609 ASIG5V.n2199 VSS 0.916891f
C1610 ASIG5V.n2200 VSS 0.462297f
C1611 ASIG5V.n2201 VSS 0.050509f
C1612 ASIG5V.n2202 VSS 0.050509f
C1613 ASIG5V.n2203 VSS 0.044113f
C1614 ASIG5V.n2204 VSS 0.052746f
C1615 ASIG5V.n2205 VSS 0.056379f
C1616 ASIG5V.n2206 VSS 0.047722f
C1617 ASIG5V.n2207 VSS 0.065343f
C1618 ASIG5V.n2208 VSS 0.045974f
C1619 ASIG5V.n2209 VSS 0.074818f
C1620 ASIG5V.n2210 VSS 0.045974f
C1621 ASIG5V.n2211 VSS 0.074818f
C1622 ASIG5V.n2212 VSS 0.408363f
C1623 ASIG5V.n2213 VSS 0.924595f
C1624 ASIG5V.n2214 VSS 0.093144f
C1625 ASIG5V.n2215 VSS 0.082599f
C1626 ASIG5V.n2216 VSS 0.093144f
C1627 ASIG5V.n2217 VSS 0.082599f
C1628 ASIG5V.n2218 VSS 0.052133f
C1629 ASIG5V.n2219 VSS 0.0621f
C1630 ASIG5V.n2220 VSS 0.0621f
C1631 ASIG5V.n2221 VSS 0.955416f
C1632 ASIG5V.n2263 VSS 0.036092f
C1633 ASIG5V.n2264 VSS 0.036092f
C1634 ASIG5V.n2265 VSS 0.056945f
C1635 ASIG5V.n2266 VSS 0.056945f
C1636 ASIG5V.n2267 VSS 0.056945f
C1637 ASIG5V.n2268 VSS 0.056945f
C1638 ASIG5V.n2269 VSS 0.056945f
C1639 ASIG5V.n2270 VSS 0.056945f
C1640 ASIG5V.n2271 VSS 0.056945f
C1641 ASIG5V.n2272 VSS 0.056945f
C1642 ASIG5V.n2273 VSS 0.056945f
C1643 ASIG5V.n2274 VSS 0.056945f
C1644 ASIG5V.n2275 VSS 0.056945f
C1645 ASIG5V.n2276 VSS 0.056945f
C1646 ASIG5V.n2277 VSS 0.056945f
C1647 ASIG5V.n2278 VSS 0.056945f
C1648 ASIG5V.n2279 VSS 0.056945f
C1649 ASIG5V.n2280 VSS 0.056945f
C1650 ASIG5V.n2281 VSS 0.056945f
C1651 ASIG5V.n2282 VSS 0.056945f
C1652 ASIG5V.n2283 VSS 0.056945f
C1653 ASIG5V.n2284 VSS 0.056945f
C1654 ASIG5V.n2285 VSS 0.056945f
C1655 ASIG5V.n2286 VSS 0.056945f
C1656 ASIG5V.n2287 VSS 0.056945f
C1657 ASIG5V.n2288 VSS 0.056945f
C1658 ASIG5V.n2289 VSS 0.056945f
C1659 ASIG5V.n2290 VSS 0.056945f
C1660 ASIG5V.n2291 VSS 0.056945f
C1661 ASIG5V.n2292 VSS 0.056945f
C1662 ASIG5V.n2293 VSS 0.056945f
C1663 ASIG5V.n2294 VSS 0.056945f
C1664 ASIG5V.n2295 VSS 0.056945f
C1665 ASIG5V.n2296 VSS 0.056945f
C1666 ASIG5V.n2297 VSS 0.056945f
C1667 ASIG5V.n2298 VSS 0.056945f
C1668 ASIG5V.n2299 VSS 0.056945f
C1669 ASIG5V.n2300 VSS 0.056945f
C1670 ASIG5V.n2301 VSS 0.056945f
C1671 ASIG5V.n2302 VSS 0.056945f
C1672 ASIG5V.n2303 VSS 0.056945f
C1673 ASIG5V.n2304 VSS 0.056945f
C1674 ASIG5V.n2305 VSS 0.036092f
C1675 ASIG5V.n2307 VSS 0.056945f
C1676 ASIG5V.n2308 VSS 0.056945f
C1677 ASIG5V.n2309 VSS 0.056945f
C1678 ASIG5V.n2310 VSS 0.056945f
C1679 ASIG5V.n2311 VSS 0.056945f
C1680 ASIG5V.n2312 VSS 0.056945f
C1681 ASIG5V.n2314 VSS 0.056945f
C1682 ASIG5V.n2315 VSS 0.056945f
C1683 ASIG5V.n2316 VSS 0.056945f
C1684 ASIG5V.n2318 VSS 0.056945f
C1685 ASIG5V.n2319 VSS 0.056945f
C1686 ASIG5V.n2320 VSS 0.056945f
C1687 ASIG5V.n2321 VSS 0.056945f
C1688 ASIG5V.n2322 VSS 0.056945f
C1689 ASIG5V.n2323 VSS 0.056945f
C1690 ASIG5V.n2324 VSS 0.056945f
C1691 ASIG5V.n2326 VSS 0.056945f
C1692 ASIG5V.n2327 VSS 0.056945f
C1693 ASIG5V.n2328 VSS 0.056945f
C1694 ASIG5V.n2330 VSS 0.056945f
C1695 ASIG5V.n2331 VSS 0.056945f
C1696 ASIG5V.n2332 VSS 0.056945f
C1697 ASIG5V.n2333 VSS 0.056945f
C1698 ASIG5V.n2334 VSS 0.056945f
C1699 ASIG5V.n2335 VSS 0.056945f
C1700 ASIG5V.n2336 VSS 0.056945f
C1701 ASIG5V.n2338 VSS 0.056945f
C1702 ASIG5V.n2339 VSS 0.056945f
C1703 ASIG5V.n2340 VSS 0.056945f
C1704 ASIG5V.n2342 VSS 0.056945f
C1705 ASIG5V.n2343 VSS 0.056945f
C1706 ASIG5V.n2344 VSS 0.056945f
C1707 ASIG5V.n2345 VSS 0.056945f
C1708 ASIG5V.n2346 VSS 0.056945f
C1709 ASIG5V.n2347 VSS 0.056945f
C1710 ASIG5V.n2348 VSS 0.056945f
C1711 ASIG5V.n2350 VSS 0.056945f
C1712 ASIG5V.n2351 VSS 0.056945f
C1713 ASIG5V.n2352 VSS 0.056945f
C1714 ASIG5V.n2354 VSS 0.056945f
C1715 ASIG5V.n2355 VSS 0.056945f
C1716 ASIG5V.n2356 VSS 0.056945f
C1717 ASIG5V.n2357 VSS 0.056945f
C1718 ASIG5V.n2358 VSS 0.056945f
C1719 ASIG5V.n2359 VSS 0.056945f
C1720 ASIG5V.n2360 VSS 0.056945f
C1721 ASIG5V.n2362 VSS 0.056945f
C1722 ASIG5V.n2363 VSS 0.056945f
C1723 ASIG5V.n2364 VSS 0.056945f
C1724 ASIG5V.n2366 VSS 0.056945f
C1725 ASIG5V.n2367 VSS 0.056945f
C1726 ASIG5V.n2368 VSS 0.056945f
C1727 ASIG5V.n2369 VSS 0.056945f
C1728 ASIG5V.n2370 VSS 0.056945f
C1729 ASIG5V.n2371 VSS 0.056945f
C1730 ASIG5V.n2372 VSS 0.056945f
C1731 ASIG5V.n2374 VSS 0.056945f
C1732 ASIG5V.n2375 VSS 0.056945f
C1733 ASIG5V.n2376 VSS 0.056945f
C1734 ASIG5V.n2378 VSS 0.056945f
C1735 ASIG5V.n2379 VSS 0.056945f
C1736 ASIG5V.n2380 VSS 0.056945f
C1737 ASIG5V.n2381 VSS 0.056945f
C1738 ASIG5V.n2382 VSS 0.056945f
C1739 ASIG5V.n2383 VSS 0.056945f
C1740 ASIG5V.n2384 VSS 0.056945f
C1741 ASIG5V.n2386 VSS 0.056945f
C1742 ASIG5V.n2387 VSS 0.056945f
C1743 ASIG5V.n2388 VSS 0.056945f
C1744 ASIG5V.n2390 VSS 0.056945f
C1745 ASIG5V.n2391 VSS 0.056945f
C1746 ASIG5V.n2392 VSS 0.056945f
C1747 ASIG5V.n2393 VSS 0.056945f
C1748 ASIG5V.n2394 VSS 0.056945f
C1749 ASIG5V.n2395 VSS 0.056945f
C1750 ASIG5V.n2396 VSS 0.056945f
C1751 ASIG5V.n2398 VSS 0.056945f
C1752 ASIG5V.n2399 VSS 0.056945f
C1753 ASIG5V.n2400 VSS 0.056945f
C1754 ASIG5V.n2402 VSS 0.056945f
C1755 ASIG5V.n2403 VSS 0.056945f
C1756 ASIG5V.n2404 VSS 0.056945f
C1757 ASIG5V.n2405 VSS 0.056945f
C1758 ASIG5V.n2406 VSS 0.056945f
C1759 ASIG5V.n2407 VSS 0.056945f
C1760 ASIG5V.n2408 VSS 0.056945f
C1761 ASIG5V.n2410 VSS 0.056945f
C1762 ASIG5V.n2411 VSS 0.056945f
C1763 ASIG5V.n2412 VSS 0.056945f
C1764 ASIG5V.n2414 VSS 0.056945f
C1765 ASIG5V.n2415 VSS 0.056945f
C1766 ASIG5V.n2416 VSS 0.056945f
C1767 ASIG5V.n2417 VSS 0.056945f
C1768 ASIG5V.n2418 VSS 0.056945f
C1769 ASIG5V.n2419 VSS 0.056945f
C1770 ASIG5V.n2420 VSS 0.056945f
C1771 ASIG5V.n2422 VSS 0.056945f
C1772 ASIG5V.n2423 VSS 0.056945f
C1773 ASIG5V.n2424 VSS 0.056945f
C1774 ASIG5V.n2426 VSS 0.056945f
C1775 ASIG5V.n2427 VSS 0.056945f
C1776 ASIG5V.n2428 VSS 0.056945f
C1777 ASIG5V.n2429 VSS 0.056945f
C1778 ASIG5V.n2430 VSS 0.056945f
C1779 ASIG5V.n2431 VSS 0.056945f
C1780 ASIG5V.n2432 VSS 0.056945f
C1781 ASIG5V.n2434 VSS 0.056945f
C1782 ASIG5V.n2435 VSS 0.056945f
C1783 ASIG5V.n2436 VSS 0.056945f
C1784 ASIG5V.n2438 VSS 0.056945f
C1785 ASIG5V.n2439 VSS 0.056945f
C1786 ASIG5V.n2440 VSS 0.056945f
C1787 ASIG5V.n2441 VSS 0.056945f
C1788 ASIG5V.n2442 VSS 0.056945f
C1789 ASIG5V.n2443 VSS 0.056945f
C1790 ASIG5V.n2444 VSS 0.056945f
C1791 ASIG5V.n2446 VSS 0.056945f
C1792 ASIG5V.n2447 VSS 0.056945f
C1793 ASIG5V.n2448 VSS 0.056945f
C1794 ASIG5V.n2450 VSS 0.056945f
C1795 ASIG5V.n2451 VSS 0.056945f
C1796 ASIG5V.n2452 VSS 0.056945f
C1797 ASIG5V.n2453 VSS 0.056945f
C1798 ASIG5V.n2454 VSS 0.056945f
C1799 ASIG5V.n2455 VSS 0.056945f
C1800 ASIG5V.n2456 VSS 0.056945f
C1801 ASIG5V.n2458 VSS 0.056945f
C1802 ASIG5V.n2459 VSS 0.056945f
C1803 ASIG5V.n2460 VSS 0.056945f
C1804 ASIG5V.n2462 VSS 0.056945f
C1805 ASIG5V.n2463 VSS 0.056945f
C1806 ASIG5V.n2464 VSS 0.056945f
C1807 ASIG5V.n2465 VSS 0.056945f
C1808 ASIG5V.n2466 VSS 0.056945f
C1809 ASIG5V.n2467 VSS 0.056945f
C1810 ASIG5V.n2468 VSS 0.056945f
C1811 ASIG5V.n2470 VSS 0.056945f
C1812 ASIG5V.n2471 VSS 0.056945f
C1813 ASIG5V.n2472 VSS 0.056945f
C1814 ASIG5V.n2474 VSS 0.056945f
C1815 ASIG5V.n2475 VSS 0.056945f
C1816 ASIG5V.n2476 VSS 0.056945f
C1817 ASIG5V.n2477 VSS 0.056945f
C1818 ASIG5V.n2478 VSS 0.056945f
C1819 ASIG5V.n2479 VSS 0.056945f
C1820 ASIG5V.n2480 VSS 0.056945f
C1821 ASIG5V.n2482 VSS 0.056945f
C1822 ASIG5V.n2483 VSS 0.056945f
C1823 ASIG5V.n2484 VSS 0.056945f
C1824 ASIG5V.n2486 VSS 0.056945f
C1825 ASIG5V.n2487 VSS 0.056945f
C1826 ASIG5V.n2488 VSS 0.056945f
C1827 ASIG5V.n2489 VSS 0.056945f
C1828 ASIG5V.n2490 VSS 0.056945f
C1829 ASIG5V.n2491 VSS 0.056945f
C1830 ASIG5V.n2492 VSS 0.056945f
C1831 ASIG5V.n2494 VSS 0.056945f
C1832 ASIG5V.n2495 VSS 0.056945f
C1833 ASIG5V.n2496 VSS 0.056945f
C1834 ASIG5V.n2498 VSS 0.056945f
C1835 ASIG5V.n2499 VSS 0.056945f
C1836 ASIG5V.n2500 VSS 0.056945f
C1837 ASIG5V.n2501 VSS 0.056945f
C1838 ASIG5V.n2502 VSS 0.056945f
C1839 ASIG5V.n2503 VSS 0.056945f
C1840 ASIG5V.n2504 VSS 0.056945f
C1841 ASIG5V.n2506 VSS 0.056945f
C1842 ASIG5V.n2507 VSS 0.056945f
C1843 ASIG5V.n2508 VSS 0.056945f
C1844 ASIG5V.n2510 VSS 0.056945f
C1845 ASIG5V.n2511 VSS 0.056945f
C1846 ASIG5V.n2512 VSS 0.056945f
C1847 ASIG5V.n2513 VSS 0.056945f
C1848 ASIG5V.n2514 VSS 0.056945f
C1849 ASIG5V.n2515 VSS 0.056945f
C1850 ASIG5V.n2516 VSS 0.056945f
C1851 ASIG5V.n2518 VSS 0.056945f
C1852 ASIG5V.n2519 VSS 0.056945f
C1853 ASIG5V.n2520 VSS 0.056945f
C1854 ASIG5V.n2522 VSS 0.056945f
C1855 ASIG5V.n2523 VSS 0.056945f
C1856 ASIG5V.n2524 VSS 0.056945f
C1857 ASIG5V.n2525 VSS 0.056945f
C1858 ASIG5V.n2526 VSS 0.056945f
C1859 ASIG5V.n2527 VSS 0.056945f
C1860 ASIG5V.n2528 VSS 0.056945f
C1861 ASIG5V.n2530 VSS 0.056945f
C1862 ASIG5V.n2531 VSS 0.056945f
C1863 ASIG5V.n2532 VSS 0.056945f
C1864 ASIG5V.n2534 VSS 0.056945f
C1865 ASIG5V.n2535 VSS 0.056945f
C1866 ASIG5V.n2536 VSS 0.056945f
C1867 ASIG5V.n2537 VSS 0.056945f
C1868 ASIG5V.n2538 VSS 0.056945f
C1869 ASIG5V.n2539 VSS 0.056945f
C1870 ASIG5V.n2540 VSS 0.056945f
C1871 ASIG5V.n2542 VSS 0.056945f
C1872 ASIG5V.n2543 VSS 0.056945f
C1873 ASIG5V.n2544 VSS 0.056945f
C1874 ASIG5V.n2546 VSS 0.056945f
C1875 ASIG5V.n2547 VSS 0.056945f
C1876 ASIG5V.n2548 VSS 0.056945f
C1877 ASIG5V.n2549 VSS 0.056945f
C1878 ASIG5V.n2550 VSS 0.056945f
C1879 ASIG5V.n2551 VSS 0.056945f
C1880 ASIG5V.n2552 VSS 0.056945f
C1881 ASIG5V.n2554 VSS 0.036092f
C1882 ASIG5V.n2555 VSS 0.824431f
C1883 ASIG5V.n2556 VSS 0.816725f
C1884 ASIG5V.n2557 VSS 0.408363f
C1885 ASIG5V.n2558 VSS 0.070297f
C1886 ASIG5V.n2559 VSS 0.070297f
C1887 ASIG5V.n2560 VSS 0.062748f
C1888 ASIG5V.n2561 VSS 0.07229f
C1889 ASIG5V.n2562 VSS 0.083142f
C1890 ASIG5V.n2563 VSS 0.052133f
C1891 ASIG5V.n2564 VSS 0.06118f
C1892 ASIG5V.n2565 VSS 0.0621f
C1893 ASIG5V.n2566 VSS 0.108961f
C1894 ASIG5V.n2567 VSS 0.0621f
C1895 ASIG5V.n2568 VSS 0.108961f
C1896 ASIG5V.n2569 VSS 0.955415f
C1897 ASIG5V.n2611 VSS 0.036092f
C1898 ASIG5V.n2612 VSS 0.847545f
C1899 ASIG5V.n2613 VSS 0.045974f
C1900 ASIG5V.n2614 VSS 0.036092f
C1901 ASIG5V.n2615 VSS 0.577872f
C1902 ASIG5V.n2616 VSS 0.547052f
C1903 ASIG5V.n2617 VSS 0.056945f
C1904 ASIG5V.n2618 VSS 0.056945f
C1905 ASIG5V.n2619 VSS 0.056945f
C1906 ASIG5V.n2620 VSS 0.056945f
C1907 ASIG5V.n2621 VSS 0.056945f
C1908 ASIG5V.n2622 VSS 0.056945f
C1909 ASIG5V.n2623 VSS 0.056945f
C1910 ASIG5V.n2624 VSS 0.056945f
C1911 ASIG5V.n2625 VSS 0.056945f
C1912 ASIG5V.n2626 VSS 0.056945f
C1913 ASIG5V.n2627 VSS 0.056945f
C1914 ASIG5V.n2628 VSS 0.056945f
C1915 ASIG5V.n2629 VSS 0.056945f
C1916 ASIG5V.n2630 VSS 0.056945f
C1917 ASIG5V.n2631 VSS 0.056945f
C1918 ASIG5V.n2632 VSS 0.056945f
C1919 ASIG5V.n2633 VSS 0.056945f
C1920 ASIG5V.n2634 VSS 0.056945f
C1921 ASIG5V.n2635 VSS 0.056945f
C1922 ASIG5V.n2636 VSS 0.056945f
C1923 ASIG5V.n2637 VSS 0.056945f
C1924 ASIG5V.n2638 VSS 0.056945f
C1925 ASIG5V.n2639 VSS 0.056945f
C1926 ASIG5V.n2640 VSS 0.056945f
C1927 ASIG5V.n2641 VSS 0.056945f
C1928 ASIG5V.n2642 VSS 0.056945f
C1929 ASIG5V.n2643 VSS 0.056945f
C1930 ASIG5V.n2644 VSS 0.056945f
C1931 ASIG5V.n2645 VSS 0.056945f
C1932 ASIG5V.n2646 VSS 0.056945f
C1933 ASIG5V.n2647 VSS 0.056945f
C1934 ASIG5V.n2648 VSS 0.056945f
C1935 ASIG5V.n2649 VSS 0.056945f
C1936 ASIG5V.n2650 VSS 0.056945f
C1937 ASIG5V.n2651 VSS 0.056945f
C1938 ASIG5V.n2652 VSS 0.056945f
C1939 ASIG5V.n2653 VSS 0.056945f
C1940 ASIG5V.n2654 VSS 0.056945f
C1941 ASIG5V.n2655 VSS 0.056945f
C1942 ASIG5V.n2656 VSS 0.056945f
C1943 ASIG5V.n2657 VSS 0.036092f
C1944 ASIG5V.n2659 VSS 0.056945f
C1945 ASIG5V.n2660 VSS 0.056945f
C1946 ASIG5V.n2661 VSS 0.056945f
C1947 ASIG5V.n2662 VSS 0.056945f
C1948 ASIG5V.n2663 VSS 0.056945f
C1949 ASIG5V.n2664 VSS 0.056945f
C1950 ASIG5V.n2666 VSS 0.056945f
C1951 ASIG5V.n2667 VSS 0.056945f
C1952 ASIG5V.n2668 VSS 0.056945f
C1953 ASIG5V.n2670 VSS 0.056945f
C1954 ASIG5V.n2671 VSS 0.056945f
C1955 ASIG5V.n2672 VSS 0.056945f
C1956 ASIG5V.n2673 VSS 0.056945f
C1957 ASIG5V.n2674 VSS 0.056945f
C1958 ASIG5V.n2675 VSS 0.056945f
C1959 ASIG5V.n2676 VSS 0.056945f
C1960 ASIG5V.n2678 VSS 0.056945f
C1961 ASIG5V.n2679 VSS 0.056945f
C1962 ASIG5V.n2680 VSS 0.056945f
C1963 ASIG5V.n2682 VSS 0.056945f
C1964 ASIG5V.n2683 VSS 0.056945f
C1965 ASIG5V.n2684 VSS 0.056945f
C1966 ASIG5V.n2685 VSS 0.056945f
C1967 ASIG5V.n2686 VSS 0.056945f
C1968 ASIG5V.n2687 VSS 0.056945f
C1969 ASIG5V.n2688 VSS 0.056945f
C1970 ASIG5V.n2690 VSS 0.056945f
C1971 ASIG5V.n2691 VSS 0.056945f
C1972 ASIG5V.n2692 VSS 0.056945f
C1973 ASIG5V.n2694 VSS 0.056945f
C1974 ASIG5V.n2695 VSS 0.056945f
C1975 ASIG5V.n2696 VSS 0.056945f
C1976 ASIG5V.n2697 VSS 0.056945f
C1977 ASIG5V.n2698 VSS 0.056945f
C1978 ASIG5V.n2699 VSS 0.056945f
C1979 ASIG5V.n2700 VSS 0.056945f
C1980 ASIG5V.n2702 VSS 0.056945f
C1981 ASIG5V.n2703 VSS 0.056945f
C1982 ASIG5V.n2704 VSS 0.056945f
C1983 ASIG5V.n2706 VSS 0.056945f
C1984 ASIG5V.n2707 VSS 0.056945f
C1985 ASIG5V.n2708 VSS 0.056945f
C1986 ASIG5V.n2709 VSS 0.056945f
C1987 ASIG5V.n2710 VSS 0.056945f
C1988 ASIG5V.n2711 VSS 0.056945f
C1989 ASIG5V.n2712 VSS 0.056945f
C1990 ASIG5V.n2714 VSS 0.056945f
C1991 ASIG5V.n2715 VSS 0.056945f
C1992 ASIG5V.n2716 VSS 0.056945f
C1993 ASIG5V.n2718 VSS 0.056945f
C1994 ASIG5V.n2719 VSS 0.056945f
C1995 ASIG5V.n2720 VSS 0.056945f
C1996 ASIG5V.n2721 VSS 0.056945f
C1997 ASIG5V.n2722 VSS 0.056945f
C1998 ASIG5V.n2723 VSS 0.056945f
C1999 ASIG5V.n2724 VSS 0.056945f
C2000 ASIG5V.n2726 VSS 0.056945f
C2001 ASIG5V.n2727 VSS 0.056945f
C2002 ASIG5V.n2728 VSS 0.056945f
C2003 ASIG5V.n2730 VSS 0.056945f
C2004 ASIG5V.n2731 VSS 0.056945f
C2005 ASIG5V.n2732 VSS 0.056945f
C2006 ASIG5V.n2733 VSS 0.056945f
C2007 ASIG5V.n2734 VSS 0.056945f
C2008 ASIG5V.n2735 VSS 0.056945f
C2009 ASIG5V.n2736 VSS 0.056945f
C2010 ASIG5V.n2738 VSS 0.056945f
C2011 ASIG5V.n2739 VSS 0.056945f
C2012 ASIG5V.n2740 VSS 0.056945f
C2013 ASIG5V.n2742 VSS 0.056945f
C2014 ASIG5V.n2743 VSS 0.056945f
C2015 ASIG5V.n2744 VSS 0.056945f
C2016 ASIG5V.n2745 VSS 0.056945f
C2017 ASIG5V.n2746 VSS 0.056945f
C2018 ASIG5V.n2747 VSS 0.056945f
C2019 ASIG5V.n2748 VSS 0.056945f
C2020 ASIG5V.n2750 VSS 0.056945f
C2021 ASIG5V.n2751 VSS 0.056945f
C2022 ASIG5V.n2752 VSS 0.056945f
C2023 ASIG5V.n2754 VSS 0.056945f
C2024 ASIG5V.n2755 VSS 0.056945f
C2025 ASIG5V.n2756 VSS 0.056945f
C2026 ASIG5V.n2757 VSS 0.056945f
C2027 ASIG5V.n2758 VSS 0.056945f
C2028 ASIG5V.n2759 VSS 0.056945f
C2029 ASIG5V.n2760 VSS 0.056945f
C2030 ASIG5V.n2762 VSS 0.056945f
C2031 ASIG5V.n2763 VSS 0.056945f
C2032 ASIG5V.n2764 VSS 0.056945f
C2033 ASIG5V.n2766 VSS 0.056945f
C2034 ASIG5V.n2767 VSS 0.056945f
C2035 ASIG5V.n2768 VSS 0.056945f
C2036 ASIG5V.n2769 VSS 0.056945f
C2037 ASIG5V.n2770 VSS 0.056945f
C2038 ASIG5V.n2771 VSS 0.056945f
C2039 ASIG5V.n2772 VSS 0.056945f
C2040 ASIG5V.n2774 VSS 0.056945f
C2041 ASIG5V.n2775 VSS 0.056945f
C2042 ASIG5V.n2776 VSS 0.056945f
C2043 ASIG5V.n2778 VSS 0.056945f
C2044 ASIG5V.n2779 VSS 0.056945f
C2045 ASIG5V.n2780 VSS 0.056945f
C2046 ASIG5V.n2781 VSS 0.056945f
C2047 ASIG5V.n2782 VSS 0.056945f
C2048 ASIG5V.n2783 VSS 0.056945f
C2049 ASIG5V.n2784 VSS 0.056945f
C2050 ASIG5V.n2786 VSS 0.056945f
C2051 ASIG5V.n2787 VSS 0.056945f
C2052 ASIG5V.n2788 VSS 0.056945f
C2053 ASIG5V.n2790 VSS 0.056945f
C2054 ASIG5V.n2791 VSS 0.056945f
C2055 ASIG5V.n2792 VSS 0.056945f
C2056 ASIG5V.n2793 VSS 0.056945f
C2057 ASIG5V.n2794 VSS 0.056945f
C2058 ASIG5V.n2795 VSS 0.056945f
C2059 ASIG5V.n2796 VSS 0.056945f
C2060 ASIG5V.n2798 VSS 0.056945f
C2061 ASIG5V.n2799 VSS 0.056945f
C2062 ASIG5V.n2800 VSS 0.056945f
C2063 ASIG5V.n2802 VSS 0.056945f
C2064 ASIG5V.n2803 VSS 0.056945f
C2065 ASIG5V.n2804 VSS 0.056945f
C2066 ASIG5V.n2805 VSS 0.056945f
C2067 ASIG5V.n2806 VSS 0.056945f
C2068 ASIG5V.n2807 VSS 0.056945f
C2069 ASIG5V.n2808 VSS 0.056945f
C2070 ASIG5V.n2810 VSS 0.056945f
C2071 ASIG5V.n2811 VSS 0.056945f
C2072 ASIG5V.n2812 VSS 0.056945f
C2073 ASIG5V.n2814 VSS 0.056945f
C2074 ASIG5V.n2815 VSS 0.056945f
C2075 ASIG5V.n2816 VSS 0.056945f
C2076 ASIG5V.n2817 VSS 0.056945f
C2077 ASIG5V.n2818 VSS 0.056945f
C2078 ASIG5V.n2819 VSS 0.056945f
C2079 ASIG5V.n2820 VSS 0.056945f
C2080 ASIG5V.n2822 VSS 0.056945f
C2081 ASIG5V.n2823 VSS 0.056945f
C2082 ASIG5V.n2824 VSS 0.056945f
C2083 ASIG5V.n2826 VSS 0.056945f
C2084 ASIG5V.n2827 VSS 0.056945f
C2085 ASIG5V.n2828 VSS 0.056945f
C2086 ASIG5V.n2829 VSS 0.056945f
C2087 ASIG5V.n2830 VSS 0.056945f
C2088 ASIG5V.n2831 VSS 0.056945f
C2089 ASIG5V.n2832 VSS 0.056945f
C2090 ASIG5V.n2834 VSS 0.056945f
C2091 ASIG5V.n2835 VSS 0.056945f
C2092 ASIG5V.n2836 VSS 0.056945f
C2093 ASIG5V.n2838 VSS 0.056945f
C2094 ASIG5V.n2839 VSS 0.056945f
C2095 ASIG5V.n2840 VSS 0.056945f
C2096 ASIG5V.n2841 VSS 0.056945f
C2097 ASIG5V.n2842 VSS 0.056945f
C2098 ASIG5V.n2843 VSS 0.056945f
C2099 ASIG5V.n2844 VSS 0.056945f
C2100 ASIG5V.n2846 VSS 0.056945f
C2101 ASIG5V.n2847 VSS 0.056945f
C2102 ASIG5V.n2848 VSS 0.056945f
C2103 ASIG5V.n2850 VSS 0.056945f
C2104 ASIG5V.n2851 VSS 0.056945f
C2105 ASIG5V.n2852 VSS 0.056945f
C2106 ASIG5V.n2853 VSS 0.056945f
C2107 ASIG5V.n2854 VSS 0.056945f
C2108 ASIG5V.n2855 VSS 0.056945f
C2109 ASIG5V.n2856 VSS 0.056945f
C2110 ASIG5V.n2858 VSS 0.056945f
C2111 ASIG5V.n2859 VSS 0.056945f
C2112 ASIG5V.n2860 VSS 0.056945f
C2113 ASIG5V.n2862 VSS 0.056945f
C2114 ASIG5V.n2863 VSS 0.056945f
C2115 ASIG5V.n2864 VSS 0.056945f
C2116 ASIG5V.n2865 VSS 0.056945f
C2117 ASIG5V.n2866 VSS 0.056945f
C2118 ASIG5V.n2867 VSS 0.056945f
C2119 ASIG5V.n2868 VSS 0.056945f
C2120 ASIG5V.n2870 VSS 0.056945f
C2121 ASIG5V.n2871 VSS 0.056945f
C2122 ASIG5V.n2872 VSS 0.056945f
C2123 ASIG5V.n2874 VSS 0.056945f
C2124 ASIG5V.n2875 VSS 0.056945f
C2125 ASIG5V.n2876 VSS 0.056945f
C2126 ASIG5V.n2877 VSS 0.056945f
C2127 ASIG5V.n2878 VSS 0.056945f
C2128 ASIG5V.n2879 VSS 0.056945f
C2129 ASIG5V.n2880 VSS 0.056945f
C2130 ASIG5V.n2882 VSS 0.056945f
C2131 ASIG5V.n2883 VSS 0.056945f
C2132 ASIG5V.n2884 VSS 0.056945f
C2133 ASIG5V.n2886 VSS 0.056945f
C2134 ASIG5V.n2887 VSS 0.056945f
C2135 ASIG5V.n2888 VSS 0.056945f
C2136 ASIG5V.n2889 VSS 0.056945f
C2137 ASIG5V.n2890 VSS 0.056945f
C2138 ASIG5V.n2891 VSS 0.056945f
C2139 ASIG5V.n2892 VSS 0.056945f
C2140 ASIG5V.n2894 VSS 0.056945f
C2141 ASIG5V.n2895 VSS 0.056945f
C2142 ASIG5V.n2896 VSS 0.056945f
C2143 ASIG5V.n2898 VSS 0.056945f
C2144 ASIG5V.n2899 VSS 0.056945f
C2145 ASIG5V.n2900 VSS 0.056945f
C2146 ASIG5V.n2901 VSS 0.056945f
C2147 ASIG5V.n2902 VSS 0.066995f
C2148 ASIG5V.n2903 VSS 0.045974f
C2149 ASIG5V.n2904 VSS 0.076709f
C2150 ASIG5V.n2905 VSS 0.045974f
C2151 ASIG5V.n2906 VSS 1.0941f
C2152 ASIG5V.n2907 VSS 0.955415f
C2153 ASIG5V.n2908 VSS 0.045974f
C2154 ASIG5V.n2909 VSS 0.047722f
C2155 ASIG5V.n2910 VSS 0.066995f
C2156 ASIG5V.n2911 VSS 0.076709f
C2157 ASIG5V.n2912 VSS 0.076709f
C2158 ASIG5V.n2913 VSS 0.801315f
C2159 ASIG5V.n2955 VSS 0.036092f
C2160 ASIG5V.n2956 VSS 0.801315f
C2161 ASIG5V.n2957 VSS 0.036092f
C2162 ASIG5V.n2958 VSS 0.955415f
C2163 ASIG5V.n2959 VSS 0.056945f
C2164 ASIG5V.n2960 VSS 0.056945f
C2165 ASIG5V.n2961 VSS 0.056945f
C2166 ASIG5V.n2962 VSS 0.056945f
C2167 ASIG5V.n2963 VSS 0.056945f
C2168 ASIG5V.n2964 VSS 0.056945f
C2169 ASIG5V.n2965 VSS 0.056945f
C2170 ASIG5V.n2966 VSS 0.056945f
C2171 ASIG5V.n2967 VSS 0.056945f
C2172 ASIG5V.n2968 VSS 0.056945f
C2173 ASIG5V.n2969 VSS 0.056945f
C2174 ASIG5V.n2970 VSS 0.056945f
C2175 ASIG5V.n2971 VSS 0.056945f
C2176 ASIG5V.n2972 VSS 0.056945f
C2177 ASIG5V.n2973 VSS 0.056945f
C2178 ASIG5V.n2974 VSS 0.056945f
C2179 ASIG5V.n2975 VSS 0.056945f
C2180 ASIG5V.n2976 VSS 0.056945f
C2181 ASIG5V.n2977 VSS 0.056945f
C2182 ASIG5V.n2978 VSS 0.056945f
C2183 ASIG5V.n2979 VSS 0.056945f
C2184 ASIG5V.n2980 VSS 0.056945f
C2185 ASIG5V.n2981 VSS 0.056945f
C2186 ASIG5V.n2982 VSS 0.056945f
C2187 ASIG5V.n2983 VSS 0.056945f
C2188 ASIG5V.n2984 VSS 0.056945f
C2189 ASIG5V.n2985 VSS 0.056945f
C2190 ASIG5V.n2986 VSS 0.056945f
C2191 ASIG5V.n2987 VSS 0.056945f
C2192 ASIG5V.n2988 VSS 0.056945f
C2193 ASIG5V.n2989 VSS 0.056945f
C2194 ASIG5V.n2990 VSS 0.056945f
C2195 ASIG5V.n2991 VSS 0.056945f
C2196 ASIG5V.n2992 VSS 0.056945f
C2197 ASIG5V.n2993 VSS 0.056945f
C2198 ASIG5V.n2994 VSS 0.056945f
C2199 ASIG5V.n2995 VSS 0.056945f
C2200 ASIG5V.n2996 VSS 0.056945f
C2201 ASIG5V.n2997 VSS 0.056945f
C2202 ASIG5V.n2998 VSS 0.056945f
C2203 ASIG5V.n3000 VSS 0.056945f
C2204 ASIG5V.n3001 VSS 0.056945f
C2205 ASIG5V.n3002 VSS 0.07229f
C2206 ASIG5V.n3004 VSS 0.493967f
C2207 ASIG5V.n3005 VSS 0.087753f
C2208 ASIG5V.n3006 VSS 0.074298f
C2209 ASIG5V.n3008 VSS 0.074298f
C2210 ASIG5V.n3009 VSS 0.314214f
C2211 ASIG5V.n3012 VSS 0.314214f
C2212 ASIG5V.n3013 VSS 0.074298f
C2213 ASIG5V.n3015 VSS 0.074298f
C2214 ASIG5V.n3018 VSS 0.087753f
C2215 ASIG5V.n3019 VSS 0.087753f
C2216 ASIG5V.n3023 VSS 0.314214f
C2217 ASIG5V.n3024 VSS 0.074298f
C2218 ASIG5V.n3026 VSS 0.074298f
C2219 ASIG5V.n3029 VSS 0.087753f
C2220 ASIG5V.n3030 VSS 0.087753f
C2221 ASIG5V.n3034 VSS 0.314214f
C2222 ASIG5V.n3035 VSS 0.074298f
C2223 ASIG5V.n3037 VSS 0.074298f
C2224 ASIG5V.n3040 VSS 0.087753f
C2225 ASIG5V.n3041 VSS 0.087753f
C2226 ASIG5V.n3045 VSS 0.314214f
C2227 ASIG5V.n3046 VSS 0.074298f
C2228 ASIG5V.n3048 VSS 0.074298f
C2229 ASIG5V.n3051 VSS 0.087753f
C2230 ASIG5V.n3052 VSS 0.087753f
C2231 ASIG5V.n3056 VSS 0.314214f
C2232 ASIG5V.n3057 VSS 0.074298f
C2233 ASIG5V.n3059 VSS 0.074298f
C2234 ASIG5V.n3062 VSS 0.087753f
C2235 ASIG5V.n3063 VSS 0.087753f
C2236 ASIG5V.n3067 VSS 0.314214f
C2237 ASIG5V.n3068 VSS 0.074298f
C2238 ASIG5V.n3070 VSS 0.074298f
C2239 ASIG5V.n3073 VSS 0.087753f
C2240 ASIG5V.n3074 VSS 0.087753f
C2241 ASIG5V.n3079 VSS 0.074298f
C2242 ASIG5V.n3080 VSS 0.074298f
C2243 ASIG5V.n3081 VSS 12.9443f
C2244 ASIG5V.n3083 VSS 0.309175f
C2245 ASIG5V.n3086 VSS 0.074298f
C2246 ASIG5V.n3087 VSS 12.9443f
C2247 ASIG5V.n3088 VSS 0.309175f
C2248 ASIG5V.n3091 VSS 0.087753f
C2249 ASIG5V.n3093 VSS 0.074298f
C2250 ASIG5V.n3094 VSS 12.9443f
C2251 ASIG5V.n3095 VSS 0.309175f
C2252 ASIG5V.n3098 VSS 0.087753f
C2253 ASIG5V.n3100 VSS 0.074298f
C2254 ASIG5V.n3101 VSS 12.9443f
C2255 ASIG5V.n3102 VSS 0.309175f
C2256 ASIG5V.n3105 VSS 0.087753f
C2257 ASIG5V.n3107 VSS 0.074298f
C2258 ASIG5V.n3108 VSS 12.9443f
C2259 ASIG5V.n3109 VSS 0.309175f
C2260 ASIG5V.n3112 VSS 0.087753f
C2261 ASIG5V.n3114 VSS 0.074298f
C2262 ASIG5V.n3115 VSS 12.9443f
C2263 ASIG5V.n3116 VSS 0.309175f
C2264 ASIG5V.n3119 VSS 0.087753f
C2265 ASIG5V.n3121 VSS 0.074298f
C2266 ASIG5V.n3122 VSS 12.9443f
C2267 ASIG5V.n3126 VSS 0.074298f
C2268 ASIG5V.n3127 VSS 0.314214f
C2269 ASIG5V.n3131 VSS 0.074298f
C2270 ASIG5V.n3132 VSS 0.314214f
C2271 ASIG5V.n3136 VSS 0.074298f
C2272 ASIG5V.n3137 VSS 0.314214f
C2273 ASIG5V.n3141 VSS 0.074298f
C2274 ASIG5V.n3142 VSS 0.314214f
C2275 ASIG5V.n3146 VSS 0.074298f
C2276 ASIG5V.n3147 VSS 0.314214f
C2277 ASIG5V.n3151 VSS 0.074298f
C2278 ASIG5V.n3152 VSS 0.074298f
C2279 ASIG5V.n3153 VSS 0.314214f
C2280 ASIG5V.n3157 VSS 0.074298f
C2281 ASIG5V.n3158 VSS 0.074298f
C2282 ASIG5V.n3159 VSS 0.087753f
C2283 ASIG5V.n3161 VSS 0.074298f
C2284 ASIG5V.n3163 VSS 0.090985f
C2285 ASIG5V.n3164 VSS 0.120921f
C2286 ASIG5V.n3165 VSS 0.108961f
C2287 ASIG5V.n3166 VSS 0.11658f
C2288 ASIG5V.n3167 VSS 0.108961f
C2289 ASIG5V.n3168 VSS 0.11658f
C2290 ASIG5V.n3169 VSS 0.955415f
C2291 ASIG5V.n3170 VSS 0.670332f
C2292 ASIG5V.n3171 VSS 0.076709f
C2293 ASIG5V.n3172 VSS 0.045974f
C2294 ASIG5V.n3173 VSS 0.076709f
C2295 ASIG5V.n3174 VSS 0.045974f
C2296 ASIG5V.n3175 VSS 0.052746f
C2297 ASIG5V.n3176 VSS 0.045974f
C2298 ASIG5V.n3177 VSS 0.045974f
C2299 ASIG5V.n3178 VSS 0.708856f
C2300 ASIG5V.n3220 VSS 0.036092f
C2301 ASIG5V.n3221 VSS 0.708856f
C2302 ASIG5V.n3222 VSS 0.036092f
C2303 ASIG5V.n3223 VSS 0.955415f
C2304 ASIG5V.n3224 VSS 0.056945f
C2305 ASIG5V.n3225 VSS 0.056945f
C2306 ASIG5V.n3226 VSS 0.056945f
C2307 ASIG5V.n3227 VSS 0.056945f
C2308 ASIG5V.n3228 VSS 0.056945f
C2309 ASIG5V.n3229 VSS 0.056945f
C2310 ASIG5V.n3230 VSS 0.056945f
C2311 ASIG5V.n3231 VSS 0.056945f
C2312 ASIG5V.n3232 VSS 0.056945f
C2313 ASIG5V.n3233 VSS 0.056945f
C2314 ASIG5V.n3234 VSS 0.056945f
C2315 ASIG5V.n3235 VSS 0.056945f
C2316 ASIG5V.n3236 VSS 0.056945f
C2317 ASIG5V.n3237 VSS 0.056945f
C2318 ASIG5V.n3238 VSS 0.056945f
C2319 ASIG5V.n3239 VSS 0.056945f
C2320 ASIG5V.n3240 VSS 0.056945f
C2321 ASIG5V.n3241 VSS 0.056945f
C2322 ASIG5V.n3242 VSS 0.056945f
C2323 ASIG5V.n3243 VSS 0.056945f
C2324 ASIG5V.n3244 VSS 0.056945f
C2325 ASIG5V.n3245 VSS 0.056945f
C2326 ASIG5V.n3246 VSS 0.056945f
C2327 ASIG5V.n3247 VSS 0.056945f
C2328 ASIG5V.n3248 VSS 0.056945f
C2329 ASIG5V.n3249 VSS 0.056945f
C2330 ASIG5V.n3250 VSS 0.056945f
C2331 ASIG5V.n3251 VSS 0.056945f
C2332 ASIG5V.n3252 VSS 0.056945f
C2333 ASIG5V.n3253 VSS 0.056945f
C2334 ASIG5V.n3254 VSS 0.056945f
C2335 ASIG5V.n3255 VSS 0.056945f
C2336 ASIG5V.n3256 VSS 0.056945f
C2337 ASIG5V.n3257 VSS 0.056945f
C2338 ASIG5V.n3258 VSS 0.056945f
C2339 ASIG5V.n3259 VSS 0.056945f
C2340 ASIG5V.n3260 VSS 0.056945f
C2341 ASIG5V.n3261 VSS 0.056945f
C2342 ASIG5V.n3262 VSS 0.056945f
C2343 ASIG5V.n3263 VSS 0.056945f
C2344 ASIG5V.n3265 VSS 0.056945f
C2345 ASIG5V.n3266 VSS 0.056945f
C2346 ASIG5V.n3267 VSS 0.07229f
C2347 ASIG5V.n3268 VSS 0.096659f
C2348 ASIG5V.n3269 VSS 0.108961f
C2349 ASIG5V.n3270 VSS 1.0941f
C2350 ASIG5V.n3271 VSS 0.076709f
C2351 ASIG5V.n3272 VSS 0.076709f
C2352 ASIG5V.n3273 VSS 0.052746f
C2353 ASIG5V.n3274 VSS 0.045974f
C2354 ASIG5V.n3275 VSS 0.045974f
C2355 ASIG5V.n3276 VSS 1.0941f
C2356 ASIG5V.n3277 VSS 0.816725f
C2357 ASIG5V.n3278 VSS 0.685742f
C2358 ASIG5V.n3279 VSS 0.0621f
C2359 ASIG5V.n3280 VSS 0.0621f
C2360 ASIG5V.n3281 VSS 0.108961f
C2361 ASIG5V.n3282 VSS 0.056945f
C2362 ASIG5V.n3283 VSS 0.056945f
C2363 ASIG5V.n3285 VSS 0.056945f
C2364 ASIG5V.n3286 VSS 0.056945f
C2365 ASIG5V.n3287 VSS 0.056945f
C2366 ASIG5V.n3288 VSS 0.056945f
C2367 ASIG5V.n3291 VSS 0.056945f
C2368 ASIG5V.n3292 VSS 0.056945f
C2369 ASIG5V.n3293 VSS 0.056945f
C2370 ASIG5V.n3294 VSS 0.056945f
C2371 ASIG5V.n3297 VSS 0.056945f
C2372 ASIG5V.n3298 VSS 0.056945f
C2373 ASIG5V.n3299 VSS 0.056945f
C2374 ASIG5V.n3300 VSS 0.056945f
C2375 ASIG5V.n3303 VSS 0.056945f
C2376 ASIG5V.n3304 VSS 0.056945f
C2377 ASIG5V.n3305 VSS 0.056945f
C2378 ASIG5V.n3306 VSS 0.056945f
C2379 ASIG5V.n3309 VSS 0.056945f
C2380 ASIG5V.n3310 VSS 0.056945f
C2381 ASIG5V.n3311 VSS 0.056945f
C2382 ASIG5V.n3312 VSS 0.056945f
C2383 ASIG5V.n3315 VSS 0.056945f
C2384 ASIG5V.n3316 VSS 0.056945f
C2385 ASIG5V.n3317 VSS 0.056945f
C2386 ASIG5V.n3318 VSS 0.056945f
C2387 ASIG5V.n3321 VSS 0.056945f
C2388 ASIG5V.n3322 VSS 0.056945f
C2389 ASIG5V.n3323 VSS 0.056945f
C2390 ASIG5V.n3324 VSS 0.056945f
C2391 ASIG5V.n3327 VSS 0.056945f
C2392 ASIG5V.n3328 VSS 0.056945f
C2393 ASIG5V.n3329 VSS 0.056945f
C2394 ASIG5V.n3330 VSS 0.056945f
C2395 ASIG5V.n3333 VSS 0.056945f
C2396 ASIG5V.n3334 VSS 0.056945f
C2397 ASIG5V.n3335 VSS 0.056945f
C2398 ASIG5V.n3336 VSS 0.056945f
C2399 ASIG5V.n3339 VSS 0.056945f
C2400 ASIG5V.n3340 VSS 0.056945f
C2401 ASIG5V.n3341 VSS 0.056945f
C2402 ASIG5V.n3342 VSS 0.056945f
C2403 ASIG5V.n3345 VSS 0.056945f
C2404 ASIG5V.n3346 VSS 0.056945f
C2405 ASIG5V.n3347 VSS 0.056945f
C2406 ASIG5V.n3348 VSS 0.056945f
C2407 ASIG5V.n3351 VSS 0.056945f
C2408 ASIG5V.n3352 VSS 0.056945f
C2409 ASIG5V.n3353 VSS 0.056945f
C2410 ASIG5V.n3354 VSS 0.056945f
C2411 ASIG5V.n3357 VSS 0.056945f
C2412 ASIG5V.n3358 VSS 0.056945f
C2413 ASIG5V.n3359 VSS 0.056945f
C2414 ASIG5V.n3360 VSS 0.056945f
C2415 ASIG5V.n3363 VSS 0.056945f
C2416 ASIG5V.n3364 VSS 0.056945f
C2417 ASIG5V.n3365 VSS 0.056945f
C2418 ASIG5V.n3366 VSS 0.056945f
C2419 ASIG5V.n3369 VSS 0.056945f
C2420 ASIG5V.n3370 VSS 0.056945f
C2421 ASIG5V.n3371 VSS 0.056945f
C2422 ASIG5V.n3372 VSS 0.056945f
C2423 ASIG5V.n3375 VSS 0.056945f
C2424 ASIG5V.n3376 VSS 0.056945f
C2425 ASIG5V.n3377 VSS 0.056945f
C2426 ASIG5V.n3378 VSS 0.056945f
C2427 ASIG5V.n3381 VSS 0.056945f
C2428 ASIG5V.n3382 VSS 0.056945f
C2429 ASIG5V.n3383 VSS 0.056945f
C2430 ASIG5V.n3384 VSS 0.056945f
C2431 ASIG5V.n3387 VSS 0.056945f
C2432 ASIG5V.n3388 VSS 0.056945f
C2433 ASIG5V.n3389 VSS 0.056945f
C2434 ASIG5V.n3390 VSS 0.056945f
C2435 ASIG5V.n3393 VSS 0.056945f
C2436 ASIG5V.n3394 VSS 0.056945f
C2437 ASIG5V.n3395 VSS 0.056945f
C2438 ASIG5V.n3396 VSS 0.056945f
C2439 ASIG5V.n3399 VSS 0.056945f
C2440 ASIG5V.n3400 VSS 0.056945f
C2441 ASIG5V.n3401 VSS 0.056945f
C2442 ASIG5V.n3402 VSS 0.056945f
C2443 ASIG5V.n3405 VSS 0.036092f
C2444 ASIG5V.n3406 VSS 0.036092f
C2445 ASIG5V.n3407 VSS 0.047722f
C2446 ASIG5V.n3408 VSS 0.056945f
C2447 ASIG5V.n3409 VSS 0.056945f
C2448 ASIG5V.n3410 VSS 0.056945f
C2449 ASIG5V.n3412 VSS 0.056945f
C2450 ASIG5V.n3414 VSS 0.056945f
C2451 ASIG5V.n3415 VSS 0.056945f
C2452 ASIG5V.n3416 VSS 0.056945f
C2453 ASIG5V.n3417 VSS 0.056945f
C2454 ASIG5V.n3418 VSS 0.056945f
C2455 ASIG5V.n3419 VSS 0.056945f
C2456 ASIG5V.n3420 VSS 0.056945f
C2457 ASIG5V.n3422 VSS 0.056945f
C2458 ASIG5V.n3424 VSS 0.056945f
C2459 ASIG5V.n3425 VSS 0.056945f
C2460 ASIG5V.n3426 VSS 0.056945f
C2461 ASIG5V.n3427 VSS 0.056945f
C2462 ASIG5V.n3428 VSS 0.056945f
C2463 ASIG5V.n3429 VSS 0.056945f
C2464 ASIG5V.n3430 VSS 0.056945f
C2465 ASIG5V.n3432 VSS 0.056945f
C2466 ASIG5V.n3434 VSS 0.056945f
C2467 ASIG5V.n3435 VSS 0.056945f
C2468 ASIG5V.n3436 VSS 0.056945f
C2469 ASIG5V.n3437 VSS 0.056945f
C2470 ASIG5V.n3438 VSS 0.056945f
C2471 ASIG5V.n3439 VSS 0.056945f
C2472 ASIG5V.n3440 VSS 0.056945f
C2473 ASIG5V.n3442 VSS 0.056945f
C2474 ASIG5V.n3444 VSS 0.056945f
C2475 ASIG5V.n3445 VSS 0.056945f
C2476 ASIG5V.n3446 VSS 0.056945f
C2477 ASIG5V.n3447 VSS 0.056945f
C2478 ASIG5V.n3448 VSS 0.056945f
C2479 ASIG5V.n3449 VSS 0.056945f
C2480 ASIG5V.n3450 VSS 0.056945f
C2481 ASIG5V.n3452 VSS 0.056945f
C2482 ASIG5V.n3454 VSS 0.056945f
C2483 ASIG5V.n3455 VSS 0.056945f
C2484 ASIG5V.n3456 VSS 0.056945f
C2485 ASIG5V.n3457 VSS 0.056945f
C2486 ASIG5V.n3458 VSS 0.056945f
C2487 ASIG5V.n3459 VSS 0.056945f
C2488 ASIG5V.n3460 VSS 0.056945f
C2489 ASIG5V.n3462 VSS 0.056945f
C2490 ASIG5V.n3464 VSS 0.056945f
C2491 ASIG5V.n3465 VSS 0.056945f
C2492 ASIG5V.n3466 VSS 0.056945f
C2493 ASIG5V.n3467 VSS 0.056945f
C2494 ASIG5V.n3468 VSS 0.056945f
C2495 ASIG5V.n3469 VSS 0.056945f
C2496 ASIG5V.n3470 VSS 0.056945f
C2497 ASIG5V.n3472 VSS 0.056945f
C2498 ASIG5V.n3474 VSS 0.056945f
C2499 ASIG5V.n3475 VSS 0.056945f
C2500 ASIG5V.n3476 VSS 0.056945f
C2501 ASIG5V.n3477 VSS 0.056945f
C2502 ASIG5V.n3478 VSS 0.056945f
C2503 ASIG5V.n3479 VSS 0.056945f
C2504 ASIG5V.n3480 VSS 0.056945f
C2505 ASIG5V.n3482 VSS 0.056945f
C2506 ASIG5V.n3484 VSS 0.056945f
C2507 ASIG5V.n3485 VSS 0.056945f
C2508 ASIG5V.n3486 VSS 0.056945f
C2509 ASIG5V.n3487 VSS 0.056945f
C2510 ASIG5V.n3488 VSS 0.056945f
C2511 ASIG5V.n3489 VSS 0.056945f
C2512 ASIG5V.n3490 VSS 0.056945f
C2513 ASIG5V.n3492 VSS 0.056945f
C2514 ASIG5V.n3494 VSS 0.056945f
C2515 ASIG5V.n3495 VSS 0.056945f
C2516 ASIG5V.n3496 VSS 0.056945f
C2517 ASIG5V.n3497 VSS 0.056945f
C2518 ASIG5V.n3498 VSS 0.056945f
C2519 ASIG5V.n3499 VSS 0.056945f
C2520 ASIG5V.n3500 VSS 0.056945f
C2521 ASIG5V.n3502 VSS 0.056945f
C2522 ASIG5V.n3504 VSS 0.056945f
C2523 ASIG5V.n3505 VSS 0.056945f
C2524 ASIG5V.n3506 VSS 0.056945f
C2525 ASIG5V.n3507 VSS 0.056945f
C2526 ASIG5V.n3508 VSS 0.056945f
C2527 ASIG5V.n3509 VSS 0.056945f
C2528 ASIG5V.n3510 VSS 0.056945f
C2529 ASIG5V.n3512 VSS 0.056945f
C2530 ASIG5V.n3514 VSS 0.056945f
C2531 ASIG5V.n3515 VSS 0.056945f
C2532 ASIG5V.n3516 VSS 0.056945f
C2533 ASIG5V.n3517 VSS 0.056945f
C2534 ASIG5V.n3518 VSS 0.056945f
C2535 ASIG5V.n3519 VSS 0.056945f
C2536 ASIG5V.n3520 VSS 0.056945f
C2537 ASIG5V.n3522 VSS 0.056945f
C2538 ASIG5V.n3524 VSS 0.056945f
C2539 ASIG5V.n3525 VSS 0.056945f
C2540 ASIG5V.n3526 VSS 0.056945f
C2541 ASIG5V.n3527 VSS 0.056945f
C2542 ASIG5V.n3528 VSS 0.056945f
C2543 ASIG5V.n3529 VSS 0.056945f
C2544 ASIG5V.n3530 VSS 0.056945f
C2545 ASIG5V.n3532 VSS 0.056945f
C2546 ASIG5V.n3534 VSS 0.056945f
C2547 ASIG5V.n3535 VSS 0.056945f
C2548 ASIG5V.n3536 VSS 0.056945f
C2549 ASIG5V.n3537 VSS 0.056945f
C2550 ASIG5V.n3538 VSS 0.056945f
C2551 ASIG5V.n3539 VSS 0.056945f
C2552 ASIG5V.n3540 VSS 0.056945f
C2553 ASIG5V.n3542 VSS 0.056945f
C2554 ASIG5V.n3544 VSS 0.056945f
C2555 ASIG5V.n3545 VSS 0.056945f
C2556 ASIG5V.n3546 VSS 0.056945f
C2557 ASIG5V.n3547 VSS 0.056945f
C2558 ASIG5V.n3548 VSS 0.056945f
C2559 ASIG5V.n3549 VSS 0.056945f
C2560 ASIG5V.n3550 VSS 0.056945f
C2561 ASIG5V.n3552 VSS 0.056945f
C2562 ASIG5V.n3554 VSS 0.056945f
C2563 ASIG5V.n3555 VSS 0.056945f
C2564 ASIG5V.n3556 VSS 0.056945f
C2565 ASIG5V.n3557 VSS 0.056945f
C2566 ASIG5V.n3558 VSS 0.056945f
C2567 ASIG5V.n3559 VSS 0.056945f
C2568 ASIG5V.n3560 VSS 0.056945f
C2569 ASIG5V.n3562 VSS 0.056945f
C2570 ASIG5V.n3564 VSS 0.056945f
C2571 ASIG5V.n3565 VSS 0.056945f
C2572 ASIG5V.n3566 VSS 0.056945f
C2573 ASIG5V.n3567 VSS 0.056945f
C2574 ASIG5V.n3568 VSS 0.056945f
C2575 ASIG5V.n3569 VSS 0.056945f
C2576 ASIG5V.n3570 VSS 0.056945f
C2577 ASIG5V.n3572 VSS 0.056945f
C2578 ASIG5V.n3574 VSS 0.056945f
C2579 ASIG5V.n3575 VSS 0.056945f
C2580 ASIG5V.n3576 VSS 0.056945f
C2581 ASIG5V.n3577 VSS 0.056945f
C2582 ASIG5V.n3578 VSS 0.056945f
C2583 ASIG5V.n3579 VSS 0.056945f
C2584 ASIG5V.n3580 VSS 0.056945f
C2585 ASIG5V.n3582 VSS 0.056945f
C2586 ASIG5V.n3584 VSS 0.056945f
C2587 ASIG5V.n3585 VSS 0.056945f
C2588 ASIG5V.n3586 VSS 0.056945f
C2589 ASIG5V.n3587 VSS 0.056945f
C2590 ASIG5V.n3588 VSS 0.056945f
C2591 ASIG5V.n3589 VSS 0.056945f
C2592 ASIG5V.n3590 VSS 0.056945f
C2593 ASIG5V.n3592 VSS 0.056945f
C2594 ASIG5V.n3594 VSS 0.056945f
C2595 ASIG5V.n3595 VSS 0.056945f
C2596 ASIG5V.n3596 VSS 0.056945f
C2597 ASIG5V.n3597 VSS 0.056945f
C2598 ASIG5V.n3598 VSS 0.056945f
C2599 ASIG5V.n3599 VSS 0.056945f
C2600 ASIG5V.n3600 VSS 0.056945f
C2601 ASIG5V.n3602 VSS 0.056945f
C2602 ASIG5V.n3604 VSS 0.056945f
C2603 ASIG5V.n3605 VSS 0.056945f
C2604 ASIG5V.n3606 VSS 0.056945f
C2605 ASIG5V.n3607 VSS 0.056945f
C2606 ASIG5V.n3608 VSS 0.056945f
C2607 ASIG5V.n3609 VSS 0.056945f
C2608 ASIG5V.n3610 VSS 0.056945f
C2609 ASIG5V.n3612 VSS 0.056945f
C2610 ASIG5V.n3614 VSS 0.036092f
C2611 ASIG5V.n3615 VSS 0.036092f
C2612 ASIG5V.n3616 VSS 0.052133f
C2613 ASIG5V.n3617 VSS 0.09726f
C2614 ASIG5V.n3618 VSS 0.108961f
C2615 ASIG5V.n3619 VSS 0.091386f
C2616 ASIG5V.n3620 VSS 0.955415f
C2617 ASIG5V.n3621 VSS 0.070496f
C2618 ASIG5V.n3622 VSS 0.070496f
C2619 ASIG5V.n3623 VSS 0.047722f
C2620 ASIG5V.n3624 VSS 0.066995f
C2621 ASIG5V.n3625 VSS 0.076709f
C2622 ASIG5V.n3626 VSS 0.045974f
C2623 ASIG5V.n3627 VSS 0.076709f
C2624 ASIG5V.n3628 VSS 0.045974f
C2625 ASIG5V.n3629 VSS 0.346723f
C2626 ASIG5V.n3671 VSS 0.056945f
C2627 ASIG5V.n3672 VSS 0.0621f
C2628 ASIG5V.n3673 VSS 0.036092f
C2629 ASIG5V.n3674 VSS 0.747381f
C2630 ASIG5V.n3716 VSS 0.056945f
C2631 ASIG5V.n3717 VSS 0.056945f
C2632 ASIG5V.n3718 VSS 0.056945f
C2633 ASIG5V.n3719 VSS 0.056945f
C2634 ASIG5V.n3720 VSS 0.056945f
C2635 ASIG5V.n3721 VSS 0.056945f
C2636 ASIG5V.n3722 VSS 0.056945f
C2637 ASIG5V.n3723 VSS 0.056945f
C2638 ASIG5V.n3724 VSS 0.056945f
C2639 ASIG5V.n3725 VSS 0.056945f
C2640 ASIG5V.n3726 VSS 0.056945f
C2641 ASIG5V.n3727 VSS 0.056945f
C2642 ASIG5V.n3728 VSS 0.056945f
C2643 ASIG5V.n3729 VSS 0.056945f
C2644 ASIG5V.n3730 VSS 0.056945f
C2645 ASIG5V.n3731 VSS 0.056945f
C2646 ASIG5V.n3732 VSS 0.056945f
C2647 ASIG5V.n3733 VSS 0.056945f
C2648 ASIG5V.n3734 VSS 0.056945f
C2649 ASIG5V.n3735 VSS 0.056945f
C2650 ASIG5V.n3736 VSS 0.056945f
C2651 ASIG5V.n3737 VSS 0.056945f
C2652 ASIG5V.n3738 VSS 0.056945f
C2653 ASIG5V.n3739 VSS 0.056945f
C2654 ASIG5V.n3740 VSS 0.056945f
C2655 ASIG5V.n3741 VSS 0.056945f
C2656 ASIG5V.n3742 VSS 0.056945f
C2657 ASIG5V.n3743 VSS 0.056945f
C2658 ASIG5V.n3744 VSS 0.056945f
C2659 ASIG5V.n3745 VSS 0.056945f
C2660 ASIG5V.n3746 VSS 0.056945f
C2661 ASIG5V.n3747 VSS 0.056945f
C2662 ASIG5V.n3748 VSS 0.056945f
C2663 ASIG5V.n3749 VSS 0.056945f
C2664 ASIG5V.n3750 VSS 0.056945f
C2665 ASIG5V.n3751 VSS 0.056945f
C2666 ASIG5V.n3752 VSS 0.056945f
C2667 ASIG5V.n3753 VSS 0.056945f
C2668 ASIG5V.n3754 VSS 0.056945f
C2669 ASIG5V.n3755 VSS 0.056945f
C2670 ASIG5V.n3756 VSS 0.056945f
C2671 ASIG5V.n3757 VSS 0.056945f
C2672 ASIG5V.n3758 VSS 0.056945f
C2673 ASIG5V.n3759 VSS 0.056945f
C2674 ASIG5V.n3760 VSS 0.056945f
C2675 ASIG5V.n3761 VSS 0.056945f
C2676 ASIG5V.n3762 VSS 0.056945f
C2677 ASIG5V.n3763 VSS 0.056945f
C2678 ASIG5V.n3764 VSS 0.056945f
C2679 ASIG5V.n3765 VSS 0.056945f
C2680 ASIG5V.n3766 VSS 0.056945f
C2681 ASIG5V.n3767 VSS 0.056945f
C2682 ASIG5V.n3768 VSS 0.056945f
C2683 ASIG5V.n3769 VSS 0.056945f
C2684 ASIG5V.n3770 VSS 0.056945f
C2685 ASIG5V.n3771 VSS 0.056945f
C2686 ASIG5V.n3772 VSS 0.056945f
C2687 ASIG5V.n3773 VSS 0.056945f
C2688 ASIG5V.n3774 VSS 0.056945f
C2689 ASIG5V.n3775 VSS 0.056945f
C2690 ASIG5V.n3776 VSS 0.056945f
C2691 ASIG5V.n3777 VSS 0.064317f
C2692 ASIG5V.n3778 VSS 0.108961f
C2693 ASIG5V.n3779 VSS 0.0621f
C2694 ASIG5V.n3780 VSS 0.955415f
C2695 ASIG5V.n3781 VSS 1.0941f
C2696 ASIG5V.n3782 VSS 0.0621f
C2697 ASIG5V.n3783 VSS 0.052133f
C2698 ASIG5V.n3784 VSS 0.09726f
C2699 ASIG5V.n3785 VSS 0.108961f
C2700 ASIG5V.n3786 VSS 0.108961f
C2701 ASIG5V.n3787 VSS 0.470002f
C2702 ASIG5V.n3829 VSS 0.036092f
C2703 ASIG5V.n3830 VSS 0.331313f
C2704 ASIG5V.n3831 VSS 0.045974f
C2705 ASIG5V.n3833 VSS 0.056945f
C2706 ASIG5V.n3834 VSS 0.056945f
C2707 ASIG5V.n3835 VSS 0.045974f
C2708 ASIG5V.n3836 VSS 0.056945f
C2709 ASIG5V.n3837 VSS 0.066995f
C2710 ASIG5V.n3838 VSS 0.076709f
C2711 ASIG5V.n3839 VSS 0.046187f
C2712 ASIG5V.n3840 VSS 0.955415f
C2713 ASIG5V.n3841 VSS 0.103317f
C2714 ASIG5V.n3842 VSS 0.103317f
C2715 ASIG5V.n3843 VSS 0.201323f
C2716 ASIG5V.n3844 VSS 0.161825f
C2717 ASIG5V.n3845 VSS 0.161825f
C2718 ASIG5V.n3847 VSS 0.955416f
C2719 ASIG5V.n3848 VSS 0.955416f
C2720 ASIG5V.n3849 VSS 0.955416f
C2721 ASIG5V.n3850 VSS 0.955416f
C2722 ASIG5V.n3851 VSS 1.01706f
C2723 ASIG5V.n3852 VSS 0.108041f
C2724 ASIG5V.n3853 VSS 0.108041f
C2725 ASIG5V.n3855 VSS 0.955416f
C2726 ASIG5V.n3856 VSS 0.161825f
C2727 ASIG5V.n3857 VSS 0.955416f
C2728 ASIG5V.n3858 VSS 0.955416f
C2729 ASIG5V.n3859 VSS 0.117005f
C2730 ASIG5V.n3860 VSS 0.117005f
C2731 ASIG5V.n3861 VSS 0.117005f
C2732 ASIG5V.n3862 VSS 0.117005f
C2733 ASIG5V.n3863 VSS 0.117005f
C2734 ASIG5V.n3864 VSS 0.117005f
C2735 ASIG5V.n3865 VSS 0.117005f
C2736 ASIG5V.n3866 VSS 0.117005f
C2737 ASIG5V.n3867 VSS 0.117005f
C2738 ASIG5V.n3868 VSS 0.117005f
C2739 ASIG5V.n3869 VSS 0.117005f
C2740 ASIG5V.n3870 VSS 0.117005f
C2741 ASIG5V.n3871 VSS 0.117005f
C2742 ASIG5V.n3872 VSS 0.117005f
C2743 ASIG5V.n3873 VSS 0.117005f
C2744 ASIG5V.n3874 VSS 0.117005f
C2745 ASIG5V.n3875 VSS 0.117005f
C2746 ASIG5V.n3876 VSS 0.117005f
C2747 ASIG5V.n3877 VSS 0.117005f
C2748 ASIG5V.n3878 VSS 0.117005f
C2749 ASIG5V.n3879 VSS 0.117005f
C2750 ASIG5V.n3880 VSS 0.117005f
C2751 ASIG5V.n3881 VSS 0.117005f
C2752 ASIG5V.n3882 VSS 0.117005f
C2753 ASIG5V.n3883 VSS 0.117005f
C2754 ASIG5V.n3884 VSS 0.117005f
C2755 ASIG5V.n3885 VSS 0.117005f
C2756 ASIG5V.n3886 VSS 0.117005f
C2757 ASIG5V.n3887 VSS 0.117005f
C2758 ASIG5V.n3888 VSS 0.117005f
C2759 ASIG5V.n3889 VSS 0.117005f
C2760 ASIG5V.n3890 VSS 0.117005f
C2761 ASIG5V.n3891 VSS 0.117005f
C2762 ASIG5V.n3892 VSS 0.117005f
C2763 ASIG5V.n3893 VSS 0.117005f
C2764 ASIG5V.n3894 VSS 0.117005f
C2765 ASIG5V.n3895 VSS 0.117005f
C2766 ASIG5V.n3896 VSS 0.117005f
C2767 ASIG5V.n3897 VSS 0.117005f
C2768 ASIG5V.n3898 VSS 0.117005f
C2769 ASIG5V.n3899 VSS 0.117005f
C2770 ASIG5V.n3900 VSS 0.117005f
C2771 ASIG5V.n3901 VSS 0.117005f
C2772 ASIG5V.n3902 VSS 0.117005f
C2773 ASIG5V.n3903 VSS 0.117005f
C2774 ASIG5V.n3904 VSS 0.117005f
C2775 ASIG5V.n3905 VSS 0.117005f
C2776 ASIG5V.n3906 VSS 0.117005f
C2777 ASIG5V.n3908 VSS 0.117005f
C2778 ASIG5V.n3909 VSS 0.19202f
C2779 ASIG5V.n3911 VSS 0.117005f
C2780 ASIG5V.n3913 VSS 0.117005f
C2781 ASIG5V.n3915 VSS 0.117005f
C2782 ASIG5V.n3917 VSS 0.117005f
C2783 ASIG5V.n3919 VSS 0.117005f
C2784 ASIG5V.n3921 VSS 0.117005f
C2785 ASIG5V.n3923 VSS 0.117005f
C2786 ASIG5V.n3925 VSS 0.117005f
C2787 ASIG5V.n3927 VSS 0.117005f
C2788 ASIG5V.n3929 VSS 0.117005f
C2789 ASIG5V.n3931 VSS 0.117005f
C2790 ASIG5V.n3933 VSS 0.117005f
C2791 ASIG5V.n3935 VSS 0.117005f
C2792 ASIG5V.n3937 VSS 0.117005f
C2793 ASIG5V.n3939 VSS 0.117005f
C2794 ASIG5V.n3941 VSS 0.117005f
C2795 ASIG5V.n3943 VSS 0.117005f
C2796 ASIG5V.n3945 VSS 0.117005f
C2797 ASIG5V.n3947 VSS 0.117005f
C2798 ASIG5V.n3949 VSS 0.117005f
C2799 ASIG5V.n3951 VSS 0.117005f
C2800 ASIG5V.n3953 VSS 0.117005f
C2801 ASIG5V.n3955 VSS 0.117005f
C2802 ASIG5V.n3957 VSS 0.117005f
C2803 ASIG5V.n3959 VSS 0.117005f
C2804 ASIG5V.n3961 VSS 0.117005f
C2805 ASIG5V.n3963 VSS 0.117005f
C2806 ASIG5V.n3965 VSS 0.117005f
C2807 ASIG5V.n3967 VSS 0.117005f
C2808 ASIG5V.n3969 VSS 0.117005f
C2809 ASIG5V.n3971 VSS 0.117005f
C2810 ASIG5V.n3973 VSS 0.117005f
C2811 ASIG5V.n3975 VSS 0.117005f
C2812 ASIG5V.n3977 VSS 0.117005f
C2813 ASIG5V.n3979 VSS 0.117005f
C2814 ASIG5V.n3981 VSS 0.117005f
C2815 ASIG5V.n3983 VSS 0.117005f
C2816 ASIG5V.n3985 VSS 0.117005f
C2817 ASIG5V.n3987 VSS 0.117005f
C2818 ASIG5V.n3989 VSS 0.117005f
C2819 ASIG5V.n3991 VSS 0.117005f
C2820 ASIG5V.n3993 VSS 0.117005f
C2821 ASIG5V.n3995 VSS 0.117005f
C2822 ASIG5V.n3997 VSS 0.117005f
C2823 ASIG5V.n3999 VSS 0.117005f
C2824 ASIG5V.n4001 VSS 0.117005f
C2825 ASIG5V.n4003 VSS 0.117005f
C2826 ASIG5V.n4051 VSS 0.955416f
C2827 ASIG5V.n4053 VSS 0.117005f
C2828 ASIG5V.n4054 VSS 0.117005f
C2829 ASIG5V.n4055 VSS 0.117005f
C2830 ASIG5V.n4056 VSS 0.117005f
C2831 ASIG5V.n4057 VSS 0.117005f
C2832 ASIG5V.n4058 VSS 0.117005f
C2833 ASIG5V.n4059 VSS 0.117005f
C2834 ASIG5V.n4060 VSS 0.117005f
C2835 ASIG5V.n4061 VSS 0.117005f
C2836 ASIG5V.n4062 VSS 0.117005f
C2837 ASIG5V.n4063 VSS 0.117005f
C2838 ASIG5V.n4064 VSS 0.117005f
C2839 ASIG5V.n4065 VSS 0.117005f
C2840 ASIG5V.n4066 VSS 0.117005f
C2841 ASIG5V.n4067 VSS 0.117005f
C2842 ASIG5V.n4068 VSS 0.117005f
C2843 ASIG5V.n4069 VSS 0.117005f
C2844 ASIG5V.n4070 VSS 0.117005f
C2845 ASIG5V.n4071 VSS 0.117005f
C2846 ASIG5V.n4072 VSS 0.117005f
C2847 ASIG5V.n4073 VSS 0.117005f
C2848 ASIG5V.n4074 VSS 0.117005f
C2849 ASIG5V.n4075 VSS 0.117005f
C2850 ASIG5V.n4076 VSS 0.117005f
C2851 ASIG5V.n4077 VSS 0.117005f
C2852 ASIG5V.n4078 VSS 0.117005f
C2853 ASIG5V.n4079 VSS 0.117005f
C2854 ASIG5V.n4080 VSS 0.117005f
C2855 ASIG5V.n4081 VSS 0.117005f
C2856 ASIG5V.n4082 VSS 0.117005f
C2857 ASIG5V.n4083 VSS 0.117005f
C2858 ASIG5V.n4084 VSS 0.117005f
C2859 ASIG5V.n4085 VSS 0.117005f
C2860 ASIG5V.n4086 VSS 0.117005f
C2861 ASIG5V.n4087 VSS 0.117005f
C2862 ASIG5V.n4088 VSS 0.117005f
C2863 ASIG5V.n4089 VSS 0.117005f
C2864 ASIG5V.n4090 VSS 0.117005f
C2865 ASIG5V.n4091 VSS 0.117005f
C2866 ASIG5V.n4092 VSS 0.117005f
C2867 ASIG5V.n4093 VSS 0.117005f
C2868 ASIG5V.n4094 VSS 0.117005f
C2869 ASIG5V.n4095 VSS 0.117005f
C2870 ASIG5V.n4096 VSS 0.117005f
C2871 ASIG5V.n4097 VSS 0.117005f
C2872 ASIG5V.n4098 VSS 0.117005f
C2873 ASIG5V.n4099 VSS 0.117005f
C2874 ASIG5V.n4100 VSS 0.117005f
C2875 ASIG5V.n4101 VSS 0.161825f
C2876 ASIG5V.n4102 VSS 0.117005f
C2877 ASIG5V.n4103 VSS 0.117005f
C2878 ASIG5V.n4104 VSS 0.117005f
C2879 ASIG5V.n4105 VSS 0.117005f
C2880 ASIG5V.n4106 VSS 0.117005f
C2881 ASIG5V.n4107 VSS 0.117005f
C2882 ASIG5V.n4108 VSS 0.117005f
C2883 ASIG5V.n4109 VSS 0.117005f
C2884 ASIG5V.n4110 VSS 0.117005f
C2885 ASIG5V.n4111 VSS 0.117005f
C2886 ASIG5V.n4112 VSS 0.117005f
C2887 ASIG5V.n4113 VSS 0.117005f
C2888 ASIG5V.n4114 VSS 0.117005f
C2889 ASIG5V.n4115 VSS 0.117005f
C2890 ASIG5V.n4116 VSS 0.117005f
C2891 ASIG5V.n4117 VSS 0.117005f
C2892 ASIG5V.n4118 VSS 0.117005f
C2893 ASIG5V.n4119 VSS 0.117005f
C2894 ASIG5V.n4120 VSS 0.117005f
C2895 ASIG5V.n4121 VSS 0.117005f
C2896 ASIG5V.n4122 VSS 0.117005f
C2897 ASIG5V.n4123 VSS 0.117005f
C2898 ASIG5V.n4124 VSS 0.117005f
C2899 ASIG5V.n4125 VSS 0.117005f
C2900 ASIG5V.n4126 VSS 0.117005f
C2901 ASIG5V.n4127 VSS 0.117005f
C2902 ASIG5V.n4128 VSS 0.117005f
C2903 ASIG5V.n4129 VSS 0.117005f
C2904 ASIG5V.n4130 VSS 0.117005f
C2905 ASIG5V.n4131 VSS 0.117005f
C2906 ASIG5V.n4132 VSS 0.117005f
C2907 ASIG5V.n4133 VSS 0.117005f
C2908 ASIG5V.n4134 VSS 0.117005f
C2909 ASIG5V.n4135 VSS 0.117005f
C2910 ASIG5V.n4136 VSS 0.117005f
C2911 ASIG5V.n4137 VSS 0.117005f
C2912 ASIG5V.n4138 VSS 0.117005f
C2913 ASIG5V.n4139 VSS 0.117005f
C2914 ASIG5V.n4140 VSS 0.117005f
C2915 ASIG5V.n4141 VSS 0.117005f
C2916 ASIG5V.n4142 VSS 0.117005f
C2917 ASIG5V.n4143 VSS 0.117005f
C2918 ASIG5V.n4144 VSS 0.117005f
C2919 ASIG5V.n4145 VSS 0.117005f
C2920 ASIG5V.n4146 VSS 0.117005f
C2921 ASIG5V.n4147 VSS 0.117005f
C2922 ASIG5V.n4148 VSS 0.117005f
C2923 ASIG5V.n4149 VSS 0.117005f
C2924 ASIG5V.n4150 VSS 0.117005f
C2925 ASIG5V.n4151 VSS 0.117005f
C2926 ASIG5V.n4152 VSS 0.117005f
C2927 ASIG5V.n4153 VSS 0.117005f
C2928 ASIG5V.n4154 VSS 0.117005f
C2929 ASIG5V.n4155 VSS 0.117005f
C2930 ASIG5V.n4156 VSS 0.117005f
C2931 ASIG5V.n4157 VSS 0.117005f
C2932 ASIG5V.n4158 VSS 0.117005f
C2933 ASIG5V.n4159 VSS 0.117005f
C2934 ASIG5V.n4160 VSS 0.117005f
C2935 ASIG5V.n4161 VSS 0.117005f
C2936 ASIG5V.n4162 VSS 0.117005f
C2937 ASIG5V.n4163 VSS 0.117005f
C2938 ASIG5V.n4164 VSS 0.117005f
C2939 ASIG5V.n4165 VSS 0.117005f
C2940 ASIG5V.n4166 VSS 0.117005f
C2941 ASIG5V.n4167 VSS 0.117005f
C2942 ASIG5V.n4168 VSS 0.117005f
C2943 ASIG5V.n4169 VSS 0.117005f
C2944 ASIG5V.n4170 VSS 0.117005f
C2945 ASIG5V.n4171 VSS 0.117005f
C2946 ASIG5V.n4172 VSS 0.117005f
C2947 ASIG5V.n4173 VSS 0.117005f
C2948 ASIG5V.n4174 VSS 0.117005f
C2949 ASIG5V.n4175 VSS 0.117005f
C2950 ASIG5V.n4176 VSS 0.117005f
C2951 ASIG5V.n4177 VSS 0.117005f
C2952 ASIG5V.n4178 VSS 0.117005f
C2953 ASIG5V.n4179 VSS 0.117005f
C2954 ASIG5V.n4180 VSS 0.117005f
C2955 ASIG5V.n4181 VSS 0.117005f
C2956 ASIG5V.n4182 VSS 0.117005f
C2957 ASIG5V.n4183 VSS 0.117005f
C2958 ASIG5V.n4184 VSS 0.117005f
C2959 ASIG5V.n4185 VSS 0.117005f
C2960 ASIG5V.n4186 VSS 0.117005f
C2961 ASIG5V.n4187 VSS 0.117005f
C2962 ASIG5V.n4188 VSS 0.117005f
C2963 ASIG5V.n4189 VSS 0.117005f
C2964 ASIG5V.n4190 VSS 0.117005f
C2965 ASIG5V.n4191 VSS 0.117005f
C2966 ASIG5V.n4192 VSS 0.117005f
C2967 ASIG5V.n4193 VSS 0.117005f
C2968 ASIG5V.n4194 VSS 0.117005f
C2969 ASIG5V.n4195 VSS 0.117005f
C2970 ASIG5V.n4196 VSS 0.117005f
C2971 ASIG5V.n4197 VSS 0.117005f
C2972 ASIG5V.n4198 VSS 0.117005f
C2973 ASIG5V.n4199 VSS 0.117005f
C2974 ASIG5V.n4200 VSS 0.117005f
C2975 ASIG5V.n4201 VSS 0.117005f
C2976 ASIG5V.n4202 VSS 0.117005f
C2977 ASIG5V.n4203 VSS 0.117005f
C2978 ASIG5V.n4204 VSS 0.117005f
C2979 ASIG5V.n4205 VSS 0.117005f
C2980 ASIG5V.n4206 VSS 0.117005f
C2981 ASIG5V.n4207 VSS 0.117005f
C2982 ASIG5V.n4208 VSS 0.117005f
C2983 ASIG5V.n4209 VSS 0.117005f
C2984 ASIG5V.n4210 VSS 0.117005f
C2985 ASIG5V.n4211 VSS 0.117005f
C2986 ASIG5V.n4212 VSS 0.117005f
C2987 ASIG5V.n4213 VSS 0.117005f
C2988 ASIG5V.n4214 VSS 0.117005f
C2989 ASIG5V.n4215 VSS 0.117005f
C2990 ASIG5V.n4216 VSS 0.117005f
C2991 ASIG5V.n4217 VSS 0.117005f
C2992 ASIG5V.n4218 VSS 0.117005f
C2993 ASIG5V.n4219 VSS 0.117005f
C2994 ASIG5V.n4220 VSS 0.117005f
C2995 ASIG5V.n4221 VSS 0.117005f
C2996 ASIG5V.n4222 VSS 0.117005f
C2997 ASIG5V.n4223 VSS 0.117005f
C2998 ASIG5V.n4224 VSS 0.117005f
C2999 ASIG5V.n4225 VSS 0.117005f
C3000 ASIG5V.n4226 VSS 0.117005f
C3001 ASIG5V.n4227 VSS 0.117005f
C3002 ASIG5V.n4228 VSS 0.117005f
C3003 ASIG5V.n4229 VSS 0.117005f
C3004 ASIG5V.n4230 VSS 0.117005f
C3005 ASIG5V.n4231 VSS 0.117005f
C3006 ASIG5V.n4232 VSS 0.117005f
C3007 ASIG5V.n4233 VSS 0.117005f
C3008 ASIG5V.n4234 VSS 0.117005f
C3009 ASIG5V.n4235 VSS 0.117005f
C3010 ASIG5V.n4236 VSS 0.117005f
C3011 ASIG5V.n4237 VSS 0.117005f
C3012 ASIG5V.n4238 VSS 0.117005f
C3013 ASIG5V.n4239 VSS 0.117005f
C3014 ASIG5V.n4240 VSS 0.117005f
C3015 ASIG5V.n4241 VSS 0.117005f
C3016 ASIG5V.n4242 VSS 0.117005f
C3017 ASIG5V.n4243 VSS 0.117005f
C3018 ASIG5V.n4244 VSS 0.117005f
C3019 ASIG5V.n4245 VSS 0.117005f
C3020 ASIG5V.n4246 VSS 0.106625f
C3021 ASIG5V.n4247 VSS 0.192509f
C3022 ASIG5V.n4248 VSS 0.243192f
C3023 ASIG5V.n4249 VSS 0.040338f
C3024 ASIG5V.n4250 VSS 0.046187f
C3025 ASIG5V.n4251 VSS 0.066335f
C3026 ASIG5V.n4252 VSS 0.092943f
C3027 ASIG5V.n4253 VSS 0.066335f
C3028 ASIG5V.n4254 VSS 0.092943f
C3029 ASIG5V.n4255 VSS 2.37313f
C3030 ASIG5V.n4256 VSS 0.161825f
C3031 ASIG5V.n4257 VSS 0.161825f
C3032 ASIG5V.n4259 VSS 0.196332f
C3033 ASIG5V.n4260 VSS 1.34837f
C3034 ASIG5V.n4261 VSS 0.067466f
C3035 ASIG5V.n4262 VSS 0.067466f
C3036 ASIG5V.n4263 VSS 0.086338f
C3037 ASIG5V.n4264 VSS 0.373154f
C3038 ASIG5V.n4265 VSS 0.088632f
C3039 ASIG5V.n4266 VSS 0.099295f
C3040 ASIG5V.n4267 VSS 0.099295f
C3041 ASIG5V.n4268 VSS 1.0941f
C3042 ASIG5V.n4309 VSS 0.036092f
C3043 ASIG5V.n4310 VSS 0.056945f
C3044 ASIG5V.n4311 VSS 0.056945f
C3045 ASIG5V.n4312 VSS 0.056945f
C3046 ASIG5V.n4313 VSS 0.056945f
C3047 ASIG5V.n4314 VSS 0.056945f
C3048 ASIG5V.n4315 VSS 0.056945f
C3049 ASIG5V.n4316 VSS 0.056945f
C3050 ASIG5V.n4317 VSS 0.056945f
C3051 ASIG5V.n4318 VSS 0.056945f
C3052 ASIG5V.n4319 VSS 0.056945f
C3053 ASIG5V.n4320 VSS 0.056945f
C3054 ASIG5V.n4321 VSS 0.056945f
C3055 ASIG5V.n4322 VSS 0.056945f
C3056 ASIG5V.n4323 VSS 0.056945f
C3057 ASIG5V.n4324 VSS 0.056945f
C3058 ASIG5V.n4325 VSS 0.056945f
C3059 ASIG5V.n4326 VSS 0.056945f
C3060 ASIG5V.n4327 VSS 0.056945f
C3061 ASIG5V.n4328 VSS 0.056945f
C3062 ASIG5V.n4329 VSS 0.056945f
C3063 ASIG5V.n4330 VSS 0.056945f
C3064 ASIG5V.n4331 VSS 0.056945f
C3065 ASIG5V.n4332 VSS 0.056945f
C3066 ASIG5V.n4333 VSS 0.056945f
C3067 ASIG5V.n4334 VSS 0.056945f
C3068 ASIG5V.n4335 VSS 0.056945f
C3069 ASIG5V.n4336 VSS 0.056945f
C3070 ASIG5V.n4337 VSS 0.056945f
C3071 ASIG5V.n4338 VSS 0.056945f
C3072 ASIG5V.n4339 VSS 0.056945f
C3073 ASIG5V.n4340 VSS 0.056945f
C3074 ASIG5V.n4341 VSS 0.056945f
C3075 ASIG5V.n4342 VSS 0.056945f
C3076 ASIG5V.n4343 VSS 0.056945f
C3077 ASIG5V.n4344 VSS 0.056945f
C3078 ASIG5V.n4345 VSS 0.056945f
C3079 ASIG5V.n4346 VSS 0.056945f
C3080 ASIG5V.n4347 VSS 0.056945f
C3081 ASIG5V.n4348 VSS 0.056945f
C3082 ASIG5V.n4349 VSS 0.056945f
C3083 ASIG5V.n4350 VSS 0.056945f
C3084 ASIG5V.n4351 VSS 0.056945f
C3085 ASIG5V.n4352 VSS 0.056945f
C3086 ASIG5V.n4353 VSS 0.056945f
C3087 ASIG5V.n4354 VSS 0.056945f
C3088 ASIG5V.n4355 VSS 0.056945f
C3089 ASIG5V.n4356 VSS 0.056945f
C3090 ASIG5V.n4357 VSS 0.056945f
C3091 ASIG5V.n4358 VSS 0.056945f
C3092 ASIG5V.n4359 VSS 0.056945f
C3093 ASIG5V.n4360 VSS 0.056945f
C3094 ASIG5V.n4361 VSS 0.056945f
C3095 ASIG5V.n4362 VSS 0.056945f
C3096 ASIG5V.n4363 VSS 0.056945f
C3097 ASIG5V.n4364 VSS 0.056945f
C3098 ASIG5V.n4365 VSS 0.056945f
C3099 ASIG5V.n4366 VSS 0.056945f
C3100 ASIG5V.n4367 VSS 0.056945f
C3101 ASIG5V.n4368 VSS 0.056945f
C3102 ASIG5V.n4369 VSS 0.056945f
C3103 ASIG5V.n4370 VSS 0.056945f
C3104 ASIG5V.n4371 VSS 0.056945f
C3105 ASIG5V.n4372 VSS 0.056945f
C3106 ASIG5V.n4373 VSS 0.056945f
C3107 ASIG5V.n4374 VSS 0.056945f
C3108 ASIG5V.n4375 VSS 0.056945f
C3109 ASIG5V.n4376 VSS 0.056945f
C3110 ASIG5V.n4377 VSS 0.056945f
C3111 ASIG5V.n4378 VSS 0.056945f
C3112 ASIG5V.n4379 VSS 0.056945f
C3113 ASIG5V.n4380 VSS 0.056945f
C3114 ASIG5V.n4381 VSS 0.056945f
C3115 ASIG5V.n4382 VSS 0.056945f
C3116 ASIG5V.n4383 VSS 0.056945f
C3117 ASIG5V.n4384 VSS 0.056945f
C3118 ASIG5V.n4385 VSS 0.056945f
C3119 ASIG5V.n4386 VSS 0.056945f
C3120 ASIG5V.n4387 VSS 0.056945f
C3121 ASIG5V.n4388 VSS 0.056945f
C3122 ASIG5V.n4389 VSS 0.056945f
C3123 ASIG5V.n4390 VSS 0.056945f
C3124 ASIG5V.n4391 VSS 0.056945f
C3125 ASIG5V.n4392 VSS 0.056945f
C3126 ASIG5V.n4393 VSS 0.056945f
C3127 ASIG5V.n4394 VSS 0.056945f
C3128 ASIG5V.n4395 VSS 0.056945f
C3129 ASIG5V.n4396 VSS 0.056945f
C3130 ASIG5V.n4397 VSS 0.056945f
C3131 ASIG5V.n4398 VSS 0.056945f
C3132 ASIG5V.n4399 VSS 0.056945f
C3133 ASIG5V.n4400 VSS 0.056945f
C3134 ASIG5V.n4401 VSS 0.056945f
C3135 ASIG5V.n4402 VSS 0.056945f
C3136 ASIG5V.n4403 VSS 0.056945f
C3137 ASIG5V.n4404 VSS 0.056945f
C3138 ASIG5V.n4405 VSS 0.056945f
C3139 ASIG5V.n4406 VSS 0.056945f
C3140 ASIG5V.n4407 VSS 0.056945f
C3141 ASIG5V.n4408 VSS 0.056945f
C3142 ASIG5V.n4409 VSS 0.056945f
C3143 ASIG5V.n4410 VSS 0.056945f
C3144 ASIG5V.n4411 VSS 0.056945f
C3145 ASIG5V.n4412 VSS 0.056945f
C3146 ASIG5V.n4413 VSS 0.056945f
C3147 ASIG5V.n4414 VSS 0.056945f
C3148 ASIG5V.n4415 VSS 0.056945f
C3149 ASIG5V.n4416 VSS 0.056945f
C3150 ASIG5V.n4417 VSS 0.056945f
C3151 ASIG5V.n4418 VSS 0.056945f
C3152 ASIG5V.n4419 VSS 0.056945f
C3153 ASIG5V.n4420 VSS 0.056945f
C3154 ASIG5V.n4421 VSS 0.056945f
C3155 ASIG5V.n4422 VSS 0.056945f
C3156 ASIG5V.n4423 VSS 0.056945f
C3157 ASIG5V.n4424 VSS 0.056945f
C3158 ASIG5V.n4425 VSS 0.056945f
C3159 ASIG5V.n4426 VSS 0.056945f
C3160 ASIG5V.n4427 VSS 0.056945f
C3161 ASIG5V.n4428 VSS 0.056945f
C3162 ASIG5V.n4429 VSS 0.056945f
C3163 ASIG5V.n4430 VSS 0.056945f
C3164 ASIG5V.n4431 VSS 0.056945f
C3165 ASIG5V.n4432 VSS 0.056945f
C3166 ASIG5V.n4433 VSS 0.056945f
C3167 ASIG5V.n4434 VSS 0.056945f
C3168 ASIG5V.n4435 VSS 0.056945f
C3169 ASIG5V.n4436 VSS 0.056945f
C3170 ASIG5V.n4437 VSS 0.056945f
C3171 ASIG5V.n4438 VSS 0.056945f
C3172 ASIG5V.n4439 VSS 0.056945f
C3173 ASIG5V.n4440 VSS 0.056945f
C3174 ASIG5V.n4441 VSS 0.056945f
C3175 ASIG5V.n4442 VSS 0.056945f
C3176 ASIG5V.n4443 VSS 0.056945f
C3177 ASIG5V.n4444 VSS 0.056945f
C3178 ASIG5V.n4445 VSS 0.056945f
C3179 ASIG5V.n4446 VSS 0.056945f
C3180 ASIG5V.n4447 VSS 0.056945f
C3181 ASIG5V.n4448 VSS 0.056945f
C3182 ASIG5V.n4449 VSS 0.056945f
C3183 ASIG5V.n4450 VSS 0.056945f
C3184 ASIG5V.n4451 VSS 0.056945f
C3185 ASIG5V.n4452 VSS 0.056945f
C3186 ASIG5V.n4453 VSS 0.056945f
C3187 ASIG5V.n4454 VSS 0.056945f
C3188 ASIG5V.n4455 VSS 0.056945f
C3189 ASIG5V.n4456 VSS 0.056945f
C3190 ASIG5V.n4457 VSS 0.056945f
C3191 ASIG5V.n4458 VSS 0.056945f
C3192 ASIG5V.n4459 VSS 0.056945f
C3193 ASIG5V.n4460 VSS 0.056945f
C3194 ASIG5V.n4461 VSS 0.056945f
C3195 ASIG5V.n4462 VSS 0.056945f
C3196 ASIG5V.n4463 VSS 0.056945f
C3197 ASIG5V.n4464 VSS 0.056945f
C3198 ASIG5V.n4465 VSS 0.056945f
C3199 ASIG5V.n4466 VSS 0.056945f
C3200 ASIG5V.n4467 VSS 0.056945f
C3201 ASIG5V.n4468 VSS 0.056945f
C3202 ASIG5V.n4469 VSS 0.056945f
C3203 ASIG5V.n4470 VSS 0.056945f
C3204 ASIG5V.n4471 VSS 0.056945f
C3205 ASIG5V.n4472 VSS 0.056945f
C3206 ASIG5V.n4473 VSS 0.056945f
C3207 ASIG5V.n4474 VSS 0.056945f
C3208 ASIG5V.n4475 VSS 0.056945f
C3209 ASIG5V.n4476 VSS 0.056945f
C3210 ASIG5V.n4477 VSS 0.056945f
C3211 ASIG5V.n4478 VSS 0.056945f
C3212 ASIG5V.n4479 VSS 0.056945f
C3213 ASIG5V.n4480 VSS 0.056945f
C3214 ASIG5V.n4481 VSS 0.056945f
C3215 ASIG5V.n4482 VSS 0.056945f
C3216 ASIG5V.n4483 VSS 0.056945f
C3217 ASIG5V.n4484 VSS 0.056945f
C3218 ASIG5V.n4485 VSS 0.056945f
C3219 ASIG5V.n4486 VSS 0.056945f
C3220 ASIG5V.n4487 VSS 0.056945f
C3221 ASIG5V.n4488 VSS 0.056945f
C3222 ASIG5V.n4489 VSS 0.056945f
C3223 ASIG5V.n4490 VSS 0.056945f
C3224 ASIG5V.n4491 VSS 0.056945f
C3225 ASIG5V.n4492 VSS 0.056945f
C3226 ASIG5V.n4493 VSS 0.056945f
C3227 ASIG5V.n4494 VSS 0.056945f
C3228 ASIG5V.n4495 VSS 0.056945f
C3229 ASIG5V.n4496 VSS 0.056945f
C3230 ASIG5V.n4497 VSS 0.056945f
C3231 ASIG5V.n4498 VSS 0.056945f
C3232 ASIG5V.n4499 VSS 0.056945f
C3233 ASIG5V.n4500 VSS 0.056945f
C3234 ASIG5V.n4501 VSS 0.056945f
C3235 ASIG5V.n4502 VSS 0.056945f
C3236 ASIG5V.n4503 VSS 0.056945f
C3237 ASIG5V.n4504 VSS 0.056945f
C3238 ASIG5V.n4505 VSS 0.056945f
C3239 ASIG5V.n4506 VSS 0.056945f
C3240 ASIG5V.n4507 VSS 0.056945f
C3241 ASIG5V.n4508 VSS 0.056945f
C3242 ASIG5V.n4509 VSS 0.056945f
C3243 ASIG5V.n4510 VSS 0.056945f
C3244 ASIG5V.n4511 VSS 0.056945f
C3245 ASIG5V.n4512 VSS 0.056945f
C3246 ASIG5V.n4513 VSS 0.056945f
C3247 ASIG5V.n4514 VSS 0.056945f
C3248 ASIG5V.n4515 VSS 0.056945f
C3249 ASIG5V.n4516 VSS 0.056945f
C3250 ASIG5V.n4517 VSS 0.056945f
C3251 ASIG5V.n4518 VSS 0.056945f
C3252 ASIG5V.n4519 VSS 0.056945f
C3253 ASIG5V.n4520 VSS 0.056945f
C3254 ASIG5V.n4521 VSS 0.056945f
C3255 ASIG5V.n4522 VSS 0.056945f
C3256 ASIG5V.n4523 VSS 0.056945f
C3257 ASIG5V.n4524 VSS 0.056945f
C3258 ASIG5V.n4525 VSS 0.056945f
C3259 ASIG5V.n4526 VSS 0.056945f
C3260 ASIG5V.n4527 VSS 0.056945f
C3261 ASIG5V.n4528 VSS 0.056945f
C3262 ASIG5V.n4529 VSS 0.056945f
C3263 ASIG5V.n4530 VSS 0.056945f
C3264 ASIG5V.n4531 VSS 0.056945f
C3265 ASIG5V.n4532 VSS 0.056945f
C3266 ASIG5V.n4533 VSS 0.056945f
C3267 ASIG5V.n4534 VSS 0.056945f
C3268 ASIG5V.n4535 VSS 0.056945f
C3269 ASIG5V.n4536 VSS 0.056945f
C3270 ASIG5V.n4537 VSS 0.056945f
C3271 ASIG5V.n4538 VSS 0.056945f
C3272 ASIG5V.n4539 VSS 0.056945f
C3273 ASIG5V.n4540 VSS 0.056945f
C3274 ASIG5V.n4541 VSS 0.056945f
C3275 ASIG5V.n4542 VSS 0.056945f
C3276 ASIG5V.n4543 VSS 0.056945f
C3277 ASIG5V.n4544 VSS 0.056945f
C3278 ASIG5V.n4545 VSS 0.056945f
C3279 ASIG5V.n4546 VSS 0.056945f
C3280 ASIG5V.n4547 VSS 0.056945f
C3281 ASIG5V.n4548 VSS 0.056945f
C3282 ASIG5V.n4549 VSS 0.056945f
C3283 ASIG5V.n4550 VSS 0.056945f
C3284 ASIG5V.n4551 VSS 0.056945f
C3285 ASIG5V.n4552 VSS 0.056945f
C3286 ASIG5V.n4554 VSS 0.670332f
C3287 ASIG5V.n4555 VSS 0.909185f
C3288 ASIG5V.n4556 VSS 0.955415f
C3289 ASIG5V.n4557 VSS 0.076709f
C3290 ASIG5V.n4558 VSS 0.051589f
C3291 ASIG5V.n4559 VSS 0.051589f
C3292 ASIG5V.n4560 VSS 0.045056f
C3293 ASIG5V.n4561 VSS 0.063474f
C3294 ASIG5V.n4562 VSS 0.063474f
C3295 ASIG5V.n4563 VSS 0.055436f
C3296 ASIG5V.n4564 VSS 0.052746f
C3297 ASIG5V.n4565 VSS 0.047722f
C3298 ASIG5V.n4566 VSS 0.036092f
C3299 ASIG5V.n4567 VSS 0.036092f
C3300 ASIG5V.n4568 VSS 0.809021f
C3301 ASIG5V.n4569 VSS 0.909185f
C3302 ASIG5V.n4570 VSS 0.059753f
C3303 ASIG5V.n4571 VSS 0.059753f
C3304 ASIG5V.n4572 VSS 0.053336f
C3305 ASIG5V.n4573 VSS 0.07229f
C3306 ASIG5V.n4574 VSS 0.09726f
C3307 ASIG5V.n4575 VSS 0.092554f
C3308 ASIG5V.n4576 VSS 0.103688f
C3309 ASIG5V.n4577 VSS 0.103688f
C3310 ASIG5V.n4578 VSS 0.108961f
C3311 ASIG5V.n4579 VSS 0.072055f
C3312 ASIG5V.n4580 VSS 0.072055f
C3313 ASIG5V.n4581 VSS 0.0621f
C3314 ASIG5V.n4582 VSS 0.091386f
C3315 ASIG5V.n4583 VSS 0.081573f
C3316 ASIG5V.n4584 VSS 0.07229f
C3317 ASIG5V.n4585 VSS 0.052133f
C3318 ASIG5V.n4586 VSS 0.056945f
C3319 ASIG5V.n4587 VSS 0.056945f
C3320 ASIG5V.n4588 VSS 0.056945f
C3321 ASIG5V.n4589 VSS 0.056945f
C3322 ASIG5V.n4590 VSS 0.056945f
C3323 ASIG5V.n4591 VSS 0.056945f
C3324 ASIG5V.n4592 VSS 0.056945f
C3325 ASIG5V.n4593 VSS 0.056945f
C3326 ASIG5V.n4594 VSS 0.056945f
C3327 ASIG5V.n4595 VSS 0.056945f
C3328 ASIG5V.n4596 VSS 0.056945f
C3329 ASIG5V.n4597 VSS 0.056945f
C3330 ASIG5V.n4598 VSS 0.056945f
C3331 ASIG5V.n4599 VSS 0.056945f
C3332 ASIG5V.n4600 VSS 0.056945f
C3333 ASIG5V.n4601 VSS 0.056945f
C3334 ASIG5V.n4602 VSS 0.056945f
C3335 ASIG5V.n4603 VSS 0.056945f
C3336 ASIG5V.n4604 VSS 0.056945f
C3337 ASIG5V.n4605 VSS 0.056945f
C3338 ASIG5V.n4606 VSS 0.056945f
C3339 ASIG5V.n4607 VSS 0.056945f
C3340 ASIG5V.n4608 VSS 0.056945f
C3341 ASIG5V.n4609 VSS 0.056945f
C3342 ASIG5V.n4610 VSS 0.056945f
C3343 ASIG5V.n4611 VSS 0.056945f
C3344 ASIG5V.n4612 VSS 0.056945f
C3345 ASIG5V.n4613 VSS 0.056945f
C3346 ASIG5V.n4614 VSS 0.056945f
C3347 ASIG5V.n4615 VSS 0.056945f
C3348 ASIG5V.n4616 VSS 0.056945f
C3349 ASIG5V.n4617 VSS 0.056945f
C3350 ASIG5V.n4618 VSS 0.056945f
C3351 ASIG5V.n4619 VSS 0.056945f
C3352 ASIG5V.n4620 VSS 0.056945f
C3353 ASIG5V.n4621 VSS 0.056945f
C3354 ASIG5V.n4622 VSS 0.056945f
C3355 ASIG5V.n4623 VSS 0.056945f
C3356 ASIG5V.n4624 VSS 0.056945f
C3357 ASIG5V.n4625 VSS 0.056945f
C3358 ASIG5V.n4626 VSS 0.056945f
C3359 ASIG5V.n4627 VSS 0.056945f
C3360 ASIG5V.n4628 VSS 0.056945f
C3361 ASIG5V.n4629 VSS 0.056945f
C3362 ASIG5V.n4630 VSS 0.056945f
C3363 ASIG5V.n4631 VSS 0.056945f
C3364 ASIG5V.n4632 VSS 0.056945f
C3365 ASIG5V.n4633 VSS 0.056945f
C3366 ASIG5V.n4634 VSS 0.056945f
C3367 ASIG5V.n4635 VSS 0.056945f
C3368 ASIG5V.n4636 VSS 0.056945f
C3369 ASIG5V.n4637 VSS 0.056945f
C3370 ASIG5V.n4638 VSS 0.056945f
C3371 ASIG5V.n4639 VSS 0.056945f
C3372 ASIG5V.n4640 VSS 0.056945f
C3373 ASIG5V.n4641 VSS 0.056945f
C3374 ASIG5V.n4642 VSS 0.056945f
C3375 ASIG5V.n4643 VSS 0.056945f
C3376 ASIG5V.n4644 VSS 0.056945f
C3377 ASIG5V.n4645 VSS 0.056945f
C3378 ASIG5V.n4646 VSS 0.056945f
C3379 ASIG5V.n4647 VSS 0.056945f
C3380 ASIG5V.n4648 VSS 0.056945f
C3381 ASIG5V.n4649 VSS 0.056945f
C3382 ASIG5V.n4650 VSS 0.056945f
C3383 ASIG5V.n4651 VSS 0.056945f
C3384 ASIG5V.n4652 VSS 0.056945f
C3385 ASIG5V.n4653 VSS 0.056945f
C3386 ASIG5V.n4654 VSS 0.056945f
C3387 ASIG5V.n4655 VSS 0.056945f
C3388 ASIG5V.n4656 VSS 0.056945f
C3389 ASIG5V.n4657 VSS 0.056945f
C3390 ASIG5V.n4658 VSS 0.056945f
C3391 ASIG5V.n4659 VSS 0.056945f
C3392 ASIG5V.n4660 VSS 0.056945f
C3393 ASIG5V.n4661 VSS 0.056945f
C3394 ASIG5V.n4662 VSS 0.056945f
C3395 ASIG5V.n4663 VSS 0.056945f
C3396 ASIG5V.n4664 VSS 0.056945f
C3397 ASIG5V.n4665 VSS 0.056945f
C3398 ASIG5V.n4666 VSS 0.056945f
C3399 ASIG5V.n4667 VSS 0.056945f
C3400 ASIG5V.n4668 VSS 0.056945f
C3401 ASIG5V.n4669 VSS 0.056945f
C3402 ASIG5V.n4670 VSS 0.056945f
C3403 ASIG5V.n4671 VSS 0.056945f
C3404 ASIG5V.n4672 VSS 0.056945f
C3405 ASIG5V.n4673 VSS 0.056945f
C3406 ASIG5V.n4674 VSS 0.056945f
C3407 ASIG5V.n4675 VSS 0.056945f
C3408 ASIG5V.n4676 VSS 0.056945f
C3409 ASIG5V.n4677 VSS 0.056945f
C3410 ASIG5V.n4678 VSS 0.056945f
C3411 ASIG5V.n4679 VSS 0.056945f
C3412 ASIG5V.n4680 VSS 0.056945f
C3413 ASIG5V.n4681 VSS 0.056945f
C3414 ASIG5V.n4682 VSS 0.056945f
C3415 ASIG5V.n4683 VSS 0.056945f
C3416 ASIG5V.n4684 VSS 0.056945f
C3417 ASIG5V.n4685 VSS 0.056945f
C3418 ASIG5V.n4686 VSS 0.056945f
C3419 ASIG5V.n4687 VSS 0.056945f
C3420 ASIG5V.n4688 VSS 0.056945f
C3421 ASIG5V.n4689 VSS 0.056945f
C3422 ASIG5V.n4690 VSS 0.056945f
C3423 ASIG5V.n4691 VSS 0.056945f
C3424 ASIG5V.n4692 VSS 0.056945f
C3425 ASIG5V.n4693 VSS 0.056945f
C3426 ASIG5V.n4694 VSS 0.056945f
C3427 ASIG5V.n4695 VSS 0.056945f
C3428 ASIG5V.n4696 VSS 0.056945f
C3429 ASIG5V.n4697 VSS 0.056945f
C3430 ASIG5V.n4698 VSS 0.056945f
C3431 ASIG5V.n4699 VSS 0.056945f
C3432 ASIG5V.n4700 VSS 0.056945f
C3433 ASIG5V.n4701 VSS 0.056945f
C3434 ASIG5V.n4702 VSS 0.056945f
C3435 ASIG5V.n4703 VSS 0.056945f
C3436 ASIG5V.n4704 VSS 0.056945f
C3437 ASIG5V.n4705 VSS 0.056945f
C3438 ASIG5V.n4706 VSS 0.056945f
C3439 ASIG5V.n4707 VSS 0.056945f
C3440 ASIG5V.n4708 VSS 0.056945f
C3441 ASIG5V.n4709 VSS 0.056945f
C3442 ASIG5V.n4710 VSS 0.056945f
C3443 ASIG5V.n4711 VSS 0.056945f
C3444 ASIG5V.n4712 VSS 0.056945f
C3445 ASIG5V.n4713 VSS 0.056945f
C3446 ASIG5V.n4714 VSS 0.056945f
C3447 ASIG5V.n4715 VSS 0.056945f
C3448 ASIG5V.n4716 VSS 0.056945f
C3449 ASIG5V.n4717 VSS 0.056945f
C3450 ASIG5V.n4718 VSS 0.056945f
C3451 ASIG5V.n4719 VSS 0.056945f
C3452 ASIG5V.n4720 VSS 0.056945f
C3453 ASIG5V.n4721 VSS 0.056945f
C3454 ASIG5V.n4722 VSS 0.056945f
C3455 ASIG5V.n4723 VSS 0.056945f
C3456 ASIG5V.n4724 VSS 0.056945f
C3457 ASIG5V.n4725 VSS 0.056945f
C3458 ASIG5V.n4726 VSS 0.056945f
C3459 ASIG5V.n4727 VSS 0.056945f
C3460 ASIG5V.n4728 VSS 0.056945f
C3461 ASIG5V.n4729 VSS 0.056945f
C3462 ASIG5V.n4730 VSS 0.056945f
C3463 ASIG5V.n4731 VSS 0.056945f
C3464 ASIG5V.n4732 VSS 0.056945f
C3465 ASIG5V.n4733 VSS 0.056945f
C3466 ASIG5V.n4734 VSS 0.056945f
C3467 ASIG5V.n4735 VSS 0.056945f
C3468 ASIG5V.n4736 VSS 0.056945f
C3469 ASIG5V.n4737 VSS 0.056945f
C3470 ASIG5V.n4738 VSS 0.056945f
C3471 ASIG5V.n4739 VSS 0.056945f
C3472 ASIG5V.n4740 VSS 0.056945f
C3473 ASIG5V.n4741 VSS 0.056945f
C3474 ASIG5V.n4742 VSS 0.056945f
C3475 ASIG5V.n4743 VSS 0.056945f
C3476 ASIG5V.n4744 VSS 0.056945f
C3477 ASIG5V.n4745 VSS 0.056945f
C3478 ASIG5V.n4746 VSS 0.056945f
C3479 ASIG5V.n4747 VSS 0.056945f
C3480 ASIG5V.n4748 VSS 0.056945f
C3481 ASIG5V.n4749 VSS 0.056945f
C3482 ASIG5V.n4750 VSS 0.056945f
C3483 ASIG5V.n4751 VSS 0.056945f
C3484 ASIG5V.n4752 VSS 0.056945f
C3485 ASIG5V.n4753 VSS 0.056945f
C3486 ASIG5V.n4754 VSS 0.056945f
C3487 ASIG5V.n4755 VSS 0.056945f
C3488 ASIG5V.n4756 VSS 0.056945f
C3489 ASIG5V.n4757 VSS 0.056945f
C3490 ASIG5V.n4758 VSS 0.056945f
C3491 ASIG5V.n4759 VSS 0.056945f
C3492 ASIG5V.n4760 VSS 0.056945f
C3493 ASIG5V.n4761 VSS 0.056945f
C3494 ASIG5V.n4762 VSS 0.056945f
C3495 ASIG5V.n4763 VSS 0.056945f
C3496 ASIG5V.n4764 VSS 0.056945f
C3497 ASIG5V.n4765 VSS 0.056945f
C3498 ASIG5V.n4766 VSS 0.056945f
C3499 ASIG5V.n4767 VSS 0.056945f
C3500 ASIG5V.n4768 VSS 0.056945f
C3501 ASIG5V.n4769 VSS 0.056945f
C3502 ASIG5V.n4770 VSS 0.036092f
C3503 ASIG5V.n4771 VSS 0.036092f
C3504 ASIG5V.n4772 VSS 0.955416f
C3505 ASIG5V.n4773 VSS 0.036092f
C3506 ASIG5V.n4775 VSS 0.346723f
C3507 ASIG5V.n4776 VSS 0.824431f
C3508 ASIG5V.n4777 VSS 0.878365f
C3509 ASIG5V.n4778 VSS 0.044567f
C3510 ASIG5V.n4779 VSS 0.044567f
C3511 ASIG5V.n4780 VSS 0.038923f
C3512 ASIG5V.n4781 VSS 0.052746f
C3513 ASIG5V.n4782 VSS 0.061569f
C3514 ASIG5V.n4783 VSS 0.066287f
C3515 ASIG5V.n4784 VSS 0.075898f
C3516 ASIG5V.n4785 VSS 0.075898f
C3517 ASIG5V.n4786 VSS 0.955415f
C3518 ASIG5V.n4787 VSS 1.0941f
C3519 ASIG5V.n4788 VSS 0.108961f
C3520 ASIG5V.n4789 VSS 0.084357f
C3521 ASIG5V.n4790 VSS 0.084357f
C3522 ASIG5V.n4791 VSS 0.075298f
C3523 ASIG5V.n4792 VSS 0.07229f
C3524 ASIG5V.n4793 VSS 0.086279f
C3525 ASIG5V.n4794 VSS 0.09726f
C3526 ASIG5V.n4795 VSS 0.070592f
C3527 ASIG5V.n4796 VSS 0.079084f
C3528 ASIG5V.n4797 VSS 0.079084f
C3529 ASIG5V.n4798 VSS 0.547052f
C3530 ASIG5V.n4799 VSS 0.955415f
C3531 ASIG5V.n4800 VSS 0.039165f
C3532 ASIG5V.n4801 VSS 0.039165f
C3533 ASIG5V.n4802 VSS 0.034205f
C3534 ASIG5V.n4803 VSS 0.066995f
C3535 ASIG5V.n4804 VSS 0.060154f
C3536 ASIG5V.n4805 VSS 0.068876f
C3537 ASIG5V.n4806 VSS 0.068876f
C3538 ASIG5V.n4807 VSS 0.955415f
C3539 ASIG5V.n4808 VSS 0.385247f
C3540 ASIG5V.n4809 VSS 0.096659f
C3541 ASIG5V.n4810 VSS 0.0621f
C3542 ASIG5V.n4811 VSS 0.066782f
C3543 ASIG5V.n4812 VSS 0.059611f
C3544 ASIG5V.n4813 VSS 0.066782f
C3545 ASIG5V.n4814 VSS 0.0621f
C3546 ASIG5V.n4815 VSS 0.036092f
C3547 ASIG5V.n4816 VSS 0.052133f
C3548 ASIG5V.n4817 VSS 0.056945f
C3549 ASIG5V.n4818 VSS 0.056945f
C3550 ASIG5V.n4819 VSS 0.056945f
C3551 ASIG5V.n4820 VSS 0.056945f
C3552 ASIG5V.n4822 VSS 0.056945f
C3553 ASIG5V.n4823 VSS 0.056945f
C3554 ASIG5V.n4824 VSS 0.056945f
C3555 ASIG5V.n4826 VSS 0.056945f
C3556 ASIG5V.n4827 VSS 0.056945f
C3557 ASIG5V.n4828 VSS 0.056945f
C3558 ASIG5V.n4829 VSS 0.056945f
C3559 ASIG5V.n4830 VSS 0.056945f
C3560 ASIG5V.n4831 VSS 0.056945f
C3561 ASIG5V.n4832 VSS 0.056945f
C3562 ASIG5V.n4834 VSS 0.056945f
C3563 ASIG5V.n4835 VSS 0.056945f
C3564 ASIG5V.n4836 VSS 0.056945f
C3565 ASIG5V.n4838 VSS 0.056945f
C3566 ASIG5V.n4839 VSS 0.056945f
C3567 ASIG5V.n4840 VSS 0.056945f
C3568 ASIG5V.n4841 VSS 0.056945f
C3569 ASIG5V.n4842 VSS 0.056945f
C3570 ASIG5V.n4843 VSS 0.056945f
C3571 ASIG5V.n4844 VSS 0.056945f
C3572 ASIG5V.n4846 VSS 0.056945f
C3573 ASIG5V.n4847 VSS 0.056945f
C3574 ASIG5V.n4848 VSS 0.056945f
C3575 ASIG5V.n4850 VSS 0.056945f
C3576 ASIG5V.n4851 VSS 0.056945f
C3577 ASIG5V.n4852 VSS 0.056945f
C3578 ASIG5V.n4853 VSS 0.056945f
C3579 ASIG5V.n4854 VSS 0.056945f
C3580 ASIG5V.n4855 VSS 0.056945f
C3581 ASIG5V.n4856 VSS 0.056945f
C3582 ASIG5V.n4858 VSS 0.056945f
C3583 ASIG5V.n4859 VSS 0.056945f
C3584 ASIG5V.n4860 VSS 0.056945f
C3585 ASIG5V.n4862 VSS 0.056945f
C3586 ASIG5V.n4863 VSS 0.056945f
C3587 ASIG5V.n4864 VSS 0.056945f
C3588 ASIG5V.n4865 VSS 0.056945f
C3589 ASIG5V.n4866 VSS 0.056945f
C3590 ASIG5V.n4867 VSS 0.056945f
C3591 ASIG5V.n4868 VSS 0.056945f
C3592 ASIG5V.n4870 VSS 0.056945f
C3593 ASIG5V.n4871 VSS 0.056945f
C3594 ASIG5V.n4872 VSS 0.056945f
C3595 ASIG5V.n4874 VSS 0.056945f
C3596 ASIG5V.n4875 VSS 0.056945f
C3597 ASIG5V.n4876 VSS 0.056945f
C3598 ASIG5V.n4877 VSS 0.056945f
C3599 ASIG5V.n4878 VSS 0.056945f
C3600 ASIG5V.n4879 VSS 0.056945f
C3601 ASIG5V.n4880 VSS 0.056945f
C3602 ASIG5V.n4882 VSS 0.056945f
C3603 ASIG5V.n4883 VSS 0.056945f
C3604 ASIG5V.n4884 VSS 0.056945f
C3605 ASIG5V.n4886 VSS 0.056945f
C3606 ASIG5V.n4887 VSS 0.056945f
C3607 ASIG5V.n4888 VSS 0.056945f
C3608 ASIG5V.n4889 VSS 0.056945f
C3609 ASIG5V.n4890 VSS 0.056945f
C3610 ASIG5V.n4891 VSS 0.056945f
C3611 ASIG5V.n4892 VSS 0.056945f
C3612 ASIG5V.n4894 VSS 0.056945f
C3613 ASIG5V.n4895 VSS 0.056945f
C3614 ASIG5V.n4896 VSS 0.056945f
C3615 ASIG5V.n4898 VSS 0.056945f
C3616 ASIG5V.n4899 VSS 0.056945f
C3617 ASIG5V.n4900 VSS 0.056945f
C3618 ASIG5V.n4901 VSS 0.056945f
C3619 ASIG5V.n4902 VSS 0.056945f
C3620 ASIG5V.n4903 VSS 0.056945f
C3621 ASIG5V.n4904 VSS 0.056945f
C3622 ASIG5V.n4906 VSS 0.056945f
C3623 ASIG5V.n4907 VSS 0.056945f
C3624 ASIG5V.n4908 VSS 0.056945f
C3625 ASIG5V.n4910 VSS 0.056945f
C3626 ASIG5V.n4911 VSS 0.056945f
C3627 ASIG5V.n4912 VSS 0.056945f
C3628 ASIG5V.n4913 VSS 0.056945f
C3629 ASIG5V.n4914 VSS 0.056945f
C3630 ASIG5V.n4915 VSS 0.056945f
C3631 ASIG5V.n4916 VSS 0.056945f
C3632 ASIG5V.n4918 VSS 0.056945f
C3633 ASIG5V.n4919 VSS 0.056945f
C3634 ASIG5V.n4920 VSS 0.056945f
C3635 ASIG5V.n4922 VSS 0.056945f
C3636 ASIG5V.n4923 VSS 0.056945f
C3637 ASIG5V.n4924 VSS 0.056945f
C3638 ASIG5V.n4925 VSS 0.056945f
C3639 ASIG5V.n4926 VSS 0.056945f
C3640 ASIG5V.n4927 VSS 0.056945f
C3641 ASIG5V.n4928 VSS 0.056945f
C3642 ASIG5V.n4930 VSS 0.056945f
C3643 ASIG5V.n4931 VSS 0.056945f
C3644 ASIG5V.n4932 VSS 0.056945f
C3645 ASIG5V.n4934 VSS 0.056945f
C3646 ASIG5V.n4935 VSS 0.056945f
C3647 ASIG5V.n4936 VSS 0.056945f
C3648 ASIG5V.n4937 VSS 0.056945f
C3649 ASIG5V.n4938 VSS 0.056945f
C3650 ASIG5V.n4939 VSS 0.056945f
C3651 ASIG5V.n4940 VSS 0.056945f
C3652 ASIG5V.n4942 VSS 0.056945f
C3653 ASIG5V.n4943 VSS 0.056945f
C3654 ASIG5V.n4944 VSS 0.056945f
C3655 ASIG5V.n4946 VSS 0.056945f
C3656 ASIG5V.n4947 VSS 0.056945f
C3657 ASIG5V.n4948 VSS 0.056945f
C3658 ASIG5V.n4949 VSS 0.056945f
C3659 ASIG5V.n4950 VSS 0.056945f
C3660 ASIG5V.n4951 VSS 0.056945f
C3661 ASIG5V.n4952 VSS 0.056945f
C3662 ASIG5V.n4954 VSS 0.056945f
C3663 ASIG5V.n4955 VSS 0.056945f
C3664 ASIG5V.n4956 VSS 0.056945f
C3665 ASIG5V.n4958 VSS 0.056945f
C3666 ASIG5V.n4959 VSS 0.056945f
C3667 ASIG5V.n4960 VSS 0.056945f
C3668 ASIG5V.n4961 VSS 0.056945f
C3669 ASIG5V.n4962 VSS 0.056945f
C3670 ASIG5V.n4963 VSS 0.056945f
C3671 ASIG5V.n4964 VSS 0.056945f
C3672 ASIG5V.n4966 VSS 0.056945f
C3673 ASIG5V.n4967 VSS 0.056945f
C3674 ASIG5V.n4968 VSS 0.056945f
C3675 ASIG5V.n4970 VSS 0.056945f
C3676 ASIG5V.n4971 VSS 0.056945f
C3677 ASIG5V.n4972 VSS 0.056945f
C3678 ASIG5V.n4973 VSS 0.056945f
C3679 ASIG5V.n4974 VSS 0.056945f
C3680 ASIG5V.n4975 VSS 0.056945f
C3681 ASIG5V.n4976 VSS 0.056945f
C3682 ASIG5V.n4978 VSS 0.056945f
C3683 ASIG5V.n4979 VSS 0.056945f
C3684 ASIG5V.n4980 VSS 0.056945f
C3685 ASIG5V.n4982 VSS 0.056945f
C3686 ASIG5V.n4983 VSS 0.056945f
C3687 ASIG5V.n4984 VSS 0.056945f
C3688 ASIG5V.n4985 VSS 0.056945f
C3689 ASIG5V.n4986 VSS 0.056945f
C3690 ASIG5V.n4987 VSS 0.056945f
C3691 ASIG5V.n4988 VSS 0.056945f
C3692 ASIG5V.n4990 VSS 0.056945f
C3693 ASIG5V.n4991 VSS 0.056945f
C3694 ASIG5V.n4992 VSS 0.056945f
C3695 ASIG5V.n4994 VSS 0.056945f
C3696 ASIG5V.n4995 VSS 0.056945f
C3697 ASIG5V.n4996 VSS 0.056945f
C3698 ASIG5V.n4997 VSS 0.056945f
C3699 ASIG5V.n4998 VSS 0.056945f
C3700 ASIG5V.n4999 VSS 0.056945f
C3701 ASIG5V.n5000 VSS 0.056945f
C3702 ASIG5V.n5002 VSS 0.056945f
C3703 ASIG5V.n5003 VSS 0.056945f
C3704 ASIG5V.n5004 VSS 0.056945f
C3705 ASIG5V.n5006 VSS 0.056945f
C3706 ASIG5V.n5007 VSS 0.056945f
C3707 ASIG5V.n5008 VSS 0.056945f
C3708 ASIG5V.n5009 VSS 0.056945f
C3709 ASIG5V.n5010 VSS 0.056945f
C3710 ASIG5V.n5011 VSS 0.056945f
C3711 ASIG5V.n5012 VSS 0.056945f
C3712 ASIG5V.n5014 VSS 0.056945f
C3713 ASIG5V.n5015 VSS 0.056945f
C3714 ASIG5V.n5016 VSS 0.056945f
C3715 ASIG5V.n5018 VSS 0.056945f
C3716 ASIG5V.n5019 VSS 0.056945f
C3717 ASIG5V.n5020 VSS 0.056945f
C3718 ASIG5V.n5021 VSS 0.056945f
C3719 ASIG5V.n5022 VSS 0.056945f
C3720 ASIG5V.n5023 VSS 0.056945f
C3721 ASIG5V.n5024 VSS 0.056945f
C3722 ASIG5V.n5026 VSS 0.056945f
C3723 ASIG5V.n5027 VSS 0.056945f
C3724 ASIG5V.n5028 VSS 0.056945f
C3725 ASIG5V.n5030 VSS 0.056945f
C3726 ASIG5V.n5031 VSS 0.056945f
C3727 ASIG5V.n5032 VSS 0.056945f
C3728 ASIG5V.n5033 VSS 0.056945f
C3729 ASIG5V.n5034 VSS 0.056945f
C3730 ASIG5V.n5035 VSS 0.056945f
C3731 ASIG5V.n5036 VSS 0.056945f
C3732 ASIG5V.n5038 VSS 0.056945f
C3733 ASIG5V.n5039 VSS 0.056945f
C3734 ASIG5V.n5040 VSS 0.056945f
C3735 ASIG5V.n5042 VSS 0.056945f
C3736 ASIG5V.n5043 VSS 0.056945f
C3737 ASIG5V.n5044 VSS 0.056945f
C3738 ASIG5V.n5045 VSS 0.056945f
C3739 ASIG5V.n5046 VSS 0.056945f
C3740 ASIG5V.n5047 VSS 0.056945f
C3741 ASIG5V.n5048 VSS 0.056945f
C3742 ASIG5V.n5050 VSS 0.056945f
C3743 ASIG5V.n5051 VSS 0.056945f
C3744 ASIG5V.n5052 VSS 0.056945f
C3745 ASIG5V.n5054 VSS 0.056945f
C3746 ASIG5V.n5055 VSS 0.056945f
C3747 ASIG5V.n5056 VSS 0.056945f
C3748 ASIG5V.n5057 VSS 0.056945f
C3749 ASIG5V.n5058 VSS 0.047722f
C3750 ASIG5V.n5059 VSS 0.056945f
C3751 ASIG5V.n5060 VSS 0.056945f
C3752 ASIG5V.n5061 VSS 0.056945f
C3753 ASIG5V.n5063 VSS 0.036092f
C3754 ASIG5V.n5064 VSS 0.947711f
C3755 ASIG5V.n5065 VSS 0.392953f
C3756 ASIG5V.n5066 VSS 0.046187f
C3757 ASIG5V.n5067 VSS 0.046187f
C3758 ASIG5V.n5068 VSS 0.040338f
C3759 ASIG5V.n5069 VSS 0.066995f
C3760 ASIG5V.n5070 VSS 0.047722f
C3761 ASIG5V.n5071 VSS 0.066995f
C3762 ASIG5V.n5072 VSS 0.076709f
C3763 ASIG5V.n5073 VSS 0.076709f
C3764 ASIG5V.n5074 VSS 0.932301f
C3765 ASIG5V.n5116 VSS 0.036092f
C3766 ASIG5V.n5117 VSS 0.955415f
C3767 ASIG5V.n5118 VSS 0.108961f
C3768 ASIG5V.n5119 VSS 0.108961f
C3769 ASIG5V.n5120 VSS 0.07229f
C3770 ASIG5V.n5121 VSS 0.0621f
C3771 ASIG5V.n5122 VSS 0.0621f
C3772 ASIG5V.n5123 VSS 0.292788f
C3773 ASIG5V.n5165 VSS 0.036092f
C3774 ASIG5V.n5166 VSS 0.154098f
C3775 ASIG5V.n5167 VSS 0.045974f
C3776 ASIG5V.n5168 VSS 0.036092f
C3777 ASIG5V.n5169 VSS 1.05558f
C3778 ASIG5V.n5170 VSS 0.701152f
C3779 ASIG5V.n5171 VSS 0.056945f
C3780 ASIG5V.n5172 VSS 0.056945f
C3781 ASIG5V.n5173 VSS 0.056945f
C3782 ASIG5V.n5174 VSS 0.056945f
C3783 ASIG5V.n5175 VSS 0.056945f
C3784 ASIG5V.n5176 VSS 0.056945f
C3785 ASIG5V.n5177 VSS 0.056945f
C3786 ASIG5V.n5178 VSS 0.056945f
C3787 ASIG5V.n5179 VSS 0.056945f
C3788 ASIG5V.n5180 VSS 0.056945f
C3789 ASIG5V.n5181 VSS 0.056945f
C3790 ASIG5V.n5182 VSS 0.056945f
C3791 ASIG5V.n5183 VSS 0.056945f
C3792 ASIG5V.n5184 VSS 0.056945f
C3793 ASIG5V.n5185 VSS 0.056945f
C3794 ASIG5V.n5186 VSS 0.056945f
C3795 ASIG5V.n5187 VSS 0.056945f
C3796 ASIG5V.n5188 VSS 0.056945f
C3797 ASIG5V.n5189 VSS 0.056945f
C3798 ASIG5V.n5190 VSS 0.056945f
C3799 ASIG5V.n5191 VSS 0.056945f
C3800 ASIG5V.n5192 VSS 0.056945f
C3801 ASIG5V.n5193 VSS 0.056945f
C3802 ASIG5V.n5194 VSS 0.056945f
C3803 ASIG5V.n5195 VSS 0.056945f
C3804 ASIG5V.n5196 VSS 0.056945f
C3805 ASIG5V.n5197 VSS 0.056945f
C3806 ASIG5V.n5198 VSS 0.056945f
C3807 ASIG5V.n5199 VSS 0.056945f
C3808 ASIG5V.n5200 VSS 0.056945f
C3809 ASIG5V.n5201 VSS 0.056945f
C3810 ASIG5V.n5202 VSS 0.056945f
C3811 ASIG5V.n5203 VSS 0.056945f
C3812 ASIG5V.n5204 VSS 0.056945f
C3813 ASIG5V.n5205 VSS 0.056945f
C3814 ASIG5V.n5206 VSS 0.056945f
C3815 ASIG5V.n5207 VSS 0.056945f
C3816 ASIG5V.n5208 VSS 0.056945f
C3817 ASIG5V.n5209 VSS 0.056945f
C3818 ASIG5V.n5210 VSS 0.056945f
C3819 ASIG5V.n5212 VSS 0.056945f
C3820 ASIG5V.n5213 VSS 0.056945f
C3821 ASIG5V.n5214 VSS 0.036092f
C3822 ASIG5V.n5215 VSS 0.052133f
C3823 ASIG5V.n5216 VSS 0.056945f
C3824 ASIG5V.n5217 VSS 0.056945f
C3825 ASIG5V.n5218 VSS 0.056945f
C3826 ASIG5V.n5219 VSS 0.056945f
C3827 ASIG5V.n5221 VSS 0.056945f
C3828 ASIG5V.n5222 VSS 0.056945f
C3829 ASIG5V.n5223 VSS 0.056945f
C3830 ASIG5V.n5225 VSS 0.056945f
C3831 ASIG5V.n5226 VSS 0.056945f
C3832 ASIG5V.n5227 VSS 0.056945f
C3833 ASIG5V.n5228 VSS 0.056945f
C3834 ASIG5V.n5229 VSS 0.056945f
C3835 ASIG5V.n5230 VSS 0.056945f
C3836 ASIG5V.n5231 VSS 0.056945f
C3837 ASIG5V.n5233 VSS 0.056945f
C3838 ASIG5V.n5234 VSS 0.056945f
C3839 ASIG5V.n5235 VSS 0.056945f
C3840 ASIG5V.n5237 VSS 0.056945f
C3841 ASIG5V.n5238 VSS 0.056945f
C3842 ASIG5V.n5239 VSS 0.056945f
C3843 ASIG5V.n5240 VSS 0.056945f
C3844 ASIG5V.n5241 VSS 0.056945f
C3845 ASIG5V.n5242 VSS 0.056945f
C3846 ASIG5V.n5243 VSS 0.056945f
C3847 ASIG5V.n5245 VSS 0.056945f
C3848 ASIG5V.n5246 VSS 0.056945f
C3849 ASIG5V.n5247 VSS 0.056945f
C3850 ASIG5V.n5249 VSS 0.056945f
C3851 ASIG5V.n5250 VSS 0.056945f
C3852 ASIG5V.n5251 VSS 0.056945f
C3853 ASIG5V.n5252 VSS 0.056945f
C3854 ASIG5V.n5253 VSS 0.056945f
C3855 ASIG5V.n5254 VSS 0.056945f
C3856 ASIG5V.n5255 VSS 0.056945f
C3857 ASIG5V.n5257 VSS 0.056945f
C3858 ASIG5V.n5258 VSS 0.056945f
C3859 ASIG5V.n5259 VSS 0.056945f
C3860 ASIG5V.n5261 VSS 0.056945f
C3861 ASIG5V.n5262 VSS 0.056945f
C3862 ASIG5V.n5263 VSS 0.056945f
C3863 ASIG5V.n5264 VSS 0.056945f
C3864 ASIG5V.n5265 VSS 0.056945f
C3865 ASIG5V.n5266 VSS 0.056945f
C3866 ASIG5V.n5267 VSS 0.056945f
C3867 ASIG5V.n5269 VSS 0.056945f
C3868 ASIG5V.n5270 VSS 0.056945f
C3869 ASIG5V.n5271 VSS 0.056945f
C3870 ASIG5V.n5273 VSS 0.056945f
C3871 ASIG5V.n5274 VSS 0.056945f
C3872 ASIG5V.n5275 VSS 0.056945f
C3873 ASIG5V.n5276 VSS 0.056945f
C3874 ASIG5V.n5277 VSS 0.056945f
C3875 ASIG5V.n5278 VSS 0.056945f
C3876 ASIG5V.n5279 VSS 0.056945f
C3877 ASIG5V.n5281 VSS 0.056945f
C3878 ASIG5V.n5282 VSS 0.056945f
C3879 ASIG5V.n5283 VSS 0.056945f
C3880 ASIG5V.n5285 VSS 0.056945f
C3881 ASIG5V.n5286 VSS 0.056945f
C3882 ASIG5V.n5287 VSS 0.056945f
C3883 ASIG5V.n5288 VSS 0.056945f
C3884 ASIG5V.n5289 VSS 0.056945f
C3885 ASIG5V.n5290 VSS 0.056945f
C3886 ASIG5V.n5291 VSS 0.056945f
C3887 ASIG5V.n5293 VSS 0.056945f
C3888 ASIG5V.n5294 VSS 0.056945f
C3889 ASIG5V.n5295 VSS 0.056945f
C3890 ASIG5V.n5297 VSS 0.056945f
C3891 ASIG5V.n5298 VSS 0.056945f
C3892 ASIG5V.n5299 VSS 0.056945f
C3893 ASIG5V.n5300 VSS 0.056945f
C3894 ASIG5V.n5301 VSS 0.056945f
C3895 ASIG5V.n5302 VSS 0.056945f
C3896 ASIG5V.n5303 VSS 0.056945f
C3897 ASIG5V.n5305 VSS 0.056945f
C3898 ASIG5V.n5306 VSS 0.056945f
C3899 ASIG5V.n5307 VSS 0.056945f
C3900 ASIG5V.n5309 VSS 0.056945f
C3901 ASIG5V.n5310 VSS 0.056945f
C3902 ASIG5V.n5311 VSS 0.056945f
C3903 ASIG5V.n5312 VSS 0.056945f
C3904 ASIG5V.n5313 VSS 0.056945f
C3905 ASIG5V.n5314 VSS 0.056945f
C3906 ASIG5V.n5315 VSS 0.056945f
C3907 ASIG5V.n5317 VSS 0.056945f
C3908 ASIG5V.n5318 VSS 0.056945f
C3909 ASIG5V.n5319 VSS 0.056945f
C3910 ASIG5V.n5321 VSS 0.056945f
C3911 ASIG5V.n5322 VSS 0.056945f
C3912 ASIG5V.n5323 VSS 0.056945f
C3913 ASIG5V.n5324 VSS 0.056945f
C3914 ASIG5V.n5325 VSS 0.056945f
C3915 ASIG5V.n5326 VSS 0.056945f
C3916 ASIG5V.n5327 VSS 0.056945f
C3917 ASIG5V.n5329 VSS 0.056945f
C3918 ASIG5V.n5330 VSS 0.056945f
C3919 ASIG5V.n5331 VSS 0.056945f
C3920 ASIG5V.n5333 VSS 0.056945f
C3921 ASIG5V.n5334 VSS 0.056945f
C3922 ASIG5V.n5335 VSS 0.056945f
C3923 ASIG5V.n5336 VSS 0.056945f
C3924 ASIG5V.n5337 VSS 0.056945f
C3925 ASIG5V.n5338 VSS 0.056945f
C3926 ASIG5V.n5339 VSS 0.056945f
C3927 ASIG5V.n5341 VSS 0.056945f
C3928 ASIG5V.n5342 VSS 0.056945f
C3929 ASIG5V.n5343 VSS 0.056945f
C3930 ASIG5V.n5345 VSS 0.056945f
C3931 ASIG5V.n5346 VSS 0.056945f
C3932 ASIG5V.n5347 VSS 0.056945f
C3933 ASIG5V.n5348 VSS 0.056945f
C3934 ASIG5V.n5349 VSS 0.056945f
C3935 ASIG5V.n5350 VSS 0.056945f
C3936 ASIG5V.n5351 VSS 0.056945f
C3937 ASIG5V.n5353 VSS 0.056945f
C3938 ASIG5V.n5354 VSS 0.056945f
C3939 ASIG5V.n5355 VSS 0.056945f
C3940 ASIG5V.n5357 VSS 0.056945f
C3941 ASIG5V.n5358 VSS 0.056945f
C3942 ASIG5V.n5359 VSS 0.056945f
C3943 ASIG5V.n5360 VSS 0.056945f
C3944 ASIG5V.n5361 VSS 0.056945f
C3945 ASIG5V.n5362 VSS 0.056945f
C3946 ASIG5V.n5363 VSS 0.056945f
C3947 ASIG5V.n5365 VSS 0.056945f
C3948 ASIG5V.n5366 VSS 0.056945f
C3949 ASIG5V.n5367 VSS 0.056945f
C3950 ASIG5V.n5369 VSS 0.056945f
C3951 ASIG5V.n5370 VSS 0.056945f
C3952 ASIG5V.n5371 VSS 0.056945f
C3953 ASIG5V.n5372 VSS 0.056945f
C3954 ASIG5V.n5373 VSS 0.056945f
C3955 ASIG5V.n5374 VSS 0.056945f
C3956 ASIG5V.n5375 VSS 0.056945f
C3957 ASIG5V.n5377 VSS 0.056945f
C3958 ASIG5V.n5378 VSS 0.056945f
C3959 ASIG5V.n5379 VSS 0.056945f
C3960 ASIG5V.n5381 VSS 0.056945f
C3961 ASIG5V.n5382 VSS 0.056945f
C3962 ASIG5V.n5383 VSS 0.056945f
C3963 ASIG5V.n5384 VSS 0.056945f
C3964 ASIG5V.n5385 VSS 0.056945f
C3965 ASIG5V.n5386 VSS 0.056945f
C3966 ASIG5V.n5387 VSS 0.056945f
C3967 ASIG5V.n5389 VSS 0.056945f
C3968 ASIG5V.n5390 VSS 0.056945f
C3969 ASIG5V.n5391 VSS 0.056945f
C3970 ASIG5V.n5393 VSS 0.056945f
C3971 ASIG5V.n5394 VSS 0.056945f
C3972 ASIG5V.n5395 VSS 0.056945f
C3973 ASIG5V.n5396 VSS 0.056945f
C3974 ASIG5V.n5397 VSS 0.056945f
C3975 ASIG5V.n5398 VSS 0.056945f
C3976 ASIG5V.n5399 VSS 0.056945f
C3977 ASIG5V.n5401 VSS 0.056945f
C3978 ASIG5V.n5402 VSS 0.056945f
C3979 ASIG5V.n5403 VSS 0.056945f
C3980 ASIG5V.n5405 VSS 0.056945f
C3981 ASIG5V.n5406 VSS 0.056945f
C3982 ASIG5V.n5407 VSS 0.056945f
C3983 ASIG5V.n5408 VSS 0.056945f
C3984 ASIG5V.n5409 VSS 0.056945f
C3985 ASIG5V.n5410 VSS 0.056945f
C3986 ASIG5V.n5411 VSS 0.056945f
C3987 ASIG5V.n5413 VSS 0.056945f
C3988 ASIG5V.n5414 VSS 0.056945f
C3989 ASIG5V.n5415 VSS 0.056945f
C3990 ASIG5V.n5417 VSS 0.056945f
C3991 ASIG5V.n5418 VSS 0.056945f
C3992 ASIG5V.n5419 VSS 0.056945f
C3993 ASIG5V.n5420 VSS 0.056945f
C3994 ASIG5V.n5421 VSS 0.056945f
C3995 ASIG5V.n5422 VSS 0.056945f
C3996 ASIG5V.n5423 VSS 0.056945f
C3997 ASIG5V.n5425 VSS 0.056945f
C3998 ASIG5V.n5426 VSS 0.056945f
C3999 ASIG5V.n5427 VSS 0.056945f
C4000 ASIG5V.n5429 VSS 0.056945f
C4001 ASIG5V.n5430 VSS 0.056945f
C4002 ASIG5V.n5431 VSS 0.056945f
C4003 ASIG5V.n5432 VSS 0.056945f
C4004 ASIG5V.n5433 VSS 0.056945f
C4005 ASIG5V.n5434 VSS 0.056945f
C4006 ASIG5V.n5435 VSS 0.056945f
C4007 ASIG5V.n5437 VSS 0.056945f
C4008 ASIG5V.n5438 VSS 0.056945f
C4009 ASIG5V.n5439 VSS 0.056945f
C4010 ASIG5V.n5441 VSS 0.056945f
C4011 ASIG5V.n5442 VSS 0.056945f
C4012 ASIG5V.n5443 VSS 0.056945f
C4013 ASIG5V.n5444 VSS 0.056945f
C4014 ASIG5V.n5445 VSS 0.056945f
C4015 ASIG5V.n5446 VSS 0.056945f
C4016 ASIG5V.n5447 VSS 0.056945f
C4017 ASIG5V.n5449 VSS 0.056945f
C4018 ASIG5V.n5450 VSS 0.056945f
C4019 ASIG5V.n5451 VSS 0.056945f
C4020 ASIG5V.n5453 VSS 0.056945f
C4021 ASIG5V.n5454 VSS 0.056945f
C4022 ASIG5V.n5455 VSS 0.056945f
C4023 ASIG5V.n5456 VSS 0.056945f
C4024 ASIG5V.n5457 VSS 0.047887f
C4025 ASIG5V.n5458 VSS 0.066995f
C4026 ASIG5V.n5459 VSS 0.054831f
C4027 ASIG5V.n5460 VSS 0.054831f
C4028 ASIG5V.n5461 VSS 0.045974f
C4029 ASIG5V.n5462 VSS 0.076709f
C4030 ASIG5V.n5463 VSS 0.047808f
C4031 ASIG5V.n5464 VSS 0.97853f
C4032 ASIG5V.n5506 VSS 0.269673f
C4033 ASIG5V.n5507 VSS 0.056945f
C4034 ASIG5V.n5508 VSS 0.0621f
C4035 ASIG5V.n5509 VSS 0.036092f
C4036 ASIG5V.n5510 VSS 0.955415f
C4037 ASIG5V.n5511 VSS 0.824431f
C4038 ASIG5V.n5553 VSS 0.924595f
C4039 ASIG5V.n5554 VSS 0.045974f
C4040 ASIG5V.n5555 VSS 0.056945f
C4041 ASIG5V.n5556 VSS 0.056945f
C4042 ASIG5V.n5557 VSS 0.047722f
C4043 ASIG5V.n5558 VSS 0.047808f
C4044 ASIG5V.n5559 VSS 0.076709f
C4045 ASIG5V.n5560 VSS 0.067255f
C4046 ASIG5V.n5561 VSS 0.041754f
C4047 ASIG5V.n5562 VSS 0.052746f
C4048 ASIG5V.n5563 VSS 0.052746f
C4049 ASIG5V.n5564 VSS 0.045974f
C4050 ASIG5V.n5565 VSS 0.076709f
C4051 ASIG5V.n5566 VSS 0.045974f
C4052 ASIG5V.n5567 VSS 0.577872f
C4053 ASIG5V.n5568 VSS 0.716561f
C4054 ASIG5V.n5569 VSS 0.0621f
C4055 ASIG5V.n5570 VSS 0.108961f
C4056 ASIG5V.n5571 VSS 0.0621f
C4057 ASIG5V.n5572 VSS 0.108961f
C4058 ASIG5V.n5573 VSS 0.056945f
C4059 ASIG5V.n5574 VSS 0.056945f
C4060 ASIG5V.n5576 VSS 0.056945f
C4061 ASIG5V.n5577 VSS 0.056945f
C4062 ASIG5V.n5578 VSS 0.056945f
C4063 ASIG5V.n5579 VSS 0.056945f
C4064 ASIG5V.n5582 VSS 0.056945f
C4065 ASIG5V.n5583 VSS 0.056945f
C4066 ASIG5V.n5584 VSS 0.056945f
C4067 ASIG5V.n5585 VSS 0.056945f
C4068 ASIG5V.n5588 VSS 0.056945f
C4069 ASIG5V.n5589 VSS 0.056945f
C4070 ASIG5V.n5590 VSS 0.056945f
C4071 ASIG5V.n5591 VSS 0.056945f
C4072 ASIG5V.n5594 VSS 0.056945f
C4073 ASIG5V.n5595 VSS 0.056945f
C4074 ASIG5V.n5596 VSS 0.056945f
C4075 ASIG5V.n5597 VSS 0.056945f
C4076 ASIG5V.n5600 VSS 0.056945f
C4077 ASIG5V.n5601 VSS 0.056945f
C4078 ASIG5V.n5602 VSS 0.056945f
C4079 ASIG5V.n5603 VSS 0.056945f
C4080 ASIG5V.n5606 VSS 0.056945f
C4081 ASIG5V.n5607 VSS 0.056945f
C4082 ASIG5V.n5608 VSS 0.056945f
C4083 ASIG5V.n5609 VSS 0.056945f
C4084 ASIG5V.n5612 VSS 0.056945f
C4085 ASIG5V.n5613 VSS 0.056945f
C4086 ASIG5V.n5614 VSS 0.056945f
C4087 ASIG5V.n5615 VSS 0.056945f
C4088 ASIG5V.n5618 VSS 0.056945f
C4089 ASIG5V.n5619 VSS 0.056945f
C4090 ASIG5V.n5620 VSS 0.056945f
C4091 ASIG5V.n5621 VSS 0.056945f
C4092 ASIG5V.n5624 VSS 0.056945f
C4093 ASIG5V.n5625 VSS 0.056945f
C4094 ASIG5V.n5626 VSS 0.056945f
C4095 ASIG5V.n5627 VSS 0.056945f
C4096 ASIG5V.n5630 VSS 0.056945f
C4097 ASIG5V.n5631 VSS 0.056945f
C4098 ASIG5V.n5632 VSS 0.056945f
C4099 ASIG5V.n5633 VSS 0.056945f
C4100 ASIG5V.n5636 VSS 0.056945f
C4101 ASIG5V.n5637 VSS 0.056945f
C4102 ASIG5V.n5638 VSS 0.056945f
C4103 ASIG5V.n5639 VSS 0.056945f
C4104 ASIG5V.n5642 VSS 0.056945f
C4105 ASIG5V.n5643 VSS 0.056945f
C4106 ASIG5V.n5644 VSS 0.056945f
C4107 ASIG5V.n5645 VSS 0.056945f
C4108 ASIG5V.n5648 VSS 0.056945f
C4109 ASIG5V.n5649 VSS 0.056945f
C4110 ASIG5V.n5650 VSS 0.056945f
C4111 ASIG5V.n5651 VSS 0.056945f
C4112 ASIG5V.n5654 VSS 0.056945f
C4113 ASIG5V.n5655 VSS 0.056945f
C4114 ASIG5V.n5656 VSS 0.056945f
C4115 ASIG5V.n5657 VSS 0.056945f
C4116 ASIG5V.n5660 VSS 0.056945f
C4117 ASIG5V.n5661 VSS 0.056945f
C4118 ASIG5V.n5662 VSS 0.056945f
C4119 ASIG5V.n5663 VSS 0.056945f
C4120 ASIG5V.n5666 VSS 0.056945f
C4121 ASIG5V.n5667 VSS 0.056945f
C4122 ASIG5V.n5668 VSS 0.056945f
C4123 ASIG5V.n5669 VSS 0.056945f
C4124 ASIG5V.n5672 VSS 0.056945f
C4125 ASIG5V.n5673 VSS 0.056945f
C4126 ASIG5V.n5674 VSS 0.056945f
C4127 ASIG5V.n5675 VSS 0.056945f
C4128 ASIG5V.n5678 VSS 0.056945f
C4129 ASIG5V.n5679 VSS 0.056945f
C4130 ASIG5V.n5680 VSS 0.056945f
C4131 ASIG5V.n5681 VSS 0.056945f
C4132 ASIG5V.n5684 VSS 0.056945f
C4133 ASIG5V.n5685 VSS 0.056945f
C4134 ASIG5V.n5686 VSS 0.056945f
C4135 ASIG5V.n5687 VSS 0.056945f
C4136 ASIG5V.n5690 VSS 0.056945f
C4137 ASIG5V.n5691 VSS 0.056945f
C4138 ASIG5V.n5692 VSS 0.056945f
C4139 ASIG5V.n5693 VSS 0.056945f
C4140 ASIG5V.n5696 VSS 0.036092f
C4141 ASIG5V.n5697 VSS 0.036092f
C4142 ASIG5V.n5698 VSS 0.047722f
C4143 ASIG5V.n5699 VSS 0.056945f
C4144 ASIG5V.n5700 VSS 0.056945f
C4145 ASIG5V.n5701 VSS 0.056945f
C4146 ASIG5V.n5703 VSS 0.056945f
C4147 ASIG5V.n5705 VSS 0.056945f
C4148 ASIG5V.n5706 VSS 0.056945f
C4149 ASIG5V.n5707 VSS 0.056945f
C4150 ASIG5V.n5708 VSS 0.056945f
C4151 ASIG5V.n5709 VSS 0.056945f
C4152 ASIG5V.n5710 VSS 0.056945f
C4153 ASIG5V.n5711 VSS 0.056945f
C4154 ASIG5V.n5713 VSS 0.056945f
C4155 ASIG5V.n5715 VSS 0.056945f
C4156 ASIG5V.n5716 VSS 0.056945f
C4157 ASIG5V.n5717 VSS 0.056945f
C4158 ASIG5V.n5718 VSS 0.056945f
C4159 ASIG5V.n5719 VSS 0.056945f
C4160 ASIG5V.n5720 VSS 0.056945f
C4161 ASIG5V.n5721 VSS 0.056945f
C4162 ASIG5V.n5723 VSS 0.056945f
C4163 ASIG5V.n5725 VSS 0.056945f
C4164 ASIG5V.n5726 VSS 0.056945f
C4165 ASIG5V.n5727 VSS 0.056945f
C4166 ASIG5V.n5728 VSS 0.056945f
C4167 ASIG5V.n5729 VSS 0.056945f
C4168 ASIG5V.n5730 VSS 0.056945f
C4169 ASIG5V.n5731 VSS 0.056945f
C4170 ASIG5V.n5733 VSS 0.056945f
C4171 ASIG5V.n5735 VSS 0.056945f
C4172 ASIG5V.n5736 VSS 0.056945f
C4173 ASIG5V.n5737 VSS 0.056945f
C4174 ASIG5V.n5738 VSS 0.056945f
C4175 ASIG5V.n5739 VSS 0.056945f
C4176 ASIG5V.n5740 VSS 0.056945f
C4177 ASIG5V.n5741 VSS 0.056945f
C4178 ASIG5V.n5743 VSS 0.056945f
C4179 ASIG5V.n5745 VSS 0.056945f
C4180 ASIG5V.n5746 VSS 0.056945f
C4181 ASIG5V.n5747 VSS 0.056945f
C4182 ASIG5V.n5748 VSS 0.056945f
C4183 ASIG5V.n5749 VSS 0.056945f
C4184 ASIG5V.n5750 VSS 0.056945f
C4185 ASIG5V.n5751 VSS 0.056945f
C4186 ASIG5V.n5753 VSS 0.056945f
C4187 ASIG5V.n5755 VSS 0.056945f
C4188 ASIG5V.n5756 VSS 0.056945f
C4189 ASIG5V.n5757 VSS 0.056945f
C4190 ASIG5V.n5758 VSS 0.056945f
C4191 ASIG5V.n5759 VSS 0.056945f
C4192 ASIG5V.n5760 VSS 0.056945f
C4193 ASIG5V.n5761 VSS 0.056945f
C4194 ASIG5V.n5763 VSS 0.056945f
C4195 ASIG5V.n5765 VSS 0.056945f
C4196 ASIG5V.n5766 VSS 0.056945f
C4197 ASIG5V.n5767 VSS 0.056945f
C4198 ASIG5V.n5768 VSS 0.056945f
C4199 ASIG5V.n5769 VSS 0.056945f
C4200 ASIG5V.n5770 VSS 0.056945f
C4201 ASIG5V.n5771 VSS 0.056945f
C4202 ASIG5V.n5773 VSS 0.056945f
C4203 ASIG5V.n5775 VSS 0.056945f
C4204 ASIG5V.n5776 VSS 0.056945f
C4205 ASIG5V.n5777 VSS 0.056945f
C4206 ASIG5V.n5778 VSS 0.056945f
C4207 ASIG5V.n5779 VSS 0.056945f
C4208 ASIG5V.n5780 VSS 0.056945f
C4209 ASIG5V.n5781 VSS 0.056945f
C4210 ASIG5V.n5783 VSS 0.056945f
C4211 ASIG5V.n5785 VSS 0.056945f
C4212 ASIG5V.n5786 VSS 0.056945f
C4213 ASIG5V.n5787 VSS 0.056945f
C4214 ASIG5V.n5788 VSS 0.056945f
C4215 ASIG5V.n5789 VSS 0.056945f
C4216 ASIG5V.n5790 VSS 0.056945f
C4217 ASIG5V.n5791 VSS 0.056945f
C4218 ASIG5V.n5793 VSS 0.056945f
C4219 ASIG5V.n5795 VSS 0.056945f
C4220 ASIG5V.n5796 VSS 0.056945f
C4221 ASIG5V.n5797 VSS 0.056945f
C4222 ASIG5V.n5798 VSS 0.056945f
C4223 ASIG5V.n5799 VSS 0.056945f
C4224 ASIG5V.n5800 VSS 0.056945f
C4225 ASIG5V.n5801 VSS 0.056945f
C4226 ASIG5V.n5803 VSS 0.056945f
C4227 ASIG5V.n5805 VSS 0.056945f
C4228 ASIG5V.n5806 VSS 0.056945f
C4229 ASIG5V.n5807 VSS 0.056945f
C4230 ASIG5V.n5808 VSS 0.056945f
C4231 ASIG5V.n5809 VSS 0.056945f
C4232 ASIG5V.n5810 VSS 0.056945f
C4233 ASIG5V.n5811 VSS 0.056945f
C4234 ASIG5V.n5813 VSS 0.056945f
C4235 ASIG5V.n5815 VSS 0.056945f
C4236 ASIG5V.n5816 VSS 0.056945f
C4237 ASIG5V.n5817 VSS 0.056945f
C4238 ASIG5V.n5818 VSS 0.056945f
C4239 ASIG5V.n5819 VSS 0.056945f
C4240 ASIG5V.n5820 VSS 0.056945f
C4241 ASIG5V.n5821 VSS 0.056945f
C4242 ASIG5V.n5823 VSS 0.056945f
C4243 ASIG5V.n5825 VSS 0.056945f
C4244 ASIG5V.n5826 VSS 0.056945f
C4245 ASIG5V.n5827 VSS 0.056945f
C4246 ASIG5V.n5828 VSS 0.056945f
C4247 ASIG5V.n5829 VSS 0.056945f
C4248 ASIG5V.n5830 VSS 0.056945f
C4249 ASIG5V.n5831 VSS 0.056945f
C4250 ASIG5V.n5833 VSS 0.056945f
C4251 ASIG5V.n5835 VSS 0.056945f
C4252 ASIG5V.n5836 VSS 0.056945f
C4253 ASIG5V.n5837 VSS 0.056945f
C4254 ASIG5V.n5838 VSS 0.056945f
C4255 ASIG5V.n5839 VSS 0.056945f
C4256 ASIG5V.n5840 VSS 0.056945f
C4257 ASIG5V.n5841 VSS 0.056945f
C4258 ASIG5V.n5843 VSS 0.056945f
C4259 ASIG5V.n5845 VSS 0.056945f
C4260 ASIG5V.n5846 VSS 0.056945f
C4261 ASIG5V.n5847 VSS 0.056945f
C4262 ASIG5V.n5848 VSS 0.056945f
C4263 ASIG5V.n5849 VSS 0.056945f
C4264 ASIG5V.n5850 VSS 0.056945f
C4265 ASIG5V.n5851 VSS 0.056945f
C4266 ASIG5V.n5853 VSS 0.056945f
C4267 ASIG5V.n5855 VSS 0.056945f
C4268 ASIG5V.n5856 VSS 0.056945f
C4269 ASIG5V.n5857 VSS 0.056945f
C4270 ASIG5V.n5858 VSS 0.056945f
C4271 ASIG5V.n5859 VSS 0.056945f
C4272 ASIG5V.n5860 VSS 0.056945f
C4273 ASIG5V.n5861 VSS 0.056945f
C4274 ASIG5V.n5863 VSS 0.056945f
C4275 ASIG5V.n5865 VSS 0.056945f
C4276 ASIG5V.n5866 VSS 0.056945f
C4277 ASIG5V.n5867 VSS 0.056945f
C4278 ASIG5V.n5868 VSS 0.056945f
C4279 ASIG5V.n5869 VSS 0.056945f
C4280 ASIG5V.n5870 VSS 0.056945f
C4281 ASIG5V.n5871 VSS 0.056945f
C4282 ASIG5V.n5873 VSS 0.056945f
C4283 ASIG5V.n5875 VSS 0.056945f
C4284 ASIG5V.n5876 VSS 0.056945f
C4285 ASIG5V.n5877 VSS 0.056945f
C4286 ASIG5V.n5878 VSS 0.056945f
C4287 ASIG5V.n5879 VSS 0.056945f
C4288 ASIG5V.n5880 VSS 0.056945f
C4289 ASIG5V.n5881 VSS 0.056945f
C4290 ASIG5V.n5883 VSS 0.056945f
C4291 ASIG5V.n5885 VSS 0.056945f
C4292 ASIG5V.n5886 VSS 0.056945f
C4293 ASIG5V.n5887 VSS 0.056945f
C4294 ASIG5V.n5888 VSS 0.056945f
C4295 ASIG5V.n5889 VSS 0.056945f
C4296 ASIG5V.n5890 VSS 0.056945f
C4297 ASIG5V.n5891 VSS 0.056945f
C4298 ASIG5V.n5893 VSS 0.056945f
C4299 ASIG5V.n5895 VSS 0.056945f
C4300 ASIG5V.n5896 VSS 0.056945f
C4301 ASIG5V.n5897 VSS 0.056945f
C4302 ASIG5V.n5898 VSS 0.056945f
C4303 ASIG5V.n5899 VSS 0.056945f
C4304 ASIG5V.n5900 VSS 0.056945f
C4305 ASIG5V.n5901 VSS 0.056945f
C4306 ASIG5V.n5903 VSS 0.056945f
C4307 ASIG5V.n5905 VSS 0.036092f
C4308 ASIG5V.n5906 VSS 0.036092f
C4309 ASIG5V.n5907 VSS 0.052133f
C4310 ASIG5V.n5908 VSS 0.07229f
C4311 ASIG5V.n5909 VSS 0.07229f
C4312 ASIG5V.n5910 VSS 0.0621f
C4313 ASIG5V.n5911 VSS 0.0621f
C4314 ASIG5V.n5912 VSS 0.955415f
C4315 ASIG5V.n5954 VSS 0.662626f
C4316 ASIG5V.n5955 VSS 0.056945f
C4317 ASIG5V.n5956 VSS 0.036092f
C4318 ASIG5V.n5957 VSS 0.470002f
C4319 ASIG5V.n5999 VSS 0.662626f
C4320 ASIG5V.n6000 VSS 0.045974f
C4321 ASIG5V.n6001 VSS 0.056945f
C4322 ASIG5V.n6002 VSS 0.056945f
C4323 ASIG5V.n6003 VSS 0.056945f
C4324 ASIG5V.n6004 VSS 0.056945f
C4325 ASIG5V.n6005 VSS 0.056945f
C4326 ASIG5V.n6006 VSS 0.056945f
C4327 ASIG5V.n6007 VSS 0.056945f
C4328 ASIG5V.n6008 VSS 0.056945f
C4329 ASIG5V.n6009 VSS 0.056945f
C4330 ASIG5V.n6010 VSS 0.056945f
C4331 ASIG5V.n6011 VSS 0.056945f
C4332 ASIG5V.n6012 VSS 0.056945f
C4333 ASIG5V.n6013 VSS 0.056945f
C4334 ASIG5V.n6014 VSS 0.056945f
C4335 ASIG5V.n6015 VSS 0.056945f
C4336 ASIG5V.n6016 VSS 0.056945f
C4337 ASIG5V.n6017 VSS 0.056945f
C4338 ASIG5V.n6018 VSS 0.056945f
C4339 ASIG5V.n6019 VSS 0.056945f
C4340 ASIG5V.n6020 VSS 0.056945f
C4341 ASIG5V.n6021 VSS 0.056945f
C4342 ASIG5V.n6022 VSS 0.056945f
C4343 ASIG5V.n6023 VSS 0.056945f
C4344 ASIG5V.n6024 VSS 0.056945f
C4345 ASIG5V.n6025 VSS 0.056945f
C4346 ASIG5V.n6026 VSS 0.056945f
C4347 ASIG5V.n6027 VSS 0.056945f
C4348 ASIG5V.n6028 VSS 0.056945f
C4349 ASIG5V.n6029 VSS 0.056945f
C4350 ASIG5V.n6030 VSS 0.056945f
C4351 ASIG5V.n6031 VSS 0.056945f
C4352 ASIG5V.n6032 VSS 0.056945f
C4353 ASIG5V.n6033 VSS 0.056945f
C4354 ASIG5V.n6034 VSS 0.056945f
C4355 ASIG5V.n6035 VSS 0.056945f
C4356 ASIG5V.n6036 VSS 0.056945f
C4357 ASIG5V.n6037 VSS 0.056945f
C4358 ASIG5V.n6038 VSS 0.056945f
C4359 ASIG5V.n6039 VSS 0.056945f
C4360 ASIG5V.n6040 VSS 0.056945f
C4361 ASIG5V.n6041 VSS 0.056945f
C4362 ASIG5V.n6042 VSS 0.056945f
C4363 ASIG5V.n6043 VSS 0.056945f
C4364 ASIG5V.n6044 VSS 0.056945f
C4365 ASIG5V.n6045 VSS 0.056945f
C4366 ASIG5V.n6046 VSS 0.056945f
C4367 ASIG5V.n6047 VSS 0.056945f
C4368 ASIG5V.n6048 VSS 0.056945f
C4369 ASIG5V.n6049 VSS 0.056945f
C4370 ASIG5V.n6050 VSS 0.056945f
C4371 ASIG5V.n6051 VSS 0.056945f
C4372 ASIG5V.n6052 VSS 0.056945f
C4373 ASIG5V.n6053 VSS 0.056945f
C4374 ASIG5V.n6054 VSS 0.056945f
C4375 ASIG5V.n6055 VSS 0.056945f
C4376 ASIG5V.n6056 VSS 0.056945f
C4377 ASIG5V.n6057 VSS 0.056945f
C4378 ASIG5V.n6058 VSS 0.056945f
C4379 ASIG5V.n6059 VSS 0.056945f
C4380 ASIG5V.n6060 VSS 0.056945f
C4381 ASIG5V.n6061 VSS 0.056945f
C4382 ASIG5V.n6062 VSS 0.056945f
C4383 ASIG5V.n6063 VSS 0.052133f
C4384 ASIG5V.n6064 VSS 0.056945f
C4385 ASIG5V.n6065 VSS 0.056945f
C4386 ASIG5V.n6066 VSS 0.056945f
C4387 ASIG5V.n6067 VSS 0.056945f
C4388 ASIG5V.n6068 VSS 0.056945f
C4389 ASIG5V.n6069 VSS 0.056945f
C4390 ASIG5V.n6070 VSS 0.056945f
C4391 ASIG5V.n6071 VSS 0.056945f
C4392 ASIG5V.n6072 VSS 0.056945f
C4393 ASIG5V.n6073 VSS 0.056945f
C4394 ASIG5V.n6074 VSS 0.056945f
C4395 ASIG5V.n6075 VSS 0.056945f
C4396 ASIG5V.n6076 VSS 0.056945f
C4397 ASIG5V.n6077 VSS 0.056945f
C4398 ASIG5V.n6078 VSS 0.056945f
C4399 ASIG5V.n6079 VSS 0.056945f
C4400 ASIG5V.n6080 VSS 0.056945f
C4401 ASIG5V.n6081 VSS 0.056945f
C4402 ASIG5V.n6082 VSS 0.056945f
C4403 ASIG5V.n6083 VSS 0.056945f
C4404 ASIG5V.n6084 VSS 0.056945f
C4405 ASIG5V.n6085 VSS 0.056945f
C4406 ASIG5V.n6086 VSS 0.056945f
C4407 ASIG5V.n6087 VSS 0.056945f
C4408 ASIG5V.n6088 VSS 0.056945f
C4409 ASIG5V.n6089 VSS 0.056945f
C4410 ASIG5V.n6090 VSS 0.056945f
C4411 ASIG5V.n6091 VSS 0.056945f
C4412 ASIG5V.n6092 VSS 0.056945f
C4413 ASIG5V.n6093 VSS 0.056945f
C4414 ASIG5V.n6094 VSS 0.056945f
C4415 ASIG5V.n6095 VSS 0.056945f
C4416 ASIG5V.n6096 VSS 0.056945f
C4417 ASIG5V.n6097 VSS 0.056945f
C4418 ASIG5V.n6098 VSS 0.056945f
C4419 ASIG5V.n6099 VSS 0.056945f
C4420 ASIG5V.n6100 VSS 0.056945f
C4421 ASIG5V.n6101 VSS 0.056945f
C4422 ASIG5V.n6102 VSS 0.056945f
C4423 ASIG5V.n6103 VSS 0.056945f
C4424 ASIG5V.n6104 VSS 0.056945f
C4425 ASIG5V.n6105 VSS 0.056945f
C4426 ASIG5V.n6106 VSS 0.056945f
C4427 ASIG5V.n6107 VSS 0.056945f
C4428 ASIG5V.n6108 VSS 0.056945f
C4429 ASIG5V.n6109 VSS 0.056945f
C4430 ASIG5V.n6110 VSS 0.056945f
C4431 ASIG5V.n6111 VSS 0.056945f
C4432 ASIG5V.n6112 VSS 0.056945f
C4433 ASIG5V.n6113 VSS 0.056945f
C4434 ASIG5V.n6114 VSS 0.056945f
C4435 ASIG5V.n6115 VSS 0.056945f
C4436 ASIG5V.n6116 VSS 0.056945f
C4437 ASIG5V.n6117 VSS 0.056945f
C4438 ASIG5V.n6118 VSS 0.056945f
C4439 ASIG5V.n6119 VSS 0.056945f
C4440 ASIG5V.n6120 VSS 0.056945f
C4441 ASIG5V.n6121 VSS 0.056945f
C4442 ASIG5V.n6122 VSS 0.056945f
C4443 ASIG5V.n6123 VSS 0.056945f
C4444 ASIG5V.n6124 VSS 0.056945f
C4445 ASIG5V.n6125 VSS 0.056945f
C4446 ASIG5V.n6126 VSS 0.056945f
C4447 ASIG5V.n6127 VSS 0.056945f
C4448 ASIG5V.n6128 VSS 0.056945f
C4449 ASIG5V.n6129 VSS 0.056945f
C4450 ASIG5V.n6130 VSS 0.056945f
C4451 ASIG5V.n6131 VSS 0.056945f
C4452 ASIG5V.n6132 VSS 0.056945f
C4453 ASIG5V.n6133 VSS 0.056945f
C4454 ASIG5V.n6134 VSS 0.056945f
C4455 ASIG5V.n6135 VSS 0.056945f
C4456 ASIG5V.n6136 VSS 0.056945f
C4457 ASIG5V.n6137 VSS 0.056945f
C4458 ASIG5V.n6138 VSS 0.056945f
C4459 ASIG5V.n6139 VSS 0.056945f
C4460 ASIG5V.n6140 VSS 0.056945f
C4461 ASIG5V.n6141 VSS 0.056945f
C4462 ASIG5V.n6142 VSS 0.056945f
C4463 ASIG5V.n6143 VSS 0.056945f
C4464 ASIG5V.n6144 VSS 0.056945f
C4465 ASIG5V.n6145 VSS 0.056945f
C4466 ASIG5V.n6146 VSS 0.056945f
C4467 ASIG5V.n6147 VSS 0.056945f
C4468 ASIG5V.n6148 VSS 0.056945f
C4469 ASIG5V.n6149 VSS 0.056945f
C4470 ASIG5V.n6150 VSS 0.056945f
C4471 ASIG5V.n6151 VSS 0.056945f
C4472 ASIG5V.n6152 VSS 0.056945f
C4473 ASIG5V.n6153 VSS 0.056945f
C4474 ASIG5V.n6154 VSS 0.056945f
C4475 ASIG5V.n6155 VSS 0.056945f
C4476 ASIG5V.n6156 VSS 0.056945f
C4477 ASIG5V.n6157 VSS 0.056945f
C4478 ASIG5V.n6158 VSS 0.056945f
C4479 ASIG5V.n6159 VSS 0.056945f
C4480 ASIG5V.n6160 VSS 0.056945f
C4481 ASIG5V.n6161 VSS 0.056945f
C4482 ASIG5V.n6162 VSS 0.056945f
C4483 ASIG5V.n6163 VSS 0.056945f
C4484 ASIG5V.n6164 VSS 0.056945f
C4485 ASIG5V.n6165 VSS 0.056945f
C4486 ASIG5V.n6166 VSS 0.056945f
C4487 ASIG5V.n6167 VSS 0.056945f
C4488 ASIG5V.n6168 VSS 0.056945f
C4489 ASIG5V.n6169 VSS 0.056945f
C4490 ASIG5V.n6170 VSS 0.056945f
C4491 ASIG5V.n6171 VSS 0.056945f
C4492 ASIG5V.n6172 VSS 0.056945f
C4493 ASIG5V.n6173 VSS 0.056945f
C4494 ASIG5V.n6174 VSS 0.056945f
C4495 ASIG5V.n6175 VSS 0.056945f
C4496 ASIG5V.n6176 VSS 0.056945f
C4497 ASIG5V.n6177 VSS 0.056945f
C4498 ASIG5V.n6178 VSS 0.056945f
C4499 ASIG5V.n6179 VSS 0.056945f
C4500 ASIG5V.n6180 VSS 0.056945f
C4501 ASIG5V.n6181 VSS 0.056945f
C4502 ASIG5V.n6182 VSS 0.056945f
C4503 ASIG5V.n6183 VSS 0.056945f
C4504 ASIG5V.n6184 VSS 0.056945f
C4505 ASIG5V.n6185 VSS 0.056945f
C4506 ASIG5V.n6186 VSS 0.056945f
C4507 ASIG5V.n6187 VSS 0.056945f
C4508 ASIG5V.n6188 VSS 0.056945f
C4509 ASIG5V.n6189 VSS 0.056945f
C4510 ASIG5V.n6190 VSS 0.056945f
C4511 ASIG5V.n6191 VSS 0.056945f
C4512 ASIG5V.n6192 VSS 0.056945f
C4513 ASIG5V.n6193 VSS 0.056945f
C4514 ASIG5V.n6194 VSS 0.056945f
C4515 ASIG5V.n6195 VSS 0.056945f
C4516 ASIG5V.n6196 VSS 0.056945f
C4517 ASIG5V.n6197 VSS 0.056945f
C4518 ASIG5V.n6198 VSS 0.056945f
C4519 ASIG5V.n6199 VSS 0.056945f
C4520 ASIG5V.n6200 VSS 0.056945f
C4521 ASIG5V.n6201 VSS 0.056945f
C4522 ASIG5V.n6202 VSS 0.056945f
C4523 ASIG5V.n6203 VSS 0.056945f
C4524 ASIG5V.n6204 VSS 0.056945f
C4525 ASIG5V.n6205 VSS 0.056945f
C4526 ASIG5V.n6206 VSS 0.056945f
C4527 ASIG5V.n6207 VSS 0.056945f
C4528 ASIG5V.n6208 VSS 0.056945f
C4529 ASIG5V.n6209 VSS 0.056945f
C4530 ASIG5V.n6210 VSS 0.056945f
C4531 ASIG5V.n6211 VSS 0.056945f
C4532 ASIG5V.n6212 VSS 0.056945f
C4533 ASIG5V.n6213 VSS 0.056945f
C4534 ASIG5V.n6214 VSS 0.056945f
C4535 ASIG5V.n6215 VSS 0.056945f
C4536 ASIG5V.n6216 VSS 0.056945f
C4537 ASIG5V.n6217 VSS 0.056945f
C4538 ASIG5V.n6218 VSS 0.056945f
C4539 ASIG5V.n6219 VSS 0.056945f
C4540 ASIG5V.n6220 VSS 0.056945f
C4541 ASIG5V.n6221 VSS 0.056945f
C4542 ASIG5V.n6222 VSS 0.056945f
C4543 ASIG5V.n6223 VSS 0.056945f
C4544 ASIG5V.n6224 VSS 0.056945f
C4545 ASIG5V.n6225 VSS 0.056945f
C4546 ASIG5V.n6226 VSS 0.056945f
C4547 ASIG5V.n6227 VSS 0.056945f
C4548 ASIG5V.n6228 VSS 0.056945f
C4549 ASIG5V.n6229 VSS 0.056945f
C4550 ASIG5V.n6230 VSS 0.056945f
C4551 ASIG5V.n6231 VSS 0.056945f
C4552 ASIG5V.n6232 VSS 0.056945f
C4553 ASIG5V.n6233 VSS 0.056945f
C4554 ASIG5V.n6234 VSS 0.056945f
C4555 ASIG5V.n6235 VSS 0.056945f
C4556 ASIG5V.n6236 VSS 0.056945f
C4557 ASIG5V.n6237 VSS 0.056945f
C4558 ASIG5V.n6238 VSS 0.056945f
C4559 ASIG5V.n6239 VSS 0.056945f
C4560 ASIG5V.n6240 VSS 0.056945f
C4561 ASIG5V.n6241 VSS 0.056945f
C4562 ASIG5V.n6242 VSS 0.056945f
C4563 ASIG5V.n6243 VSS 0.056945f
C4564 ASIG5V.n6244 VSS 0.056945f
C4565 ASIG5V.n6245 VSS 0.056945f
C4566 ASIG5V.n6246 VSS 0.056945f
C4567 ASIG5V.n6247 VSS 0.047722f
C4568 ASIG5V.n6248 VSS 0.072117f
C4569 ASIG5V.n6249 VSS 0.076709f
C4570 ASIG5V.n6250 VSS 0.042946f
C4571 ASIG5V.n6251 VSS 0.072117f
C4572 ASIG5V.n6252 VSS 1.0941f
C4573 ASIG5V.n6253 VSS 0.678036f
C4574 ASIG5V.n6254 VSS 0.074278f
C4575 ASIG5V.n6255 VSS 0.074278f
C4576 ASIG5V.n6256 VSS 0.064871f
C4577 ASIG5V.n6257 VSS 0.062984f
C4578 ASIG5V.n6258 VSS 0.052746f
C4579 ASIG5V.n6259 VSS 0.052746f
C4580 ASIG5V.n6260 VSS 0.045974f
C4581 ASIG5V.n6261 VSS 0.076709f
C4582 ASIG5V.n6262 VSS 0.045974f
C4583 ASIG5V.n6263 VSS 0.955415f
C4584 ASIG5V.n6264 VSS 1.0941f
C4585 ASIG5V.n6306 VSS 0.886071f
C4586 ASIG5V.n6307 VSS 0.056945f
C4587 ASIG5V.n6308 VSS 0.0621f
C4588 ASIG5V.n6309 VSS 0.036092f
C4589 ASIG5V.n6310 VSS 0.662626f
C4590 ASIG5V.n6352 VSS 0.886071f
C4591 ASIG5V.n6353 VSS 0.056945f
C4592 ASIG5V.n6354 VSS 0.056945f
C4593 ASIG5V.n6355 VSS 0.056945f
C4594 ASIG5V.n6356 VSS 0.056945f
C4595 ASIG5V.n6357 VSS 0.056945f
C4596 ASIG5V.n6358 VSS 0.056945f
C4597 ASIG5V.n6359 VSS 0.056945f
C4598 ASIG5V.n6360 VSS 0.056945f
C4599 ASIG5V.n6361 VSS 0.056945f
C4600 ASIG5V.n6362 VSS 0.056945f
C4601 ASIG5V.n6363 VSS 0.056945f
C4602 ASIG5V.n6364 VSS 0.056945f
C4603 ASIG5V.n6365 VSS 0.056945f
C4604 ASIG5V.n6366 VSS 0.056945f
C4605 ASIG5V.n6367 VSS 0.056945f
C4606 ASIG5V.n6368 VSS 0.056945f
C4607 ASIG5V.n6369 VSS 0.056945f
C4608 ASIG5V.n6370 VSS 0.056945f
C4609 ASIG5V.n6371 VSS 0.056945f
C4610 ASIG5V.n6372 VSS 0.056945f
C4611 ASIG5V.n6373 VSS 0.056945f
C4612 ASIG5V.n6374 VSS 0.056945f
C4613 ASIG5V.n6375 VSS 0.056945f
C4614 ASIG5V.n6376 VSS 0.056945f
C4615 ASIG5V.n6377 VSS 0.056945f
C4616 ASIG5V.n6378 VSS 0.056945f
C4617 ASIG5V.n6379 VSS 0.056945f
C4618 ASIG5V.n6380 VSS 0.056945f
C4619 ASIG5V.n6381 VSS 0.056945f
C4620 ASIG5V.n6382 VSS 0.056945f
C4621 ASIG5V.n6383 VSS 0.056945f
C4622 ASIG5V.n6384 VSS 0.056945f
C4623 ASIG5V.n6385 VSS 0.056945f
C4624 ASIG5V.n6386 VSS 0.056945f
C4625 ASIG5V.n6387 VSS 0.056945f
C4626 ASIG5V.n6388 VSS 0.056945f
C4627 ASIG5V.n6389 VSS 0.056945f
C4628 ASIG5V.n6390 VSS 0.056945f
C4629 ASIG5V.n6391 VSS 0.056945f
C4630 ASIG5V.n6392 VSS 0.056945f
C4631 ASIG5V.n6393 VSS 0.056945f
C4632 ASIG5V.n6394 VSS 0.056945f
C4633 ASIG5V.n6395 VSS 0.056945f
C4634 ASIG5V.n6396 VSS 0.056945f
C4635 ASIG5V.n6397 VSS 0.056945f
C4636 ASIG5V.n6398 VSS 0.056945f
C4637 ASIG5V.n6399 VSS 0.056945f
C4638 ASIG5V.n6400 VSS 0.056945f
C4639 ASIG5V.n6401 VSS 0.056945f
C4640 ASIG5V.n6402 VSS 0.056945f
C4641 ASIG5V.n6403 VSS 0.056945f
C4642 ASIG5V.n6404 VSS 0.056945f
C4643 ASIG5V.n6405 VSS 0.056945f
C4644 ASIG5V.n6406 VSS 0.056945f
C4645 ASIG5V.n6407 VSS 0.056945f
C4646 ASIG5V.n6408 VSS 0.056945f
C4647 ASIG5V.n6409 VSS 0.056945f
C4648 ASIG5V.n6410 VSS 0.056945f
C4649 ASIG5V.n6411 VSS 0.056945f
C4650 ASIG5V.n6412 VSS 0.056945f
C4651 ASIG5V.n6413 VSS 0.056945f
C4652 ASIG5V.n6414 VSS 0.056945f
C4653 ASIG5V.n6415 VSS 0.054905f
C4654 ASIG5V.n6416 VSS 0.548344f
C4655 ASIG5V.n6417 VSS 0.108961f
C4656 ASIG5V.n6418 VSS 0.059753f
C4657 ASIG5V.n6419 VSS 0.059753f
C4658 ASIG5V.n6420 VSS 0.053336f
C4659 ASIG5V.n6421 VSS 0.09726f
C4660 ASIG5V.n6422 VSS 0.09726f
C4661 ASIG5V.n6423 VSS 0.108961f
C4662 ASIG5V.n6424 VSS 0.108961f
C4663 ASIG5V.n6425 VSS 0.108961f
C4664 ASIG5V.n6426 VSS 0.06151f
C4665 ASIG5V.n6427 VSS 0.06151f
C4666 ASIG5V.n6428 VSS 0.0621f
C4667 ASIG5V.n6429 VSS 0.108961f
C4668 ASIG5V.n6430 VSS 0.073812f
C4669 ASIG5V.n6431 VSS 0.955415f
C4670 ASIG5V.n6432 VSS 0.223443f
C4671 ASIG5V.n6433 VSS 0.076709f
C4672 ASIG5V.n6434 VSS 0.045974f
C4673 ASIG5V.n6435 VSS 0.076709f
C4674 ASIG5V.n6436 VSS 0.045974f
C4675 ASIG5V.n6437 VSS 0.049969f
C4676 ASIG5V.n6438 VSS 0.049969f
C4677 ASIG5V.n6439 VSS 0.043641f
C4678 ASIG5V.n6440 VSS 0.066995f
C4679 ASIG5V.n6441 VSS 0.047722f
C4680 ASIG5V.n6442 VSS 0.066995f
C4681 ASIG5V.n6443 VSS 0.076709f
C4682 ASIG5V.n6444 VSS 0.076709f
C4683 ASIG5V.n6445 VSS 1.0864f
C4684 ASIG5V.n6487 VSS 0.036092f
C4685 ASIG5V.n6488 VSS 1.03247f
C4686 ASIG5V.n6489 VSS 0.036092f
C4687 ASIG5V.n6490 VSS 0.056945f
C4688 ASIG5V.n6491 VSS 0.056945f
C4689 ASIG5V.n6492 VSS 0.056945f
C4690 ASIG5V.n6493 VSS 0.056945f
C4691 ASIG5V.n6494 VSS 0.056945f
C4692 ASIG5V.n6495 VSS 0.056945f
C4693 ASIG5V.n6496 VSS 0.056945f
C4694 ASIG5V.n6497 VSS 0.056945f
C4695 ASIG5V.n6498 VSS 0.056945f
C4696 ASIG5V.n6499 VSS 0.056945f
C4697 ASIG5V.n6500 VSS 0.056945f
C4698 ASIG5V.n6501 VSS 0.056945f
C4699 ASIG5V.n6502 VSS 0.056945f
C4700 ASIG5V.n6503 VSS 0.056945f
C4701 ASIG5V.n6504 VSS 0.056945f
C4702 ASIG5V.n6505 VSS 0.056945f
C4703 ASIG5V.n6506 VSS 0.056945f
C4704 ASIG5V.n6507 VSS 0.056945f
C4705 ASIG5V.n6508 VSS 0.056945f
C4706 ASIG5V.n6509 VSS 0.056945f
C4707 ASIG5V.n6510 VSS 0.056945f
C4708 ASIG5V.n6511 VSS 0.056945f
C4709 ASIG5V.n6512 VSS 0.056945f
C4710 ASIG5V.n6513 VSS 0.056945f
C4711 ASIG5V.n6514 VSS 0.056945f
C4712 ASIG5V.n6515 VSS 0.056945f
C4713 ASIG5V.n6516 VSS 0.056945f
C4714 ASIG5V.n6517 VSS 0.056945f
C4715 ASIG5V.n6518 VSS 0.056945f
C4716 ASIG5V.n6519 VSS 0.056945f
C4717 ASIG5V.n6520 VSS 0.056945f
C4718 ASIG5V.n6521 VSS 0.056945f
C4719 ASIG5V.n6522 VSS 0.056945f
C4720 ASIG5V.n6523 VSS 0.056945f
C4721 ASIG5V.n6524 VSS 0.056945f
C4722 ASIG5V.n6525 VSS 0.056945f
C4723 ASIG5V.n6526 VSS 0.056945f
C4724 ASIG5V.n6527 VSS 0.056945f
C4725 ASIG5V.n6528 VSS 0.056945f
C4726 ASIG5V.n6529 VSS 0.056945f
C4727 ASIG5V.n6531 VSS 0.056945f
C4728 ASIG5V.n6532 VSS 0.056945f
C4729 ASIG5V.n6533 VSS 0.07229f
C4730 ASIG5V.n6534 VSS 0.087848f
C4731 ASIG5V.n6535 VSS 0.065886f
C4732 ASIG5V.n6536 VSS 0.073812f
C4733 ASIG5V.n6537 VSS 0.108961f
C4734 ASIG5V.n6538 VSS 0.0621f
C4735 ASIG5V.n6539 VSS 0.089629f
C4736 ASIG5V.n6540 VSS 0.07229f
C4737 ASIG5V.n6541 VSS 0.0621f
C4738 ASIG5V.n6542 VSS 0.108961f
C4739 ASIG5V.n6543 VSS 0.0621f
C4740 ASIG5V.n6544 VSS 1.00935f
C4741 ASIG5V.n6545 VSS 0.955415f
C4742 ASIG5V.n6587 VSS 0.947711f
C4743 ASIG5V.n6588 VSS 0.056945f
C4744 ASIG5V.n6589 VSS 0.036092f
C4745 ASIG5V.n6590 VSS 0.909185f
C4746 ASIG5V.n6632 VSS 0.809021f
C4747 ASIG5V.n6633 VSS 0.045974f
C4748 ASIG5V.n6634 VSS 0.056945f
C4749 ASIG5V.n6635 VSS 0.056945f
C4750 ASIG5V.n6636 VSS 0.056945f
C4751 ASIG5V.n6637 VSS 0.056945f
C4752 ASIG5V.n6638 VSS 0.056945f
C4753 ASIG5V.n6639 VSS 0.056945f
C4754 ASIG5V.n6640 VSS 0.056945f
C4755 ASIG5V.n6641 VSS 0.056945f
C4756 ASIG5V.n6642 VSS 0.056945f
C4757 ASIG5V.n6643 VSS 0.056945f
C4758 ASIG5V.n6644 VSS 0.056945f
C4759 ASIG5V.n6645 VSS 0.056945f
C4760 ASIG5V.n6646 VSS 0.056945f
C4761 ASIG5V.n6647 VSS 0.056945f
C4762 ASIG5V.n6648 VSS 0.056945f
C4763 ASIG5V.n6649 VSS 0.056945f
C4764 ASIG5V.n6650 VSS 0.056945f
C4765 ASIG5V.n6651 VSS 0.056945f
C4766 ASIG5V.n6652 VSS 0.056945f
C4767 ASIG5V.n6653 VSS 0.056945f
C4768 ASIG5V.n6654 VSS 0.056945f
C4769 ASIG5V.n6655 VSS 0.056945f
C4770 ASIG5V.n6656 VSS 0.056945f
C4771 ASIG5V.n6657 VSS 0.056945f
C4772 ASIG5V.n6658 VSS 0.056945f
C4773 ASIG5V.n6659 VSS 0.056945f
C4774 ASIG5V.n6660 VSS 0.056945f
C4775 ASIG5V.n6661 VSS 0.056945f
C4776 ASIG5V.n6662 VSS 0.056945f
C4777 ASIG5V.n6663 VSS 0.056945f
C4778 ASIG5V.n6664 VSS 0.056945f
C4779 ASIG5V.n6665 VSS 0.056945f
C4780 ASIG5V.n6666 VSS 0.056945f
C4781 ASIG5V.n6667 VSS 0.056945f
C4782 ASIG5V.n6668 VSS 0.056945f
C4783 ASIG5V.n6669 VSS 0.056945f
C4784 ASIG5V.n6670 VSS 0.056945f
C4785 ASIG5V.n6671 VSS 0.056945f
C4786 ASIG5V.n6672 VSS 0.056945f
C4787 ASIG5V.n6673 VSS 0.056945f
C4788 ASIG5V.n6674 VSS 0.056945f
C4789 ASIG5V.n6675 VSS 0.056945f
C4790 ASIG5V.n6676 VSS 0.056945f
C4791 ASIG5V.n6677 VSS 0.056945f
C4792 ASIG5V.n6678 VSS 0.056945f
C4793 ASIG5V.n6679 VSS 0.056945f
C4794 ASIG5V.n6680 VSS 0.056945f
C4795 ASIG5V.n6681 VSS 0.056945f
C4796 ASIG5V.n6682 VSS 0.056945f
C4797 ASIG5V.n6683 VSS 0.056945f
C4798 ASIG5V.n6684 VSS 0.056945f
C4799 ASIG5V.n6685 VSS 0.056945f
C4800 ASIG5V.n6686 VSS 0.056945f
C4801 ASIG5V.n6687 VSS 0.056945f
C4802 ASIG5V.n6688 VSS 0.056945f
C4803 ASIG5V.n6689 VSS 0.056945f
C4804 ASIG5V.n6690 VSS 0.056945f
C4805 ASIG5V.n6691 VSS 0.056945f
C4806 ASIG5V.n6692 VSS 0.056945f
C4807 ASIG5V.n6693 VSS 0.056945f
C4808 ASIG5V.n6694 VSS 0.056945f
C4809 ASIG5V.n6695 VSS 0.056945f
C4810 ASIG5V.n6696 VSS 0.052133f
C4811 ASIG5V.n6697 VSS 0.056945f
C4812 ASIG5V.n6698 VSS 0.056945f
C4813 ASIG5V.n6699 VSS 0.056945f
C4814 ASIG5V.n6700 VSS 0.056945f
C4815 ASIG5V.n6701 VSS 0.056945f
C4816 ASIG5V.n6702 VSS 0.056945f
C4817 ASIG5V.n6703 VSS 0.056945f
C4818 ASIG5V.n6704 VSS 0.056945f
C4819 ASIG5V.n6705 VSS 0.056945f
C4820 ASIG5V.n6706 VSS 0.056945f
C4821 ASIG5V.n6707 VSS 0.056945f
C4822 ASIG5V.n6708 VSS 0.056945f
C4823 ASIG5V.n6709 VSS 0.056945f
C4824 ASIG5V.n6710 VSS 0.056945f
C4825 ASIG5V.n6711 VSS 0.056945f
C4826 ASIG5V.n6712 VSS 0.056945f
C4827 ASIG5V.n6713 VSS 0.056945f
C4828 ASIG5V.n6714 VSS 0.056945f
C4829 ASIG5V.n6715 VSS 0.056945f
C4830 ASIG5V.n6716 VSS 0.056945f
C4831 ASIG5V.n6717 VSS 0.056945f
C4832 ASIG5V.n6718 VSS 0.056945f
C4833 ASIG5V.n6719 VSS 0.056945f
C4834 ASIG5V.n6720 VSS 0.056945f
C4835 ASIG5V.n6721 VSS 0.056945f
C4836 ASIG5V.n6722 VSS 0.056945f
C4837 ASIG5V.n6723 VSS 0.056945f
C4838 ASIG5V.n6724 VSS 0.056945f
C4839 ASIG5V.n6725 VSS 0.056945f
C4840 ASIG5V.n6726 VSS 0.056945f
C4841 ASIG5V.n6727 VSS 0.056945f
C4842 ASIG5V.n6728 VSS 0.056945f
C4843 ASIG5V.n6729 VSS 0.056945f
C4844 ASIG5V.n6730 VSS 0.056945f
C4845 ASIG5V.n6731 VSS 0.056945f
C4846 ASIG5V.n6732 VSS 0.056945f
C4847 ASIG5V.n6733 VSS 0.056945f
C4848 ASIG5V.n6734 VSS 0.056945f
C4849 ASIG5V.n6735 VSS 0.056945f
C4850 ASIG5V.n6736 VSS 0.056945f
C4851 ASIG5V.n6737 VSS 0.056945f
C4852 ASIG5V.n6738 VSS 0.056945f
C4853 ASIG5V.n6739 VSS 0.056945f
C4854 ASIG5V.n6740 VSS 0.056945f
C4855 ASIG5V.n6741 VSS 0.056945f
C4856 ASIG5V.n6742 VSS 0.056945f
C4857 ASIG5V.n6743 VSS 0.056945f
C4858 ASIG5V.n6744 VSS 0.056945f
C4859 ASIG5V.n6745 VSS 0.056945f
C4860 ASIG5V.n6746 VSS 0.056945f
C4861 ASIG5V.n6747 VSS 0.056945f
C4862 ASIG5V.n6748 VSS 0.056945f
C4863 ASIG5V.n6749 VSS 0.056945f
C4864 ASIG5V.n6750 VSS 0.056945f
C4865 ASIG5V.n6751 VSS 0.056945f
C4866 ASIG5V.n6752 VSS 0.056945f
C4867 ASIG5V.n6753 VSS 0.056945f
C4868 ASIG5V.n6754 VSS 0.056945f
C4869 ASIG5V.n6755 VSS 0.056945f
C4870 ASIG5V.n6756 VSS 0.056945f
C4871 ASIG5V.n6757 VSS 0.056945f
C4872 ASIG5V.n6758 VSS 0.056945f
C4873 ASIG5V.n6759 VSS 0.056945f
C4874 ASIG5V.n6760 VSS 0.056945f
C4875 ASIG5V.n6761 VSS 0.056945f
C4876 ASIG5V.n6762 VSS 0.056945f
C4877 ASIG5V.n6763 VSS 0.056945f
C4878 ASIG5V.n6764 VSS 0.056945f
C4879 ASIG5V.n6765 VSS 0.056945f
C4880 ASIG5V.n6766 VSS 0.056945f
C4881 ASIG5V.n6767 VSS 0.056945f
C4882 ASIG5V.n6768 VSS 0.056945f
C4883 ASIG5V.n6769 VSS 0.056945f
C4884 ASIG5V.n6770 VSS 0.056945f
C4885 ASIG5V.n6771 VSS 0.056945f
C4886 ASIG5V.n6772 VSS 0.056945f
C4887 ASIG5V.n6773 VSS 0.056945f
C4888 ASIG5V.n6774 VSS 0.056945f
C4889 ASIG5V.n6775 VSS 0.056945f
C4890 ASIG5V.n6776 VSS 0.056945f
C4891 ASIG5V.n6777 VSS 0.056945f
C4892 ASIG5V.n6778 VSS 0.056945f
C4893 ASIG5V.n6779 VSS 0.056945f
C4894 ASIG5V.n6780 VSS 0.056945f
C4895 ASIG5V.n6781 VSS 0.056945f
C4896 ASIG5V.n6782 VSS 0.056945f
C4897 ASIG5V.n6783 VSS 0.056945f
C4898 ASIG5V.n6784 VSS 0.056945f
C4899 ASIG5V.n6785 VSS 0.056945f
C4900 ASIG5V.n6786 VSS 0.056945f
C4901 ASIG5V.n6787 VSS 0.056945f
C4902 ASIG5V.n6788 VSS 0.056945f
C4903 ASIG5V.n6789 VSS 0.056945f
C4904 ASIG5V.n6790 VSS 0.056945f
C4905 ASIG5V.n6791 VSS 0.056945f
C4906 ASIG5V.n6792 VSS 0.056945f
C4907 ASIG5V.n6793 VSS 0.056945f
C4908 ASIG5V.n6794 VSS 0.056945f
C4909 ASIG5V.n6795 VSS 0.056945f
C4910 ASIG5V.n6796 VSS 0.056945f
C4911 ASIG5V.n6797 VSS 0.056945f
C4912 ASIG5V.n6798 VSS 0.056945f
C4913 ASIG5V.n6799 VSS 0.056945f
C4914 ASIG5V.n6800 VSS 0.056945f
C4915 ASIG5V.n6801 VSS 0.056945f
C4916 ASIG5V.n6802 VSS 0.056945f
C4917 ASIG5V.n6803 VSS 0.056945f
C4918 ASIG5V.n6804 VSS 0.056945f
C4919 ASIG5V.n6805 VSS 0.056945f
C4920 ASIG5V.n6806 VSS 0.056945f
C4921 ASIG5V.n6807 VSS 0.056945f
C4922 ASIG5V.n6808 VSS 0.056945f
C4923 ASIG5V.n6809 VSS 0.056945f
C4924 ASIG5V.n6810 VSS 0.056945f
C4925 ASIG5V.n6811 VSS 0.056945f
C4926 ASIG5V.n6812 VSS 0.056945f
C4927 ASIG5V.n6813 VSS 0.056945f
C4928 ASIG5V.n6814 VSS 0.056945f
C4929 ASIG5V.n6815 VSS 0.056945f
C4930 ASIG5V.n6816 VSS 0.056945f
C4931 ASIG5V.n6817 VSS 0.056945f
C4932 ASIG5V.n6818 VSS 0.056945f
C4933 ASIG5V.n6819 VSS 0.056945f
C4934 ASIG5V.n6820 VSS 0.056945f
C4935 ASIG5V.n6821 VSS 0.056945f
C4936 ASIG5V.n6822 VSS 0.056945f
C4937 ASIG5V.n6823 VSS 0.056945f
C4938 ASIG5V.n6824 VSS 0.056945f
C4939 ASIG5V.n6825 VSS 0.056945f
C4940 ASIG5V.n6826 VSS 0.056945f
C4941 ASIG5V.n6827 VSS 0.056945f
C4942 ASIG5V.n6828 VSS 0.056945f
C4943 ASIG5V.n6829 VSS 0.056945f
C4944 ASIG5V.n6830 VSS 0.056945f
C4945 ASIG5V.n6831 VSS 0.056945f
C4946 ASIG5V.n6832 VSS 0.056945f
C4947 ASIG5V.n6833 VSS 0.056945f
C4948 ASIG5V.n6834 VSS 0.056945f
C4949 ASIG5V.n6835 VSS 0.056945f
C4950 ASIG5V.n6836 VSS 0.056945f
C4951 ASIG5V.n6837 VSS 0.056945f
C4952 ASIG5V.n6838 VSS 0.056945f
C4953 ASIG5V.n6839 VSS 0.056945f
C4954 ASIG5V.n6840 VSS 0.056945f
C4955 ASIG5V.n6841 VSS 0.056945f
C4956 ASIG5V.n6842 VSS 0.056945f
C4957 ASIG5V.n6843 VSS 0.056945f
C4958 ASIG5V.n6844 VSS 0.056945f
C4959 ASIG5V.n6845 VSS 0.056945f
C4960 ASIG5V.n6846 VSS 0.056945f
C4961 ASIG5V.n6847 VSS 0.056945f
C4962 ASIG5V.n6848 VSS 0.056945f
C4963 ASIG5V.n6849 VSS 0.056945f
C4964 ASIG5V.n6850 VSS 0.056945f
C4965 ASIG5V.n6851 VSS 0.056945f
C4966 ASIG5V.n6852 VSS 0.056945f
C4967 ASIG5V.n6853 VSS 0.056945f
C4968 ASIG5V.n6854 VSS 0.056945f
C4969 ASIG5V.n6855 VSS 0.056945f
C4970 ASIG5V.n6856 VSS 0.056945f
C4971 ASIG5V.n6857 VSS 0.056945f
C4972 ASIG5V.n6858 VSS 0.056945f
C4973 ASIG5V.n6859 VSS 0.056945f
C4974 ASIG5V.n6860 VSS 0.056945f
C4975 ASIG5V.n6861 VSS 0.056945f
C4976 ASIG5V.n6862 VSS 0.056945f
C4977 ASIG5V.n6863 VSS 0.056945f
C4978 ASIG5V.n6864 VSS 0.056945f
C4979 ASIG5V.n6865 VSS 0.056945f
C4980 ASIG5V.n6866 VSS 0.056945f
C4981 ASIG5V.n6867 VSS 0.056945f
C4982 ASIG5V.n6868 VSS 0.056945f
C4983 ASIG5V.n6869 VSS 0.056945f
C4984 ASIG5V.n6870 VSS 0.056945f
C4985 ASIG5V.n6871 VSS 0.056945f
C4986 ASIG5V.n6872 VSS 0.056945f
C4987 ASIG5V.n6873 VSS 0.056945f
C4988 ASIG5V.n6874 VSS 0.056945f
C4989 ASIG5V.n6875 VSS 0.056945f
C4990 ASIG5V.n6876 VSS 0.056945f
C4991 ASIG5V.n6877 VSS 0.056945f
C4992 ASIG5V.n6878 VSS 0.056945f
C4993 ASIG5V.n6879 VSS 0.056945f
C4994 ASIG5V.n6880 VSS 0.047722f
C4995 ASIG5V.n6881 VSS 0.051049f
C4996 ASIG5V.n6882 VSS 0.051049f
C4997 ASIG5V.n6883 VSS 0.076709f
C4998 ASIG5V.n6884 VSS 0.064014f
C4999 ASIG5V.n6885 VSS 0.044584f
C5000 ASIG5V.n6886 VSS 0.052746f
C5001 ASIG5V.n6887 VSS 0.052746f
C5002 ASIG5V.n6888 VSS 0.045974f
C5003 ASIG5V.n6889 VSS 0.076709f
C5004 ASIG5V.n6890 VSS 0.045974f
C5005 ASIG5V.n6891 VSS 0.608692f
C5006 ASIG5V.n6892 VSS 0.747381f
C5007 ASIG5V.n6893 VSS 0.0621f
C5008 ASIG5V.n6894 VSS 0.108961f
C5009 ASIG5V.n6895 VSS 0.0621f
C5010 ASIG5V.n6896 VSS 0.108961f
C5011 ASIG5V.n6897 VSS 0.056945f
C5012 ASIG5V.n6898 VSS 0.056945f
C5013 ASIG5V.n6900 VSS 0.056945f
C5014 ASIG5V.n6901 VSS 0.056945f
C5015 ASIG5V.n6902 VSS 0.056945f
C5016 ASIG5V.n6903 VSS 0.056945f
C5017 ASIG5V.n6906 VSS 0.056945f
C5018 ASIG5V.n6907 VSS 0.056945f
C5019 ASIG5V.n6908 VSS 0.056945f
C5020 ASIG5V.n6909 VSS 0.056945f
C5021 ASIG5V.n6912 VSS 0.056945f
C5022 ASIG5V.n6913 VSS 0.056945f
C5023 ASIG5V.n6914 VSS 0.056945f
C5024 ASIG5V.n6915 VSS 0.056945f
C5025 ASIG5V.n6918 VSS 0.056945f
C5026 ASIG5V.n6919 VSS 0.056945f
C5027 ASIG5V.n6920 VSS 0.056945f
C5028 ASIG5V.n6921 VSS 0.056945f
C5029 ASIG5V.n6924 VSS 0.056945f
C5030 ASIG5V.n6925 VSS 0.056945f
C5031 ASIG5V.n6926 VSS 0.056945f
C5032 ASIG5V.n6927 VSS 0.056945f
C5033 ASIG5V.n6930 VSS 0.056945f
C5034 ASIG5V.n6931 VSS 0.056945f
C5035 ASIG5V.n6932 VSS 0.056945f
C5036 ASIG5V.n6933 VSS 0.056945f
C5037 ASIG5V.n6936 VSS 0.056945f
C5038 ASIG5V.n6937 VSS 0.056945f
C5039 ASIG5V.n6938 VSS 0.056945f
C5040 ASIG5V.n6939 VSS 0.056945f
C5041 ASIG5V.n6942 VSS 0.056945f
C5042 ASIG5V.n6943 VSS 0.056945f
C5043 ASIG5V.n6944 VSS 0.056945f
C5044 ASIG5V.n6945 VSS 0.056945f
C5045 ASIG5V.n6948 VSS 0.056945f
C5046 ASIG5V.n6949 VSS 0.056945f
C5047 ASIG5V.n6950 VSS 0.056945f
C5048 ASIG5V.n6951 VSS 0.056945f
C5049 ASIG5V.n6954 VSS 0.056945f
C5050 ASIG5V.n6955 VSS 0.056945f
C5051 ASIG5V.n6956 VSS 0.056945f
C5052 ASIG5V.n6957 VSS 0.056945f
C5053 ASIG5V.n6960 VSS 0.056945f
C5054 ASIG5V.n6961 VSS 0.056945f
C5055 ASIG5V.n6962 VSS 0.056945f
C5056 ASIG5V.n6963 VSS 0.056945f
C5057 ASIG5V.n6966 VSS 0.056945f
C5058 ASIG5V.n6967 VSS 0.056945f
C5059 ASIG5V.n6968 VSS 0.056945f
C5060 ASIG5V.n6969 VSS 0.056945f
C5061 ASIG5V.n6972 VSS 0.056945f
C5062 ASIG5V.n6973 VSS 0.056945f
C5063 ASIG5V.n6974 VSS 0.056945f
C5064 ASIG5V.n6975 VSS 0.056945f
C5065 ASIG5V.n6978 VSS 0.056945f
C5066 ASIG5V.n6979 VSS 0.056945f
C5067 ASIG5V.n6980 VSS 0.056945f
C5068 ASIG5V.n6981 VSS 0.056945f
C5069 ASIG5V.n6984 VSS 0.056945f
C5070 ASIG5V.n6985 VSS 0.056945f
C5071 ASIG5V.n6986 VSS 0.056945f
C5072 ASIG5V.n6987 VSS 0.056945f
C5073 ASIG5V.n6990 VSS 0.056945f
C5074 ASIG5V.n6991 VSS 0.056945f
C5075 ASIG5V.n6992 VSS 0.056945f
C5076 ASIG5V.n6993 VSS 0.056945f
C5077 ASIG5V.n6996 VSS 0.056945f
C5078 ASIG5V.n6997 VSS 0.056945f
C5079 ASIG5V.n6998 VSS 0.056945f
C5080 ASIG5V.n6999 VSS 0.056945f
C5081 ASIG5V.n7002 VSS 0.056945f
C5082 ASIG5V.n7003 VSS 0.056945f
C5083 ASIG5V.n7004 VSS 0.056945f
C5084 ASIG5V.n7005 VSS 0.056945f
C5085 ASIG5V.n7008 VSS 0.056945f
C5086 ASIG5V.n7009 VSS 0.056945f
C5087 ASIG5V.n7010 VSS 0.056945f
C5088 ASIG5V.n7011 VSS 0.056945f
C5089 ASIG5V.n7014 VSS 0.056945f
C5090 ASIG5V.n7015 VSS 0.056945f
C5091 ASIG5V.n7016 VSS 0.056945f
C5092 ASIG5V.n7017 VSS 0.056945f
C5093 ASIG5V.n7020 VSS 0.036092f
C5094 ASIG5V.n7021 VSS 0.036092f
C5095 ASIG5V.n7022 VSS 0.047722f
C5096 ASIG5V.n7023 VSS 0.056945f
C5097 ASIG5V.n7024 VSS 0.056945f
C5098 ASIG5V.n7025 VSS 0.056945f
C5099 ASIG5V.n7027 VSS 0.056945f
C5100 ASIG5V.n7029 VSS 0.056945f
C5101 ASIG5V.n7030 VSS 0.056945f
C5102 ASIG5V.n7031 VSS 0.056945f
C5103 ASIG5V.n7032 VSS 0.056945f
C5104 ASIG5V.n7033 VSS 0.056945f
C5105 ASIG5V.n7034 VSS 0.056945f
C5106 ASIG5V.n7035 VSS 0.056945f
C5107 ASIG5V.n7037 VSS 0.056945f
C5108 ASIG5V.n7039 VSS 0.056945f
C5109 ASIG5V.n7040 VSS 0.056945f
C5110 ASIG5V.n7041 VSS 0.056945f
C5111 ASIG5V.n7042 VSS 0.056945f
C5112 ASIG5V.n7043 VSS 0.056945f
C5113 ASIG5V.n7044 VSS 0.056945f
C5114 ASIG5V.n7045 VSS 0.056945f
C5115 ASIG5V.n7047 VSS 0.056945f
C5116 ASIG5V.n7049 VSS 0.056945f
C5117 ASIG5V.n7050 VSS 0.056945f
C5118 ASIG5V.n7051 VSS 0.056945f
C5119 ASIG5V.n7052 VSS 0.056945f
C5120 ASIG5V.n7053 VSS 0.056945f
C5121 ASIG5V.n7054 VSS 0.056945f
C5122 ASIG5V.n7055 VSS 0.056945f
C5123 ASIG5V.n7057 VSS 0.056945f
C5124 ASIG5V.n7059 VSS 0.056945f
C5125 ASIG5V.n7060 VSS 0.056945f
C5126 ASIG5V.n7061 VSS 0.056945f
C5127 ASIG5V.n7062 VSS 0.056945f
C5128 ASIG5V.n7063 VSS 0.056945f
C5129 ASIG5V.n7064 VSS 0.056945f
C5130 ASIG5V.n7065 VSS 0.056945f
C5131 ASIG5V.n7067 VSS 0.056945f
C5132 ASIG5V.n7069 VSS 0.056945f
C5133 ASIG5V.n7070 VSS 0.056945f
C5134 ASIG5V.n7071 VSS 0.056945f
C5135 ASIG5V.n7072 VSS 0.056945f
C5136 ASIG5V.n7073 VSS 0.056945f
C5137 ASIG5V.n7074 VSS 0.056945f
C5138 ASIG5V.n7075 VSS 0.056945f
C5139 ASIG5V.n7077 VSS 0.056945f
C5140 ASIG5V.n7079 VSS 0.056945f
C5141 ASIG5V.n7080 VSS 0.056945f
C5142 ASIG5V.n7081 VSS 0.056945f
C5143 ASIG5V.n7082 VSS 0.056945f
C5144 ASIG5V.n7083 VSS 0.056945f
C5145 ASIG5V.n7084 VSS 0.056945f
C5146 ASIG5V.n7085 VSS 0.056945f
C5147 ASIG5V.n7087 VSS 0.056945f
C5148 ASIG5V.n7089 VSS 0.056945f
C5149 ASIG5V.n7090 VSS 0.056945f
C5150 ASIG5V.n7091 VSS 0.056945f
C5151 ASIG5V.n7092 VSS 0.056945f
C5152 ASIG5V.n7093 VSS 0.056945f
C5153 ASIG5V.n7094 VSS 0.056945f
C5154 ASIG5V.n7095 VSS 0.056945f
C5155 ASIG5V.n7097 VSS 0.056945f
C5156 ASIG5V.n7099 VSS 0.056945f
C5157 ASIG5V.n7100 VSS 0.056945f
C5158 ASIG5V.n7101 VSS 0.056945f
C5159 ASIG5V.n7102 VSS 0.056945f
C5160 ASIG5V.n7103 VSS 0.056945f
C5161 ASIG5V.n7104 VSS 0.056945f
C5162 ASIG5V.n7105 VSS 0.056945f
C5163 ASIG5V.n7107 VSS 0.056945f
C5164 ASIG5V.n7109 VSS 0.056945f
C5165 ASIG5V.n7110 VSS 0.056945f
C5166 ASIG5V.n7111 VSS 0.056945f
C5167 ASIG5V.n7112 VSS 0.056945f
C5168 ASIG5V.n7113 VSS 0.056945f
C5169 ASIG5V.n7114 VSS 0.056945f
C5170 ASIG5V.n7115 VSS 0.056945f
C5171 ASIG5V.n7117 VSS 0.056945f
C5172 ASIG5V.n7119 VSS 0.056945f
C5173 ASIG5V.n7120 VSS 0.056945f
C5174 ASIG5V.n7121 VSS 0.056945f
C5175 ASIG5V.n7122 VSS 0.056945f
C5176 ASIG5V.n7123 VSS 0.056945f
C5177 ASIG5V.n7124 VSS 0.056945f
C5178 ASIG5V.n7125 VSS 0.056945f
C5179 ASIG5V.n7127 VSS 0.056945f
C5180 ASIG5V.n7129 VSS 0.056945f
C5181 ASIG5V.n7130 VSS 0.056945f
C5182 ASIG5V.n7131 VSS 0.056945f
C5183 ASIG5V.n7132 VSS 0.056945f
C5184 ASIG5V.n7133 VSS 0.056945f
C5185 ASIG5V.n7134 VSS 0.056945f
C5186 ASIG5V.n7135 VSS 0.056945f
C5187 ASIG5V.n7137 VSS 0.056945f
C5188 ASIG5V.n7139 VSS 0.056945f
C5189 ASIG5V.n7140 VSS 0.056945f
C5190 ASIG5V.n7141 VSS 0.056945f
C5191 ASIG5V.n7142 VSS 0.056945f
C5192 ASIG5V.n7143 VSS 0.056945f
C5193 ASIG5V.n7144 VSS 0.056945f
C5194 ASIG5V.n7145 VSS 0.056945f
C5195 ASIG5V.n7147 VSS 0.056945f
C5196 ASIG5V.n7149 VSS 0.056945f
C5197 ASIG5V.n7150 VSS 0.056945f
C5198 ASIG5V.n7151 VSS 0.056945f
C5199 ASIG5V.n7152 VSS 0.056945f
C5200 ASIG5V.n7153 VSS 0.056945f
C5201 ASIG5V.n7154 VSS 0.056945f
C5202 ASIG5V.n7155 VSS 0.056945f
C5203 ASIG5V.n7157 VSS 0.056945f
C5204 ASIG5V.n7159 VSS 0.056945f
C5205 ASIG5V.n7160 VSS 0.056945f
C5206 ASIG5V.n7161 VSS 0.056945f
C5207 ASIG5V.n7162 VSS 0.056945f
C5208 ASIG5V.n7163 VSS 0.056945f
C5209 ASIG5V.n7164 VSS 0.056945f
C5210 ASIG5V.n7165 VSS 0.056945f
C5211 ASIG5V.n7167 VSS 0.056945f
C5212 ASIG5V.n7169 VSS 0.056945f
C5213 ASIG5V.n7170 VSS 0.056945f
C5214 ASIG5V.n7171 VSS 0.056945f
C5215 ASIG5V.n7172 VSS 0.056945f
C5216 ASIG5V.n7173 VSS 0.056945f
C5217 ASIG5V.n7174 VSS 0.056945f
C5218 ASIG5V.n7175 VSS 0.056945f
C5219 ASIG5V.n7177 VSS 0.056945f
C5220 ASIG5V.n7179 VSS 0.056945f
C5221 ASIG5V.n7180 VSS 0.056945f
C5222 ASIG5V.n7181 VSS 0.056945f
C5223 ASIG5V.n7182 VSS 0.056945f
C5224 ASIG5V.n7183 VSS 0.056945f
C5225 ASIG5V.n7184 VSS 0.056945f
C5226 ASIG5V.n7185 VSS 0.056945f
C5227 ASIG5V.n7187 VSS 0.056945f
C5228 ASIG5V.n7189 VSS 0.056945f
C5229 ASIG5V.n7190 VSS 0.056945f
C5230 ASIG5V.n7191 VSS 0.056945f
C5231 ASIG5V.n7192 VSS 0.056945f
C5232 ASIG5V.n7193 VSS 0.056945f
C5233 ASIG5V.n7194 VSS 0.056945f
C5234 ASIG5V.n7195 VSS 0.056945f
C5235 ASIG5V.n7197 VSS 0.056945f
C5236 ASIG5V.n7199 VSS 0.056945f
C5237 ASIG5V.n7200 VSS 0.056945f
C5238 ASIG5V.n7201 VSS 0.056945f
C5239 ASIG5V.n7202 VSS 0.056945f
C5240 ASIG5V.n7203 VSS 0.056945f
C5241 ASIG5V.n7204 VSS 0.056945f
C5242 ASIG5V.n7205 VSS 0.056945f
C5243 ASIG5V.n7207 VSS 0.056945f
C5244 ASIG5V.n7209 VSS 0.056945f
C5245 ASIG5V.n7210 VSS 0.056945f
C5246 ASIG5V.n7211 VSS 0.056945f
C5247 ASIG5V.n7212 VSS 0.056945f
C5248 ASIG5V.n7213 VSS 0.056945f
C5249 ASIG5V.n7214 VSS 0.056945f
C5250 ASIG5V.n7215 VSS 0.056945f
C5251 ASIG5V.n7217 VSS 0.056945f
C5252 ASIG5V.n7219 VSS 0.056945f
C5253 ASIG5V.n7220 VSS 0.056945f
C5254 ASIG5V.n7221 VSS 0.056945f
C5255 ASIG5V.n7222 VSS 0.056945f
C5256 ASIG5V.n7223 VSS 0.056945f
C5257 ASIG5V.n7224 VSS 0.056945f
C5258 ASIG5V.n7225 VSS 0.056945f
C5259 ASIG5V.n7227 VSS 0.056945f
C5260 ASIG5V.n7229 VSS 0.036092f
C5261 ASIG5V.n7230 VSS 0.036092f
C5262 ASIG5V.n7231 VSS 0.052133f
C5263 ASIG5V.n7232 VSS 0.09726f
C5264 ASIG5V.n7233 VSS 0.108961f
C5265 ASIG5V.n7234 VSS 0.069023f
C5266 ASIG5V.n7235 VSS 0.077327f
C5267 ASIG5V.n7236 VSS 0.077327f
C5268 ASIG5V.n7237 VSS 0.108961f
C5269 ASIG5V.n7238 VSS 1.0941f
C5270 ASIG5V.n7239 VSS 0.955415f
C5271 ASIG5V.n7240 VSS 0.662626f
C5272 ASIG5V.n7241 VSS 0.098416f
C5273 ASIG5V.n7242 VSS 0.098416f
C5274 ASIG5V.n7243 VSS 0.087848f
C5275 ASIG5V.n7244 VSS 0.07229f
C5276 ASIG5V.n7247 VSS 0.314214f
C5277 ASIG5V.n7248 VSS 0.074298f
C5278 ASIG5V.n7250 VSS 0.074298f
C5279 ASIG5V.n7253 VSS 0.087753f
C5280 ASIG5V.n7254 VSS 0.087753f
C5281 ASIG5V.t2 VSS 7.07689f
C5282 ASIG5V.n7258 VSS 0.314214f
C5283 ASIG5V.n7259 VSS 0.074298f
C5284 ASIG5V.n7261 VSS 0.074298f
C5285 ASIG5V.n7264 VSS 0.087753f
C5286 ASIG5V.n7265 VSS 0.087753f
C5287 ASIG5V.t3 VSS 7.07689f
C5288 ASIG5V.n7269 VSS 0.314214f
C5289 ASIG5V.n7270 VSS 0.074298f
C5290 ASIG5V.n7271 VSS 0.074298f
C5291 ASIG5V.n7272 VSS 0.087753f
C5292 ASIG5V.n7274 VSS 0.309175f
C5293 ASIG5V.n7277 VSS 0.087753f
C5294 ASIG5V.n7279 VSS 0.074298f
C5295 ASIG5V.n7283 VSS 0.309175f
C5296 ASIG5V.n7284 VSS 0.087753f
C5297 ASIG5V.n7286 VSS 0.074298f
C5298 ASIG5V.n7287 VSS 0.314214f
C5299 ASIG5V.t7 VSS 7.07689f
C5300 ASIG5V.n7290 VSS 0.074298f
C5301 ASIG5V.n7291 VSS 0.074298f
C5302 ASIG5V.n7292 VSS 0.087753f
C5303 ASIG5V.n7294 VSS 0.845738f
C5304 ASIG5V.n7297 VSS 0.087753f
C5305 ASIG5V.n7299 VSS 0.074298f
C5306 ASIG5V.n7303 VSS 0.309175f
C5307 ASIG5V.n7304 VSS 0.087753f
C5308 ASIG5V.n7306 VSS 0.074298f
C5309 ASIG5V.n7307 VSS 0.314214f
C5310 ASIG5V.n7310 VSS 0.314214f
C5311 ASIG5V.n7311 VSS 0.074298f
C5312 ASIG5V.n7312 VSS 0.074298f
C5313 ASIG5V.n7313 VSS 0.087753f
C5314 ASIG5V.n7315 VSS 0.309175f
C5315 ASIG5V.n7318 VSS 0.087753f
C5316 ASIG5V.n7320 VSS 0.074298f
C5317 ASIG5V.n7326 VSS 0.074298f
C5318 ASIG5V.n7328 VSS 0.314214f
C5319 ASIG5V.n7330 VSS 0.074298f
C5320 ASIG5V.n7332 VSS 0.314214f
C5321 ASIG5V.n7334 VSS 0.074298f
C5322 ASIG5V.n7337 VSS 0.074298f
C5323 ASIG5V.n7338 VSS 0.309175f
C5324 ASIG5V.n7339 VSS 0.021962f
C5325 ASIG5V.n7340 VSS 0.548344f
C5326 ASIG5V.n7341 VSS 0.536863f
C5327 ASIG5V.n7344 VSS 0.087753f
C5328 ASIG5V.n7346 VSS 0.074298f
C5329 ASIG5V.n7349 VSS 0.074298f
C5330 ASIG5V.n7351 VSS 0.074298f
C5331 ASIG5V.n7354 VSS 0.087753f
C5332 ASIG5V.n7355 VSS 0.087753f
C5333 ASIG5V.n7357 VSS 0.074298f
C5334 ASIG5V.n7361 VSS 0.087753f
C5335 ASIG5V.n7363 VSS 0.074298f
C5336 ASIG5V.n7366 VSS 0.087753f
C5337 ASIG5V.n7367 VSS 0.074298f
C5338 ASIG5V.n7369 VSS 0.314214f
C5339 ASIG5V.n7370 VSS 0.074298f
C5340 ASIG5V.n7373 VSS 0.074298f
C5341 ASIG5V.n7375 VSS 0.087753f
C5342 ASIG5V.n7377 VSS 0.309175f
C5343 ASIG5V.n7378 VSS 0.309175f
C5344 ASIG5V.n7379 VSS 0.314214f
C5345 ASIG5V.n7381 VSS 0.074298f
C5346 ASIG5V.n7383 VSS 0.087753f
C5347 ASIG5V.n7385 VSS 0.309175f
C5348 ASIG5V.n7386 VSS 0.314214f
C5349 ASIG5V.n7387 VSS 0.314214f
C5350 ASIG5V.n7388 VSS 0.074298f
C5351 ASIG5V.n7390 VSS 0.250522f
C5352 ASIG5V.n7391 VSS 0.309175f
C5353 ASIG5V.n7392 VSS 0.309175f
C5354 ASIG5V.n7395 VSS 0.087753f
C5355 ASIG5V.n7397 VSS 0.087753f
C5356 ASIG5V.n7399 VSS 0.074298f
C5357 ASIG5V.n7401 VSS 0.250522f
C5358 ASIG5V.n7402 VSS 0.074298f
C5359 ASIG5V.n7404 VSS 0.314214f
C5360 ASIG5V.n7406 VSS 0.087753f
C5361 ASIG5V.n7408 VSS 0.074298f
C5362 ASIG5V.n7410 VSS 0.314214f
C5363 ASIG5V.n7411 VSS 0.074298f
C5364 ASIG5V.n7413 VSS 0.314214f
C5365 ASIG5V.n7414 VSS 0.314214f
C5366 ASIG5V.n7416 VSS 0.074298f
C5367 ASIG5V.n7418 VSS 0.074298f
C5368 ASIG5V.n7420 VSS 0.074298f
C5369 ASIG5V.n7422 VSS 0.087753f
C5370 ASIG5V.n7424 VSS 0.087753f
C5371 ASIG5V.n7426 VSS 0.309175f
C5372 ASIG5V.n7427 VSS 0.309175f
C5373 ASIG5V.n7429 VSS 0.074298f
C5374 ASIG5V.n7431 VSS 0.074298f
C5375 ASIG5V.n7433 VSS 0.087753f
C5376 ASIG5V.n7435 VSS 0.087753f
C5377 ASIG5V.n7437 VSS 0.309175f
C5378 ASIG5V.n7438 VSS 0.309175f
C5379 ASIG5V.n7440 VSS 0.074298f
C5380 ASIG5V.n7442 VSS 0.074298f
C5381 ASIG5V.n7444 VSS 0.087753f
C5382 ASIG5V.n7446 VSS 0.087753f
C5383 ASIG5V.n7448 VSS 0.309175f
C5384 ASIG5V.n7449 VSS 0.309175f
C5385 ASIG5V.n7451 VSS 0.074298f
C5386 ASIG5V.n7453 VSS 0.074298f
C5387 ASIG5V.n7455 VSS 0.087753f
C5388 ASIG5V.n7457 VSS 0.087753f
C5389 ASIG5V.n7459 VSS 0.845738f
C5390 ASIG5V.n7460 VSS 0.087753f
C5391 ASIG5V.n7461 VSS 0.074298f
C5392 ASIG5V.n7464 VSS 0.314214f
C5393 ASIG5V.n7465 VSS 0.074298f
C5394 ASIG5V.n7466 VSS 0.074298f
C5395 ASIG5V.n7467 VSS 0.087753f
C5396 ASIG5V.n7469 VSS 0.087753f
C5397 ASIG5V.n7470 VSS 0.074298f
C5398 ASIG5V.n7472 VSS 0.074298f
C5399 ASIG5V.n7474 VSS 0.074298f
C5400 ASIG5V.n7475 VSS 0.309175f
C5401 ASIG5V.n7476 VSS 0.309175f
C5402 ASIG5V.n7479 VSS 0.087753f
C5403 ASIG5V.n7481 VSS 0.074298f
C5404 ASIG5V.n7482 VSS 0.309175f
C5405 ASIG5V.n7483 VSS 0.309175f
C5406 ASIG5V.n7486 VSS 0.087753f
C5407 ASIG5V.n7488 VSS 0.074298f
C5408 ASIG5V.n7489 VSS 0.309175f
C5409 ASIG5V.n7490 VSS 0.309175f
C5410 ASIG5V.n7493 VSS 0.087753f
C5411 ASIG5V.n7495 VSS 0.074298f
C5412 ASIG5V.n7496 VSS 0.309175f
C5413 ASIG5V.n7497 VSS 0.309175f
C5414 ASIG5V.n7500 VSS 0.087753f
C5415 ASIG5V.n7502 VSS 0.074298f
C5416 ASIG5V.n7503 VSS 0.309175f
C5417 ASIG5V.n7507 VSS 0.074298f
C5418 ASIG5V.n7508 VSS 0.314214f
C5419 ASIG5V.n7512 VSS 0.074298f
C5420 ASIG5V.n7513 VSS 0.314214f
C5421 ASIG5V.n7517 VSS 0.074298f
C5422 ASIG5V.n7518 VSS 0.314214f
C5423 ASIG5V.n7522 VSS 0.074298f
C5424 ASIG5V.n7523 VSS 0.314214f
C5425 ASIG5V.n7527 VSS 0.074298f
C5426 ASIG5V.n7528 VSS 0.314214f
C5427 ASIG5V.n7532 VSS 0.074298f
C5428 ASIG5V.n7533 VSS 0.074298f
C5429 ASIG5V.n7537 VSS 0.087753f
C5430 ASIG5V.n7538 VSS 0.074298f
C5431 ASIG5V.n7540 VSS 0.087753f
C5432 ASIG5V.n7541 VSS 0.074298f
C5433 ASIG5V.n7544 VSS 0.074298f
C5434 ASIG5V.n7546 VSS 0.087753f
C5435 ASIG5V.n7547 VSS 0.074298f
C5436 ASIG5V.n7549 VSS 0.087753f
C5437 ASIG5V.n7550 VSS 0.074298f
C5438 ASIG5V.n7552 VSS 0.314214f
C5439 ASIG5V.n7554 VSS 0.087753f
C5440 ASIG5V.n7555 VSS 0.074298f
C5441 ASIG5V.n7557 VSS 0.314214f
C5442 ASIG5V.n7559 VSS 0.087753f
C5443 ASIG5V.n7560 VSS 0.074298f
C5444 ASIG5V.n7562 VSS 0.074298f
C5445 ASIG5V.n7566 VSS 0.309175f
C5446 ASIG5V.n7567 VSS 0.087753f
C5447 ASIG5V.n7569 VSS 0.074298f
C5448 ASIG5V.n7570 VSS 0.074298f
C5449 ASIG5V.n7575 VSS 0.087753f
C5450 ASIG5V.n7577 VSS 0.074298f
C5451 ASIG5V.n7581 VSS 0.074298f
C5452 ASIG5V.n7582 VSS 0.074298f
C5453 ASIG5V.n7585 VSS 0.074298f
C5454 ASIG5V.n7587 VSS 0.087753f
C5455 ASIG5V.n7588 VSS 0.087753f
C5456 ASIG5V.n7590 VSS 0.309175f
C5457 ASIG5V.n7591 VSS 0.250522f
C5458 ASIG5V.n7592 VSS 0.845738f
C5459 ASIG5V.n7593 VSS 0.845738f
C5460 ASIG5V.n7595 VSS 0.074298f
C5461 ASIG5V.n7598 VSS 0.087753f
C5462 ASIG5V.n7601 VSS 0.087753f
C5463 ASIG5V.n7602 VSS 0.074298f
C5464 ASIG5V.n7604 VSS 0.250522f
C5465 ASIG5V.t6 VSS 7.07689f
C5466 ASIG5V.n7607 VSS 0.845738f
C5467 ASIG5V.n7609 VSS 0.074298f
C5468 ASIG5V.n7610 VSS 0.087753f
C5469 ASIG5V.n7612 VSS 0.074298f
C5470 ASIG5V.n7613 VSS 0.074298f
C5471 ASIG5V.n7615 VSS 0.250522f
C5472 ASIG5V.n7617 VSS 0.309175f
C5473 ASIG5V.n7618 VSS 0.087753f
C5474 ASIG5V.n7620 VSS 0.074298f
C5475 ASIG5V.n7623 VSS 0.087753f
C5476 ASIG5V.n7624 VSS 0.309175f
C5477 ASIG5V.n7626 VSS 0.074298f
C5478 ASIG5V.n7628 VSS 0.074298f
C5479 ASIG5V.n7630 VSS 0.087753f
C5480 ASIG5V.n7631 VSS 0.074298f
C5481 ASIG5V.n7633 VSS 0.309175f
C5482 ASIG5V.n7635 VSS 0.314214f
C5483 ASIG5V.n7636 VSS 0.309175f
C5484 ASIG5V.n7637 VSS 0.314214f
C5485 ASIG5V.n7639 VSS 0.074298f
C5486 ASIG5V.n7641 VSS 0.087753f
C5487 ASIG5V.n7643 VSS 0.309175f
C5488 ASIG5V.n7644 VSS 0.250522f
C5489 ASIG5V.t0 VSS 7.07689f
C5490 ASIG5V.n7645 VSS 0.309175f
C5491 ASIG5V.n7646 VSS 0.250522f
C5492 ASIG5V.n7648 VSS 0.074298f
C5493 ASIG5V.n7650 VSS 0.087753f
C5494 ASIG5V.n7652 VSS 0.309175f
C5495 ASIG5V.n7653 VSS 0.314214f
C5496 ASIG5V.n7655 VSS 0.309175f
C5497 ASIG5V.n7656 VSS 0.314214f
C5498 ASIG5V.n7657 VSS 0.074298f
C5499 ASIG5V.n7660 VSS 0.074298f
C5500 ASIG5V.n7662 VSS 0.087753f
C5501 ASIG5V.n7664 VSS 0.309175f
C5502 ASIG5V.n7666 VSS 0.309175f
C5503 ASIG5V.n7667 VSS 0.314214f
C5504 ASIG5V.n7668 VSS 0.074298f
C5505 ASIG5V.n7671 VSS 0.074298f
C5506 ASIG5V.n7673 VSS 0.087753f
C5507 ASIG5V.n7675 VSS 0.845738f
C5508 ASIG5V.n7677 VSS 0.845738f
C5509 ASIG5V.n7678 VSS 0.314214f
C5510 ASIG5V.n7679 VSS 0.074298f
C5511 ASIG5V.n7682 VSS 0.074298f
C5512 ASIG5V.n7684 VSS 0.087753f
C5513 ASIG5V.n7686 VSS 0.309175f
C5514 ASIG5V.n7688 VSS 0.309175f
C5515 ASIG5V.n7690 VSS 0.074298f
C5516 ASIG5V.n7693 VSS 0.074298f
C5517 ASIG5V.n7695 VSS 0.087753f
C5518 ASIG5V.n7697 VSS 0.309175f
C5519 ASIG5V.n7698 VSS 0.309175f
C5520 ASIG5V.n7700 VSS 0.074298f
C5521 ASIG5V.n7702 VSS 0.087753f
C5522 ASIG5V.n7704 VSS 0.309175f
C5523 ASIG5V.n7705 VSS 0.309175f
C5524 ASIG5V.n7708 VSS 0.074298f
C5525 ASIG5V.n7710 VSS 0.087753f
C5526 ASIG5V.n7712 VSS 0.536863f
C5527 ASIG5V.n7713 VSS 0.314214f
C5528 ASIG5V.n7714 VSS 0.050199f
C5529 ASIG5V.n7715 VSS 0.108961f
C5530 ASIG5V.n7716 VSS 0.0621f
C5531 ASIG5V.n7717 VSS 0.056945f
C5532 ASIG5V.n7718 VSS 0.056945f
C5533 ASIG5V.n7719 VSS 0.056945f
C5534 ASIG5V.n7720 VSS 0.056945f
C5535 ASIG5V.n7721 VSS 0.056945f
C5536 ASIG5V.n7722 VSS 0.056945f
C5537 ASIG5V.n7723 VSS 0.056945f
C5538 ASIG5V.n7724 VSS 0.056945f
C5539 ASIG5V.n7725 VSS 0.056945f
C5540 ASIG5V.n7726 VSS 0.056945f
C5541 ASIG5V.n7727 VSS 0.056945f
C5542 ASIG5V.n7728 VSS 0.056945f
C5543 ASIG5V.n7729 VSS 0.056945f
C5544 ASIG5V.n7730 VSS 0.056945f
C5545 ASIG5V.n7731 VSS 0.056945f
C5546 ASIG5V.n7732 VSS 0.056945f
C5547 ASIG5V.n7733 VSS 0.056945f
C5548 ASIG5V.n7734 VSS 0.056945f
C5549 ASIG5V.n7735 VSS 0.056945f
C5550 ASIG5V.n7736 VSS 0.056945f
C5551 ASIG5V.n7737 VSS 0.056945f
C5552 ASIG5V.n7738 VSS 0.056945f
C5553 ASIG5V.n7739 VSS 0.056945f
C5554 ASIG5V.n7740 VSS 0.056945f
C5555 ASIG5V.n7741 VSS 0.056945f
C5556 ASIG5V.n7742 VSS 0.056945f
C5557 ASIG5V.n7743 VSS 0.056945f
C5558 ASIG5V.n7744 VSS 0.056945f
C5559 ASIG5V.n7745 VSS 0.056945f
C5560 ASIG5V.n7746 VSS 0.056945f
C5561 ASIG5V.n7747 VSS 0.056945f
C5562 ASIG5V.n7748 VSS 0.056945f
C5563 ASIG5V.n7749 VSS 0.056945f
C5564 ASIG5V.n7750 VSS 0.056945f
C5565 ASIG5V.n7751 VSS 0.056945f
C5566 ASIG5V.n7752 VSS 0.056945f
C5567 ASIG5V.n7753 VSS 0.056945f
C5568 ASIG5V.n7754 VSS 0.056945f
C5569 ASIG5V.n7755 VSS 0.056945f
C5570 ASIG5V.n7756 VSS 0.056945f
C5571 ASIG5V.n7757 VSS 0.056945f
C5572 ASIG5V.n7758 VSS 0.056945f
C5573 ASIG5V.n7759 VSS 0.056945f
C5574 ASIG5V.n7760 VSS 0.056945f
C5575 ASIG5V.n7761 VSS 0.056945f
C5576 ASIG5V.n7762 VSS 0.056945f
C5577 ASIG5V.n7763 VSS 0.056945f
C5578 ASIG5V.n7764 VSS 0.056945f
C5579 ASIG5V.n7765 VSS 0.056945f
C5580 ASIG5V.n7766 VSS 0.056945f
C5581 ASIG5V.n7767 VSS 0.056945f
C5582 ASIG5V.n7768 VSS 0.056945f
C5583 ASIG5V.n7769 VSS 0.056945f
C5584 ASIG5V.n7770 VSS 0.056945f
C5585 ASIG5V.n7771 VSS 0.056945f
C5586 ASIG5V.n7772 VSS 0.056945f
C5587 ASIG5V.n7773 VSS 0.056945f
C5588 ASIG5V.n7774 VSS 0.056945f
C5589 ASIG5V.n7775 VSS 0.056945f
C5590 ASIG5V.n7776 VSS 0.056945f
C5591 ASIG5V.n7777 VSS 0.056945f
C5592 ASIG5V.n7778 VSS 0.056945f
C5593 ASIG5V.n7779 VSS 0.056945f
C5594 ASIG5V.n7780 VSS 0.056945f
C5595 ASIG5V.n7781 VSS 0.056945f
C5596 ASIG5V.n7782 VSS 0.056945f
C5597 ASIG5V.n7783 VSS 0.056945f
C5598 ASIG5V.n7784 VSS 0.056945f
C5599 ASIG5V.n7785 VSS 0.056945f
C5600 ASIG5V.n7786 VSS 0.056945f
C5601 ASIG5V.n7787 VSS 0.056945f
C5602 ASIG5V.n7788 VSS 0.056945f
C5603 ASIG5V.n7789 VSS 0.056945f
C5604 ASIG5V.n7790 VSS 0.056945f
C5605 ASIG5V.n7791 VSS 0.056945f
C5606 ASIG5V.n7792 VSS 0.056945f
C5607 ASIG5V.n7793 VSS 0.056945f
C5608 ASIG5V.n7794 VSS 0.056945f
C5609 ASIG5V.n7795 VSS 0.056945f
C5610 ASIG5V.n7796 VSS 0.056945f
C5611 ASIG5V.n7797 VSS 0.056945f
C5612 ASIG5V.n7798 VSS 0.056945f
C5613 ASIG5V.n7799 VSS 0.056945f
C5614 ASIG5V.n7800 VSS 0.056945f
C5615 ASIG5V.n7801 VSS 0.056945f
C5616 ASIG5V.n7802 VSS 0.056945f
C5617 ASIG5V.n7803 VSS 0.056945f
C5618 ASIG5V.n7804 VSS 0.056945f
C5619 ASIG5V.n7805 VSS 0.056945f
C5620 ASIG5V.n7806 VSS 0.056945f
C5621 ASIG5V.n7807 VSS 0.056945f
C5622 ASIG5V.n7808 VSS 0.056945f
C5623 ASIG5V.n7809 VSS 0.056945f
C5624 ASIG5V.n7810 VSS 0.056945f
C5625 ASIG5V.n7811 VSS 0.056945f
C5626 ASIG5V.n7812 VSS 0.056945f
C5627 ASIG5V.n7813 VSS 0.056945f
C5628 ASIG5V.n7814 VSS 0.056945f
C5629 ASIG5V.n7815 VSS 0.056945f
C5630 ASIG5V.n7816 VSS 0.056945f
C5631 ASIG5V.n7817 VSS 0.056945f
C5632 ASIG5V.n7818 VSS 0.056945f
C5633 ASIG5V.n7819 VSS 0.056945f
C5634 ASIG5V.n7820 VSS 0.056945f
C5635 ASIG5V.n7821 VSS 0.056945f
C5636 ASIG5V.n7822 VSS 0.056945f
C5637 ASIG5V.n7823 VSS 0.056945f
C5638 ASIG5V.n7824 VSS 0.056945f
C5639 ASIG5V.n7825 VSS 0.056945f
C5640 ASIG5V.n7826 VSS 0.056945f
C5641 ASIG5V.n7827 VSS 0.056945f
C5642 ASIG5V.n7828 VSS 0.056945f
C5643 ASIG5V.n7829 VSS 0.056945f
C5644 ASIG5V.n7830 VSS 0.056945f
C5645 ASIG5V.n7831 VSS 0.056945f
C5646 ASIG5V.n7832 VSS 0.056945f
C5647 ASIG5V.n7833 VSS 0.056945f
C5648 ASIG5V.n7834 VSS 0.056945f
C5649 ASIG5V.n7835 VSS 0.056945f
C5650 ASIG5V.n7836 VSS 0.056945f
C5651 ASIG5V.n7837 VSS 0.056945f
C5652 ASIG5V.n7838 VSS 0.056945f
C5653 ASIG5V.n7839 VSS 0.056945f
C5654 ASIG5V.n7840 VSS 0.056945f
C5655 ASIG5V.n7841 VSS 0.056945f
C5656 ASIG5V.n7842 VSS 0.056945f
C5657 ASIG5V.n7843 VSS 0.056945f
C5658 ASIG5V.n7844 VSS 0.056945f
C5659 ASIG5V.n7845 VSS 0.056945f
C5660 ASIG5V.n7846 VSS 0.056945f
C5661 ASIG5V.n7847 VSS 0.056945f
C5662 ASIG5V.n7848 VSS 0.056945f
C5663 ASIG5V.n7849 VSS 0.056945f
C5664 ASIG5V.n7850 VSS 0.056945f
C5665 ASIG5V.n7851 VSS 0.056945f
C5666 ASIG5V.n7852 VSS 0.056945f
C5667 ASIG5V.n7853 VSS 0.056945f
C5668 ASIG5V.n7854 VSS 0.056945f
C5669 ASIG5V.n7855 VSS 0.056945f
C5670 ASIG5V.n7856 VSS 0.056945f
C5671 ASIG5V.n7857 VSS 0.056945f
C5672 ASIG5V.n7858 VSS 0.056945f
C5673 ASIG5V.n7859 VSS 0.056945f
C5674 ASIG5V.n7860 VSS 0.056945f
C5675 ASIG5V.n7861 VSS 0.056945f
C5676 ASIG5V.n7862 VSS 0.056945f
C5677 ASIG5V.n7863 VSS 0.056945f
C5678 ASIG5V.n7864 VSS 0.056945f
C5679 ASIG5V.n7865 VSS 0.056945f
C5680 ASIG5V.n7866 VSS 0.056945f
C5681 ASIG5V.n7867 VSS 0.056945f
C5682 ASIG5V.n7868 VSS 0.056945f
C5683 ASIG5V.n7869 VSS 0.056945f
C5684 ASIG5V.n7870 VSS 0.056945f
C5685 ASIG5V.n7871 VSS 0.056945f
C5686 ASIG5V.n7872 VSS 0.056945f
C5687 ASIG5V.n7873 VSS 0.056945f
C5688 ASIG5V.n7874 VSS 0.056945f
C5689 ASIG5V.n7875 VSS 0.056945f
C5690 ASIG5V.n7876 VSS 0.056945f
C5691 ASIG5V.n7877 VSS 0.056945f
C5692 ASIG5V.n7878 VSS 0.056945f
C5693 ASIG5V.n7879 VSS 0.056945f
C5694 ASIG5V.n7880 VSS 0.056945f
C5695 ASIG5V.n7881 VSS 0.056945f
C5696 ASIG5V.n7882 VSS 0.056945f
C5697 ASIG5V.n7883 VSS 0.056945f
C5698 ASIG5V.n7884 VSS 0.056945f
C5699 ASIG5V.n7885 VSS 0.056945f
C5700 ASIG5V.n7886 VSS 0.056945f
C5701 ASIG5V.n7887 VSS 0.056945f
C5702 ASIG5V.n7888 VSS 0.056945f
C5703 ASIG5V.n7889 VSS 0.056945f
C5704 ASIG5V.n7890 VSS 0.056945f
C5705 ASIG5V.n7891 VSS 0.056945f
C5706 ASIG5V.n7892 VSS 0.056945f
C5707 ASIG5V.n7893 VSS 0.056945f
C5708 ASIG5V.n7894 VSS 0.056945f
C5709 ASIG5V.n7895 VSS 0.056945f
C5710 ASIG5V.n7896 VSS 0.056945f
C5711 ASIG5V.n7897 VSS 0.056945f
C5712 ASIG5V.n7898 VSS 0.056945f
C5713 ASIG5V.n7899 VSS 0.056945f
C5714 ASIG5V.n7900 VSS 0.056945f
C5715 ASIG5V.n7901 VSS 0.056945f
C5716 ASIG5V.n7902 VSS 0.056945f
C5717 ASIG5V.n7903 VSS 0.056945f
C5718 ASIG5V.n7904 VSS 0.056945f
C5719 ASIG5V.n7905 VSS 0.056945f
C5720 ASIG5V.n7906 VSS 0.056945f
C5721 ASIG5V.n7907 VSS 0.056945f
C5722 ASIG5V.n7908 VSS 0.056945f
C5723 ASIG5V.n7909 VSS 0.056945f
C5724 ASIG5V.n7910 VSS 0.056945f
C5725 ASIG5V.n7911 VSS 0.056945f
C5726 ASIG5V.n7912 VSS 0.056945f
C5727 ASIG5V.n7913 VSS 0.056945f
C5728 ASIG5V.n7914 VSS 0.056945f
C5729 ASIG5V.n7915 VSS 0.056945f
C5730 ASIG5V.n7916 VSS 0.056945f
C5731 ASIG5V.n7917 VSS 0.056945f
C5732 ASIG5V.n7918 VSS 0.056945f
C5733 ASIG5V.n7919 VSS 0.056945f
C5734 ASIG5V.n7920 VSS 0.056945f
C5735 ASIG5V.n7921 VSS 0.056945f
C5736 ASIG5V.n7922 VSS 0.056945f
C5737 ASIG5V.n7923 VSS 0.056945f
C5738 ASIG5V.n7924 VSS 0.056945f
C5739 ASIG5V.n7925 VSS 0.056945f
C5740 ASIG5V.n7926 VSS 0.056945f
C5741 ASIG5V.n7927 VSS 0.056945f
C5742 ASIG5V.n7928 VSS 0.056945f
C5743 ASIG5V.n7929 VSS 0.056945f
C5744 ASIG5V.n7930 VSS 0.056945f
C5745 ASIG5V.n7931 VSS 0.056945f
C5746 ASIG5V.n7932 VSS 0.056945f
C5747 ASIG5V.n7933 VSS 0.056945f
C5748 ASIG5V.n7934 VSS 0.056945f
C5749 ASIG5V.n7935 VSS 0.056945f
C5750 ASIG5V.n7936 VSS 0.056945f
C5751 ASIG5V.n7937 VSS 0.056945f
C5752 ASIG5V.n7938 VSS 0.056945f
C5753 ASIG5V.n7939 VSS 0.056945f
C5754 ASIG5V.n7940 VSS 0.056945f
C5755 ASIG5V.n7941 VSS 0.056945f
C5756 ASIG5V.n7942 VSS 0.056945f
C5757 ASIG5V.n7943 VSS 0.056945f
C5758 ASIG5V.n7944 VSS 0.056945f
C5759 ASIG5V.n7945 VSS 0.056945f
C5760 ASIG5V.n7946 VSS 0.056945f
C5761 ASIG5V.n7947 VSS 0.056945f
C5762 ASIG5V.n7948 VSS 0.056945f
C5763 ASIG5V.n7949 VSS 0.056945f
C5764 ASIG5V.n7950 VSS 0.056945f
C5765 ASIG5V.n7951 VSS 0.056945f
C5766 ASIG5V.n7952 VSS 0.056945f
C5767 ASIG5V.n7953 VSS 0.056945f
C5768 ASIG5V.n7954 VSS 0.056945f
C5769 ASIG5V.n7955 VSS 0.056945f
C5770 ASIG5V.n7956 VSS 0.056945f
C5771 ASIG5V.n7957 VSS 0.056945f
C5772 ASIG5V.n7958 VSS 0.056945f
C5773 ASIG5V.n7959 VSS 0.056945f
C5774 ASIG5V.n7960 VSS 0.052133f
C5775 ASIG5V.n7961 VSS 0.09726f
C5776 ASIG5V.n7962 VSS 0.108961f
C5777 ASIG5V.n7963 VSS 1.07099f
C5778 ASIG5V.n7964 VSS 0.086279f
C5779 ASIG5V.n7965 VSS 0.096659f
C5780 ASIG5V.n7966 VSS 0.096659f
C5781 ASIG5V.n7967 VSS 0.108961f
C5782 ASIG5V.n7968 VSS 0.079084f
C5783 ASIG5V.n7969 VSS 0.079084f
C5784 ASIG5V.n7970 VSS 0.070592f
C5785 ASIG5V.n7971 VSS 0.07229f
C5786 ASIG5V.n7972 VSS 0.075298f
C5787 ASIG5V.n7973 VSS 0.084357f
C5788 ASIG5V.n7974 VSS 0.084357f
C5789 ASIG5V.n7975 VSS 0.108961f
C5790 ASIG5V.n7976 VSS 1.0941f
C5791 ASIG5V.n7977 VSS 0.955415f
C5792 ASIG5V.n7978 VSS 0.654922f
C5793 ASIG5V.n7979 VSS 0.091386f
C5794 ASIG5V.n7980 VSS 0.091386f
C5795 ASIG5V.n7981 VSS 0.080004f
C5796 ASIG5V.n7982 VSS 0.548344f
C5797 ASIG5V.n7983 VSS 0.536863f
C5798 ASIG5V.n7985 VSS 0.087753f
C5799 ASIG5V.n7987 VSS 0.087753f
C5800 ASIG5V.n7988 VSS 0.314214f
C5801 ASIG5V.n7989 VSS 0.074298f
C5802 ASIG5V.n7991 VSS 0.314214f
C5803 ASIG5V.n7992 VSS 0.074298f
C5804 ASIG5V.n7994 VSS 0.314214f
C5805 ASIG5V.n7995 VSS 0.309175f
C5806 ASIG5V.n7996 VSS 0.309175f
C5807 ASIG5V.n7998 VSS 0.074298f
C5808 ASIG5V.n8000 VSS 0.087753f
C5809 ASIG5V.n8002 VSS 0.087753f
C5810 ASIG5V.n8003 VSS 0.074298f
C5811 ASIG5V.n8005 VSS 0.314214f
C5812 ASIG5V.n8006 VSS 0.309175f
C5813 ASIG5V.n8007 VSS 0.309175f
C5814 ASIG5V.n8009 VSS 0.074298f
C5815 ASIG5V.n8011 VSS 0.087753f
C5816 ASIG5V.n8013 VSS 0.087753f
C5817 ASIG5V.n8014 VSS 0.074298f
C5818 ASIG5V.n8016 VSS 0.314214f
C5819 ASIG5V.n8017 VSS 0.309175f
C5820 ASIG5V.n8018 VSS 0.309175f
C5821 ASIG5V.n8020 VSS 0.074298f
C5822 ASIG5V.n8022 VSS 0.087753f
C5823 ASIG5V.n8024 VSS 0.087753f
C5824 ASIG5V.n8025 VSS 0.074298f
C5825 ASIG5V.n8027 VSS 0.314214f
C5826 ASIG5V.n8028 VSS 0.845738f
C5827 ASIG5V.n8029 VSS 0.845738f
C5828 ASIG5V.n8031 VSS 0.074298f
C5829 ASIG5V.n8033 VSS 0.087753f
C5830 ASIG5V.n8035 VSS 0.087753f
C5831 ASIG5V.n8036 VSS 0.074298f
C5832 ASIG5V.n8038 VSS 0.314214f
C5833 ASIG5V.n8039 VSS 0.309175f
C5834 ASIG5V.n8040 VSS 0.309175f
C5835 ASIG5V.n8042 VSS 0.074298f
C5836 ASIG5V.n8044 VSS 0.087753f
C5837 ASIG5V.n8046 VSS 0.087753f
C5838 ASIG5V.n8047 VSS 0.074298f
C5839 ASIG5V.n8049 VSS 0.314214f
C5840 ASIG5V.n8050 VSS 0.309175f
C5841 ASIG5V.n8051 VSS 0.309175f
C5842 ASIG5V.n8053 VSS 0.074298f
C5843 ASIG5V.n8056 VSS 0.087753f
C5844 ASIG5V.n8059 VSS 0.087753f
C5845 ASIG5V.n8060 VSS 0.074298f
C5846 ASIG5V.n8062 VSS 0.314214f
C5847 ASIG5V.n8064 VSS 0.087753f
C5848 ASIG5V.n8066 VSS 0.074298f
C5849 ASIG5V.n8068 VSS 0.314214f
C5850 ASIG5V.n8069 VSS 0.074298f
C5851 ASIG5V.n8071 VSS 0.314214f
C5852 ASIG5V.n8073 VSS 0.087753f
C5853 ASIG5V.n8075 VSS 0.074298f
C5854 ASIG5V.n8077 VSS 0.314214f
C5855 ASIG5V.n8078 VSS 0.074298f
C5856 ASIG5V.n8080 VSS 0.250522f
C5857 ASIG5V.t1 VSS 7.07689f
C5858 ASIG5V.n8082 VSS 0.087753f
C5859 ASIG5V.n8084 VSS 0.074298f
C5860 ASIG5V.n8086 VSS 0.250522f
C5861 ASIG5V.n8087 VSS 0.074298f
C5862 ASIG5V.n8089 VSS 0.314214f
C5863 ASIG5V.n8091 VSS 0.087753f
C5864 ASIG5V.n8093 VSS 0.074298f
C5865 ASIG5V.n8095 VSS 0.314214f
C5866 ASIG5V.n8096 VSS 0.074298f
C5867 ASIG5V.n8098 VSS 0.314214f
C5868 ASIG5V.n8100 VSS 0.314214f
C5869 ASIG5V.n8103 VSS 0.074298f
C5870 ASIG5V.n8105 VSS 0.087753f
C5871 ASIG5V.n8107 VSS 0.309175f
C5872 ASIG5V.n8109 VSS 0.309175f
C5873 ASIG5V.n8111 VSS 0.087753f
C5874 ASIG5V.n8114 VSS 0.074298f
C5875 ASIG5V.n8115 VSS 0.314214f
C5876 ASIG5V.n8116 VSS 0.309175f
C5877 ASIG5V.n8117 VSS 0.309175f
C5878 ASIG5V.n8120 VSS 0.074298f
C5879 ASIG5V.n8122 VSS 0.087753f
C5880 ASIG5V.n8124 VSS 0.845738f
C5881 ASIG5V.n8125 VSS 0.314214f
C5882 ASIG5V.n8126 VSS 0.314214f
C5883 ASIG5V.n8127 VSS 0.074298f
C5884 ASIG5V.n8128 VSS 0.314214f
C5885 ASIG5V.n8129 VSS 0.845738f
C5886 ASIG5V.n8130 VSS 0.845738f
C5887 ASIG5V.n8131 VSS 0.314214f
C5888 ASIG5V.n8133 VSS 0.074298f
C5889 ASIG5V.n8135 VSS 0.087753f
C5890 ASIG5V.n8137 VSS 0.309175f
C5891 ASIG5V.n8138 VSS 0.314214f
C5892 ASIG5V.n8139 VSS 0.314214f
C5893 ASIG5V.n8140 VSS 0.074298f
C5894 ASIG5V.n8141 VSS 0.250522f
C5895 ASIG5V.n8142 VSS 0.309175f
C5896 ASIG5V.n8143 VSS 0.309175f
C5897 ASIG5V.n8144 VSS 0.314214f
C5898 ASIG5V.n8146 VSS 0.074298f
C5899 ASIG5V.n8148 VSS 0.087753f
C5900 ASIG5V.n8150 VSS 0.309175f
C5901 ASIG5V.n8151 VSS 0.250522f
C5902 ASIG5V.t5 VSS 7.07689f
C5903 ASIG5V.n8152 VSS 0.250522f
C5904 ASIG5V.n8153 VSS 0.074298f
C5905 ASIG5V.n8154 VSS 0.314214f
C5906 ASIG5V.n8155 VSS 0.309175f
C5907 ASIG5V.n8156 VSS 0.309175f
C5908 ASIG5V.n8157 VSS 0.250522f
C5909 ASIG5V.n8158 VSS 0.074298f
C5910 ASIG5V.n8160 VSS 0.314214f
C5911 ASIG5V.n8161 VSS 0.309175f
C5912 ASIG5V.n8162 VSS 0.309175f
C5913 ASIG5V.n8163 VSS 0.250522f
C5914 ASIG5V.n8164 VSS 0.074298f
C5915 ASIG5V.n8166 VSS 0.314214f
C5916 ASIG5V.n8167 VSS 0.536863f
C5917 ASIG5V.n8168 VSS 0.050199f
C5918 ASIG5V.n8169 VSS 0.056238f
C5919 ASIG5V.n8170 VSS 0.056238f
C5920 ASIG5V.n8171 VSS 0.955415f
C5921 ASIG5V.n8213 VSS 0.608692f
C5922 ASIG5V.n8214 VSS 0.056945f
C5923 ASIG5V.n8215 VSS 0.0621f
C5924 ASIG5V.n8216 VSS 0.036092f
C5925 ASIG5V.n8217 VSS 0.554757f
C5926 ASIG5V.n8259 VSS 0.608692f
C5927 ASIG5V.n8260 VSS 0.045974f
C5928 ASIG5V.n8261 VSS 0.056945f
C5929 ASIG5V.n8262 VSS 0.056945f
C5930 ASIG5V.n8263 VSS 0.047722f
C5931 ASIG5V.n8264 VSS 0.075358f
C5932 ASIG5V.n8265 VSS 0.076709f
C5933 ASIG5V.n8266 VSS 0.039705f
C5934 ASIG5V.n8267 VSS 0.075358f
C5935 ASIG5V.n8268 VSS 1.0941f
C5936 ASIG5V.n8269 VSS 0.639512f
C5937 ASIG5V.n8270 VSS 0.071037f
C5938 ASIG5V.n8271 VSS 0.071037f
C5939 ASIG5V.n8272 VSS 0.062041f
C5940 ASIG5V.n8273 VSS 0.065815f
C5941 ASIG5V.n8274 VSS 0.052746f
C5942 ASIG5V.n8275 VSS 0.076709f
C5943 ASIG5V.n8276 VSS 0.955415f
C5944 ASIG5V.n8277 VSS 1.0941f
C5945 ASIG5V.n8319 VSS 0.056945f
C5946 ASIG5V.n8320 VSS 0.0621f
C5947 ASIG5V.n8321 VSS 0.0621f
C5948 ASIG5V.n8322 VSS 0.09726f
C5949 ASIG5V.n8323 VSS 0.108961f
C5950 ASIG5V.n8324 VSS 0.0621f
C5951 ASIG5V.n8325 VSS 0.056945f
C5952 ASIG5V.n8326 VSS 0.056945f
C5953 ASIG5V.n8327 VSS 0.056945f
C5954 ASIG5V.n8328 VSS 0.056945f
C5955 ASIG5V.n8329 VSS 0.056945f
C5956 ASIG5V.n8330 VSS 0.056945f
C5957 ASIG5V.n8331 VSS 0.056945f
C5958 ASIG5V.n8332 VSS 0.056945f
C5959 ASIG5V.n8333 VSS 0.056945f
C5960 ASIG5V.n8334 VSS 0.056945f
C5961 ASIG5V.n8335 VSS 0.056945f
C5962 ASIG5V.n8336 VSS 0.056945f
C5963 ASIG5V.n8337 VSS 0.056945f
C5964 ASIG5V.n8338 VSS 0.056945f
C5965 ASIG5V.n8339 VSS 0.056945f
C5966 ASIG5V.n8340 VSS 0.056945f
C5967 ASIG5V.n8341 VSS 0.056945f
C5968 ASIG5V.n8342 VSS 0.056945f
C5969 ASIG5V.n8343 VSS 0.056945f
C5970 ASIG5V.n8344 VSS 0.056945f
C5971 ASIG5V.n8345 VSS 0.056945f
C5972 ASIG5V.n8346 VSS 0.056945f
C5973 ASIG5V.n8347 VSS 0.056945f
C5974 ASIG5V.n8348 VSS 0.056945f
C5975 ASIG5V.n8349 VSS 0.056945f
C5976 ASIG5V.n8350 VSS 0.056945f
C5977 ASIG5V.n8351 VSS 0.056945f
C5978 ASIG5V.n8352 VSS 0.056945f
C5979 ASIG5V.n8353 VSS 0.056945f
C5980 ASIG5V.n8354 VSS 0.056945f
C5981 ASIG5V.n8355 VSS 0.056945f
C5982 ASIG5V.n8356 VSS 0.056945f
C5983 ASIG5V.n8357 VSS 0.056945f
C5984 ASIG5V.n8358 VSS 0.056945f
C5985 ASIG5V.n8359 VSS 0.056945f
C5986 ASIG5V.n8360 VSS 0.056945f
C5987 ASIG5V.n8361 VSS 0.056945f
C5988 ASIG5V.n8362 VSS 0.056945f
C5989 ASIG5V.n8363 VSS 0.056945f
C5990 ASIG5V.n8364 VSS 0.056945f
C5991 ASIG5V.n8365 VSS 0.056945f
C5992 ASIG5V.n8366 VSS 0.056945f
C5993 ASIG5V.n8367 VSS 0.056945f
C5994 ASIG5V.n8368 VSS 0.056945f
C5995 ASIG5V.n8369 VSS 0.056945f
C5996 ASIG5V.n8370 VSS 0.056945f
C5997 ASIG5V.n8371 VSS 0.056945f
C5998 ASIG5V.n8372 VSS 0.056945f
C5999 ASIG5V.n8373 VSS 0.056945f
C6000 ASIG5V.n8374 VSS 0.056945f
C6001 ASIG5V.n8375 VSS 0.056945f
C6002 ASIG5V.n8376 VSS 0.056945f
C6003 ASIG5V.n8377 VSS 0.056945f
C6004 ASIG5V.n8378 VSS 0.056945f
C6005 ASIG5V.n8379 VSS 0.056945f
C6006 ASIG5V.n8380 VSS 0.056945f
C6007 ASIG5V.n8381 VSS 0.056945f
C6008 ASIG5V.n8382 VSS 0.056945f
C6009 ASIG5V.n8383 VSS 0.056945f
C6010 ASIG5V.n8384 VSS 0.056945f
C6011 ASIG5V.n8385 VSS 0.056945f
C6012 ASIG5V.n8386 VSS 0.056945f
C6013 ASIG5V.n8387 VSS 0.056945f
C6014 ASIG5V.n8388 VSS 0.056945f
C6015 ASIG5V.n8389 VSS 0.056945f
C6016 ASIG5V.n8390 VSS 0.056945f
C6017 ASIG5V.n8391 VSS 0.056945f
C6018 ASIG5V.n8392 VSS 0.056945f
C6019 ASIG5V.n8393 VSS 0.056945f
C6020 ASIG5V.n8394 VSS 0.056945f
C6021 ASIG5V.n8395 VSS 0.056945f
C6022 ASIG5V.n8396 VSS 0.056945f
C6023 ASIG5V.n8397 VSS 0.056945f
C6024 ASIG5V.n8398 VSS 0.056945f
C6025 ASIG5V.n8399 VSS 0.056945f
C6026 ASIG5V.n8400 VSS 0.056945f
C6027 ASIG5V.n8401 VSS 0.056945f
C6028 ASIG5V.n8402 VSS 0.056945f
C6029 ASIG5V.n8403 VSS 0.056945f
C6030 ASIG5V.n8404 VSS 0.056945f
C6031 ASIG5V.n8405 VSS 0.056945f
C6032 ASIG5V.n8406 VSS 0.056945f
C6033 ASIG5V.n8407 VSS 0.056945f
C6034 ASIG5V.n8408 VSS 0.056945f
C6035 ASIG5V.n8409 VSS 0.056945f
C6036 ASIG5V.n8410 VSS 0.056945f
C6037 ASIG5V.n8411 VSS 0.056945f
C6038 ASIG5V.n8412 VSS 0.056945f
C6039 ASIG5V.n8413 VSS 0.056945f
C6040 ASIG5V.n8414 VSS 0.056945f
C6041 ASIG5V.n8415 VSS 0.056945f
C6042 ASIG5V.n8416 VSS 0.056945f
C6043 ASIG5V.n8417 VSS 0.056945f
C6044 ASIG5V.n8418 VSS 0.056945f
C6045 ASIG5V.n8419 VSS 0.056945f
C6046 ASIG5V.n8420 VSS 0.056945f
C6047 ASIG5V.n8421 VSS 0.056945f
C6048 ASIG5V.n8422 VSS 0.056945f
C6049 ASIG5V.n8423 VSS 0.056945f
C6050 ASIG5V.n8424 VSS 0.056945f
C6051 ASIG5V.n8425 VSS 0.056945f
C6052 ASIG5V.n8426 VSS 0.056945f
C6053 ASIG5V.n8427 VSS 0.056945f
C6054 ASIG5V.n8428 VSS 0.056945f
C6055 ASIG5V.n8429 VSS 0.056945f
C6056 ASIG5V.n8430 VSS 0.056945f
C6057 ASIG5V.n8431 VSS 0.056945f
C6058 ASIG5V.n8432 VSS 0.056945f
C6059 ASIG5V.n8433 VSS 0.056945f
C6060 ASIG5V.n8434 VSS 0.056945f
C6061 ASIG5V.n8435 VSS 0.056945f
C6062 ASIG5V.n8436 VSS 0.056945f
C6063 ASIG5V.n8437 VSS 0.056945f
C6064 ASIG5V.n8438 VSS 0.056945f
C6065 ASIG5V.n8439 VSS 0.056945f
C6066 ASIG5V.n8440 VSS 0.056945f
C6067 ASIG5V.n8441 VSS 0.056945f
C6068 ASIG5V.n8442 VSS 0.056945f
C6069 ASIG5V.n8443 VSS 0.056945f
C6070 ASIG5V.n8444 VSS 0.056945f
C6071 ASIG5V.n8445 VSS 0.056945f
C6072 ASIG5V.n8446 VSS 0.056945f
C6073 ASIG5V.n8447 VSS 0.056945f
C6074 ASIG5V.n8448 VSS 0.056945f
C6075 ASIG5V.n8449 VSS 0.056945f
C6076 ASIG5V.n8450 VSS 0.056945f
C6077 ASIG5V.n8451 VSS 0.056945f
C6078 ASIG5V.n8452 VSS 0.056945f
C6079 ASIG5V.n8453 VSS 0.056945f
C6080 ASIG5V.n8454 VSS 0.056945f
C6081 ASIG5V.n8455 VSS 0.056945f
C6082 ASIG5V.n8456 VSS 0.056945f
C6083 ASIG5V.n8457 VSS 0.056945f
C6084 ASIG5V.n8458 VSS 0.056945f
C6085 ASIG5V.n8459 VSS 0.056945f
C6086 ASIG5V.n8460 VSS 0.056945f
C6087 ASIG5V.n8461 VSS 0.056945f
C6088 ASIG5V.n8462 VSS 0.056945f
C6089 ASIG5V.n8463 VSS 0.056945f
C6090 ASIG5V.n8464 VSS 0.056945f
C6091 ASIG5V.n8465 VSS 0.056945f
C6092 ASIG5V.n8466 VSS 0.056945f
C6093 ASIG5V.n8467 VSS 0.056945f
C6094 ASIG5V.n8468 VSS 0.056945f
C6095 ASIG5V.n8469 VSS 0.056945f
C6096 ASIG5V.n8470 VSS 0.056945f
C6097 ASIG5V.n8471 VSS 0.056945f
C6098 ASIG5V.n8472 VSS 0.056945f
C6099 ASIG5V.n8473 VSS 0.056945f
C6100 ASIG5V.n8474 VSS 0.056945f
C6101 ASIG5V.n8475 VSS 0.056945f
C6102 ASIG5V.n8476 VSS 0.056945f
C6103 ASIG5V.n8477 VSS 0.056945f
C6104 ASIG5V.n8478 VSS 0.056945f
C6105 ASIG5V.n8479 VSS 0.056945f
C6106 ASIG5V.n8480 VSS 0.056945f
C6107 ASIG5V.n8481 VSS 0.056945f
C6108 ASIG5V.n8482 VSS 0.056945f
C6109 ASIG5V.n8483 VSS 0.056945f
C6110 ASIG5V.n8484 VSS 0.056945f
C6111 ASIG5V.n8485 VSS 0.056945f
C6112 ASIG5V.n8486 VSS 0.056945f
C6113 ASIG5V.n8487 VSS 0.056945f
C6114 ASIG5V.n8488 VSS 0.056945f
C6115 ASIG5V.n8489 VSS 0.056945f
C6116 ASIG5V.n8490 VSS 0.056945f
C6117 ASIG5V.n8491 VSS 0.056945f
C6118 ASIG5V.n8492 VSS 0.056945f
C6119 ASIG5V.n8493 VSS 0.056945f
C6120 ASIG5V.n8494 VSS 0.056945f
C6121 ASIG5V.n8495 VSS 0.056945f
C6122 ASIG5V.n8496 VSS 0.056945f
C6123 ASIG5V.n8497 VSS 0.056945f
C6124 ASIG5V.n8498 VSS 0.056945f
C6125 ASIG5V.n8499 VSS 0.056945f
C6126 ASIG5V.n8500 VSS 0.056945f
C6127 ASIG5V.n8501 VSS 0.056945f
C6128 ASIG5V.n8502 VSS 0.056945f
C6129 ASIG5V.n8503 VSS 0.056945f
C6130 ASIG5V.n8504 VSS 0.056945f
C6131 ASIG5V.n8505 VSS 0.056945f
C6132 ASIG5V.n8506 VSS 0.056945f
C6133 ASIG5V.n8507 VSS 0.056945f
C6134 ASIG5V.n8508 VSS 0.056945f
C6135 ASIG5V.n8509 VSS 0.056945f
C6136 ASIG5V.n8510 VSS 0.056945f
C6137 ASIG5V.n8511 VSS 0.056945f
C6138 ASIG5V.n8512 VSS 0.056945f
C6139 ASIG5V.n8513 VSS 0.056945f
C6140 ASIG5V.n8514 VSS 0.056945f
C6141 ASIG5V.n8515 VSS 0.056945f
C6142 ASIG5V.n8516 VSS 0.056945f
C6143 ASIG5V.n8517 VSS 0.056945f
C6144 ASIG5V.n8518 VSS 0.056945f
C6145 ASIG5V.n8519 VSS 0.056945f
C6146 ASIG5V.n8520 VSS 0.056945f
C6147 ASIG5V.n8521 VSS 0.056945f
C6148 ASIG5V.n8522 VSS 0.056945f
C6149 ASIG5V.n8523 VSS 0.056945f
C6150 ASIG5V.n8524 VSS 0.056945f
C6151 ASIG5V.n8525 VSS 0.056945f
C6152 ASIG5V.n8526 VSS 0.056945f
C6153 ASIG5V.n8527 VSS 0.056945f
C6154 ASIG5V.n8528 VSS 0.056945f
C6155 ASIG5V.n8529 VSS 0.056945f
C6156 ASIG5V.n8530 VSS 0.056945f
C6157 ASIG5V.n8531 VSS 0.056945f
C6158 ASIG5V.n8532 VSS 0.056945f
C6159 ASIG5V.n8533 VSS 0.056945f
C6160 ASIG5V.n8534 VSS 0.056945f
C6161 ASIG5V.n8535 VSS 0.056945f
C6162 ASIG5V.n8536 VSS 0.056945f
C6163 ASIG5V.n8537 VSS 0.056945f
C6164 ASIG5V.n8538 VSS 0.056945f
C6165 ASIG5V.n8539 VSS 0.056945f
C6166 ASIG5V.n8540 VSS 0.056945f
C6167 ASIG5V.n8541 VSS 0.056945f
C6168 ASIG5V.n8542 VSS 0.056945f
C6169 ASIG5V.n8543 VSS 0.056945f
C6170 ASIG5V.n8544 VSS 0.056945f
C6171 ASIG5V.n8545 VSS 0.056945f
C6172 ASIG5V.n8546 VSS 0.056945f
C6173 ASIG5V.n8547 VSS 0.056945f
C6174 ASIG5V.n8548 VSS 0.056945f
C6175 ASIG5V.n8549 VSS 0.056945f
C6176 ASIG5V.n8550 VSS 0.056945f
C6177 ASIG5V.n8551 VSS 0.056945f
C6178 ASIG5V.n8552 VSS 0.056945f
C6179 ASIG5V.n8553 VSS 0.056945f
C6180 ASIG5V.n8554 VSS 0.056945f
C6181 ASIG5V.n8555 VSS 0.056945f
C6182 ASIG5V.n8556 VSS 0.056945f
C6183 ASIG5V.n8557 VSS 0.056945f
C6184 ASIG5V.n8558 VSS 0.056945f
C6185 ASIG5V.n8559 VSS 0.056945f
C6186 ASIG5V.n8560 VSS 0.056945f
C6187 ASIG5V.n8561 VSS 0.056945f
C6188 ASIG5V.n8562 VSS 0.056945f
C6189 ASIG5V.n8563 VSS 0.056945f
C6190 ASIG5V.n8564 VSS 0.056945f
C6191 ASIG5V.n8565 VSS 0.056945f
C6192 ASIG5V.n8566 VSS 0.056945f
C6193 ASIG5V.n8567 VSS 0.056945f
C6194 ASIG5V.n8568 VSS 0.052133f
C6195 ASIG5V.n8569 VSS 0.07229f
C6196 ASIG5V.n8570 VSS 0.095691f
C6197 ASIG5V.n8571 VSS 0.107203f
C6198 ASIG5V.n8572 VSS 0.107203f
C6199 ASIG5V.n8573 VSS 0.108961f
C6200 ASIG5V.n8574 VSS 0.06854f
C6201 ASIG5V.n8575 VSS 0.06854f
C6202 ASIG5V.n8576 VSS 0.06118f
C6203 ASIG5V.n8577 VSS 0.09726f
C6204 ASIG5V.n8578 VSS 0.108961f
C6205 ASIG5V.n8579 VSS 0.080842f
C6206 ASIG5V.n8580 VSS 0.080842f
C6207 ASIG5V.n8581 VSS 0.108961f
C6208 ASIG5V.n8582 VSS 0.955415f
C6209 ASIG5V.n8583 VSS 0.793611f
C6210 ASIG5V.n8584 VSS 0.094901f
C6211 ASIG5V.n8585 VSS 0.094901f
C6212 ASIG5V.n8586 VSS 0.08471f
C6213 ASIG5V.n8587 VSS 0.07229f
C6214 ASIG5V.n8588 VSS 0.052133f
C6215 ASIG5V.n8590 VSS 0.056945f
C6216 ASIG5V.n8591 VSS 0.056945f
C6217 ASIG5V.n8592 VSS 0.056945f
C6218 ASIG5V.n8593 VSS 0.056945f
C6219 ASIG5V.n8594 VSS 0.056945f
C6220 ASIG5V.n8595 VSS 0.056945f
C6221 ASIG5V.n8596 VSS 0.056945f
C6222 ASIG5V.n8597 VSS 0.056945f
C6223 ASIG5V.n8598 VSS 0.056945f
C6224 ASIG5V.n8599 VSS 0.056945f
C6225 ASIG5V.n8600 VSS 0.056945f
C6226 ASIG5V.n8601 VSS 0.056945f
C6227 ASIG5V.n8602 VSS 0.056945f
C6228 ASIG5V.n8603 VSS 0.056945f
C6229 ASIG5V.n8604 VSS 0.056945f
C6230 ASIG5V.n8605 VSS 0.056945f
C6231 ASIG5V.n8606 VSS 0.056945f
C6232 ASIG5V.n8607 VSS 0.056945f
C6233 ASIG5V.n8608 VSS 0.056945f
C6234 ASIG5V.n8609 VSS 0.056945f
C6235 ASIG5V.n8610 VSS 0.056945f
C6236 ASIG5V.n8611 VSS 0.056945f
C6237 ASIG5V.n8612 VSS 0.056945f
C6238 ASIG5V.n8613 VSS 0.056945f
C6239 ASIG5V.n8614 VSS 0.056945f
C6240 ASIG5V.n8615 VSS 0.056945f
C6241 ASIG5V.n8616 VSS 0.056945f
C6242 ASIG5V.n8617 VSS 0.056945f
C6243 ASIG5V.n8618 VSS 0.056945f
C6244 ASIG5V.n8619 VSS 0.056945f
C6245 ASIG5V.n8620 VSS 0.056945f
C6246 ASIG5V.n8621 VSS 0.056945f
C6247 ASIG5V.n8622 VSS 0.056945f
C6248 ASIG5V.n8623 VSS 0.056945f
C6249 ASIG5V.n8624 VSS 0.056945f
C6250 ASIG5V.n8625 VSS 0.056945f
C6251 ASIG5V.n8626 VSS 0.056945f
C6252 ASIG5V.n8627 VSS 0.056945f
C6253 ASIG5V.n8628 VSS 0.056945f
C6254 ASIG5V.n8629 VSS 0.056945f
C6255 ASIG5V.n8630 VSS 0.056945f
C6256 ASIG5V.n8631 VSS 0.056945f
C6257 ASIG5V.n8632 VSS 0.036092f
C6258 ASIG5V.n8633 VSS 0.036092f
C6259 ASIG5V.n8634 VSS 0.047722f
C6260 ASIG5V.n8635 VSS 0.056945f
C6261 ASIG5V.n8636 VSS 0.056945f
C6262 ASIG5V.n8637 VSS 0.056945f
C6263 ASIG5V.n8639 VSS 0.056945f
C6264 ASIG5V.n8640 VSS 0.056945f
C6265 ASIG5V.n8641 VSS 0.056945f
C6266 ASIG5V.n8642 VSS 0.056945f
C6267 ASIG5V.n8644 VSS 0.056945f
C6268 ASIG5V.n8645 VSS 0.056945f
C6269 ASIG5V.n8646 VSS 0.056945f
C6270 ASIG5V.n8647 VSS 0.056945f
C6271 ASIG5V.n8648 VSS 0.056945f
C6272 ASIG5V.n8649 VSS 0.056945f
C6273 ASIG5V.n8651 VSS 0.056945f
C6274 ASIG5V.n8652 VSS 0.056945f
C6275 ASIG5V.n8653 VSS 0.056945f
C6276 ASIG5V.n8654 VSS 0.056945f
C6277 ASIG5V.n8656 VSS 0.056945f
C6278 ASIG5V.n8657 VSS 0.056945f
C6279 ASIG5V.n8658 VSS 0.056945f
C6280 ASIG5V.n8659 VSS 0.056945f
C6281 ASIG5V.n8660 VSS 0.056945f
C6282 ASIG5V.n8661 VSS 0.056945f
C6283 ASIG5V.n8663 VSS 0.056945f
C6284 ASIG5V.n8664 VSS 0.056945f
C6285 ASIG5V.n8665 VSS 0.056945f
C6286 ASIG5V.n8666 VSS 0.056945f
C6287 ASIG5V.n8668 VSS 0.056945f
C6288 ASIG5V.n8669 VSS 0.056945f
C6289 ASIG5V.n8670 VSS 0.056945f
C6290 ASIG5V.n8671 VSS 0.056945f
C6291 ASIG5V.n8672 VSS 0.056945f
C6292 ASIG5V.n8673 VSS 0.056945f
C6293 ASIG5V.n8675 VSS 0.056945f
C6294 ASIG5V.n8676 VSS 0.056945f
C6295 ASIG5V.n8677 VSS 0.056945f
C6296 ASIG5V.n8678 VSS 0.056945f
C6297 ASIG5V.n8680 VSS 0.056945f
C6298 ASIG5V.n8681 VSS 0.056945f
C6299 ASIG5V.n8682 VSS 0.056945f
C6300 ASIG5V.n8683 VSS 0.056945f
C6301 ASIG5V.n8684 VSS 0.056945f
C6302 ASIG5V.n8685 VSS 0.056945f
C6303 ASIG5V.n8687 VSS 0.056945f
C6304 ASIG5V.n8688 VSS 0.056945f
C6305 ASIG5V.n8689 VSS 0.056945f
C6306 ASIG5V.n8690 VSS 0.056945f
C6307 ASIG5V.n8692 VSS 0.056945f
C6308 ASIG5V.n8693 VSS 0.056945f
C6309 ASIG5V.n8694 VSS 0.056945f
C6310 ASIG5V.n8695 VSS 0.056945f
C6311 ASIG5V.n8696 VSS 0.056945f
C6312 ASIG5V.n8697 VSS 0.056945f
C6313 ASIG5V.n8699 VSS 0.056945f
C6314 ASIG5V.n8700 VSS 0.056945f
C6315 ASIG5V.n8701 VSS 0.056945f
C6316 ASIG5V.n8702 VSS 0.056945f
C6317 ASIG5V.n8704 VSS 0.056945f
C6318 ASIG5V.n8705 VSS 0.056945f
C6319 ASIG5V.n8706 VSS 0.056945f
C6320 ASIG5V.n8707 VSS 0.056945f
C6321 ASIG5V.n8708 VSS 0.056945f
C6322 ASIG5V.n8709 VSS 0.056945f
C6323 ASIG5V.n8711 VSS 0.056945f
C6324 ASIG5V.n8712 VSS 0.056945f
C6325 ASIG5V.n8713 VSS 0.056945f
C6326 ASIG5V.n8714 VSS 0.056945f
C6327 ASIG5V.n8716 VSS 0.056945f
C6328 ASIG5V.n8717 VSS 0.056945f
C6329 ASIG5V.n8718 VSS 0.056945f
C6330 ASIG5V.n8719 VSS 0.056945f
C6331 ASIG5V.n8720 VSS 0.056945f
C6332 ASIG5V.n8721 VSS 0.056945f
C6333 ASIG5V.n8723 VSS 0.056945f
C6334 ASIG5V.n8724 VSS 0.056945f
C6335 ASIG5V.n8725 VSS 0.056945f
C6336 ASIG5V.n8726 VSS 0.056945f
C6337 ASIG5V.n8728 VSS 0.056945f
C6338 ASIG5V.n8729 VSS 0.056945f
C6339 ASIG5V.n8730 VSS 0.056945f
C6340 ASIG5V.n8731 VSS 0.056945f
C6341 ASIG5V.n8732 VSS 0.056945f
C6342 ASIG5V.n8733 VSS 0.056945f
C6343 ASIG5V.n8735 VSS 0.056945f
C6344 ASIG5V.n8736 VSS 0.056945f
C6345 ASIG5V.n8737 VSS 0.056945f
C6346 ASIG5V.n8738 VSS 0.056945f
C6347 ASIG5V.n8740 VSS 0.056945f
C6348 ASIG5V.n8741 VSS 0.056945f
C6349 ASIG5V.n8742 VSS 0.056945f
C6350 ASIG5V.n8743 VSS 0.056945f
C6351 ASIG5V.n8744 VSS 0.056945f
C6352 ASIG5V.n8745 VSS 0.056945f
C6353 ASIG5V.n8747 VSS 0.056945f
C6354 ASIG5V.n8748 VSS 0.056945f
C6355 ASIG5V.n8749 VSS 0.056945f
C6356 ASIG5V.n8750 VSS 0.056945f
C6357 ASIG5V.n8752 VSS 0.056945f
C6358 ASIG5V.n8753 VSS 0.056945f
C6359 ASIG5V.n8754 VSS 0.056945f
C6360 ASIG5V.n8755 VSS 0.056945f
C6361 ASIG5V.n8756 VSS 0.056945f
C6362 ASIG5V.n8757 VSS 0.056945f
C6363 ASIG5V.n8759 VSS 0.056945f
C6364 ASIG5V.n8760 VSS 0.056945f
C6365 ASIG5V.n8761 VSS 0.056945f
C6366 ASIG5V.n8762 VSS 0.056945f
C6367 ASIG5V.n8764 VSS 0.056945f
C6368 ASIG5V.n8765 VSS 0.056945f
C6369 ASIG5V.n8766 VSS 0.056945f
C6370 ASIG5V.n8767 VSS 0.056945f
C6371 ASIG5V.n8768 VSS 0.056945f
C6372 ASIG5V.n8769 VSS 0.056945f
C6373 ASIG5V.n8771 VSS 0.056945f
C6374 ASIG5V.n8772 VSS 0.056945f
C6375 ASIG5V.n8773 VSS 0.056945f
C6376 ASIG5V.n8774 VSS 0.056945f
C6377 ASIG5V.n8776 VSS 0.056945f
C6378 ASIG5V.n8777 VSS 0.056945f
C6379 ASIG5V.n8778 VSS 0.056945f
C6380 ASIG5V.n8779 VSS 0.056945f
C6381 ASIG5V.n8780 VSS 0.056945f
C6382 ASIG5V.n8781 VSS 0.056945f
C6383 ASIG5V.n8783 VSS 0.056945f
C6384 ASIG5V.n8784 VSS 0.056945f
C6385 ASIG5V.n8785 VSS 0.056945f
C6386 ASIG5V.n8786 VSS 0.056945f
C6387 ASIG5V.n8788 VSS 0.056945f
C6388 ASIG5V.n8789 VSS 0.056945f
C6389 ASIG5V.n8790 VSS 0.056945f
C6390 ASIG5V.n8791 VSS 0.056945f
C6391 ASIG5V.n8792 VSS 0.056945f
C6392 ASIG5V.n8793 VSS 0.056945f
C6393 ASIG5V.n8795 VSS 0.056945f
C6394 ASIG5V.n8796 VSS 0.056945f
C6395 ASIG5V.n8797 VSS 0.056945f
C6396 ASIG5V.n8798 VSS 0.056945f
C6397 ASIG5V.n8800 VSS 0.056945f
C6398 ASIG5V.n8801 VSS 0.056945f
C6399 ASIG5V.n8802 VSS 0.056945f
C6400 ASIG5V.n8803 VSS 0.056945f
C6401 ASIG5V.n8804 VSS 0.056945f
C6402 ASIG5V.n8805 VSS 0.056945f
C6403 ASIG5V.n8807 VSS 0.056945f
C6404 ASIG5V.n8808 VSS 0.056945f
C6405 ASIG5V.n8809 VSS 0.056945f
C6406 ASIG5V.n8810 VSS 0.056945f
C6407 ASIG5V.n8812 VSS 0.056945f
C6408 ASIG5V.n8813 VSS 0.056945f
C6409 ASIG5V.n8814 VSS 0.056945f
C6410 ASIG5V.n8815 VSS 0.056945f
C6411 ASIG5V.n8816 VSS 0.056945f
C6412 ASIG5V.n8817 VSS 0.056945f
C6413 ASIG5V.n8819 VSS 0.056945f
C6414 ASIG5V.n8820 VSS 0.056945f
C6415 ASIG5V.n8821 VSS 0.056945f
C6416 ASIG5V.n8822 VSS 0.056945f
C6417 ASIG5V.n8824 VSS 0.056945f
C6418 ASIG5V.n8825 VSS 0.056945f
C6419 ASIG5V.n8826 VSS 0.056945f
C6420 ASIG5V.n8827 VSS 0.056945f
C6421 ASIG5V.n8828 VSS 0.056945f
C6422 ASIG5V.n8829 VSS 0.056945f
C6423 ASIG5V.n8831 VSS 0.056945f
C6424 ASIG5V.n8832 VSS 0.056945f
C6425 ASIG5V.n8833 VSS 0.056945f
C6426 ASIG5V.n8834 VSS 0.056945f
C6427 ASIG5V.n8836 VSS 0.056945f
C6428 ASIG5V.n8837 VSS 0.056945f
C6429 ASIG5V.n8838 VSS 0.056945f
C6430 ASIG5V.n8839 VSS 0.056945f
C6431 ASIG5V.n8840 VSS 0.056945f
C6432 ASIG5V.n8841 VSS 0.056945f
C6433 ASIG5V.n8843 VSS 0.056945f
C6434 ASIG5V.n8844 VSS 0.056945f
C6435 ASIG5V.n8845 VSS 0.056945f
C6436 ASIG5V.n8846 VSS 0.056945f
C6437 ASIG5V.n8848 VSS 0.056945f
C6438 ASIG5V.n8849 VSS 0.056945f
C6439 ASIG5V.n8850 VSS 0.056945f
C6440 ASIG5V.n8851 VSS 0.056945f
C6441 ASIG5V.n8852 VSS 0.056945f
C6442 ASIG5V.n8853 VSS 0.056945f
C6443 ASIG5V.n8855 VSS 0.056945f
C6444 ASIG5V.n8856 VSS 0.056945f
C6445 ASIG5V.n8857 VSS 0.056945f
C6446 ASIG5V.n8858 VSS 0.056945f
C6447 ASIG5V.n8860 VSS 0.056945f
C6448 ASIG5V.n8861 VSS 0.056945f
C6449 ASIG5V.n8862 VSS 0.056945f
C6450 ASIG5V.n8863 VSS 0.056945f
C6451 ASIG5V.n8864 VSS 0.056945f
C6452 ASIG5V.n8865 VSS 0.056945f
C6453 ASIG5V.n8867 VSS 0.056945f
C6454 ASIG5V.n8868 VSS 0.056945f
C6455 ASIG5V.n8869 VSS 0.056945f
C6456 ASIG5V.n8870 VSS 0.056945f
C6457 ASIG5V.n8872 VSS 0.056945f
C6458 ASIG5V.n8873 VSS 0.056945f
C6459 ASIG5V.n8874 VSS 0.056945f
C6460 ASIG5V.n8875 VSS 0.056945f
C6461 ASIG5V.n8876 VSS 0.056945f
C6462 ASIG5V.n8877 VSS 0.056945f
C6463 ASIG5V.n8878 VSS 0.036092f
C6464 ASIG5V.n8879 VSS 0.036092f
C6465 ASIG5V.n8881 VSS 0.608692f
C6466 ASIG5V.n8882 VSS 0.647216f
C6467 ASIG5V.n8883 VSS 0.068336f
C6468 ASIG5V.n8884 VSS 0.068336f
C6469 ASIG5V.n8885 VSS 0.059682f
C6470 ASIG5V.n8886 VSS 0.066995f
C6471 ASIG5V.n8887 VSS 0.034677f
C6472 ASIG5V.n8888 VSS 0.039705f
C6473 ASIG5V.n8889 VSS 0.045974f
C6474 ASIG5V.n8890 VSS 0.036092f
C6475 ASIG5V.n8891 VSS 0.036092f
C6476 ASIG5V.n8892 VSS 0.886071f
C6477 ASIG5V.n8893 VSS 0.036092f
C6478 ASIG5V.n8895 VSS 0.955416f
C6479 ASIG5V.n8896 VSS 0.485412f
C6480 ASIG5V.n8897 VSS 0.108961f
C6481 ASIG5V.n8898 VSS 0.108961f
C6482 ASIG5V.n8899 VSS 0.09726f
C6483 ASIG5V.n8900 VSS 0.080004f
C6484 ASIG5V.n8901 VSS 0.548344f
C6485 ASIG5V.n8902 VSS 0.026668f
C6486 ASIG5V.n8903 VSS 0.065025f
C6487 ASIG5V.n8904 VSS 0.065025f
C6488 ASIG5V.n8905 VSS 0.662626f
C6489 ASIG5V.n8906 VSS 0.778201f
C6490 ASIG5V.n8907 VSS 0.044026f
C6491 ASIG5V.n8908 VSS 0.044026f
C6492 ASIG5V.n8909 VSS 0.038451f
C6493 ASIG5V.n8910 VSS 0.066995f
C6494 ASIG5V.n8911 VSS 0.055908f
C6495 ASIG5V.n8912 VSS 0.064014f
C6496 ASIG5V.n8913 VSS 0.045974f
C6497 ASIG5V.n8914 VSS 0.036092f
C6498 ASIG5V.n8915 VSS 0.036092f
C6499 ASIG5V.n8916 VSS 0.331313f
C6500 ASIG5V.n8917 VSS 0.036092f
C6501 ASIG5V.n8919 VSS 0.192624f
C6502 ASIG5V.n8920 VSS 0.909185f
C6503 ASIG5V.n8921 VSS 0.086114f
C6504 ASIG5V.n8922 VSS 0.086114f
C6505 ASIG5V.n8923 VSS 0.076867f
C6506 ASIG5V.n8924 VSS 0.09726f
C6507 ASIG5V.n8925 VSS 0.080004f
C6508 ASIG5V.n8926 VSS 0.089629f
C6509 ASIG5V.n8927 VSS 0.0621f
C6510 ASIG5V.n8928 VSS 0.036092f
C6511 ASIG5V.n8929 VSS 0.052133f
C6512 ASIG5V.n8930 VSS 0.056945f
C6513 ASIG5V.n8931 VSS 0.056945f
C6514 ASIG5V.n8932 VSS 0.056945f
C6515 ASIG5V.n8933 VSS 0.056945f
C6516 ASIG5V.n8935 VSS 0.056945f
C6517 ASIG5V.n8936 VSS 0.056945f
C6518 ASIG5V.n8937 VSS 0.056945f
C6519 ASIG5V.n8939 VSS 0.056945f
C6520 ASIG5V.n8940 VSS 0.056945f
C6521 ASIG5V.n8941 VSS 0.056945f
C6522 ASIG5V.n8942 VSS 0.056945f
C6523 ASIG5V.n8943 VSS 0.056945f
C6524 ASIG5V.n8944 VSS 0.056945f
C6525 ASIG5V.n8945 VSS 0.056945f
C6526 ASIG5V.n8947 VSS 0.056945f
C6527 ASIG5V.n8948 VSS 0.056945f
C6528 ASIG5V.n8949 VSS 0.056945f
C6529 ASIG5V.n8951 VSS 0.056945f
C6530 ASIG5V.n8952 VSS 0.056945f
C6531 ASIG5V.n8953 VSS 0.056945f
C6532 ASIG5V.n8954 VSS 0.056945f
C6533 ASIG5V.n8955 VSS 0.056945f
C6534 ASIG5V.n8956 VSS 0.056945f
C6535 ASIG5V.n8957 VSS 0.056945f
C6536 ASIG5V.n8959 VSS 0.056945f
C6537 ASIG5V.n8960 VSS 0.056945f
C6538 ASIG5V.n8961 VSS 0.056945f
C6539 ASIG5V.n8963 VSS 0.056945f
C6540 ASIG5V.n8964 VSS 0.056945f
C6541 ASIG5V.n8965 VSS 0.056945f
C6542 ASIG5V.n8966 VSS 0.056945f
C6543 ASIG5V.n8967 VSS 0.056945f
C6544 ASIG5V.n8968 VSS 0.056945f
C6545 ASIG5V.n8969 VSS 0.056945f
C6546 ASIG5V.n8971 VSS 0.056945f
C6547 ASIG5V.n8972 VSS 0.056945f
C6548 ASIG5V.n8973 VSS 0.056945f
C6549 ASIG5V.n8975 VSS 0.056945f
C6550 ASIG5V.n8976 VSS 0.056945f
C6551 ASIG5V.n8977 VSS 0.056945f
C6552 ASIG5V.n8978 VSS 0.056945f
C6553 ASIG5V.n8979 VSS 0.056945f
C6554 ASIG5V.n8980 VSS 0.056945f
C6555 ASIG5V.n8981 VSS 0.056945f
C6556 ASIG5V.n8983 VSS 0.056945f
C6557 ASIG5V.n8984 VSS 0.056945f
C6558 ASIG5V.n8985 VSS 0.056945f
C6559 ASIG5V.n8987 VSS 0.056945f
C6560 ASIG5V.n8988 VSS 0.056945f
C6561 ASIG5V.n8989 VSS 0.056945f
C6562 ASIG5V.n8990 VSS 0.056945f
C6563 ASIG5V.n8991 VSS 0.056945f
C6564 ASIG5V.n8992 VSS 0.056945f
C6565 ASIG5V.n8993 VSS 0.056945f
C6566 ASIG5V.n8995 VSS 0.056945f
C6567 ASIG5V.n8996 VSS 0.056945f
C6568 ASIG5V.n8997 VSS 0.056945f
C6569 ASIG5V.n8999 VSS 0.056945f
C6570 ASIG5V.n9000 VSS 0.056945f
C6571 ASIG5V.n9001 VSS 0.056945f
C6572 ASIG5V.n9002 VSS 0.056945f
C6573 ASIG5V.n9003 VSS 0.056945f
C6574 ASIG5V.n9004 VSS 0.056945f
C6575 ASIG5V.n9005 VSS 0.056945f
C6576 ASIG5V.n9007 VSS 0.056945f
C6577 ASIG5V.n9008 VSS 0.056945f
C6578 ASIG5V.n9009 VSS 0.056945f
C6579 ASIG5V.n9011 VSS 0.056945f
C6580 ASIG5V.n9012 VSS 0.056945f
C6581 ASIG5V.n9013 VSS 0.056945f
C6582 ASIG5V.n9014 VSS 0.056945f
C6583 ASIG5V.n9015 VSS 0.056945f
C6584 ASIG5V.n9016 VSS 0.056945f
C6585 ASIG5V.n9017 VSS 0.056945f
C6586 ASIG5V.n9019 VSS 0.056945f
C6587 ASIG5V.n9020 VSS 0.056945f
C6588 ASIG5V.n9021 VSS 0.056945f
C6589 ASIG5V.n9023 VSS 0.056945f
C6590 ASIG5V.n9024 VSS 0.056945f
C6591 ASIG5V.n9025 VSS 0.056945f
C6592 ASIG5V.n9026 VSS 0.056945f
C6593 ASIG5V.n9027 VSS 0.056945f
C6594 ASIG5V.n9028 VSS 0.056945f
C6595 ASIG5V.n9029 VSS 0.056945f
C6596 ASIG5V.n9031 VSS 0.056945f
C6597 ASIG5V.n9032 VSS 0.056945f
C6598 ASIG5V.n9033 VSS 0.056945f
C6599 ASIG5V.n9035 VSS 0.056945f
C6600 ASIG5V.n9036 VSS 0.056945f
C6601 ASIG5V.n9037 VSS 0.056945f
C6602 ASIG5V.n9038 VSS 0.056945f
C6603 ASIG5V.n9039 VSS 0.056945f
C6604 ASIG5V.n9040 VSS 0.056945f
C6605 ASIG5V.n9041 VSS 0.056945f
C6606 ASIG5V.n9043 VSS 0.056945f
C6607 ASIG5V.n9044 VSS 0.056945f
C6608 ASIG5V.n9045 VSS 0.056945f
C6609 ASIG5V.n9047 VSS 0.056945f
C6610 ASIG5V.n9048 VSS 0.056945f
C6611 ASIG5V.n9049 VSS 0.056945f
C6612 ASIG5V.n9050 VSS 0.056945f
C6613 ASIG5V.n9051 VSS 0.056945f
C6614 ASIG5V.n9052 VSS 0.056945f
C6615 ASIG5V.n9053 VSS 0.056945f
C6616 ASIG5V.n9055 VSS 0.056945f
C6617 ASIG5V.n9056 VSS 0.056945f
C6618 ASIG5V.n9057 VSS 0.056945f
C6619 ASIG5V.n9059 VSS 0.056945f
C6620 ASIG5V.n9060 VSS 0.056945f
C6621 ASIG5V.n9061 VSS 0.056945f
C6622 ASIG5V.n9062 VSS 0.056945f
C6623 ASIG5V.n9063 VSS 0.056945f
C6624 ASIG5V.n9064 VSS 0.056945f
C6625 ASIG5V.n9065 VSS 0.056945f
C6626 ASIG5V.n9067 VSS 0.056945f
C6627 ASIG5V.n9068 VSS 0.056945f
C6628 ASIG5V.n9069 VSS 0.056945f
C6629 ASIG5V.n9071 VSS 0.056945f
C6630 ASIG5V.n9072 VSS 0.056945f
C6631 ASIG5V.n9073 VSS 0.056945f
C6632 ASIG5V.n9074 VSS 0.056945f
C6633 ASIG5V.n9075 VSS 0.056945f
C6634 ASIG5V.n9076 VSS 0.056945f
C6635 ASIG5V.n9077 VSS 0.056945f
C6636 ASIG5V.n9079 VSS 0.056945f
C6637 ASIG5V.n9080 VSS 0.056945f
C6638 ASIG5V.n9081 VSS 0.056945f
C6639 ASIG5V.n9083 VSS 0.056945f
C6640 ASIG5V.n9084 VSS 0.056945f
C6641 ASIG5V.n9085 VSS 0.056945f
C6642 ASIG5V.n9086 VSS 0.056945f
C6643 ASIG5V.n9087 VSS 0.056945f
C6644 ASIG5V.n9088 VSS 0.056945f
C6645 ASIG5V.n9089 VSS 0.056945f
C6646 ASIG5V.n9091 VSS 0.056945f
C6647 ASIG5V.n9092 VSS 0.056945f
C6648 ASIG5V.n9093 VSS 0.056945f
C6649 ASIG5V.n9095 VSS 0.056945f
C6650 ASIG5V.n9096 VSS 0.056945f
C6651 ASIG5V.n9097 VSS 0.056945f
C6652 ASIG5V.n9098 VSS 0.056945f
C6653 ASIG5V.n9099 VSS 0.056945f
C6654 ASIG5V.n9100 VSS 0.056945f
C6655 ASIG5V.n9101 VSS 0.056945f
C6656 ASIG5V.n9103 VSS 0.056945f
C6657 ASIG5V.n9104 VSS 0.056945f
C6658 ASIG5V.n9105 VSS 0.056945f
C6659 ASIG5V.n9107 VSS 0.056945f
C6660 ASIG5V.n9108 VSS 0.056945f
C6661 ASIG5V.n9109 VSS 0.056945f
C6662 ASIG5V.n9110 VSS 0.056945f
C6663 ASIG5V.n9111 VSS 0.056945f
C6664 ASIG5V.n9112 VSS 0.056945f
C6665 ASIG5V.n9113 VSS 0.056945f
C6666 ASIG5V.n9115 VSS 0.056945f
C6667 ASIG5V.n9116 VSS 0.056945f
C6668 ASIG5V.n9117 VSS 0.056945f
C6669 ASIG5V.n9119 VSS 0.056945f
C6670 ASIG5V.n9120 VSS 0.056945f
C6671 ASIG5V.n9121 VSS 0.056945f
C6672 ASIG5V.n9122 VSS 0.056945f
C6673 ASIG5V.n9123 VSS 0.056945f
C6674 ASIG5V.n9124 VSS 0.056945f
C6675 ASIG5V.n9125 VSS 0.056945f
C6676 ASIG5V.n9127 VSS 0.056945f
C6677 ASIG5V.n9128 VSS 0.056945f
C6678 ASIG5V.n9129 VSS 0.056945f
C6679 ASIG5V.n9131 VSS 0.056945f
C6680 ASIG5V.n9132 VSS 0.056945f
C6681 ASIG5V.n9133 VSS 0.056945f
C6682 ASIG5V.n9134 VSS 0.056945f
C6683 ASIG5V.n9135 VSS 0.056945f
C6684 ASIG5V.n9136 VSS 0.056945f
C6685 ASIG5V.n9137 VSS 0.056945f
C6686 ASIG5V.n9139 VSS 0.056945f
C6687 ASIG5V.n9140 VSS 0.056945f
C6688 ASIG5V.n9141 VSS 0.056945f
C6689 ASIG5V.n9143 VSS 0.056945f
C6690 ASIG5V.n9144 VSS 0.056945f
C6691 ASIG5V.n9145 VSS 0.056945f
C6692 ASIG5V.n9146 VSS 0.056945f
C6693 ASIG5V.n9147 VSS 0.056945f
C6694 ASIG5V.n9148 VSS 0.056945f
C6695 ASIG5V.n9149 VSS 0.056945f
C6696 ASIG5V.n9151 VSS 0.056945f
C6697 ASIG5V.n9152 VSS 0.056945f
C6698 ASIG5V.n9153 VSS 0.056945f
C6699 ASIG5V.n9155 VSS 0.056945f
C6700 ASIG5V.n9156 VSS 0.056945f
C6701 ASIG5V.n9157 VSS 0.056945f
C6702 ASIG5V.n9158 VSS 0.056945f
C6703 ASIG5V.n9159 VSS 0.056945f
C6704 ASIG5V.n9160 VSS 0.056945f
C6705 ASIG5V.n9161 VSS 0.056945f
C6706 ASIG5V.n9163 VSS 0.056945f
C6707 ASIG5V.n9164 VSS 0.056945f
C6708 ASIG5V.n9165 VSS 0.056945f
C6709 ASIG5V.n9167 VSS 0.056945f
C6710 ASIG5V.n9168 VSS 0.056945f
C6711 ASIG5V.n9169 VSS 0.056945f
C6712 ASIG5V.n9170 VSS 0.056945f
C6713 ASIG5V.n9171 VSS 0.056945f
C6714 ASIG5V.n9172 VSS 0.056945f
C6715 ASIG5V.n9173 VSS 0.056945f
C6716 ASIG5V.n9175 VSS 0.036092f
C6717 ASIG5V.n9176 VSS 0.084754f
C6718 ASIG5V.n9177 VSS 0.878365f
C6719 ASIG5V.n9178 VSS 0.056991f
C6720 ASIG5V.n9179 VSS 0.056991f
C6721 ASIG5V.n9180 VSS 0.049774f
C6722 ASIG5V.n9181 VSS 0.052746f
C6723 ASIG5V.n9182 VSS 0.050718f
C6724 ASIG5V.n9183 VSS 0.058072f
C6725 ASIG5V.n9184 VSS 0.058072f
C6726 ASIG5V.n9185 VSS 0.739676f
C6727 ASIG5V.n9186 VSS 1.0941f
C6728 ASIG5V.n9187 VSS 0.108961f
C6729 ASIG5V.n9188 VSS 0.101931f
C6730 ASIG5V.n9189 VSS 0.101931f
C6731 ASIG5V.n9190 VSS 0.051768f
C6732 ASIG5V.n9191 VSS 0.07229f
C6733 ASIG5V.n9192 VSS 0.052133f
C6734 ASIG5V.n9193 VSS 0.056945f
C6735 ASIG5V.n9194 VSS 0.056945f
C6736 ASIG5V.n9195 VSS 0.056945f
C6737 ASIG5V.n9196 VSS 0.056945f
C6738 ASIG5V.n9197 VSS 0.056945f
C6739 ASIG5V.n9198 VSS 0.056945f
C6740 ASIG5V.n9199 VSS 0.056945f
C6741 ASIG5V.n9200 VSS 0.056945f
C6742 ASIG5V.n9201 VSS 0.056945f
C6743 ASIG5V.n9202 VSS 0.056945f
C6744 ASIG5V.n9203 VSS 0.056945f
C6745 ASIG5V.n9204 VSS 0.056945f
C6746 ASIG5V.n9205 VSS 0.056945f
C6747 ASIG5V.n9206 VSS 0.056945f
C6748 ASIG5V.n9207 VSS 0.056945f
C6749 ASIG5V.n9208 VSS 0.056945f
C6750 ASIG5V.n9209 VSS 0.056945f
C6751 ASIG5V.n9210 VSS 0.056945f
C6752 ASIG5V.n9211 VSS 0.056945f
C6753 ASIG5V.n9212 VSS 0.056945f
C6754 ASIG5V.n9213 VSS 0.056945f
C6755 ASIG5V.n9214 VSS 0.056945f
C6756 ASIG5V.n9215 VSS 0.056945f
C6757 ASIG5V.n9216 VSS 0.056945f
C6758 ASIG5V.n9217 VSS 0.056945f
C6759 ASIG5V.n9218 VSS 0.056945f
C6760 ASIG5V.n9219 VSS 0.056945f
C6761 ASIG5V.n9220 VSS 0.056945f
C6762 ASIG5V.n9221 VSS 0.056945f
C6763 ASIG5V.n9222 VSS 0.056945f
C6764 ASIG5V.n9223 VSS 0.056945f
C6765 ASIG5V.n9224 VSS 0.056945f
C6766 ASIG5V.n9225 VSS 0.056945f
C6767 ASIG5V.n9226 VSS 0.056945f
C6768 ASIG5V.n9227 VSS 0.056945f
C6769 ASIG5V.n9228 VSS 0.056945f
C6770 ASIG5V.n9229 VSS 0.056945f
C6771 ASIG5V.n9230 VSS 0.056945f
C6772 ASIG5V.n9231 VSS 0.056945f
C6773 ASIG5V.n9232 VSS 0.056945f
C6774 ASIG5V.n9233 VSS 0.056945f
C6775 ASIG5V.n9234 VSS 0.056945f
C6776 ASIG5V.n9235 VSS 0.056945f
C6777 ASIG5V.n9236 VSS 0.056945f
C6778 ASIG5V.n9237 VSS 0.056945f
C6779 ASIG5V.n9238 VSS 0.056945f
C6780 ASIG5V.n9239 VSS 0.056945f
C6781 ASIG5V.n9240 VSS 0.056945f
C6782 ASIG5V.n9241 VSS 0.056945f
C6783 ASIG5V.n9242 VSS 0.056945f
C6784 ASIG5V.n9243 VSS 0.056945f
C6785 ASIG5V.n9244 VSS 0.056945f
C6786 ASIG5V.n9245 VSS 0.056945f
C6787 ASIG5V.n9246 VSS 0.056945f
C6788 ASIG5V.n9247 VSS 0.056945f
C6789 ASIG5V.n9248 VSS 0.056945f
C6790 ASIG5V.n9249 VSS 0.056945f
C6791 ASIG5V.n9250 VSS 0.056945f
C6792 ASIG5V.n9251 VSS 0.056945f
C6793 ASIG5V.n9252 VSS 0.056945f
C6794 ASIG5V.n9253 VSS 0.056945f
C6795 ASIG5V.n9254 VSS 0.056945f
C6796 ASIG5V.n9255 VSS 0.056945f
C6797 ASIG5V.n9256 VSS 0.056945f
C6798 ASIG5V.n9257 VSS 0.056945f
C6799 ASIG5V.n9258 VSS 0.056945f
C6800 ASIG5V.n9259 VSS 0.056945f
C6801 ASIG5V.n9260 VSS 0.056945f
C6802 ASIG5V.n9261 VSS 0.056945f
C6803 ASIG5V.n9262 VSS 0.056945f
C6804 ASIG5V.n9263 VSS 0.056945f
C6805 ASIG5V.n9264 VSS 0.056945f
C6806 ASIG5V.n9265 VSS 0.056945f
C6807 ASIG5V.n9266 VSS 0.056945f
C6808 ASIG5V.n9267 VSS 0.056945f
C6809 ASIG5V.n9268 VSS 0.056945f
C6810 ASIG5V.n9269 VSS 0.056945f
C6811 ASIG5V.n9270 VSS 0.056945f
C6812 ASIG5V.n9271 VSS 0.056945f
C6813 ASIG5V.n9272 VSS 0.056945f
C6814 ASIG5V.n9273 VSS 0.056945f
C6815 ASIG5V.n9274 VSS 0.056945f
C6816 ASIG5V.n9275 VSS 0.056945f
C6817 ASIG5V.n9276 VSS 0.056945f
C6818 ASIG5V.n9277 VSS 0.056945f
C6819 ASIG5V.n9278 VSS 0.056945f
C6820 ASIG5V.n9279 VSS 0.056945f
C6821 ASIG5V.n9280 VSS 0.056945f
C6822 ASIG5V.n9281 VSS 0.056945f
C6823 ASIG5V.n9282 VSS 0.056945f
C6824 ASIG5V.n9283 VSS 0.056945f
C6825 ASIG5V.n9284 VSS 0.056945f
C6826 ASIG5V.n9285 VSS 0.056945f
C6827 ASIG5V.n9286 VSS 0.056945f
C6828 ASIG5V.n9287 VSS 0.056945f
C6829 ASIG5V.n9288 VSS 0.056945f
C6830 ASIG5V.n9289 VSS 0.056945f
C6831 ASIG5V.n9290 VSS 0.056945f
C6832 ASIG5V.n9291 VSS 0.056945f
C6833 ASIG5V.n9292 VSS 0.056945f
C6834 ASIG5V.n9293 VSS 0.056945f
C6835 ASIG5V.n9294 VSS 0.056945f
C6836 ASIG5V.n9295 VSS 0.056945f
C6837 ASIG5V.n9296 VSS 0.056945f
C6838 ASIG5V.n9297 VSS 0.056945f
C6839 ASIG5V.n9298 VSS 0.056945f
C6840 ASIG5V.n9299 VSS 0.056945f
C6841 ASIG5V.n9300 VSS 0.056945f
C6842 ASIG5V.n9301 VSS 0.056945f
C6843 ASIG5V.n9302 VSS 0.056945f
C6844 ASIG5V.n9303 VSS 0.056945f
C6845 ASIG5V.n9304 VSS 0.056945f
C6846 ASIG5V.n9305 VSS 0.056945f
C6847 ASIG5V.n9306 VSS 0.056945f
C6848 ASIG5V.n9307 VSS 0.056945f
C6849 ASIG5V.n9308 VSS 0.056945f
C6850 ASIG5V.n9309 VSS 0.056945f
C6851 ASIG5V.n9310 VSS 0.056945f
C6852 ASIG5V.n9311 VSS 0.056945f
C6853 ASIG5V.n9312 VSS 0.056945f
C6854 ASIG5V.n9313 VSS 0.056945f
C6855 ASIG5V.n9314 VSS 0.056945f
C6856 ASIG5V.n9315 VSS 0.056945f
C6857 ASIG5V.n9316 VSS 0.056945f
C6858 ASIG5V.n9317 VSS 0.056945f
C6859 ASIG5V.n9318 VSS 0.056945f
C6860 ASIG5V.n9319 VSS 0.056945f
C6861 ASIG5V.n9320 VSS 0.056945f
C6862 ASIG5V.n9321 VSS 0.056945f
C6863 ASIG5V.n9322 VSS 0.056945f
C6864 ASIG5V.n9323 VSS 0.056945f
C6865 ASIG5V.n9324 VSS 0.056945f
C6866 ASIG5V.n9325 VSS 0.056945f
C6867 ASIG5V.n9326 VSS 0.056945f
C6868 ASIG5V.n9327 VSS 0.056945f
C6869 ASIG5V.n9328 VSS 0.056945f
C6870 ASIG5V.n9329 VSS 0.056945f
C6871 ASIG5V.n9330 VSS 0.056945f
C6872 ASIG5V.n9331 VSS 0.056945f
C6873 ASIG5V.n9332 VSS 0.056945f
C6874 ASIG5V.n9333 VSS 0.056945f
C6875 ASIG5V.n9334 VSS 0.056945f
C6876 ASIG5V.n9335 VSS 0.056945f
C6877 ASIG5V.n9336 VSS 0.056945f
C6878 ASIG5V.n9337 VSS 0.056945f
C6879 ASIG5V.n9338 VSS 0.056945f
C6880 ASIG5V.n9339 VSS 0.056945f
C6881 ASIG5V.n9340 VSS 0.056945f
C6882 ASIG5V.n9341 VSS 0.056945f
C6883 ASIG5V.n9342 VSS 0.056945f
C6884 ASIG5V.n9343 VSS 0.056945f
C6885 ASIG5V.n9344 VSS 0.056945f
C6886 ASIG5V.n9345 VSS 0.056945f
C6887 ASIG5V.n9346 VSS 0.056945f
C6888 ASIG5V.n9347 VSS 0.056945f
C6889 ASIG5V.n9348 VSS 0.056945f
C6890 ASIG5V.n9349 VSS 0.056945f
C6891 ASIG5V.n9350 VSS 0.056945f
C6892 ASIG5V.n9351 VSS 0.056945f
C6893 ASIG5V.n9352 VSS 0.056945f
C6894 ASIG5V.n9353 VSS 0.056945f
C6895 ASIG5V.n9354 VSS 0.056945f
C6896 ASIG5V.n9355 VSS 0.056945f
C6897 ASIG5V.n9356 VSS 0.056945f
C6898 ASIG5V.n9357 VSS 0.056945f
C6899 ASIG5V.n9358 VSS 0.056945f
C6900 ASIG5V.n9359 VSS 0.056945f
C6901 ASIG5V.n9360 VSS 0.056945f
C6902 ASIG5V.n9361 VSS 0.056945f
C6903 ASIG5V.n9362 VSS 0.056945f
C6904 ASIG5V.n9363 VSS 0.056945f
C6905 ASIG5V.n9364 VSS 0.056945f
C6906 ASIG5V.n9365 VSS 0.056945f
C6907 ASIG5V.n9366 VSS 0.056945f
C6908 ASIG5V.n9367 VSS 0.056945f
C6909 ASIG5V.n9368 VSS 0.056945f
C6910 ASIG5V.n9369 VSS 0.056945f
C6911 ASIG5V.n9370 VSS 0.056945f
C6912 ASIG5V.n9371 VSS 0.056945f
C6913 ASIG5V.n9372 VSS 0.056945f
C6914 ASIG5V.n9373 VSS 0.056945f
C6915 ASIG5V.n9374 VSS 0.056945f
C6916 ASIG5V.n9375 VSS 0.056945f
C6917 ASIG5V.n9376 VSS 0.047722f
C6918 ASIG5V.n9377 VSS 0.036092f
C6919 ASIG5V.n9378 VSS 0.036092f
C6920 ASIG5V.n9379 VSS 0.500822f
C6921 ASIG5V.n9380 VSS 0.036092f
C6922 ASIG5V.n9382 VSS 0.639512f
C6923 ASIG5V.n9383 VSS 0.523937f
C6924 ASIG5V.n9384 VSS 0.065094f
C6925 ASIG5V.n9385 VSS 0.065094f
C6926 ASIG5V.n9386 VSS 0.056851f
C6927 ASIG5V.n9387 VSS 0.066995f
C6928 ASIG5V.n9388 VSS 0.037508f
C6929 ASIG5V.n9389 VSS 0.042946f
C6930 ASIG5V.n9390 VSS 0.045974f
C6931 ASIG5V.n9391 VSS 0.036092f
C6932 ASIG5V.n9392 VSS 0.036092f
C6933 ASIG5V.n9393 VSS 0.916891f
C6934 ASIG5V.n9394 VSS 0.036092f
C6935 ASIG5V.n9396 VSS 0.955415f
C6936 ASIG5V.n9397 VSS 0.431477f
C6937 ASIG5V.n9398 VSS 0.103688f
C6938 ASIG5V.n9399 VSS 0.103688f
C6939 ASIG5V.n9400 VSS 0.092554f
C6940 ASIG5V.n9401 VSS 0.09726f
C6941 ASIG5V.n9402 VSS 0.064317f
C6942 ASIG5V.n9403 VSS 0.072055f
C6943 ASIG5V.n9404 VSS 0.072055f
C6944 ASIG5V.n9405 VSS 0.654922f
C6945 ASIG5V.n9406 VSS 0.816725f
C6946 ASIG5V.n9407 VSS 0.040785f
C6947 ASIG5V.n9408 VSS 0.040785f
C6948 ASIG5V.n9409 VSS 0.03562f
C6949 ASIG5V.n9410 VSS 0.066995f
C6950 ASIG5V.n9411 VSS 0.058738f
C6951 ASIG5V.n9412 VSS 0.067255f
C6952 ASIG5V.n9413 VSS 0.045974f
C6953 ASIG5V.n9414 VSS 0.036092f
C6954 ASIG5V.n9415 VSS 0.036092f
C6955 ASIG5V.n9416 VSS 0.300493f
C6956 ASIG5V.n9417 VSS 0.036092f
C6957 ASIG5V.n9419 VSS 0.932301f
C6958 ASIG5V.n9420 VSS 0.847545f
C6959 ASIG5V.n9421 VSS 0.076709f
C6960 ASIG5V.n9422 VSS 0.060233f
C6961 ASIG5V.n9423 VSS 0.060233f
C6962 ASIG5V.n9424 VSS 0.052605f
C6963 ASIG5V.n9425 VSS 0.052746f
C6964 ASIG5V.n9426 VSS 0.047722f
C6965 ASIG5V.n9427 VSS 0.056945f
C6966 ASIG5V.n9428 VSS 0.056945f
C6967 ASIG5V.n9429 VSS 0.056945f
C6968 ASIG5V.n9431 VSS 0.036092f
C6969 ASIG5V.n9432 VSS 0.839841f
C6970 ASIG5V.n9433 VSS 1.05558f
C6971 ASIG5V.n9434 VSS 0.066782f
C6972 ASIG5V.n9435 VSS 0.066782f
C6973 ASIG5V.n9436 VSS 0.059611f
C6974 ASIG5V.n9437 VSS 0.09726f
C6975 ASIG5V.n9438 VSS 0.09726f
C6976 ASIG5V.n9439 VSS 0.108961f
C6977 ASIG5V.n9440 VSS 0.108961f
C6978 ASIG5V.n9441 VSS 0.932301f
C6979 ASIG5V.n9442 VSS 0.036092f
C6980 ASIG5V.n9443 VSS 0.056945f
C6981 ASIG5V.n9444 VSS 0.056945f
C6982 ASIG5V.n9445 VSS 0.056945f
C6983 ASIG5V.n9446 VSS 0.056945f
C6984 ASIG5V.n9447 VSS 0.056945f
C6985 ASIG5V.n9448 VSS 0.056945f
C6986 ASIG5V.n9449 VSS 0.056945f
C6987 ASIG5V.n9450 VSS 0.056945f
C6988 ASIG5V.n9451 VSS 0.056945f
C6989 ASIG5V.n9452 VSS 0.056945f
C6990 ASIG5V.n9453 VSS 0.056945f
C6991 ASIG5V.n9454 VSS 0.056945f
C6992 ASIG5V.n9455 VSS 0.056945f
C6993 ASIG5V.n9456 VSS 0.056945f
C6994 ASIG5V.n9457 VSS 0.056945f
C6995 ASIG5V.n9458 VSS 0.056945f
C6996 ASIG5V.n9459 VSS 0.056945f
C6997 ASIG5V.n9460 VSS 0.056945f
C6998 ASIG5V.n9461 VSS 0.056945f
C6999 ASIG5V.n9462 VSS 0.056945f
C7000 ASIG5V.n9463 VSS 0.056945f
C7001 ASIG5V.n9464 VSS 0.056945f
C7002 ASIG5V.n9465 VSS 0.056945f
C7003 ASIG5V.n9466 VSS 0.056945f
C7004 ASIG5V.n9467 VSS 0.056945f
C7005 ASIG5V.n9468 VSS 0.056945f
C7006 ASIG5V.n9469 VSS 0.056945f
C7007 ASIG5V.n9470 VSS 0.056945f
C7008 ASIG5V.n9471 VSS 0.056945f
C7009 ASIG5V.n9472 VSS 0.056945f
C7010 ASIG5V.n9473 VSS 0.056945f
C7011 ASIG5V.n9474 VSS 0.056945f
C7012 ASIG5V.n9475 VSS 0.056945f
C7013 ASIG5V.n9476 VSS 0.056945f
C7014 ASIG5V.n9477 VSS 0.056945f
C7015 ASIG5V.n9478 VSS 0.056945f
C7016 ASIG5V.n9479 VSS 0.056945f
C7017 ASIG5V.n9480 VSS 0.056945f
C7018 ASIG5V.n9481 VSS 0.056945f
C7019 ASIG5V.n9482 VSS 0.056945f
C7020 ASIG5V.n9484 VSS 0.056945f
C7021 ASIG5V.n9485 VSS 0.056945f
C7022 ASIG5V.n9486 VSS 0.036092f
C7023 ASIG5V.n9487 VSS 0.052133f
C7024 ASIG5V.n9488 VSS 0.056945f
C7025 ASIG5V.n9489 VSS 0.056945f
C7026 ASIG5V.n9490 VSS 0.056945f
C7027 ASIG5V.n9491 VSS 0.056945f
C7028 ASIG5V.n9493 VSS 0.056945f
C7029 ASIG5V.n9494 VSS 0.056945f
C7030 ASIG5V.n9495 VSS 0.056945f
C7031 ASIG5V.n9497 VSS 0.056945f
C7032 ASIG5V.n9498 VSS 0.056945f
C7033 ASIG5V.n9499 VSS 0.056945f
C7034 ASIG5V.n9500 VSS 0.056945f
C7035 ASIG5V.n9501 VSS 0.056945f
C7036 ASIG5V.n9502 VSS 0.056945f
C7037 ASIG5V.n9503 VSS 0.056945f
C7038 ASIG5V.n9505 VSS 0.056945f
C7039 ASIG5V.n9506 VSS 0.056945f
C7040 ASIG5V.n9507 VSS 0.056945f
C7041 ASIG5V.n9509 VSS 0.056945f
C7042 ASIG5V.n9510 VSS 0.056945f
C7043 ASIG5V.n9511 VSS 0.056945f
C7044 ASIG5V.n9512 VSS 0.056945f
C7045 ASIG5V.n9513 VSS 0.056945f
C7046 ASIG5V.n9514 VSS 0.056945f
C7047 ASIG5V.n9515 VSS 0.056945f
C7048 ASIG5V.n9517 VSS 0.056945f
C7049 ASIG5V.n9518 VSS 0.056945f
C7050 ASIG5V.n9519 VSS 0.056945f
C7051 ASIG5V.n9521 VSS 0.056945f
C7052 ASIG5V.n9522 VSS 0.056945f
C7053 ASIG5V.n9523 VSS 0.056945f
C7054 ASIG5V.n9524 VSS 0.056945f
C7055 ASIG5V.n9525 VSS 0.056945f
C7056 ASIG5V.n9526 VSS 0.056945f
C7057 ASIG5V.n9527 VSS 0.056945f
C7058 ASIG5V.n9529 VSS 0.056945f
C7059 ASIG5V.n9530 VSS 0.056945f
C7060 ASIG5V.n9531 VSS 0.056945f
C7061 ASIG5V.n9533 VSS 0.056945f
C7062 ASIG5V.n9534 VSS 0.056945f
C7063 ASIG5V.n9535 VSS 0.056945f
C7064 ASIG5V.n9536 VSS 0.056945f
C7065 ASIG5V.n9537 VSS 0.056945f
C7066 ASIG5V.n9538 VSS 0.056945f
C7067 ASIG5V.n9539 VSS 0.056945f
C7068 ASIG5V.n9541 VSS 0.056945f
C7069 ASIG5V.n9542 VSS 0.056945f
C7070 ASIG5V.n9543 VSS 0.056945f
C7071 ASIG5V.n9545 VSS 0.056945f
C7072 ASIG5V.n9546 VSS 0.056945f
C7073 ASIG5V.n9547 VSS 0.056945f
C7074 ASIG5V.n9548 VSS 0.056945f
C7075 ASIG5V.n9549 VSS 0.056945f
C7076 ASIG5V.n9550 VSS 0.056945f
C7077 ASIG5V.n9551 VSS 0.056945f
C7078 ASIG5V.n9553 VSS 0.056945f
C7079 ASIG5V.n9554 VSS 0.056945f
C7080 ASIG5V.n9555 VSS 0.056945f
C7081 ASIG5V.n9557 VSS 0.056945f
C7082 ASIG5V.n9558 VSS 0.056945f
C7083 ASIG5V.n9559 VSS 0.056945f
C7084 ASIG5V.n9560 VSS 0.056945f
C7085 ASIG5V.n9561 VSS 0.056945f
C7086 ASIG5V.n9562 VSS 0.056945f
C7087 ASIG5V.n9563 VSS 0.056945f
C7088 ASIG5V.n9565 VSS 0.056945f
C7089 ASIG5V.n9566 VSS 0.056945f
C7090 ASIG5V.n9567 VSS 0.056945f
C7091 ASIG5V.n9569 VSS 0.056945f
C7092 ASIG5V.n9570 VSS 0.056945f
C7093 ASIG5V.n9571 VSS 0.056945f
C7094 ASIG5V.n9572 VSS 0.056945f
C7095 ASIG5V.n9573 VSS 0.056945f
C7096 ASIG5V.n9574 VSS 0.056945f
C7097 ASIG5V.n9575 VSS 0.056945f
C7098 ASIG5V.n9577 VSS 0.056945f
C7099 ASIG5V.n9578 VSS 0.056945f
C7100 ASIG5V.n9579 VSS 0.056945f
C7101 ASIG5V.n9581 VSS 0.056945f
C7102 ASIG5V.n9582 VSS 0.056945f
C7103 ASIG5V.n9583 VSS 0.056945f
C7104 ASIG5V.n9584 VSS 0.056945f
C7105 ASIG5V.n9585 VSS 0.056945f
C7106 ASIG5V.n9586 VSS 0.056945f
C7107 ASIG5V.n9587 VSS 0.056945f
C7108 ASIG5V.n9589 VSS 0.056945f
C7109 ASIG5V.n9590 VSS 0.056945f
C7110 ASIG5V.n9591 VSS 0.056945f
C7111 ASIG5V.n9593 VSS 0.056945f
C7112 ASIG5V.n9594 VSS 0.056945f
C7113 ASIG5V.n9595 VSS 0.056945f
C7114 ASIG5V.n9596 VSS 0.056945f
C7115 ASIG5V.n9597 VSS 0.056945f
C7116 ASIG5V.n9598 VSS 0.056945f
C7117 ASIG5V.n9599 VSS 0.056945f
C7118 ASIG5V.n9601 VSS 0.056945f
C7119 ASIG5V.n9602 VSS 0.056945f
C7120 ASIG5V.n9603 VSS 0.056945f
C7121 ASIG5V.n9605 VSS 0.056945f
C7122 ASIG5V.n9606 VSS 0.056945f
C7123 ASIG5V.n9607 VSS 0.056945f
C7124 ASIG5V.n9608 VSS 0.056945f
C7125 ASIG5V.n9609 VSS 0.056945f
C7126 ASIG5V.n9610 VSS 0.056945f
C7127 ASIG5V.n9611 VSS 0.056945f
C7128 ASIG5V.n9613 VSS 0.056945f
C7129 ASIG5V.n9614 VSS 0.056945f
C7130 ASIG5V.n9615 VSS 0.056945f
C7131 ASIG5V.n9617 VSS 0.056945f
C7132 ASIG5V.n9618 VSS 0.056945f
C7133 ASIG5V.n9619 VSS 0.056945f
C7134 ASIG5V.n9620 VSS 0.056945f
C7135 ASIG5V.n9621 VSS 0.056945f
C7136 ASIG5V.n9622 VSS 0.056945f
C7137 ASIG5V.n9623 VSS 0.056945f
C7138 ASIG5V.n9625 VSS 0.056945f
C7139 ASIG5V.n9626 VSS 0.056945f
C7140 ASIG5V.n9627 VSS 0.056945f
C7141 ASIG5V.n9629 VSS 0.056945f
C7142 ASIG5V.n9630 VSS 0.056945f
C7143 ASIG5V.n9631 VSS 0.056945f
C7144 ASIG5V.n9632 VSS 0.056945f
C7145 ASIG5V.n9633 VSS 0.056945f
C7146 ASIG5V.n9634 VSS 0.056945f
C7147 ASIG5V.n9635 VSS 0.056945f
C7148 ASIG5V.n9637 VSS 0.056945f
C7149 ASIG5V.n9638 VSS 0.056945f
C7150 ASIG5V.n9639 VSS 0.056945f
C7151 ASIG5V.n9641 VSS 0.056945f
C7152 ASIG5V.n9642 VSS 0.056945f
C7153 ASIG5V.n9643 VSS 0.056945f
C7154 ASIG5V.n9644 VSS 0.056945f
C7155 ASIG5V.n9645 VSS 0.056945f
C7156 ASIG5V.n9646 VSS 0.056945f
C7157 ASIG5V.n9647 VSS 0.056945f
C7158 ASIG5V.n9649 VSS 0.056945f
C7159 ASIG5V.n9650 VSS 0.056945f
C7160 ASIG5V.n9651 VSS 0.056945f
C7161 ASIG5V.n9653 VSS 0.056945f
C7162 ASIG5V.n9654 VSS 0.056945f
C7163 ASIG5V.n9655 VSS 0.056945f
C7164 ASIG5V.n9656 VSS 0.056945f
C7165 ASIG5V.n9657 VSS 0.056945f
C7166 ASIG5V.n9658 VSS 0.056945f
C7167 ASIG5V.n9659 VSS 0.056945f
C7168 ASIG5V.n9661 VSS 0.056945f
C7169 ASIG5V.n9662 VSS 0.056945f
C7170 ASIG5V.n9663 VSS 0.056945f
C7171 ASIG5V.n9665 VSS 0.056945f
C7172 ASIG5V.n9666 VSS 0.056945f
C7173 ASIG5V.n9667 VSS 0.056945f
C7174 ASIG5V.n9668 VSS 0.056945f
C7175 ASIG5V.n9669 VSS 0.056945f
C7176 ASIG5V.n9670 VSS 0.056945f
C7177 ASIG5V.n9671 VSS 0.056945f
C7178 ASIG5V.n9673 VSS 0.056945f
C7179 ASIG5V.n9674 VSS 0.056945f
C7180 ASIG5V.n9675 VSS 0.056945f
C7181 ASIG5V.n9677 VSS 0.056945f
C7182 ASIG5V.n9678 VSS 0.056945f
C7183 ASIG5V.n9679 VSS 0.056945f
C7184 ASIG5V.n9680 VSS 0.056945f
C7185 ASIG5V.n9681 VSS 0.056945f
C7186 ASIG5V.n9682 VSS 0.056945f
C7187 ASIG5V.n9683 VSS 0.056945f
C7188 ASIG5V.n9685 VSS 0.056945f
C7189 ASIG5V.n9686 VSS 0.056945f
C7190 ASIG5V.n9687 VSS 0.056945f
C7191 ASIG5V.n9689 VSS 0.056945f
C7192 ASIG5V.n9690 VSS 0.056945f
C7193 ASIG5V.n9691 VSS 0.056945f
C7194 ASIG5V.n9692 VSS 0.056945f
C7195 ASIG5V.n9693 VSS 0.056945f
C7196 ASIG5V.n9694 VSS 0.056945f
C7197 ASIG5V.n9695 VSS 0.056945f
C7198 ASIG5V.n9697 VSS 0.056945f
C7199 ASIG5V.n9698 VSS 0.056945f
C7200 ASIG5V.n9699 VSS 0.056945f
C7201 ASIG5V.n9701 VSS 0.056945f
C7202 ASIG5V.n9702 VSS 0.056945f
C7203 ASIG5V.n9703 VSS 0.056945f
C7204 ASIG5V.n9704 VSS 0.056945f
C7205 ASIG5V.n9705 VSS 0.056945f
C7206 ASIG5V.n9706 VSS 0.056945f
C7207 ASIG5V.n9707 VSS 0.056945f
C7208 ASIG5V.n9709 VSS 0.056945f
C7209 ASIG5V.n9710 VSS 0.056945f
C7210 ASIG5V.n9711 VSS 0.056945f
C7211 ASIG5V.n9713 VSS 0.056945f
C7212 ASIG5V.n9714 VSS 0.056945f
C7213 ASIG5V.n9715 VSS 0.056945f
C7214 ASIG5V.n9716 VSS 0.056945f
C7215 ASIG5V.n9717 VSS 0.056945f
C7216 ASIG5V.n9718 VSS 0.056945f
C7217 ASIG5V.n9719 VSS 0.056945f
C7218 ASIG5V.n9721 VSS 0.056945f
C7219 ASIG5V.n9722 VSS 0.056945f
C7220 ASIG5V.n9723 VSS 0.056945f
C7221 ASIG5V.n9725 VSS 0.056945f
C7222 ASIG5V.n9726 VSS 0.056945f
C7223 ASIG5V.n9727 VSS 0.056945f
C7224 ASIG5V.n9728 VSS 0.056945f
C7225 ASIG5V.n9729 VSS 0.056945f
C7226 ASIG5V.n9730 VSS 0.056945f
C7227 ASIG5V.n9731 VSS 0.056945f
C7228 ASIG5V.n9733 VSS 0.036092f
C7229 ASIG5V.n9734 VSS 0.531642f
C7230 ASIG5V.n9735 VSS 0.585576f
C7231 ASIG5V.n9736 VSS 0.05321f
C7232 ASIG5V.n9737 VSS 0.05321f
C7233 ASIG5V.n9738 VSS 0.046472f
C7234 ASIG5V.n9739 VSS 0.052746f
C7235 ASIG5V.n9740 VSS 0.05402f
C7236 ASIG5V.n9741 VSS 0.061853f
C7237 ASIG5V.n9742 VSS 0.061853f
C7238 ASIG5V.n9743 VSS 0.446887f
C7239 ASIG5V.n9744 VSS 1.0941f
C7240 ASIG5V.n9745 VSS 0.108961f
C7241 ASIG5V.n9746 VSS 0.108961f
C7242 ASIG5V.n9747 VSS 0.054905f
C7243 ASIG5V.n9748 VSS 0.548344f
C7244 ASIG5V.n9750 VSS 0.087753f
C7245 ASIG5V.n9752 VSS 0.536863f
C7246 ASIG5V.n9753 VSS 0.493967f
C7247 ASIG5V.n9754 VSS 0.309175f
C7248 ASIG5V.n9755 VSS 0.493967f
C7249 ASIG5V.n9757 VSS 0.074298f
C7250 ASIG5V.n9759 VSS 0.087753f
C7251 ASIG5V.n9760 VSS 0.087753f
C7252 ASIG5V.n9762 VSS 0.309175f
C7253 ASIG5V.n9763 VSS 0.314214f
C7254 ASIG5V.n9764 VSS 0.309175f
C7255 ASIG5V.n9765 VSS 0.309175f
C7256 ASIG5V.n9767 VSS 0.087753f
C7257 ASIG5V.n9769 VSS 0.087753f
C7258 ASIG5V.n9770 VSS 0.074298f
C7259 ASIG5V.n9772 VSS 0.493967f
C7260 ASIG5V.n9773 VSS 0.074298f
C7261 ASIG5V.n9775 VSS 0.314214f
C7262 ASIG5V.n9776 VSS 0.309175f
C7263 ASIG5V.n9777 VSS 0.309175f
C7264 ASIG5V.n9779 VSS 0.087753f
C7265 ASIG5V.n9781 VSS 0.087753f
C7266 ASIG5V.n9782 VSS 0.074298f
C7267 ASIG5V.n9784 VSS 0.493967f
C7268 ASIG5V.n9785 VSS 0.074298f
C7269 ASIG5V.n9787 VSS 0.314214f
C7270 ASIG5V.n9788 VSS 0.845738f
C7271 ASIG5V.n9789 VSS 0.845738f
C7272 ASIG5V.n9791 VSS 0.087753f
C7273 ASIG5V.n9793 VSS 0.087753f
C7274 ASIG5V.n9794 VSS 0.074298f
C7275 ASIG5V.n9796 VSS 0.493967f
C7276 ASIG5V.n9797 VSS 0.074298f
C7277 ASIG5V.n9799 VSS 0.314214f
C7278 ASIG5V.n9800 VSS 0.309175f
C7279 ASIG5V.n9801 VSS 0.309175f
C7280 ASIG5V.n9803 VSS 0.087753f
C7281 ASIG5V.n9805 VSS 0.087753f
C7282 ASIG5V.n9806 VSS 0.074298f
C7283 ASIG5V.n9808 VSS 0.493967f
C7284 ASIG5V.n9809 VSS 0.074298f
C7285 ASIG5V.n9811 VSS 0.314214f
C7286 ASIG5V.n9812 VSS 0.309175f
C7287 ASIG5V.n9813 VSS 0.309175f
C7288 ASIG5V.n9815 VSS 0.087753f
C7289 ASIG5V.n9817 VSS 0.087753f
C7290 ASIG5V.n9818 VSS 0.074298f
C7291 ASIG5V.n9820 VSS 0.493967f
C7292 ASIG5V.n9821 VSS 0.074298f
C7293 ASIG5V.n9823 VSS 0.314214f
C7294 ASIG5V.n9824 VSS 0.309175f
C7295 ASIG5V.n9825 VSS 0.309175f
C7296 ASIG5V.n9828 VSS 0.087753f
C7297 ASIG5V.n9830 VSS 0.087753f
C7298 ASIG5V.n9832 VSS 0.074298f
C7299 ASIG5V.n9834 VSS 0.493967f
C7300 ASIG5V.n9835 VSS 0.074298f
C7301 ASIG5V.n9837 VSS 0.314214f
C7302 ASIG5V.n9839 VSS 0.087753f
C7303 ASIG5V.n9841 VSS 0.074298f
C7304 ASIG5V.n9843 VSS 0.314214f
C7305 ASIG5V.n9844 VSS 0.074298f
C7306 ASIG5V.n9846 VSS 0.314214f
C7307 ASIG5V.n9848 VSS 0.087753f
C7308 ASIG5V.n9850 VSS 0.074298f
C7309 ASIG5V.n9852 VSS 0.314214f
C7310 ASIG5V.n9853 VSS 0.074298f
C7311 ASIG5V.n9855 VSS 0.314214f
C7312 ASIG5V.n9857 VSS 0.087753f
C7313 ASIG5V.n9859 VSS 0.074298f
C7314 ASIG5V.n9861 VSS 0.314214f
C7315 ASIG5V.n9862 VSS 0.074298f
C7316 ASIG5V.n9864 VSS 0.250522f
C7317 ASIG5V.t4 VSS 7.07689f
C7318 ASIG5V.n9866 VSS 0.087753f
C7319 ASIG5V.n9868 VSS 0.074298f
C7320 ASIG5V.n9870 VSS 0.250522f
C7321 ASIG5V.n9871 VSS 0.074298f
C7322 ASIG5V.n9873 VSS 0.314214f
C7323 ASIG5V.n9875 VSS 0.087753f
C7324 ASIG5V.n9877 VSS 0.074298f
C7325 ASIG5V.n9879 VSS 0.314214f
C7326 ASIG5V.n9880 VSS 0.074298f
C7327 ASIG5V.n9882 VSS 0.314214f
C7328 ASIG5V.n9883 VSS 0.074298f
C7329 ASIG5V.n9885 VSS 0.314214f
C7330 ASIG5V.n9887 VSS 0.087753f
C7331 ASIG5V.n9889 VSS 0.087753f
C7332 ASIG5V.n9891 VSS 0.309175f
C7333 ASIG5V.n9892 VSS 0.314214f
C7334 ASIG5V.n9893 VSS 0.074298f
C7335 ASIG5V.n9895 VSS 0.074298f
C7336 ASIG5V.n9898 VSS 0.087753f
C7337 ASIG5V.n9899 VSS 0.087753f
C7338 ASIG5V.n9901 VSS 12.9443f
C7339 ASIG5V.n9902 VSS 0.493967f
C7340 ASIG5V.n9903 VSS 0.074298f
C7341 ASIG5V.n9905 VSS 0.314214f
C7342 ASIG5V.n9906 VSS 0.309175f
C7343 ASIG5V.n9907 VSS 0.309175f
C7344 ASIG5V.n9908 VSS 0.493967f
C7345 ASIG5V.n9909 VSS 0.074298f
C7346 ASIG5V.n9911 VSS 0.314214f
C7347 ASIG5V.n9912 VSS 0.309175f
C7348 ASIG5V.n9913 VSS 0.309175f
C7349 ASIG5V.n9914 VSS 0.493967f
C7350 ASIG5V.n9915 VSS 0.074298f
C7351 ASIG5V.n9917 VSS 0.314214f
C7352 ASIG5V.n9918 VSS 0.309175f
C7353 ASIG5V.n9919 VSS 0.309175f
C7354 ASIG5V.n9920 VSS 0.493967f
C7355 ASIG5V.n9921 VSS 0.074298f
C7356 ASIG5V.n9923 VSS 0.314214f
C7357 ASIG5V.n9924 VSS 0.845738f
C7358 ASIG5V.n9925 VSS 0.845738f
C7359 ASIG5V.n9926 VSS 0.493967f
C7360 ASIG5V.n9927 VSS 0.074298f
C7361 ASIG5V.n9929 VSS 0.314214f
C7362 ASIG5V.n9930 VSS 0.309175f
C7363 ASIG5V.n9931 VSS 0.309175f
C7364 ASIG5V.n9932 VSS 0.493967f
C7365 ASIG5V.n9933 VSS 0.074298f
C7366 ASIG5V.n9935 VSS 0.314214f
C7367 ASIG5V.n9936 VSS 0.309175f
C7368 ASIG5V.n9937 VSS 0.309175f
C7369 ASIG5V.n9938 VSS 0.493967f
C7370 ASIG5V.n9939 VSS 0.074298f
C7371 ASIG5V.n9941 VSS 0.314214f
C7372 ASIG5V.n9942 VSS 0.309175f
C7373 ASIG5V.n9943 VSS 0.309175f
C7374 ASIG5V.n9945 VSS 0.314214f
C7375 ASIG5V.n9948 VSS 0.074298f
C7376 ASIG5V.n9950 VSS 0.087753f
C7377 ASIG5V.n9952 VSS 0.536863f
C7378 ASIG5V.n9953 VSS 0.548344f
C7379 ASIG5V.n9954 VSS 0.072161f
C7380 ASIG5V.n9955 VSS 0.094901f
C7381 ASIG5V.n9956 VSS 0.108961f
C7382 ASIG5V.n9957 VSS 0.292788f
C7383 ASIG5V.n9958 VSS 0.094901f
C7384 ASIG5V.n9959 VSS 0.0621f
C7385 ASIG5V.n9960 VSS 0.06854f
C7386 ASIG5V.n9961 VSS 0.07229f
C7387 ASIG5V.n9962 VSS 0.0621f
C7388 ASIG5V.n9963 VSS 0.108961f
C7389 ASIG5V.n9964 VSS 0.0621f
C7390 ASIG5V.n9965 VSS 0.955415f
C7391 ASIG5V.n9966 VSS 0.670332f
C7392 ASIG5V.n9967 VSS 0.045974f
C7393 ASIG5V.n9968 VSS 0.045974f
C7394 ASIG5V.n9969 VSS 0.047722f
C7395 ASIG5V.n9970 VSS 0.066995f
C7396 ASIG5V.n9971 VSS 0.076709f
C7397 ASIG5V.n9972 VSS 0.076709f
C7398 ASIG5V.n9973 VSS 1.02476f
C7399 ASIG5V.n10015 VSS 0.036092f
C7400 ASIG5V.n10016 VSS 0.955415f
C7401 ASIG5V.n10017 VSS 0.056238f
C7402 ASIG5V.n10018 VSS 0.108961f
C7403 ASIG5V.n10019 VSS 0.056238f
C7404 ASIG5V.n10020 VSS 0.108961f
C7405 ASIG5V.n10021 VSS 0.050199f
C7406 ASIG5V.n10022 VSS 0.07229f
C7407 ASIG5V.n10023 VSS 0.0621f
C7408 ASIG5V.n10024 VSS 0.0621f
C7409 ASIG5V.n10025 VSS 0.385247f
C7410 ASIG5V.n10067 VSS 0.036092f
C7411 ASIG5V.n10068 VSS 0.246558f
C7412 ASIG5V.n10069 VSS 0.045974f
C7413 ASIG5V.n10071 VSS 0.056945f
C7414 ASIG5V.n10072 VSS 0.056945f
C7415 ASIG5V.n10073 VSS 0.056945f
C7416 ASIG5V.n10074 VSS 0.056945f
C7417 ASIG5V.n10075 VSS 0.056945f
C7418 ASIG5V.n10076 VSS 0.96312f
C7419 ASIG5V.n10116 VSS 0.036092f
C7420 ASIG5V.n10117 VSS 0.056945f
C7421 ASIG5V.n10118 VSS 0.056945f
C7422 ASIG5V.n10119 VSS 0.052133f
C7423 ASIG5V.n10120 VSS 0.056945f
C7424 ASIG5V.n10121 VSS 0.056945f
C7425 ASIG5V.n10122 VSS 0.056945f
C7426 ASIG5V.n10123 VSS 0.056945f
C7427 ASIG5V.n10124 VSS 0.056945f
C7428 ASIG5V.n10125 VSS 0.056945f
C7429 ASIG5V.n10126 VSS 0.056945f
C7430 ASIG5V.n10127 VSS 0.056945f
C7431 ASIG5V.n10128 VSS 0.056945f
C7432 ASIG5V.n10129 VSS 0.056945f
C7433 ASIG5V.n10130 VSS 0.056945f
C7434 ASIG5V.n10131 VSS 0.056945f
C7435 ASIG5V.n10132 VSS 0.056945f
C7436 ASIG5V.n10133 VSS 0.056945f
C7437 ASIG5V.n10134 VSS 0.056945f
C7438 ASIG5V.n10135 VSS 0.056945f
C7439 ASIG5V.n10136 VSS 0.056945f
C7440 ASIG5V.n10137 VSS 0.056945f
C7441 ASIG5V.n10138 VSS 0.056945f
C7442 ASIG5V.n10139 VSS 0.056945f
C7443 ASIG5V.n10140 VSS 0.056945f
C7444 ASIG5V.n10141 VSS 0.056945f
C7445 ASIG5V.n10142 VSS 0.056945f
C7446 ASIG5V.n10143 VSS 0.056945f
C7447 ASIG5V.n10144 VSS 0.056945f
C7448 ASIG5V.n10145 VSS 0.056945f
C7449 ASIG5V.n10146 VSS 0.056945f
C7450 ASIG5V.n10147 VSS 0.056945f
C7451 ASIG5V.n10148 VSS 0.056945f
C7452 ASIG5V.n10149 VSS 0.056945f
C7453 ASIG5V.n10150 VSS 0.056945f
C7454 ASIG5V.n10151 VSS 0.056945f
C7455 ASIG5V.n10152 VSS 0.056945f
C7456 ASIG5V.n10153 VSS 0.056945f
C7457 ASIG5V.n10154 VSS 0.056945f
C7458 ASIG5V.n10155 VSS 0.056945f
C7459 ASIG5V.n10156 VSS 0.056945f
C7460 ASIG5V.n10157 VSS 0.056945f
C7461 ASIG5V.n10158 VSS 0.056945f
C7462 ASIG5V.n10159 VSS 0.056945f
C7463 ASIG5V.n10160 VSS 0.056945f
C7464 ASIG5V.n10161 VSS 0.056945f
C7465 ASIG5V.n10162 VSS 0.056945f
C7466 ASIG5V.n10163 VSS 0.056945f
C7467 ASIG5V.n10164 VSS 0.056945f
C7468 ASIG5V.n10165 VSS 0.056945f
C7469 ASIG5V.n10166 VSS 0.056945f
C7470 ASIG5V.n10167 VSS 0.056945f
C7471 ASIG5V.n10168 VSS 0.056945f
C7472 ASIG5V.n10169 VSS 0.056945f
C7473 ASIG5V.n10170 VSS 0.056945f
C7474 ASIG5V.n10171 VSS 0.056945f
C7475 ASIG5V.n10172 VSS 0.056945f
C7476 ASIG5V.n10173 VSS 0.056945f
C7477 ASIG5V.n10174 VSS 0.056945f
C7478 ASIG5V.n10175 VSS 0.056945f
C7479 ASIG5V.n10176 VSS 0.056945f
C7480 ASIG5V.n10177 VSS 0.056945f
C7481 ASIG5V.n10178 VSS 0.056945f
C7482 ASIG5V.n10179 VSS 0.056945f
C7483 ASIG5V.n10180 VSS 0.056945f
C7484 ASIG5V.n10181 VSS 0.056945f
C7485 ASIG5V.n10182 VSS 0.056945f
C7486 ASIG5V.n10183 VSS 0.056945f
C7487 ASIG5V.n10184 VSS 0.056945f
C7488 ASIG5V.n10185 VSS 0.056945f
C7489 ASIG5V.n10186 VSS 0.056945f
C7490 ASIG5V.n10187 VSS 0.056945f
C7491 ASIG5V.n10188 VSS 0.056945f
C7492 ASIG5V.n10189 VSS 0.056945f
C7493 ASIG5V.n10190 VSS 0.056945f
C7494 ASIG5V.n10191 VSS 0.056945f
C7495 ASIG5V.n10192 VSS 0.056945f
C7496 ASIG5V.n10193 VSS 0.056945f
C7497 ASIG5V.n10194 VSS 0.056945f
C7498 ASIG5V.n10195 VSS 0.056945f
C7499 ASIG5V.n10196 VSS 0.056945f
C7500 ASIG5V.n10197 VSS 0.056945f
C7501 ASIG5V.n10198 VSS 0.056945f
C7502 ASIG5V.n10199 VSS 0.056945f
C7503 ASIG5V.n10200 VSS 0.056945f
C7504 ASIG5V.n10201 VSS 0.056945f
C7505 ASIG5V.n10202 VSS 0.056945f
C7506 ASIG5V.n10203 VSS 0.056945f
C7507 ASIG5V.n10204 VSS 0.056945f
C7508 ASIG5V.n10205 VSS 0.056945f
C7509 ASIG5V.n10206 VSS 0.056945f
C7510 ASIG5V.n10207 VSS 0.056945f
C7511 ASIG5V.n10208 VSS 0.056945f
C7512 ASIG5V.n10209 VSS 0.056945f
C7513 ASIG5V.n10210 VSS 0.056945f
C7514 ASIG5V.n10211 VSS 0.056945f
C7515 ASIG5V.n10212 VSS 0.056945f
C7516 ASIG5V.n10213 VSS 0.056945f
C7517 ASIG5V.n10214 VSS 0.056945f
C7518 ASIG5V.n10215 VSS 0.056945f
C7519 ASIG5V.n10216 VSS 0.056945f
C7520 ASIG5V.n10217 VSS 0.056945f
C7521 ASIG5V.n10218 VSS 0.056945f
C7522 ASIG5V.n10219 VSS 0.056945f
C7523 ASIG5V.n10220 VSS 0.056945f
C7524 ASIG5V.n10221 VSS 0.056945f
C7525 ASIG5V.n10222 VSS 0.056945f
C7526 ASIG5V.n10223 VSS 0.056945f
C7527 ASIG5V.n10224 VSS 0.056945f
C7528 ASIG5V.n10225 VSS 0.056945f
C7529 ASIG5V.n10226 VSS 0.056945f
C7530 ASIG5V.n10227 VSS 0.056945f
C7531 ASIG5V.n10228 VSS 0.056945f
C7532 ASIG5V.n10229 VSS 0.056945f
C7533 ASIG5V.n10230 VSS 0.056945f
C7534 ASIG5V.n10231 VSS 0.056945f
C7535 ASIG5V.n10232 VSS 0.056945f
C7536 ASIG5V.n10233 VSS 0.056945f
C7537 ASIG5V.n10234 VSS 0.056945f
C7538 ASIG5V.n10235 VSS 0.056945f
C7539 ASIG5V.n10236 VSS 0.056945f
C7540 ASIG5V.n10237 VSS 0.056945f
C7541 ASIG5V.n10238 VSS 0.056945f
C7542 ASIG5V.n10239 VSS 0.056945f
C7543 ASIG5V.n10240 VSS 0.056945f
C7544 ASIG5V.n10241 VSS 0.056945f
C7545 ASIG5V.n10242 VSS 0.056945f
C7546 ASIG5V.n10243 VSS 0.056945f
C7547 ASIG5V.n10244 VSS 0.056945f
C7548 ASIG5V.n10245 VSS 0.056945f
C7549 ASIG5V.n10246 VSS 0.056945f
C7550 ASIG5V.n10247 VSS 0.056945f
C7551 ASIG5V.n10248 VSS 0.056945f
C7552 ASIG5V.n10249 VSS 0.056945f
C7553 ASIG5V.n10250 VSS 0.056945f
C7554 ASIG5V.n10251 VSS 0.056945f
C7555 ASIG5V.n10252 VSS 0.056945f
C7556 ASIG5V.n10253 VSS 0.056945f
C7557 ASIG5V.n10254 VSS 0.056945f
C7558 ASIG5V.n10255 VSS 0.056945f
C7559 ASIG5V.n10256 VSS 0.056945f
C7560 ASIG5V.n10257 VSS 0.056945f
C7561 ASIG5V.n10258 VSS 0.056945f
C7562 ASIG5V.n10259 VSS 0.056945f
C7563 ASIG5V.n10260 VSS 0.056945f
C7564 ASIG5V.n10261 VSS 0.056945f
C7565 ASIG5V.n10262 VSS 0.056945f
C7566 ASIG5V.n10263 VSS 0.056945f
C7567 ASIG5V.n10264 VSS 0.056945f
C7568 ASIG5V.n10265 VSS 0.056945f
C7569 ASIG5V.n10266 VSS 0.056945f
C7570 ASIG5V.n10267 VSS 0.056945f
C7571 ASIG5V.n10268 VSS 0.056945f
C7572 ASIG5V.n10269 VSS 0.056945f
C7573 ASIG5V.n10270 VSS 0.056945f
C7574 ASIG5V.n10271 VSS 0.056945f
C7575 ASIG5V.n10272 VSS 0.056945f
C7576 ASIG5V.n10273 VSS 0.056945f
C7577 ASIG5V.n10274 VSS 0.056945f
C7578 ASIG5V.n10275 VSS 0.056945f
C7579 ASIG5V.n10276 VSS 0.056945f
C7580 ASIG5V.n10277 VSS 0.056945f
C7581 ASIG5V.n10278 VSS 0.056945f
C7582 ASIG5V.n10279 VSS 0.056945f
C7583 ASIG5V.n10280 VSS 0.056945f
C7584 ASIG5V.n10281 VSS 0.056945f
C7585 ASIG5V.n10282 VSS 0.056945f
C7586 ASIG5V.n10283 VSS 0.056945f
C7587 ASIG5V.n10284 VSS 0.056945f
C7588 ASIG5V.n10285 VSS 0.056945f
C7589 ASIG5V.n10286 VSS 0.056945f
C7590 ASIG5V.n10287 VSS 0.056945f
C7591 ASIG5V.n10288 VSS 0.056945f
C7592 ASIG5V.n10289 VSS 0.056945f
C7593 ASIG5V.n10290 VSS 0.056945f
C7594 ASIG5V.n10291 VSS 0.056945f
C7595 ASIG5V.n10292 VSS 0.056945f
C7596 ASIG5V.n10293 VSS 0.056945f
C7597 ASIG5V.n10294 VSS 0.056945f
C7598 ASIG5V.n10295 VSS 0.056945f
C7599 ASIG5V.n10296 VSS 0.056945f
C7600 ASIG5V.n10297 VSS 0.056945f
C7601 ASIG5V.n10298 VSS 0.056945f
C7602 ASIG5V.n10299 VSS 0.056945f
C7603 ASIG5V.n10300 VSS 0.056945f
C7604 ASIG5V.n10301 VSS 0.056945f
C7605 ASIG5V.n10302 VSS 0.056945f
C7606 ASIG5V.n10303 VSS 0.056945f
C7607 ASIG5V.n10304 VSS 0.056945f
C7608 ASIG5V.n10305 VSS 0.056945f
C7609 ASIG5V.n10306 VSS 0.056945f
C7610 ASIG5V.n10307 VSS 0.056945f
C7611 ASIG5V.n10308 VSS 0.056945f
C7612 ASIG5V.n10309 VSS 0.056945f
C7613 ASIG5V.n10310 VSS 0.056945f
C7614 ASIG5V.n10311 VSS 0.056945f
C7615 ASIG5V.n10312 VSS 0.056945f
C7616 ASIG5V.n10313 VSS 0.056945f
C7617 ASIG5V.n10314 VSS 0.056945f
C7618 ASIG5V.n10315 VSS 0.056945f
C7619 ASIG5V.n10316 VSS 0.056945f
C7620 ASIG5V.n10317 VSS 0.056945f
C7621 ASIG5V.n10318 VSS 0.056945f
C7622 ASIG5V.n10319 VSS 0.056945f
C7623 ASIG5V.n10320 VSS 0.056945f
C7624 ASIG5V.n10321 VSS 0.056945f
C7625 ASIG5V.n10322 VSS 0.056945f
C7626 ASIG5V.n10323 VSS 0.056945f
C7627 ASIG5V.n10324 VSS 0.056945f
C7628 ASIG5V.n10325 VSS 0.056945f
C7629 ASIG5V.n10326 VSS 0.056945f
C7630 ASIG5V.n10327 VSS 0.056945f
C7631 ASIG5V.n10328 VSS 0.056945f
C7632 ASIG5V.n10329 VSS 0.056945f
C7633 ASIG5V.n10330 VSS 0.056945f
C7634 ASIG5V.n10331 VSS 0.056945f
C7635 ASIG5V.n10332 VSS 0.056945f
C7636 ASIG5V.n10333 VSS 0.056945f
C7637 ASIG5V.n10334 VSS 0.056945f
C7638 ASIG5V.n10335 VSS 0.056945f
C7639 ASIG5V.n10336 VSS 0.056945f
C7640 ASIG5V.n10337 VSS 0.056945f
C7641 ASIG5V.n10338 VSS 0.056945f
C7642 ASIG5V.n10339 VSS 0.056945f
C7643 ASIG5V.n10340 VSS 0.056945f
C7644 ASIG5V.n10341 VSS 0.056945f
C7645 ASIG5V.n10342 VSS 0.056945f
C7646 ASIG5V.n10343 VSS 0.056945f
C7647 ASIG5V.n10344 VSS 0.056945f
C7648 ASIG5V.n10345 VSS 0.056945f
C7649 ASIG5V.n10346 VSS 0.056945f
C7650 ASIG5V.n10347 VSS 0.056945f
C7651 ASIG5V.n10348 VSS 0.056945f
C7652 ASIG5V.n10349 VSS 0.056945f
C7653 ASIG5V.n10350 VSS 0.056945f
C7654 ASIG5V.n10351 VSS 0.056945f
C7655 ASIG5V.n10352 VSS 0.056945f
C7656 ASIG5V.n10353 VSS 0.056945f
C7657 ASIG5V.n10354 VSS 0.056945f
C7658 ASIG5V.n10356 VSS 0.701152f
C7659 ASIG5V.n10358 VSS 0.056945f
C7660 ASIG5V.n10359 VSS 0.056945f
C7661 ASIG5V.n10360 VSS 0.056945f
C7662 ASIG5V.n10361 VSS 0.056945f
C7663 ASIG5V.n10362 VSS 0.047722f
C7664 ASIG5V.n10363 VSS 0.05375f
C7665 ASIG5V.n10364 VSS 0.05375f
C7666 ASIG5V.n10365 VSS 0.076709f
C7667 ASIG5V.n10366 VSS 0.061313f
C7668 ASIG5V.n10367 VSS 0.046943f
C7669 ASIG5V.n10368 VSS 0.052746f
C7670 ASIG5V.n10369 VSS 0.052746f
C7671 ASIG5V.n10370 VSS 0.045974f
C7672 ASIG5V.n10371 VSS 0.076709f
C7673 ASIG5V.n10372 VSS 0.045974f
C7674 ASIG5V.n10373 VSS 0.323607f
C7675 ASIG5V.n10415 VSS 0.036092f
C7676 ASIG5V.n10416 VSS 0.323607f
C7677 ASIG5V.n10418 VSS 0.056945f
C7678 ASIG5V.n10419 VSS 0.056945f
C7679 ASIG5V.n10420 VSS 0.056945f
C7680 ASIG5V.n10421 VSS 0.056945f
C7681 ASIG5V.n10422 VSS 0.056945f
C7682 ASIG5V.n10423 VSS 0.793611f
C7683 ASIG5V.n10463 VSS 0.036092f
C7684 ASIG5V.n10464 VSS 0.056945f
C7685 ASIG5V.n10465 VSS 0.056945f
C7686 ASIG5V.n10466 VSS 0.069023f
C7687 ASIG5V.n10467 VSS 0.09726f
C7688 ASIG5V.n10468 VSS 0.0621f
C7689 ASIG5V.n10469 VSS 0.108961f
C7690 ASIG5V.n10470 VSS 0.108961f
C7691 ASIG5V.n10471 VSS 0.97853f
C7692 ASIG5V.n10472 VSS 1.07099f
C7693 ASIG5V.n10473 VSS 0.098416f
C7694 ASIG5V.n10474 VSS 0.098416f
C7695 ASIG5V.n10475 VSS 0.087848f
C7696 ASIG5V.n10476 VSS 0.09726f
C7697 ASIG5V.n10477 VSS 0.108961f
C7698 ASIG5V.n10478 VSS 0.077327f
C7699 ASIG5V.n10479 VSS 0.077327f
C7700 ASIG5V.n10480 VSS 0.0621f
C7701 ASIG5V.n10481 VSS 0.106324f
C7702 ASIG5V.n10482 VSS 0.955415f
C7703 ASIG5V.n10483 VSS 1.0941f
C7704 ASIG5V.n10484 VSS 0.068336f
C7705 ASIG5V.n10485 VSS 0.049969f
C7706 ASIG5V.n10486 VSS 0.068336f
C7707 ASIG5V.n10487 VSS 0.049969f
C7708 ASIG5V.n10488 VSS 0.059682f
C7709 ASIG5V.n10489 VSS 0.106625f
C7710 ASIG5V.n10490 VSS 0.070117f
C7711 ASIG5V.n10491 VSS 0.070117f
C7712 ASIG5V.n10492 VSS 0.955416f
C7713 ASIG5V.n10493 VSS 0.955416f
C7714 ASIG5V.n10494 VSS 2.43477f
C7715 ASIG5V.n10495 VSS 0.955416f
C7716 ASIG5V.n10496 VSS 1.20198f
C7717 ASIG5V.n10497 VSS 0.161825f
C7718 ASIG5V.n10498 VSS 0.117005f
C7719 ASIG5V.n10499 VSS 0.117005f
C7720 ASIG5V.n10500 VSS 0.117005f
C7721 ASIG5V.n10501 VSS 0.117005f
C7722 ASIG5V.n10502 VSS 0.117005f
C7723 ASIG5V.n10503 VSS 0.117005f
C7724 ASIG5V.n10504 VSS 0.117005f
C7725 ASIG5V.n10505 VSS 0.117005f
C7726 ASIG5V.n10506 VSS 0.117005f
C7727 ASIG5V.n10507 VSS 0.117005f
C7728 ASIG5V.n10508 VSS 0.117005f
C7729 ASIG5V.n10509 VSS 0.117005f
C7730 ASIG5V.n10510 VSS 0.117005f
C7731 ASIG5V.n10511 VSS 0.117005f
C7732 ASIG5V.n10512 VSS 0.117005f
C7733 ASIG5V.n10513 VSS 0.117005f
C7734 ASIG5V.n10514 VSS 0.117005f
C7735 ASIG5V.n10515 VSS 0.117005f
C7736 ASIG5V.n10516 VSS 0.117005f
C7737 ASIG5V.n10517 VSS 0.117005f
C7738 ASIG5V.n10518 VSS 0.117005f
C7739 ASIG5V.n10519 VSS 0.117005f
C7740 ASIG5V.n10520 VSS 0.117005f
C7741 ASIG5V.n10521 VSS 0.117005f
C7742 ASIG5V.n10522 VSS 0.117005f
C7743 ASIG5V.n10523 VSS 0.117005f
C7744 ASIG5V.n10524 VSS 0.117005f
C7745 ASIG5V.n10525 VSS 0.117005f
C7746 ASIG5V.n10526 VSS 0.117005f
C7747 ASIG5V.n10527 VSS 0.117005f
C7748 ASIG5V.n10528 VSS 0.117005f
C7749 ASIG5V.n10529 VSS 0.117005f
C7750 ASIG5V.n10530 VSS 0.117005f
C7751 ASIG5V.n10531 VSS 0.117005f
C7752 ASIG5V.n10532 VSS 0.117005f
C7753 ASIG5V.n10533 VSS 0.117005f
C7754 ASIG5V.n10534 VSS 0.117005f
C7755 ASIG5V.n10535 VSS 0.117005f
C7756 ASIG5V.n10536 VSS 0.117005f
C7757 ASIG5V.n10537 VSS 0.117005f
C7758 ASIG5V.n10538 VSS 0.117005f
C7759 ASIG5V.n10539 VSS 0.117005f
C7760 ASIG5V.n10540 VSS 0.117005f
C7761 ASIG5V.n10541 VSS 0.117005f
C7762 ASIG5V.n10542 VSS 0.117005f
C7763 ASIG5V.n10543 VSS 0.117005f
C7764 ASIG5V.n10544 VSS 0.117005f
C7765 ASIG5V.n10545 VSS 0.117005f
C7766 ASIG5V.n10546 VSS 0.955416f
C7767 ASIG5V.n10548 VSS 0.092943f
C7768 ASIG5V.n10551 VSS 0.117005f
C7769 ASIG5V.n10554 VSS 0.117005f
C7770 ASIG5V.n10557 VSS 0.117005f
C7771 ASIG5V.n10560 VSS 0.117005f
C7772 ASIG5V.n10563 VSS 0.117005f
C7773 ASIG5V.n10566 VSS 0.117005f
C7774 ASIG5V.n10569 VSS 0.117005f
C7775 ASIG5V.n10572 VSS 0.117005f
C7776 ASIG5V.n10575 VSS 0.117005f
C7777 ASIG5V.n10578 VSS 0.117005f
C7778 ASIG5V.n10581 VSS 0.117005f
C7779 ASIG5V.n10584 VSS 0.117005f
C7780 ASIG5V.n10587 VSS 0.117005f
C7781 ASIG5V.n10590 VSS 0.117005f
C7782 ASIG5V.n10593 VSS 0.117005f
C7783 ASIG5V.n10596 VSS 0.117005f
C7784 ASIG5V.n10599 VSS 0.117005f
C7785 ASIG5V.n10602 VSS 0.117005f
C7786 ASIG5V.n10605 VSS 0.117005f
C7787 ASIG5V.n10608 VSS 0.117005f
C7788 ASIG5V.n10611 VSS 0.117005f
C7789 ASIG5V.n10614 VSS 0.117005f
C7790 ASIG5V.n10617 VSS 0.117005f
C7791 ASIG5V.n10620 VSS 0.117005f
C7792 ASIG5V.n10623 VSS 0.117005f
C7793 ASIG5V.n10626 VSS 0.117005f
C7794 ASIG5V.n10629 VSS 0.117005f
C7795 ASIG5V.n10632 VSS 0.117005f
C7796 ASIG5V.n10635 VSS 0.117005f
C7797 ASIG5V.n10638 VSS 0.117005f
C7798 ASIG5V.n10641 VSS 0.117005f
C7799 ASIG5V.n10644 VSS 0.117005f
C7800 ASIG5V.n10647 VSS 0.117005f
C7801 ASIG5V.n10650 VSS 0.117005f
C7802 ASIG5V.n10653 VSS 0.117005f
C7803 ASIG5V.n10656 VSS 0.117005f
C7804 ASIG5V.n10659 VSS 0.117005f
C7805 ASIG5V.n10662 VSS 0.117005f
C7806 ASIG5V.n10665 VSS 0.117005f
C7807 ASIG5V.n10668 VSS 0.117005f
C7808 ASIG5V.n10671 VSS 0.117005f
C7809 ASIG5V.n10674 VSS 0.117005f
C7810 ASIG5V.n10677 VSS 0.117005f
C7811 ASIG5V.n10680 VSS 0.117005f
C7812 ASIG5V.n10683 VSS 0.117005f
C7813 ASIG5V.n10686 VSS 0.117005f
C7814 ASIG5V.n10689 VSS 0.117005f
C7815 ASIG5V.n10692 VSS 0.161825f
C7816 ASIG5V.n10693 VSS 0.086338f
C7817 ASIG5V.n10694 VSS 0.067466f
C7818 ASIG5V.n10697 VSS 0.955416f
C7819 ASIG5V.n10698 VSS 0.108041f
C7820 ASIG5V.n10699 VSS 0.110346f
C7821 ASIG5V.n10700 VSS 0.067466f
C7822 ASIG5V.n10701 VSS 0.955416f
C7823 ASIG5V.n10703 VSS 0.955415f
C7824 ASIG5V.n10704 VSS 1.33296f
C7825 ASIG5V.n10705 VSS 0.108041f
C7826 ASIG5V.n10706 VSS 0.110346f
C7827 ASIG5V.n10707 VSS 0.106324f
C7828 ASIG5V.n10708 VSS 0.094907f
C7829 ASIG5V.n10709 VSS 0.379429f
C7830 ASIG5V.n10710 VSS 0.201323f
C7831 ASIG5V.n10711 VSS 0.196332f
C7832 ASIG5V.n10712 VSS 0.955416f
C7833 ASIG5V.n10713 VSS 0.161825f
C7834 ASIG5V.n10714 VSS 0.161825f
C7835 ASIG5V.n10715 VSS 0.161825f
C7836 ASIG5V.n10716 VSS 0.161825f
C7837 ASIG5V.n10717 VSS 0.117005f
C7838 ASIG5V.n10718 VSS 0.117005f
C7839 ASIG5V.n10719 VSS 0.117005f
C7840 ASIG5V.n10720 VSS 0.117005f
C7841 ASIG5V.n10721 VSS 0.117005f
C7842 ASIG5V.n10722 VSS 0.117005f
C7843 ASIG5V.n10723 VSS 0.117005f
C7844 ASIG5V.n10724 VSS 0.117005f
C7845 ASIG5V.n10725 VSS 0.117005f
C7846 ASIG5V.n10726 VSS 0.117005f
C7847 ASIG5V.n10727 VSS 0.117005f
C7848 ASIG5V.n10728 VSS 0.117005f
C7849 ASIG5V.n10729 VSS 0.117005f
C7850 ASIG5V.n10730 VSS 0.117005f
C7851 ASIG5V.n10731 VSS 0.117005f
C7852 ASIG5V.n10732 VSS 0.117005f
C7853 ASIG5V.n10733 VSS 0.117005f
C7854 ASIG5V.n10734 VSS 0.117005f
C7855 ASIG5V.n10735 VSS 0.117005f
C7856 ASIG5V.n10736 VSS 0.117005f
C7857 ASIG5V.n10737 VSS 0.117005f
C7858 ASIG5V.n10738 VSS 0.117005f
C7859 ASIG5V.n10739 VSS 0.117005f
C7860 ASIG5V.n10740 VSS 0.117005f
C7861 ASIG5V.n10741 VSS 0.117005f
C7862 ASIG5V.n10742 VSS 0.117005f
C7863 ASIG5V.n10743 VSS 0.117005f
C7864 ASIG5V.n10744 VSS 0.117005f
C7865 ASIG5V.n10745 VSS 0.117005f
C7866 ASIG5V.n10746 VSS 0.117005f
C7867 ASIG5V.n10747 VSS 0.117005f
C7868 ASIG5V.n10748 VSS 0.117005f
C7869 ASIG5V.n10749 VSS 0.117005f
C7870 ASIG5V.n10750 VSS 0.117005f
C7871 ASIG5V.n10751 VSS 0.117005f
C7872 ASIG5V.n10752 VSS 0.117005f
C7873 ASIG5V.n10753 VSS 0.117005f
C7874 ASIG5V.n10754 VSS 0.117005f
C7875 ASIG5V.n10755 VSS 0.117005f
C7876 ASIG5V.n10756 VSS 0.117005f
C7877 ASIG5V.n10757 VSS 0.117005f
C7878 ASIG5V.n10758 VSS 0.117005f
C7879 ASIG5V.n10759 VSS 0.117005f
C7880 ASIG5V.n10760 VSS 0.117005f
C7881 ASIG5V.n10761 VSS 0.117005f
C7882 ASIG5V.n10762 VSS 0.117005f
C7883 ASIG5V.n10763 VSS 0.117005f
C7884 ASIG5V.n10764 VSS 0.117005f
C7885 ASIG5V.n10765 VSS 0.117005f
C7886 ASIG5V.n10766 VSS 0.117005f
C7887 ASIG5V.n10767 VSS 0.117005f
C7888 ASIG5V.n10768 VSS 0.117005f
C7889 ASIG5V.n10769 VSS 0.117005f
C7890 ASIG5V.n10770 VSS 0.117005f
C7891 ASIG5V.n10771 VSS 0.117005f
C7892 ASIG5V.n10772 VSS 0.117005f
C7893 ASIG5V.n10773 VSS 0.117005f
C7894 ASIG5V.n10774 VSS 0.117005f
C7895 ASIG5V.n10775 VSS 0.117005f
C7896 ASIG5V.n10776 VSS 0.117005f
C7897 ASIG5V.n10777 VSS 0.117005f
C7898 ASIG5V.n10778 VSS 0.117005f
C7899 ASIG5V.n10779 VSS 0.117005f
C7900 ASIG5V.n10780 VSS 0.117005f
C7901 ASIG5V.n10781 VSS 0.117005f
C7902 ASIG5V.n10782 VSS 0.117005f
C7903 ASIG5V.n10783 VSS 0.117005f
C7904 ASIG5V.n10784 VSS 0.117005f
C7905 ASIG5V.n10785 VSS 0.117005f
C7906 ASIG5V.n10786 VSS 0.117005f
C7907 ASIG5V.n10787 VSS 0.117005f
C7908 ASIG5V.n10788 VSS 0.117005f
C7909 ASIG5V.n10789 VSS 0.117005f
C7910 ASIG5V.n10790 VSS 0.117005f
C7911 ASIG5V.n10791 VSS 0.117005f
C7912 ASIG5V.n10792 VSS 0.117005f
C7913 ASIG5V.n10793 VSS 0.117005f
C7914 ASIG5V.n10794 VSS 0.117005f
C7915 ASIG5V.n10795 VSS 0.117005f
C7916 ASIG5V.n10796 VSS 0.117005f
C7917 ASIG5V.n10797 VSS 0.117005f
C7918 ASIG5V.n10798 VSS 0.117005f
C7919 ASIG5V.n10799 VSS 0.117005f
C7920 ASIG5V.n10800 VSS 0.117005f
C7921 ASIG5V.n10801 VSS 0.117005f
C7922 ASIG5V.n10802 VSS 0.117005f
C7923 ASIG5V.n10803 VSS 0.117005f
C7924 ASIG5V.n10804 VSS 0.117005f
C7925 ASIG5V.n10805 VSS 0.117005f
C7926 ASIG5V.n10806 VSS 0.117005f
C7927 ASIG5V.n10807 VSS 0.117005f
C7928 ASIG5V.n10808 VSS 0.117005f
C7929 ASIG5V.n10809 VSS 0.117005f
C7930 ASIG5V.n10810 VSS 0.117005f
C7931 ASIG5V.n10811 VSS 0.117005f
C7932 ASIG5V.n10812 VSS 0.117005f
C7933 ASIG5V.n10813 VSS 0.092943f
C7934 ASIG5V.n10814 VSS 0.117005f
C7935 ASIG5V.n10815 VSS 0.117005f
C7936 ASIG5V.n10816 VSS 0.117005f
C7937 ASIG5V.n10817 VSS 0.117005f
C7938 ASIG5V.n10818 VSS 0.117005f
C7939 ASIG5V.n10819 VSS 0.117005f
C7940 ASIG5V.n10820 VSS 0.117005f
C7941 ASIG5V.n10821 VSS 0.117005f
C7942 ASIG5V.n10822 VSS 0.117005f
C7943 ASIG5V.n10823 VSS 0.117005f
C7944 ASIG5V.n10824 VSS 0.117005f
C7945 ASIG5V.n10825 VSS 0.117005f
C7946 ASIG5V.n10826 VSS 0.117005f
C7947 ASIG5V.n10827 VSS 0.117005f
C7948 ASIG5V.n10828 VSS 0.117005f
C7949 ASIG5V.n10829 VSS 0.117005f
C7950 ASIG5V.n10830 VSS 0.117005f
C7951 ASIG5V.n10831 VSS 0.117005f
C7952 ASIG5V.n10832 VSS 0.117005f
C7953 ASIG5V.n10833 VSS 0.117005f
C7954 ASIG5V.n10834 VSS 0.117005f
C7955 ASIG5V.n10835 VSS 0.117005f
C7956 ASIG5V.n10836 VSS 0.117005f
C7957 ASIG5V.n10837 VSS 0.117005f
C7958 ASIG5V.n10838 VSS 0.117005f
C7959 ASIG5V.n10839 VSS 0.117005f
C7960 ASIG5V.n10840 VSS 0.117005f
C7961 ASIG5V.n10841 VSS 0.117005f
C7962 ASIG5V.n10842 VSS 0.117005f
C7963 ASIG5V.n10843 VSS 0.117005f
C7964 ASIG5V.n10844 VSS 0.117005f
C7965 ASIG5V.n10845 VSS 0.117005f
C7966 ASIG5V.n10846 VSS 0.117005f
C7967 ASIG5V.n10847 VSS 0.117005f
C7968 ASIG5V.n10848 VSS 0.117005f
C7969 ASIG5V.n10849 VSS 0.117005f
C7970 ASIG5V.n10850 VSS 0.117005f
C7971 ASIG5V.n10851 VSS 0.117005f
C7972 ASIG5V.n10852 VSS 0.117005f
C7973 ASIG5V.n10853 VSS 0.117005f
C7974 ASIG5V.n10854 VSS 0.117005f
C7975 ASIG5V.n10855 VSS 0.117005f
C7976 ASIG5V.n10856 VSS 0.117005f
C7977 ASIG5V.n10857 VSS 0.117005f
C7978 ASIG5V.n10858 VSS 0.117005f
C7979 ASIG5V.n10859 VSS 0.117005f
C7980 ASIG5V.n10860 VSS 0.117005f
C7981 ASIG5V.n10861 VSS 0.117005f
C7982 ASIG5V.n10862 VSS 0.117005f
C7983 ASIG5V.n10863 VSS 0.117005f
C7984 ASIG5V.n10864 VSS 0.117005f
C7985 ASIG5V.n10865 VSS 0.117005f
C7986 ASIG5V.n10866 VSS 0.117005f
C7987 ASIG5V.n10867 VSS 0.117005f
C7988 ASIG5V.n10868 VSS 0.117005f
C7989 ASIG5V.n10869 VSS 0.117005f
C7990 ASIG5V.n10870 VSS 0.117005f
C7991 ASIG5V.n10871 VSS 0.117005f
C7992 ASIG5V.n10872 VSS 0.117005f
C7993 ASIG5V.n10873 VSS 0.117005f
C7994 ASIG5V.n10874 VSS 0.117005f
C7995 ASIG5V.n10875 VSS 0.117005f
C7996 ASIG5V.n10876 VSS 0.117005f
C7997 ASIG5V.n10877 VSS 0.117005f
C7998 ASIG5V.n10878 VSS 0.117005f
C7999 ASIG5V.n10879 VSS 0.117005f
C8000 ASIG5V.n10880 VSS 0.117005f
C8001 ASIG5V.n10881 VSS 0.117005f
C8002 ASIG5V.n10882 VSS 0.117005f
C8003 ASIG5V.n10883 VSS 0.117005f
C8004 ASIG5V.n10884 VSS 0.117005f
C8005 ASIG5V.n10885 VSS 0.117005f
C8006 ASIG5V.n10886 VSS 0.117005f
C8007 ASIG5V.n10887 VSS 0.117005f
C8008 ASIG5V.n10888 VSS 0.117005f
C8009 ASIG5V.n10889 VSS 0.117005f
C8010 ASIG5V.n10890 VSS 0.117005f
C8011 ASIG5V.n10891 VSS 0.117005f
C8012 ASIG5V.n10892 VSS 0.117005f
C8013 ASIG5V.n10893 VSS 0.117005f
C8014 ASIG5V.n10894 VSS 0.117005f
C8015 ASIG5V.n10895 VSS 0.117005f
C8016 ASIG5V.n10896 VSS 0.117005f
C8017 ASIG5V.n10897 VSS 0.117005f
C8018 ASIG5V.n10898 VSS 0.117005f
C8019 ASIG5V.n10899 VSS 0.117005f
C8020 ASIG5V.n10900 VSS 0.117005f
C8021 ASIG5V.n10901 VSS 0.117005f
C8022 ASIG5V.n10902 VSS 0.117005f
C8023 ASIG5V.n10903 VSS 0.117005f
C8024 ASIG5V.n10904 VSS 0.117005f
C8025 ASIG5V.n10905 VSS 0.117005f
C8026 ASIG5V.n10906 VSS 0.117005f
C8027 ASIG5V.n10907 VSS 0.117005f
C8028 ASIG5V.n10908 VSS 0.117005f
C8029 ASIG5V.n10909 VSS 0.117005f
C8030 ASIG5V.n10910 VSS 0.117005f
C8031 ASIG5V.n10911 VSS 0.955416f
C8032 ASIG5V.n10912 VSS 0.19202f
C8033 ASIG5V.n10913 VSS 0.192509f
C8034 ASIG5V.n10914 VSS 0.246495f
C8035 ASIG5V.n10915 VSS 0.043641f
C8036 ASIG5V.n10916 VSS 0.066995f
C8037 ASIG5V.n10917 VSS 0.076709f
C8038 ASIG5V.n10918 VSS 0.076709f
C8039 ASIG5V.n10919 VSS 0.955415f
C8040 ASIG5V.n10920 VSS 1.0941f
C8041 ASIG5V.n10921 VSS 0.108961f
C8042 ASIG5V.n10922 VSS 0.086114f
C8043 ASIG5V.n10923 VSS 0.086114f
C8044 ASIG5V.n10924 VSS 0.076867f
C8045 ASIG5V.n10925 VSS 0.07229f
C8046 ASIG5V.n10926 VSS 0.052133f
C8047 ASIG5V.n10927 VSS 0.056945f
C8048 ASIG5V.n10928 VSS 0.056945f
C8049 ASIG5V.n10929 VSS 0.056945f
C8050 ASIG5V.n10930 VSS 0.056945f
C8051 ASIG5V.n10931 VSS 0.056945f
C8052 ASIG5V.n10932 VSS 0.056945f
C8053 ASIG5V.n10933 VSS 0.056945f
C8054 ASIG5V.n10934 VSS 0.056945f
C8055 ASIG5V.n10935 VSS 0.056945f
C8056 ASIG5V.n10936 VSS 0.056945f
C8057 ASIG5V.n10937 VSS 0.056945f
C8058 ASIG5V.n10938 VSS 0.056945f
C8059 ASIG5V.n10939 VSS 0.056945f
C8060 ASIG5V.n10940 VSS 0.056945f
C8061 ASIG5V.n10941 VSS 0.056945f
C8062 ASIG5V.n10942 VSS 0.056945f
C8063 ASIG5V.n10943 VSS 0.056945f
C8064 ASIG5V.n10944 VSS 0.056945f
C8065 ASIG5V.n10945 VSS 0.056945f
C8066 ASIG5V.n10946 VSS 0.056945f
C8067 ASIG5V.n10947 VSS 0.056945f
C8068 ASIG5V.n10948 VSS 0.056945f
C8069 ASIG5V.n10949 VSS 0.056945f
C8070 ASIG5V.n10950 VSS 0.056945f
C8071 ASIG5V.n10951 VSS 0.056945f
C8072 ASIG5V.n10952 VSS 0.056945f
C8073 ASIG5V.n10953 VSS 0.056945f
C8074 ASIG5V.n10954 VSS 0.056945f
C8075 ASIG5V.n10955 VSS 0.056945f
C8076 ASIG5V.n10956 VSS 0.056945f
C8077 ASIG5V.n10957 VSS 0.056945f
C8078 ASIG5V.n10958 VSS 0.056945f
C8079 ASIG5V.n10959 VSS 0.056945f
C8080 ASIG5V.n10960 VSS 0.056945f
C8081 ASIG5V.n10961 VSS 0.056945f
C8082 ASIG5V.n10962 VSS 0.056945f
C8083 ASIG5V.n10963 VSS 0.056945f
C8084 ASIG5V.n10964 VSS 0.056945f
C8085 ASIG5V.n10965 VSS 0.056945f
C8086 ASIG5V.n10966 VSS 0.056945f
C8087 ASIG5V.n10967 VSS 0.056945f
C8088 ASIG5V.n10968 VSS 0.056945f
C8089 ASIG5V.n10969 VSS 0.056945f
C8090 ASIG5V.n10970 VSS 0.056945f
C8091 ASIG5V.n10971 VSS 0.056945f
C8092 ASIG5V.n10972 VSS 0.056945f
C8093 ASIG5V.n10973 VSS 0.056945f
C8094 ASIG5V.n10974 VSS 0.056945f
C8095 ASIG5V.n10975 VSS 0.056945f
C8096 ASIG5V.n10976 VSS 0.056945f
C8097 ASIG5V.n10977 VSS 0.056945f
C8098 ASIG5V.n10978 VSS 0.056945f
C8099 ASIG5V.n10979 VSS 0.056945f
C8100 ASIG5V.n10980 VSS 0.056945f
C8101 ASIG5V.n10981 VSS 0.056945f
C8102 ASIG5V.n10982 VSS 0.056945f
C8103 ASIG5V.n10983 VSS 0.056945f
C8104 ASIG5V.n10984 VSS 0.056945f
C8105 ASIG5V.n10985 VSS 0.056945f
C8106 ASIG5V.n10986 VSS 0.056945f
C8107 ASIG5V.n10987 VSS 0.056945f
C8108 ASIG5V.n10988 VSS 0.056945f
C8109 ASIG5V.n10989 VSS 0.056945f
C8110 ASIG5V.n10990 VSS 0.056945f
C8111 ASIG5V.n10991 VSS 0.056945f
C8112 ASIG5V.n10992 VSS 0.056945f
C8113 ASIG5V.n10993 VSS 0.056945f
C8114 ASIG5V.n10994 VSS 0.056945f
C8115 ASIG5V.n10995 VSS 0.056945f
C8116 ASIG5V.n10996 VSS 0.056945f
C8117 ASIG5V.n10997 VSS 0.056945f
C8118 ASIG5V.n10998 VSS 0.056945f
C8119 ASIG5V.n10999 VSS 0.056945f
C8120 ASIG5V.n11000 VSS 0.056945f
C8121 ASIG5V.n11001 VSS 0.056945f
C8122 ASIG5V.n11002 VSS 0.056945f
C8123 ASIG5V.n11003 VSS 0.056945f
C8124 ASIG5V.n11004 VSS 0.056945f
C8125 ASIG5V.n11005 VSS 0.056945f
C8126 ASIG5V.n11006 VSS 0.056945f
C8127 ASIG5V.n11007 VSS 0.056945f
C8128 ASIG5V.n11008 VSS 0.056945f
C8129 ASIG5V.n11009 VSS 0.056945f
C8130 ASIG5V.n11010 VSS 0.056945f
C8131 ASIG5V.n11011 VSS 0.056945f
C8132 ASIG5V.n11012 VSS 0.056945f
C8133 ASIG5V.n11013 VSS 0.056945f
C8134 ASIG5V.n11014 VSS 0.056945f
C8135 ASIG5V.n11015 VSS 0.056945f
C8136 ASIG5V.n11016 VSS 0.056945f
C8137 ASIG5V.n11017 VSS 0.056945f
C8138 ASIG5V.n11018 VSS 0.056945f
C8139 ASIG5V.n11019 VSS 0.056945f
C8140 ASIG5V.n11020 VSS 0.056945f
C8141 ASIG5V.n11021 VSS 0.056945f
C8142 ASIG5V.n11022 VSS 0.056945f
C8143 ASIG5V.n11023 VSS 0.056945f
C8144 ASIG5V.n11024 VSS 0.056945f
C8145 ASIG5V.n11025 VSS 0.056945f
C8146 ASIG5V.n11026 VSS 0.056945f
C8147 ASIG5V.n11027 VSS 0.056945f
C8148 ASIG5V.n11028 VSS 0.056945f
C8149 ASIG5V.n11029 VSS 0.056945f
C8150 ASIG5V.n11030 VSS 0.056945f
C8151 ASIG5V.n11031 VSS 0.056945f
C8152 ASIG5V.n11032 VSS 0.056945f
C8153 ASIG5V.n11033 VSS 0.056945f
C8154 ASIG5V.n11034 VSS 0.056945f
C8155 ASIG5V.n11035 VSS 0.056945f
C8156 ASIG5V.n11036 VSS 0.056945f
C8157 ASIG5V.n11037 VSS 0.056945f
C8158 ASIG5V.n11038 VSS 0.056945f
C8159 ASIG5V.n11039 VSS 0.056945f
C8160 ASIG5V.n11040 VSS 0.056945f
C8161 ASIG5V.n11041 VSS 0.056945f
C8162 ASIG5V.n11042 VSS 0.056945f
C8163 ASIG5V.n11043 VSS 0.056945f
C8164 ASIG5V.n11044 VSS 0.056945f
C8165 ASIG5V.n11045 VSS 0.056945f
C8166 ASIG5V.n11046 VSS 0.056945f
C8167 ASIG5V.n11047 VSS 0.056945f
C8168 ASIG5V.n11048 VSS 0.056945f
C8169 ASIG5V.n11049 VSS 0.056945f
C8170 ASIG5V.n11050 VSS 0.056945f
C8171 ASIG5V.n11051 VSS 0.056945f
C8172 ASIG5V.n11052 VSS 0.056945f
C8173 ASIG5V.n11053 VSS 0.056945f
C8174 ASIG5V.n11054 VSS 0.056945f
C8175 ASIG5V.n11055 VSS 0.056945f
C8176 ASIG5V.n11056 VSS 0.056945f
C8177 ASIG5V.n11057 VSS 0.056945f
C8178 ASIG5V.n11058 VSS 0.056945f
C8179 ASIG5V.n11059 VSS 0.056945f
C8180 ASIG5V.n11060 VSS 0.056945f
C8181 ASIG5V.n11061 VSS 0.056945f
C8182 ASIG5V.n11062 VSS 0.056945f
C8183 ASIG5V.n11063 VSS 0.056945f
C8184 ASIG5V.n11064 VSS 0.056945f
C8185 ASIG5V.n11065 VSS 0.056945f
C8186 ASIG5V.n11066 VSS 0.056945f
C8187 ASIG5V.n11067 VSS 0.056945f
C8188 ASIG5V.n11068 VSS 0.056945f
C8189 ASIG5V.n11069 VSS 0.056945f
C8190 ASIG5V.n11070 VSS 0.056945f
C8191 ASIG5V.n11071 VSS 0.056945f
C8192 ASIG5V.n11072 VSS 0.056945f
C8193 ASIG5V.n11073 VSS 0.056945f
C8194 ASIG5V.n11074 VSS 0.056945f
C8195 ASIG5V.n11075 VSS 0.056945f
C8196 ASIG5V.n11076 VSS 0.056945f
C8197 ASIG5V.n11077 VSS 0.056945f
C8198 ASIG5V.n11078 VSS 0.056945f
C8199 ASIG5V.n11079 VSS 0.056945f
C8200 ASIG5V.n11080 VSS 0.056945f
C8201 ASIG5V.n11081 VSS 0.056945f
C8202 ASIG5V.n11082 VSS 0.056945f
C8203 ASIG5V.n11083 VSS 0.056945f
C8204 ASIG5V.n11084 VSS 0.056945f
C8205 ASIG5V.n11085 VSS 0.056945f
C8206 ASIG5V.n11086 VSS 0.056945f
C8207 ASIG5V.n11087 VSS 0.056945f
C8208 ASIG5V.n11088 VSS 0.056945f
C8209 ASIG5V.n11089 VSS 0.056945f
C8210 ASIG5V.n11090 VSS 0.056945f
C8211 ASIG5V.n11091 VSS 0.056945f
C8212 ASIG5V.n11092 VSS 0.056945f
C8213 ASIG5V.n11093 VSS 0.056945f
C8214 ASIG5V.n11094 VSS 0.056945f
C8215 ASIG5V.n11095 VSS 0.056945f
C8216 ASIG5V.n11096 VSS 0.056945f
C8217 ASIG5V.n11097 VSS 0.056945f
C8218 ASIG5V.n11098 VSS 0.056945f
C8219 ASIG5V.n11099 VSS 0.056945f
C8220 ASIG5V.n11100 VSS 0.056945f
C8221 ASIG5V.n11101 VSS 0.056945f
C8222 ASIG5V.n11102 VSS 0.056945f
C8223 ASIG5V.n11103 VSS 0.056945f
C8224 ASIG5V.n11104 VSS 0.056945f
C8225 ASIG5V.n11105 VSS 0.056945f
C8226 ASIG5V.n11106 VSS 0.056945f
C8227 ASIG5V.n11107 VSS 0.056945f
C8228 ASIG5V.n11108 VSS 0.056945f
C8229 ASIG5V.n11109 VSS 0.056945f
C8230 ASIG5V.n11110 VSS 0.056945f
C8231 ASIG5V.n11111 VSS 0.056945f
C8232 ASIG5V.n11112 VSS 0.056945f
C8233 ASIG5V.n11113 VSS 0.056945f
C8234 ASIG5V.n11114 VSS 0.056945f
C8235 ASIG5V.n11115 VSS 0.056945f
C8236 ASIG5V.n11116 VSS 0.056945f
C8237 ASIG5V.n11117 VSS 0.056945f
C8238 ASIG5V.n11118 VSS 0.056945f
C8239 ASIG5V.n11119 VSS 0.056945f
C8240 ASIG5V.n11120 VSS 0.056945f
C8241 ASIG5V.n11121 VSS 0.056945f
C8242 ASIG5V.n11122 VSS 0.056945f
C8243 ASIG5V.n11123 VSS 0.056945f
C8244 ASIG5V.n11124 VSS 0.056945f
C8245 ASIG5V.n11125 VSS 0.056945f
C8246 ASIG5V.n11126 VSS 0.056945f
C8247 ASIG5V.n11127 VSS 0.056945f
C8248 ASIG5V.n11128 VSS 0.056945f
C8249 ASIG5V.n11129 VSS 0.056945f
C8250 ASIG5V.n11130 VSS 0.056945f
C8251 ASIG5V.n11131 VSS 0.056945f
C8252 ASIG5V.n11132 VSS 0.056945f
C8253 ASIG5V.n11133 VSS 0.056945f
C8254 ASIG5V.n11134 VSS 0.056945f
C8255 ASIG5V.n11135 VSS 0.056945f
C8256 ASIG5V.n11136 VSS 0.056945f
C8257 ASIG5V.n11137 VSS 0.056945f
C8258 ASIG5V.n11138 VSS 0.056945f
C8259 ASIG5V.n11139 VSS 0.056945f
C8260 ASIG5V.n11140 VSS 0.056945f
C8261 ASIG5V.n11141 VSS 0.056945f
C8262 ASIG5V.n11142 VSS 0.056945f
C8263 ASIG5V.n11143 VSS 0.056945f
C8264 ASIG5V.n11144 VSS 0.056945f
C8265 ASIG5V.n11145 VSS 0.056945f
C8266 ASIG5V.n11146 VSS 0.056945f
C8267 ASIG5V.n11147 VSS 0.056945f
C8268 ASIG5V.n11148 VSS 0.056945f
C8269 ASIG5V.n11149 VSS 0.056945f
C8270 ASIG5V.n11150 VSS 0.056945f
C8271 ASIG5V.n11151 VSS 0.056945f
C8272 ASIG5V.n11152 VSS 0.056945f
C8273 ASIG5V.n11153 VSS 0.056945f
C8274 ASIG5V.n11154 VSS 0.056945f
C8275 ASIG5V.n11155 VSS 0.056945f
C8276 ASIG5V.n11156 VSS 0.056945f
C8277 ASIG5V.n11157 VSS 0.056945f
C8278 ASIG5V.n11158 VSS 0.056945f
C8279 ASIG5V.n11159 VSS 0.056945f
C8280 ASIG5V.n11160 VSS 0.056945f
C8281 ASIG5V.n11161 VSS 0.056945f
C8282 ASIG5V.n11163 VSS 0.932301f
C8283 ASIG5V.n11165 VSS 0.056945f
C8284 ASIG5V.n11166 VSS 0.056945f
C8285 ASIG5V.n11167 VSS 0.056945f
C8286 ASIG5V.n11168 VSS 0.056945f
C8287 ASIG5V.n11169 VSS 0.047722f
C8288 ASIG5V.n11170 VSS 0.036092f
C8289 ASIG5V.n11171 VSS 0.036092f
C8290 ASIG5V.n11172 VSS 0.793611f
C8291 ASIG5V.n11173 VSS 0.932301f
C8292 ASIG5V.n11174 VSS 0.046728f
C8293 ASIG5V.n11175 VSS 0.046728f
C8294 ASIG5V.n11176 VSS 0.04081f
C8295 ASIG5V.n11177 VSS 0.066995f
C8296 ASIG5V.n11178 VSS 0.053548f
C8297 ASIG5V.n11179 VSS 0.061313f
C8298 ASIG5V.n11180 VSS 0.045974f
C8299 ASIG5V.n11181 VSS 0.036092f
C8300 ASIG5V.n11182 VSS 0.036092f
C8301 ASIG5V.n11183 VSS 0.839841f
C8302 ASIG5V.n11184 VSS 0.96312f
C8303 ASIG5V.n11185 VSS 0.065025f
C8304 ASIG5V.n11186 VSS 0.065025f
C8305 ASIG5V.n11187 VSS 0.058042f
C8306 ASIG5V.n11188 VSS 0.09726f
C8307 ASIG5V.n11189 VSS 0.09726f
C8308 ASIG5V.n11190 VSS 0.108961f
C8309 ASIG5V.n11191 VSS 0.108961f
C8310 ASIG5V.n11192 VSS 1.02476f
C8311 ASIG5V.n11193 VSS 0.036092f
C8312 ASIG5V.n11194 VSS 0.056945f
C8313 ASIG5V.n11195 VSS 0.056945f
C8314 ASIG5V.n11196 VSS 0.056945f
C8315 ASIG5V.n11197 VSS 0.056945f
C8316 ASIG5V.n11198 VSS 0.056945f
C8317 ASIG5V.n11199 VSS 0.056945f
C8318 ASIG5V.n11200 VSS 0.056945f
C8319 ASIG5V.n11201 VSS 0.056945f
C8320 ASIG5V.n11202 VSS 0.056945f
C8321 ASIG5V.n11203 VSS 0.056945f
C8322 ASIG5V.n11204 VSS 0.056945f
C8323 ASIG5V.n11205 VSS 0.056945f
C8324 ASIG5V.n11206 VSS 0.056945f
C8325 ASIG5V.n11207 VSS 0.056945f
C8326 ASIG5V.n11208 VSS 0.056945f
C8327 ASIG5V.n11209 VSS 0.056945f
C8328 ASIG5V.n11210 VSS 0.056945f
C8329 ASIG5V.n11211 VSS 0.056945f
C8330 ASIG5V.n11212 VSS 0.056945f
C8331 ASIG5V.n11213 VSS 0.056945f
C8332 ASIG5V.n11214 VSS 0.056945f
C8333 ASIG5V.n11215 VSS 0.056945f
C8334 ASIG5V.n11216 VSS 0.056945f
C8335 ASIG5V.n11217 VSS 0.056945f
C8336 ASIG5V.n11218 VSS 0.056945f
C8337 ASIG5V.n11219 VSS 0.056945f
C8338 ASIG5V.n11220 VSS 0.056945f
C8339 ASIG5V.n11221 VSS 0.056945f
C8340 ASIG5V.n11222 VSS 0.056945f
C8341 ASIG5V.n11223 VSS 0.056945f
C8342 ASIG5V.n11224 VSS 0.056945f
C8343 ASIG5V.n11225 VSS 0.056945f
C8344 ASIG5V.n11226 VSS 0.056945f
C8345 ASIG5V.n11227 VSS 0.056945f
C8346 ASIG5V.n11228 VSS 0.056945f
C8347 ASIG5V.n11229 VSS 0.056945f
C8348 ASIG5V.n11230 VSS 0.056945f
C8349 ASIG5V.n11231 VSS 0.056945f
C8350 ASIG5V.n11232 VSS 0.056945f
C8351 ASIG5V.n11233 VSS 0.056945f
C8352 ASIG5V.n11235 VSS 0.056945f
C8353 ASIG5V.n11236 VSS 0.056945f
C8354 ASIG5V.n11237 VSS 0.036092f
C8355 ASIG5V.n11238 VSS 0.052133f
C8356 ASIG5V.n11239 VSS 0.056945f
C8357 ASIG5V.n11240 VSS 0.056945f
C8358 ASIG5V.n11241 VSS 0.056945f
C8359 ASIG5V.n11242 VSS 0.056945f
C8360 ASIG5V.n11244 VSS 0.056945f
C8361 ASIG5V.n11245 VSS 0.056945f
C8362 ASIG5V.n11246 VSS 0.056945f
C8363 ASIG5V.n11248 VSS 0.056945f
C8364 ASIG5V.n11249 VSS 0.056945f
C8365 ASIG5V.n11250 VSS 0.056945f
C8366 ASIG5V.n11251 VSS 0.056945f
C8367 ASIG5V.n11252 VSS 0.056945f
C8368 ASIG5V.n11253 VSS 0.056945f
C8369 ASIG5V.n11254 VSS 0.056945f
C8370 ASIG5V.n11256 VSS 0.056945f
C8371 ASIG5V.n11257 VSS 0.056945f
C8372 ASIG5V.n11258 VSS 0.056945f
C8373 ASIG5V.n11260 VSS 0.056945f
C8374 ASIG5V.n11261 VSS 0.056945f
C8375 ASIG5V.n11262 VSS 0.056945f
C8376 ASIG5V.n11263 VSS 0.056945f
C8377 ASIG5V.n11264 VSS 0.056945f
C8378 ASIG5V.n11265 VSS 0.056945f
C8379 ASIG5V.n11266 VSS 0.056945f
C8380 ASIG5V.n11268 VSS 0.056945f
C8381 ASIG5V.n11269 VSS 0.056945f
C8382 ASIG5V.n11270 VSS 0.056945f
C8383 ASIG5V.n11272 VSS 0.056945f
C8384 ASIG5V.n11273 VSS 0.056945f
C8385 ASIG5V.n11274 VSS 0.056945f
C8386 ASIG5V.n11275 VSS 0.056945f
C8387 ASIG5V.n11276 VSS 0.056945f
C8388 ASIG5V.n11277 VSS 0.056945f
C8389 ASIG5V.n11278 VSS 0.056945f
C8390 ASIG5V.n11280 VSS 0.056945f
C8391 ASIG5V.n11281 VSS 0.056945f
C8392 ASIG5V.n11282 VSS 0.056945f
C8393 ASIG5V.n11284 VSS 0.056945f
C8394 ASIG5V.n11285 VSS 0.056945f
C8395 ASIG5V.n11286 VSS 0.056945f
C8396 ASIG5V.n11287 VSS 0.056945f
C8397 ASIG5V.n11288 VSS 0.056945f
C8398 ASIG5V.n11289 VSS 0.056945f
C8399 ASIG5V.n11290 VSS 0.056945f
C8400 ASIG5V.n11292 VSS 0.056945f
C8401 ASIG5V.n11293 VSS 0.056945f
C8402 ASIG5V.n11294 VSS 0.056945f
C8403 ASIG5V.n11296 VSS 0.056945f
C8404 ASIG5V.n11297 VSS 0.056945f
C8405 ASIG5V.n11298 VSS 0.056945f
C8406 ASIG5V.n11299 VSS 0.056945f
C8407 ASIG5V.n11300 VSS 0.056945f
C8408 ASIG5V.n11301 VSS 0.056945f
C8409 ASIG5V.n11302 VSS 0.056945f
C8410 ASIG5V.n11304 VSS 0.056945f
C8411 ASIG5V.n11305 VSS 0.056945f
C8412 ASIG5V.n11306 VSS 0.056945f
C8413 ASIG5V.n11308 VSS 0.056945f
C8414 ASIG5V.n11309 VSS 0.056945f
C8415 ASIG5V.n11310 VSS 0.056945f
C8416 ASIG5V.n11311 VSS 0.056945f
C8417 ASIG5V.n11312 VSS 0.056945f
C8418 ASIG5V.n11313 VSS 0.056945f
C8419 ASIG5V.n11314 VSS 0.056945f
C8420 ASIG5V.n11316 VSS 0.056945f
C8421 ASIG5V.n11317 VSS 0.056945f
C8422 ASIG5V.n11318 VSS 0.056945f
C8423 ASIG5V.n11320 VSS 0.056945f
C8424 ASIG5V.n11321 VSS 0.056945f
C8425 ASIG5V.n11322 VSS 0.056945f
C8426 ASIG5V.n11323 VSS 0.056945f
C8427 ASIG5V.n11324 VSS 0.056945f
C8428 ASIG5V.n11325 VSS 0.056945f
C8429 ASIG5V.n11326 VSS 0.056945f
C8430 ASIG5V.n11328 VSS 0.056945f
C8431 ASIG5V.n11329 VSS 0.056945f
C8432 ASIG5V.n11330 VSS 0.056945f
C8433 ASIG5V.n11332 VSS 0.056945f
C8434 ASIG5V.n11333 VSS 0.056945f
C8435 ASIG5V.n11334 VSS 0.056945f
C8436 ASIG5V.n11335 VSS 0.056945f
C8437 ASIG5V.n11336 VSS 0.056945f
C8438 ASIG5V.n11337 VSS 0.056945f
C8439 ASIG5V.n11338 VSS 0.056945f
C8440 ASIG5V.n11340 VSS 0.056945f
C8441 ASIG5V.n11341 VSS 0.056945f
C8442 ASIG5V.n11342 VSS 0.056945f
C8443 ASIG5V.n11344 VSS 0.056945f
C8444 ASIG5V.n11345 VSS 0.056945f
C8445 ASIG5V.n11346 VSS 0.056945f
C8446 ASIG5V.n11347 VSS 0.056945f
C8447 ASIG5V.n11348 VSS 0.056945f
C8448 ASIG5V.n11349 VSS 0.056945f
C8449 ASIG5V.n11350 VSS 0.056945f
C8450 ASIG5V.n11352 VSS 0.056945f
C8451 ASIG5V.n11353 VSS 0.056945f
C8452 ASIG5V.n11354 VSS 0.056945f
C8453 ASIG5V.n11356 VSS 0.056945f
C8454 ASIG5V.n11357 VSS 0.056945f
C8455 ASIG5V.n11358 VSS 0.056945f
C8456 ASIG5V.n11359 VSS 0.056945f
C8457 ASIG5V.n11360 VSS 0.056945f
C8458 ASIG5V.n11361 VSS 0.056945f
C8459 ASIG5V.n11362 VSS 0.056945f
C8460 ASIG5V.n11364 VSS 0.056945f
C8461 ASIG5V.n11365 VSS 0.056945f
C8462 ASIG5V.n11366 VSS 0.056945f
C8463 ASIG5V.n11368 VSS 0.056945f
C8464 ASIG5V.n11369 VSS 0.056945f
C8465 ASIG5V.n11370 VSS 0.056945f
C8466 ASIG5V.n11371 VSS 0.056945f
C8467 ASIG5V.n11372 VSS 0.056945f
C8468 ASIG5V.n11373 VSS 0.056945f
C8469 ASIG5V.n11374 VSS 0.056945f
C8470 ASIG5V.n11376 VSS 0.056945f
C8471 ASIG5V.n11377 VSS 0.056945f
C8472 ASIG5V.n11378 VSS 0.056945f
C8473 ASIG5V.n11380 VSS 0.056945f
C8474 ASIG5V.n11381 VSS 0.056945f
C8475 ASIG5V.n11382 VSS 0.056945f
C8476 ASIG5V.n11383 VSS 0.056945f
C8477 ASIG5V.n11384 VSS 0.056945f
C8478 ASIG5V.n11385 VSS 0.056945f
C8479 ASIG5V.n11386 VSS 0.056945f
C8480 ASIG5V.n11388 VSS 0.056945f
C8481 ASIG5V.n11389 VSS 0.056945f
C8482 ASIG5V.n11390 VSS 0.056945f
C8483 ASIG5V.n11392 VSS 0.056945f
C8484 ASIG5V.n11393 VSS 0.056945f
C8485 ASIG5V.n11394 VSS 0.056945f
C8486 ASIG5V.n11395 VSS 0.056945f
C8487 ASIG5V.n11396 VSS 0.056945f
C8488 ASIG5V.n11397 VSS 0.056945f
C8489 ASIG5V.n11398 VSS 0.056945f
C8490 ASIG5V.n11400 VSS 0.056945f
C8491 ASIG5V.n11401 VSS 0.056945f
C8492 ASIG5V.n11402 VSS 0.056945f
C8493 ASIG5V.n11404 VSS 0.056945f
C8494 ASIG5V.n11405 VSS 0.056945f
C8495 ASIG5V.n11406 VSS 0.056945f
C8496 ASIG5V.n11407 VSS 0.056945f
C8497 ASIG5V.n11408 VSS 0.056945f
C8498 ASIG5V.n11409 VSS 0.056945f
C8499 ASIG5V.n11410 VSS 0.056945f
C8500 ASIG5V.n11412 VSS 0.056945f
C8501 ASIG5V.n11413 VSS 0.056945f
C8502 ASIG5V.n11414 VSS 0.056945f
C8503 ASIG5V.n11416 VSS 0.056945f
C8504 ASIG5V.n11417 VSS 0.056945f
C8505 ASIG5V.n11418 VSS 0.056945f
C8506 ASIG5V.n11419 VSS 0.056945f
C8507 ASIG5V.n11420 VSS 0.056945f
C8508 ASIG5V.n11421 VSS 0.056945f
C8509 ASIG5V.n11422 VSS 0.056945f
C8510 ASIG5V.n11424 VSS 0.056945f
C8511 ASIG5V.n11425 VSS 0.056945f
C8512 ASIG5V.n11426 VSS 0.056945f
C8513 ASIG5V.n11428 VSS 0.056945f
C8514 ASIG5V.n11429 VSS 0.056945f
C8515 ASIG5V.n11430 VSS 0.056945f
C8516 ASIG5V.n11431 VSS 0.056945f
C8517 ASIG5V.n11432 VSS 0.056945f
C8518 ASIG5V.n11433 VSS 0.056945f
C8519 ASIG5V.n11434 VSS 0.056945f
C8520 ASIG5V.n11436 VSS 0.056945f
C8521 ASIG5V.n11437 VSS 0.056945f
C8522 ASIG5V.n11438 VSS 0.056945f
C8523 ASIG5V.n11440 VSS 0.056945f
C8524 ASIG5V.n11441 VSS 0.056945f
C8525 ASIG5V.n11442 VSS 0.056945f
C8526 ASIG5V.n11443 VSS 0.056945f
C8527 ASIG5V.n11444 VSS 0.056945f
C8528 ASIG5V.n11445 VSS 0.056945f
C8529 ASIG5V.n11446 VSS 0.056945f
C8530 ASIG5V.n11448 VSS 0.056945f
C8531 ASIG5V.n11449 VSS 0.056945f
C8532 ASIG5V.n11450 VSS 0.056945f
C8533 ASIG5V.n11452 VSS 0.056945f
C8534 ASIG5V.n11453 VSS 0.056945f
C8535 ASIG5V.n11454 VSS 0.056945f
C8536 ASIG5V.n11455 VSS 0.056945f
C8537 ASIG5V.n11456 VSS 0.056945f
C8538 ASIG5V.n11457 VSS 0.056945f
C8539 ASIG5V.n11458 VSS 0.056945f
C8540 ASIG5V.n11460 VSS 0.056945f
C8541 ASIG5V.n11461 VSS 0.056945f
C8542 ASIG5V.n11462 VSS 0.056945f
C8543 ASIG5V.n11464 VSS 0.056945f
C8544 ASIG5V.n11465 VSS 0.056945f
C8545 ASIG5V.n11466 VSS 0.056945f
C8546 ASIG5V.n11467 VSS 0.056945f
C8547 ASIG5V.n11468 VSS 0.056945f
C8548 ASIG5V.n11469 VSS 0.056945f
C8549 ASIG5V.n11470 VSS 0.056945f
C8550 ASIG5V.n11472 VSS 0.056945f
C8551 ASIG5V.n11473 VSS 0.056945f
C8552 ASIG5V.n11474 VSS 0.056945f
C8553 ASIG5V.n11476 VSS 0.056945f
C8554 ASIG5V.n11477 VSS 0.056945f
C8555 ASIG5V.n11478 VSS 0.056945f
C8556 ASIG5V.n11479 VSS 0.056945f
C8557 ASIG5V.n11480 VSS 0.056945f
C8558 ASIG5V.n11481 VSS 0.056945f
C8559 ASIG5V.n11482 VSS 0.056945f
C8560 ASIG5V.n11484 VSS 0.036092f
C8561 ASIG5V.n11485 VSS 0.531642f
C8562 ASIG5V.n11486 VSS 0.493117f
C8563 ASIG5V.n11487 VSS 0.05429f
C8564 ASIG5V.n11488 VSS 0.05429f
C8565 ASIG5V.n11489 VSS 0.047415f
C8566 ASIG5V.n11490 VSS 0.052746f
C8567 ASIG5V.n11491 VSS 0.053077f
C8568 ASIG5V.n11492 VSS 0.060773f
C8569 ASIG5V.n11493 VSS 0.060773f
C8570 ASIG5V.n11494 VSS 0.354427f
C8571 ASIG5V.n11495 VSS 1.0941f
C8572 ASIG5V.n11496 VSS 0.107203f
C8573 ASIG5V.n11497 VSS 0.107203f
C8574 ASIG5V.n11498 VSS 0.095691f
C8575 ASIG5V.n11499 VSS 0.09726f
C8576 ASIG5V.n11500 VSS 0.06118f
C8577 ASIG5V.n11501 VSS 0.06854f
C8578 ASIG5V.n11502 VSS 0.0621f
C8579 ASIG5V.n11503 VSS 0.036092f
C8580 ASIG5V.n11504 VSS 0.052133f
C8581 ASIG5V.n11505 VSS 0.056945f
C8582 ASIG5V.n11506 VSS 0.056945f
C8583 ASIG5V.n11507 VSS 0.056945f
C8584 ASIG5V.n11508 VSS 0.056945f
C8585 ASIG5V.n11510 VSS 0.056945f
C8586 ASIG5V.n11511 VSS 0.056945f
C8587 ASIG5V.n11512 VSS 0.056945f
C8588 ASIG5V.n11514 VSS 0.056945f
C8589 ASIG5V.n11515 VSS 0.056945f
C8590 ASIG5V.n11516 VSS 0.056945f
C8591 ASIG5V.n11517 VSS 0.056945f
C8592 ASIG5V.n11518 VSS 0.056945f
C8593 ASIG5V.n11519 VSS 0.056945f
C8594 ASIG5V.n11520 VSS 0.056945f
C8595 ASIG5V.n11522 VSS 0.056945f
C8596 ASIG5V.n11523 VSS 0.056945f
C8597 ASIG5V.n11524 VSS 0.056945f
C8598 ASIG5V.n11526 VSS 0.056945f
C8599 ASIG5V.n11527 VSS 0.056945f
C8600 ASIG5V.n11528 VSS 0.056945f
C8601 ASIG5V.n11529 VSS 0.056945f
C8602 ASIG5V.n11530 VSS 0.056945f
C8603 ASIG5V.n11531 VSS 0.056945f
C8604 ASIG5V.n11532 VSS 0.056945f
C8605 ASIG5V.n11534 VSS 0.056945f
C8606 ASIG5V.n11535 VSS 0.056945f
C8607 ASIG5V.n11536 VSS 0.056945f
C8608 ASIG5V.n11538 VSS 0.056945f
C8609 ASIG5V.n11539 VSS 0.056945f
C8610 ASIG5V.n11540 VSS 0.056945f
C8611 ASIG5V.n11541 VSS 0.056945f
C8612 ASIG5V.n11542 VSS 0.056945f
C8613 ASIG5V.n11543 VSS 0.056945f
C8614 ASIG5V.n11544 VSS 0.056945f
C8615 ASIG5V.n11546 VSS 0.056945f
C8616 ASIG5V.n11547 VSS 0.056945f
C8617 ASIG5V.n11548 VSS 0.056945f
C8618 ASIG5V.n11550 VSS 0.056945f
C8619 ASIG5V.n11551 VSS 0.056945f
C8620 ASIG5V.n11552 VSS 0.056945f
C8621 ASIG5V.n11553 VSS 0.056945f
C8622 ASIG5V.n11554 VSS 0.056945f
C8623 ASIG5V.n11555 VSS 0.056945f
C8624 ASIG5V.n11556 VSS 0.056945f
C8625 ASIG5V.n11558 VSS 0.056945f
C8626 ASIG5V.n11559 VSS 0.056945f
C8627 ASIG5V.n11560 VSS 0.056945f
C8628 ASIG5V.n11562 VSS 0.056945f
C8629 ASIG5V.n11563 VSS 0.056945f
C8630 ASIG5V.n11564 VSS 0.056945f
C8631 ASIG5V.n11565 VSS 0.056945f
C8632 ASIG5V.n11566 VSS 0.056945f
C8633 ASIG5V.n11567 VSS 0.056945f
C8634 ASIG5V.n11568 VSS 0.056945f
C8635 ASIG5V.n11570 VSS 0.056945f
C8636 ASIG5V.n11571 VSS 0.056945f
C8637 ASIG5V.n11572 VSS 0.056945f
C8638 ASIG5V.n11574 VSS 0.056945f
C8639 ASIG5V.n11575 VSS 0.056945f
C8640 ASIG5V.n11576 VSS 0.056945f
C8641 ASIG5V.n11577 VSS 0.056945f
C8642 ASIG5V.n11578 VSS 0.056945f
C8643 ASIG5V.n11579 VSS 0.056945f
C8644 ASIG5V.n11580 VSS 0.056945f
C8645 ASIG5V.n11582 VSS 0.056945f
C8646 ASIG5V.n11583 VSS 0.056945f
C8647 ASIG5V.n11584 VSS 0.056945f
C8648 ASIG5V.n11586 VSS 0.056945f
C8649 ASIG5V.n11587 VSS 0.056945f
C8650 ASIG5V.n11588 VSS 0.056945f
C8651 ASIG5V.n11589 VSS 0.056945f
C8652 ASIG5V.n11590 VSS 0.056945f
C8653 ASIG5V.n11591 VSS 0.056945f
C8654 ASIG5V.n11592 VSS 0.056945f
C8655 ASIG5V.n11594 VSS 0.056945f
C8656 ASIG5V.n11595 VSS 0.056945f
C8657 ASIG5V.n11596 VSS 0.056945f
C8658 ASIG5V.n11598 VSS 0.056945f
C8659 ASIG5V.n11599 VSS 0.056945f
C8660 ASIG5V.n11600 VSS 0.056945f
C8661 ASIG5V.n11601 VSS 0.056945f
C8662 ASIG5V.n11602 VSS 0.056945f
C8663 ASIG5V.n11603 VSS 0.056945f
C8664 ASIG5V.n11604 VSS 0.056945f
C8665 ASIG5V.n11606 VSS 0.056945f
C8666 ASIG5V.n11607 VSS 0.056945f
C8667 ASIG5V.n11608 VSS 0.056945f
C8668 ASIG5V.n11610 VSS 0.056945f
C8669 ASIG5V.n11611 VSS 0.056945f
C8670 ASIG5V.n11612 VSS 0.056945f
C8671 ASIG5V.n11613 VSS 0.056945f
C8672 ASIG5V.n11614 VSS 0.056945f
C8673 ASIG5V.n11615 VSS 0.056945f
C8674 ASIG5V.n11616 VSS 0.056945f
C8675 ASIG5V.n11618 VSS 0.056945f
C8676 ASIG5V.n11619 VSS 0.056945f
C8677 ASIG5V.n11620 VSS 0.056945f
C8678 ASIG5V.n11622 VSS 0.056945f
C8679 ASIG5V.n11623 VSS 0.056945f
C8680 ASIG5V.n11624 VSS 0.056945f
C8681 ASIG5V.n11625 VSS 0.056945f
C8682 ASIG5V.n11626 VSS 0.056945f
C8683 ASIG5V.n11627 VSS 0.056945f
C8684 ASIG5V.n11628 VSS 0.056945f
C8685 ASIG5V.n11630 VSS 0.056945f
C8686 ASIG5V.n11631 VSS 0.056945f
C8687 ASIG5V.n11632 VSS 0.056945f
C8688 ASIG5V.n11634 VSS 0.056945f
C8689 ASIG5V.n11635 VSS 0.056945f
C8690 ASIG5V.n11636 VSS 0.056945f
C8691 ASIG5V.n11637 VSS 0.056945f
C8692 ASIG5V.n11638 VSS 0.056945f
C8693 ASIG5V.n11639 VSS 0.056945f
C8694 ASIG5V.n11640 VSS 0.056945f
C8695 ASIG5V.n11642 VSS 0.056945f
C8696 ASIG5V.n11643 VSS 0.056945f
C8697 ASIG5V.n11644 VSS 0.056945f
C8698 ASIG5V.n11646 VSS 0.056945f
C8699 ASIG5V.n11647 VSS 0.056945f
C8700 ASIG5V.n11648 VSS 0.056945f
C8701 ASIG5V.n11649 VSS 0.056945f
C8702 ASIG5V.n11650 VSS 0.056945f
C8703 ASIG5V.n11651 VSS 0.056945f
C8704 ASIG5V.n11652 VSS 0.056945f
C8705 ASIG5V.n11654 VSS 0.056945f
C8706 ASIG5V.n11655 VSS 0.056945f
C8707 ASIG5V.n11656 VSS 0.056945f
C8708 ASIG5V.n11658 VSS 0.056945f
C8709 ASIG5V.n11659 VSS 0.056945f
C8710 ASIG5V.n11660 VSS 0.056945f
C8711 ASIG5V.n11661 VSS 0.056945f
C8712 ASIG5V.n11662 VSS 0.056945f
C8713 ASIG5V.n11663 VSS 0.056945f
C8714 ASIG5V.n11664 VSS 0.056945f
C8715 ASIG5V.n11666 VSS 0.056945f
C8716 ASIG5V.n11667 VSS 0.056945f
C8717 ASIG5V.n11668 VSS 0.056945f
C8718 ASIG5V.n11670 VSS 0.056945f
C8719 ASIG5V.n11671 VSS 0.056945f
C8720 ASIG5V.n11672 VSS 0.056945f
C8721 ASIG5V.n11673 VSS 0.056945f
C8722 ASIG5V.n11674 VSS 0.056945f
C8723 ASIG5V.n11675 VSS 0.056945f
C8724 ASIG5V.n11676 VSS 0.056945f
C8725 ASIG5V.n11678 VSS 0.056945f
C8726 ASIG5V.n11679 VSS 0.056945f
C8727 ASIG5V.n11680 VSS 0.056945f
C8728 ASIG5V.n11682 VSS 0.056945f
C8729 ASIG5V.n11683 VSS 0.056945f
C8730 ASIG5V.n11684 VSS 0.056945f
C8731 ASIG5V.n11685 VSS 0.056945f
C8732 ASIG5V.n11686 VSS 0.056945f
C8733 ASIG5V.n11687 VSS 0.056945f
C8734 ASIG5V.n11688 VSS 0.056945f
C8735 ASIG5V.n11690 VSS 0.056945f
C8736 ASIG5V.n11691 VSS 0.056945f
C8737 ASIG5V.n11692 VSS 0.056945f
C8738 ASIG5V.n11694 VSS 0.056945f
C8739 ASIG5V.n11695 VSS 0.056945f
C8740 ASIG5V.n11696 VSS 0.056945f
C8741 ASIG5V.n11697 VSS 0.056945f
C8742 ASIG5V.n11698 VSS 0.056945f
C8743 ASIG5V.n11699 VSS 0.056945f
C8744 ASIG5V.n11700 VSS 0.056945f
C8745 ASIG5V.n11702 VSS 0.056945f
C8746 ASIG5V.n11703 VSS 0.056945f
C8747 ASIG5V.n11704 VSS 0.056945f
C8748 ASIG5V.n11706 VSS 0.056945f
C8749 ASIG5V.n11707 VSS 0.056945f
C8750 ASIG5V.n11708 VSS 0.056945f
C8751 ASIG5V.n11709 VSS 0.056945f
C8752 ASIG5V.n11710 VSS 0.056945f
C8753 ASIG5V.n11711 VSS 0.056945f
C8754 ASIG5V.n11712 VSS 0.056945f
C8755 ASIG5V.n11714 VSS 0.056945f
C8756 ASIG5V.n11715 VSS 0.056945f
C8757 ASIG5V.n11716 VSS 0.056945f
C8758 ASIG5V.n11718 VSS 0.056945f
C8759 ASIG5V.n11719 VSS 0.056945f
C8760 ASIG5V.n11720 VSS 0.056945f
C8761 ASIG5V.n11721 VSS 0.056945f
C8762 ASIG5V.n11722 VSS 0.056945f
C8763 ASIG5V.n11723 VSS 0.056945f
C8764 ASIG5V.n11724 VSS 0.056945f
C8765 ASIG5V.n11726 VSS 0.056945f
C8766 ASIG5V.n11727 VSS 0.056945f
C8767 ASIG5V.n11728 VSS 0.056945f
C8768 ASIG5V.n11730 VSS 0.056945f
C8769 ASIG5V.n11731 VSS 0.056945f
C8770 ASIG5V.n11732 VSS 0.056945f
C8771 ASIG5V.n11733 VSS 0.056945f
C8772 ASIG5V.n11734 VSS 0.056945f
C8773 ASIG5V.n11735 VSS 0.056945f
C8774 ASIG5V.n11736 VSS 0.056945f
C8775 ASIG5V.n11738 VSS 0.056945f
C8776 ASIG5V.n11739 VSS 0.056945f
C8777 ASIG5V.n11740 VSS 0.056945f
C8778 ASIG5V.n11742 VSS 0.056945f
C8779 ASIG5V.n11743 VSS 0.056945f
C8780 ASIG5V.n11744 VSS 0.056945f
C8781 ASIG5V.n11745 VSS 0.056945f
C8782 ASIG5V.n11746 VSS 0.056945f
C8783 ASIG5V.n11747 VSS 0.056945f
C8784 ASIG5V.n11748 VSS 0.056945f
C8785 ASIG5V.n11750 VSS 0.036092f
C8786 ASIG5V.n11751 VSS 0.947711f
C8787 ASIG5V.n11752 VSS 0.300493f
C8788 ASIG5V.n11753 VSS 0.047268f
C8789 ASIG5V.n11754 VSS 0.047268f
C8790 ASIG5V.n11755 VSS 0.041282f
C8791 ASIG5V.n11756 VSS 0.052746f
C8792 ASIG5V.n11757 VSS 0.05921f
C8793 ASIG5V.n11758 VSS 0.067796f
C8794 ASIG5V.n11759 VSS 0.067796f
C8795 ASIG5V.n11760 VSS 0.076709f
C8796 ASIG5V.n11761 VSS 0.040245f
C8797 ASIG5V.n11762 VSS 0.040245f
C8798 ASIG5V.n11763 VSS 0.035149f
C8799 ASIG5V.n11764 VSS 0.052746f
C8800 ASIG5V.n11765 VSS 0.047722f
C8801 ASIG5V.n11766 VSS 0.056945f
C8802 ASIG5V.n11767 VSS 0.056945f
C8803 ASIG5V.n11768 VSS 0.056945f
C8804 ASIG5V.n11770 VSS 0.036092f
C8805 ASIG5V.n11771 VSS 0.685742f
C8806 ASIG5V.n11772 VSS 0.516232f
C8807 ASIG5V.n11773 VSS 0.080842f
C8808 ASIG5V.n11774 VSS 0.080842f
C8809 ASIG5V.n11775 VSS 0.072161f
C8810 ASIG5V.n11776 VSS 0.07229f
C8811 ASIG5V.n11777 VSS 0.073729f
C8812 ASIG5V.n11778 VSS 0.09726f
C8813 ASIG5V.n11779 VSS 0.108961f
C8814 ASIG5V.n11780 VSS 0.108961f
C8815 ASIG5V.n11781 VSS 1.0941f
C8816 ASIG5V.n11782 VSS 0.955415f
C8817 ASIG5V.n11783 VSS 0.071577f
C8818 ASIG5V.n11784 VSS 0.071577f
C8819 ASIG5V.n11785 VSS 0.062513f
C8820 ASIG5V.n11786 VSS 0.052746f
C8821 ASIG5V.n11787 VSS 0.037979f
C8822 ASIG5V.n11788 VSS 0.066995f
C8823 ASIG5V.n11789 VSS 0.076709f
C8824 ASIG5V.n11790 VSS 0.076709f
C8825 ASIG5V.n11791 VSS 0.955415f
C8826 ASIG5V.n11792 VSS 1.0941f
C8827 ASIG5V.n11793 VSS 0.105446f
C8828 ASIG5V.n11794 VSS 0.105446f
C8829 ASIG5V.n11795 VSS 0.094123f
C8830 ASIG5V.n11796 VSS 0.07229f
C8831 ASIG5V.n11797 VSS 0.047061f
C8832 ASIG5V.n11798 VSS 0.548344f
C8833 ASIG5V.n11799 VSS 0.053336f
C8834 ASIG5V.n11800 VSS 0.108961f
C8835 ASIG5V.n11801 VSS 0.108961f
C8836 ASIG5V.n11802 VSS 0.108961f
C8837 ASIG5V.n11803 VSS 0.063267f
C8838 ASIG5V.n11804 VSS 0.063267f
C8839 ASIG5V.n11805 VSS 0.056474f
C8840 ASIG5V.n11806 VSS 0.07229f
C8841 ASIG5V.n11807 VSS 0.052133f
C8842 ASIG5V.n11808 VSS 0.056945f
C8843 ASIG5V.n11809 VSS 0.056945f
C8844 ASIG5V.n11810 VSS 0.056945f
C8845 ASIG5V.n11811 VSS 0.056945f
C8846 ASIG5V.n11812 VSS 0.056945f
C8847 ASIG5V.n11813 VSS 0.056945f
C8848 ASIG5V.n11814 VSS 0.056945f
C8849 ASIG5V.n11815 VSS 0.056945f
C8850 ASIG5V.n11816 VSS 0.056945f
C8851 ASIG5V.n11817 VSS 0.056945f
C8852 ASIG5V.n11818 VSS 0.056945f
C8853 ASIG5V.n11819 VSS 0.056945f
C8854 ASIG5V.n11820 VSS 0.056945f
C8855 ASIG5V.n11821 VSS 0.056945f
C8856 ASIG5V.n11822 VSS 0.056945f
C8857 ASIG5V.n11823 VSS 0.056945f
C8858 ASIG5V.n11824 VSS 0.056945f
C8859 ASIG5V.n11825 VSS 0.056945f
C8860 ASIG5V.n11826 VSS 0.056945f
C8861 ASIG5V.n11827 VSS 0.056945f
C8862 ASIG5V.n11828 VSS 0.056945f
C8863 ASIG5V.n11829 VSS 0.056945f
C8864 ASIG5V.n11830 VSS 0.056945f
C8865 ASIG5V.n11831 VSS 0.056945f
C8866 ASIG5V.n11832 VSS 0.056945f
C8867 ASIG5V.n11833 VSS 0.056945f
C8868 ASIG5V.n11834 VSS 0.056945f
C8869 ASIG5V.n11835 VSS 0.056945f
C8870 ASIG5V.n11836 VSS 0.056945f
C8871 ASIG5V.n11837 VSS 0.056945f
C8872 ASIG5V.n11838 VSS 0.056945f
C8873 ASIG5V.n11839 VSS 0.056945f
C8874 ASIG5V.n11840 VSS 0.056945f
C8875 ASIG5V.n11841 VSS 0.056945f
C8876 ASIG5V.n11842 VSS 0.056945f
C8877 ASIG5V.n11843 VSS 0.056945f
C8878 ASIG5V.n11844 VSS 0.056945f
C8879 ASIG5V.n11845 VSS 0.056945f
C8880 ASIG5V.n11846 VSS 0.056945f
C8881 ASIG5V.n11847 VSS 0.056945f
C8882 ASIG5V.n11848 VSS 0.056945f
C8883 ASIG5V.n11849 VSS 0.056945f
C8884 ASIG5V.n11850 VSS 0.056945f
C8885 ASIG5V.n11851 VSS 0.056945f
C8886 ASIG5V.n11852 VSS 0.056945f
C8887 ASIG5V.n11853 VSS 0.056945f
C8888 ASIG5V.n11854 VSS 0.056945f
C8889 ASIG5V.n11855 VSS 0.056945f
C8890 ASIG5V.n11856 VSS 0.056945f
C8891 ASIG5V.n11857 VSS 0.056945f
C8892 ASIG5V.n11858 VSS 0.056945f
C8893 ASIG5V.n11859 VSS 0.056945f
C8894 ASIG5V.n11860 VSS 0.056945f
C8895 ASIG5V.n11861 VSS 0.056945f
C8896 ASIG5V.n11862 VSS 0.056945f
C8897 ASIG5V.n11863 VSS 0.056945f
C8898 ASIG5V.n11864 VSS 0.056945f
C8899 ASIG5V.n11865 VSS 0.056945f
C8900 ASIG5V.n11866 VSS 0.056945f
C8901 ASIG5V.n11867 VSS 0.056945f
C8902 ASIG5V.n11868 VSS 0.056945f
C8903 ASIG5V.n11869 VSS 0.056945f
C8904 ASIG5V.n11870 VSS 0.056945f
C8905 ASIG5V.n11871 VSS 0.056945f
C8906 ASIG5V.n11872 VSS 0.056945f
C8907 ASIG5V.n11873 VSS 0.056945f
C8908 ASIG5V.n11874 VSS 0.056945f
C8909 ASIG5V.n11875 VSS 0.056945f
C8910 ASIG5V.n11876 VSS 0.056945f
C8911 ASIG5V.n11877 VSS 0.056945f
C8912 ASIG5V.n11878 VSS 0.056945f
C8913 ASIG5V.n11879 VSS 0.056945f
C8914 ASIG5V.n11880 VSS 0.056945f
C8915 ASIG5V.n11881 VSS 0.056945f
C8916 ASIG5V.n11882 VSS 0.056945f
C8917 ASIG5V.n11883 VSS 0.056945f
C8918 ASIG5V.n11884 VSS 0.056945f
C8919 ASIG5V.n11885 VSS 0.056945f
C8920 ASIG5V.n11886 VSS 0.056945f
C8921 ASIG5V.n11887 VSS 0.056945f
C8922 ASIG5V.n11888 VSS 0.056945f
C8923 ASIG5V.n11889 VSS 0.056945f
C8924 ASIG5V.n11890 VSS 0.056945f
C8925 ASIG5V.n11891 VSS 0.056945f
C8926 ASIG5V.n11892 VSS 0.056945f
C8927 ASIG5V.n11893 VSS 0.056945f
C8928 ASIG5V.n11894 VSS 0.056945f
C8929 ASIG5V.n11895 VSS 0.056945f
C8930 ASIG5V.n11896 VSS 0.056945f
C8931 ASIG5V.n11897 VSS 0.056945f
C8932 ASIG5V.n11898 VSS 0.056945f
C8933 ASIG5V.n11899 VSS 0.056945f
C8934 ASIG5V.n11900 VSS 0.056945f
C8935 ASIG5V.n11901 VSS 0.056945f
C8936 ASIG5V.n11902 VSS 0.056945f
C8937 ASIG5V.n11903 VSS 0.056945f
C8938 ASIG5V.n11904 VSS 0.056945f
C8939 ASIG5V.n11905 VSS 0.056945f
C8940 ASIG5V.n11906 VSS 0.056945f
C8941 ASIG5V.n11907 VSS 0.056945f
C8942 ASIG5V.n11908 VSS 0.056945f
C8943 ASIG5V.n11909 VSS 0.056945f
C8944 ASIG5V.n11910 VSS 0.056945f
C8945 ASIG5V.n11911 VSS 0.056945f
C8946 ASIG5V.n11912 VSS 0.056945f
C8947 ASIG5V.n11913 VSS 0.056945f
C8948 ASIG5V.n11914 VSS 0.056945f
C8949 ASIG5V.n11915 VSS 0.056945f
C8950 ASIG5V.n11916 VSS 0.056945f
C8951 ASIG5V.n11917 VSS 0.056945f
C8952 ASIG5V.n11918 VSS 0.056945f
C8953 ASIG5V.n11919 VSS 0.056945f
C8954 ASIG5V.n11920 VSS 0.056945f
C8955 ASIG5V.n11921 VSS 0.056945f
C8956 ASIG5V.n11922 VSS 0.056945f
C8957 ASIG5V.n11923 VSS 0.056945f
C8958 ASIG5V.n11924 VSS 0.056945f
C8959 ASIG5V.n11925 VSS 0.056945f
C8960 ASIG5V.n11926 VSS 0.056945f
C8961 ASIG5V.n11927 VSS 0.056945f
C8962 ASIG5V.n11928 VSS 0.056945f
C8963 ASIG5V.n11929 VSS 0.056945f
C8964 ASIG5V.n11930 VSS 0.056945f
C8965 ASIG5V.n11931 VSS 0.056945f
C8966 ASIG5V.n11932 VSS 0.056945f
C8967 ASIG5V.n11933 VSS 0.056945f
C8968 ASIG5V.n11934 VSS 0.056945f
C8969 ASIG5V.n11935 VSS 0.056945f
C8970 ASIG5V.n11936 VSS 0.056945f
C8971 ASIG5V.n11937 VSS 0.056945f
C8972 ASIG5V.n11938 VSS 0.056945f
C8973 ASIG5V.n11939 VSS 0.056945f
C8974 ASIG5V.n11940 VSS 0.056945f
C8975 ASIG5V.n11941 VSS 0.056945f
C8976 ASIG5V.n11942 VSS 0.056945f
C8977 ASIG5V.n11943 VSS 0.056945f
C8978 ASIG5V.n11944 VSS 0.056945f
C8979 ASIG5V.n11945 VSS 0.056945f
C8980 ASIG5V.n11946 VSS 0.056945f
C8981 ASIG5V.n11947 VSS 0.056945f
C8982 ASIG5V.n11948 VSS 0.056945f
C8983 ASIG5V.n11949 VSS 0.056945f
C8984 ASIG5V.n11950 VSS 0.056945f
C8985 ASIG5V.n11951 VSS 0.056945f
C8986 ASIG5V.n11952 VSS 0.056945f
C8987 ASIG5V.n11953 VSS 0.056945f
C8988 ASIG5V.n11954 VSS 0.056945f
C8989 ASIG5V.n11955 VSS 0.056945f
C8990 ASIG5V.n11956 VSS 0.056945f
C8991 ASIG5V.n11957 VSS 0.056945f
C8992 ASIG5V.n11958 VSS 0.056945f
C8993 ASIG5V.n11959 VSS 0.056945f
C8994 ASIG5V.n11960 VSS 0.056945f
C8995 ASIG5V.n11961 VSS 0.056945f
C8996 ASIG5V.n11962 VSS 0.056945f
C8997 ASIG5V.n11963 VSS 0.056945f
C8998 ASIG5V.n11964 VSS 0.056945f
C8999 ASIG5V.n11965 VSS 0.056945f
C9000 ASIG5V.n11966 VSS 0.056945f
C9001 ASIG5V.n11967 VSS 0.056945f
C9002 ASIG5V.n11968 VSS 0.056945f
C9003 ASIG5V.n11969 VSS 0.056945f
C9004 ASIG5V.n11970 VSS 0.056945f
C9005 ASIG5V.n11971 VSS 0.056945f
C9006 ASIG5V.n11972 VSS 0.056945f
C9007 ASIG5V.n11973 VSS 0.056945f
C9008 ASIG5V.n11974 VSS 0.056945f
C9009 ASIG5V.n11975 VSS 0.056945f
C9010 ASIG5V.n11976 VSS 0.056945f
C9011 ASIG5V.n11977 VSS 0.056945f
C9012 ASIG5V.n11978 VSS 0.056945f
C9013 ASIG5V.n11979 VSS 0.056945f
C9014 ASIG5V.n11980 VSS 0.056945f
C9015 ASIG5V.n11981 VSS 0.056945f
C9016 ASIG5V.n11982 VSS 0.056945f
C9017 ASIG5V.n11983 VSS 0.056945f
C9018 ASIG5V.n11984 VSS 0.056945f
C9019 ASIG5V.n11985 VSS 0.056945f
C9020 ASIG5V.n11986 VSS 0.056945f
C9021 ASIG5V.n11987 VSS 0.056945f
C9022 ASIG5V.n11988 VSS 0.056945f
C9023 ASIG5V.n11989 VSS 0.056945f
C9024 ASIG5V.n11990 VSS 0.056945f
C9025 ASIG5V.n11991 VSS 0.047722f
C9026 ASIG5V.n11992 VSS 0.036092f
C9027 ASIG5V.n11993 VSS 0.036092f
C9028 ASIG5V.n11994 VSS 0.562462f
C9029 ASIG5V.n11995 VSS 0.036092f
C9030 ASIG5V.n11997 VSS 0.701152f
C9031 ASIG5V.n11998 VSS 0.277378f
C9032 ASIG5V.n11999 VSS 0.057532f
C9033 ASIG5V.n12000 VSS 0.057532f
C9034 ASIG5V.n12001 VSS 0.050246f
C9035 ASIG5V.n12002 VSS 0.066995f
C9036 ASIG5V.n12003 VSS 0.044113f
C9037 ASIG5V.n12004 VSS 0.050509f
C9038 ASIG5V.n12005 VSS 0.045974f
C9039 ASIG5V.n12006 VSS 0.036092f
C9040 ASIG5V.n12007 VSS 0.036092f
C9041 ASIG5V.n12008 VSS 0.955415f
C9042 ASIG5V.n12009 VSS 0.036092f
C9043 ASIG5V.n12011 VSS 0.932301f
C9044 ASIG5V.n12012 VSS 0.246558f
C9045 ASIG5V.n12013 VSS 0.087871f
C9046 ASIG5V.n12014 VSS 0.087871f
C9047 ASIG5V.n12015 VSS 0.078436f
C9048 ASIG5V.n12016 VSS 0.09726f
C9049 ASIG5V.n12017 VSS 0.078436f
C9050 ASIG5V.n12018 VSS 0.087871f
C9051 ASIG5V.n12019 VSS 0.0621f
C9052 ASIG5V.n12020 VSS 0.036092f
C9053 ASIG5V.n12021 VSS 0.052133f
C9054 ASIG5V.n12022 VSS 0.056945f
C9055 ASIG5V.n12023 VSS 0.056945f
C9056 ASIG5V.n12024 VSS 0.056945f
C9057 ASIG5V.n12025 VSS 0.056945f
C9058 ASIG5V.n12027 VSS 0.056945f
C9059 ASIG5V.n12028 VSS 0.056945f
C9060 ASIG5V.n12029 VSS 0.056945f
C9061 ASIG5V.n12031 VSS 0.056945f
C9062 ASIG5V.n12032 VSS 0.056945f
C9063 ASIG5V.n12033 VSS 0.056945f
C9064 ASIG5V.n12034 VSS 0.056945f
C9065 ASIG5V.n12035 VSS 0.056945f
C9066 ASIG5V.n12036 VSS 0.056945f
C9067 ASIG5V.n12037 VSS 0.056945f
C9068 ASIG5V.n12039 VSS 0.056945f
C9069 ASIG5V.n12040 VSS 0.056945f
C9070 ASIG5V.n12041 VSS 0.056945f
C9071 ASIG5V.n12043 VSS 0.056945f
C9072 ASIG5V.n12044 VSS 0.056945f
C9073 ASIG5V.n12045 VSS 0.056945f
C9074 ASIG5V.n12046 VSS 0.056945f
C9075 ASIG5V.n12047 VSS 0.056945f
C9076 ASIG5V.n12048 VSS 0.056945f
C9077 ASIG5V.n12049 VSS 0.056945f
C9078 ASIG5V.n12051 VSS 0.056945f
C9079 ASIG5V.n12052 VSS 0.056945f
C9080 ASIG5V.n12053 VSS 0.056945f
C9081 ASIG5V.n12055 VSS 0.056945f
C9082 ASIG5V.n12056 VSS 0.056945f
C9083 ASIG5V.n12057 VSS 0.056945f
C9084 ASIG5V.n12058 VSS 0.056945f
C9085 ASIG5V.n12059 VSS 0.056945f
C9086 ASIG5V.n12060 VSS 0.056945f
C9087 ASIG5V.n12061 VSS 0.056945f
C9088 ASIG5V.n12063 VSS 0.056945f
C9089 ASIG5V.n12064 VSS 0.056945f
C9090 ASIG5V.n12065 VSS 0.056945f
C9091 ASIG5V.n12067 VSS 0.056945f
C9092 ASIG5V.n12068 VSS 0.056945f
C9093 ASIG5V.n12069 VSS 0.056945f
C9094 ASIG5V.n12070 VSS 0.056945f
C9095 ASIG5V.n12071 VSS 0.056945f
C9096 ASIG5V.n12072 VSS 0.056945f
C9097 ASIG5V.n12073 VSS 0.056945f
C9098 ASIG5V.n12075 VSS 0.056945f
C9099 ASIG5V.n12076 VSS 0.056945f
C9100 ASIG5V.n12077 VSS 0.056945f
C9101 ASIG5V.n12079 VSS 0.056945f
C9102 ASIG5V.n12080 VSS 0.056945f
C9103 ASIG5V.n12081 VSS 0.056945f
C9104 ASIG5V.n12082 VSS 0.056945f
C9105 ASIG5V.n12083 VSS 0.056945f
C9106 ASIG5V.n12084 VSS 0.056945f
C9107 ASIG5V.n12085 VSS 0.056945f
C9108 ASIG5V.n12087 VSS 0.056945f
C9109 ASIG5V.n12088 VSS 0.056945f
C9110 ASIG5V.n12089 VSS 0.056945f
C9111 ASIG5V.n12091 VSS 0.056945f
C9112 ASIG5V.n12092 VSS 0.056945f
C9113 ASIG5V.n12093 VSS 0.056945f
C9114 ASIG5V.n12094 VSS 0.056945f
C9115 ASIG5V.n12095 VSS 0.056945f
C9116 ASIG5V.n12096 VSS 0.056945f
C9117 ASIG5V.n12097 VSS 0.056945f
C9118 ASIG5V.n12099 VSS 0.056945f
C9119 ASIG5V.n12100 VSS 0.056945f
C9120 ASIG5V.n12101 VSS 0.056945f
C9121 ASIG5V.n12103 VSS 0.056945f
C9122 ASIG5V.n12104 VSS 0.056945f
C9123 ASIG5V.n12105 VSS 0.056945f
C9124 ASIG5V.n12106 VSS 0.056945f
C9125 ASIG5V.n12107 VSS 0.056945f
C9126 ASIG5V.n12108 VSS 0.056945f
C9127 ASIG5V.n12109 VSS 0.056945f
C9128 ASIG5V.n12111 VSS 0.056945f
C9129 ASIG5V.n12112 VSS 0.056945f
C9130 ASIG5V.n12113 VSS 0.056945f
C9131 ASIG5V.n12115 VSS 0.056945f
C9132 ASIG5V.n12116 VSS 0.056945f
C9133 ASIG5V.n12117 VSS 0.056945f
C9134 ASIG5V.n12118 VSS 0.056945f
C9135 ASIG5V.n12119 VSS 0.056945f
C9136 ASIG5V.n12120 VSS 0.056945f
C9137 ASIG5V.n12121 VSS 0.056945f
C9138 ASIG5V.n12123 VSS 0.056945f
C9139 ASIG5V.n12124 VSS 0.056945f
C9140 ASIG5V.n12125 VSS 0.056945f
C9141 ASIG5V.n12127 VSS 0.056945f
C9142 ASIG5V.n12128 VSS 0.056945f
C9143 ASIG5V.n12129 VSS 0.056945f
C9144 ASIG5V.n12130 VSS 0.056945f
C9145 ASIG5V.n12131 VSS 0.056945f
C9146 ASIG5V.n12132 VSS 0.056945f
C9147 ASIG5V.n12133 VSS 0.056945f
C9148 ASIG5V.n12135 VSS 0.056945f
C9149 ASIG5V.n12136 VSS 0.056945f
C9150 ASIG5V.n12137 VSS 0.056945f
C9151 ASIG5V.n12139 VSS 0.056945f
C9152 ASIG5V.n12140 VSS 0.056945f
C9153 ASIG5V.n12141 VSS 0.056945f
C9154 ASIG5V.n12142 VSS 0.056945f
C9155 ASIG5V.n12143 VSS 0.056945f
C9156 ASIG5V.n12144 VSS 0.056945f
C9157 ASIG5V.n12145 VSS 0.056945f
C9158 ASIG5V.n12147 VSS 0.056945f
C9159 ASIG5V.n12148 VSS 0.056945f
C9160 ASIG5V.n12149 VSS 0.056945f
C9161 ASIG5V.n12151 VSS 0.056945f
C9162 ASIG5V.n12152 VSS 0.056945f
C9163 ASIG5V.n12153 VSS 0.056945f
C9164 ASIG5V.n12154 VSS 0.056945f
C9165 ASIG5V.n12155 VSS 0.056945f
C9166 ASIG5V.n12156 VSS 0.056945f
C9167 ASIG5V.n12157 VSS 0.056945f
C9168 ASIG5V.n12159 VSS 0.056945f
C9169 ASIG5V.n12160 VSS 0.056945f
C9170 ASIG5V.n12161 VSS 0.056945f
C9171 ASIG5V.n12163 VSS 0.056945f
C9172 ASIG5V.n12164 VSS 0.056945f
C9173 ASIG5V.n12165 VSS 0.056945f
C9174 ASIG5V.n12166 VSS 0.056945f
C9175 ASIG5V.n12167 VSS 0.056945f
C9176 ASIG5V.n12168 VSS 0.056945f
C9177 ASIG5V.n12169 VSS 0.056945f
C9178 ASIG5V.n12171 VSS 0.056945f
C9179 ASIG5V.n12172 VSS 0.056945f
C9180 ASIG5V.n12173 VSS 0.056945f
C9181 ASIG5V.n12175 VSS 0.056945f
C9182 ASIG5V.n12176 VSS 0.056945f
C9183 ASIG5V.n12177 VSS 0.056945f
C9184 ASIG5V.n12178 VSS 0.056945f
C9185 ASIG5V.n12179 VSS 0.056945f
C9186 ASIG5V.n12180 VSS 0.056945f
C9187 ASIG5V.n12181 VSS 0.056945f
C9188 ASIG5V.n12183 VSS 0.056945f
C9189 ASIG5V.n12184 VSS 0.056945f
C9190 ASIG5V.n12185 VSS 0.056945f
C9191 ASIG5V.n12187 VSS 0.056945f
C9192 ASIG5V.n12188 VSS 0.056945f
C9193 ASIG5V.n12189 VSS 0.056945f
C9194 ASIG5V.n12190 VSS 0.056945f
C9195 ASIG5V.n12191 VSS 0.056945f
C9196 ASIG5V.n12192 VSS 0.056945f
C9197 ASIG5V.n12193 VSS 0.056945f
C9198 ASIG5V.n12195 VSS 0.056945f
C9199 ASIG5V.n12196 VSS 0.056945f
C9200 ASIG5V.n12197 VSS 0.056945f
C9201 ASIG5V.n12199 VSS 0.056945f
C9202 ASIG5V.n12200 VSS 0.056945f
C9203 ASIG5V.n12201 VSS 0.056945f
C9204 ASIG5V.n12202 VSS 0.056945f
C9205 ASIG5V.n12203 VSS 0.056945f
C9206 ASIG5V.n12204 VSS 0.056945f
C9207 ASIG5V.n12205 VSS 0.056945f
C9208 ASIG5V.n12207 VSS 0.056945f
C9209 ASIG5V.n12208 VSS 0.056945f
C9210 ASIG5V.n12209 VSS 0.056945f
C9211 ASIG5V.n12211 VSS 0.056945f
C9212 ASIG5V.n12212 VSS 0.056945f
C9213 ASIG5V.n12213 VSS 0.056945f
C9214 ASIG5V.n12214 VSS 0.056945f
C9215 ASIG5V.n12215 VSS 0.056945f
C9216 ASIG5V.n12216 VSS 0.056945f
C9217 ASIG5V.n12217 VSS 0.056945f
C9218 ASIG5V.n12219 VSS 0.056945f
C9219 ASIG5V.n12220 VSS 0.056945f
C9220 ASIG5V.n12221 VSS 0.056945f
C9221 ASIG5V.n12223 VSS 0.056945f
C9222 ASIG5V.n12224 VSS 0.056945f
C9223 ASIG5V.n12225 VSS 0.056945f
C9224 ASIG5V.n12226 VSS 0.056945f
C9225 ASIG5V.n12227 VSS 0.056945f
C9226 ASIG5V.n12228 VSS 0.056945f
C9227 ASIG5V.n12229 VSS 0.056945f
C9228 ASIG5V.n12231 VSS 0.056945f
C9229 ASIG5V.n12232 VSS 0.056945f
C9230 ASIG5V.n12233 VSS 0.056945f
C9231 ASIG5V.n12235 VSS 0.056945f
C9232 ASIG5V.n12236 VSS 0.056945f
C9233 ASIG5V.n12237 VSS 0.056945f
C9234 ASIG5V.n12238 VSS 0.056945f
C9235 ASIG5V.n12239 VSS 0.056945f
C9236 ASIG5V.n12240 VSS 0.056945f
C9237 ASIG5V.n12241 VSS 0.056945f
C9238 ASIG5V.n12243 VSS 0.056945f
C9239 ASIG5V.n12244 VSS 0.056945f
C9240 ASIG5V.n12245 VSS 0.056945f
C9241 ASIG5V.n12247 VSS 0.056945f
C9242 ASIG5V.n12248 VSS 0.056945f
C9243 ASIG5V.n12249 VSS 0.056945f
C9244 ASIG5V.n12250 VSS 0.056945f
C9245 ASIG5V.n12251 VSS 0.056945f
C9246 ASIG5V.n12252 VSS 0.056945f
C9247 ASIG5V.n12253 VSS 0.056945f
C9248 ASIG5V.n12255 VSS 0.056945f
C9249 ASIG5V.n12256 VSS 0.056945f
C9250 ASIG5V.n12257 VSS 0.056945f
C9251 ASIG5V.n12259 VSS 0.056945f
C9252 ASIG5V.n12260 VSS 0.056945f
C9253 ASIG5V.n12261 VSS 0.056945f
C9254 ASIG5V.n12262 VSS 0.056945f
C9255 ASIG5V.n12263 VSS 0.056945f
C9256 ASIG5V.n12264 VSS 0.056945f
C9257 ASIG5V.n12265 VSS 0.056945f
C9258 ASIG5V.n12267 VSS 0.036092f
C9259 ASIG5V.n12268 VSS 0.439183f
C9260 ASIG5V.n12269 VSS 0.924595f
C9261 ASIG5V.n12270 VSS 0.043486f
C9262 ASIG5V.n12271 VSS 0.043486f
C9263 ASIG5V.n12272 VSS 0.037979f
C9264 ASIG5V.n12273 VSS 0.052746f
C9265 ASIG5V.n12274 VSS 0.062513f
C9266 ASIG5V.n12275 VSS 0.065343f
C9267 ASIG5V.n12276 VSS 0.074818f
C9268 ASIG5V.n12277 VSS 0.074818f
C9269 ASIG5V.n12278 VSS 0.955415f
C9270 ASIG5V.n12279 VSS 0.485412f
C9271 ASIG5V.n12280 VSS 0.100173f
C9272 ASIG5V.n12281 VSS 0.100173f
C9273 ASIG5V.n12282 VSS 0.089417f
C9274 ASIG5V.n12283 VSS 0.07229f
C9275 ASIG5V.n12284 VSS 0.056474f
C9276 ASIG5V.n12285 VSS 0.09726f
C9277 ASIG5V.n12286 VSS 0.108961f
C9278 ASIG5V.n12287 VSS 0.108961f
C9279 ASIG5V.n12288 VSS 0.608692f
C9280 ASIG5V.n12289 VSS 0.955415f
C9281 ASIG5V.n12290 VSS 0.076709f
C9282 ASIG5V.n12291 VSS 0.067796f
C9283 ASIG5V.n12292 VSS 0.067796f
C9284 ASIG5V.n12293 VSS 0.05921f
C9285 ASIG5V.n12294 VSS 0.052746f
C9286 ASIG5V.n12295 VSS 0.047722f
C9287 ASIG5V.n12296 VSS 0.056945f
C9288 ASIG5V.n12297 VSS 0.056945f
C9289 ASIG5V.n12298 VSS 0.056945f
C9290 ASIG5V.n12300 VSS 0.036092f
C9291 ASIG5V.n12301 VSS 0.778201f
C9292 ASIG5V.n12302 VSS 0.770496f
C9293 ASIG5V.n12303 VSS 0.057995f
C9294 ASIG5V.n12304 VSS 0.057995f
C9295 ASIG5V.n12305 VSS 0.051768f
C9296 ASIG5V.n12306 VSS 0.07229f
C9297 ASIG5V.n12307 VSS 0.094123f
C9298 ASIG5V.n12308 VSS 0.105446f
C9299 ASIG5V.n12309 VSS 0.105446f
C9300 ASIG5V.n12310 VSS 0.770496f
C9301 ASIG5V.n12311 VSS 0.955415f
C9302 ASIG5V.n12312 VSS 0.076709f
C9303 ASIG5V.n12313 VSS 0.060773f
C9304 ASIG5V.n12314 VSS 0.060773f
C9305 ASIG5V.n12315 VSS 0.053077f
C9306 ASIG5V.n12316 VSS 0.052746f
C9307 ASIG5V.n12317 VSS 0.047722f
C9308 ASIG5V.n12318 VSS 0.056945f
C9309 ASIG5V.n12319 VSS 0.056945f
C9310 ASIG5V.n12320 VSS 0.056945f
C9311 ASIG5V.n12322 VSS 0.036092f
C9312 ASIG5V.n12323 VSS 0.362133f
C9313 ASIG5V.n12324 VSS 0.99394f
C9314 ASIG5V.n12325 VSS 0.070297f
C9315 ASIG5V.n12326 VSS 0.070297f
C9316 ASIG5V.n12327 VSS 0.059611f
C9317 ASIG5V.n12328 VSS 0.513832f
C9318 ASIG5V.n12329 VSS 0.06131f
C9319 ASIG5V.n12330 VSS 0.083142f
C9320 ASIG5V.n12331 VSS 0.093144f
C9321 ASIG5V.n12332 VSS 0.093144f
C9322 ASIG5V.n12333 VSS 0.108961f
C9323 ASIG5V.n12334 VSS 0.082599f
C9324 ASIG5V.n12335 VSS 0.082599f
C9325 ASIG5V.n12336 VSS 0.073729f
C9326 ASIG5V.n12337 VSS 0.07229f
C9327 ASIG5V.n12338 VSS 0.052133f
C9328 ASIG5V.n12339 VSS 0.056945f
C9329 ASIG5V.n12340 VSS 0.056945f
C9330 ASIG5V.n12341 VSS 0.056945f
C9331 ASIG5V.n12342 VSS 0.056945f
C9332 ASIG5V.n12343 VSS 0.056945f
C9333 ASIG5V.n12344 VSS 0.056945f
C9334 ASIG5V.n12345 VSS 0.056945f
C9335 ASIG5V.n12346 VSS 0.056945f
C9336 ASIG5V.n12347 VSS 0.056945f
C9337 ASIG5V.n12348 VSS 0.056945f
C9338 ASIG5V.n12349 VSS 0.056945f
C9339 ASIG5V.n12350 VSS 0.056945f
C9340 ASIG5V.n12351 VSS 0.056945f
C9341 ASIG5V.n12352 VSS 0.056945f
C9342 ASIG5V.n12353 VSS 0.056945f
C9343 ASIG5V.n12354 VSS 0.056945f
C9344 ASIG5V.n12355 VSS 0.056945f
C9345 ASIG5V.n12356 VSS 0.056945f
C9346 ASIG5V.n12357 VSS 0.056945f
C9347 ASIG5V.n12358 VSS 0.056945f
C9348 ASIG5V.n12359 VSS 0.056945f
C9349 ASIG5V.n12360 VSS 0.056945f
C9350 ASIG5V.n12361 VSS 0.056945f
C9351 ASIG5V.n12362 VSS 0.056945f
C9352 ASIG5V.n12363 VSS 0.056945f
C9353 ASIG5V.n12364 VSS 0.056945f
C9354 ASIG5V.n12365 VSS 0.056945f
C9355 ASIG5V.n12366 VSS 0.056945f
C9356 ASIG5V.n12367 VSS 0.056945f
C9357 ASIG5V.n12368 VSS 0.056945f
C9358 ASIG5V.n12369 VSS 0.056945f
C9359 ASIG5V.n12370 VSS 0.056945f
C9360 ASIG5V.n12371 VSS 0.056945f
C9361 ASIG5V.n12372 VSS 0.056945f
C9362 ASIG5V.n12373 VSS 0.056945f
C9363 ASIG5V.n12374 VSS 0.056945f
C9364 ASIG5V.n12375 VSS 0.056945f
C9365 ASIG5V.n12376 VSS 0.056945f
C9366 ASIG5V.n12377 VSS 0.056945f
C9367 ASIG5V.n12378 VSS 0.056945f
C9368 ASIG5V.n12379 VSS 0.056945f
C9369 ASIG5V.n12380 VSS 0.056945f
C9370 ASIG5V.n12381 VSS 0.056945f
C9371 ASIG5V.n12382 VSS 0.056945f
C9372 ASIG5V.n12383 VSS 0.056945f
C9373 ASIG5V.n12384 VSS 0.056945f
C9374 ASIG5V.n12385 VSS 0.056945f
C9375 ASIG5V.n12386 VSS 0.056945f
C9376 ASIG5V.n12387 VSS 0.056945f
C9377 ASIG5V.n12388 VSS 0.056945f
C9378 ASIG5V.n12389 VSS 0.056945f
C9379 ASIG5V.n12390 VSS 0.056945f
C9380 ASIG5V.n12391 VSS 0.056945f
C9381 ASIG5V.n12392 VSS 0.056945f
C9382 ASIG5V.n12393 VSS 0.056945f
C9383 ASIG5V.n12394 VSS 0.056945f
C9384 ASIG5V.n12395 VSS 0.056945f
C9385 ASIG5V.n12396 VSS 0.056945f
C9386 ASIG5V.n12397 VSS 0.056945f
C9387 ASIG5V.n12398 VSS 0.056945f
C9388 ASIG5V.n12399 VSS 0.056945f
C9389 ASIG5V.n12400 VSS 0.056945f
C9390 ASIG5V.n12401 VSS 0.056945f
C9391 ASIG5V.n12402 VSS 0.056945f
C9392 ASIG5V.n12403 VSS 0.056945f
C9393 ASIG5V.n12404 VSS 0.056945f
C9394 ASIG5V.n12405 VSS 0.056945f
C9395 ASIG5V.n12406 VSS 0.056945f
C9396 ASIG5V.n12407 VSS 0.056945f
C9397 ASIG5V.n12408 VSS 0.056945f
C9398 ASIG5V.n12409 VSS 0.056945f
C9399 ASIG5V.n12410 VSS 0.056945f
C9400 ASIG5V.n12411 VSS 0.056945f
C9401 ASIG5V.n12412 VSS 0.056945f
C9402 ASIG5V.n12413 VSS 0.056945f
C9403 ASIG5V.n12414 VSS 0.056945f
C9404 ASIG5V.n12415 VSS 0.056945f
C9405 ASIG5V.n12416 VSS 0.056945f
C9406 ASIG5V.n12417 VSS 0.056945f
C9407 ASIG5V.n12418 VSS 0.056945f
C9408 ASIG5V.n12419 VSS 0.056945f
C9409 ASIG5V.n12420 VSS 0.056945f
C9410 ASIG5V.n12421 VSS 0.056945f
C9411 ASIG5V.n12422 VSS 0.056945f
C9412 ASIG5V.n12423 VSS 0.056945f
C9413 ASIG5V.n12424 VSS 0.056945f
C9414 ASIG5V.n12425 VSS 0.056945f
C9415 ASIG5V.n12426 VSS 0.056945f
C9416 ASIG5V.n12427 VSS 0.056945f
C9417 ASIG5V.n12428 VSS 0.056945f
C9418 ASIG5V.n12429 VSS 0.056945f
C9419 ASIG5V.n12430 VSS 0.056945f
C9420 ASIG5V.n12431 VSS 0.056945f
C9421 ASIG5V.n12432 VSS 0.056945f
C9422 ASIG5V.n12433 VSS 0.056945f
C9423 ASIG5V.n12434 VSS 0.056945f
C9424 ASIG5V.n12435 VSS 0.056945f
C9425 ASIG5V.n12436 VSS 0.056945f
C9426 ASIG5V.n12437 VSS 0.056945f
C9427 ASIG5V.n12438 VSS 0.056945f
C9428 ASIG5V.n12439 VSS 0.056945f
C9429 ASIG5V.n12440 VSS 0.056945f
C9430 ASIG5V.n12441 VSS 0.056945f
C9431 ASIG5V.n12442 VSS 0.056945f
C9432 ASIG5V.n12443 VSS 0.056945f
C9433 ASIG5V.n12444 VSS 0.056945f
C9434 ASIG5V.n12445 VSS 0.056945f
C9435 ASIG5V.n12446 VSS 0.056945f
C9436 ASIG5V.n12447 VSS 0.056945f
C9437 ASIG5V.n12448 VSS 0.056945f
C9438 ASIG5V.n12449 VSS 0.056945f
C9439 ASIG5V.n12450 VSS 0.056945f
C9440 ASIG5V.n12451 VSS 0.056945f
C9441 ASIG5V.n12452 VSS 0.056945f
C9442 ASIG5V.n12453 VSS 0.056945f
C9443 ASIG5V.n12454 VSS 0.056945f
C9444 ASIG5V.n12455 VSS 0.056945f
C9445 ASIG5V.n12456 VSS 0.056945f
C9446 ASIG5V.n12457 VSS 0.056945f
C9447 ASIG5V.n12458 VSS 0.056945f
C9448 ASIG5V.n12459 VSS 0.056945f
C9449 ASIG5V.n12460 VSS 0.056945f
C9450 ASIG5V.n12461 VSS 0.056945f
C9451 ASIG5V.n12462 VSS 0.056945f
C9452 ASIG5V.n12463 VSS 0.056945f
C9453 ASIG5V.n12464 VSS 0.056945f
C9454 ASIG5V.n12465 VSS 0.056945f
C9455 ASIG5V.n12466 VSS 0.056945f
C9456 ASIG5V.n12467 VSS 0.056945f
C9457 ASIG5V.n12468 VSS 0.056945f
C9458 ASIG5V.n12469 VSS 0.056945f
C9459 ASIG5V.n12470 VSS 0.056945f
C9460 ASIG5V.n12471 VSS 0.056945f
C9461 ASIG5V.n12472 VSS 0.056945f
C9462 ASIG5V.n12473 VSS 0.056945f
C9463 ASIG5V.n12474 VSS 0.056945f
C9464 ASIG5V.n12475 VSS 0.056945f
C9465 ASIG5V.n12476 VSS 0.056945f
C9466 ASIG5V.n12477 VSS 0.056945f
C9467 ASIG5V.n12478 VSS 0.056945f
C9468 ASIG5V.n12479 VSS 0.056945f
C9469 ASIG5V.n12480 VSS 0.056945f
C9470 ASIG5V.n12481 VSS 0.056945f
C9471 ASIG5V.n12482 VSS 0.056945f
C9472 ASIG5V.n12483 VSS 0.056945f
C9473 ASIG5V.n12484 VSS 0.056945f
C9474 ASIG5V.n12485 VSS 0.056945f
C9475 ASIG5V.n12486 VSS 0.056945f
C9476 ASIG5V.n12487 VSS 0.056945f
C9477 ASIG5V.n12488 VSS 0.056945f
C9478 ASIG5V.n12489 VSS 0.056945f
C9479 ASIG5V.n12490 VSS 0.056945f
C9480 ASIG5V.n12491 VSS 0.056945f
C9481 ASIG5V.n12492 VSS 0.056945f
C9482 ASIG5V.n12493 VSS 0.056945f
C9483 ASIG5V.n12494 VSS 0.056945f
C9484 ASIG5V.n12495 VSS 0.056945f
C9485 ASIG5V.n12496 VSS 0.056945f
C9486 ASIG5V.n12497 VSS 0.056945f
C9487 ASIG5V.n12498 VSS 0.056945f
C9488 ASIG5V.n12499 VSS 0.056945f
C9489 ASIG5V.n12500 VSS 0.056945f
C9490 ASIG5V.n12501 VSS 0.056945f
C9491 ASIG5V.n12502 VSS 0.056945f
C9492 ASIG5V.n12503 VSS 0.056945f
C9493 ASIG5V.n12504 VSS 0.056945f
C9494 ASIG5V.n12505 VSS 0.056945f
C9495 ASIG5V.n12506 VSS 0.056945f
C9496 ASIG5V.n12507 VSS 0.056945f
C9497 ASIG5V.n12508 VSS 0.056945f
C9498 ASIG5V.n12509 VSS 0.056945f
C9499 ASIG5V.n12510 VSS 0.056945f
C9500 ASIG5V.n12511 VSS 0.056945f
C9501 ASIG5V.n12512 VSS 0.056945f
C9502 ASIG5V.n12513 VSS 0.056945f
C9503 ASIG5V.n12514 VSS 0.056945f
C9504 ASIG5V.n12515 VSS 0.056945f
C9505 ASIG5V.n12516 VSS 0.056945f
C9506 ASIG5V.n12517 VSS 0.056945f
C9507 ASIG5V.n12518 VSS 0.056945f
C9508 ASIG5V.n12519 VSS 0.056945f
C9509 ASIG5V.n12520 VSS 0.056945f
C9510 ASIG5V.n12521 VSS 0.056945f
C9511 ASIG5V.n12522 VSS 0.047722f
C9512 ASIG5V.n12523 VSS 0.036092f
C9513 ASIG5V.n12524 VSS 0.036092f
C9514 ASIG5V.n12525 VSS 0.955415f
C9515 ASIG5V.n12526 VSS 0.036092f
C9516 ASIG5V.n12528 VSS 0.192624f
C9517 ASIG5V.n12529 VSS 0.886071f
C9518 ASIG5V.n12530 VSS 0.061313f
C9519 ASIG5V.n12531 VSS 0.061313f
C9520 ASIG5V.n12532 VSS 0.053548f
C9521 ASIG5V.n12533 VSS 0.066995f
C9522 ASIG5V.n12534 VSS 0.04081f
C9523 ASIG5V.n12535 VSS 0.046728f
C9524 ASIG5V.n12536 VSS 0.046728f
C9525 ASIG5V.n12537 VSS 0.392953f
C9526 DVSS.n0 VSS 0.039859f
C9527 DVSS.n1 VSS 1.32112f
C9528 DVSS.n2 VSS 0.184347f
C9529 DVSS.n3 VSS 0.154453f
C9530 DVSS.n4 VSS 0.154453f
C9531 DVSS.n5 VSS 0.154453f
C9532 DVSS.n17 VSS 0.099554f
C9533 DVSS.n19 VSS 0.176874f
C9534 DVSS.n20 VSS 0.353747f
C9535 DVSS.n21 VSS 0.353747f
C9536 DVSS.n22 VSS 0.353747f
C9537 DVSS.n23 VSS 0.353747f
C9538 DVSS.n24 VSS 0.154453f
C9539 DVSS.n25 VSS 0.022779f
C9540 DVSS.n26 VSS 0.022779f
C9541 DVSS.n27 VSS 0.022779f
C9542 DVSS.n28 VSS 0.022779f
C9543 DVSS.n29 VSS 0.022779f
C9544 DVSS.n30 VSS 0.022779f
C9545 DVSS.n31 VSS 0.022779f
C9546 DVSS.n32 VSS 0.022779f
C9547 DVSS.n33 VSS 0.022779f
C9548 DVSS.n34 VSS 0.022779f
C9549 DVSS.n35 VSS 0.022779f
C9550 DVSS.n36 VSS 0.022779f
C9551 DVSS.n37 VSS 0.022779f
C9552 DVSS.n38 VSS 0.022779f
C9553 DVSS.n39 VSS 0.022779f
C9554 DVSS.n40 VSS 0.022779f
C9555 DVSS.n41 VSS 0.022779f
C9556 DVSS.n42 VSS 0.022779f
C9557 DVSS.n43 VSS 0.022779f
C9558 DVSS.n44 VSS 0.022779f
C9559 DVSS.n45 VSS 0.022779f
C9560 DVSS.n46 VSS 0.022779f
C9561 DVSS.n47 VSS 0.022779f
C9562 DVSS.n48 VSS 0.026154f
C9563 DVSS.n49 VSS 0.176874f
C9564 DVSS.n50 VSS 0.176874f
C9565 DVSS.n51 VSS 0.036489f
C9566 DVSS.n52 VSS 0.154453f
C9567 DVSS.n53 VSS 0.353747f
C9568 DVSS.n54 VSS 0.353747f
C9569 DVSS.n55 VSS 0.353747f
C9570 DVSS.n56 VSS 0.353747f
C9571 DVSS.n57 VSS 0.323853f
C9572 DVSS.n58 VSS 0.323853f
C9573 DVSS.n59 VSS 0.675109f
C9574 DVSS.n60 VSS 0.353747f
C9575 DVSS.n61 VSS 0.353747f
C9576 DVSS.n62 VSS 0.163172f
C9577 DVSS.n63 VSS 0.425991f
C9578 DVSS.n64 VSS 0.206768f
C9579 DVSS.n65 VSS 0.323853f
C9580 DVSS.n66 VSS 0.353747f
C9581 DVSS.n67 VSS 0.353747f
C9582 DVSS.n68 VSS 0.353747f
C9583 DVSS.n69 VSS 0.353747f
C9584 DVSS.n70 VSS 0.287731f
C9585 DVSS.n71 VSS 0.154453f
C9586 DVSS.n72 VSS 0.353747f
C9587 DVSS.n73 VSS 0.353747f
C9588 DVSS.n74 VSS 0.154453f
C9589 DVSS.n75 VSS 0.310152f
C9590 DVSS.n76 VSS 0.353747f
C9591 DVSS.n77 VSS 0.353747f
C9592 DVSS.n78 VSS 0.267802f
C9593 DVSS.n79 VSS 0.353747f
C9594 DVSS.n80 VSS 0.353747f
C9595 DVSS.n81 VSS 0.227943f
C9596 DVSS.n82 VSS 0.154453f
C9597 DVSS.n83 VSS 0.353747f
C9598 DVSS.n84 VSS 0.779994f
C9599 DVSS.n85 VSS 0.154453f
C9600 DVSS.n86 VSS 0.052308f
C9601 DVSS.n87 VSS 0.052308f
C9602 DVSS.n88 VSS 0.052308f
C9603 DVSS.n89 VSS 0.052308f
C9604 DVSS.n90 VSS 0.052308f
C9605 DVSS.n91 VSS 0.052308f
C9606 DVSS.n92 VSS 0.052308f
C9607 DVSS.n93 VSS 0.052308f
C9608 DVSS.n94 VSS 0.052308f
C9609 DVSS.n95 VSS 0.052308f
C9610 DVSS.n96 VSS 0.052308f
C9611 DVSS.n98 VSS 0.779994f
C9612 DVSS.n99 VSS 0.176874f
C9613 DVSS.n100 VSS 0.145734f
C9614 DVSS.n101 VSS 0.052308f
C9615 DVSS.n102 VSS 0.052308f
C9616 DVSS.n103 VSS 0.052308f
C9617 DVSS.n104 VSS 0.052308f
C9618 DVSS.n105 VSS 0.052308f
C9619 DVSS.n106 VSS 0.052308f
C9620 DVSS.n107 VSS 0.052308f
C9621 DVSS.n108 VSS 0.052308f
C9622 DVSS.n109 VSS 0.052308f
C9623 DVSS.n110 VSS 0.052308f
C9624 DVSS.n111 VSS 0.052308f
C9625 DVSS.n112 VSS 0.438291f
C9626 DVSS.n113 VSS 0.154453f
C9627 DVSS.n115 VSS 0.052308f
C9628 DVSS.n117 VSS 0.052308f
C9629 DVSS.n119 VSS 0.052308f
C9630 DVSS.n121 VSS 0.052308f
C9631 DVSS.n123 VSS 0.052308f
C9632 DVSS.n125 VSS 0.052308f
C9633 DVSS.n127 VSS 0.052308f
C9634 DVSS.n129 VSS 0.052308f
C9635 DVSS.n131 VSS 0.052308f
C9636 DVSS.n133 VSS 0.052308f
C9637 DVSS.n134 VSS 0.353747f
C9638 DVSS.n135 VSS 0.154453f
C9639 DVSS.n136 VSS 0.353747f
C9640 DVSS.n137 VSS 0.353747f
C9641 DVSS.n138 VSS 0.353747f
C9642 DVSS.n139 VSS 0.310152f
C9643 DVSS.n140 VSS 0.353747f
C9644 DVSS.n141 VSS 0.353747f
C9645 DVSS.n142 VSS 0.353747f
C9646 DVSS.n143 VSS 0.176874f
C9647 DVSS.n155 VSS 0.438291f
C9648 DVSS.n156 VSS 0.026154f
C9649 DVSS.n157 VSS 0.176874f
C9650 DVSS.n158 VSS 0.042395f
C9651 DVSS.n159 VSS 0.353747f
C9652 DVSS.n160 VSS 0.353747f
C9653 DVSS.n161 VSS 0.353747f
C9654 DVSS.n162 VSS 0.425991f
C9655 DVSS.n163 VSS 0.353747f
C9656 DVSS.n164 VSS 0.353747f
C9657 DVSS.n165 VSS 0.154453f
C9658 DVSS.n170 VSS 0.051254f
C9659 DVSS.n175 VSS 0.052308f
C9660 DVSS.n176 VSS 0.022779f
C9661 DVSS.n177 VSS 0.249729f
C9662 DVSS.n178 VSS 0.026998f
C9663 DVSS.n179 VSS 0.03206f
C9664 DVSS.n180 VSS 0.022779f
C9665 DVSS.n181 VSS 0.026154f
C9666 DVSS.n183 VSS 0.176874f
C9667 DVSS.n184 VSS 0.176874f
C9668 DVSS.n185 VSS 0.041973f
C9669 DVSS.n186 VSS 0.154453f
C9670 DVSS.n187 VSS 0.041973f
C9671 DVSS.n188 VSS 0.030583f
C9672 DVSS.n189 VSS 0.353747f
C9673 DVSS.n190 VSS 0.353747f
C9674 DVSS.n191 VSS 0.353747f
C9675 DVSS.n192 VSS 0.353747f
C9676 DVSS.n193 VSS 0.353747f
C9677 DVSS.n194 VSS 0.353747f
C9678 DVSS.n195 VSS 0.353747f
C9679 DVSS.n196 VSS 0.353747f
C9680 DVSS.n197 VSS 0.353747f
C9681 DVSS.n198 VSS 0.353747f
C9682 DVSS.n199 VSS 0.353747f
C9683 DVSS.n200 VSS 0.353747f
C9684 DVSS.n201 VSS 0.353747f
C9685 DVSS.n202 VSS 0.353747f
C9686 DVSS.n203 VSS 0.353747f
C9687 DVSS.n204 VSS 0.154453f
C9688 DVSS.n209 VSS 0.051254f
C9689 DVSS.n214 VSS 0.052308f
C9690 DVSS.n215 VSS 0.022779f
C9691 DVSS.n216 VSS 0.249729f
C9692 DVSS.n217 VSS 0.026998f
C9693 DVSS.n218 VSS 0.03206f
C9694 DVSS.n219 VSS 0.022779f
C9695 DVSS.n220 VSS 0.026154f
C9696 DVSS.n222 VSS 0.176874f
C9697 DVSS.n223 VSS 0.176874f
C9698 DVSS.n224 VSS 0.041973f
C9699 DVSS.n225 VSS 0.154453f
C9700 DVSS.n226 VSS 0.041973f
C9701 DVSS.n227 VSS 0.030583f
C9702 DVSS.n228 VSS 0.353747f
C9703 DVSS.n229 VSS 0.353747f
C9704 DVSS.n230 VSS 0.353747f
C9705 DVSS.n231 VSS 0.313888f
C9706 DVSS.n232 VSS 0.313888f
C9707 DVSS.n233 VSS 0.216732f
C9708 DVSS.n234 VSS 0.425991f
C9709 DVSS.n235 VSS 0.216732f
C9710 DVSS.n236 VSS 0.353747f
C9711 DVSS.n237 VSS 0.675109f
C9712 DVSS.n238 VSS 0.313888f
C9713 DVSS.n239 VSS 0.353747f
C9714 DVSS.n240 VSS 0.353747f
C9715 DVSS.n241 VSS 0.353747f
C9716 DVSS.n242 VSS 0.353747f
C9717 DVSS.n243 VSS 0.154453f
C9718 DVSS.n244 VSS 0.154453f
C9719 DVSS.n245 VSS 0.154453f
C9720 DVSS.n246 VSS 0.353747f
C9721 DVSS.n247 VSS 0.353747f
C9722 DVSS.n248 VSS 0.353747f
C9723 DVSS.n249 VSS 0.353747f
C9724 DVSS.n250 VSS 0.353747f
C9725 DVSS.n251 VSS 0.353747f
C9726 DVSS.n252 VSS 0.353747f
C9727 DVSS.n253 VSS 0.353747f
C9728 DVSS.n254 VSS 0.353747f
C9729 DVSS.n255 VSS 0.353747f
C9730 DVSS.n256 VSS 0.353747f
C9731 DVSS.n257 VSS 0.353747f
C9732 DVSS.n258 VSS 0.353747f
C9733 DVSS.n259 VSS 0.353747f
C9734 DVSS.n260 VSS 0.353747f
C9735 DVSS.n261 VSS 0.353747f
C9736 DVSS.n262 VSS 0.353747f
C9737 DVSS.n263 VSS 0.353747f
C9738 DVSS.n264 VSS 0.353747f
C9739 DVSS.n265 VSS 0.154453f
C9740 DVSS.n266 VSS 0.154453f
C9741 DVSS.n267 VSS 0.176874f
C9742 DVSS.n268 VSS 0.031427f
C9743 DVSS.n269 VSS 0.425991f
C9744 DVSS.n270 VSS 0.675109f
C9745 DVSS.n271 VSS 0.163172f
C9746 DVSS.n273 VSS 0.052308f
C9747 DVSS.n285 VSS 0.176874f
C9748 DVSS.n286 VSS 0.154453f
C9749 DVSS.n287 VSS 0.176874f
C9750 DVSS.n288 VSS 0.287731f
C9751 DVSS.n289 VSS 0.052308f
C9752 DVSS.n290 VSS 0.052308f
C9753 DVSS.n291 VSS 0.052308f
C9754 DVSS.n292 VSS 0.052308f
C9755 DVSS.n293 VSS 0.052308f
C9756 DVSS.n294 VSS 0.052308f
C9757 DVSS.n295 VSS 0.052308f
C9758 DVSS.n296 VSS 0.052308f
C9759 DVSS.n297 VSS 0.052308f
C9760 DVSS.n298 VSS 0.052308f
C9761 DVSS.n299 VSS 0.052308f
C9762 DVSS.n300 VSS 0.154453f
C9763 DVSS.n302 VSS 0.052308f
C9764 DVSS.n304 VSS 0.052308f
C9765 DVSS.n306 VSS 0.052308f
C9766 DVSS.n308 VSS 0.052308f
C9767 DVSS.n310 VSS 0.052308f
C9768 DVSS.n312 VSS 0.052308f
C9769 DVSS.n314 VSS 0.052308f
C9770 DVSS.n316 VSS 0.052308f
C9771 DVSS.n318 VSS 0.052308f
C9772 DVSS.n320 VSS 0.052308f
C9773 DVSS.n322 VSS 0.052308f
C9774 DVSS.n325 VSS 0.393287f
C9775 DVSS.n326 VSS 0.048189f
C9776 DVSS.n327 VSS 0.048189f
C9777 DVSS.n328 VSS 0.052308f
C9778 DVSS.n330 VSS 0.046402f
C9779 DVSS.n331 VSS 0.05737f
C9780 DVSS.n332 VSS 0.029924f
C9781 DVSS.n334 VSS 0.045559f
C9782 DVSS.n336 VSS -1.4011f
C9783 DVSS.n337 VSS 0.028052f
C9784 DVSS.n338 VSS 0.041971f
C9785 DVSS.n339 VSS 0.022779f
C9786 DVSS.n340 VSS 0.176874f
C9787 DVSS.n341 VSS 0.176874f
C9788 DVSS.n342 VSS 0.154453f
C9789 DVSS.n343 VSS 0.176874f
C9790 DVSS.n344 VSS 0.022779f
C9791 DVSS.n345 VSS 0.022779f
C9792 DVSS.n346 VSS 0.022779f
C9793 DVSS.n347 VSS 0.022779f
C9794 DVSS.n348 VSS 0.022779f
C9795 DVSS.n349 VSS 0.022779f
C9796 DVSS.n350 VSS 0.022779f
C9797 DVSS.n351 VSS 0.022779f
C9798 DVSS.n352 VSS 0.022779f
C9799 DVSS.n353 VSS 0.022779f
C9800 DVSS.n354 VSS 0.022779f
C9801 DVSS.n355 VSS 0.022779f
C9802 DVSS.n356 VSS 0.022779f
C9803 DVSS.n357 VSS 0.022779f
C9804 DVSS.n358 VSS 0.022779f
C9805 DVSS.n359 VSS 0.022779f
C9806 DVSS.n360 VSS 0.022779f
C9807 DVSS.n361 VSS 0.022779f
C9808 DVSS.n362 VSS 0.022779f
C9809 DVSS.n363 VSS 0.022779f
C9810 DVSS.n364 VSS 0.022779f
C9811 DVSS.n365 VSS 0.029924f
C9812 DVSS.n366 VSS 0.031005f
C9813 DVSS.n367 VSS 0.031427f
C9814 DVSS.n368 VSS 0.052308f
C9815 DVSS.n369 VSS 0.031427f
C9816 DVSS.n370 VSS 0.052308f
C9817 DVSS.n372 VSS 0.026354f
C9818 DVSS.n373 VSS 0.043865f
C9819 DVSS.n374 VSS 0.035198f
C9820 DVSS.n375 VSS 0.021932f
C9821 DVSS.n377 VSS 0.048189f
C9822 DVSS.n378 VSS 0.047218f
C9823 DVSS.n379 VSS 6.77029f
C9824 DVSS.n380 VSS 1.13994f
C9825 DVSS.n381 VSS 78.2638f
C9826 DVSS.n382 VSS 0.047218f
C9827 DVSS.n383 VSS 0.038912f
C9828 DVSS.n384 VSS 0.048189f
C9829 DVSS.n386 VSS 0.030953f
C9830 DVSS.n388 VSS 0.043865f
C9831 DVSS.n392 VSS 0.176874f
C9832 DVSS.n393 VSS 0.176874f
C9833 DVSS.n394 VSS 0.287731f
C9834 DVSS.n395 VSS 0.052308f
C9835 DVSS.n396 VSS 0.052308f
C9836 DVSS.n397 VSS 0.052308f
C9837 DVSS.n398 VSS 0.052308f
C9838 DVSS.n399 VSS 0.052308f
C9839 DVSS.n400 VSS 0.052308f
C9840 DVSS.n401 VSS 0.052308f
C9841 DVSS.n402 VSS 0.052308f
C9842 DVSS.n403 VSS 0.052308f
C9843 DVSS.n404 VSS 0.052308f
C9844 DVSS.n405 VSS 0.052308f
C9845 DVSS.n407 VSS 0.176874f
C9846 DVSS.n408 VSS 0.176874f
C9847 DVSS.n409 VSS 0.287731f
C9848 DVSS.n410 VSS 0.052308f
C9849 DVSS.n411 VSS 0.052308f
C9850 DVSS.n412 VSS 0.052308f
C9851 DVSS.n413 VSS 0.052308f
C9852 DVSS.n414 VSS 0.052308f
C9853 DVSS.n415 VSS 0.052308f
C9854 DVSS.n416 VSS 0.052308f
C9855 DVSS.n417 VSS 0.052308f
C9856 DVSS.n418 VSS 0.052308f
C9857 DVSS.n419 VSS 0.052308f
C9858 DVSS.n420 VSS 0.052308f
C9859 DVSS.n421 VSS 0.031427f
C9860 DVSS.n424 VSS 0.052308f
C9861 DVSS.n426 VSS 0.052308f
C9862 DVSS.n428 VSS 0.052308f
C9863 DVSS.n430 VSS 0.052308f
C9864 DVSS.n432 VSS 0.052308f
C9865 DVSS.n434 VSS 0.052308f
C9866 DVSS.n436 VSS 0.052308f
C9867 DVSS.n438 VSS 0.052308f
C9868 DVSS.n440 VSS 0.052308f
C9869 DVSS.n442 VSS 0.052308f
C9870 DVSS.n443 VSS 0.310152f
C9871 DVSS.n453 VSS 0.176874f
C9872 DVSS.n456 VSS 0.052308f
C9873 DVSS.n457 VSS 0.176874f
C9874 DVSS.n458 VSS 0.099554f
C9875 DVSS.n459 VSS 0.099554f
C9876 DVSS.n460 VSS 0.154453f
C9877 DVSS.n462 VSS 0.052308f
C9878 DVSS.n464 VSS 0.052308f
C9879 DVSS.n466 VSS 0.052308f
C9880 DVSS.n468 VSS 0.052308f
C9881 DVSS.n470 VSS 0.052308f
C9882 DVSS.n472 VSS 0.052308f
C9883 DVSS.n474 VSS 0.052308f
C9884 DVSS.n476 VSS 0.052308f
C9885 DVSS.n478 VSS 0.052308f
C9886 DVSS.n480 VSS 0.052308f
C9887 DVSS.n481 VSS 0.353747f
C9888 DVSS.n482 VSS 0.154453f
C9889 DVSS.n483 VSS 0.353747f
C9890 DVSS.n484 VSS 0.353747f
C9891 DVSS.n485 VSS 0.353747f
C9892 DVSS.n486 VSS 0.425991f
C9893 DVSS.n487 VSS 0.353747f
C9894 DVSS.n488 VSS 0.216732f
C9895 DVSS.n489 VSS 0.353747f
C9896 DVSS.n490 VSS 0.353747f
C9897 DVSS.n491 VSS 0.353747f
C9898 DVSS.n492 VSS 0.353747f
C9899 DVSS.n493 VSS 0.353747f
C9900 DVSS.n494 VSS 0.353747f
C9901 DVSS.n495 VSS 0.176874f
C9902 DVSS.n496 VSS 0.353747f
C9903 DVSS.n497 VSS 0.353747f
C9904 DVSS.n498 VSS 0.353747f
C9905 DVSS.n499 VSS 0.176874f
C9906 DVSS.n500 VSS 0.154453f
C9907 DVSS.n502 VSS 0.176874f
C9908 DVSS.n503 VSS 0.239153f
C9909 DVSS.n504 VSS 0.043865f
C9910 DVSS.n505 VSS 0.043865f
C9911 DVSS.n506 VSS 0.043865f
C9912 DVSS.n507 VSS 0.043865f
C9913 DVSS.n508 VSS 0.043865f
C9914 DVSS.n509 VSS 0.043865f
C9915 DVSS.n510 VSS 0.043865f
C9916 DVSS.n511 VSS 0.043865f
C9917 DVSS.n512 VSS 0.043865f
C9918 DVSS.n513 VSS 0.043865f
C9919 DVSS.n514 VSS 0.043865f
C9920 DVSS.n515 VSS 0.026354f
C9921 DVSS.n516 VSS 0.154453f
C9922 DVSS.n518 VSS 0.043865f
C9923 DVSS.n520 VSS 0.043865f
C9924 DVSS.n522 VSS 0.043865f
C9925 DVSS.n524 VSS 0.043865f
C9926 DVSS.n526 VSS 0.043865f
C9927 DVSS.n528 VSS 0.043865f
C9928 DVSS.n530 VSS 0.043865f
C9929 DVSS.n532 VSS 0.043865f
C9930 DVSS.n534 VSS 0.043865f
C9931 DVSS.n536 VSS 0.043865f
C9932 DVSS.n537 VSS 0.353747f
C9933 DVSS.n538 VSS 0.353747f
C9934 DVSS.n539 VSS 0.353747f
C9935 DVSS.n540 VSS 0.353747f
C9936 DVSS.n541 VSS 0.336309f
C9937 DVSS.n542 VSS 0.353747f
C9938 DVSS.n543 VSS 0.353747f
C9939 DVSS.n544 VSS 0.353747f
C9940 DVSS.n545 VSS 0.353747f
C9941 DVSS.n546 VSS 0.353747f
C9942 DVSS.n547 VSS 0.353747f
C9943 DVSS.n548 VSS 0.353747f
C9944 DVSS.n549 VSS 0.353747f
C9945 DVSS.n550 VSS 0.353747f
C9946 DVSS.n551 VSS 0.353747f
C9947 DVSS.n552 VSS 0.353747f
C9948 DVSS.n553 VSS 0.353747f
C9949 DVSS.n554 VSS 0.353747f
C9950 DVSS.n555 VSS 0.353747f
C9951 DVSS.n556 VSS 0.353747f
C9952 DVSS.n557 VSS 0.353747f
C9953 DVSS.n558 VSS 0.353747f
C9954 DVSS.n559 VSS 0.154453f
C9955 DVSS.n560 VSS 0.04298f
C9956 DVSS.n561 VSS 0.025647f
C9957 DVSS.n566 VSS 0.019102f
C9958 DVSS.n567 VSS 0.209418f
C9959 DVSS.n568 VSS 0.02264f
C9960 DVSS.n569 VSS 0.026885f
C9961 DVSS.n570 VSS 0.019102f
C9962 DVSS.n575 VSS 0.239153f
C9963 DVSS.n576 VSS 0.043865f
C9964 DVSS.n577 VSS 0.043865f
C9965 DVSS.n578 VSS 0.043865f
C9966 DVSS.n579 VSS 0.043865f
C9967 DVSS.n580 VSS 0.043865f
C9968 DVSS.n581 VSS 0.043865f
C9969 DVSS.n582 VSS 0.043865f
C9970 DVSS.n583 VSS 0.353747f
C9971 DVSS.n584 VSS 0.353747f
C9972 DVSS.n585 VSS 0.353747f
C9973 DVSS.n586 VSS 0.353747f
C9974 DVSS.n587 VSS 0.154453f
C9975 DVSS.n588 VSS 0.04298f
C9976 DVSS.n589 VSS 0.025647f
C9977 DVSS.n594 VSS 0.019102f
C9978 DVSS.n595 VSS 0.209418f
C9979 DVSS.n596 VSS 0.02264f
C9980 DVSS.n597 VSS 0.026885f
C9981 DVSS.n598 VSS 0.019102f
C9982 DVSS.n603 VSS 0.021932f
C9983 DVSS.n605 VSS 0.176874f
C9984 DVSS.n606 VSS 0.035198f
C9985 DVSS.n607 VSS 0.341291f
C9986 DVSS.n608 VSS 0.035198f
C9987 DVSS.n609 VSS 0.043865f
C9988 DVSS.n610 VSS 0.043865f
C9989 DVSS.n611 VSS 0.043865f
C9990 DVSS.n612 VSS 0.043865f
C9991 DVSS.n613 VSS 0.043865f
C9992 DVSS.n614 VSS 0.043865f
C9993 DVSS.n616 VSS 0.043865f
C9994 DVSS.n617 VSS 0.353747f
C9995 DVSS.n618 VSS 0.353747f
C9996 DVSS.n619 VSS 0.353747f
C9997 DVSS.n620 VSS 0.353747f
C9998 DVSS.n621 VSS 0.353747f
C9999 DVSS.n622 VSS 0.353747f
C10000 DVSS.n623 VSS 0.353747f
C10001 DVSS.n624 VSS 0.303924f
C10002 DVSS.n625 VSS 0.303924f
C10003 DVSS.n626 VSS 0.675109f
C10004 DVSS.n627 VSS 0.353747f
C10005 DVSS.n628 VSS 0.353747f
C10006 DVSS.n629 VSS 0.226697f
C10007 DVSS.n630 VSS 0.425991f
C10008 DVSS.n631 VSS 0.226697f
C10009 DVSS.n632 VSS 0.303924f
C10010 DVSS.n633 VSS 0.353747f
C10011 DVSS.n634 VSS 0.353747f
C10012 DVSS.n635 VSS 0.353747f
C10013 DVSS.n636 VSS 0.353747f
C10014 DVSS.n637 VSS 0.353747f
C10015 DVSS.n638 VSS 0.353747f
C10016 DVSS.n639 VSS 0.353747f
C10017 DVSS.n640 VSS 0.353747f
C10018 DVSS.n641 VSS 0.353747f
C10019 DVSS.n642 VSS 0.353747f
C10020 DVSS.n643 VSS 0.353747f
C10021 DVSS.n644 VSS 0.341291f
C10022 DVSS.n645 VSS 0.353747f
C10023 DVSS.n646 VSS 0.353747f
C10024 DVSS.n647 VSS 0.154453f
C10025 DVSS.n648 VSS 0.026354f
C10026 DVSS.n662 VSS 0.176874f
C10027 DVSS.n663 VSS 0.341291f
C10028 DVSS.n664 VSS 0.043865f
C10029 DVSS.n665 VSS 0.043865f
C10030 DVSS.n666 VSS 0.043865f
C10031 DVSS.n667 VSS 0.043865f
C10032 DVSS.n668 VSS 0.043865f
C10033 DVSS.n669 VSS 0.043865f
C10034 DVSS.n670 VSS 0.043865f
C10035 DVSS.n671 VSS 0.043865f
C10036 DVSS.n672 VSS 0.043865f
C10037 DVSS.n673 VSS 0.043865f
C10038 DVSS.n674 VSS 0.043865f
C10039 DVSS.n675 VSS 0.154453f
C10040 DVSS.n677 VSS 0.043865f
C10041 DVSS.n679 VSS 0.043865f
C10042 DVSS.n681 VSS 0.043865f
C10043 DVSS.n683 VSS 0.043865f
C10044 DVSS.n685 VSS 0.043865f
C10045 DVSS.n687 VSS 0.043865f
C10046 DVSS.n689 VSS 0.043865f
C10047 DVSS.n691 VSS 0.043865f
C10048 DVSS.n693 VSS 0.043865f
C10049 DVSS.n695 VSS 0.043865f
C10050 DVSS.n697 VSS 0.043865f
C10051 DVSS.n700 VSS 0.048189f
C10052 DVSS.n701 VSS 0.052308f
C10053 DVSS.n702 VSS 0.046402f
C10054 DVSS.n704 VSS 0.052308f
C10055 DVSS.n705 VSS 0.036911f
C10056 DVSS.n707 VSS 0.048189f
C10057 DVSS.n708 VSS 0.052308f
C10058 DVSS.n709 VSS 0.046402f
C10059 DVSS.n711 VSS 0.052308f
C10060 DVSS.n712 VSS 0.036911f
C10061 DVSS.n714 VSS 0.029924f
C10062 DVSS.n715 VSS 0.045559f
C10063 DVSS.n716 VSS 0.05737f
C10064 DVSS.n718 VSS 0.045559f
C10065 DVSS.n719 VSS 0.022779f
C10066 DVSS.n721 VSS 0.041971f
C10067 DVSS.n722 VSS 0.026154f
C10068 DVSS.n723 VSS 0.176874f
C10069 DVSS.n724 VSS 0.176874f
C10070 DVSS.n725 VSS 0.176874f
C10071 DVSS.n726 VSS 0.154453f
C10072 DVSS.n727 VSS 0.022779f
C10073 DVSS.n728 VSS 0.022779f
C10074 DVSS.n729 VSS 0.022779f
C10075 DVSS.n730 VSS 0.022779f
C10076 DVSS.n731 VSS 0.022779f
C10077 DVSS.n732 VSS 0.022779f
C10078 DVSS.n733 VSS 0.022779f
C10079 DVSS.n734 VSS 0.022779f
C10080 DVSS.n735 VSS 0.022779f
C10081 DVSS.n736 VSS 0.022779f
C10082 DVSS.n737 VSS 0.022779f
C10083 DVSS.n738 VSS 0.282749f
C10084 DVSS.n739 VSS 0.022779f
C10085 DVSS.n740 VSS 0.022779f
C10086 DVSS.n741 VSS 0.022779f
C10087 DVSS.n742 VSS 0.022779f
C10088 DVSS.n743 VSS 0.022779f
C10089 DVSS.n744 VSS 0.022779f
C10090 DVSS.n745 VSS 0.022779f
C10091 DVSS.n746 VSS 0.022779f
C10092 DVSS.n747 VSS 0.022779f
C10093 DVSS.n748 VSS 0.022779f
C10094 DVSS.n749 VSS 0.023834f
C10095 DVSS.n750 VSS 16.32f
C10096 DVSS.n751 VSS -1.4011f
C10097 DVSS.n752 VSS 0.028052f
C10098 DVSS.n753 VSS 0.041971f
C10099 DVSS.n754 VSS 0.022779f
C10100 DVSS.n755 VSS 0.176874f
C10101 DVSS.n756 VSS 0.176874f
C10102 DVSS.n757 VSS 0.176874f
C10103 DVSS.n758 VSS 0.315134f
C10104 DVSS.n759 VSS 0.022779f
C10105 DVSS.n760 VSS 0.022779f
C10106 DVSS.n761 VSS 0.022779f
C10107 DVSS.n762 VSS 0.022779f
C10108 DVSS.n763 VSS 0.022779f
C10109 DVSS.n764 VSS 0.022779f
C10110 DVSS.n765 VSS 0.022779f
C10111 DVSS.n766 VSS 0.022779f
C10112 DVSS.n767 VSS 0.022779f
C10113 DVSS.n768 VSS 0.022779f
C10114 DVSS.n769 VSS 0.022779f
C10115 DVSS.n770 VSS 0.154453f
C10116 DVSS.n771 VSS 0.022779f
C10117 DVSS.n772 VSS 0.022779f
C10118 DVSS.n773 VSS 0.022779f
C10119 DVSS.n774 VSS 0.022779f
C10120 DVSS.n775 VSS 0.022779f
C10121 DVSS.n776 VSS 0.022779f
C10122 DVSS.n777 VSS 0.022779f
C10123 DVSS.n778 VSS 0.022779f
C10124 DVSS.n779 VSS 0.022779f
C10125 DVSS.n780 VSS 0.022779f
C10126 DVSS.n781 VSS 0.078891f
C10127 DVSS.n784 VSS 0.049144f
C10128 DVSS.n785 VSS 0.022779f
C10129 DVSS.n786 VSS 0.031005f
C10130 DVSS.n789 VSS 0.041973f
C10131 DVSS.n791 VSS 0.026154f
C10132 DVSS.n793 VSS 0.048189f
C10133 DVSS.n795 VSS 0.041973f
C10134 DVSS.n796 VSS 0.031427f
C10135 DVSS.n799 VSS 0.041973f
C10136 DVSS.n801 VSS 0.026154f
C10137 DVSS.n803 VSS 0.048189f
C10138 DVSS.n805 VSS 0.041973f
C10139 DVSS.n807 VSS 0.176874f
C10140 DVSS.n808 VSS 0.176874f
C10141 DVSS.n809 VSS 0.154453f
C10142 DVSS.n810 VSS 0.282749f
C10143 DVSS.n811 VSS 0.052308f
C10144 DVSS.n822 VSS 0.099554f
C10145 DVSS.n824 VSS 0.154453f
C10146 DVSS.n825 VSS 0.353747f
C10147 DVSS.n826 VSS 0.353747f
C10148 DVSS.n827 VSS 0.353747f
C10149 DVSS.n828 VSS 0.353747f
C10150 DVSS.n829 VSS 0.353747f
C10151 DVSS.n830 VSS 0.226697f
C10152 DVSS.n831 VSS 0.353747f
C10153 DVSS.n832 VSS 0.353747f
C10154 DVSS.n833 VSS 0.353747f
C10155 DVSS.n834 VSS 0.353747f
C10156 DVSS.n835 VSS 0.176874f
C10157 DVSS.n836 VSS 0.353747f
C10158 DVSS.n837 VSS 0.353747f
C10159 DVSS.n838 VSS 0.353747f
C10160 DVSS.n839 VSS 0.176874f
C10161 DVSS.n841 VSS 0.052308f
C10162 DVSS.n842 VSS 0.052308f
C10163 DVSS.n843 VSS 0.052308f
C10164 DVSS.n844 VSS 0.052308f
C10165 DVSS.n845 VSS 0.052308f
C10166 DVSS.n846 VSS 0.052308f
C10167 DVSS.n847 VSS 0.052308f
C10168 DVSS.n848 VSS 0.052308f
C10169 DVSS.n849 VSS 0.052308f
C10170 DVSS.n850 VSS 0.052308f
C10171 DVSS.n851 VSS 0.052308f
C10172 DVSS.n852 VSS 0.099554f
C10173 DVSS.n853 VSS 0.154453f
C10174 DVSS.n856 VSS 0.052308f
C10175 DVSS.n859 VSS 0.052308f
C10176 DVSS.n862 VSS 0.052308f
C10177 DVSS.n865 VSS 0.052308f
C10178 DVSS.n868 VSS 0.052308f
C10179 DVSS.n871 VSS 0.052308f
C10180 DVSS.n874 VSS 0.052308f
C10181 DVSS.n877 VSS 0.052308f
C10182 DVSS.n880 VSS 0.052308f
C10183 DVSS.n883 VSS 0.052308f
C10184 DVSS.n886 VSS 0.353747f
C10185 DVSS.n887 VSS 0.353747f
C10186 DVSS.n888 VSS 0.353747f
C10187 DVSS.n889 VSS 0.353747f
C10188 DVSS.n890 VSS 0.353747f
C10189 DVSS.n891 VSS 0.353747f
C10190 DVSS.n892 VSS 0.353747f
C10191 DVSS.n893 VSS 0.353747f
C10192 DVSS.n894 VSS 0.353747f
C10193 DVSS.n895 VSS 0.353747f
C10194 DVSS.n896 VSS 0.353747f
C10195 DVSS.n897 VSS 0.353747f
C10196 DVSS.n898 VSS 0.176874f
C10197 DVSS.n899 VSS 0.353747f
C10198 DVSS.n900 VSS 0.353747f
C10199 DVSS.n901 VSS 0.353747f
C10200 DVSS.n902 VSS 0.176874f
C10201 DVSS.n904 VSS 0.052308f
C10202 DVSS.n905 VSS 0.052308f
C10203 DVSS.n906 VSS 0.052308f
C10204 DVSS.n907 VSS 0.052308f
C10205 DVSS.n908 VSS 0.052308f
C10206 DVSS.n909 VSS 0.052308f
C10207 DVSS.n910 VSS 0.052308f
C10208 DVSS.n911 VSS 0.052308f
C10209 DVSS.n912 VSS 0.052308f
C10210 DVSS.n913 VSS 0.052308f
C10211 DVSS.n914 VSS 0.052308f
C10212 DVSS.n915 VSS 0.099554f
C10213 DVSS.n916 VSS 0.154453f
C10214 DVSS.n919 VSS 0.052308f
C10215 DVSS.n922 VSS 0.052308f
C10216 DVSS.n925 VSS 0.052308f
C10217 DVSS.n928 VSS 0.052308f
C10218 DVSS.n931 VSS 0.052308f
C10219 DVSS.n934 VSS 0.052308f
C10220 DVSS.n937 VSS 0.052308f
C10221 DVSS.n940 VSS 0.052308f
C10222 DVSS.n943 VSS 0.052308f
C10223 DVSS.n946 VSS 0.052308f
C10224 DVSS.n949 VSS 0.425991f
C10225 DVSS.n950 VSS 0.425991f
C10226 DVSS.n951 VSS 0.675109f
C10227 DVSS.n952 VSS 0.353747f
C10228 DVSS.n953 VSS 0.353747f
C10229 DVSS.n954 VSS 0.353747f
C10230 DVSS.n955 VSS 0.353747f
C10231 DVSS.n956 VSS 0.353747f
C10232 DVSS.n957 VSS 0.154453f
C10233 DVSS.n958 VSS 0.353747f
C10234 DVSS.n959 VSS 0.353747f
C10235 DVSS.n960 VSS 0.282749f
C10236 DVSS.n961 VSS 0.353747f
C10237 DVSS.n962 VSS 1.31155f
C10238 DVSS.n963 VSS 0.353747f
C10239 DVSS.n964 VSS 0.176874f
C10240 DVSS.n977 VSS 0.176874f
C10241 DVSS.n978 VSS 0.176874f
C10242 DVSS.n979 VSS 0.670635f
C10243 DVSS.n980 VSS 0.052308f
C10244 DVSS.n981 VSS 0.052308f
C10245 DVSS.n982 VSS 0.052308f
C10246 DVSS.n983 VSS 0.052308f
C10247 DVSS.n984 VSS 0.052308f
C10248 DVSS.n985 VSS 0.052308f
C10249 DVSS.n986 VSS 0.052308f
C10250 DVSS.n987 VSS 0.052308f
C10251 DVSS.n988 VSS 0.052308f
C10252 DVSS.n989 VSS 0.052308f
C10253 DVSS.n990 VSS 0.052308f
C10254 DVSS.n991 VSS 0.099554f
C10255 DVSS.n992 VSS 0.154453f
C10256 DVSS.n994 VSS 0.052308f
C10257 DVSS.n996 VSS 0.052308f
C10258 DVSS.n998 VSS 0.052308f
C10259 DVSS.n1000 VSS 0.052308f
C10260 DVSS.n1002 VSS 0.052308f
C10261 DVSS.n1004 VSS 0.052308f
C10262 DVSS.n1006 VSS 0.052308f
C10263 DVSS.n1008 VSS 0.052308f
C10264 DVSS.n1010 VSS 0.052308f
C10265 DVSS.n1012 VSS 0.052308f
C10266 DVSS.n1013 VSS 0.353747f
C10267 DVSS.n1014 VSS 0.154453f
C10268 DVSS.n1015 VSS 0.353747f
C10269 DVSS.n1016 VSS 0.353747f
C10270 DVSS.n1017 VSS 0.282749f
C10271 DVSS.n1018 VSS 0.353747f
C10272 DVSS.n1019 VSS 0.353747f
C10273 DVSS.n1020 VSS 0.353747f
C10274 DVSS.n1021 VSS 0.353747f
C10275 DVSS.n1022 VSS 0.353747f
C10276 DVSS.n1023 VSS 0.154453f
C10277 DVSS.n1024 VSS 0.154453f
C10278 DVSS.n1025 VSS 0.353747f
C10279 DVSS.n1026 VSS 0.353747f
C10280 DVSS.n1027 VSS 0.282749f
C10281 DVSS.n1028 VSS 0.353747f
C10282 DVSS.n1029 VSS 0.353747f
C10283 DVSS.n1030 VSS 0.236662f
C10284 DVSS.n1031 VSS 0.293959f
C10285 DVSS.n1032 VSS 0.236662f
C10286 DVSS.n1033 VSS 0.255346f
C10287 DVSS.n1034 VSS 0.353747f
C10288 DVSS.n1035 VSS 0.425991f
C10289 DVSS.n1036 VSS 0.353747f
C10290 DVSS.n1037 VSS 0.154453f
C10291 DVSS.n1038 VSS 0.154453f
C10292 DVSS.n1039 VSS 0.282749f
C10293 DVSS.n1040 VSS 0.353747f
C10294 DVSS.n1041 VSS 0.353747f
C10295 DVSS.n1042 VSS 0.353747f
C10296 DVSS.n1043 VSS 0.353747f
C10297 DVSS.n1044 VSS 0.353747f
C10298 DVSS.n1045 VSS 0.353747f
C10299 DVSS.n1046 VSS 0.353747f
C10300 DVSS.n1047 VSS 0.353747f
C10301 DVSS.n1048 VSS 0.353747f
C10302 DVSS.n1049 VSS 0.353747f
C10303 DVSS.n1050 VSS 0.353747f
C10304 DVSS.n1051 VSS 0.353747f
C10305 DVSS.n1052 VSS 0.353747f
C10306 DVSS.n1053 VSS 0.353747f
C10307 DVSS.n1054 VSS 0.353747f
C10308 DVSS.n1055 VSS 0.353747f
C10309 DVSS.n1056 VSS 0.353747f
C10310 DVSS.n1057 VSS 0.315134f
C10311 DVSS.n1058 VSS 0.353747f
C10312 DVSS.n1059 VSS 0.353747f
C10313 DVSS.n1060 VSS 0.154453f
C10314 DVSS.n1061 VSS 0.154453f
C10315 DVSS.n1066 VSS 0.051254f
C10316 DVSS.n1071 VSS 0.052308f
C10317 DVSS.n1072 VSS 0.022779f
C10318 DVSS.n1073 VSS 0.249729f
C10319 DVSS.n1074 VSS 0.026998f
C10320 DVSS.n1075 VSS 0.03206f
C10321 DVSS.n1076 VSS 0.026154f
C10322 DVSS.n1078 VSS 0.176874f
C10323 DVSS.n1080 VSS 0.009955f
C10324 DVSS.n1081 VSS 1.18511f
C10325 DVSS.n1082 VSS 0.021932f
C10326 DVSS.n1083 VSS 0.021932f
C10327 DVSS.n1084 VSS 0.009955f
C10328 DVSS.n1085 VSS 0.009955f
C10329 DVSS.n1086 VSS 0.009955f
C10330 DVSS.n1087 VSS 0.009955f
C10331 DVSS.n1088 VSS 0.186081f
C10332 DVSS.n1089 VSS 1.02218f
C10333 DVSS.t37 VSS 25.4676f
C10334 DVSS.n1090 VSS 0.101916f
C10335 DVSS.n1091 VSS 1.00578f
C10336 DVSS.n1092 VSS 0.101916f
C10337 DVSS.n1093 VSS 1.18511f
C10338 DVSS.n1094 VSS 1.02218f
C10339 DVSS.n1095 VSS 0.102784f
C10340 DVSS.n1096 VSS 0.094754f
C10341 DVSS.n1098 VSS 0.026154f
C10342 DVSS.n1100 VSS 0.033721f
C10343 DVSS.n1101 VSS 0.029107f
C10344 DVSS.n1103 VSS 0.033721f
C10345 DVSS.n1104 VSS 0.30411f
C10346 DVSS.n1105 VSS 0.082541f
C10347 DVSS.n1106 VSS 0.082541f
C10348 DVSS.n1107 VSS 0.082541f
C10349 DVSS.n1108 VSS 0.134274f
C10350 DVSS.n1109 VSS 0.052308f
C10351 DVSS.n1111 VSS 0.052308f
C10352 DVSS.n1112 VSS 0.052308f
C10353 DVSS.n1113 VSS 0.052308f
C10354 DVSS.n1114 VSS 0.072078f
C10355 DVSS.n1116 VSS 0.163463f
C10356 DVSS.n1119 VSS 0.052308f
C10357 DVSS.n1121 VSS 0.029951f
C10358 DVSS.n1124 VSS 0.052308f
C10359 DVSS.n1128 VSS 0.033721f
C10360 DVSS.n1129 VSS 0.033721f
C10361 DVSS.n1131 VSS 0.033721f
C10362 DVSS.n1134 VSS 0.045559f
C10363 DVSS.n1135 VSS 0.169158f
C10364 DVSS.n1138 VSS 0.033721f
C10365 DVSS.n1139 VSS 0.033721f
C10366 DVSS.n1142 VSS 0.038205f
C10367 DVSS.n1143 VSS 0.141853f
C10368 DVSS.n1145 VSS 0.029505f
C10369 DVSS.n1146 VSS 0.101916f
C10370 DVSS.n1147 VSS 1.00578f
C10371 DVSS.n1148 VSS 1.02218f
C10372 DVSS.n1149 VSS 0.094754f
C10373 DVSS.n1150 VSS 0.663966f
C10374 DVSS.n1151 VSS 0.102784f
C10375 DVSS.n1152 VSS 0.023201f
C10376 DVSS.n1155 VSS 0.033721f
C10377 DVSS.n1156 VSS 0.029107f
C10378 DVSS.n1158 VSS 0.30411f
C10379 DVSS.n1159 VSS 0.033721f
C10380 DVSS.n1160 VSS 0.029951f
C10381 DVSS.n1161 VSS 0.082541f
C10382 DVSS.n1162 VSS 0.082541f
C10383 DVSS.n1163 VSS 0.082541f
C10384 DVSS.n1164 VSS 0.147063f
C10385 DVSS.n1165 VSS 0.052308f
C10386 DVSS.n1167 VSS 0.052308f
C10387 DVSS.n1169 VSS 0.052308f
C10388 DVSS.n1170 VSS 0.052308f
C10389 DVSS.n1171 VSS 0.072078f
C10390 DVSS.n1173 VSS 0.163463f
C10391 DVSS.n1176 VSS 0.052308f
C10392 DVSS.n1179 VSS 0.052308f
C10393 DVSS.n1183 VSS 0.033721f
C10394 DVSS.n1184 VSS 0.033721f
C10395 DVSS.n1186 VSS 0.033721f
C10396 DVSS.n1188 VSS 0.182276f
C10397 DVSS.n1190 VSS 0.176874f
C10398 DVSS.n1191 VSS 0.176874f
C10399 DVSS.n1192 VSS 0.052308f
C10400 DVSS.n1193 VSS 0.052308f
C10401 DVSS.n1194 VSS 0.052308f
C10402 DVSS.n1195 VSS 0.051254f
C10403 DVSS.n1196 VSS 0.030583f
C10404 DVSS.n1197 VSS 0.052308f
C10405 DVSS.n1198 VSS 0.052308f
C10406 DVSS.n1199 VSS 0.052308f
C10407 DVSS.n1200 VSS 0.052308f
C10408 DVSS.n1201 VSS 0.022779f
C10409 DVSS.n1202 VSS 0.154453f
C10410 DVSS.n1203 VSS 0.026998f
C10411 DVSS.n1205 VSS 0.03206f
C10412 DVSS.n1207 VSS 0.052308f
C10413 DVSS.n1209 VSS 0.052308f
C10414 DVSS.n1211 VSS 0.052308f
C10415 DVSS.n1213 VSS 0.052308f
C10416 DVSS.n1214 VSS 0.026154f
C10417 DVSS.n1215 VSS 0.179554f
C10418 DVSS.n1216 VSS 0.179554f
C10419 DVSS.n1217 VSS 0.009955f
C10420 DVSS.n1218 VSS 0.019909f
C10421 DVSS.n1219 VSS 0.019909f
C10422 DVSS.n1220 VSS 0.02531f
C10423 DVSS.n1222 VSS 0.033721f
C10424 DVSS.n1225 VSS 0.033721f
C10425 DVSS.n1227 VSS 0.02531f
C10426 DVSS.n1229 VSS 0.033721f
C10427 DVSS.n1232 VSS 0.033721f
C10428 DVSS.n1234 VSS 0.021225f
C10429 DVSS.n1236 VSS 0.033721f
C10430 DVSS.n1237 VSS 0.033721f
C10431 DVSS.n1238 VSS 0.021225f
C10432 DVSS.n1240 VSS 0.033721f
C10433 DVSS.n1241 VSS 0.033721f
C10434 DVSS.n1242 VSS 0.02531f
C10435 DVSS.n1244 VSS 0.033721f
C10436 DVSS.n1247 VSS 0.033721f
C10437 DVSS.n1249 VSS 0.02531f
C10438 DVSS.n1251 VSS 0.033721f
C10439 DVSS.n1254 VSS 0.033721f
C10440 DVSS.n1256 VSS 0.07353f
C10441 DVSS.n1257 VSS 0.023623f
C10442 DVSS.n1258 VSS 0.033721f
C10443 DVSS.n1259 VSS 0.026154f
C10444 DVSS.n1260 VSS 0.30411f
C10445 DVSS.n1261 VSS 0.30411f
C10446 DVSS.n1262 VSS 0.023623f
C10447 DVSS.n1263 VSS 0.033721f
C10448 DVSS.n1264 VSS 0.026154f
C10449 DVSS.n1265 VSS 0.306139f
C10450 DVSS.n1267 VSS 0.01981f
C10451 DVSS.n1268 VSS 0.306139f
C10452 DVSS.n1270 VSS 0.021932f
C10453 DVSS.n1271 VSS 0.029505f
C10454 DVSS.n1272 VSS 1.02218f
C10455 DVSS.n1273 VSS 1.75989f
C10456 DVSS.n1274 VSS 0.02529f
C10457 DVSS.n1276 VSS 0.01981f
C10458 DVSS.n1277 VSS 0.029505f
C10459 DVSS.n1279 VSS 0.021932f
C10460 DVSS.n1280 VSS 0.306139f
C10461 DVSS.n1281 VSS 0.306139f
C10462 DVSS.n1282 VSS 0.023623f
C10463 DVSS.n1283 VSS 0.033721f
C10464 DVSS.n1284 VSS 0.026154f
C10465 DVSS.n1285 VSS 0.30411f
C10466 DVSS.n1286 VSS 0.30411f
C10467 DVSS.n1287 VSS 0.023623f
C10468 DVSS.n1288 VSS 0.033721f
C10469 DVSS.n1289 VSS 0.026154f
C10470 DVSS.n1290 VSS 0.07353f
C10471 DVSS.n1291 VSS 0.094754f
C10472 DVSS.n1292 VSS 0.186081f
C10473 DVSS.n1293 VSS 0.136683f
C10474 DVSS.n1294 VSS 0.009955f
C10475 DVSS.n1295 VSS 0.102784f
C10476 DVSS.n1296 VSS 0.026154f
C10477 DVSS.n1297 VSS 0.022779f
C10478 DVSS.n1299 VSS 0.052308f
C10479 DVSS.n1301 VSS 0.052308f
C10480 DVSS.n1303 VSS 0.052308f
C10481 DVSS.n1311 VSS 0.176874f
C10482 DVSS.n1314 VSS 0.052308f
C10483 DVSS.n1315 VSS 0.176874f
C10484 DVSS.n1316 VSS 0.249729f
C10485 DVSS.n1317 VSS 0.246354f
C10486 DVSS.n1318 VSS 0.07353f
C10487 DVSS.n1319 VSS 0.045559f
C10488 DVSS.n1320 VSS 0.033721f
C10489 DVSS.n1323 VSS 0.033721f
C10490 DVSS.n1324 VSS 0.306139f
C10491 DVSS.n1326 VSS 0.082541f
C10492 DVSS.n1327 VSS 0.082541f
C10493 DVSS.n1328 VSS 0.147063f
C10494 DVSS.n1329 VSS 0.052308f
C10495 DVSS.n1330 VSS 0.052308f
C10496 DVSS.n1331 VSS 0.022779f
C10497 DVSS.n1332 VSS 0.052308f
C10498 DVSS.n1333 VSS 0.052308f
C10499 DVSS.n1334 VSS 0.072078f
C10500 DVSS.n1335 VSS 0.163463f
C10501 DVSS.n1337 VSS 0.052308f
C10502 DVSS.n1339 VSS 0.029951f
C10503 DVSS.n1341 VSS 0.029107f
C10504 DVSS.n1344 VSS 0.165082f
C10505 DVSS.n1345 VSS 0.072078f
C10506 DVSS.n1346 VSS 0.165082f
C10507 DVSS.n1347 VSS 0.165082f
C10508 DVSS.n1348 VSS 0.165082f
C10509 DVSS.n1349 VSS 0.165082f
C10510 DVSS.n1350 VSS 0.165082f
C10511 DVSS.n1351 VSS 0.165082f
C10512 DVSS.n1352 VSS 0.165082f
C10513 DVSS.n1353 VSS 0.165082f
C10514 DVSS.n1354 VSS 0.165082f
C10515 DVSS.n1355 VSS 0.165082f
C10516 DVSS.n1356 VSS 0.165082f
C10517 DVSS.n1357 VSS 0.165082f
C10518 DVSS.n1358 VSS 0.165082f
C10519 DVSS.n1359 VSS 0.165082f
C10520 DVSS.n1360 VSS 0.165082f
C10521 DVSS.n1361 VSS 0.165082f
C10522 DVSS.n1362 VSS 0.043865f
C10523 DVSS.n1363 VSS 0.043865f
C10524 DVSS.n1364 VSS 0.019102f
C10525 DVSS.n1365 VSS 0.043865f
C10526 DVSS.n1366 VSS 0.043865f
C10527 DVSS.n1367 VSS 0.072078f
C10528 DVSS.n1368 VSS 0.137077f
C10529 DVSS.n1369 VSS 0.043865f
C10530 DVSS.n1370 VSS 0.025116f
C10531 DVSS.n1371 VSS 0.024409f
C10532 DVSS.n1372 VSS 0.043865f
C10533 DVSS.n1377 VSS 0.082541f
C10534 DVSS.n1379 VSS 0.306139f
C10535 DVSS.n1380 VSS 0.033721f
C10536 DVSS.n1382 VSS 0.206588f
C10537 DVSS.n1383 VSS 0.038205f
C10538 DVSS.n1385 VSS 0.033721f
C10539 DVSS.n1387 VSS 0.139023f
C10540 DVSS.n1388 VSS 0.072078f
C10541 DVSS.n1392 VSS 0.111605f
C10542 DVSS.n1393 VSS 0.165082f
C10543 DVSS.n1394 VSS 0.165082f
C10544 DVSS.n1395 VSS 0.165082f
C10545 DVSS.n1396 VSS 0.165082f
C10546 DVSS.n1397 VSS 0.165082f
C10547 DVSS.n1398 VSS 0.082541f
C10548 DVSS.n1401 VSS 0.019102f
C10549 DVSS.n1404 VSS 0.072078f
C10550 DVSS.n1405 VSS 0.021932f
C10551 DVSS.n1406 VSS 0.043865f
C10552 DVSS.n1408 VSS 0.043865f
C10553 DVSS.n1409 VSS 0.043865f
C10554 DVSS.n1411 VSS 0.043865f
C10555 DVSS.n1412 VSS 0.043865f
C10556 DVSS.n1414 VSS 0.156944f
C10557 DVSS.n1415 VSS 0.137077f
C10558 DVSS.n1417 VSS 0.023201f
C10559 DVSS.n1421 VSS 0.033721f
C10560 DVSS.n1422 VSS 0.029107f
C10561 DVSS.n1423 VSS 0.033721f
C10562 DVSS.n1424 VSS 0.029951f
C10563 DVSS.n1425 VSS 0.082541f
C10564 DVSS.n1426 VSS 0.082541f
C10565 DVSS.n1427 VSS 0.082541f
C10566 DVSS.n1428 VSS 0.134274f
C10567 DVSS.n1430 VSS 0.052308f
C10568 DVSS.n1432 VSS 0.052308f
C10569 DVSS.n1434 VSS 0.052308f
C10570 DVSS.n1435 VSS 0.052308f
C10571 DVSS.n1436 VSS 0.072078f
C10572 DVSS.n1438 VSS 0.179554f
C10573 DVSS.n1439 VSS 0.009955f
C10574 DVSS.n1440 VSS 0.180752f
C10575 DVSS.n1441 VSS 0.019909f
C10576 DVSS.n1442 VSS 0.019909f
C10577 DVSS.n1443 VSS 0.184214f
C10578 DVSS.n1444 VSS 0.180752f
C10579 DVSS.n1446 VSS 0.306139f
C10580 DVSS.n1448 VSS 0.033721f
C10581 DVSS.n1449 VSS 0.161143f
C10582 DVSS.n1450 VSS 0.045718f
C10583 DVSS.n1451 VSS 0.797916f
C10584 DVSS.n1452 VSS 0.922342f
C10585 DVSS.t3 VSS 13.811f
C10586 DVSS.n1453 VSS 0.04802f
C10587 DVSS.n1454 VSS 0.952584f
C10588 DVSS.n1455 VSS 0.04802f
C10589 DVSS.n1456 VSS 0.922342f
C10590 DVSS.n1457 VSS 0.797916f
C10591 DVSS.n1458 VSS 0.184214f
C10592 DVSS.n1459 VSS 0.045718f
C10593 DVSS.n1460 VSS 0.033721f
C10594 DVSS.n1461 VSS 0.157979f
C10595 DVSS.n1463 VSS 0.045559f
C10596 DVSS.n1465 VSS 0.161143f
C10597 DVSS.n1466 VSS 0.033721f
C10598 DVSS.n1467 VSS 0.132478f
C10599 DVSS.n1469 VSS 0.038205f
C10600 DVSS.n1471 VSS 0.135131f
C10601 DVSS.n1472 VSS 0.029505f
C10602 DVSS.n1473 VSS 0.507231f
C10603 DVSS.n1474 VSS 0.77032f
C10604 DVSS.n1475 VSS 0.045718f
C10605 DVSS.n1476 VSS 0.952584f
C10606 DVSS.n1477 VSS 0.507231f
C10607 DVSS.n1478 VSS 0.797916f
C10608 DVSS.n1479 VSS 0.328284f
C10609 DVSS.n1480 VSS 0.211948f
C10610 DVSS.n1482 VSS 0.045559f
C10611 DVSS.n1484 VSS 0.157979f
C10612 DVSS.n1486 VSS 0.033721f
C10613 DVSS.n1488 VSS 0.033721f
C10614 DVSS.n1489 VSS 0.033721f
C10615 DVSS.n1490 VSS 0.161143f
C10616 DVSS.n1492 VSS 0.132478f
C10617 DVSS.n1494 VSS 0.033721f
C10618 DVSS.n1496 VSS 0.033721f
C10619 DVSS.n1497 VSS 0.135131f
C10620 DVSS.n1499 VSS 0.132478f
C10621 DVSS.n1501 VSS 0.033721f
C10622 DVSS.n1503 VSS 0.033721f
C10623 DVSS.n1506 VSS 0.033721f
C10624 DVSS.n1507 VSS 0.135131f
C10625 DVSS.n1509 VSS 0.038205f
C10626 DVSS.n1511 VSS 0.033721f
C10627 DVSS.n1513 VSS 0.267267f
C10628 DVSS.n1515 VSS 0.033721f
C10629 DVSS.n1516 VSS 0.157979f
C10630 DVSS.n1518 VSS 0.135131f
C10631 DVSS.n1521 VSS 0.019909f
C10632 DVSS.n1522 VSS 0.019909f
C10633 DVSS.n1523 VSS 0.249392f
C10634 DVSS.n1526 VSS 0.019909f
C10635 DVSS.n1527 VSS 0.019909f
C10636 DVSS.n1528 VSS 0.249392f
C10637 DVSS.n1529 VSS 0.009955f
C10638 DVSS.n1533 VSS 0.032106f
C10639 DVSS.n1534 VSS 0.032106f
C10640 DVSS.n1536 VSS 0.032106f
C10641 DVSS.n1538 VSS 0.74982f
C10642 DVSS.t22 VSS 0.394423f
C10643 DVSS.n1539 VSS 0.635269f
C10644 DVSS.n1541 VSS 0.045559f
C10645 DVSS.n1544 VSS 0.009955f
C10646 DVSS.n1545 VSS 0.179554f
C10647 DVSS.n1546 VSS 0.160088f
C10648 DVSS.n1547 VSS 0.009955f
C10649 DVSS.n1548 VSS 0.019909f
C10650 DVSS.n1549 VSS 0.019909f
C10651 DVSS.n1550 VSS 1.42561f
C10652 DVSS.n1552 VSS 0.032106f
C10653 DVSS.n1553 VSS 0.753194f
C10654 DVSS.n1555 VSS 0.045559f
C10655 DVSS.n1557 VSS 1.58907f
C10656 DVSS.n1559 VSS 0.032106f
C10657 DVSS.n1560 VSS 0.753194f
C10658 DVSS.n1563 VSS 0.363609f
C10659 DVSS.n1564 VSS 0.082541f
C10660 DVSS.n1565 VSS 0.068009f
C10661 DVSS.n1566 VSS 0.052308f
C10662 DVSS.n1567 VSS 0.052308f
C10663 DVSS.n1568 VSS 0.052308f
C10664 DVSS.n1569 VSS 0.052308f
C10665 DVSS.n1570 VSS 0.052308f
C10666 DVSS.n1571 VSS 0.072078f
C10667 DVSS.n1573 VSS 0.052308f
C10668 DVSS.n1575 VSS 0.052308f
C10669 DVSS.n1577 VSS 0.052308f
C10670 DVSS.n1579 VSS 0.052308f
C10671 DVSS.n1585 VSS 0.165082f
C10672 DVSS.n1586 VSS 0.072078f
C10673 DVSS.n1587 VSS 0.165082f
C10674 DVSS.n1588 VSS 0.165082f
C10675 DVSS.n1589 VSS 0.165082f
C10676 DVSS.n1590 VSS 0.144737f
C10677 DVSS.n1591 VSS 0.165082f
C10678 DVSS.n1592 VSS 0.165082f
C10679 DVSS.n1593 VSS 0.165082f
C10680 DVSS.n1594 VSS 0.082541f
C10681 DVSS.n1599 VSS 0.438291f
C10682 DVSS.n1601 VSS 0.134274f
C10683 DVSS.n1602 VSS 0.052308f
C10684 DVSS.n1603 VSS 0.052308f
C10685 DVSS.n1604 VSS 0.052308f
C10686 DVSS.n1605 VSS 0.052308f
C10687 DVSS.n1606 VSS 0.165082f
C10688 DVSS.n1607 VSS 0.165082f
C10689 DVSS.n1608 VSS 0.165082f
C10690 DVSS.n1609 VSS 0.144737f
C10691 DVSS.n1610 VSS 0.165082f
C10692 DVSS.n1611 VSS 0.165082f
C10693 DVSS.n1612 VSS 0.165082f
C10694 DVSS.n1613 VSS 0.165082f
C10695 DVSS.n1614 VSS 0.165082f
C10696 DVSS.n1615 VSS 0.165082f
C10697 DVSS.n1616 VSS 0.165082f
C10698 DVSS.n1617 VSS 0.165082f
C10699 DVSS.n1618 VSS 0.165082f
C10700 DVSS.n1619 VSS 0.165082f
C10701 DVSS.n1620 VSS 0.165082f
C10702 DVSS.n1621 VSS 0.165082f
C10703 DVSS.n1622 VSS 0.165082f
C10704 DVSS.n1623 VSS 0.144737f
C10705 DVSS.n1624 VSS 0.165082f
C10706 DVSS.n1625 VSS 0.165082f
C10707 DVSS.n1626 VSS 0.165082f
C10708 DVSS.n1627 VSS 0.165082f
C10709 DVSS.n1628 VSS 0.165082f
C10710 DVSS.n1629 VSS 0.165082f
C10711 DVSS.n1630 VSS 0.165082f
C10712 DVSS.n1631 VSS 0.165082f
C10713 DVSS.n1632 VSS 0.165082f
C10714 DVSS.n1633 VSS 0.165082f
C10715 DVSS.n1634 VSS 0.165082f
C10716 DVSS.n1635 VSS 0.165082f
C10717 DVSS.n1636 VSS 0.165082f
C10718 DVSS.n1637 VSS 0.165082f
C10719 DVSS.n1638 VSS 0.165082f
C10720 DVSS.n1639 VSS 0.165082f
C10721 DVSS.n1640 VSS 0.165082f
C10722 DVSS.n1641 VSS 0.165082f
C10723 DVSS.n1642 VSS 0.165082f
C10724 DVSS.n1643 VSS 0.165082f
C10725 DVSS.n1644 VSS 0.165082f
C10726 DVSS.n1645 VSS 0.165082f
C10727 DVSS.n1646 VSS 0.165082f
C10728 DVSS.n1647 VSS 0.165082f
C10729 DVSS.n1648 VSS 0.165082f
C10730 DVSS.n1649 VSS 0.165082f
C10731 DVSS.n1650 VSS 0.165082f
C10732 DVSS.n1651 VSS 0.165082f
C10733 DVSS.n1652 VSS 0.165082f
C10734 DVSS.n1653 VSS 0.165082f
C10735 DVSS.n1654 VSS 0.165082f
C10736 DVSS.n1655 VSS 0.165082f
C10737 DVSS.n1656 VSS 0.165082f
C10738 DVSS.n1657 VSS 0.165082f
C10739 DVSS.n1658 VSS 0.165082f
C10740 DVSS.n1659 VSS 0.165082f
C10741 DVSS.n1660 VSS 0.165082f
C10742 DVSS.n1661 VSS 0.165082f
C10743 DVSS.n1662 VSS 0.165082f
C10744 DVSS.n1663 VSS 0.165082f
C10745 DVSS.n1664 VSS 0.165082f
C10746 DVSS.n1665 VSS 0.072078f
C10747 DVSS.n1666 VSS 0.165082f
C10748 DVSS.n1667 VSS 0.072078f
C10749 DVSS.n1668 VSS 0.165082f
C10750 DVSS.n1669 VSS 0.165082f
C10751 DVSS.n1670 VSS 0.165082f
C10752 DVSS.n1671 VSS 0.165082f
C10753 DVSS.n1672 VSS 0.165082f
C10754 DVSS.n1673 VSS 0.165082f
C10755 DVSS.n1674 VSS 0.165082f
C10756 DVSS.n1675 VSS 0.165082f
C10757 DVSS.n1676 VSS 0.165082f
C10758 DVSS.n1677 VSS 0.165082f
C10759 DVSS.n1678 VSS 0.165082f
C10760 DVSS.n1679 VSS 0.165082f
C10761 DVSS.n1680 VSS 0.165082f
C10762 DVSS.n1681 VSS 0.165082f
C10763 DVSS.n1682 VSS 0.165082f
C10764 DVSS.n1683 VSS 0.165082f
C10765 DVSS.n1684 VSS 0.165082f
C10766 DVSS.n1685 VSS 0.165082f
C10767 DVSS.n1686 VSS 0.165082f
C10768 DVSS.n1687 VSS 0.165082f
C10769 DVSS.n1688 VSS 0.165082f
C10770 DVSS.n1689 VSS 0.165082f
C10771 DVSS.n1690 VSS 0.165082f
C10772 DVSS.n1691 VSS 0.165082f
C10773 DVSS.n1692 VSS 0.165082f
C10774 DVSS.n1693 VSS 0.165082f
C10775 DVSS.n1694 VSS 0.165082f
C10776 DVSS.n1695 VSS 0.165082f
C10777 DVSS.n1696 VSS 0.165082f
C10778 DVSS.n1697 VSS 0.072078f
C10779 DVSS.n1698 VSS 0.165082f
C10780 DVSS.n1699 VSS 0.072078f
C10781 DVSS.n1700 VSS 0.165082f
C10782 DVSS.n1701 VSS 0.165082f
C10783 DVSS.n1702 VSS 0.165082f
C10784 DVSS.n1703 VSS 0.165082f
C10785 DVSS.n1704 VSS 0.165082f
C10786 DVSS.n1705 VSS 0.165082f
C10787 DVSS.n1706 VSS 0.165082f
C10788 DVSS.n1707 VSS 0.165082f
C10789 DVSS.n1708 VSS 0.165082f
C10790 DVSS.n1709 VSS 0.165082f
C10791 DVSS.n1710 VSS 0.165082f
C10792 DVSS.n1711 VSS 0.165082f
C10793 DVSS.n1712 VSS 0.165082f
C10794 DVSS.n1713 VSS 0.072078f
C10795 DVSS.n1714 VSS 0.052308f
C10796 DVSS.n1715 VSS 0.052308f
C10797 DVSS.n1719 VSS 0.072078f
C10798 DVSS.n1720 VSS 0.082541f
C10799 DVSS.n1722 VSS 0.052308f
C10800 DVSS.n1723 VSS 0.052308f
C10801 DVSS.n1724 VSS 0.082541f
C10802 DVSS.n1725 VSS 0.052308f
C10803 DVSS.n1727 VSS 0.082541f
C10804 DVSS.n1728 VSS 0.072078f
C10805 DVSS.n1729 VSS 0.165082f
C10806 DVSS.n1730 VSS 0.165082f
C10807 DVSS.n1731 VSS 0.165082f
C10808 DVSS.n1732 VSS 0.165082f
C10809 DVSS.n1733 VSS 0.165082f
C10810 DVSS.n1734 VSS 0.165082f
C10811 DVSS.n1735 VSS 0.165082f
C10812 DVSS.n1736 VSS 0.165082f
C10813 DVSS.n1737 VSS 0.148806f
C10814 DVSS.n1738 VSS 0.148806f
C10815 DVSS.n1739 VSS 0.098817f
C10816 DVSS.n1740 VSS 0.084866f
C10817 DVSS.n1741 VSS 0.162757f
C10818 DVSS.n1742 VSS 0.319361f
C10819 DVSS.n1743 VSS 0.616179f
C10820 DVSS.n1744 VSS 0.165082f
C10821 DVSS.n1745 VSS 0.072078f
C10822 DVSS.n1746 VSS 0.082541f
C10823 DVSS.n1747 VSS 0.438291f
C10824 DVSS.n1748 VSS 0.082541f
C10825 DVSS.n1749 VSS 1.58907f
C10826 DVSS.n1750 VSS 1.58569f
C10827 DVSS.n1751 VSS 0.756569f
C10828 DVSS.n1752 VSS 0.21755f
C10829 DVSS.n1755 VSS 0.045559f
C10830 DVSS.n1756 VSS 0.058114f
C10831 DVSS.n1757 VSS 0.045559f
C10832 DVSS.n1758 VSS 0.331802f
C10833 DVSS.n1759 VSS 0.045559f
C10834 DVSS.n1762 VSS 0.082541f
C10835 DVSS.n1763 VSS 0.082541f
C10836 DVSS.n1764 VSS 0.068009f
C10837 DVSS.n1765 VSS 0.052308f
C10838 DVSS.n1766 VSS 0.052308f
C10839 DVSS.n1767 VSS 0.052308f
C10840 DVSS.n1768 VSS 0.052308f
C10841 DVSS.n1769 VSS 0.052308f
C10842 DVSS.n1770 VSS 0.072078f
C10843 DVSS.n1772 VSS 0.163885f
C10844 DVSS.n1774 VSS 0.052308f
C10845 DVSS.n1776 VSS 0.052308f
C10846 DVSS.n1778 VSS 0.052308f
C10847 DVSS.n1779 VSS 0.072078f
C10848 DVSS.n1780 VSS 0.165082f
C10849 DVSS.n1781 VSS 0.162757f
C10850 DVSS.n1782 VSS 0.165082f
C10851 DVSS.n1783 VSS 0.165082f
C10852 DVSS.n1784 VSS 0.144737f
C10853 DVSS.n1785 VSS 0.165082f
C10854 DVSS.n1786 VSS 0.165082f
C10855 DVSS.n1787 VSS 0.165082f
C10856 DVSS.n1788 VSS 0.082541f
C10857 DVSS.n1789 VSS 0.157135f
C10858 DVSS.n1794 VSS 0.361727f
C10859 DVSS.n1796 VSS 0.134274f
C10860 DVSS.n1797 VSS 0.052308f
C10861 DVSS.n1798 VSS 0.052308f
C10862 DVSS.n1799 VSS 0.052308f
C10863 DVSS.n1800 VSS 0.052308f
C10864 DVSS.n1801 VSS 0.165082f
C10865 DVSS.n1802 VSS 0.165082f
C10866 DVSS.n1803 VSS 0.165082f
C10867 DVSS.n1804 VSS 0.144737f
C10868 DVSS.n1805 VSS 0.165082f
C10869 DVSS.n1806 VSS 0.165082f
C10870 DVSS.n1807 VSS 0.165082f
C10871 DVSS.n1808 VSS 0.082541f
C10872 DVSS.n1814 VSS 0.157135f
C10873 DVSS.n1816 VSS 0.134274f
C10874 DVSS.n1817 VSS 0.052308f
C10875 DVSS.n1818 VSS 0.052308f
C10876 DVSS.n1819 VSS 0.052308f
C10877 DVSS.n1820 VSS 0.052308f
C10878 DVSS.n1821 VSS 0.052308f
C10879 DVSS.n1822 VSS 0.072078f
C10880 DVSS.n1823 VSS 0.052308f
C10881 DVSS.n1824 VSS 0.052308f
C10882 DVSS.n1825 VSS 0.052308f
C10883 DVSS.n1826 VSS 0.052308f
C10884 DVSS.n1831 VSS 0.072078f
C10885 DVSS.n1832 VSS 0.082541f
C10886 DVSS.n1835 VSS 0.066724f
C10887 DVSS.n1837 VSS 0.052308f
C10888 DVSS.n1840 VSS 0.052308f
C10889 DVSS.n1842 VSS 0.066724f
C10890 DVSS.n1844 VSS 0.052308f
C10891 DVSS.n1846 VSS 0.066724f
C10892 DVSS.n1847 VSS 0.052308f
C10893 DVSS.n1848 VSS 0.222771f
C10894 DVSS.n1849 VSS 0.361727f
C10895 DVSS.n1851 VSS 0.179185f
C10896 DVSS.n1852 VSS 0.052308f
C10897 DVSS.t5 VSS 0.394423f
C10898 DVSS.n1854 VSS 0.635269f
C10899 DVSS.n1855 VSS 0.066724f
C10900 DVSS.n1856 VSS 0.361727f
C10901 DVSS.n1857 VSS 0.052308f
C10902 DVSS.n1859 VSS 0.753194f
C10903 DVSS.n1860 VSS 0.052308f
C10904 DVSS.n1864 VSS 0.066724f
C10905 DVSS.n1866 VSS 0.043865f
C10906 DVSS.n1868 VSS 0.069335f
C10907 DVSS.n1870 VSS -0.427302f
C10908 DVSS.n1871 VSS 0.038205f
C10909 DVSS.n1872 VSS 0.035873f
C10910 DVSS.n1873 VSS 0.038205f
C10911 DVSS.n1875 VSS 0.043865f
C10912 DVSS.n1876 VSS 0.066724f
C10913 DVSS.n1877 VSS 0.043865f
C10914 DVSS.n1879 VSS 0.069335f
C10915 DVSS.n1881 VSS 0.066724f
C10916 DVSS.n1882 VSS 0.361727f
C10917 DVSS.n1883 VSS 0.052308f
C10918 DVSS.n1885 VSS 0.753194f
C10919 DVSS.n1886 VSS 0.052308f
C10920 DVSS.t4 VSS 0.330478f
C10921 DVSS.n1890 VSS 0.635269f
C10922 DVSS.n1891 VSS 0.066724f
C10923 DVSS.n1892 VSS 0.361727f
C10924 DVSS.n1893 VSS 0.052308f
C10925 DVSS.n1895 VSS 0.753194f
C10926 DVSS.n1896 VSS 0.052308f
C10927 DVSS.n1900 VSS 0.066724f
C10928 DVSS.n1901 VSS 0.361727f
C10929 DVSS.n1902 VSS 0.052308f
C10930 DVSS.n1904 VSS 0.753194f
C10931 DVSS.n1905 VSS 0.052308f
C10932 DVSS.t11 VSS 0.394423f
C10933 DVSS.n1909 VSS 0.045559f
C10934 DVSS.n1910 VSS 0.045559f
C10935 DVSS.n1911 VSS 0.045559f
C10936 DVSS.n1914 VSS 0.756569f
C10937 DVSS.n1915 VSS 0.217854f
C10938 DVSS.n1917 VSS 0.082541f
C10939 DVSS.n1918 VSS 0.082541f
C10940 DVSS.n1919 VSS 0.3147f
C10941 DVSS.n1920 VSS 0.052308f
C10942 DVSS.n1921 VSS 0.052308f
C10943 DVSS.n1922 VSS 0.052308f
C10944 DVSS.n1923 VSS 0.052308f
C10945 DVSS.n1924 VSS 0.052308f
C10946 DVSS.n1925 VSS 0.072078f
C10947 DVSS.n1927 VSS 0.163885f
C10948 DVSS.n1929 VSS 0.052308f
C10949 DVSS.n1931 VSS 0.052308f
C10950 DVSS.n1933 VSS 0.052308f
C10951 DVSS.n1934 VSS 0.072078f
C10952 DVSS.n1935 VSS 0.165082f
C10953 DVSS.n1936 VSS 0.165082f
C10954 DVSS.n1937 VSS 0.165082f
C10955 DVSS.n1938 VSS 0.165082f
C10956 DVSS.n1939 VSS 0.072078f
C10957 DVSS.n1940 VSS 0.165082f
C10958 DVSS.n1941 VSS 0.611712f
C10959 DVSS.n1942 VSS 0.165082f
C10960 DVSS.n1943 VSS 0.165082f
C10961 DVSS.n1944 VSS 0.165082f
C10962 DVSS.n1945 VSS 0.082541f
C10963 DVSS.n1946 VSS 0.165082f
C10964 DVSS.n1947 VSS 0.165082f
C10965 DVSS.n1948 VSS 0.165082f
C10966 DVSS.n1949 VSS 0.072078f
C10967 DVSS.n1950 VSS 0.082541f
C10968 DVSS.n1951 VSS 0.052308f
C10969 DVSS.n1952 VSS 0.052308f
C10970 DVSS.n1953 VSS 0.052308f
C10971 DVSS.n1954 VSS 0.052308f
C10972 DVSS.n1955 VSS 0.052308f
C10973 DVSS.n1956 VSS 0.072078f
C10974 DVSS.n1958 VSS 0.157135f
C10975 DVSS.n1960 VSS 0.052308f
C10976 DVSS.n1962 VSS 0.052308f
C10977 DVSS.n1964 VSS 0.052308f
C10978 DVSS.n1966 VSS 0.052308f
C10979 DVSS.n1967 VSS 0.165082f
C10980 DVSS.n1968 VSS 0.165082f
C10981 DVSS.n1969 VSS 0.165082f
C10982 DVSS.n1970 VSS 0.165082f
C10983 DVSS.n1971 VSS 0.082541f
C10984 DVSS.n1972 VSS 0.165082f
C10985 DVSS.n1973 VSS 0.165082f
C10986 DVSS.n1974 VSS 0.165082f
C10987 DVSS.n1975 VSS 0.072078f
C10988 DVSS.n1976 VSS 0.082541f
C10989 DVSS.n1977 VSS 0.052308f
C10990 DVSS.n1978 VSS 0.052308f
C10991 DVSS.n1979 VSS 0.052308f
C10992 DVSS.n1980 VSS 0.052308f
C10993 DVSS.n1981 VSS 0.052308f
C10994 DVSS.n1982 VSS 0.072078f
C10995 DVSS.n1984 VSS 0.157135f
C10996 DVSS.n1986 VSS 0.052308f
C10997 DVSS.n1988 VSS 0.052308f
C10998 DVSS.n1990 VSS 0.052308f
C10999 DVSS.n1992 VSS 0.052308f
C11000 DVSS.n1993 VSS 0.165082f
C11001 DVSS.n1994 VSS 0.165082f
C11002 DVSS.n1995 VSS 0.165082f
C11003 DVSS.n1996 VSS 0.165082f
C11004 DVSS.n1997 VSS 0.165082f
C11005 DVSS.n1998 VSS 0.165082f
C11006 DVSS.n1999 VSS 0.165082f
C11007 DVSS.n2000 VSS 0.165082f
C11008 DVSS.n2001 VSS 0.165082f
C11009 DVSS.n2002 VSS 0.165082f
C11010 DVSS.n2003 VSS 0.165082f
C11011 DVSS.n2004 VSS 0.165082f
C11012 DVSS.n2005 VSS 0.082541f
C11013 DVSS.n2006 VSS 0.165082f
C11014 DVSS.n2007 VSS 0.165082f
C11015 DVSS.n2008 VSS 0.165082f
C11016 DVSS.n2009 VSS 0.072078f
C11017 DVSS.n2010 VSS 0.082541f
C11018 DVSS.n2011 VSS 0.052308f
C11019 DVSS.n2012 VSS 0.052308f
C11020 DVSS.n2013 VSS 0.052308f
C11021 DVSS.n2014 VSS 0.052308f
C11022 DVSS.n2015 VSS 0.052308f
C11023 DVSS.n2016 VSS 0.072078f
C11024 DVSS.n2018 VSS 0.157135f
C11025 DVSS.n2020 VSS 0.052308f
C11026 DVSS.n2022 VSS 0.052308f
C11027 DVSS.n2024 VSS 0.052308f
C11028 DVSS.n2026 VSS 0.052308f
C11029 DVSS.n2027 VSS 0.165082f
C11030 DVSS.n2028 VSS 0.165082f
C11031 DVSS.n2029 VSS 0.165082f
C11032 DVSS.n2030 VSS 0.165082f
C11033 DVSS.n2031 VSS 0.165082f
C11034 DVSS.n2032 VSS 0.165082f
C11035 DVSS.n2033 VSS 0.165082f
C11036 DVSS.n2034 VSS 0.165082f
C11037 DVSS.n2035 VSS 0.165082f
C11038 DVSS.n2036 VSS 0.165082f
C11039 DVSS.n2037 VSS 0.165082f
C11040 DVSS.n2038 VSS 0.165082f
C11041 DVSS.n2039 VSS 0.082541f
C11042 DVSS.n2040 VSS 0.165082f
C11043 DVSS.n2041 VSS 0.165082f
C11044 DVSS.n2042 VSS 0.165082f
C11045 DVSS.n2043 VSS 0.072078f
C11046 DVSS.n2044 VSS 0.082541f
C11047 DVSS.n2045 VSS 0.019102f
C11048 DVSS.n2046 VSS 0.019102f
C11049 DVSS.n2047 VSS 0.019102f
C11050 DVSS.n2048 VSS 0.019102f
C11051 DVSS.n2049 VSS 0.019102f
C11052 DVSS.n2050 VSS 0.10928f
C11053 DVSS.n2051 VSS 0.019102f
C11054 DVSS.n2052 VSS 0.019102f
C11055 DVSS.n2053 VSS 0.019102f
C11056 DVSS.n2054 VSS 0.019102f
C11057 DVSS.n2055 VSS 0.019102f
C11058 DVSS.n2056 VSS 0.021932f
C11059 DVSS.n2057 VSS 0.038205f
C11060 DVSS.n2058 VSS 0.026905f
C11061 DVSS.n2059 VSS 0.021932f
C11062 DVSS.n2060 VSS 0.082541f
C11063 DVSS.n2061 VSS 0.082541f
C11064 DVSS.n2062 VSS 0.111605f
C11065 DVSS.n2063 VSS 0.019102f
C11066 DVSS.n2064 VSS 0.019102f
C11067 DVSS.n2065 VSS 0.019102f
C11068 DVSS.n2066 VSS 0.019102f
C11069 DVSS.n2067 VSS 0.019102f
C11070 DVSS.n2068 VSS 0.072078f
C11071 DVSS.n2069 VSS 0.019102f
C11072 DVSS.n2070 VSS 0.019102f
C11073 DVSS.n2071 VSS 0.019102f
C11074 DVSS.n2072 VSS 0.019102f
C11075 DVSS.n2073 VSS 0.021932f
C11076 DVSS.n2074 VSS 0.035873f
C11077 DVSS.n2075 VSS 0.024232f
C11078 DVSS.n2076 VSS 0.066505f
C11079 DVSS.n2077 VSS 0.031887f
C11080 DVSS.n2079 VSS 0.065379f
C11081 DVSS.n2080 VSS 0.066724f
C11082 DVSS.n2082 VSS 0.043865f
C11083 DVSS.n2085 VSS 0.052308f
C11084 DVSS.n2086 VSS 0.754249f
C11085 DVSS.n2088 VSS 0.066724f
C11086 DVSS.n2089 VSS 0.052308f
C11087 DVSS.t18 VSS 0.394423f
C11088 DVSS.n2090 VSS 0.635269f
C11089 DVSS.n2093 VSS 0.052308f
C11090 DVSS.n2094 VSS 0.754249f
C11091 DVSS.n2096 VSS 0.066724f
C11092 DVSS.n2098 VSS 0.052308f
C11093 DVSS.n2101 VSS 0.052308f
C11094 DVSS.n2102 VSS 0.754249f
C11095 DVSS.n2104 VSS 0.066724f
C11096 DVSS.n2105 VSS 0.052308f
C11097 DVSS.n2108 VSS 0.045559f
C11098 DVSS.n2109 VSS 0.058114f
C11099 DVSS.n2112 VSS 0.21755f
C11100 DVSS.n2114 VSS 0.045559f
C11101 DVSS.n2115 VSS 0.045559f
C11102 DVSS.n2116 VSS 0.331802f
C11103 DVSS.n2119 VSS 0.779994f
C11104 DVSS.n2120 VSS 0.176874f
C11105 DVSS.n2121 VSS 0.145734f
C11106 DVSS.n2122 VSS 0.052308f
C11107 DVSS.n2123 VSS 0.052308f
C11108 DVSS.n2124 VSS 0.052308f
C11109 DVSS.n2125 VSS 0.052308f
C11110 DVSS.n2126 VSS 0.052308f
C11111 DVSS.n2127 VSS 0.052308f
C11112 DVSS.n2128 VSS 0.052308f
C11113 DVSS.n2129 VSS 0.052308f
C11114 DVSS.n2130 VSS 0.052308f
C11115 DVSS.n2131 VSS 0.052308f
C11116 DVSS.n2132 VSS 0.052308f
C11117 DVSS.n2133 VSS 0.140683f
C11118 DVSS.n2134 VSS 0.154453f
C11119 DVSS.n2136 VSS 0.052308f
C11120 DVSS.n2138 VSS 0.052308f
C11121 DVSS.n2140 VSS 0.052308f
C11122 DVSS.n2142 VSS 0.052308f
C11123 DVSS.n2144 VSS 0.052308f
C11124 DVSS.n2146 VSS 0.052308f
C11125 DVSS.n2148 VSS 0.052308f
C11126 DVSS.n2150 VSS 0.052308f
C11127 DVSS.n2152 VSS 0.052308f
C11128 DVSS.n2154 VSS 0.052308f
C11129 DVSS.n2155 VSS 0.353747f
C11130 DVSS.n2156 VSS 0.353747f
C11131 DVSS.n2157 VSS 0.318871f
C11132 DVSS.n2158 VSS 0.310152f
C11133 DVSS.n2159 VSS 0.353747f
C11134 DVSS.n2160 VSS 0.353747f
C11135 DVSS.n2161 VSS 0.353747f
C11136 DVSS.n2162 VSS 0.176874f
C11137 DVSS.n2174 VSS 0.133934f
C11138 DVSS.n2176 VSS 0.044926f
C11139 DVSS.n2177 VSS 0.287731f
C11140 DVSS.n2178 VSS 0.052308f
C11141 DVSS.n2179 VSS 0.052308f
C11142 DVSS.n2180 VSS 0.052308f
C11143 DVSS.n2181 VSS 0.052308f
C11144 DVSS.n2182 VSS 0.052308f
C11145 DVSS.n2183 VSS 0.052308f
C11146 DVSS.n2184 VSS 0.052308f
C11147 DVSS.n2185 VSS 0.052308f
C11148 DVSS.n2186 VSS 0.052308f
C11149 DVSS.n2187 VSS 0.052308f
C11150 DVSS.n2188 VSS 0.052308f
C11151 DVSS.n2189 VSS 0.353747f
C11152 DVSS.n2190 VSS 0.353747f
C11153 DVSS.n2191 VSS 0.353747f
C11154 DVSS.n2192 VSS 0.310152f
C11155 DVSS.n2193 VSS 0.353747f
C11156 DVSS.n2194 VSS 0.353747f
C11157 DVSS.n2195 VSS 0.353747f
C11158 DVSS.n2196 VSS 0.176874f
C11159 DVSS.n2208 VSS 0.133934f
C11160 DVSS.n2210 VSS 0.044926f
C11161 DVSS.n2211 VSS 0.287731f
C11162 DVSS.n2212 VSS 0.052308f
C11163 DVSS.n2213 VSS 0.052308f
C11164 DVSS.n2214 VSS 0.052308f
C11165 DVSS.n2215 VSS 0.052308f
C11166 DVSS.n2216 VSS 0.052308f
C11167 DVSS.n2217 VSS 0.052308f
C11168 DVSS.n2218 VSS 0.052308f
C11169 DVSS.n2219 VSS 0.052308f
C11170 DVSS.n2220 VSS 0.052308f
C11171 DVSS.n2221 VSS 0.052308f
C11172 DVSS.n2222 VSS 0.052308f
C11173 DVSS.n2223 VSS 0.353747f
C11174 DVSS.n2224 VSS 0.353747f
C11175 DVSS.n2225 VSS 0.353747f
C11176 DVSS.n2226 VSS 0.353747f
C11177 DVSS.n2227 VSS 0.353747f
C11178 DVSS.n2228 VSS 0.353747f
C11179 DVSS.n2229 VSS 0.353747f
C11180 DVSS.n2230 VSS 0.353747f
C11181 DVSS.n2231 VSS 0.353747f
C11182 DVSS.n2232 VSS 0.353747f
C11183 DVSS.n2233 VSS 0.353747f
C11184 DVSS.n2234 VSS 0.310152f
C11185 DVSS.n2235 VSS 0.353747f
C11186 DVSS.n2236 VSS 0.353747f
C11187 DVSS.n2237 VSS 0.353747f
C11188 DVSS.n2238 VSS 0.176874f
C11189 DVSS.n2250 VSS 0.133934f
C11190 DVSS.n2252 VSS 0.044926f
C11191 DVSS.n2253 VSS 0.287731f
C11192 DVSS.n2254 VSS 0.052308f
C11193 DVSS.n2255 VSS 0.052308f
C11194 DVSS.n2256 VSS 0.052308f
C11195 DVSS.n2257 VSS 0.052308f
C11196 DVSS.n2258 VSS 0.052308f
C11197 DVSS.n2259 VSS 0.052308f
C11198 DVSS.n2260 VSS 0.052308f
C11199 DVSS.n2261 VSS 0.052308f
C11200 DVSS.n2262 VSS 0.052308f
C11201 DVSS.n2263 VSS 0.052308f
C11202 DVSS.n2264 VSS 0.052308f
C11203 DVSS.n2265 VSS 0.353747f
C11204 DVSS.n2266 VSS 0.353747f
C11205 DVSS.n2267 VSS 0.353747f
C11206 DVSS.n2268 VSS 0.353747f
C11207 DVSS.n2269 VSS 0.353747f
C11208 DVSS.n2270 VSS 0.353747f
C11209 DVSS.n2271 VSS 0.353747f
C11210 DVSS.n2272 VSS 0.353747f
C11211 DVSS.n2273 VSS 0.353747f
C11212 DVSS.n2274 VSS 0.353747f
C11213 DVSS.n2275 VSS 0.353747f
C11214 DVSS.n2276 VSS 0.336309f
C11215 DVSS.n2277 VSS 0.353747f
C11216 DVSS.n2278 VSS 0.353747f
C11217 DVSS.n2279 VSS 0.353747f
C11218 DVSS.n2280 VSS 0.176874f
C11219 DVSS.n2281 VSS 0.03166f
C11220 DVSS.n2282 VSS 0.019102f
C11221 DVSS.n2283 VSS 0.019102f
C11222 DVSS.n2284 VSS 0.019102f
C11223 DVSS.n2285 VSS 0.019102f
C11224 DVSS.n2286 VSS 0.019102f
C11225 DVSS.n2287 VSS 0.019102f
C11226 DVSS.n2288 VSS 0.019102f
C11227 DVSS.n2289 VSS 0.019102f
C11228 DVSS.n2290 VSS 0.019102f
C11229 DVSS.n2291 VSS 0.019102f
C11230 DVSS.n2292 VSS 0.019102f
C11231 DVSS.n2293 VSS 0.019102f
C11232 DVSS.n2294 VSS 0.019102f
C11233 DVSS.n2295 VSS 0.019102f
C11234 DVSS.n2296 VSS 0.019102f
C11235 DVSS.n2297 VSS 0.019102f
C11236 DVSS.n2298 VSS 0.019102f
C11237 DVSS.n2299 VSS 0.019102f
C11238 DVSS.n2300 VSS 0.019102f
C11239 DVSS.n2301 VSS 0.019102f
C11240 DVSS.n2302 VSS 0.019102f
C11241 DVSS.n2303 VSS 0.019102f
C11242 DVSS.n2305 VSS 0.037674f
C11243 DVSS.n2306 VSS 0.234171f
C11244 DVSS.n2307 VSS 0.353747f
C11245 DVSS.n2308 VSS 0.353747f
C11246 DVSS.n2309 VSS 0.353747f
C11247 DVSS.n2310 VSS 0.176874f
C11248 DVSS.n2311 VSS 0.03166f
C11249 DVSS.n2312 VSS 0.019102f
C11250 DVSS.n2313 VSS 0.019102f
C11251 DVSS.n2314 VSS 0.019102f
C11252 DVSS.n2315 VSS 0.019102f
C11253 DVSS.n2316 VSS 0.019102f
C11254 DVSS.n2317 VSS 0.019102f
C11255 DVSS.n2318 VSS 0.019102f
C11256 DVSS.n2319 VSS 0.019102f
C11257 DVSS.n2320 VSS 0.019102f
C11258 DVSS.n2321 VSS 0.019102f
C11259 DVSS.n2322 VSS 0.019102f
C11260 DVSS.n2323 VSS 0.019102f
C11261 DVSS.n2324 VSS 0.019102f
C11262 DVSS.n2325 VSS 0.019102f
C11263 DVSS.n2326 VSS 0.019102f
C11264 DVSS.n2327 VSS 0.019102f
C11265 DVSS.n2328 VSS 0.019102f
C11266 DVSS.n2329 VSS 0.019102f
C11267 DVSS.n2330 VSS 0.019102f
C11268 DVSS.n2331 VSS 0.019102f
C11269 DVSS.n2332 VSS 0.019102f
C11270 DVSS.n2333 VSS 0.019102f
C11271 DVSS.n2335 VSS 0.037674f
C11272 DVSS.n2336 VSS 0.353747f
C11273 DVSS.n2337 VSS 0.353747f
C11274 DVSS.n2338 VSS 0.353747f
C11275 DVSS.n2339 VSS 0.353747f
C11276 DVSS.n2340 VSS 0.353747f
C11277 DVSS.n2341 VSS 0.353747f
C11278 DVSS.n2342 VSS 0.353747f
C11279 DVSS.n2343 VSS 0.353747f
C11280 DVSS.n2344 VSS 0.353747f
C11281 DVSS.n2345 VSS 0.353747f
C11282 DVSS.n2346 VSS 0.353747f
C11283 DVSS.n2347 VSS 0.353747f
C11284 DVSS.n2348 VSS 0.176874f
C11285 DVSS.n2349 VSS 0.353747f
C11286 DVSS.n2350 VSS 0.353747f
C11287 DVSS.n2351 VSS 0.353747f
C11288 DVSS.n2352 VSS 0.176874f
C11289 DVSS.n2353 VSS 0.052308f
C11290 DVSS.n2354 VSS 0.052308f
C11291 DVSS.n2355 VSS 0.052308f
C11292 DVSS.n2356 VSS 0.052308f
C11293 DVSS.n2357 VSS 0.052308f
C11294 DVSS.n2358 VSS 0.052308f
C11295 DVSS.n2359 VSS 0.052308f
C11296 DVSS.n2360 VSS 0.052308f
C11297 DVSS.n2361 VSS 0.052308f
C11298 DVSS.n2362 VSS 0.052308f
C11299 DVSS.n2363 VSS 0.052308f
C11300 DVSS.n2364 VSS 0.133934f
C11301 DVSS.n2365 VSS 0.154453f
C11302 DVSS.n2368 VSS 0.052308f
C11303 DVSS.n2371 VSS 0.052308f
C11304 DVSS.n2374 VSS 0.052308f
C11305 DVSS.n2377 VSS 0.052308f
C11306 DVSS.n2380 VSS 0.052308f
C11307 DVSS.n2383 VSS 0.052308f
C11308 DVSS.n2386 VSS 0.052308f
C11309 DVSS.n2389 VSS 0.052308f
C11310 DVSS.n2392 VSS 0.052308f
C11311 DVSS.n2395 VSS 0.052308f
C11312 DVSS.n2398 VSS 0.052308f
C11313 DVSS.n2400 VSS 0.044926f
C11314 DVSS.n2401 VSS 0.353747f
C11315 DVSS.n2402 VSS 0.353747f
C11316 DVSS.n2403 VSS 0.353747f
C11317 DVSS.n2404 VSS 0.353747f
C11318 DVSS.n2405 VSS 0.353747f
C11319 DVSS.n2406 VSS 0.353747f
C11320 DVSS.n2407 VSS 0.353747f
C11321 DVSS.n2408 VSS 0.353747f
C11322 DVSS.n2409 VSS 0.353747f
C11323 DVSS.n2410 VSS 0.353747f
C11324 DVSS.n2411 VSS 0.353747f
C11325 DVSS.n2412 VSS 0.353747f
C11326 DVSS.n2413 VSS 0.176874f
C11327 DVSS.n2414 VSS 0.353747f
C11328 DVSS.n2415 VSS 0.353747f
C11329 DVSS.n2416 VSS 0.353747f
C11330 DVSS.n2417 VSS 0.176874f
C11331 DVSS.n2418 VSS 0.052308f
C11332 DVSS.n2419 VSS 0.052308f
C11333 DVSS.n2420 VSS 0.052308f
C11334 DVSS.n2421 VSS 0.052308f
C11335 DVSS.n2422 VSS 0.052308f
C11336 DVSS.n2423 VSS 0.052308f
C11337 DVSS.n2424 VSS 0.052308f
C11338 DVSS.n2425 VSS 0.052308f
C11339 DVSS.n2426 VSS 0.052308f
C11340 DVSS.n2427 VSS 0.052308f
C11341 DVSS.n2428 VSS 0.052308f
C11342 DVSS.n2429 VSS 0.133934f
C11343 DVSS.n2430 VSS 0.154453f
C11344 DVSS.n2432 VSS 0.052308f
C11345 DVSS.n2435 VSS 0.052308f
C11346 DVSS.n2438 VSS 0.052308f
C11347 DVSS.n2441 VSS 0.052308f
C11348 DVSS.n2444 VSS 0.052308f
C11349 DVSS.n2447 VSS 0.052308f
C11350 DVSS.n2450 VSS 0.052308f
C11351 DVSS.n2453 VSS 0.052308f
C11352 DVSS.n2456 VSS 0.052308f
C11353 DVSS.n2459 VSS 0.052308f
C11354 DVSS.n2462 VSS 0.052308f
C11355 DVSS.n2464 VSS 0.044926f
C11356 DVSS.n2465 VSS 0.353747f
C11357 DVSS.n2466 VSS 0.353747f
C11358 DVSS.n2467 VSS 0.353747f
C11359 DVSS.n2468 VSS 0.353747f
C11360 DVSS.n2469 VSS 0.176874f
C11361 DVSS.n2470 VSS 0.353747f
C11362 DVSS.n2471 VSS 0.353747f
C11363 DVSS.n2472 VSS 0.353747f
C11364 DVSS.n2473 VSS 0.176874f
C11365 DVSS.n2474 VSS 0.052308f
C11366 DVSS.n2475 VSS 0.052308f
C11367 DVSS.n2476 VSS 0.052308f
C11368 DVSS.n2477 VSS 0.052308f
C11369 DVSS.n2478 VSS 0.052308f
C11370 DVSS.n2479 VSS 0.052308f
C11371 DVSS.n2480 VSS 0.052308f
C11372 DVSS.n2481 VSS 0.052308f
C11373 DVSS.n2482 VSS 0.052308f
C11374 DVSS.n2483 VSS 0.052308f
C11375 DVSS.n2484 VSS 0.052308f
C11376 DVSS.n2485 VSS 0.042673f
C11377 DVSS.n2486 VSS 0.154453f
C11378 DVSS.n2489 VSS 0.052308f
C11379 DVSS.n2492 VSS 0.052308f
C11380 DVSS.n2495 VSS 0.052308f
C11381 DVSS.n2498 VSS 0.052308f
C11382 DVSS.n2501 VSS 0.052308f
C11383 DVSS.n2504 VSS 0.052308f
C11384 DVSS.n2507 VSS 0.052308f
C11385 DVSS.n2510 VSS 0.052308f
C11386 DVSS.n2513 VSS 0.052308f
C11387 DVSS.n2516 VSS 0.052308f
C11388 DVSS.n2519 VSS 0.052308f
C11389 DVSS.n2521 VSS 0.044926f
C11390 DVSS.n2522 VSS 0.353747f
C11391 DVSS.n2523 VSS 0.353747f
C11392 DVSS.n2524 VSS 0.353747f
C11393 DVSS.n2525 VSS 0.353747f
C11394 DVSS.n2526 VSS 0.176874f
C11395 DVSS.n2527 VSS 0.353747f
C11396 DVSS.n2528 VSS 0.672799f
C11397 DVSS.n2529 VSS 0.353747f
C11398 DVSS.n2530 VSS 0.176874f
C11399 DVSS.n2531 VSS 0.052308f
C11400 DVSS.n2532 VSS 0.052308f
C11401 DVSS.n2533 VSS 0.052308f
C11402 DVSS.n2534 VSS 0.052308f
C11403 DVSS.n2535 VSS 0.052308f
C11404 DVSS.n2536 VSS 0.052308f
C11405 DVSS.n2537 VSS 0.052308f
C11406 DVSS.n2538 VSS 0.052308f
C11407 DVSS.n2539 VSS 0.052308f
C11408 DVSS.n2540 VSS 0.052308f
C11409 DVSS.n2541 VSS 0.052308f
C11410 DVSS.n2542 VSS 0.140683f
C11411 DVSS.n2543 VSS 0.154453f
C11412 DVSS.n2546 VSS 0.052308f
C11413 DVSS.n2549 VSS 0.052308f
C11414 DVSS.n2552 VSS 0.052308f
C11415 DVSS.n2555 VSS 0.052308f
C11416 DVSS.n2558 VSS 0.052308f
C11417 DVSS.n2561 VSS 0.052308f
C11418 DVSS.n2564 VSS 0.052308f
C11419 DVSS.n2567 VSS 0.052308f
C11420 DVSS.n2570 VSS 0.052308f
C11421 DVSS.n2573 VSS 0.052308f
C11422 DVSS.n2576 VSS 0.052308f
C11423 DVSS.n2579 VSS 0.041971f
C11424 DVSS.n2581 VSS 0.045559f
C11425 DVSS.t0 VSS 0.394423f
C11426 DVSS.n2582 VSS 0.331802f
C11427 DVSS.n2584 VSS 0.045559f
C11428 DVSS.n2585 VSS 0.058114f
C11429 DVSS.n2588 VSS 0.041971f
C11430 DVSS.n2590 VSS 0.045559f
C11431 DVSS.t20 VSS 0.394423f
C11432 DVSS.n2593 VSS 0.052308f
C11433 DVSS.n2594 VSS 0.754249f
C11434 DVSS.n2596 VSS 0.066724f
C11435 DVSS.n2597 VSS 0.052308f
C11436 DVSS.n2600 VSS 0.052308f
C11437 DVSS.n2601 VSS 0.754249f
C11438 DVSS.n2603 VSS 0.066724f
C11439 DVSS.n2604 VSS 0.052308f
C11440 DVSS.t17 VSS 0.330478f
C11441 DVSS.n2605 VSS 0.635269f
C11442 DVSS.n2608 VSS 0.052308f
C11443 DVSS.n2609 VSS 0.754249f
C11444 DVSS.n2611 VSS 0.066724f
C11445 DVSS.n2612 VSS 0.052308f
C11446 DVSS.n2615 VSS 0.069335f
C11447 DVSS.n2617 VSS 0.066724f
C11448 DVSS.n2619 VSS 0.043865f
C11449 DVSS.n2620 VSS 0.043865f
C11450 DVSS.n2621 VSS 0.065379f
C11451 DVSS.n2622 VSS 0.038205f
C11452 DVSS.n2623 VSS 0.035873f
C11453 DVSS.n2624 VSS -0.427302f
C11454 DVSS.n2625 VSS 0.038205f
C11455 DVSS.n2626 VSS 0.035873f
C11456 DVSS.n2627 VSS 0.038205f
C11457 DVSS.n2628 VSS 0.035873f
C11458 DVSS.n2629 VSS 0.038205f
C11459 DVSS.n2630 VSS 0.035873f
C11460 DVSS.n2631 VSS 0.038205f
C11461 DVSS.n2632 VSS 0.035873f
C11462 DVSS.n2633 VSS 0.038205f
C11463 DVSS.n2634 VSS 0.033714f
C11464 DVSS.n2635 VSS 0.038205f
C11465 DVSS.n2636 VSS 0.026905f
C11466 DVSS.n2637 VSS 0.038205f
C11467 DVSS.n2638 VSS 0.035873f
C11468 DVSS.t34 VSS 0.330478f
C11469 DVSS.n2639 VSS 0.125906f
C11470 DVSS.n2640 VSS 0.038205f
C11471 DVSS.n2641 VSS 0.035873f
C11472 DVSS.n2642 VSS 0.038205f
C11473 DVSS.n2643 VSS 0.035873f
C11474 DVSS.n2644 VSS 0.038205f
C11475 DVSS.n2645 VSS 0.035873f
C11476 DVSS.n2646 VSS 0.038205f
C11477 DVSS.n2647 VSS 0.035873f
C11478 DVSS.n2648 VSS 0.038205f
C11479 DVSS.n2649 VSS 0.035873f
C11480 DVSS.n2650 VSS 0.066505f
C11481 DVSS.n2651 VSS 0.031887f
C11482 DVSS.n2653 VSS 0.066724f
C11483 DVSS.n2655 VSS 0.052308f
C11484 DVSS.n2656 VSS 0.052308f
C11485 DVSS.t30 VSS 0.330478f
C11486 DVSS.n2660 VSS 0.635269f
C11487 DVSS.n2661 VSS 0.066724f
C11488 DVSS.n2663 VSS 0.052308f
C11489 DVSS.n2664 VSS 0.052308f
C11490 DVSS.n2668 VSS 0.066724f
C11491 DVSS.n2670 VSS 0.052308f
C11492 DVSS.n2671 VSS 0.052308f
C11493 DVSS.n2676 VSS 0.222771f
C11494 DVSS.n2678 VSS 0.066724f
C11495 DVSS.n2679 VSS 0.052308f
C11496 DVSS.n2680 VSS 0.179185f
C11497 DVSS.n2682 VSS 0.09309f
C11498 DVSS.n2684 VSS 0.066724f
C11499 DVSS.n2685 VSS 0.052308f
C11500 DVSS.n2686 VSS 0.335771f
C11501 DVSS.n2687 VSS 0.756156f
C11502 DVSS.n2689 VSS 0.242143f
C11503 DVSS.n2691 VSS 0.066724f
C11504 DVSS.n2692 VSS 0.052308f
C11505 DVSS.n2693 VSS 0.186719f
C11506 DVSS.n2694 VSS 0.396845f
C11507 DVSS.n2696 VSS 0.066724f
C11508 DVSS.n2698 VSS 0.043865f
C11509 DVSS.n2699 VSS 0.021932f
C11510 DVSS.n2700 VSS 0.021932f
C11511 DVSS.n2701 VSS 0.049824f
C11512 DVSS.n2704 VSS 0.069335f
C11513 DVSS.n2706 VSS 0.066724f
C11514 DVSS.n2708 VSS 0.043865f
C11515 DVSS.n2712 VSS 0.066724f
C11516 DVSS.n2714 VSS 0.066724f
C11517 DVSS.n2716 VSS 0.052308f
C11518 DVSS.t27 VSS 0.394423f
C11519 DVSS.n2717 VSS 0.635269f
C11520 DVSS.n2721 VSS 0.066724f
C11521 DVSS.n2723 VSS 0.066724f
C11522 DVSS.n2725 VSS 0.052308f
C11523 DVSS.n2729 VSS 0.066724f
C11524 DVSS.n2731 VSS 0.066724f
C11525 DVSS.n2733 VSS 0.052308f
C11526 DVSS.n2734 VSS 0.052308f
C11527 DVSS.n2735 VSS 0.222771f
C11528 DVSS.n2736 VSS 0.052308f
C11529 DVSS.n2738 VSS 0.179185f
C11530 DVSS.n2739 VSS 0.052308f
C11531 DVSS.n2740 VSS 0.09309f
C11532 DVSS.n2741 VSS 0.052308f
C11533 DVSS.n2743 VSS 0.335771f
C11534 DVSS.n2744 VSS 0.756156f
C11535 DVSS.n2745 VSS 0.052308f
C11536 DVSS.n2746 VSS 0.242143f
C11537 DVSS.n2747 VSS 0.052308f
C11538 DVSS.n2749 VSS 0.186719f
C11539 DVSS.n2750 VSS 0.043865f
C11540 DVSS.n2751 VSS 0.396845f
C11541 DVSS.n2753 VSS 0.043865f
C11542 DVSS.n2754 VSS 0.065379f
C11543 DVSS.n2755 VSS 36.516f
C11544 DVSS.n2756 VSS 2.56489f
C11545 DVSS.n2757 VSS 47.205f
C11546 DVSS.n2758 VSS 48.8624f
C11547 DVSS.n2759 VSS 0.028093f
C11548 DVSS.n2761 VSS 0.021932f
C11549 DVSS.n2762 VSS 0.036967f
C11550 DVSS.n2763 VSS 0.032106f
C11551 DVSS.n2764 VSS 0.019102f
C11552 DVSS.n2766 VSS 0.032106f
C11553 DVSS.n2768 VSS 0.026154f
C11554 DVSS.n2770 VSS 0.044082f
C11555 DVSS.n2771 VSS 0.032106f
C11556 DVSS.n2772 VSS 0.032106f
C11557 DVSS.n2773 VSS 0.022779f
C11558 DVSS.n2775 VSS 0.032106f
C11559 DVSS.n2777 VSS 0.289551f
C11560 DVSS.n2778 VSS 0.022779f
C11561 DVSS.n2781 VSS 0.075348f
C11562 DVSS.n2782 VSS 0.075348f
C11563 DVSS.n2783 VSS 0.122573f
C11564 DVSS.n2785 VSS 0.060323f
C11565 DVSS.n2786 VSS 0.439768f
C11566 DVSS.n2787 VSS 0.052308f
C11567 DVSS.n2788 VSS 0.052308f
C11568 DVSS.n2789 VSS 0.065797f
C11569 DVSS.n2791 VSS 0.052308f
C11570 DVSS.n2794 VSS 0.150696f
C11571 DVSS.n2795 VSS 0.150696f
C11572 DVSS.n2796 VSS 0.150696f
C11573 DVSS.n2797 VSS 0.150696f
C11574 DVSS.n2798 VSS 0.150696f
C11575 DVSS.n2799 VSS 0.150696f
C11576 DVSS.n2800 VSS 0.150696f
C11577 DVSS.n2801 VSS 0.150696f
C11578 DVSS.n2802 VSS 0.150696f
C11579 DVSS.n2803 VSS 0.150696f
C11580 DVSS.n2804 VSS 0.150696f
C11581 DVSS.n2805 VSS 0.150696f
C11582 DVSS.n2806 VSS 0.150696f
C11583 DVSS.n2807 VSS 0.150696f
C11584 DVSS.n2808 VSS 0.150696f
C11585 DVSS.n2809 VSS 0.150696f
C11586 DVSS.n2810 VSS 0.150696f
C11587 DVSS.n2811 VSS 0.150696f
C11588 DVSS.n2812 VSS 0.150696f
C11589 DVSS.n2813 VSS 0.150696f
C11590 DVSS.n2814 VSS 0.150696f
C11591 DVSS.n2815 VSS 0.150696f
C11592 DVSS.n2816 VSS 0.150696f
C11593 DVSS.n2817 VSS 0.060323f
C11594 DVSS.n2818 VSS 0.439768f
C11595 DVSS.n2819 VSS 0.052308f
C11596 DVSS.n2820 VSS 0.052308f
C11597 DVSS.n2821 VSS 0.022779f
C11598 DVSS.n2822 VSS 0.065797f
C11599 DVSS.n2823 VSS 0.041129f
C11600 DVSS.n2824 VSS 0.052308f
C11601 DVSS.n2825 VSS 0.052308f
C11602 DVSS.n2826 VSS 0.044082f
C11603 DVSS.n2827 VSS 0.026154f
C11604 DVSS.n2830 VSS 0.075348f
C11605 DVSS.n2831 VSS 0.026154f
C11606 DVSS.n2833 VSS 0.075348f
C11607 DVSS.n2837 VSS 0.150696f
C11608 DVSS.n2838 VSS 0.150696f
C11609 DVSS.n2839 VSS 0.150696f
C11610 DVSS.n2840 VSS 0.150696f
C11611 DVSS.n2841 VSS 0.150696f
C11612 DVSS.n2842 VSS 0.150696f
C11613 DVSS.n2843 VSS 0.150696f
C11614 DVSS.n2844 VSS 0.150696f
C11615 DVSS.n2845 VSS 0.150696f
C11616 DVSS.n2846 VSS 0.150696f
C11617 DVSS.n2847 VSS 0.150696f
C11618 DVSS.n2848 VSS 0.060323f
C11619 DVSS.n2849 VSS 0.439768f
C11620 DVSS.n2850 VSS 0.052308f
C11621 DVSS.n2851 VSS 0.052308f
C11622 DVSS.n2852 VSS 0.022779f
C11623 DVSS.n2853 VSS 0.065797f
C11624 DVSS.n2854 VSS 0.041129f
C11625 DVSS.n2855 VSS 0.052308f
C11626 DVSS.n2856 VSS 0.052308f
C11627 DVSS.n2857 VSS 0.044082f
C11628 DVSS.n2858 VSS 0.026154f
C11629 DVSS.n2863 VSS 0.075348f
C11630 DVSS.n2864 VSS 0.026154f
C11631 DVSS.n2865 VSS 0.075348f
C11632 DVSS.n2866 VSS 0.150696f
C11633 DVSS.n2867 VSS 0.150696f
C11634 DVSS.n2868 VSS 0.150696f
C11635 DVSS.n2869 VSS 0.150696f
C11636 DVSS.n2870 VSS 0.150696f
C11637 DVSS.n2871 VSS 0.135839f
C11638 DVSS.n2872 VSS 0.150696f
C11639 DVSS.n2873 VSS 0.150696f
C11640 DVSS.n2874 VSS 0.150696f
C11641 DVSS.n2875 VSS 0.077471f
C11642 DVSS.n2876 VSS 0.150696f
C11643 DVSS.n2877 VSS 0.060323f
C11644 DVSS.n2878 VSS 0.439768f
C11645 DVSS.n2879 VSS 0.052308f
C11646 DVSS.n2880 VSS 0.052308f
C11647 DVSS.n2881 VSS 0.022779f
C11648 DVSS.n2882 VSS 0.065797f
C11649 DVSS.n2883 VSS 0.041129f
C11650 DVSS.n2884 VSS 0.052308f
C11651 DVSS.n2885 VSS 0.052308f
C11652 DVSS.n2886 VSS 0.044082f
C11653 DVSS.n2887 VSS 0.026154f
C11654 DVSS.n2890 VSS 0.331907f
C11655 DVSS.n2893 VSS 0.032106f
C11656 DVSS.n2895 VSS 0.032106f
C11657 DVSS.n2897 VSS 0.032106f
C11658 DVSS.n2899 VSS 0.032106f
C11659 DVSS.n2901 VSS 0.032106f
C11660 DVSS.n2903 VSS 0.032106f
C11661 DVSS.n2905 VSS 0.026154f
C11662 DVSS.n2906 VSS 0.120696f
C11663 DVSS.n2907 VSS 0.120696f
C11664 DVSS.n2909 VSS 0.026154f
C11665 DVSS.n2910 VSS 0.127236f
C11666 DVSS.n2911 VSS 0.041971f
C11667 DVSS.n2912 VSS 0.21755f
C11668 DVSS.n2914 VSS 0.026154f
C11669 DVSS.n2915 VSS 0.746867f
C11670 DVSS.n2916 VSS 0.026154f
C11671 DVSS.n2917 VSS 0.022779f
C11672 DVSS.n2918 VSS 0.058114f
C11673 DVSS.n2919 VSS 0.044926f
C11674 DVSS.n2920 VSS 0.331802f
C11675 DVSS.n2922 VSS 0.082541f
C11676 DVSS.n2923 VSS 0.363609f
C11677 DVSS.n2924 VSS 0.082541f
C11678 DVSS.n2925 VSS 0.068009f
C11679 DVSS.n2926 VSS 0.052308f
C11680 DVSS.n2927 VSS 0.052308f
C11681 DVSS.n2929 VSS 0.052308f
C11682 DVSS.n2930 VSS 0.022779f
C11683 DVSS.n2931 VSS 0.072078f
C11684 DVSS.n2932 VSS 0.022779f
C11685 DVSS.n2935 VSS 0.052308f
C11686 DVSS.n2938 VSS 0.052308f
C11687 DVSS.n2941 VSS 0.363609f
C11688 DVSS.n2942 VSS 0.082541f
C11689 DVSS.n2943 VSS 0.068009f
C11690 DVSS.n2944 VSS 0.022779f
C11691 DVSS.n2945 VSS 0.022779f
C11692 DVSS.n2946 VSS 0.047879f
C11693 DVSS.n2947 VSS 0.052308f
C11694 DVSS.n2948 VSS 0.052308f
C11695 DVSS.n2949 VSS 0.072078f
C11696 DVSS.n2951 VSS 0.052308f
C11697 DVSS.n2953 VSS 0.052308f
C11698 DVSS.n2954 VSS 0.022779f
C11699 DVSS.n2955 VSS 0.022779f
C11700 DVSS.n2956 VSS 0.026154f
C11701 DVSS.n2959 VSS 0.082541f
C11702 DVSS.n2960 VSS 0.058114f
C11703 DVSS.n2962 VSS 0.331802f
C11704 DVSS.n2965 VSS 0.045559f
C11705 DVSS.n2966 VSS 0.045559f
C11706 DVSS.n2968 VSS 0.170965f
C11707 DVSS.n2969 VSS 0.058114f
C11708 DVSS.n2971 VSS 0.331802f
C11709 DVSS.n2974 VSS 0.045559f
C11710 DVSS.n2975 VSS 0.045559f
C11711 DVSS.n2977 VSS 36.516f
C11712 DVSS.n2978 VSS 0.170965f
C11713 DVSS.n2979 VSS 0.21755f
C11714 DVSS.n2980 VSS 0.21755f
C11715 DVSS.n2982 VSS 0.058114f
C11716 DVSS.n2985 VSS 0.045559f
C11717 DVSS.n2986 VSS 0.045559f
C11718 DVSS.t26 VSS 0.394423f
C11719 DVSS.n2987 VSS 0.32373f
C11720 DVSS.n2989 VSS 0.045559f
C11721 DVSS.n2991 VSS 0.048967f
C11722 DVSS.n2993 VSS 0.026154f
C11723 DVSS.n2994 VSS 0.082541f
C11724 DVSS.n2995 VSS 0.082541f
C11725 DVSS.n2996 VSS 0.082541f
C11726 DVSS.n2997 VSS 0.3147f
C11727 DVSS.n2998 VSS 0.022779f
C11728 DVSS.n2999 VSS 0.022779f
C11729 DVSS.n3000 VSS 0.047879f
C11730 DVSS.n3001 VSS 0.052308f
C11731 DVSS.n3002 VSS 0.052308f
C11732 DVSS.n3003 VSS 0.072078f
C11733 DVSS.n3005 VSS 0.439557f
C11734 DVSS.n3008 VSS 0.052308f
C11735 DVSS.n3011 VSS 0.052308f
C11736 DVSS.n3012 VSS 0.022779f
C11737 DVSS.n3013 VSS 0.026154f
C11738 DVSS.n3014 VSS 0.058114f
C11739 DVSS.n3015 VSS 0.048967f
C11740 DVSS.n3016 VSS 0.217854f
C11741 DVSS.n3017 VSS 0.026154f
C11742 DVSS.n3018 VSS 0.026154f
C11743 DVSS.n3020 VSS 0.746867f
C11744 DVSS.n3021 VSS 0.022779f
C11745 DVSS.n3022 VSS 0.058114f
C11746 DVSS.n3023 VSS 0.044926f
C11747 DVSS.t31 VSS 0.394423f
C11748 DVSS.n3025 VSS 0.32373f
C11749 DVSS.n3026 VSS 0.022779f
C11750 DVSS.n3027 VSS 0.082541f
C11751 DVSS.n3028 VSS 0.082541f
C11752 DVSS.n3029 VSS 0.082541f
C11753 DVSS.n3030 VSS 0.3147f
C11754 DVSS.n3031 VSS 0.052308f
C11755 DVSS.n3032 VSS 0.052308f
C11756 DVSS.n3034 VSS 0.052308f
C11757 DVSS.n3035 VSS 0.072078f
C11758 DVSS.n3036 VSS 0.165082f
C11759 DVSS.n3037 VSS 0.165082f
C11760 DVSS.n3038 VSS 0.165082f
C11761 DVSS.n3039 VSS 0.165082f
C11762 DVSS.n3040 VSS 0.165082f
C11763 DVSS.n3041 VSS 0.165082f
C11764 DVSS.n3042 VSS 0.165082f
C11765 DVSS.n3043 VSS 0.010297f
C11766 DVSS.n3044 VSS 0.020594f
C11767 DVSS.n3045 VSS 0.020594f
C11768 DVSS.n3046 VSS 0.010297f
C11769 DVSS.n3047 VSS 0.010297f
C11770 DVSS.n3048 VSS 0.072078f
C11771 DVSS.n3049 VSS 0.010297f
C11772 DVSS.n3050 VSS 0.010297f
C11773 DVSS.n3051 VSS 0.010297f
C11774 DVSS.n3052 VSS 0.020594f
C11775 DVSS.n3053 VSS 0.020594f
C11776 DVSS.n3054 VSS 0.128462f
C11777 DVSS.n3055 VSS 0.010297f
C11778 DVSS.n3056 VSS 0.129624f
C11779 DVSS.n3057 VSS 0.010297f
C11780 DVSS.n3058 VSS 0.010297f
C11781 DVSS.n3059 VSS 0.016193f
C11782 DVSS.n3060 VSS 0.020594f
C11783 DVSS.n3061 VSS 0.020594f
C11784 DVSS.n3062 VSS 0.072078f
C11785 DVSS.n3063 VSS 0.010297f
C11786 DVSS.n3064 VSS 0.010297f
C11787 DVSS.n3065 VSS 0.010297f
C11788 DVSS.n3066 VSS 0.292547f
C11789 DVSS.n3067 VSS 0.010297f
C11790 DVSS.n3068 VSS 0.020594f
C11791 DVSS.n3069 VSS 0.165082f
C11792 DVSS.n3070 VSS 0.165082f
C11793 DVSS.n3071 VSS 0.165082f
C11794 DVSS.n3072 VSS 0.165082f
C11795 DVSS.n3073 VSS 0.165082f
C11796 DVSS.n3074 VSS 0.131949f
C11797 DVSS.n3075 VSS 0.165082f
C11798 DVSS.n3076 VSS 0.611712f
C11799 DVSS.n3077 VSS 0.165082f
C11800 DVSS.n3078 VSS 0.072078f
C11801 DVSS.n3079 VSS 0.165082f
C11802 DVSS.n3080 VSS 0.072078f
C11803 DVSS.n3081 VSS 0.165082f
C11804 DVSS.n3082 VSS 0.165082f
C11805 DVSS.n3083 VSS 0.165082f
C11806 DVSS.n3084 VSS 0.165082f
C11807 DVSS.n3085 VSS 0.165082f
C11808 DVSS.n3086 VSS 0.165082f
C11809 DVSS.n3087 VSS 0.165082f
C11810 DVSS.n3088 VSS 0.165082f
C11811 DVSS.n3089 VSS 0.165082f
C11812 DVSS.n3090 VSS 0.165082f
C11813 DVSS.n3091 VSS 0.165082f
C11814 DVSS.n3092 VSS 0.165082f
C11815 DVSS.n3093 VSS 0.165082f
C11816 DVSS.n3094 VSS 0.165082f
C11817 DVSS.n3095 VSS 0.165082f
C11818 DVSS.n3096 VSS 0.165082f
C11819 DVSS.n3097 VSS 0.165082f
C11820 DVSS.n3098 VSS 0.165082f
C11821 DVSS.n3099 VSS 0.165082f
C11822 DVSS.n3100 VSS 0.026154f
C11823 DVSS.n3101 VSS 0.026154f
C11824 DVSS.n3102 VSS 0.041129f
C11825 DVSS.n3103 VSS 0.052308f
C11826 DVSS.n3104 VSS 0.052308f
C11827 DVSS.n3105 VSS 0.072078f
C11828 DVSS.n3106 VSS 0.439557f
C11829 DVSS.n3107 VSS 0.052308f
C11830 DVSS.n3108 VSS 0.052308f
C11831 DVSS.n3109 VSS 0.026154f
C11832 DVSS.n3110 VSS 0.026154f
C11833 DVSS.n3111 VSS 0.026154f
C11834 DVSS.n3112 VSS 0.082541f
C11835 DVSS.n3113 VSS 0.74307f
C11836 DVSS.n3117 VSS 0.082541f
C11837 DVSS.n3118 VSS 0.072078f
C11838 DVSS.n3119 VSS 0.165082f
C11839 DVSS.n3120 VSS 0.165082f
C11840 DVSS.n3121 VSS 0.165082f
C11841 DVSS.n3122 VSS 0.072078f
C11842 DVSS.n3123 VSS 0.165082f
C11843 DVSS.n3124 VSS 0.165082f
C11844 DVSS.n3125 VSS 0.165082f
C11845 DVSS.n3126 VSS 0.165082f
C11846 DVSS.n3127 VSS 0.165082f
C11847 DVSS.n3128 VSS 0.165082f
C11848 DVSS.n3129 VSS 0.165082f
C11849 DVSS.n3130 VSS 0.165082f
C11850 DVSS.n3131 VSS 0.165082f
C11851 DVSS.n3132 VSS 0.165082f
C11852 DVSS.n3133 VSS 0.165082f
C11853 DVSS.n3134 VSS 0.165082f
C11854 DVSS.n3135 VSS 0.165082f
C11855 DVSS.n3136 VSS 0.082541f
C11856 DVSS.n3137 VSS 0.165082f
C11857 DVSS.n3138 VSS 0.165082f
C11858 DVSS.n3139 VSS 0.165082f
C11859 DVSS.n3140 VSS 0.072078f
C11860 DVSS.n3141 VSS 0.082541f
C11861 DVSS.n3142 VSS 0.026154f
C11862 DVSS.n3143 VSS 0.026154f
C11863 DVSS.n3144 VSS 0.041129f
C11864 DVSS.n3145 VSS 0.052308f
C11865 DVSS.n3146 VSS 0.052308f
C11866 DVSS.n3147 VSS 0.072078f
C11867 DVSS.n3149 VSS 0.439557f
C11868 DVSS.n3151 VSS 0.052308f
C11869 DVSS.n3153 VSS 0.052308f
C11870 DVSS.n3154 VSS 0.026154f
C11871 DVSS.n3155 VSS 0.026154f
C11872 DVSS.n3156 VSS 0.026154f
C11873 DVSS.n3157 VSS 0.74307f
C11874 DVSS.n3158 VSS 0.165082f
C11875 DVSS.n3159 VSS 0.165082f
C11876 DVSS.n3160 VSS 0.165082f
C11877 DVSS.n3161 VSS 0.165082f
C11878 DVSS.n3162 VSS 0.165082f
C11879 DVSS.n3163 VSS 0.165082f
C11880 DVSS.n3164 VSS 0.165082f
C11881 DVSS.n3165 VSS 0.165082f
C11882 DVSS.n3166 VSS 0.165082f
C11883 DVSS.n3167 VSS 0.165082f
C11884 DVSS.n3168 VSS 0.165082f
C11885 DVSS.n3169 VSS 0.165082f
C11886 DVSS.n3170 VSS 0.082541f
C11887 DVSS.n3171 VSS 0.165082f
C11888 DVSS.n3172 VSS 0.165082f
C11889 DVSS.n3173 VSS 0.165082f
C11890 DVSS.n3174 VSS 0.072078f
C11891 DVSS.n3175 VSS 0.082541f
C11892 DVSS.n3176 VSS 0.021932f
C11893 DVSS.n3177 VSS 0.021932f
C11894 DVSS.n3178 VSS 0.03449f
C11895 DVSS.n3179 VSS 0.019102f
C11896 DVSS.n3180 VSS 0.019102f
C11897 DVSS.n3181 VSS 0.10928f
C11898 DVSS.n3182 VSS 0.019102f
C11899 DVSS.n3183 VSS 0.019102f
C11900 DVSS.n3185 VSS 0.034844f
C11901 DVSS.n3186 VSS 0.021932f
C11902 DVSS.n3187 VSS 0.021932f
C11903 DVSS.n3188 VSS 0.021932f
C11904 DVSS.n3189 VSS 0.038205f
C11905 DVSS.n3190 VSS 0.05713f
C11906 DVSS.n3191 VSS 0.038205f
C11907 DVSS.n3192 VSS 0.038205f
C11908 DVSS.n3193 VSS 0.035873f
C11909 DVSS.n3194 VSS 0.038205f
C11910 DVSS.n3195 VSS 0.038205f
C11911 DVSS.n3196 VSS 0.038205f
C11912 DVSS.n3197 VSS 0.038205f
C11913 DVSS.n3198 VSS 0.038205f
C11914 DVSS.n3199 VSS 0.035873f
C11915 DVSS.n3200 VSS 0.038205f
C11916 DVSS.n3201 VSS 0.038205f
C11917 DVSS.n3202 VSS 0.038205f
C11918 DVSS.n3203 VSS 0.038205f
C11919 DVSS.n3204 VSS 0.038205f
C11920 DVSS.n3205 VSS 0.035873f
C11921 DVSS.n3206 VSS 0.038205f
C11922 DVSS.n3207 VSS 0.038205f
C11923 DVSS.n3208 VSS 0.038205f
C11924 DVSS.n3209 VSS 0.038205f
C11925 DVSS.n3210 VSS 0.038205f
C11926 DVSS.n3211 VSS 0.020096f
C11927 DVSS.n3212 VSS 0.038205f
C11928 DVSS.n3213 VSS 0.038205f
C11929 DVSS.n3214 VSS 0.038205f
C11930 DVSS.n3215 VSS 0.038205f
C11931 DVSS.n3216 VSS 0.038205f
C11932 DVSS.n3217 VSS 0.035873f
C11933 DVSS.n3218 VSS 0.038205f
C11934 DVSS.n3219 VSS 0.038205f
C11935 DVSS.n3220 VSS 0.038205f
C11936 DVSS.n3221 VSS 0.038205f
C11937 DVSS.n3222 VSS 0.038205f
C11938 DVSS.n3223 VSS 0.035873f
C11939 DVSS.n3224 VSS 0.038205f
C11940 DVSS.n3225 VSS 0.038205f
C11941 DVSS.n3226 VSS 0.038205f
C11942 DVSS.n3227 VSS 0.038205f
C11943 DVSS.n3228 VSS 0.038205f
C11944 DVSS.n3229 VSS 0.049824f
C11945 DVSS.n3231 VSS 0.043865f
C11946 DVSS.n3232 VSS 0.066724f
C11947 DVSS.n3233 VSS 0.043865f
C11948 DVSS.n3234 VSS -0.427302f
C11949 DVSS.n3236 VSS 0.069335f
C11950 DVSS.n3238 VSS 0.066724f
C11951 DVSS.n3239 VSS 0.052308f
C11952 DVSS.n3241 VSS 0.754249f
C11953 DVSS.n3242 VSS 0.052308f
C11954 DVSS.t35 VSS 0.330478f
C11955 DVSS.n3246 VSS 0.635269f
C11956 DVSS.n3247 VSS 0.066724f
C11957 DVSS.n3248 VSS 0.052308f
C11958 DVSS.n3250 VSS 0.754249f
C11959 DVSS.n3251 VSS 0.052308f
C11960 DVSS.n3256 VSS 0.020594f
C11961 DVSS.n3258 VSS 0.010297f
C11962 DVSS.n3259 VSS 0.020594f
C11963 DVSS.n3262 VSS 0.052308f
C11964 DVSS.n3264 VSS 0.066724f
C11965 DVSS.n3265 VSS 0.052308f
C11966 DVSS.t21 VSS 0.330478f
C11967 DVSS.n3266 VSS 0.635269f
C11968 DVSS.n3269 VSS 0.052308f
C11969 DVSS.n3271 VSS 0.066724f
C11970 DVSS.n3272 VSS 0.052308f
C11971 DVSS.n3275 VSS 0.069335f
C11972 DVSS.n3277 VSS 0.066724f
C11973 DVSS.n3279 VSS 0.043865f
C11974 DVSS.n3280 VSS 0.043865f
C11975 DVSS.n3281 VSS 0.065379f
C11976 DVSS.n3282 VSS 0.038205f
C11977 DVSS.n3283 VSS 0.035873f
C11978 DVSS.n3284 VSS -0.427302f
C11979 DVSS.n3285 VSS 0.038205f
C11980 DVSS.n3287 VSS 0.043865f
C11981 DVSS.n3288 VSS 0.066724f
C11982 DVSS.n3289 VSS 0.043865f
C11983 DVSS.n3292 VSS 0.052308f
C11984 DVSS.n3293 VSS 0.754249f
C11985 DVSS.n3295 VSS 0.066724f
C11986 DVSS.n3296 VSS 0.052308f
C11987 DVSS.t19 VSS 0.394423f
C11988 DVSS.n3297 VSS 0.635269f
C11989 DVSS.n3300 VSS 0.052308f
C11990 DVSS.n3301 VSS 0.754249f
C11991 DVSS.n3303 VSS 0.066724f
C11992 DVSS.n3304 VSS 0.052308f
C11993 DVSS.n3307 VSS 0.052308f
C11994 DVSS.n3310 VSS 0.066724f
C11995 DVSS.n3311 VSS 0.74307f
C11996 DVSS.n3312 VSS 0.052308f
C11997 DVSS.n3313 VSS 0.052308f
C11998 DVSS.n3314 VSS 0.066724f
C11999 DVSS.n3315 VSS 0.74307f
C12000 DVSS.n3317 VSS 0.052308f
C12001 DVSS.n3318 VSS 0.052308f
C12002 DVSS.t33 VSS 0.394423f
C12003 DVSS.n3322 VSS 0.635269f
C12004 DVSS.n3323 VSS 0.066724f
C12005 DVSS.n3324 VSS 0.026154f
C12006 DVSS.n3325 VSS 0.082541f
C12007 DVSS.n3326 VSS 0.082541f
C12008 DVSS.n3327 VSS 0.082541f
C12009 DVSS.n3328 VSS 0.072078f
C12010 DVSS.n3329 VSS 0.026154f
C12011 DVSS.n3330 VSS 0.026154f
C12012 DVSS.n3331 VSS 0.041129f
C12013 DVSS.n3332 VSS 0.144737f
C12014 DVSS.n3333 VSS 0.439557f
C12015 DVSS.n3335 VSS 0.052308f
C12016 DVSS.n3338 VSS 0.052308f
C12017 DVSS.n3339 VSS 0.052308f
C12018 DVSS.n3341 VSS 0.052308f
C12019 DVSS.n3343 VSS 0.026154f
C12020 DVSS.n3344 VSS 0.026154f
C12021 DVSS.n3346 VSS 0.186719f
C12022 DVSS.n3347 VSS 0.026154f
C12023 DVSS.n3349 VSS 0.066724f
C12024 DVSS.t2 VSS 0.394423f
C12025 DVSS.n3350 VSS 0.635269f
C12026 DVSS.n3351 VSS 0.026154f
C12027 DVSS.n3353 VSS 0.026154f
C12028 DVSS.n3354 VSS 0.026154f
C12029 DVSS.n3355 VSS 0.026154f
C12030 DVSS.n3356 VSS 0.066724f
C12031 DVSS.n3357 VSS 0.026154f
C12032 DVSS.n3359 VSS 0.066724f
C12033 DVSS.n3361 VSS 0.026154f
C12034 DVSS.n3363 VSS 0.026154f
C12035 DVSS.n3364 VSS 0.026154f
C12036 DVSS.n3365 VSS 0.026154f
C12037 DVSS.n3366 VSS 0.066724f
C12038 DVSS.n3367 VSS 0.026154f
C12039 DVSS.n3369 VSS 0.066724f
C12040 DVSS.n3370 VSS 0.026154f
C12041 DVSS.n3371 VSS 0.082541f
C12042 DVSS.n3372 VSS 0.082541f
C12043 DVSS.n3373 VSS 0.082541f
C12044 DVSS.n3374 VSS 0.072078f
C12045 DVSS.n3375 VSS 0.041129f
C12046 DVSS.n3376 VSS 0.144737f
C12047 DVSS.n3378 VSS 0.082541f
C12048 DVSS.n3379 VSS 0.082541f
C12049 DVSS.n3380 VSS 0.134274f
C12050 DVSS.n3381 VSS 0.052308f
C12051 DVSS.n3382 VSS 0.052308f
C12052 DVSS.n3383 VSS 0.052308f
C12053 DVSS.n3384 VSS 0.026154f
C12054 DVSS.n3385 VSS 0.026154f
C12055 DVSS.n3386 VSS 0.072078f
C12056 DVSS.n3387 VSS 0.026154f
C12057 DVSS.n3388 VSS 0.026154f
C12058 DVSS.n3390 VSS 0.038176f
C12059 DVSS.n3392 VSS 0.052308f
C12060 DVSS.n3393 VSS 0.072078f
C12061 DVSS.n3394 VSS 0.165082f
C12062 DVSS.n3395 VSS 0.165082f
C12063 DVSS.n3396 VSS 0.165082f
C12064 DVSS.n3397 VSS 0.165082f
C12065 DVSS.n3398 VSS 0.165082f
C12066 DVSS.n3399 VSS 0.165082f
C12067 DVSS.n3400 VSS 0.165082f
C12068 DVSS.n3401 VSS 0.082541f
C12069 DVSS.n3402 VSS 0.165082f
C12070 DVSS.n3403 VSS 0.165082f
C12071 DVSS.n3404 VSS 0.165082f
C12072 DVSS.n3405 VSS 0.082541f
C12073 DVSS.n3406 VSS 0.052308f
C12074 DVSS.n3407 VSS 0.052308f
C12075 DVSS.n3408 VSS 0.052308f
C12076 DVSS.n3409 VSS 0.026154f
C12077 DVSS.n3410 VSS 0.026154f
C12078 DVSS.n3411 VSS 0.072078f
C12079 DVSS.n3412 VSS 0.026154f
C12080 DVSS.n3413 VSS 0.026154f
C12081 DVSS.n3415 VSS 0.038176f
C12082 DVSS.n3418 VSS 0.052308f
C12083 DVSS.n3421 VSS 0.052308f
C12084 DVSS.n3423 VSS 0.439557f
C12085 DVSS.n3424 VSS 0.165082f
C12086 DVSS.n3425 VSS 0.165082f
C12087 DVSS.n3426 VSS 0.165082f
C12088 DVSS.n3427 VSS 0.165082f
C12089 DVSS.n3428 VSS 0.165082f
C12090 DVSS.n3429 VSS 0.165082f
C12091 DVSS.n3430 VSS 0.165082f
C12092 DVSS.n3431 VSS 0.165082f
C12093 DVSS.n3432 VSS 0.165082f
C12094 DVSS.n3433 VSS 0.165082f
C12095 DVSS.n3434 VSS 0.165082f
C12096 DVSS.n3435 VSS 0.165082f
C12097 DVSS.n3436 VSS 0.082541f
C12098 DVSS.n3437 VSS 0.165082f
C12099 DVSS.n3438 VSS 0.165082f
C12100 DVSS.n3439 VSS 0.165082f
C12101 DVSS.n3440 VSS 0.082541f
C12102 DVSS.n3441 VSS 0.052308f
C12103 DVSS.n3442 VSS 0.052308f
C12104 DVSS.n3443 VSS 0.052308f
C12105 DVSS.n3444 VSS 0.026154f
C12106 DVSS.n3445 VSS 0.026154f
C12107 DVSS.n3446 VSS 0.072078f
C12108 DVSS.n3447 VSS 0.026154f
C12109 DVSS.n3448 VSS 0.026154f
C12110 DVSS.n3450 VSS 0.038176f
C12111 DVSS.n3453 VSS 0.052308f
C12112 DVSS.n3456 VSS 0.052308f
C12113 DVSS.n3458 VSS 0.165082f
C12114 DVSS.n3459 VSS 0.165082f
C12115 DVSS.n3460 VSS 0.165082f
C12116 DVSS.n3461 VSS 0.165082f
C12117 DVSS.n3462 VSS 0.165082f
C12118 DVSS.n3463 VSS 0.165082f
C12119 DVSS.n3464 VSS 0.165082f
C12120 DVSS.n3465 VSS 0.165082f
C12121 DVSS.n3466 VSS 0.165082f
C12122 DVSS.n3467 VSS 0.165082f
C12123 DVSS.n3468 VSS 0.165082f
C12124 DVSS.n3469 VSS 0.165082f
C12125 DVSS.n3470 VSS 0.082541f
C12126 DVSS.n3471 VSS 0.165082f
C12127 DVSS.n3472 VSS 0.165082f
C12128 DVSS.n3473 VSS 0.165082f
C12129 DVSS.n3474 VSS 0.082541f
C12130 DVSS.n3475 VSS 0.019102f
C12131 DVSS.n3476 VSS 0.019102f
C12132 DVSS.n3478 VSS 0.021932f
C12133 DVSS.n3479 VSS 0.021932f
C12134 DVSS.n3480 VSS 0.072078f
C12135 DVSS.n3481 VSS 0.021932f
C12136 DVSS.n3482 VSS 0.021932f
C12137 DVSS.n3483 VSS 0.019102f
C12138 DVSS.n3484 VSS 0.019102f
C12139 DVSS.n3485 VSS 0.021932f
C12140 DVSS.n3486 VSS 0.038205f
C12141 DVSS.n3487 VSS 0.035873f
C12142 DVSS.n3488 VSS 0.035873f
C12143 DVSS.n3489 VSS 0.019102f
C12144 DVSS.n3490 VSS 0.038205f
C12145 DVSS.n3491 VSS 0.038205f
C12146 DVSS.n3492 VSS 0.038205f
C12147 DVSS.n3493 VSS 0.038205f
C12148 DVSS.n3494 VSS 0.035873f
C12149 DVSS.n3495 VSS 0.038205f
C12150 DVSS.n3496 VSS 0.038205f
C12151 DVSS.n3497 VSS 0.038205f
C12152 DVSS.n3498 VSS 0.038205f
C12153 DVSS.n3499 VSS 0.038205f
C12154 DVSS.t15 VSS 0.330478f
C12155 DVSS.n3500 VSS 0.125906f
C12156 DVSS.n3501 VSS 0.038205f
C12157 DVSS.n3502 VSS 0.038205f
C12158 DVSS.n3503 VSS 0.038205f
C12159 DVSS.n3504 VSS 0.038205f
C12160 DVSS.n3505 VSS 0.035873f
C12161 DVSS.n3506 VSS 0.038205f
C12162 DVSS.n3507 VSS 0.038205f
C12163 DVSS.n3508 VSS 0.038205f
C12164 DVSS.n3509 VSS 0.038205f
C12165 DVSS.n3510 VSS 0.038205f
C12166 DVSS.n3511 VSS 0.035873f
C12167 DVSS.n3512 VSS 0.020694f
C12168 DVSS.n3513 VSS 0.038205f
C12169 DVSS.n3514 VSS 0.038205f
C12170 DVSS.n3515 VSS 0.020694f
C12171 DVSS.n3516 VSS 0.021932f
C12172 DVSS.n3517 VSS 0.021932f
C12173 DVSS.n3518 VSS 0.021932f
C12174 DVSS.n3519 VSS 0.021932f
C12175 DVSS.n3520 VSS 0.021932f
C12176 DVSS.n3522 VSS 0.021932f
C12177 DVSS.n3523 VSS 0.066724f
C12178 DVSS.n3524 VSS 0.026154f
C12179 DVSS.n3526 VSS 0.026154f
C12180 DVSS.n3527 VSS 0.066724f
C12181 DVSS.t1 VSS 0.330478f
C12182 DVSS.n3528 VSS 0.635269f
C12183 DVSS.n3529 VSS 0.026154f
C12184 DVSS.n3531 VSS 0.026154f
C12185 DVSS.n3532 VSS 0.066724f
C12186 DVSS.n3533 VSS 0.010297f
C12187 DVSS.n3534 VSS 0.010297f
C12188 DVSS.n3536 VSS 0.010297f
C12189 DVSS.t8 VSS 0.394423f
C12190 DVSS.n3537 VSS 0.32373f
C12191 DVSS.n3538 VSS 0.2147f
C12192 DVSS.n3539 VSS 0.010297f
C12193 DVSS.n3540 VSS 0.253981f
C12194 DVSS.n3541 VSS 0.09309f
C12195 DVSS.n3542 VSS 0.026154f
C12196 DVSS.n3545 VSS 0.066724f
C12197 DVSS.n3546 VSS 0.026154f
C12198 DVSS.n3547 VSS 0.335771f
C12199 DVSS.n3548 VSS 0.756156f
C12200 DVSS.n3549 VSS 0.242143f
C12201 DVSS.n3550 VSS 0.026154f
C12202 DVSS.n3553 VSS 0.066724f
C12203 DVSS.n3554 VSS 0.026154f
C12204 DVSS.n3555 VSS 0.186719f
C12205 DVSS.n3556 VSS 0.021932f
C12206 DVSS.n3558 VSS 0.396845f
C12207 DVSS.n3559 VSS 0.021932f
C12208 DVSS.n3560 VSS 0.065379f
C12209 DVSS.n3561 VSS 0.049824f
C12210 DVSS.n3562 VSS 0.065379f
C12211 DVSS.n3563 VSS 0.057484f
C12212 DVSS.n3564 VSS 0.021932f
C12213 DVSS.n3566 VSS 0.021932f
C12214 DVSS.n3567 VSS 0.066724f
C12215 DVSS.n3569 VSS 0.740117f
C12216 DVSS.n3571 VSS 0.026154f
C12217 DVSS.n3572 VSS 0.026154f
C12218 DVSS.n3573 VSS 0.066724f
C12219 DVSS.n3575 VSS 0.066724f
C12220 DVSS.n3576 VSS 0.026154f
C12221 DVSS.t24 VSS 0.394423f
C12222 DVSS.n3578 VSS 0.635269f
C12223 DVSS.n3579 VSS 0.740117f
C12224 DVSS.n3581 VSS 0.026154f
C12225 DVSS.n3582 VSS 0.026154f
C12226 DVSS.n3583 VSS 0.066724f
C12227 DVSS.n3585 VSS 0.066724f
C12228 DVSS.n3586 VSS 0.026154f
C12229 DVSS.n3588 VSS 0.026154f
C12230 DVSS.n3590 VSS 0.179185f
C12231 DVSS.n3591 VSS 0.026154f
C12232 DVSS.n3593 VSS 0.331802f
C12233 DVSS.n3594 VSS 0.026154f
C12234 DVSS.n3595 VSS 0.026154f
C12235 DVSS.n3596 VSS 0.066724f
C12236 DVSS.n3597 VSS 0.026154f
C12237 DVSS.n3598 VSS 0.082541f
C12238 DVSS.n3599 VSS 0.082541f
C12239 DVSS.n3600 VSS 0.082541f
C12240 DVSS.n3601 VSS 0.134274f
C12241 DVSS.n3602 VSS 0.052308f
C12242 DVSS.n3603 VSS 0.052308f
C12243 DVSS.n3604 VSS 0.052308f
C12244 DVSS.n3605 VSS 0.165082f
C12245 DVSS.n3606 VSS 0.072078f
C12246 DVSS.n3607 VSS 0.165082f
C12247 DVSS.n3608 VSS 0.165082f
C12248 DVSS.n3609 VSS 0.165082f
C12249 DVSS.n3610 VSS 0.144737f
C12250 DVSS.n3611 VSS 0.165082f
C12251 DVSS.n3612 VSS 0.165082f
C12252 DVSS.n3613 VSS 0.165082f
C12253 DVSS.n3614 VSS 0.082541f
C12254 DVSS.n3615 VSS 0.026154f
C12255 DVSS.n3616 VSS 0.026154f
C12256 DVSS.n3619 VSS 0.052308f
C12257 DVSS.n3620 VSS 0.439768f
C12258 DVSS.n3621 VSS 0.036911f
C12259 DVSS.n3622 VSS 0.026154f
C12260 DVSS.n3623 VSS 0.026154f
C12261 DVSS.n3624 VSS 0.072078f
C12262 DVSS.n3625 VSS 0.082541f
C12263 DVSS.n3626 VSS 0.738852f
C12264 DVSS.n3627 VSS 0.134274f
C12265 DVSS.n3629 VSS 0.052308f
C12266 DVSS.n3630 VSS 0.052308f
C12267 DVSS.n3632 VSS 0.165082f
C12268 DVSS.n3633 VSS 0.165082f
C12269 DVSS.n3634 VSS 0.165082f
C12270 DVSS.n3635 VSS 0.165082f
C12271 DVSS.n3636 VSS 0.165082f
C12272 DVSS.n3637 VSS 0.165082f
C12273 DVSS.n3638 VSS 0.165082f
C12274 DVSS.n3639 VSS 0.165082f
C12275 DVSS.n3640 VSS 0.165082f
C12276 DVSS.n3641 VSS 0.165082f
C12277 DVSS.n3642 VSS 0.165082f
C12278 DVSS.n3643 VSS 0.144737f
C12279 DVSS.n3644 VSS 0.165082f
C12280 DVSS.n3645 VSS 0.165082f
C12281 DVSS.n3646 VSS 0.165082f
C12282 DVSS.n3647 VSS 0.082541f
C12283 DVSS.n3648 VSS 0.026154f
C12284 DVSS.n3649 VSS 0.026154f
C12285 DVSS.n3650 VSS 0.026154f
C12286 DVSS.n3651 VSS 0.026154f
C12287 DVSS.n3656 VSS 0.134274f
C12288 DVSS.n3657 VSS 0.052308f
C12289 DVSS.n3658 VSS 0.052308f
C12290 DVSS.n3659 VSS 0.052308f
C12291 DVSS.n3660 VSS 0.072078f
C12292 DVSS.n3661 VSS 0.052308f
C12293 DVSS.n3662 VSS 0.052308f
C12294 DVSS.n3665 VSS 0.072078f
C12295 DVSS.n3666 VSS 0.082541f
C12296 DVSS.n3667 VSS 0.066724f
C12297 DVSS.n3668 VSS 0.021932f
C12298 DVSS.n3670 VSS 0.056423f
C12299 DVSS.n3671 VSS 0.021932f
C12300 DVSS.n3672 VSS 0.021932f
C12301 DVSS.n3673 VSS 0.066724f
C12302 DVSS.n3674 VSS 0.021932f
C12303 DVSS.n3675 VSS -0.427302f
C12304 DVSS.n3676 VSS 0.021932f
C12305 DVSS.n3677 VSS 0.082541f
C12306 DVSS.n3678 VSS 0.082541f
C12307 DVSS.n3679 VSS 0.111605f
C12308 DVSS.n3680 VSS 0.038382f
C12309 DVSS.n3681 VSS 0.019102f
C12310 DVSS.n3682 VSS 0.019102f
C12311 DVSS.n3683 VSS 0.072078f
C12312 DVSS.n3684 VSS 0.019102f
C12313 DVSS.n3685 VSS 0.019102f
C12314 DVSS.n3686 VSS 0.021932f
C12315 DVSS.n3687 VSS 0.035873f
C12316 DVSS.n3688 VSS 0.019102f
C12317 DVSS.n3690 VSS 0.082541f
C12318 DVSS.n3691 VSS 0.159269f
C12319 DVSS.n3692 VSS 0.021932f
C12320 DVSS.n3693 VSS 0.021932f
C12321 DVSS.n3694 VSS 0.021932f
C12322 DVSS.n3695 VSS 0.019102f
C12323 DVSS.n3696 VSS 0.019102f
C12324 DVSS.n3697 VSS 0.072078f
C12325 DVSS.n3698 VSS 0.019102f
C12326 DVSS.n3699 VSS 0.019102f
C12327 DVSS.n3700 VSS 0.030953f
C12328 DVSS.n3701 VSS 0.021932f
C12329 DVSS.n3702 VSS 0.021932f
C12330 DVSS.n3703 VSS 0.082541f
C12331 DVSS.n3705 VSS 0.066505f
C12332 DVSS.n3706 VSS 0.021932f
C12333 DVSS.n3708 VSS 0.021932f
C12334 DVSS.n3709 VSS 0.066724f
C12335 DVSS.n3710 VSS 0.026154f
C12336 DVSS.n3712 VSS 0.738852f
C12337 DVSS.n3713 VSS 0.026154f
C12338 DVSS.n3714 VSS 0.026154f
C12339 DVSS.n3715 VSS 0.066724f
C12340 DVSS.n3716 VSS 0.242143f
C12341 DVSS.n3717 VSS 0.026154f
C12342 DVSS.n3718 VSS 0.026154f
C12343 DVSS.n3719 VSS 0.082541f
C12344 DVSS.n3720 VSS 0.082541f
C12345 DVSS.n3721 VSS 0.082541f
C12346 DVSS.n3722 VSS 0.147063f
C12347 DVSS.n3723 VSS 0.052308f
C12348 DVSS.n3724 VSS 0.052308f
C12349 DVSS.n3725 VSS 0.052308f
C12350 DVSS.n3726 VSS 0.072078f
C12351 DVSS.n3728 VSS 0.075348f
C12352 DVSS.n3729 VSS 0.075348f
C12353 DVSS.n3730 VSS 0.134247f
C12354 DVSS.n3731 VSS 0.060323f
C12355 DVSS.n3732 VSS 0.052308f
C12356 DVSS.n3733 VSS 0.052308f
C12357 DVSS.n3734 VSS 0.022779f
C12358 DVSS.n3735 VSS 0.065797f
C12359 DVSS.n3736 VSS 0.041129f
C12360 DVSS.n3738 VSS 0.052308f
C12361 DVSS.n3740 VSS 0.052308f
C12362 DVSS.n3742 VSS 0.044082f
C12363 DVSS.n3743 VSS 0.026154f
C12364 DVSS.n3744 VSS 0.026154f
C12365 DVSS.n3747 VSS 0.150696f
C12366 DVSS.n3748 VSS 0.150696f
C12367 DVSS.n3749 VSS 0.150696f
C12368 DVSS.n3750 VSS 0.150696f
C12369 DVSS.n3751 VSS 0.150696f
C12370 DVSS.n3752 VSS 0.150696f
C12371 DVSS.n3753 VSS 0.150696f
C12372 DVSS.n3754 VSS 0.150696f
C12373 DVSS.n3755 VSS 0.150696f
C12374 DVSS.n3756 VSS 0.150696f
C12375 DVSS.n3757 VSS 0.150696f
C12376 DVSS.n3758 VSS 0.150696f
C12377 DVSS.n3759 VSS 0.150696f
C12378 DVSS.n3760 VSS 0.150696f
C12379 DVSS.n3761 VSS 0.150696f
C12380 DVSS.n3762 VSS 0.150696f
C12381 DVSS.n3763 VSS 0.150696f
C12382 DVSS.n3764 VSS 0.150696f
C12383 DVSS.n3765 VSS 0.150696f
C12384 DVSS.n3766 VSS 0.150696f
C12385 DVSS.n3767 VSS 0.150696f
C12386 DVSS.n3768 VSS 0.150696f
C12387 DVSS.n3769 VSS 0.150696f
C12388 DVSS.n3770 VSS 0.050586f
C12389 DVSS.n3771 VSS 0.019102f
C12390 DVSS.n3772 VSS 0.019102f
C12391 DVSS.n3773 VSS 0.03396f
C12392 DVSS.n3774 VSS 0.019102f
C12393 DVSS.n3775 VSS 0.065797f
C12394 DVSS.n3776 VSS 0.03449f
C12395 DVSS.n3777 VSS 0.019102f
C12396 DVSS.n3778 VSS 0.019102f
C12397 DVSS.n3779 VSS 0.036967f
C12398 DVSS.n3780 VSS 0.021932f
C12399 DVSS.n3783 VSS 0.075348f
C12400 DVSS.n3786 VSS 0.032106f
C12401 DVSS.n3788 VSS 0.032106f
C12402 DVSS.n3790 VSS 0.032106f
C12403 DVSS.n3792 VSS 0.026154f
C12404 DVSS.n3793 VSS 0.044082f
C12405 DVSS.n3794 VSS 0.032106f
C12406 DVSS.n3795 VSS 0.032106f
C12407 DVSS.n3796 VSS 0.022779f
C12408 DVSS.n3798 VSS 0.120696f
C12409 DVSS.n3799 VSS 0.075348f
C12410 DVSS.n3800 VSS 0.075348f
C12411 DVSS.n3801 VSS 0.075348f
C12412 DVSS.n3802 VSS 0.134247f
C12413 DVSS.n3804 VSS 0.060323f
C12414 DVSS.n3805 VSS 0.439768f
C12415 DVSS.n3806 VSS 0.052308f
C12416 DVSS.n3807 VSS 0.052308f
C12417 DVSS.n3808 VSS 0.150696f
C12418 DVSS.n3809 VSS 0.150696f
C12419 DVSS.n3810 VSS 0.150696f
C12420 DVSS.n3811 VSS 0.120451f
C12421 DVSS.n3812 VSS 0.150696f
C12422 DVSS.n3813 VSS 0.150696f
C12423 DVSS.n3814 VSS 0.150696f
C12424 DVSS.n3815 VSS 0.075348f
C12425 DVSS.n3816 VSS 0.060323f
C12426 DVSS.n3817 VSS 0.439768f
C12427 DVSS.n3818 VSS 0.022779f
C12428 DVSS.n3819 VSS 0.041129f
C12429 DVSS.n3823 VSS 0.044082f
C12430 DVSS.n3824 VSS 0.026154f
C12431 DVSS.n3825 VSS 0.075348f
C12432 DVSS.n3826 VSS 0.026154f
C12433 DVSS.n3827 VSS 0.150696f
C12434 DVSS.n3828 VSS 0.150696f
C12435 DVSS.n3829 VSS 0.150696f
C12436 DVSS.n3830 VSS 0.120451f
C12437 DVSS.n3831 VSS 0.150696f
C12438 DVSS.n3832 VSS 0.558604f
C12439 DVSS.n3833 VSS 0.150696f
C12440 DVSS.n3834 VSS 0.075348f
C12441 DVSS.n3835 VSS 0.060323f
C12442 DVSS.n3837 VSS 0.082541f
C12443 DVSS.n3838 VSS 0.082541f
C12444 DVSS.n3839 VSS 0.3147f
C12445 DVSS.n3840 VSS 0.022779f
C12446 DVSS.n3841 VSS 0.022779f
C12447 DVSS.n3842 VSS 0.052308f
C12448 DVSS.n3843 VSS 0.052308f
C12449 DVSS.n3844 VSS 0.052308f
C12450 DVSS.n3845 VSS 0.072078f
C12451 DVSS.n3847 VSS 0.052308f
C12452 DVSS.n3849 VSS 0.052308f
C12453 DVSS.n3851 VSS 0.04366f
C12454 DVSS.n3852 VSS 0.022779f
C12455 DVSS.n3853 VSS 0.026154f
C12456 DVSS.n3856 VSS 0.082541f
C12457 DVSS.n3857 VSS 0.058114f
C12458 DVSS.t36 VSS 0.394423f
C12459 DVSS.n3858 VSS 0.026154f
C12460 DVSS.n3860 VSS 0.32751f
C12461 DVSS.n3861 VSS 0.026154f
C12462 DVSS.n3862 VSS 0.026154f
C12463 DVSS.n3863 VSS 0.066724f
C12464 DVSS.n3864 VSS 0.026154f
C12465 DVSS.n3866 VSS 0.066724f
C12466 DVSS.n3868 VSS 0.026154f
C12467 DVSS.n3870 VSS 0.066724f
C12468 DVSS.n3871 VSS 0.286603f
C12469 DVSS.n3872 VSS 0.010297f
C12470 DVSS.n3874 VSS 0.010297f
C12471 DVSS.n3875 VSS 0.2147f
C12472 DVSS.n3876 VSS 0.010297f
C12473 DVSS.n3877 VSS 0.253981f
C12474 DVSS.n3878 VSS 0.09309f
C12475 DVSS.n3879 VSS 0.026154f
C12476 DVSS.n3880 VSS 0.066724f
C12477 DVSS.t23 VSS 0.330478f
C12478 DVSS.n3882 VSS 0.635269f
C12479 DVSS.n3883 VSS 0.756156f
C12480 DVSS.n3885 VSS 0.026154f
C12481 DVSS.n3886 VSS 0.026154f
C12482 DVSS.n3887 VSS 0.082541f
C12483 DVSS.n3888 VSS 0.082541f
C12484 DVSS.n3889 VSS 0.082541f
C12485 DVSS.n3890 VSS 0.147063f
C12486 DVSS.n3891 VSS 0.052308f
C12487 DVSS.n3892 VSS 0.052308f
C12488 DVSS.n3893 VSS 0.052308f
C12489 DVSS.n3894 VSS 0.026154f
C12490 DVSS.n3895 VSS 0.165082f
C12491 DVSS.n3896 VSS 0.072078f
C12492 DVSS.n3897 VSS 0.165082f
C12493 DVSS.n3898 VSS 0.165082f
C12494 DVSS.n3899 VSS 0.165082f
C12495 DVSS.n3900 VSS 0.165082f
C12496 DVSS.n3901 VSS 0.165082f
C12497 DVSS.n3902 VSS 0.165082f
C12498 DVSS.n3903 VSS 0.165082f
C12499 DVSS.n3904 VSS 0.165082f
C12500 DVSS.n3905 VSS 0.165082f
C12501 DVSS.n3906 VSS 0.165082f
C12502 DVSS.n3907 VSS 0.165082f
C12503 DVSS.n3908 VSS 0.165082f
C12504 DVSS.n3909 VSS 0.165082f
C12505 DVSS.n3910 VSS 0.165082f
C12506 DVSS.n3911 VSS 0.165082f
C12507 DVSS.n3912 VSS 0.165082f
C12508 DVSS.n3913 VSS 0.165082f
C12509 DVSS.n3914 VSS 0.165082f
C12510 DVSS.n3915 VSS 0.165082f
C12511 DVSS.n3916 VSS 0.165082f
C12512 DVSS.n3917 VSS 0.165082f
C12513 DVSS.n3918 VSS 0.165082f
C12514 DVSS.n3919 VSS 0.165082f
C12515 DVSS.n3920 VSS 0.165082f
C12516 DVSS.n3921 VSS 0.165082f
C12517 DVSS.n3922 VSS 0.165082f
C12518 DVSS.n3923 VSS 0.165082f
C12519 DVSS.n3924 VSS 0.165082f
C12520 DVSS.n3925 VSS 0.165082f
C12521 DVSS.n3926 VSS 0.165082f
C12522 DVSS.n3927 VSS 0.165082f
C12523 DVSS.n3928 VSS 0.165082f
C12524 DVSS.n3929 VSS 0.165082f
C12525 DVSS.n3930 VSS 0.165082f
C12526 DVSS.n3931 VSS 0.052308f
C12527 DVSS.n3932 VSS 0.052308f
C12528 DVSS.n3933 VSS 0.052308f
C12529 DVSS.n3934 VSS 0.026154f
C12530 DVSS.n3935 VSS 0.026154f
C12531 DVSS.n3936 VSS 0.072078f
C12532 DVSS.n3937 VSS 0.026154f
C12533 DVSS.n3938 VSS 0.026154f
C12534 DVSS.n3939 VSS 0.038176f
C12535 DVSS.n3940 VSS 0.052308f
C12536 DVSS.n3941 VSS 0.052308f
C12537 DVSS.n3946 VSS 0.082541f
C12538 DVSS.n3947 VSS 0.072078f
C12539 DVSS.n3950 VSS 0.082541f
C12540 DVSS.n3951 VSS 0.165082f
C12541 DVSS.n3952 VSS 0.165082f
C12542 DVSS.n3953 VSS 0.165082f
C12543 DVSS.n3954 VSS 0.165082f
C12544 DVSS.n3955 VSS 0.165082f
C12545 DVSS.n3956 VSS 0.131949f
C12546 DVSS.n3957 VSS 0.165082f
C12547 DVSS.n3958 VSS 0.165082f
C12548 DVSS.n3959 VSS 0.165082f
C12549 DVSS.n3960 VSS 0.165082f
C12550 DVSS.n3961 VSS 0.165082f
C12551 DVSS.n3962 VSS 0.165082f
C12552 DVSS.n3963 VSS 0.165082f
C12553 DVSS.n3964 VSS 0.165082f
C12554 DVSS.n3965 VSS 0.159269f
C12555 DVSS.n3966 VSS 0.165082f
C12556 DVSS.n3967 VSS 0.165082f
C12557 DVSS.n3968 VSS 0.165082f
C12558 DVSS.n3969 VSS 0.082541f
C12559 DVSS.n3970 VSS 0.021932f
C12560 DVSS.n3971 VSS 0.019102f
C12561 DVSS.n3972 VSS 0.019102f
C12562 DVSS.n3974 VSS 0.021932f
C12563 DVSS.n3975 VSS 0.021932f
C12564 DVSS.n3976 VSS 0.072078f
C12565 DVSS.n3977 VSS 0.021932f
C12566 DVSS.n3978 VSS 0.021932f
C12567 DVSS.n3979 VSS 0.019102f
C12568 DVSS.n3980 VSS 0.021932f
C12569 DVSS.n3981 VSS 0.021932f
C12570 DVSS.n3982 VSS 0.03732f
C12571 DVSS.n3983 VSS 0.021932f
C12572 DVSS.n3984 VSS 0.021932f
C12573 DVSS.n3985 VSS 0.021932f
C12574 DVSS.n3986 VSS 0.021932f
C12575 DVSS.n3987 VSS 0.035873f
C12576 DVSS.n3988 VSS 0.035873f
C12577 DVSS.n3989 VSS 0.021932f
C12578 DVSS.n3990 VSS 0.035873f
C12579 DVSS.n3991 VSS 0.031887f
C12580 DVSS.n3992 VSS 0.021932f
C12581 DVSS.n3993 VSS 0.03732f
C12582 DVSS.n3994 VSS 0.111605f
C12583 DVSS.n3995 VSS 0.165082f
C12584 DVSS.n3996 VSS 0.165082f
C12585 DVSS.n3997 VSS 0.10928f
C12586 DVSS.n3998 VSS 0.066724f
C12587 DVSS.n3999 VSS 0.740117f
C12588 DVSS.n4001 VSS 0.026154f
C12589 DVSS.n4002 VSS 0.026154f
C12590 DVSS.n4003 VSS 0.066724f
C12591 DVSS.n4004 VSS 0.242143f
C12592 DVSS.n4005 VSS 0.026154f
C12593 DVSS.n4008 VSS 0.066724f
C12594 DVSS.n4009 VSS 0.026154f
C12595 DVSS.n4010 VSS 0.186719f
C12596 DVSS.n4011 VSS 0.038205f
C12597 DVSS.n4012 VSS 0.035873f
C12598 DVSS.n4013 VSS 0.038205f
C12599 DVSS.n4014 VSS 0.035873f
C12600 DVSS.n4015 VSS 0.038205f
C12601 DVSS.n4016 VSS 0.035873f
C12602 DVSS.n4017 VSS 0.038205f
C12603 DVSS.n4018 VSS 0.035873f
C12604 DVSS.n4019 VSS 0.038205f
C12605 DVSS.n4020 VSS 0.035873f
C12606 DVSS.n4021 VSS 0.038205f
C12607 DVSS.n4022 VSS 0.038205f
C12608 DVSS.t10 VSS 0.330478f
C12609 DVSS.n4023 VSS 0.125906f
C12610 DVSS.n4024 VSS 0.038205f
C12611 DVSS.n4025 VSS 0.035873f
C12612 DVSS.n4026 VSS 0.038205f
C12613 DVSS.n4027 VSS 0.035873f
C12614 DVSS.n4028 VSS 0.038205f
C12615 DVSS.n4029 VSS 0.035873f
C12616 DVSS.n4030 VSS 0.038205f
C12617 DVSS.n4031 VSS 0.035873f
C12618 DVSS.n4032 VSS 0.038205f
C12619 DVSS.n4033 VSS 0.035873f
C12620 DVSS.n4034 VSS 0.038205f
C12621 DVSS.n4035 VSS 0.035873f
C12622 DVSS.n4036 VSS 0.066505f
C12623 DVSS.n4037 VSS 0.031887f
C12624 DVSS.n4038 VSS 0.038205f
C12625 DVSS.n4039 VSS 0.035873f
C12626 DVSS.n4040 VSS 0.038205f
C12627 DVSS.n4041 VSS 0.038205f
C12628 DVSS.n4042 VSS 0.038205f
C12629 DVSS.n4043 VSS 0.035873f
C12630 DVSS.n4044 VSS 0.038205f
C12631 DVSS.n4045 VSS 0.038205f
C12632 DVSS.n4046 VSS 0.038205f
C12633 DVSS.n4047 VSS 0.035873f
C12634 DVSS.n4048 VSS 0.038205f
C12635 DVSS.n4049 VSS 0.038205f
C12636 DVSS.n4050 VSS 0.038205f
C12637 DVSS.n4051 VSS 0.035873f
C12638 DVSS.n4052 VSS 0.038205f
C12639 DVSS.n4053 VSS 0.038205f
C12640 DVSS.n4054 VSS 0.038205f
C12641 DVSS.n4055 VSS 0.035873f
C12642 DVSS.n4056 VSS 0.038205f
C12643 DVSS.n4057 VSS 0.038205f
C12644 DVSS.n4058 VSS 0.038205f
C12645 DVSS.n4059 VSS 0.035873f
C12646 DVSS.n4060 VSS 0.038205f
C12647 DVSS.n4061 VSS 0.038205f
C12648 DVSS.n4062 VSS 0.038205f
C12649 DVSS.n4063 VSS 0.026905f
C12650 DVSS.n4064 VSS 0.038205f
C12651 DVSS.n4065 VSS 0.038205f
C12652 DVSS.n4066 VSS 0.026905f
C12653 DVSS.n4067 VSS 0.020096f
C12654 DVSS.n4068 VSS 0.038205f
C12655 DVSS.n4069 VSS 0.038205f
C12656 DVSS.n4070 VSS 0.033714f
C12657 DVSS.n4071 VSS 0.038205f
C12658 DVSS.n4072 VSS 0.038205f
C12659 DVSS.n4073 VSS 0.038205f
C12660 DVSS.n4074 VSS 0.035873f
C12661 DVSS.n4075 VSS 0.038205f
C12662 DVSS.n4076 VSS 0.038205f
C12663 DVSS.n4077 VSS 0.038205f
C12664 DVSS.n4078 VSS 0.035873f
C12665 DVSS.n4079 VSS 0.038205f
C12666 DVSS.n4080 VSS 0.038205f
C12667 DVSS.n4081 VSS 0.038205f
C12668 DVSS.n4082 VSS 0.035873f
C12669 DVSS.n4083 VSS 0.038205f
C12670 DVSS.n4084 VSS 0.038205f
C12671 DVSS.n4085 VSS 0.038205f
C12672 DVSS.n4086 VSS 0.035873f
C12673 DVSS.n4087 VSS 0.038205f
C12674 DVSS.n4088 VSS 0.038205f
C12675 DVSS.n4089 VSS 0.066505f
C12676 DVSS.n4090 VSS 0.038205f
C12677 DVSS.n4091 VSS 0.035873f
C12678 DVSS.n4092 VSS 0.038205f
C12679 DVSS.n4093 VSS 0.066505f
C12680 DVSS.n4094 VSS 0.057484f
C12681 DVSS.n4096 VSS 0.021932f
C12682 DVSS.n4097 VSS 0.021932f
C12683 DVSS.n4098 VSS 0.021932f
C12684 DVSS.n4099 VSS 0.396845f
C12685 DVSS.n4101 VSS 0.021932f
C12686 DVSS.n4102 VSS 0.032014f
C12687 DVSS.n4103 VSS 0.082541f
C12688 DVSS.n4104 VSS 0.019102f
C12689 DVSS.n4105 VSS 0.082541f
C12690 DVSS.n4106 VSS 0.072078f
C12691 DVSS.n4107 VSS 0.165082f
C12692 DVSS.n4108 VSS 0.165082f
C12693 DVSS.n4109 VSS 0.165082f
C12694 DVSS.n4110 VSS 0.165082f
C12695 DVSS.n4111 VSS 0.165082f
C12696 DVSS.n4112 VSS 0.165082f
C12697 DVSS.n4113 VSS 0.165082f
C12698 DVSS.n4114 VSS 0.165082f
C12699 DVSS.n4115 VSS 0.165082f
C12700 DVSS.n4116 VSS 0.165082f
C12701 DVSS.n4117 VSS 0.165082f
C12702 DVSS.n4118 VSS 0.165082f
C12703 DVSS.n4119 VSS 0.165082f
C12704 DVSS.n4120 VSS 0.165082f
C12705 DVSS.n4121 VSS 0.165082f
C12706 DVSS.n4122 VSS 0.165082f
C12707 DVSS.n4123 VSS 0.165082f
C12708 DVSS.n4124 VSS 0.165082f
C12709 DVSS.n4125 VSS 0.165082f
C12710 DVSS.n4126 VSS 0.165082f
C12711 DVSS.n4127 VSS 0.165082f
C12712 DVSS.n4128 VSS 0.165082f
C12713 DVSS.n4129 VSS 0.165082f
C12714 DVSS.n4130 VSS 0.165082f
C12715 DVSS.n4131 VSS 0.165082f
C12716 DVSS.n4132 VSS 0.165082f
C12717 DVSS.n4133 VSS 0.165082f
C12718 DVSS.n4134 VSS 0.165082f
C12719 DVSS.n4135 VSS 0.165082f
C12720 DVSS.n4136 VSS 0.072078f
C12721 DVSS.n4137 VSS 0.082541f
C12722 DVSS.n4138 VSS 0.439557f
C12723 DVSS.n4139 VSS 0.082541f
C12724 DVSS.n4140 VSS 0.147063f
C12725 DVSS.n4141 VSS 0.165082f
C12726 DVSS.n4142 VSS 0.165082f
C12727 DVSS.n4143 VSS 0.165082f
C12728 DVSS.n4144 VSS 0.165082f
C12729 DVSS.n4145 VSS 0.165082f
C12730 DVSS.n4146 VSS 0.165082f
C12731 DVSS.n4147 VSS 0.165082f
C12732 DVSS.n4148 VSS 0.165082f
C12733 DVSS.n4149 VSS 0.165082f
C12734 DVSS.n4150 VSS 0.165082f
C12735 DVSS.n4151 VSS 0.165082f
C12736 DVSS.n4152 VSS 0.165082f
C12737 DVSS.n4153 VSS 0.165082f
C12738 DVSS.n4154 VSS 0.165082f
C12739 DVSS.n4155 VSS 0.165082f
C12740 DVSS.n4156 VSS 0.165082f
C12741 DVSS.n4157 VSS 0.165082f
C12742 DVSS.n4158 VSS 0.165082f
C12743 DVSS.n4159 VSS 0.165082f
C12744 DVSS.n4160 VSS 0.165082f
C12745 DVSS.n4161 VSS 0.165082f
C12746 DVSS.n4162 VSS 0.165082f
C12747 DVSS.n4163 VSS 0.165082f
C12748 DVSS.n4164 VSS 0.131949f
C12749 DVSS.n4165 VSS 0.165082f
C12750 DVSS.n4166 VSS 0.072078f
C12751 DVSS.n4167 VSS 0.165082f
C12752 DVSS.n4168 VSS 0.165082f
C12753 DVSS.n4169 VSS 0.165082f
C12754 DVSS.n4170 VSS 0.165082f
C12755 DVSS.n4171 VSS 0.165082f
C12756 DVSS.n4172 VSS 0.072078f
C12757 DVSS.n4174 VSS 0.026154f
C12758 DVSS.n4175 VSS 0.026154f
C12759 DVSS.n4177 VSS 0.038176f
C12760 DVSS.n4180 VSS 0.052308f
C12761 DVSS.n4183 VSS 0.052308f
C12762 DVSS.n4185 VSS 0.439557f
C12763 DVSS.n4186 VSS 0.082541f
C12764 DVSS.n4187 VSS 0.026154f
C12765 DVSS.n4188 VSS 0.026154f
C12766 DVSS.n4189 VSS 0.335771f
C12767 DVSS.n4190 VSS 0.740117f
C12768 DVSS.n4191 VSS 0.738852f
C12769 DVSS.n4192 VSS 0.026154f
C12770 DVSS.n4193 VSS 0.026154f
C12771 DVSS.n4194 VSS 0.066724f
C12772 DVSS.n4195 VSS 0.026154f
C12773 DVSS.n4197 VSS 0.066724f
C12774 DVSS.n4198 VSS 0.026154f
C12775 DVSS.n4199 VSS 0.082541f
C12776 DVSS.n4200 VSS 0.082541f
C12777 DVSS.n4201 VSS 0.082541f
C12778 DVSS.n4202 VSS 0.147063f
C12779 DVSS.n4203 VSS 0.052308f
C12780 DVSS.n4204 VSS 0.052308f
C12781 DVSS.n4205 VSS 0.052308f
C12782 DVSS.n4206 VSS 0.165082f
C12783 DVSS.n4207 VSS 0.072078f
C12784 DVSS.n4208 VSS 0.165082f
C12785 DVSS.n4209 VSS 0.165082f
C12786 DVSS.n4210 VSS 0.165082f
C12787 DVSS.n4211 VSS 0.131949f
C12788 DVSS.n4212 VSS 0.165082f
C12789 DVSS.n4213 VSS 0.165082f
C12790 DVSS.n4214 VSS 0.165082f
C12791 DVSS.n4215 VSS 0.082541f
C12792 DVSS.n4216 VSS 0.026154f
C12793 DVSS.n4217 VSS 0.439768f
C12794 DVSS.n4221 VSS 0.026154f
C12795 DVSS.n4222 VSS 0.072078f
C12796 DVSS.n4223 VSS 0.082541f
C12797 DVSS.n4224 VSS 0.147063f
C12798 DVSS.n4225 VSS 0.052308f
C12799 DVSS.n4226 VSS 0.052308f
C12800 DVSS.n4228 VSS 0.052308f
C12801 DVSS.n4229 VSS 0.165082f
C12802 DVSS.n4230 VSS 0.165082f
C12803 DVSS.n4231 VSS 0.165082f
C12804 DVSS.n4232 VSS 0.131949f
C12805 DVSS.n4233 VSS 0.165082f
C12806 DVSS.n4234 VSS 0.611712f
C12807 DVSS.n4235 VSS 0.165082f
C12808 DVSS.n4236 VSS 0.072078f
C12809 DVSS.n4237 VSS 0.165082f
C12810 DVSS.n4238 VSS 0.072078f
C12811 DVSS.n4239 VSS 0.165082f
C12812 DVSS.n4240 VSS 0.165082f
C12813 DVSS.n4241 VSS 0.165082f
C12814 DVSS.n4242 VSS 0.165082f
C12815 DVSS.n4243 VSS 0.165082f
C12816 DVSS.n4244 VSS 0.165082f
C12817 DVSS.n4245 VSS 0.165082f
C12818 DVSS.n4246 VSS 0.165082f
C12819 DVSS.n4247 VSS 0.165082f
C12820 DVSS.n4248 VSS 0.165082f
C12821 DVSS.n4249 VSS 0.165082f
C12822 DVSS.n4250 VSS 0.165082f
C12823 DVSS.n4251 VSS 0.165082f
C12824 DVSS.n4252 VSS 0.072078f
C12825 DVSS.n4254 VSS 0.052308f
C12826 DVSS.n4256 VSS 0.052308f
C12827 DVSS.n4257 VSS 0.036911f
C12828 DVSS.n4258 VSS 0.082541f
C12829 DVSS.n4259 VSS 0.026154f
C12830 DVSS.n4260 VSS 0.082541f
C12831 DVSS.n4261 VSS 0.072078f
C12832 DVSS.n4262 VSS 0.165082f
C12833 DVSS.n4263 VSS 0.165082f
C12834 DVSS.n4264 VSS 0.165082f
C12835 DVSS.n4265 VSS 0.165082f
C12836 DVSS.n4266 VSS 0.165082f
C12837 DVSS.n4267 VSS 0.165082f
C12838 DVSS.n4268 VSS 0.165082f
C12839 DVSS.n4269 VSS 0.165082f
C12840 DVSS.n4270 VSS 0.165082f
C12841 DVSS.n4271 VSS 0.165082f
C12842 DVSS.n4272 VSS 0.165082f
C12843 DVSS.n4273 VSS 0.165082f
C12844 DVSS.n4274 VSS 0.165082f
C12845 DVSS.n4275 VSS 0.165082f
C12846 DVSS.n4276 VSS 0.165082f
C12847 DVSS.n4277 VSS 0.165082f
C12848 DVSS.n4278 VSS 0.165082f
C12849 DVSS.n4279 VSS 0.165082f
C12850 DVSS.n4280 VSS 0.165082f
C12851 DVSS.n4281 VSS 0.165082f
C12852 DVSS.n4282 VSS 0.165082f
C12853 DVSS.n4283 VSS 0.165082f
C12854 DVSS.n4284 VSS 0.165082f
C12855 DVSS.n4285 VSS 0.165082f
C12856 DVSS.n4286 VSS 0.165082f
C12857 DVSS.n4287 VSS 0.072078f
C12858 DVSS.n4288 VSS 0.165082f
C12859 DVSS.n4289 VSS 0.165082f
C12860 DVSS.n4290 VSS 0.165082f
C12861 DVSS.n4291 VSS 0.165082f
C12862 DVSS.n4292 VSS 0.165082f
C12863 DVSS.n4293 VSS 0.165082f
C12864 DVSS.n4294 VSS 0.165082f
C12865 DVSS.n4295 VSS 0.165082f
C12866 DVSS.n4296 VSS 0.165082f
C12867 DVSS.n4297 VSS 0.165082f
C12868 DVSS.n4298 VSS 0.165082f
C12869 DVSS.n4299 VSS 0.165082f
C12870 DVSS.n4300 VSS 0.165082f
C12871 DVSS.n4301 VSS 0.165082f
C12872 DVSS.n4302 VSS 0.10928f
C12873 DVSS.n4303 VSS 0.165082f
C12874 DVSS.n4304 VSS 0.165082f
C12875 DVSS.n4305 VSS 0.165082f
C12876 DVSS.n4306 VSS 0.165082f
C12877 DVSS.n4307 VSS 0.165082f
C12878 DVSS.n4308 VSS 0.156944f
C12879 DVSS.n4309 VSS 0.165082f
C12880 DVSS.n4310 VSS 0.165082f
C12881 DVSS.n4311 VSS 0.165082f
C12882 DVSS.n4312 VSS 0.165082f
C12883 DVSS.n4313 VSS 0.165082f
C12884 DVSS.n4314 VSS 0.165082f
C12885 DVSS.n4315 VSS 0.165082f
C12886 DVSS.n4316 VSS 0.165082f
C12887 DVSS.n4317 VSS 0.165082f
C12888 DVSS.n4318 VSS 0.165082f
C12889 DVSS.n4319 VSS 0.165082f
C12890 DVSS.n4320 VSS 0.165082f
C12891 DVSS.n4321 VSS 0.165082f
C12892 DVSS.n4322 VSS 0.165082f
C12893 DVSS.n4323 VSS 0.165082f
C12894 DVSS.n4324 VSS 0.165082f
C12895 DVSS.n4325 VSS 0.165082f
C12896 DVSS.n4326 VSS 0.165082f
C12897 DVSS.n4327 VSS 0.165082f
C12898 DVSS.n4328 VSS 0.165082f
C12899 DVSS.n4329 VSS 0.165082f
C12900 DVSS.n4330 VSS 0.165082f
C12901 DVSS.n4331 VSS 0.165082f
C12902 DVSS.n4332 VSS 0.165082f
C12903 DVSS.n4333 VSS 0.165082f
C12904 DVSS.n4334 VSS 0.165082f
C12905 DVSS.n4335 VSS 0.165082f
C12906 DVSS.n4336 VSS 0.165082f
C12907 DVSS.n4337 VSS 0.165082f
C12908 DVSS.n4338 VSS 0.165082f
C12909 DVSS.n4339 VSS 0.165082f
C12910 DVSS.n4340 VSS 0.165082f
C12911 DVSS.n4341 VSS 0.165082f
C12912 DVSS.n4342 VSS 0.165082f
C12913 DVSS.n4343 VSS 0.165082f
C12914 DVSS.n4344 VSS 0.165082f
C12915 DVSS.n4345 VSS 0.165082f
C12916 DVSS.n4346 VSS 0.072078f
C12917 DVSS.n4347 VSS 0.165082f
C12918 DVSS.n4348 VSS 0.165082f
C12919 DVSS.n4349 VSS 0.165082f
C12920 DVSS.n4350 VSS 0.165082f
C12921 DVSS.n4351 VSS 0.165082f
C12922 DVSS.n4352 VSS 0.165082f
C12923 DVSS.n4353 VSS 0.072078f
C12924 DVSS.n4354 VSS 0.165082f
C12925 DVSS.n4355 VSS 0.165082f
C12926 DVSS.n4356 VSS 0.165082f
C12927 DVSS.n4357 VSS 0.165082f
C12928 DVSS.n4358 VSS 0.165082f
C12929 DVSS.n4359 VSS 0.165082f
C12930 DVSS.n4360 VSS 0.165082f
C12931 DVSS.n4361 VSS 0.165082f
C12932 DVSS.n4362 VSS 0.165082f
C12933 DVSS.n4363 VSS 0.165082f
C12934 DVSS.n4364 VSS 0.165082f
C12935 DVSS.n4365 VSS 0.165082f
C12936 DVSS.n4366 VSS 0.165082f
C12937 DVSS.n4367 VSS 0.165082f
C12938 DVSS.n4368 VSS 0.165082f
C12939 DVSS.n4369 VSS 0.165082f
C12940 DVSS.n4370 VSS 0.165082f
C12941 DVSS.n4371 VSS 0.165082f
C12942 DVSS.n4372 VSS 0.165082f
C12943 DVSS.n4373 VSS 0.165082f
C12944 DVSS.n4374 VSS 0.165082f
C12945 DVSS.n4375 VSS 0.165082f
C12946 DVSS.n4376 VSS 0.165082f
C12947 DVSS.n4377 VSS 0.165082f
C12948 DVSS.n4378 VSS 0.165082f
C12949 DVSS.n4379 VSS 0.131949f
C12950 DVSS.n4380 VSS 0.165082f
C12951 DVSS.n4381 VSS 0.165082f
C12952 DVSS.n4382 VSS 0.165082f
C12953 DVSS.n4383 VSS 0.165082f
C12954 DVSS.n4384 VSS 0.072078f
C12955 DVSS.n4385 VSS 0.165082f
C12956 DVSS.n4386 VSS 0.165082f
C12957 DVSS.n4387 VSS 0.165082f
C12958 DVSS.n4388 VSS 0.165082f
C12959 DVSS.n4389 VSS 0.165082f
C12960 DVSS.n4390 VSS 0.165082f
C12961 DVSS.n4391 VSS 0.165082f
C12962 DVSS.n4392 VSS 0.165082f
C12963 DVSS.n4393 VSS 0.165082f
C12964 DVSS.n4394 VSS 0.165082f
C12965 DVSS.n4395 VSS 0.165082f
C12966 DVSS.n4396 VSS 0.165082f
C12967 DVSS.n4397 VSS 0.165082f
C12968 DVSS.n4398 VSS 0.165082f
C12969 DVSS.n4399 VSS 0.165082f
C12970 DVSS.n4400 VSS 0.165082f
C12971 DVSS.n4401 VSS 0.165082f
C12972 DVSS.n4402 VSS 0.165082f
C12973 DVSS.n4403 VSS 0.165082f
C12974 DVSS.n4404 VSS 0.165082f
C12975 DVSS.n4405 VSS 0.165082f
C12976 DVSS.n4406 VSS 0.165082f
C12977 DVSS.n4407 VSS 0.165082f
C12978 DVSS.n4408 VSS 0.165082f
C12979 DVSS.n4409 VSS 0.165082f
C12980 DVSS.n4410 VSS 0.131949f
C12981 DVSS.n4411 VSS 0.165082f
C12982 DVSS.n4412 VSS 0.072078f
C12983 DVSS.n4413 VSS 0.165082f
C12984 DVSS.n4414 VSS 0.165082f
C12985 DVSS.n4415 VSS 0.165082f
C12986 DVSS.n4416 VSS 0.165082f
C12987 DVSS.n4417 VSS 0.165082f
C12988 DVSS.n4418 VSS 0.072078f
C12989 DVSS.n4420 VSS 0.439768f
C12990 DVSS.n4423 VSS 0.052308f
C12991 DVSS.n4426 VSS 0.052308f
C12992 DVSS.n4428 VSS 0.036911f
C12993 DVSS.n4429 VSS 0.082541f
C12994 DVSS.n4430 VSS 0.026154f
C12995 DVSS.n4431 VSS 0.026154f
C12996 DVSS.t28 VSS 0.330478f
C12997 DVSS.n4433 VSS 0.635269f
C12998 DVSS.n4434 VSS 0.756156f
C12999 DVSS.n4435 VSS 0.335771f
C13000 DVSS.n4436 VSS 0.026154f
C13001 DVSS.n4437 VSS 0.09309f
C13002 DVSS.n4438 VSS 0.179185f
C13003 DVSS.n4439 VSS 0.026154f
C13004 DVSS.n4440 VSS 0.222771f
C13005 DVSS.n4441 VSS 0.331802f
C13006 DVSS.n4442 VSS 0.048967f
C13007 DVSS.n4444 VSS 0.026154f
C13008 DVSS.n4445 VSS 0.026154f
C13009 DVSS.n4447 VSS 0.026154f
C13010 DVSS.n4448 VSS 0.041971f
C13011 DVSS.n4449 VSS 0.745601f
C13012 DVSS.n4450 VSS 0.022779f
C13013 DVSS.n4451 VSS 0.361112f
C13014 DVSS.n4452 VSS 0.439768f
C13015 DVSS.n4453 VSS 0.439768f
C13016 DVSS.n4454 VSS 0.022779f
C13017 DVSS.n4455 VSS 0.041129f
C13018 DVSS.n4459 VSS 0.044082f
C13019 DVSS.n4460 VSS 0.026154f
C13020 DVSS.n4461 VSS 0.329631f
C13021 DVSS.n4463 VSS 0.032106f
C13022 DVSS.n4464 VSS 0.032106f
C13023 DVSS.n4466 VSS 0.032106f
C13024 DVSS.n4468 VSS 0.032106f
C13025 DVSS.n4470 VSS 0.120696f
C13026 DVSS.n4471 VSS 0.026154f
C13027 DVSS.n4473 VSS 0.127236f
C13028 DVSS.n4474 VSS 0.127236f
C13029 DVSS.n4475 VSS 0.026154f
C13030 DVSS.n4477 VSS 0.133296f
C13031 DVSS.n4478 VSS 0.026154f
C13032 DVSS.n4479 VSS 0.28709f
C13033 DVSS.n4480 VSS 0.150696f
C13034 DVSS.n4481 VSS 0.065797f
C13035 DVSS.n4482 VSS 0.052308f
C13036 DVSS.n4484 VSS 0.052308f
C13037 DVSS.n4485 VSS 0.052308f
C13038 DVSS.n4487 VSS 0.052308f
C13039 DVSS.n4489 VSS 0.065797f
C13040 DVSS.n4490 VSS 0.075348f
C13041 DVSS.n4491 VSS 0.022779f
C13042 DVSS.n4492 VSS 0.075348f
C13043 DVSS.n4493 VSS 0.065797f
C13044 DVSS.n4494 VSS 0.150696f
C13045 DVSS.n4495 VSS 0.150696f
C13046 DVSS.n4496 VSS 0.150696f
C13047 DVSS.n4497 VSS 0.150696f
C13048 DVSS.n4498 VSS 0.150696f
C13049 DVSS.n4499 VSS 0.150696f
C13050 DVSS.n4500 VSS 0.150696f
C13051 DVSS.n4501 VSS 0.134247f
C13052 DVSS.n4502 VSS 0.150696f
C13053 DVSS.n4503 VSS 0.150696f
C13054 DVSS.n4504 VSS 0.150696f
C13055 DVSS.n4505 VSS 0.150696f
C13056 DVSS.n4506 VSS 0.150696f
C13057 DVSS.n4507 VSS 0.150696f
C13058 DVSS.n4508 VSS 0.065797f
C13059 DVSS.n4509 VSS 0.052308f
C13060 DVSS.n4511 VSS 0.052308f
C13061 DVSS.n4512 VSS 0.052308f
C13062 DVSS.n4514 VSS 0.052308f
C13063 DVSS.n4516 VSS 0.065797f
C13064 DVSS.n4517 VSS 0.075348f
C13065 DVSS.n4518 VSS 0.022779f
C13066 DVSS.n4519 VSS 0.075348f
C13067 DVSS.n4520 VSS 0.065797f
C13068 DVSS.n4521 VSS 0.150696f
C13069 DVSS.n4522 VSS 0.150696f
C13070 DVSS.n4523 VSS 0.150696f
C13071 DVSS.n4524 VSS 0.150696f
C13072 DVSS.n4525 VSS 0.150696f
C13073 DVSS.n4526 VSS 0.150696f
C13074 DVSS.n4527 VSS 0.150696f
C13075 DVSS.n4528 VSS 0.150696f
C13076 DVSS.n4529 VSS 0.150696f
C13077 DVSS.n4530 VSS 0.150696f
C13078 DVSS.n4531 VSS 0.150696f
C13079 DVSS.n4532 VSS 0.150696f
C13080 DVSS.n4533 VSS 0.150696f
C13081 DVSS.n4534 VSS 0.150696f
C13082 DVSS.n4535 VSS 0.150696f
C13083 DVSS.n4536 VSS 0.150696f
C13084 DVSS.n4537 VSS 0.150696f
C13085 DVSS.n4538 VSS 0.150696f
C13086 DVSS.n4539 VSS 0.150696f
C13087 DVSS.n4540 VSS 0.150696f
C13088 DVSS.n4541 VSS 0.150696f
C13089 DVSS.n4542 VSS 0.150696f
C13090 DVSS.n4543 VSS 0.150696f
C13091 DVSS.n4544 VSS 0.150696f
C13092 DVSS.n4545 VSS 0.150696f
C13093 DVSS.n4546 VSS 0.150696f
C13094 DVSS.n4547 VSS 0.150696f
C13095 DVSS.n4548 VSS 0.150696f
C13096 DVSS.n4549 VSS 0.150696f
C13097 DVSS.n4550 VSS 0.150696f
C13098 DVSS.n4551 VSS 0.150696f
C13099 DVSS.n4552 VSS 0.150696f
C13100 DVSS.n4553 VSS 0.150696f
C13101 DVSS.n4554 VSS 0.150696f
C13102 DVSS.n4555 VSS 0.150696f
C13103 DVSS.n4556 VSS 0.150696f
C13104 DVSS.n4557 VSS 0.150696f
C13105 DVSS.n4558 VSS 0.150696f
C13106 DVSS.n4559 VSS 0.150696f
C13107 DVSS.n4560 VSS 0.150696f
C13108 DVSS.n4561 VSS 0.150696f
C13109 DVSS.n4562 VSS 0.150696f
C13110 DVSS.n4563 VSS 0.150696f
C13111 DVSS.n4564 VSS 0.150696f
C13112 DVSS.n4565 VSS 0.150696f
C13113 DVSS.n4566 VSS 0.150696f
C13114 DVSS.n4567 VSS 0.150696f
C13115 DVSS.n4568 VSS 0.150696f
C13116 DVSS.n4569 VSS 0.150696f
C13117 DVSS.n4570 VSS 0.150696f
C13118 DVSS.n4571 VSS 0.150696f
C13119 DVSS.n4572 VSS 0.120451f
C13120 DVSS.n4573 VSS 0.150696f
C13121 DVSS.n4574 VSS 0.065797f
C13122 DVSS.n4575 VSS 0.150696f
C13123 DVSS.n4576 VSS 0.065797f
C13124 DVSS.n4577 VSS 0.150696f
C13125 DVSS.n4578 VSS 0.150696f
C13126 DVSS.n4579 VSS 0.065797f
C13127 DVSS.n4581 VSS 0.041129f
C13128 DVSS.n4584 VSS 0.052308f
C13129 DVSS.n4587 VSS 0.052308f
C13130 DVSS.n4588 VSS 0.075348f
C13131 DVSS.n4589 VSS 0.022779f
C13132 DVSS.n4590 VSS 0.026154f
C13133 DVSS.n4593 VSS 0.032106f
C13134 DVSS.n4594 VSS 0.026154f
C13135 DVSS.n4595 VSS 0.289551f
C13136 DVSS.n4596 VSS 0.289551f
C13137 DVSS.n4598 VSS 0.026154f
C13138 DVSS.n4599 VSS 0.291484f
C13139 DVSS.n4600 VSS 0.291484f
C13140 DVSS.n4601 VSS 0.032106f
C13141 DVSS.n4602 VSS 0.021932f
C13142 DVSS.n4604 VSS 0.032106f
C13143 DVSS.n4606 VSS 0.021932f
C13144 DVSS.n4607 VSS 0.065797f
C13145 DVSS.n4608 VSS 0.101879f
C13146 DVSS.n4609 VSS 0.150696f
C13147 DVSS.n4610 VSS 0.150696f
C13148 DVSS.n4611 VSS 0.150696f
C13149 DVSS.n4612 VSS 0.150696f
C13150 DVSS.n4613 VSS 0.150696f
C13151 DVSS.n4614 VSS 0.150696f
C13152 DVSS.n4615 VSS 0.150696f
C13153 DVSS.n4616 VSS 0.075348f
C13154 DVSS.n4617 VSS 0.019102f
C13155 DVSS.n4618 VSS 0.019102f
C13156 DVSS.n4620 VSS 0.021932f
C13157 DVSS.n4621 VSS 0.019102f
C13158 DVSS.n4622 VSS 0.065797f
C13159 DVSS.n4623 VSS 0.019102f
C13160 DVSS.n4624 VSS 0.019102f
C13161 DVSS.n4625 VSS 0.021932f
C13162 DVSS.n4626 VSS 0.021932f
C13163 DVSS.n4627 VSS 0.021932f
C13164 DVSS.n4628 VSS 0.01981f
C13165 DVSS.n4629 VSS 0.035873f
C13166 DVSS.n4630 VSS 0.038205f
C13167 DVSS.n4631 VSS 0.038205f
C13168 DVSS.n4632 VSS 0.038205f
C13169 DVSS.n4633 VSS 0.038205f
C13170 DVSS.n4634 VSS 0.038205f
C13171 DVSS.n4635 VSS 0.035873f
C13172 DVSS.n4636 VSS 0.038205f
C13173 DVSS.n4637 VSS 0.038205f
C13174 DVSS.n4638 VSS 0.038205f
C13175 DVSS.n4639 VSS 0.038205f
C13176 DVSS.n4640 VSS 0.038205f
C13177 DVSS.n4641 VSS 0.026905f
C13178 DVSS.n4642 VSS 0.038205f
C13179 DVSS.t13 VSS 0.330478f
C13180 DVSS.n4643 VSS 0.125906f
C13181 DVSS.n4644 VSS 0.038205f
C13182 DVSS.n4645 VSS 0.038205f
C13183 DVSS.n4646 VSS 0.038205f
C13184 DVSS.n4647 VSS 0.038205f
C13185 DVSS.n4648 VSS 0.035873f
C13186 DVSS.n4649 VSS 0.038205f
C13187 DVSS.n4650 VSS 0.038205f
C13188 DVSS.n4651 VSS 0.038205f
C13189 DVSS.n4652 VSS 0.038205f
C13190 DVSS.n4653 VSS 0.038205f
C13191 DVSS.n4654 VSS 0.035873f
C13192 DVSS.n4655 VSS 0.038205f
C13193 DVSS.n4656 VSS 0.021402f
C13194 DVSS.n4657 VSS 0.021932f
C13195 DVSS.n4658 VSS 0.021932f
C13196 DVSS.n4659 VSS 0.021932f
C13197 DVSS.n4660 VSS 0.021932f
C13198 DVSS.n4661 VSS 0.035873f
C13199 DVSS.n4662 VSS 0.021932f
C13200 DVSS.n4663 VSS 0.035873f
C13201 DVSS.n4664 VSS 0.021932f
C13202 DVSS.n4665 VSS 0.035873f
C13203 DVSS.n4666 VSS 0.035873f
C13204 DVSS.n4667 VSS 0.021402f
C13205 DVSS.n4668 VSS 0.038205f
C13206 DVSS.n4669 VSS 0.038205f
C13207 DVSS.n4670 VSS 0.035873f
C13208 DVSS.n4671 VSS 0.035873f
C13209 DVSS.n4672 VSS 0.035873f
C13210 DVSS.n4673 VSS 0.038205f
C13211 DVSS.n4674 VSS 0.038205f
C13212 DVSS.n4675 VSS 0.038205f
C13213 DVSS.n4676 VSS 0.033714f
C13214 DVSS.n4677 VSS 0.020096f
C13215 DVSS.n4678 VSS 0.026905f
C13216 DVSS.n4679 VSS 0.038205f
C13217 DVSS.n4680 VSS 0.038205f
C13218 DVSS.n4681 VSS 0.038205f
C13219 DVSS.n4682 VSS 0.035873f
C13220 DVSS.n4683 VSS 0.035873f
C13221 DVSS.n4684 VSS 0.035873f
C13222 DVSS.n4685 VSS 0.038205f
C13223 DVSS.n4686 VSS 0.038205f
C13224 DVSS.n4687 VSS 0.038205f
C13225 DVSS.n4688 VSS 0.035873f
C13226 DVSS.n4689 VSS 0.035873f
C13227 DVSS.n4690 VSS 0.035873f
C13228 DVSS.n4691 VSS 0.038205f
C13229 DVSS.n4692 VSS 0.038205f
C13230 DVSS.n4693 VSS 0.01981f
C13231 DVSS.n4694 VSS 0.035873f
C13232 DVSS.n4695 VSS 0.021932f
C13233 DVSS.n4696 VSS 0.035873f
C13234 DVSS.n4697 VSS 0.021932f
C13235 DVSS.n4698 VSS 0.035873f
C13236 DVSS.n4699 VSS 0.021932f
C13237 DVSS.n4700 VSS 0.035873f
C13238 DVSS.n4701 VSS 0.021932f
C13239 DVSS.n4702 VSS 0.031887f
C13240 DVSS.n4703 VSS 0.021932f
C13241 DVSS.n4704 VSS 0.03396f
C13242 DVSS.n4705 VSS 0.150696f
C13243 DVSS.n4706 VSS 0.150696f
C13244 DVSS.n4707 VSS 0.150696f
C13245 DVSS.n4708 VSS 0.150696f
C13246 DVSS.n4709 VSS 0.150696f
C13247 DVSS.n4710 VSS 0.150696f
C13248 DVSS.n4711 VSS 0.150696f
C13249 DVSS.n4712 VSS 0.150696f
C13250 DVSS.n4713 VSS 0.150696f
C13251 DVSS.n4714 VSS 0.150696f
C13252 DVSS.n4715 VSS 0.150696f
C13253 DVSS.n4716 VSS 0.150696f
C13254 DVSS.n4717 VSS 0.150696f
C13255 DVSS.n4718 VSS 0.150696f
C13256 DVSS.n4719 VSS 0.150696f
C13257 DVSS.n4720 VSS 0.150696f
C13258 DVSS.n4721 VSS 0.150696f
C13259 DVSS.n4722 VSS 0.150696f
C13260 DVSS.n4723 VSS 0.150696f
C13261 DVSS.n4724 VSS 0.150696f
C13262 DVSS.n4725 VSS 0.150696f
C13263 DVSS.n4726 VSS 0.150696f
C13264 DVSS.n4727 VSS 0.150696f
C13265 DVSS.n4728 VSS 0.150696f
C13266 DVSS.n4729 VSS 0.150696f
C13267 DVSS.n4730 VSS 0.150696f
C13268 DVSS.n4731 VSS 0.150696f
C13269 DVSS.n4732 VSS 0.150696f
C13270 DVSS.n4733 VSS 0.150696f
C13271 DVSS.n4734 VSS 0.150696f
C13272 DVSS.n4735 VSS 0.150696f
C13273 DVSS.n4736 VSS 0.150696f
C13274 DVSS.n4737 VSS 0.150696f
C13275 DVSS.n4738 VSS 0.150696f
C13276 DVSS.n4739 VSS 0.150696f
C13277 DVSS.n4740 VSS 0.150696f
C13278 DVSS.n4741 VSS 0.150696f
C13279 DVSS.n4742 VSS 0.150696f
C13280 DVSS.n4743 VSS 0.150696f
C13281 DVSS.n4744 VSS 0.143268f
C13282 DVSS.n4745 VSS 0.03449f
C13283 DVSS.n4746 VSS 0.075348f
C13284 DVSS.n4747 VSS 0.050586f
C13285 DVSS.n4749 VSS 0.075348f
C13286 DVSS.n4750 VSS 0.065797f
C13287 DVSS.n4751 VSS 0.150696f
C13288 DVSS.n4752 VSS 0.150696f
C13289 DVSS.n4753 VSS 0.150696f
C13290 DVSS.n4754 VSS 0.099757f
C13291 DVSS.n4755 VSS 0.075348f
C13292 DVSS.n4756 VSS 0.019102f
C13293 DVSS.n4757 VSS 0.075348f
C13294 DVSS.n4758 VSS 0.14539f
C13295 DVSS.n4759 VSS 0.150696f
C13296 DVSS.n4760 VSS 0.150696f
C13297 DVSS.n4761 VSS 0.150696f
C13298 DVSS.n4762 VSS 0.150696f
C13299 DVSS.n4763 VSS 0.150696f
C13300 DVSS.n4764 VSS 0.150696f
C13301 DVSS.n4765 VSS 0.150696f
C13302 DVSS.n4766 VSS 0.150696f
C13303 DVSS.n4767 VSS 0.150696f
C13304 DVSS.n4768 VSS 0.150696f
C13305 DVSS.n4769 VSS 0.150696f
C13306 DVSS.n4770 VSS 0.150696f
C13307 DVSS.n4771 VSS 0.150696f
C13308 DVSS.n4772 VSS 0.150696f
C13309 DVSS.n4773 VSS 0.150696f
C13310 DVSS.n4774 VSS 0.150696f
C13311 DVSS.n4775 VSS 0.150696f
C13312 DVSS.n4776 VSS 0.120451f
C13313 DVSS.n4777 VSS 0.150696f
C13314 DVSS.n4778 VSS 0.065797f
C13315 DVSS.n4779 VSS 0.150696f
C13316 DVSS.n4780 VSS 0.150696f
C13317 DVSS.n4781 VSS 0.065797f
C13318 DVSS.n4782 VSS 0.075348f
C13319 DVSS.n4783 VSS 0.022779f
C13320 DVSS.n4784 VSS 0.075348f
C13321 DVSS.n4785 VSS 0.439768f
C13322 DVSS.n4787 VSS 0.439768f
C13323 DVSS.n4790 VSS 0.052308f
C13324 DVSS.n4793 VSS 0.052308f
C13325 DVSS.n4795 VSS 0.036911f
C13326 DVSS.n4796 VSS 0.082541f
C13327 DVSS.n4797 VSS 0.026154f
C13328 DVSS.n4798 VSS 0.026154f
C13329 DVSS.n4801 VSS 0.066724f
C13330 DVSS.n4802 VSS 0.026154f
C13331 DVSS.n4803 VSS 0.186719f
C13332 DVSS.n4804 VSS 0.396845f
C13333 DVSS.n4805 VSS 0.021932f
C13334 DVSS.n4806 VSS 0.065379f
C13335 DVSS.n4807 VSS 0.056423f
C13336 DVSS.n4808 VSS 0.021932f
C13337 DVSS.n4809 VSS 0.082541f
C13338 DVSS.n4810 VSS 0.038382f
C13339 DVSS.n4811 VSS 0.021932f
C13340 DVSS.n4812 VSS 0.049824f
C13341 DVSS.n4813 VSS 0.021932f
C13342 DVSS.n4814 VSS 0.019102f
C13343 DVSS.n4816 VSS 0.030953f
C13344 DVSS.n4817 VSS 0.082541f
C13345 DVSS.n4818 VSS 0.021932f
C13346 DVSS.n4819 VSS 0.021932f
C13347 DVSS.n4821 VSS 0.065379f
C13348 DVSS.n4822 VSS 0.021932f
C13349 DVSS.n4823 VSS 0.396845f
C13350 DVSS.n4824 VSS 0.186719f
C13351 DVSS.n4825 VSS 0.066724f
C13352 DVSS.n4827 VSS 0.026154f
C13353 DVSS.t29 VSS 0.394423f
C13354 DVSS.n4829 VSS 0.635269f
C13355 DVSS.n4830 VSS 0.026154f
C13356 DVSS.n4832 VSS 0.026154f
C13357 DVSS.n4833 VSS 0.066724f
C13358 DVSS.n4835 VSS 0.066724f
C13359 DVSS.n4837 VSS 0.09309f
C13360 DVSS.n4838 VSS 0.026154f
C13361 DVSS.n4839 VSS 0.335771f
C13362 DVSS.n4840 VSS 0.756156f
C13363 DVSS.n4842 VSS 0.738852f
C13364 DVSS.n4843 VSS 0.026154f
C13365 DVSS.n4844 VSS 0.026154f
C13366 DVSS.n4845 VSS 0.242143f
C13367 DVSS.n4846 VSS 0.026154f
C13368 DVSS.n4847 VSS 0.036911f
C13369 DVSS.n4848 VSS 0.082541f
C13370 DVSS.n4849 VSS 0.439768f
C13371 DVSS.n4850 VSS 0.082541f
C13372 DVSS.n4851 VSS 0.072078f
C13373 DVSS.n4852 VSS 0.165082f
C13374 DVSS.n4853 VSS 0.165082f
C13375 DVSS.n4854 VSS 0.165082f
C13376 DVSS.n4855 VSS 0.165082f
C13377 DVSS.n4856 VSS 0.165082f
C13378 DVSS.n4857 VSS 0.165082f
C13379 DVSS.n4858 VSS 0.165082f
C13380 DVSS.n4859 VSS 0.165082f
C13381 DVSS.n4860 VSS 0.165082f
C13382 DVSS.n4861 VSS 0.165082f
C13383 DVSS.n4862 VSS 0.165082f
C13384 DVSS.n4863 VSS 0.165082f
C13385 DVSS.n4864 VSS 0.165082f
C13386 DVSS.n4865 VSS 0.165082f
C13387 DVSS.n4866 VSS 0.165082f
C13388 DVSS.n4867 VSS 0.165082f
C13389 DVSS.n4868 VSS 0.165082f
C13390 DVSS.n4869 VSS 0.165082f
C13391 DVSS.n4870 VSS 0.165082f
C13392 DVSS.n4871 VSS 0.165082f
C13393 DVSS.n4872 VSS 0.165082f
C13394 DVSS.n4873 VSS 0.165082f
C13395 DVSS.n4874 VSS 0.165082f
C13396 DVSS.n4875 VSS 0.165082f
C13397 DVSS.n4876 VSS 0.165082f
C13398 DVSS.n4877 VSS 0.165082f
C13399 DVSS.n4878 VSS 0.165082f
C13400 DVSS.n4879 VSS 0.165082f
C13401 DVSS.n4880 VSS 0.165082f
C13402 DVSS.n4881 VSS 0.072078f
C13403 DVSS.n4883 VSS 0.052308f
C13404 DVSS.n4885 VSS 0.052308f
C13405 DVSS.n4886 VSS 0.082541f
C13406 DVSS.n4887 VSS 0.026154f
C13407 DVSS.n4888 VSS 0.082541f
C13408 DVSS.n4889 VSS 0.072078f
C13409 DVSS.n4890 VSS 0.165082f
C13410 DVSS.n4891 VSS 0.165082f
C13411 DVSS.n4892 VSS 0.165082f
C13412 DVSS.n4893 VSS 0.165082f
C13413 DVSS.n4894 VSS 0.165082f
C13414 DVSS.n4895 VSS 0.165082f
C13415 DVSS.n4896 VSS 0.165082f
C13416 DVSS.n4897 VSS 0.165082f
C13417 DVSS.n4898 VSS 0.165082f
C13418 DVSS.n4899 VSS 0.165082f
C13419 DVSS.n4900 VSS 0.165082f
C13420 DVSS.n4901 VSS 0.165082f
C13421 DVSS.n4902 VSS 0.165082f
C13422 DVSS.n4903 VSS 0.148806f
C13423 DVSS.n4904 VSS 0.148806f
C13424 DVSS.n4905 VSS 0.165082f
C13425 DVSS.n4906 VSS 0.165082f
C13426 DVSS.n4907 VSS 0.022779f
C13427 DVSS.n4908 VSS 0.022779f
C13428 DVSS.n4909 VSS 0.052308f
C13429 DVSS.n4910 VSS 0.052308f
C13430 DVSS.n4911 VSS 0.052308f
C13431 DVSS.n4912 VSS 0.072078f
C13432 DVSS.n4913 VSS 0.439768f
C13433 DVSS.n4914 VSS 0.052308f
C13434 DVSS.n4915 VSS 0.052308f
C13435 DVSS.n4916 VSS 0.04366f
C13436 DVSS.n4917 VSS 0.022779f
C13437 DVSS.n4918 VSS 0.026154f
C13438 DVSS.n4922 VSS 0.082541f
C13439 DVSS.n4926 VSS 0.363609f
C13440 DVSS.n4928 VSS 0.058114f
C13441 DVSS.n4929 VSS 0.026154f
C13442 DVSS.n4931 VSS 0.026154f
C13443 DVSS.n4932 VSS 0.026154f
C13444 DVSS.n4933 VSS 0.048967f
C13445 DVSS.n4934 VSS 0.745601f
C13446 DVSS.n4935 VSS 0.072078f
C13447 DVSS.n4936 VSS 0.165082f
C13448 DVSS.n4937 VSS 0.162757f
C13449 DVSS.n4938 VSS 0.616179f
C13450 DVSS.n4939 VSS 0.319361f
C13451 DVSS.n4940 VSS 0.165082f
C13452 DVSS.n4941 VSS 0.072078f
C13453 DVSS.n4942 VSS 0.082541f
C13454 DVSS.n4943 VSS 0.022779f
C13455 DVSS.n4944 VSS 0.082541f
C13456 DVSS.n4945 VSS 0.068009f
C13457 DVSS.n4946 VSS 0.098817f
C13458 DVSS.n4947 VSS 0.084866f
C13459 DVSS.n4948 VSS 0.165082f
C13460 DVSS.n4949 VSS 0.165082f
C13461 DVSS.n4950 VSS 0.165082f
C13462 DVSS.n4951 VSS 0.165082f
C13463 DVSS.n4952 VSS 0.165082f
C13464 DVSS.n4953 VSS 0.144737f
C13465 DVSS.n4954 VSS 0.165082f
C13466 DVSS.n4955 VSS 0.072078f
C13467 DVSS.n4956 VSS 0.165082f
C13468 DVSS.n4957 VSS 0.165082f
C13469 DVSS.n4958 VSS 0.165082f
C13470 DVSS.n4959 VSS 0.165082f
C13471 DVSS.n4960 VSS 0.165082f
C13472 DVSS.n4961 VSS 0.072078f
C13473 DVSS.n4963 VSS 0.439768f
C13474 DVSS.n4966 VSS 0.052308f
C13475 DVSS.n4969 VSS 0.052308f
C13476 DVSS.n4971 VSS 0.036911f
C13477 DVSS.n4972 VSS 0.082541f
C13478 DVSS.n4973 VSS 0.026154f
C13479 DVSS.n4974 VSS 0.026154f
C13480 DVSS.n4976 VSS 0.066724f
C13481 DVSS.n4977 VSS 0.026154f
C13482 DVSS.n4978 VSS 0.222771f
C13483 DVSS.n4979 VSS 0.738852f
C13484 DVSS.n4980 VSS 0.740117f
C13485 DVSS.n4982 VSS 0.026154f
C13486 DVSS.n4983 VSS 0.026154f
C13487 DVSS.n4984 VSS 0.066724f
C13488 DVSS.n4986 VSS 0.066724f
C13489 DVSS.n4987 VSS 0.026154f
C13490 DVSS.n4989 VSS 0.222771f
C13491 DVSS.n4990 VSS 0.026154f
C13492 DVSS.n4991 VSS 0.179185f
C13493 DVSS.n4992 VSS 0.09309f
C13494 DVSS.n4993 VSS 0.026154f
C13495 DVSS.n4994 VSS 0.335771f
C13496 DVSS.n4995 VSS 0.756156f
C13497 DVSS.n4996 VSS 0.242143f
C13498 DVSS.n4997 VSS 0.026154f
C13499 DVSS.n4998 VSS 0.186719f
C13500 DVSS.n4999 VSS 0.032014f
C13501 DVSS.n5000 VSS 0.021932f
C13502 DVSS.n5001 VSS 0.396845f
C13503 DVSS.n5002 VSS 0.021932f
C13504 DVSS.n5003 VSS 0.065379f
C13505 DVSS.n5004 VSS -0.427302f
C13506 DVSS.n5005 VSS 48.8624f
C13507 DVSS.n5006 VSS 48.8624f
C13508 DVSS.n5007 VSS -0.427302f
C13509 DVSS.n5008 VSS 0.019102f
C13510 DVSS.n5010 VSS 0.082541f
C13511 DVSS.n5011 VSS 0.111605f
C13512 DVSS.n5012 VSS 0.021932f
C13513 DVSS.n5013 VSS 0.021932f
C13514 DVSS.n5014 VSS 0.03449f
C13515 DVSS.n5015 VSS 0.019102f
C13516 DVSS.n5016 VSS 0.072078f
C13517 DVSS.n5017 VSS 0.019102f
C13518 DVSS.n5018 VSS 0.019102f
C13519 DVSS.n5019 VSS 0.021932f
C13520 DVSS.n5020 VSS 0.021932f
C13521 DVSS.n5022 VSS 0.021932f
C13522 DVSS.n5024 VSS 0.021932f
C13523 DVSS.n5025 VSS 0.066724f
C13524 DVSS.n5026 VSS 0.021932f
C13525 DVSS.n5027 VSS 0.065379f
C13526 DVSS.n5028 VSS 0.021932f
C13527 DVSS.n5029 VSS 0.396845f
C13528 DVSS.n5030 VSS 0.021932f
C13529 DVSS.n5031 VSS 0.165082f
C13530 DVSS.n5032 VSS 0.165082f
C13531 DVSS.n5033 VSS 0.165082f
C13532 DVSS.n5034 VSS 0.165082f
C13533 DVSS.n5035 VSS 0.165082f
C13534 DVSS.n5036 VSS 0.165082f
C13535 DVSS.n5037 VSS 0.165082f
C13536 DVSS.n5038 VSS 0.156944f
C13537 DVSS.n5039 VSS 0.165082f
C13538 DVSS.n5040 VSS 0.165082f
C13539 DVSS.n5041 VSS 0.165082f
C13540 DVSS.n5042 VSS 0.165082f
C13541 DVSS.n5043 VSS 0.165082f
C13542 DVSS.n5044 VSS 0.165082f
C13543 DVSS.n5045 VSS 0.165082f
C13544 DVSS.n5046 VSS 0.165082f
C13545 DVSS.n5047 VSS 0.134274f
C13546 DVSS.n5048 VSS 0.165082f
C13547 DVSS.n5049 VSS 0.165082f
C13548 DVSS.n5050 VSS 0.165082f
C13549 DVSS.n5051 VSS 0.165082f
C13550 DVSS.n5052 VSS 0.165082f
C13551 DVSS.n5053 VSS 0.165082f
C13552 DVSS.n5054 VSS 0.165082f
C13553 DVSS.n5055 VSS 0.165082f
C13554 DVSS.n5056 VSS 0.165082f
C13555 DVSS.n5057 VSS 0.165082f
C13556 DVSS.n5058 VSS 0.165082f
C13557 DVSS.n5059 VSS 0.165082f
C13558 DVSS.n5060 VSS 0.165082f
C13559 DVSS.n5061 VSS 0.134274f
C13560 DVSS.n5062 VSS 0.165082f
C13561 DVSS.n5063 VSS 0.165082f
C13562 DVSS.n5064 VSS 0.165082f
C13563 DVSS.n5065 VSS 0.082541f
C13564 DVSS.n5066 VSS 0.026154f
C13565 DVSS.n5067 VSS 0.041129f
C13566 DVSS.n5068 VSS 0.072078f
C13567 DVSS.n5071 VSS 0.026154f
C13568 DVSS.n5072 VSS 0.026154f
C13569 DVSS.n5073 VSS 0.082541f
C13570 DVSS.n5074 VSS 0.072078f
C13571 DVSS.n5075 VSS 0.052308f
C13572 DVSS.n5077 VSS 0.052308f
C13573 DVSS.n5078 VSS 0.052308f
C13574 DVSS.n5080 VSS 0.052308f
C13575 DVSS.n5082 VSS 0.165082f
C13576 DVSS.n5083 VSS 0.165082f
C13577 DVSS.n5084 VSS 0.165082f
C13578 DVSS.n5085 VSS 0.165082f
C13579 DVSS.n5086 VSS 0.165082f
C13580 DVSS.n5087 VSS 0.165082f
C13581 DVSS.n5088 VSS 0.072078f
C13582 DVSS.n5089 VSS 0.165082f
C13583 DVSS.n5090 VSS 0.165082f
C13584 DVSS.n5091 VSS 0.165082f
C13585 DVSS.n5092 VSS 0.165082f
C13586 DVSS.n5093 VSS 0.165082f
C13587 DVSS.n5094 VSS 0.319361f
C13588 DVSS.n5095 VSS 0.072078f
C13589 DVSS.n5096 VSS 0.165082f
C13590 DVSS.n5097 VSS 0.072078f
C13591 DVSS.n5098 VSS 0.165082f
C13592 DVSS.n5099 VSS 0.616179f
C13593 DVSS.n5100 VSS 0.162757f
C13594 DVSS.n5101 VSS 0.084866f
C13595 DVSS.n5102 VSS 0.098817f
C13596 DVSS.n5103 VSS 0.148806f
C13597 DVSS.n5104 VSS 0.165082f
C13598 DVSS.n5105 VSS 0.148806f
C13599 DVSS.n5106 VSS 0.165082f
C13600 DVSS.n5107 VSS 0.165082f
C13601 DVSS.n5108 VSS 0.165082f
C13602 DVSS.n5109 VSS 0.165082f
C13603 DVSS.n5110 VSS 0.165082f
C13604 DVSS.n5111 VSS 0.165082f
C13605 DVSS.n5112 VSS 0.165082f
C13606 DVSS.n5113 VSS 0.072078f
C13607 DVSS.n5114 VSS 0.165082f
C13608 DVSS.n5115 VSS 0.165082f
C13609 DVSS.n5116 VSS 0.165082f
C13610 DVSS.n5117 VSS 0.165082f
C13611 DVSS.n5118 VSS 0.165082f
C13612 DVSS.n5119 VSS 0.134274f
C13613 DVSS.n5120 VSS 0.165082f
C13614 DVSS.n5121 VSS 0.165082f
C13615 DVSS.n5122 VSS 0.165082f
C13616 DVSS.n5123 VSS 0.165082f
C13617 DVSS.n5124 VSS 0.165082f
C13618 DVSS.n5125 VSS 0.165082f
C13619 DVSS.n5126 VSS 0.165082f
C13620 DVSS.n5127 VSS 0.144737f
C13621 DVSS.n5128 VSS 0.082541f
C13622 DVSS.n5129 VSS 0.728095f
C13623 DVSS.n5130 VSS 0.082541f
C13624 DVSS.n5131 VSS 0.072078f
C13625 DVSS.n5132 VSS 0.165082f
C13626 DVSS.n5133 VSS 0.165082f
C13627 DVSS.n5134 VSS 0.165082f
C13628 DVSS.n5135 VSS 0.165082f
C13629 DVSS.n5136 VSS 0.165082f
C13630 DVSS.n5137 VSS 0.165082f
C13631 DVSS.n5138 VSS 0.165082f
C13632 DVSS.n5139 VSS 0.165082f
C13633 DVSS.n5140 VSS 0.165082f
C13634 DVSS.n5141 VSS 0.165082f
C13635 DVSS.n5142 VSS 0.165082f
C13636 DVSS.n5143 VSS 0.165082f
C13637 DVSS.n5144 VSS 0.165082f
C13638 DVSS.n5145 VSS 0.165082f
C13639 DVSS.n5146 VSS 0.165082f
C13640 DVSS.n5147 VSS 0.165082f
C13641 DVSS.n5148 VSS 0.165082f
C13642 DVSS.n5149 VSS 0.165082f
C13643 DVSS.n5150 VSS 0.165082f
C13644 DVSS.n5151 VSS 0.165082f
C13645 DVSS.n5152 VSS 0.165082f
C13646 DVSS.n5153 VSS 0.165082f
C13647 DVSS.n5154 VSS 0.165082f
C13648 DVSS.n5155 VSS 0.165082f
C13649 DVSS.n5156 VSS 0.165082f
C13650 DVSS.n5157 VSS 0.165082f
C13651 DVSS.n5158 VSS 0.165082f
C13652 DVSS.n5159 VSS 0.165082f
C13653 DVSS.n5160 VSS 0.165082f
C13654 DVSS.n5161 VSS 0.072078f
C13655 DVSS.n5162 VSS 0.165082f
C13656 DVSS.n5163 VSS 0.072078f
C13657 DVSS.n5164 VSS 0.165082f
C13658 DVSS.n5165 VSS 0.165082f
C13659 DVSS.n5166 VSS 0.165082f
C13660 DVSS.n5167 VSS 0.165082f
C13661 DVSS.n5168 VSS 0.165082f
C13662 DVSS.n5169 VSS 0.165082f
C13663 DVSS.n5170 VSS 0.165082f
C13664 DVSS.n5171 VSS 0.165082f
C13665 DVSS.n5172 VSS 0.165082f
C13666 DVSS.n5173 VSS 0.165082f
C13667 DVSS.n5174 VSS 0.165082f
C13668 DVSS.n5175 VSS 0.165082f
C13669 DVSS.n5176 VSS 0.165082f
C13670 DVSS.n5177 VSS 0.165082f
C13671 DVSS.n5178 VSS 0.165082f
C13672 DVSS.n5179 VSS 0.165082f
C13673 DVSS.n5180 VSS 0.165082f
C13674 DVSS.n5181 VSS 0.165082f
C13675 DVSS.n5182 VSS 0.165082f
C13676 DVSS.n5183 VSS 0.165082f
C13677 DVSS.n5184 VSS 0.165082f
C13678 DVSS.n5185 VSS 0.165082f
C13679 DVSS.n5186 VSS 0.165082f
C13680 DVSS.n5187 VSS 0.165082f
C13681 DVSS.n5188 VSS 0.165082f
C13682 DVSS.n5189 VSS 0.165082f
C13683 DVSS.n5190 VSS 0.165082f
C13684 DVSS.n5191 VSS 0.165082f
C13685 DVSS.n5192 VSS 0.165082f
C13686 DVSS.n5193 VSS 0.072078f
C13687 DVSS.n5194 VSS 0.082541f
C13688 DVSS.n5195 VSS 0.047402f
C13689 DVSS.n5196 VSS 0.082541f
C13690 DVSS.n5197 VSS 0.034844f
C13691 DVSS.n5198 VSS 0.021932f
C13692 DVSS.n5199 VSS 0.049824f
C13693 DVSS.n5200 VSS 0.021932f
C13694 DVSS.n5201 VSS 0.035873f
C13695 DVSS.n5202 VSS 0.021932f
C13696 DVSS.n5203 VSS 0.035873f
C13697 DVSS.n5204 VSS 0.021932f
C13698 DVSS.n5205 VSS 0.035873f
C13699 DVSS.n5206 VSS 0.035873f
C13700 DVSS.n5207 VSS 0.035873f
C13701 DVSS.n5208 VSS 0.038205f
C13702 DVSS.n5209 VSS 0.038205f
C13703 DVSS.n5210 VSS 0.038205f
C13704 DVSS.n5211 VSS 0.035873f
C13705 DVSS.n5212 VSS 0.035873f
C13706 DVSS.n5213 VSS 0.035873f
C13707 DVSS.n5214 VSS 0.038205f
C13708 DVSS.n5215 VSS 0.038205f
C13709 DVSS.n5216 VSS 0.038205f
C13710 DVSS.n5217 VSS 0.033714f
C13711 DVSS.n5218 VSS 0.020096f
C13712 DVSS.n5219 VSS 0.026905f
C13713 DVSS.n5220 VSS 0.038205f
C13714 DVSS.n5221 VSS 0.038205f
C13715 DVSS.n5222 VSS 0.026905f
C13716 DVSS.n5223 VSS 0.035873f
C13717 DVSS.n5224 VSS 0.035873f
C13718 DVSS.n5225 VSS 0.038205f
C13719 DVSS.n5226 VSS 0.038205f
C13720 DVSS.n5227 VSS 0.038205f
C13721 DVSS.n5228 VSS 0.035873f
C13722 DVSS.n5229 VSS 0.035873f
C13723 DVSS.n5230 VSS 0.035873f
C13724 DVSS.n5231 VSS 0.038205f
C13725 DVSS.n5232 VSS 0.038205f
C13726 DVSS.n5233 VSS 0.020341f
C13727 DVSS.n5234 VSS 0.035873f
C13728 DVSS.n5235 VSS 0.020341f
C13729 DVSS.n5236 VSS 0.019102f
C13730 DVSS.n5237 VSS 0.082541f
C13731 DVSS.n5238 VSS 0.072078f
C13732 DVSS.n5239 VSS 0.165082f
C13733 DVSS.n5240 VSS 0.165082f
C13734 DVSS.n5241 VSS 0.165082f
C13735 DVSS.n5242 VSS 0.165082f
C13736 DVSS.n5243 VSS 0.165082f
C13737 DVSS.n5244 VSS 0.156944f
C13738 DVSS.n5245 VSS 0.165082f
C13739 DVSS.n5246 VSS 0.165082f
C13740 DVSS.n5247 VSS 0.165082f
C13741 DVSS.n5248 VSS 0.165082f
C13742 DVSS.n5249 VSS 0.165082f
C13743 DVSS.n5250 VSS 0.165082f
C13744 DVSS.n5251 VSS 0.165082f
C13745 DVSS.n5252 VSS 0.165082f
C13746 DVSS.n5253 VSS 0.165082f
C13747 DVSS.n5254 VSS 0.165082f
C13748 DVSS.n5255 VSS 0.165082f
C13749 DVSS.n5256 VSS 0.165082f
C13750 DVSS.n5257 VSS 0.165082f
C13751 DVSS.n5258 VSS 0.165082f
C13752 DVSS.n5259 VSS 0.165082f
C13753 DVSS.n5260 VSS 0.165082f
C13754 DVSS.n5261 VSS 0.165082f
C13755 DVSS.n5262 VSS 0.165082f
C13756 DVSS.n5263 VSS 0.165082f
C13757 DVSS.n5264 VSS 0.165082f
C13758 DVSS.n5265 VSS 0.165082f
C13759 DVSS.n5266 VSS 0.165082f
C13760 DVSS.n5267 VSS 0.165082f
C13761 DVSS.n5268 VSS 0.134274f
C13762 DVSS.n5269 VSS 0.072078f
C13763 DVSS.n5270 VSS 0.082541f
C13764 DVSS.n5271 VSS 0.439557f
C13765 DVSS.n5272 VSS 0.082541f
C13766 DVSS.n5273 VSS 0.072078f
C13767 DVSS.n5274 VSS 0.165082f
C13768 DVSS.n5275 VSS 0.165082f
C13769 DVSS.n5276 VSS 0.165082f
C13770 DVSS.n5277 VSS 0.165082f
C13771 DVSS.n5278 VSS 0.165082f
C13772 DVSS.n5279 VSS 0.144737f
C13773 DVSS.n5280 VSS 0.165082f
C13774 DVSS.n5281 VSS 0.165082f
C13775 DVSS.n5282 VSS 0.165082f
C13776 DVSS.n5283 VSS 0.165082f
C13777 DVSS.n5284 VSS 0.165082f
C13778 DVSS.n5285 VSS 0.165082f
C13779 DVSS.n5286 VSS 0.165082f
C13780 DVSS.n5287 VSS 0.165082f
C13781 DVSS.n5288 VSS 0.165082f
C13782 DVSS.n5289 VSS 0.165082f
C13783 DVSS.n5290 VSS 0.165082f
C13784 DVSS.n5291 VSS 0.165082f
C13785 DVSS.n5292 VSS 0.165082f
C13786 DVSS.n5293 VSS 0.165082f
C13787 DVSS.n5294 VSS 0.165082f
C13788 DVSS.n5295 VSS 0.165082f
C13789 DVSS.n5296 VSS 0.165082f
C13790 DVSS.n5297 VSS 0.165082f
C13791 DVSS.n5298 VSS 0.165082f
C13792 DVSS.n5299 VSS 0.165082f
C13793 DVSS.n5300 VSS 0.165082f
C13794 DVSS.n5301 VSS 0.165082f
C13795 DVSS.n5302 VSS 0.165082f
C13796 DVSS.n5303 VSS 0.134274f
C13797 DVSS.n5304 VSS 0.072078f
C13798 DVSS.n5305 VSS 0.082541f
C13799 DVSS.n5306 VSS 0.439557f
C13800 DVSS.n5307 VSS 0.082541f
C13801 DVSS.n5308 VSS 0.072078f
C13802 DVSS.n5309 VSS 0.165082f
C13803 DVSS.n5310 VSS 0.165082f
C13804 DVSS.n5311 VSS 0.165082f
C13805 DVSS.n5312 VSS 0.165082f
C13806 DVSS.n5313 VSS 0.165082f
C13807 DVSS.n5314 VSS 0.144737f
C13808 DVSS.n5315 VSS 0.165082f
C13809 DVSS.n5316 VSS 0.165082f
C13810 DVSS.n5317 VSS 0.165082f
C13811 DVSS.n5318 VSS 0.165082f
C13812 DVSS.n5319 VSS 0.165082f
C13813 DVSS.n5320 VSS 0.165082f
C13814 DVSS.n5321 VSS 0.165082f
C13815 DVSS.n5322 VSS 0.165082f
C13816 DVSS.n5323 VSS 0.165082f
C13817 DVSS.n5324 VSS 0.072078f
C13818 DVSS.n5325 VSS 0.165082f
C13819 DVSS.n5326 VSS 0.165082f
C13820 DVSS.n5327 VSS 0.165082f
C13821 DVSS.n5328 VSS 0.165082f
C13822 DVSS.n5329 VSS 0.165082f
C13823 DVSS.n5330 VSS 0.319361f
C13824 DVSS.n5331 VSS 0.072078f
C13825 DVSS.n5332 VSS 0.165082f
C13826 DVSS.n5333 VSS 0.072078f
C13827 DVSS.n5334 VSS 0.165082f
C13828 DVSS.n5335 VSS 0.616179f
C13829 DVSS.n5336 VSS 0.162757f
C13830 DVSS.n5337 VSS 0.084866f
C13831 DVSS.n5338 VSS 0.098817f
C13832 DVSS.n5339 VSS 0.148806f
C13833 DVSS.n5340 VSS 0.148806f
C13834 DVSS.n5341 VSS 0.165082f
C13835 DVSS.n5342 VSS 0.165082f
C13836 DVSS.n5343 VSS 0.165082f
C13837 DVSS.n5344 VSS 0.165082f
C13838 DVSS.n5345 VSS 0.165082f
C13839 DVSS.n5346 VSS 0.165082f
C13840 DVSS.n5347 VSS 0.144737f
C13841 DVSS.n5349 VSS 0.082541f
C13842 DVSS.n5352 VSS 0.052308f
C13843 DVSS.n5353 VSS 0.082541f
C13844 DVSS.n5354 VSS 0.439557f
C13845 DVSS.n5355 VSS 0.439557f
C13846 DVSS.n5357 VSS 0.052308f
C13847 DVSS.n5360 VSS 0.052308f
C13848 DVSS.n5361 VSS 0.052308f
C13849 DVSS.n5363 VSS 0.052308f
C13850 DVSS.n5365 VSS 0.728095f
C13851 DVSS.n5366 VSS 0.082541f
C13852 DVSS.n5367 VSS 0.026154f
C13853 DVSS.n5368 VSS 0.026154f
C13854 DVSS.n5371 VSS 0.026154f
C13855 DVSS.n5372 VSS 0.026154f
C13856 DVSS.n5373 VSS 0.058114f
C13857 DVSS.n5375 VSS 0.026154f
C13858 DVSS.n5376 VSS 0.041971f
C13859 DVSS.n5377 VSS 0.026154f
C13860 DVSS.n5378 VSS 0.048967f
C13861 DVSS.n5379 VSS 0.331802f
C13862 DVSS.n5380 VSS 0.222771f
C13863 DVSS.n5381 VSS 0.026154f
C13864 DVSS.n5382 VSS 0.179185f
C13865 DVSS.n5383 VSS 0.09309f
C13866 DVSS.n5384 VSS 0.026154f
C13867 DVSS.n5385 VSS 0.335771f
C13868 DVSS.n5386 VSS 0.756156f
C13869 DVSS.n5387 VSS 0.242143f
C13870 DVSS.n5388 VSS 0.026154f
C13871 DVSS.n5389 VSS 0.066724f
C13872 DVSS.n5391 VSS 0.026154f
C13873 DVSS.n5392 VSS 0.026154f
C13874 DVSS.n5393 VSS 0.082541f
C13875 DVSS.n5394 VSS 0.728095f
C13876 DVSS.n5395 VSS 0.74307f
C13877 DVSS.n5397 VSS 0.052308f
C13878 DVSS.n5398 VSS 0.052308f
C13879 DVSS.n5402 VSS 0.066724f
C13880 DVSS.n5404 VSS 0.043865f
C13881 DVSS.n5406 VSS 0.038205f
C13882 DVSS.n5407 VSS 0.035873f
C13883 DVSS.n5408 VSS 0.038205f
C13884 DVSS.n5409 VSS 0.038205f
C13885 DVSS.n5410 VSS 0.038205f
C13886 DVSS.n5411 VSS 0.038205f
C13887 DVSS.n5412 VSS 0.035873f
C13888 DVSS.n5413 VSS 0.038205f
C13889 DVSS.n5414 VSS 0.038205f
C13890 DVSS.n5415 VSS 0.038205f
C13891 DVSS.n5416 VSS 0.038205f
C13892 DVSS.n5417 VSS 0.038205f
C13893 DVSS.n5418 VSS 0.035873f
C13894 DVSS.n5419 VSS 0.038205f
C13895 DVSS.n5420 VSS 0.038205f
C13896 DVSS.n5421 VSS 0.038205f
C13897 DVSS.n5422 VSS 0.038205f
C13898 DVSS.n5423 VSS 0.038205f
C13899 DVSS.n5424 VSS 0.026905f
C13900 DVSS.n5425 VSS 0.038205f
C13901 DVSS.t6 VSS 0.330478f
C13902 DVSS.n5426 VSS 0.125906f
C13903 DVSS.n5427 VSS 0.038205f
C13904 DVSS.n5428 VSS 0.038205f
C13905 DVSS.n5429 VSS 0.038205f
C13906 DVSS.n5430 VSS 0.038205f
C13907 DVSS.n5431 VSS 0.035873f
C13908 DVSS.n5432 VSS 0.038205f
C13909 DVSS.n5433 VSS 0.038205f
C13910 DVSS.n5434 VSS 0.038205f
C13911 DVSS.n5435 VSS 0.038205f
C13912 DVSS.n5436 VSS 0.038205f
C13913 DVSS.n5437 VSS 0.035873f
C13914 DVSS.n5438 VSS 0.038205f
C13915 DVSS.n5439 VSS 0.038205f
C13916 DVSS.n5440 VSS 0.038205f
C13917 DVSS.n5441 VSS 0.038205f
C13918 DVSS.n5442 VSS 0.038205f
C13919 DVSS.n5443 VSS 0.038205f
C13920 DVSS.n5444 VSS 0.035873f
C13921 DVSS.n5445 VSS 0.038205f
C13922 DVSS.n5446 VSS 0.038205f
C13923 DVSS.n5447 VSS 0.035873f
C13924 DVSS.n5448 VSS 0.035873f
C13925 DVSS.n5449 VSS 0.035873f
C13926 DVSS.n5450 VSS 0.038205f
C13927 DVSS.n5451 VSS 0.038205f
C13928 DVSS.n5452 VSS 0.038205f
C13929 DVSS.n5453 VSS 0.035873f
C13930 DVSS.n5454 VSS 0.035873f
C13931 DVSS.n5455 VSS 0.035873f
C13932 DVSS.n5456 VSS 0.038205f
C13933 DVSS.n5457 VSS 0.038205f
C13934 DVSS.n5458 VSS 0.038205f
C13935 DVSS.n5459 VSS 0.033714f
C13936 DVSS.n5460 VSS 0.020096f
C13937 DVSS.n5461 VSS 0.026905f
C13938 DVSS.n5462 VSS 0.038205f
C13939 DVSS.n5463 VSS 0.038205f
C13940 DVSS.n5464 VSS 0.038205f
C13941 DVSS.n5465 VSS 0.035873f
C13942 DVSS.n5466 VSS 0.035873f
C13943 DVSS.n5467 VSS 0.035873f
C13944 DVSS.n5468 VSS 0.038205f
C13945 DVSS.n5469 VSS 0.038205f
C13946 DVSS.n5470 VSS 0.038205f
C13947 DVSS.n5471 VSS 0.035873f
C13948 DVSS.n5472 VSS 0.035873f
C13949 DVSS.n5473 VSS 0.035873f
C13950 DVSS.n5474 VSS 0.038205f
C13951 DVSS.n5475 VSS 0.038205f
C13952 DVSS.n5476 VSS 0.038205f
C13953 DVSS.n5477 VSS 0.035873f
C13954 DVSS.n5478 VSS 0.035873f
C13955 DVSS.n5479 VSS 0.035873f
C13956 DVSS.n5480 VSS 0.038205f
C13957 DVSS.n5481 VSS 0.038205f
C13958 DVSS.n5482 VSS 0.066505f
C13959 DVSS.n5483 VSS 0.031887f
C13960 DVSS.n5484 VSS 0.066505f
C13961 DVSS.n5485 VSS 0.069335f
C13962 DVSS.n5487 VSS 0.066505f
C13963 DVSS.n5488 VSS 0.069335f
C13964 DVSS.n5490 VSS 0.043865f
C13965 DVSS.n5491 VSS 0.065379f
C13966 DVSS.n5493 VSS 0.043865f
C13967 DVSS.n5494 VSS 0.396845f
C13968 DVSS.n5496 VSS 0.186719f
C13969 DVSS.n5498 VSS 0.066724f
C13970 DVSS.n5499 VSS 0.052308f
C13971 DVSS.n5500 VSS 0.242143f
C13972 DVSS.n5501 VSS 0.756156f
C13973 DVSS.n5503 VSS 0.335771f
C13974 DVSS.n5505 VSS 0.066724f
C13975 DVSS.n5506 VSS 0.052308f
C13976 DVSS.n5507 VSS 0.09309f
C13977 DVSS.n5509 VSS 0.179185f
C13978 DVSS.n5513 VSS 0.066724f
C13979 DVSS.n5514 VSS 0.052308f
C13980 DVSS.n5515 VSS 0.222771f
C13981 DVSS.n5516 VSS 0.754249f
C13982 DVSS.n5518 VSS 0.066724f
C13983 DVSS.n5519 VSS 0.052308f
C13984 DVSS.n5521 VSS 0.133934f
C13985 DVSS.n5523 VSS 0.066724f
C13986 DVSS.n5524 VSS 0.052308f
C13987 DVSS.n5525 VSS 0.222771f
C13988 DVSS.n5526 VSS 0.754249f
C13989 DVSS.n5528 VSS 0.179185f
C13990 DVSS.n5530 VSS 0.133934f
C13991 DVSS.n5532 VSS 0.066724f
C13992 DVSS.n5533 VSS 0.052308f
C13993 DVSS.n5534 VSS 0.09309f
C13994 DVSS.n5535 VSS 0.754249f
C13995 DVSS.n5537 VSS 0.335771f
C13996 DVSS.n5538 VSS 0.756156f
C13997 DVSS.n5540 VSS 0.133934f
C13998 DVSS.n5542 VSS 0.066724f
C13999 DVSS.n5543 VSS 0.052308f
C14000 DVSS.n5544 VSS 0.242143f
C14001 DVSS.n5545 VSS 0.754249f
C14002 DVSS.n5547 VSS 0.186719f
C14003 DVSS.n5549 VSS 0.038205f
C14004 DVSS.n5550 VSS 0.035873f
C14005 DVSS.n5551 VSS 0.023878f
C14006 DVSS.n5552 VSS 0.021932f
C14007 DVSS.n5553 VSS 0.021932f
C14008 DVSS.n5554 VSS 0.021932f
C14009 DVSS.n5555 VSS 0.021932f
C14010 DVSS.n5556 VSS 0.021932f
C14011 DVSS.n5557 VSS 0.019279f
C14012 DVSS.n5558 VSS 0.021755f
C14013 DVSS.n5559 VSS 0.021932f
C14014 DVSS.n5560 VSS 0.021932f
C14015 DVSS.n5561 VSS 0.021932f
C14016 DVSS.n5562 VSS 0.021932f
C14017 DVSS.n5563 VSS 0.021932f
C14018 DVSS.n5564 VSS 0.021402f
C14019 DVSS.n5565 VSS 0.019633f
C14020 DVSS.n5566 VSS 0.021932f
C14021 DVSS.n5567 VSS 0.021932f
C14022 DVSS.n5568 VSS 0.021932f
C14023 DVSS.n5569 VSS 0.021932f
C14024 DVSS.n5570 VSS 0.021932f
C14025 DVSS.n5571 VSS 0.021932f
C14026 DVSS.n5572 VSS 0.020694f
C14027 DVSS.n5573 VSS 0.020341f
C14028 DVSS.n5574 VSS 0.021932f
C14029 DVSS.n5575 VSS 0.021932f
C14030 DVSS.n5576 VSS 0.021932f
C14031 DVSS.n5577 VSS 0.035873f
C14032 DVSS.n5578 VSS 0.021932f
C14033 DVSS.n5579 VSS 0.035873f
C14034 DVSS.n5580 VSS 0.035873f
C14035 DVSS.n5581 VSS 0.020341f
C14036 DVSS.n5582 VSS 0.020694f
C14037 DVSS.n5583 VSS 0.035873f
C14038 DVSS.n5584 VSS 0.021932f
C14039 DVSS.n5585 VSS 0.035873f
C14040 DVSS.n5586 VSS 0.021932f
C14041 DVSS.n5587 VSS 0.035873f
C14042 DVSS.n5588 VSS 0.021932f
C14043 DVSS.n5589 VSS 0.035873f
C14044 DVSS.n5590 VSS 0.021932f
C14045 DVSS.n5591 VSS 0.035873f
C14046 DVSS.n5592 VSS 0.021932f
C14047 DVSS.n5593 VSS 0.035873f
C14048 DVSS.n5594 VSS 0.021932f
C14049 DVSS.n5595 VSS 0.035873f
C14050 DVSS.n5596 VSS 0.033714f
C14051 DVSS.n5597 VSS 0.019633f
C14052 DVSS.n5598 VSS 0.021402f
C14053 DVSS.n5599 VSS 0.020096f
C14054 DVSS.n5600 VSS 0.021932f
C14055 DVSS.n5601 VSS 0.026905f
C14056 DVSS.t12 VSS 0.330478f
C14057 DVSS.n5602 VSS 0.125906f
C14058 DVSS.n5603 VSS 0.021932f
C14059 DVSS.n5604 VSS 0.026905f
C14060 DVSS.n5605 VSS 0.021932f
C14061 DVSS.n5606 VSS 0.035873f
C14062 DVSS.n5607 VSS 0.021932f
C14063 DVSS.n5608 VSS 0.035873f
C14064 DVSS.n5609 VSS 0.021932f
C14065 DVSS.n5610 VSS 0.035873f
C14066 DVSS.n5611 VSS 0.035873f
C14067 DVSS.n5612 VSS 0.021755f
C14068 DVSS.n5613 VSS 0.019279f
C14069 DVSS.n5614 VSS 0.035873f
C14070 DVSS.n5615 VSS 0.021932f
C14071 DVSS.n5616 VSS 0.035873f
C14072 DVSS.n5617 VSS 0.021932f
C14073 DVSS.n5618 VSS 0.035873f
C14074 DVSS.n5619 VSS 0.021932f
C14075 DVSS.n5620 VSS 0.035873f
C14076 DVSS.n5621 VSS 0.021932f
C14077 DVSS.n5622 VSS 0.035873f
C14078 DVSS.n5623 VSS 0.021932f
C14079 DVSS.n5624 VSS 0.035873f
C14080 DVSS.n5625 VSS 0.035873f
C14081 DVSS.n5626 VSS 0.023878f
C14082 DVSS.n5627 VSS 0.038205f
C14083 DVSS.n5628 VSS 0.066505f
C14084 DVSS.n5629 VSS 0.031887f
C14085 DVSS.n5630 VSS 0.066505f
C14086 DVSS.n5631 VSS 0.069335f
C14087 DVSS.n5633 VSS 0.065379f
C14088 DVSS.n5635 VSS 0.043865f
C14089 DVSS.n5636 VSS 0.396845f
C14090 DVSS.n5638 VSS 0.069335f
C14091 DVSS.n5639 VSS 0.066505f
C14092 DVSS.n5640 VSS 0.049824f
C14093 DVSS.n5641 VSS 0.066505f
C14094 DVSS.n5642 VSS 0.069335f
C14095 DVSS.n5644 VSS 0.043865f
C14096 DVSS.n5645 VSS 0.396845f
C14097 DVSS.n5647 VSS 0.133934f
C14098 DVSS.n5649 VSS 0.066724f
C14099 DVSS.n5650 VSS 0.052308f
C14100 DVSS.n5651 VSS 0.186719f
C14101 DVSS.n5652 VSS 0.754249f
C14102 DVSS.n5654 VSS 0.242143f
C14103 DVSS.n5655 VSS 0.756156f
C14104 DVSS.n5657 VSS 0.133934f
C14105 DVSS.n5659 VSS 0.066724f
C14106 DVSS.n5660 VSS 0.052308f
C14107 DVSS.n5661 VSS 0.335771f
C14108 DVSS.n5662 VSS 0.754249f
C14109 DVSS.n5664 VSS 0.09309f
C14110 DVSS.n5665 VSS 0.2147f
C14111 DVSS.n5666 VSS 0.010297f
C14112 DVSS.n5667 VSS 0.088337f
C14113 DVSS.n5668 VSS 0.253981f
C14114 DVSS.n5669 VSS 0.020594f
C14115 DVSS.n5670 VSS 0.296948f
C14116 DVSS.n5671 VSS 0.296948f
C14117 DVSS.t7 VSS 0.394423f
C14118 DVSS.n5672 VSS 0.32373f
C14119 DVSS.n5673 VSS 0.010297f
C14120 DVSS.n5674 VSS 0.2147f
C14121 DVSS.n5675 VSS 0.010297f
C14122 DVSS.n5676 VSS 0.020594f
C14123 DVSS.n5677 VSS 0.253981f
C14124 DVSS.n5679 VSS 0.09309f
C14125 DVSS.n5681 VSS 0.066724f
C14126 DVSS.n5682 VSS 0.052308f
C14127 DVSS.n5683 VSS 0.335771f
C14128 DVSS.n5684 VSS 0.756156f
C14129 DVSS.n5686 VSS 0.242143f
C14130 DVSS.n5688 VSS 0.066724f
C14131 DVSS.n5689 VSS 0.052308f
C14132 DVSS.n5690 VSS 0.186719f
C14133 DVSS.n5691 VSS 0.396845f
C14134 DVSS.n5693 VSS 0.043865f
C14135 DVSS.n5694 VSS 0.065379f
C14136 DVSS.n5696 VSS 0.069335f
C14137 DVSS.n5697 VSS 0.066505f
C14138 DVSS.n5698 VSS 0.038205f
C14139 DVSS.n5699 VSS 0.035873f
C14140 DVSS.n5700 VSS 0.035873f
C14141 DVSS.n5701 VSS 0.035873f
C14142 DVSS.n5702 VSS 0.038205f
C14143 DVSS.n5703 VSS 0.038205f
C14144 DVSS.n5704 VSS 0.038205f
C14145 DVSS.n5705 VSS 0.035873f
C14146 DVSS.n5706 VSS 0.035873f
C14147 DVSS.n5707 VSS 0.035873f
C14148 DVSS.n5708 VSS 0.038205f
C14149 DVSS.n5709 VSS 0.038205f
C14150 DVSS.n5710 VSS 0.038205f
C14151 DVSS.n5711 VSS 0.035873f
C14152 DVSS.n5712 VSS 0.035873f
C14153 DVSS.n5713 VSS 0.033714f
C14154 DVSS.n5714 VSS 0.038205f
C14155 DVSS.n5715 VSS 0.038205f
C14156 DVSS.n5716 VSS 0.038205f
C14157 DVSS.n5717 VSS 0.026905f
C14158 DVSS.t14 VSS 0.330478f
C14159 DVSS.n5718 VSS 0.125906f
C14160 DVSS.n5719 VSS 0.026905f
C14161 DVSS.n5720 VSS 0.035873f
C14162 DVSS.n5721 VSS 0.038205f
C14163 DVSS.n5722 VSS 0.038205f
C14164 DVSS.n5723 VSS 0.038205f
C14165 DVSS.n5724 VSS 0.035873f
C14166 DVSS.n5725 VSS 0.035873f
C14167 DVSS.n5726 VSS 0.035873f
C14168 DVSS.n5727 VSS 0.038205f
C14169 DVSS.n5728 VSS 0.038205f
C14170 DVSS.n5729 VSS 0.038205f
C14171 DVSS.n5730 VSS 0.035873f
C14172 DVSS.n5731 VSS 0.035873f
C14173 DVSS.n5732 VSS 0.035873f
C14174 DVSS.n5733 VSS 0.038205f
C14175 DVSS.n5734 VSS 0.038205f
C14176 DVSS.n5735 VSS 0.038205f
C14177 DVSS.n5736 VSS 0.035873f
C14178 DVSS.n5737 VSS 0.035873f
C14179 DVSS.n5738 VSS 0.031887f
C14180 DVSS.n5739 VSS 0.05713f
C14181 DVSS.n5740 VSS 0.047402f
C14182 DVSS.n5741 VSS 0.082541f
C14183 DVSS.n5742 VSS 0.072078f
C14184 DVSS.n5743 VSS 0.165082f
C14185 DVSS.n5744 VSS 0.165082f
C14186 DVSS.n5745 VSS 0.165082f
C14187 DVSS.n5746 VSS 0.165082f
C14188 DVSS.n5747 VSS 0.165082f
C14189 DVSS.n5748 VSS 0.159269f
C14190 DVSS.n5749 VSS 0.165082f
C14191 DVSS.n5750 VSS 0.165082f
C14192 DVSS.n5751 VSS 0.165082f
C14193 DVSS.n5752 VSS 0.165082f
C14194 DVSS.n5753 VSS 0.165082f
C14195 DVSS.n5754 VSS 0.165082f
C14196 DVSS.n5755 VSS 0.165082f
C14197 DVSS.n5756 VSS 0.165082f
C14198 DVSS.n5757 VSS 0.165082f
C14199 DVSS.n5758 VSS 0.165082f
C14200 DVSS.n5759 VSS 0.165082f
C14201 DVSS.n5760 VSS 0.165082f
C14202 DVSS.n5761 VSS 0.165082f
C14203 DVSS.n5762 VSS 0.165082f
C14204 DVSS.n5763 VSS 0.165082f
C14205 DVSS.n5764 VSS 0.165082f
C14206 DVSS.n5765 VSS 0.165082f
C14207 DVSS.n5766 VSS 0.165082f
C14208 DVSS.n5767 VSS 0.165082f
C14209 DVSS.n5768 VSS 0.165082f
C14210 DVSS.n5769 VSS 0.165082f
C14211 DVSS.n5770 VSS 0.165082f
C14212 DVSS.n5771 VSS 0.165082f
C14213 DVSS.n5772 VSS 0.131949f
C14214 DVSS.n5775 VSS 0.082541f
C14215 DVSS.n5776 VSS 0.728095f
C14216 DVSS.n5777 VSS 0.082541f
C14217 DVSS.n5778 VSS 0.072078f
C14218 DVSS.n5779 VSS 0.165082f
C14219 DVSS.n5780 VSS 0.165082f
C14220 DVSS.n5781 VSS 0.165082f
C14221 DVSS.n5782 VSS 0.165082f
C14222 DVSS.n5783 VSS 0.165082f
C14223 DVSS.n5784 VSS 0.147063f
C14224 DVSS.n5785 VSS 0.165082f
C14225 DVSS.n5786 VSS 0.165082f
C14226 DVSS.n5787 VSS 0.165082f
C14227 DVSS.n5788 VSS 0.165082f
C14228 DVSS.n5789 VSS 0.165082f
C14229 DVSS.n5790 VSS 0.165082f
C14230 DVSS.n5791 VSS 0.165082f
C14231 DVSS.n5792 VSS 0.165082f
C14232 DVSS.n5793 VSS 0.165082f
C14233 DVSS.n5794 VSS 0.165082f
C14234 DVSS.n5795 VSS 0.165082f
C14235 DVSS.n5796 VSS 0.165082f
C14236 DVSS.n5797 VSS 0.165082f
C14237 DVSS.n5798 VSS 0.165082f
C14238 DVSS.n5799 VSS 0.165082f
C14239 DVSS.n5800 VSS 0.165082f
C14240 DVSS.n5801 VSS 0.165082f
C14241 DVSS.n5802 VSS 0.165082f
C14242 DVSS.n5803 VSS 0.165082f
C14243 DVSS.n5804 VSS 0.165082f
C14244 DVSS.n5805 VSS 0.165082f
C14245 DVSS.n5806 VSS 0.165082f
C14246 DVSS.n5807 VSS 0.165082f
C14247 DVSS.n5808 VSS 0.131949f
C14248 DVSS.n5811 VSS 0.082541f
C14249 DVSS.n5812 VSS 0.728095f
C14250 DVSS.n5813 VSS 0.082541f
C14251 DVSS.n5814 VSS 0.147063f
C14252 DVSS.n5815 VSS 0.165082f
C14253 DVSS.n5816 VSS 0.165082f
C14254 DVSS.n5817 VSS 0.165082f
C14255 DVSS.n5818 VSS 0.165082f
C14256 DVSS.n5819 VSS 0.165082f
C14257 DVSS.n5820 VSS 0.165082f
C14258 DVSS.n5821 VSS 0.165082f
C14259 DVSS.n5822 VSS 0.165082f
C14260 DVSS.n5823 VSS 0.165082f
C14261 DVSS.n5824 VSS 0.165082f
C14262 DVSS.n5825 VSS 0.165082f
C14263 DVSS.n5826 VSS 0.165082f
C14264 DVSS.n5827 VSS 0.165082f
C14265 DVSS.n5828 VSS 0.128462f
C14266 DVSS.n5829 VSS 0.082541f
C14267 DVSS.n5830 VSS 0.286652f
C14268 DVSS.n5831 VSS 0.082541f
C14269 DVSS.n5832 VSS 0.173054f
C14270 DVSS.n5833 VSS 0.173054f
C14271 DVSS.n5834 VSS 0.082541f
C14272 DVSS.n5835 VSS 0.010297f
C14273 DVSS.n5836 VSS 0.01503f
C14274 DVSS.n5837 VSS 0.082541f
C14275 DVSS.n5838 VSS 0.129624f
C14276 DVSS.n5839 VSS 0.165082f
C14277 DVSS.n5840 VSS 0.165082f
C14278 DVSS.n5841 VSS 0.165082f
C14279 DVSS.n5842 VSS 0.165082f
C14280 DVSS.n5843 VSS 0.165082f
C14281 DVSS.n5844 VSS 0.165082f
C14282 DVSS.n5845 VSS 0.165082f
C14283 DVSS.n5846 VSS 0.131949f
C14284 DVSS.n5847 VSS 0.165082f
C14285 DVSS.n5848 VSS 0.165082f
C14286 DVSS.n5849 VSS 0.165082f
C14287 DVSS.n5850 VSS 0.611712f
C14288 DVSS.n5851 VSS 0.072078f
C14289 DVSS.n5852 VSS 0.165082f
C14290 DVSS.n5853 VSS 0.165082f
C14291 DVSS.n5854 VSS 0.072078f
C14292 DVSS.n5855 VSS 0.022779f
C14293 DVSS.n5858 VSS 0.052308f
C14294 DVSS.n5861 VSS 0.052308f
C14295 DVSS.n5863 VSS 0.439557f
C14296 DVSS.n5864 VSS 0.361112f
C14297 DVSS.n5865 VSS 0.022779f
C14298 DVSS.n5866 VSS 0.026154f
C14299 DVSS.n5867 VSS 0.048967f
C14300 DVSS.n5868 VSS 0.026154f
C14301 DVSS.n5869 VSS 0.041971f
C14302 DVSS.n5870 VSS 0.21755f
C14303 DVSS.n5871 VSS 0.21755f
C14304 DVSS.n5873 VSS 0.026154f
C14305 DVSS.n5875 VSS 0.026154f
C14306 DVSS.n5876 VSS 0.041971f
C14307 DVSS.n5877 VSS 0.026154f
C14308 DVSS.n5878 VSS 0.022779f
C14309 DVSS.n5879 VSS 0.361112f
C14310 DVSS.n5880 VSS 0.741594f
C14311 DVSS.n5881 VSS 0.746445f
C14312 DVSS.n5883 VSS 0.058114f
C14313 DVSS.n5884 VSS 0.045559f
C14314 DVSS.n5885 VSS 0.045559f
C14315 DVSS.n5887 VSS 0.045559f
C14316 DVSS.n5889 VSS 0.041971f
C14317 DVSS.n5890 VSS 0.764373f
C14318 DVSS.n5891 VSS 0.764373f
C14319 DVSS.n5893 VSS 0.048967f
C14320 DVSS.n5894 VSS 0.137309f
C14321 DVSS.n5895 VSS 0.041971f
C14322 DVSS.n5896 VSS 0.170965f
C14323 DVSS.n5897 VSS -1.23794f
C14324 DVSS.n5898 VSS 22.0306f
C14325 DVSS.n5899 VSS -1.23794f
C14326 DVSS.n5900 VSS 0.170965f
C14327 DVSS.n5901 VSS 0.137309f
C14328 DVSS.n5902 VSS 0.041971f
C14329 DVSS.n5903 VSS 0.045559f
C14330 DVSS.n5904 VSS 0.048967f
C14331 DVSS.n5905 VSS 0.764373f
C14332 DVSS.n5906 VSS 0.764373f
C14333 DVSS.n5907 VSS 0.041971f
C14334 DVSS.n5908 VSS 0.045559f
C14335 DVSS.n5909 VSS 0.048967f
C14336 DVSS.n5910 VSS 0.746445f
C14337 DVSS.n5911 VSS 0.741594f
C14338 DVSS.n5912 VSS 0.082541f
C14339 DVSS.n5913 VSS 0.439557f
C14340 DVSS.n5914 VSS 0.439557f
C14341 DVSS.n5915 VSS 0.082541f
C14342 DVSS.n5916 VSS 0.022779f
C14343 DVSS.n5917 VSS 0.026154f
C14344 DVSS.n5918 VSS 0.048967f
C14345 DVSS.n5919 VSS 0.026154f
C14346 DVSS.n5920 VSS 0.041971f
C14347 DVSS.n5921 VSS 0.21755f
C14348 DVSS.n5922 VSS 0.217854f
C14349 DVSS.n5923 VSS 0.133296f
C14350 DVSS.n5924 VSS 0.026154f
C14351 DVSS.n5925 VSS 0.032106f
C14352 DVSS.n5927 VSS 0.127236f
C14353 DVSS.n5928 VSS 0.026154f
C14354 DVSS.n5930 VSS 0.075348f
C14355 DVSS.n5934 VSS 0.148574f
C14356 DVSS.n5935 VSS 0.562685f
C14357 DVSS.n5936 VSS 0.291346f
C14358 DVSS.n5937 VSS 0.065797f
C14359 DVSS.n5938 VSS 0.150696f
C14360 DVSS.n5939 VSS 0.150696f
C14361 DVSS.n5940 VSS 0.065797f
C14362 DVSS.n5941 VSS 0.075348f
C14363 DVSS.n5942 VSS 0.022779f
C14364 DVSS.n5943 VSS 0.075348f
C14365 DVSS.n5944 VSS 0.062083f
C14366 DVSS.n5945 VSS 0.090206f
C14367 DVSS.n5946 VSS 0.135839f
C14368 DVSS.n5947 VSS 0.150696f
C14369 DVSS.n5948 VSS 0.150696f
C14370 DVSS.n5949 VSS 0.150696f
C14371 DVSS.n5950 VSS 0.132125f
C14372 DVSS.n5951 VSS 0.150696f
C14373 DVSS.n5952 VSS 0.065797f
C14374 DVSS.n5953 VSS 0.150696f
C14375 DVSS.n5954 VSS 0.150696f
C14376 DVSS.n5955 VSS 0.065797f
C14377 DVSS.n5958 VSS 0.075348f
C14378 DVSS.n5959 VSS 0.022779f
C14379 DVSS.n5960 VSS 0.075348f
C14380 DVSS.n5961 VSS 0.122573f
C14381 DVSS.n5962 VSS 0.150696f
C14382 DVSS.n5963 VSS 0.150696f
C14383 DVSS.n5964 VSS 0.150696f
C14384 DVSS.n5965 VSS 0.150696f
C14385 DVSS.n5966 VSS 0.150696f
C14386 DVSS.n5967 VSS 0.132125f
C14387 DVSS.n5968 VSS 0.150696f
C14388 DVSS.n5969 VSS 0.065797f
C14389 DVSS.n5970 VSS 0.150696f
C14390 DVSS.n5971 VSS 0.150696f
C14391 DVSS.n5972 VSS 0.065797f
C14392 DVSS.n5973 VSS 0.075348f
C14393 DVSS.n5974 VSS 0.022779f
C14394 DVSS.n5975 VSS 0.075348f
C14395 DVSS.n5976 VSS 0.122573f
C14396 DVSS.n5977 VSS 0.150696f
C14397 DVSS.n5978 VSS 0.150696f
C14398 DVSS.n5979 VSS 0.150696f
C14399 DVSS.n5980 VSS 0.150696f
C14400 DVSS.n5981 VSS 0.150696f
C14401 DVSS.n5982 VSS 0.150696f
C14402 DVSS.n5983 VSS 0.150696f
C14403 DVSS.n5984 VSS 0.150696f
C14404 DVSS.n5985 VSS 0.150696f
C14405 DVSS.n5986 VSS 0.150696f
C14406 DVSS.n5987 VSS 0.150696f
C14407 DVSS.n5988 VSS 0.150696f
C14408 DVSS.n5989 VSS 0.150696f
C14409 DVSS.n5990 VSS 0.150696f
C14410 DVSS.n5991 VSS 0.150696f
C14411 DVSS.n5992 VSS 0.150696f
C14412 DVSS.n5993 VSS 0.150696f
C14413 DVSS.n5994 VSS 0.132125f
C14414 DVSS.n5995 VSS 0.150696f
C14415 DVSS.n5996 VSS 0.065797f
C14416 DVSS.n5997 VSS 0.150696f
C14417 DVSS.n5998 VSS 0.150696f
C14418 DVSS.n5999 VSS 0.065797f
C14419 DVSS.n6000 VSS 0.075348f
C14420 DVSS.n6002 VSS 0.052308f
C14421 DVSS.n6003 VSS 0.075348f
C14422 DVSS.n6004 VSS 0.041129f
C14423 DVSS.n6005 VSS 0.026154f
C14424 DVSS.n6006 VSS 0.289551f
C14425 DVSS.n6007 VSS 0.026154f
C14426 DVSS.n6008 VSS 0.291484f
C14427 DVSS.n6009 VSS 0.291484f
C14428 DVSS.n6010 VSS 0.021932f
C14429 DVSS.n6011 VSS 0.028093f
C14430 DVSS.n6012 VSS -0.499142f
C14431 DVSS.n6013 VSS 26.9724f
C14432 DVSS.n6014 VSS 8.5528f
C14433 DVSS.n6015 VSS 4.16152f
C14434 DVSS.n6016 VSS 1.22586f
C14435 DVSS.n6017 VSS 1.48043f
C14436 DVSS.n6018 VSS 0.310331f
C14437 DVSS.n6019 VSS 0.165082f
C14438 DVSS.n6020 VSS 0.165082f
C14439 DVSS.n6021 VSS 0.165082f
C14440 DVSS.n6022 VSS 0.165082f
C14441 DVSS.n6023 VSS 0.165082f
C14442 DVSS.n6024 VSS 0.165082f
C14443 DVSS.n6025 VSS 0.165082f
C14444 DVSS.n6026 VSS 0.165082f
C14445 DVSS.n6027 VSS 0.165082f
C14446 DVSS.n6028 VSS 0.105392f
C14447 DVSS.n6029 VSS 0.165082f
C14448 DVSS.n6030 VSS 0.165082f
C14449 DVSS.n6031 VSS 0.165082f
C14450 DVSS.n6032 VSS 0.072078f
C14451 DVSS.n6033 VSS 0.105506f
C14452 DVSS.n6034 VSS 0.143575f
C14453 DVSS.n6035 VSS 0.165082f
C14454 DVSS.n6036 VSS 0.165082f
C14455 DVSS.n6037 VSS 0.165082f
C14456 DVSS.n6038 VSS 0.165082f
C14457 DVSS.n6039 VSS 0.165082f
C14458 DVSS.n6040 VSS 0.165082f
C14459 DVSS.n6041 VSS 0.165082f
C14460 DVSS.n6042 VSS 0.165082f
C14461 DVSS.n6043 VSS 0.165082f
C14462 DVSS.n6044 VSS 0.165082f
C14463 DVSS.n6045 VSS 0.336866f
C14464 DVSS.n6046 VSS 0.165082f
C14465 DVSS.n6047 VSS 0.165082f
C14466 DVSS.n6048 VSS 0.310331f
C14467 DVSS.n6049 VSS 0.611712f
C14468 DVSS.n6050 VSS 0.165082f
C14469 DVSS.n6051 VSS 0.165082f
C14470 DVSS.n6052 VSS 0.165082f
C14471 DVSS.n6053 VSS 0.165082f
C14472 DVSS.n6054 VSS 0.165082f
C14473 DVSS.n6055 VSS 0.165082f
C14474 DVSS.n6056 VSS 0.165082f
C14475 DVSS.n6057 VSS 0.165082f
C14476 DVSS.n6058 VSS 0.165082f
C14477 DVSS.n6059 VSS 0.165082f
C14478 DVSS.n6060 VSS 0.165082f
C14479 DVSS.n6061 VSS 0.165082f
C14480 DVSS.n6062 VSS 0.165082f
C14481 DVSS.n6063 VSS 0.165082f
C14482 DVSS.n6064 VSS 0.165082f
C14483 DVSS.n6065 VSS 0.165082f
C14484 DVSS.n6066 VSS 0.165082f
C14485 DVSS.n6067 VSS 0.165082f
C14486 DVSS.n6068 VSS 0.114511f
C14487 DVSS.n6069 VSS 0.165082f
C14488 DVSS.n6070 VSS 0.165082f
C14489 DVSS.n6071 VSS 0.165082f
C14490 DVSS.n6072 VSS 0.165082f
C14491 DVSS.n6073 VSS 0.165082f
C14492 DVSS.n6074 VSS 0.165082f
C14493 DVSS.n6075 VSS 0.165082f
C14494 DVSS.n6076 VSS 0.165082f
C14495 DVSS.n6077 VSS 0.165082f
C14496 DVSS.n6078 VSS 0.165082f
C14497 DVSS.n6079 VSS 0.165082f
C14498 DVSS.n6080 VSS 0.165082f
C14499 DVSS.n6081 VSS 0.165082f
C14500 DVSS.n6082 VSS 0.165082f
C14501 DVSS.n6083 VSS 0.165082f
C14502 DVSS.n6084 VSS 0.165082f
C14503 DVSS.n6085 VSS 0.165082f
C14504 DVSS.n6086 VSS 0.165082f
C14505 DVSS.n6087 VSS 0.165082f
C14506 DVSS.n6088 VSS 0.165082f
C14507 DVSS.n6089 VSS 0.165082f
C14508 DVSS.n6090 VSS 0.165082f
C14509 DVSS.n6091 VSS 0.165082f
C14510 DVSS.n6092 VSS 0.165082f
C14511 DVSS.n6093 VSS 0.165082f
C14512 DVSS.n6094 VSS 0.165082f
C14513 DVSS.n6095 VSS 0.165082f
C14514 DVSS.n6096 VSS 0.165082f
C14515 DVSS.n6097 VSS 0.165082f
C14516 DVSS.n6098 VSS 0.165082f
C14517 DVSS.n6099 VSS 0.165082f
C14518 DVSS.n6100 VSS 0.165082f
C14519 DVSS.n6101 VSS 0.165082f
C14520 DVSS.n6102 VSS 0.165082f
C14521 DVSS.n6103 VSS 0.165082f
C14522 DVSS.n6104 VSS 0.165082f
C14523 DVSS.n6105 VSS 0.165082f
C14524 DVSS.n6106 VSS 0.165082f
C14525 DVSS.n6107 VSS 0.165082f
C14526 DVSS.n6108 VSS 0.165082f
C14527 DVSS.n6109 VSS 0.165082f
C14528 DVSS.n6110 VSS 0.165082f
C14529 DVSS.n6111 VSS 0.165082f
C14530 DVSS.n6112 VSS 0.165082f
C14531 DVSS.n6113 VSS 0.165082f
C14532 DVSS.n6114 VSS 0.165082f
C14533 DVSS.n6115 VSS 0.165082f
C14534 DVSS.n6116 VSS 0.165082f
C14535 DVSS.n6117 VSS 0.165082f
C14536 DVSS.n6118 VSS 0.165082f
C14537 DVSS.n6119 VSS 0.165082f
C14538 DVSS.n6120 VSS 0.165082f
C14539 DVSS.n6121 VSS 0.165082f
C14540 DVSS.n6122 VSS 0.165082f
C14541 DVSS.n6123 VSS 0.165082f
C14542 DVSS.n6124 VSS 0.165082f
C14543 DVSS.n6125 VSS 0.165082f
C14544 DVSS.n6126 VSS 0.165082f
C14545 DVSS.n6127 VSS 0.165082f
C14546 DVSS.n6128 VSS 0.165082f
C14547 DVSS.n6129 VSS 0.165082f
C14548 DVSS.n6130 VSS 0.165082f
C14549 DVSS.n6131 VSS 0.165082f
C14550 DVSS.n6132 VSS 0.165082f
C14551 DVSS.n6133 VSS 0.165082f
C14552 DVSS.n6134 VSS 0.165082f
C14553 DVSS.n6135 VSS 0.165082f
C14554 DVSS.n6136 VSS 0.165082f
C14555 DVSS.n6137 VSS 0.165082f
C14556 DVSS.n6138 VSS 0.165082f
C14557 DVSS.n6139 VSS 0.165082f
C14558 DVSS.n6140 VSS 0.165082f
C14559 DVSS.n6141 VSS 0.165082f
C14560 DVSS.n6142 VSS 0.165082f
C14561 DVSS.n6143 VSS 0.165082f
C14562 DVSS.n6144 VSS 0.165082f
C14563 DVSS.n6145 VSS 0.165082f
C14564 DVSS.n6146 VSS 0.165082f
C14565 DVSS.n6147 VSS 0.165082f
C14566 DVSS.n6148 VSS 0.165082f
C14567 DVSS.n6149 VSS 0.165082f
C14568 DVSS.n6150 VSS 0.165082f
C14569 DVSS.n6151 VSS 0.165082f
C14570 DVSS.n6152 VSS 0.148806f
C14571 DVSS.n6153 VSS 0.165082f
C14572 DVSS.n6154 VSS 0.165082f
C14573 DVSS.n6155 VSS 0.315112f
C14574 DVSS.n6156 VSS 0.165082f
C14575 DVSS.n6157 VSS 1.84499f
C14576 DVSS.n6158 VSS 1.48464f
C14577 DVSS.n6159 VSS 0.341473f
C14578 DVSS.n6160 VSS 0.165082f
C14579 DVSS.n6161 VSS 0.165082f
C14580 DVSS.n6162 VSS 0.165082f
C14581 DVSS.n6163 VSS 0.616179f
C14582 DVSS.n6164 VSS 0.162757f
C14583 DVSS.n6165 VSS 0.084866f
C14584 DVSS.n6166 VSS 0.098817f
C14585 DVSS.n6167 VSS 0.098817f
C14586 DVSS.n6168 VSS 0.148806f
C14587 DVSS.n6169 VSS 0.165082f
C14588 DVSS.n6170 VSS 0.165082f
C14589 DVSS.n6171 VSS 0.165082f
C14590 DVSS.n6172 VSS 0.165082f
C14591 DVSS.n6173 VSS 0.165082f
C14592 DVSS.n6174 VSS 0.165082f
C14593 DVSS.n6175 VSS 0.165082f
C14594 DVSS.n6176 VSS 0.165082f
C14595 DVSS.n6177 VSS 0.165082f
C14596 DVSS.n6178 VSS 0.165082f
C14597 DVSS.n6179 VSS 0.165082f
C14598 DVSS.n6180 VSS 0.165082f
C14599 DVSS.n6181 VSS 0.165082f
C14600 DVSS.n6182 VSS 0.165082f
C14601 DVSS.n6183 VSS 0.165082f
C14602 DVSS.n6184 VSS 0.165082f
C14603 DVSS.n6185 VSS 0.165082f
C14604 DVSS.n6186 VSS 0.165082f
C14605 DVSS.n6187 VSS 0.165082f
C14606 DVSS.n6188 VSS 0.165082f
C14607 DVSS.n6189 VSS 0.165082f
C14608 DVSS.n6190 VSS 0.165082f
C14609 DVSS.n6191 VSS 0.165082f
C14610 DVSS.n6192 VSS 0.165082f
C14611 DVSS.n6193 VSS 0.165082f
C14612 DVSS.n6194 VSS 0.165082f
C14613 DVSS.n6195 VSS 0.165082f
C14614 DVSS.n6196 VSS 0.165082f
C14615 DVSS.n6197 VSS 0.165082f
C14616 DVSS.n6198 VSS 0.165082f
C14617 DVSS.n6199 VSS 0.165082f
C14618 DVSS.n6200 VSS 0.165082f
C14619 DVSS.n6201 VSS 0.165082f
C14620 DVSS.n6202 VSS 0.165082f
C14621 DVSS.n6203 VSS 0.165082f
C14622 DVSS.n6204 VSS 0.165082f
C14623 DVSS.n6205 VSS 0.165082f
C14624 DVSS.n6206 VSS 0.165082f
C14625 DVSS.n6207 VSS 0.165082f
C14626 DVSS.n6208 VSS 0.165082f
C14627 DVSS.n6209 VSS 0.165082f
C14628 DVSS.n6210 VSS 0.165082f
C14629 DVSS.n6211 VSS 0.165082f
C14630 DVSS.n6212 VSS 0.165082f
C14631 DVSS.n6213 VSS 0.165082f
C14632 DVSS.n6214 VSS 0.165082f
C14633 DVSS.n6215 VSS 0.165082f
C14634 DVSS.n6216 VSS 0.165082f
C14635 DVSS.n6217 VSS 0.165082f
C14636 DVSS.n6218 VSS 0.165082f
C14637 DVSS.n6219 VSS 0.165082f
C14638 DVSS.n6220 VSS 0.165082f
C14639 DVSS.n6221 VSS 0.165082f
C14640 DVSS.n6222 VSS 0.165082f
C14641 DVSS.n6223 VSS 0.165082f
C14642 DVSS.n6224 VSS 0.165082f
C14643 DVSS.n6225 VSS 0.165082f
C14644 DVSS.n6226 VSS 0.165082f
C14645 DVSS.n6227 VSS 0.165082f
C14646 DVSS.n6228 VSS 0.165082f
C14647 DVSS.n6229 VSS 0.165082f
C14648 DVSS.n6230 VSS 0.165082f
C14649 DVSS.n6231 VSS 0.165082f
C14650 DVSS.n6232 VSS 0.165082f
C14651 DVSS.n6233 VSS 0.165082f
C14652 DVSS.n6234 VSS 0.165082f
C14653 DVSS.n6235 VSS 0.165082f
C14654 DVSS.n6236 VSS 0.165082f
C14655 DVSS.n6237 VSS 0.165082f
C14656 DVSS.n6238 VSS 0.165082f
C14657 DVSS.n6239 VSS 0.165082f
C14658 DVSS.n6240 VSS 0.165082f
C14659 DVSS.n6241 VSS 0.165082f
C14660 DVSS.n6242 VSS 0.165082f
C14661 DVSS.n6243 VSS 0.165082f
C14662 DVSS.n6244 VSS 0.165082f
C14663 DVSS.n6245 VSS 0.165082f
C14664 DVSS.n6246 VSS 0.165082f
C14665 DVSS.n6247 VSS 0.165082f
C14666 DVSS.n6248 VSS 0.165082f
C14667 DVSS.n6249 VSS 0.165082f
C14668 DVSS.n6250 VSS 0.165082f
C14669 DVSS.n6251 VSS 0.165082f
C14670 DVSS.n6252 VSS 0.165082f
C14671 DVSS.n6253 VSS 0.165082f
C14672 DVSS.n6254 VSS 0.165082f
C14673 DVSS.n6255 VSS 0.165082f
C14674 DVSS.n6256 VSS 0.165082f
C14675 DVSS.n6257 VSS 0.165082f
C14676 DVSS.n6258 VSS 0.165082f
C14677 DVSS.n6259 VSS 0.165082f
C14678 DVSS.n6260 VSS 0.165082f
C14679 DVSS.n6261 VSS 0.165082f
C14680 DVSS.n6262 VSS 0.165082f
C14681 DVSS.n6263 VSS 0.165082f
C14682 DVSS.n6264 VSS 0.165082f
C14683 DVSS.n6265 VSS 0.165082f
C14684 DVSS.n6266 VSS 0.165082f
C14685 DVSS.n6267 VSS 0.165082f
C14686 DVSS.n6268 VSS 0.165082f
C14687 DVSS.n6269 VSS 0.165082f
C14688 DVSS.n6270 VSS 0.165082f
C14689 DVSS.n6271 VSS 0.165082f
C14690 DVSS.n6272 VSS 0.165082f
C14691 DVSS.n6273 VSS 0.165082f
C14692 DVSS.n6274 VSS 0.165082f
C14693 DVSS.n6275 VSS 0.165082f
C14694 DVSS.n6276 VSS 0.165082f
C14695 DVSS.n6277 VSS 0.165082f
C14696 DVSS.n6278 VSS 0.165082f
C14697 DVSS.n6279 VSS 0.165082f
C14698 DVSS.n6280 VSS 0.165082f
C14699 DVSS.n6281 VSS 0.165082f
C14700 DVSS.n6282 VSS 0.165082f
C14701 DVSS.n6283 VSS 0.165082f
C14702 DVSS.n6284 VSS 0.165082f
C14703 DVSS.n6285 VSS 0.165082f
C14704 DVSS.n6286 VSS 0.165082f
C14705 DVSS.n6287 VSS 0.165082f
C14706 DVSS.n6288 VSS 0.165082f
C14707 DVSS.n6289 VSS 0.165082f
C14708 DVSS.n6290 VSS 0.165082f
C14709 DVSS.n6291 VSS 0.165082f
C14710 DVSS.n6292 VSS 0.165082f
C14711 DVSS.n6293 VSS 0.165082f
C14712 DVSS.n6294 VSS 0.165082f
C14713 DVSS.n6295 VSS 0.165082f
C14714 DVSS.n6296 VSS 0.165082f
C14715 DVSS.n6297 VSS 0.165082f
C14716 DVSS.n6298 VSS 0.165082f
C14717 DVSS.n6299 VSS 0.165082f
C14718 DVSS.n6300 VSS 0.165082f
C14719 DVSS.n6301 VSS 0.165082f
C14720 DVSS.n6302 VSS 0.165082f
C14721 DVSS.n6303 VSS 0.165082f
C14722 DVSS.n6304 VSS 0.165082f
C14723 DVSS.n6305 VSS 0.165082f
C14724 DVSS.n6306 VSS 0.165082f
C14725 DVSS.n6307 VSS 0.165082f
C14726 DVSS.n6308 VSS 0.165082f
C14727 DVSS.n6309 VSS 0.165082f
C14728 DVSS.n6310 VSS 0.165082f
C14729 DVSS.n6311 VSS 0.165082f
C14730 DVSS.n6312 VSS 0.165082f
C14731 DVSS.n6313 VSS 0.165082f
C14732 DVSS.n6314 VSS 0.165082f
C14733 DVSS.n6315 VSS 0.165082f
C14734 DVSS.n6316 VSS 0.165082f
C14735 DVSS.n6317 VSS 0.165082f
C14736 DVSS.n6318 VSS 0.165082f
C14737 DVSS.n6319 VSS 0.165082f
C14738 DVSS.n6320 VSS 0.165082f
C14739 DVSS.n6321 VSS 0.165082f
C14740 DVSS.n6322 VSS 0.165082f
C14741 DVSS.n6323 VSS 0.165082f
C14742 DVSS.n6324 VSS 0.165082f
C14743 DVSS.n6325 VSS 0.165082f
C14744 DVSS.n6326 VSS 0.165082f
C14745 DVSS.n6327 VSS 0.165082f
C14746 DVSS.n6328 VSS 0.165082f
C14747 DVSS.n6329 VSS 0.165082f
C14748 DVSS.n6330 VSS 0.165082f
C14749 DVSS.n6331 VSS 0.165082f
C14750 DVSS.n6332 VSS 0.165082f
C14751 DVSS.n6333 VSS 0.165082f
C14752 DVSS.n6334 VSS 0.165082f
C14753 DVSS.n6335 VSS 0.165082f
C14754 DVSS.n6336 VSS 0.165082f
C14755 DVSS.n6337 VSS 0.165082f
C14756 DVSS.n6338 VSS 0.165082f
C14757 DVSS.n6339 VSS 0.165082f
C14758 DVSS.n6340 VSS 0.165082f
C14759 DVSS.n6341 VSS 0.165082f
C14760 DVSS.n6342 VSS 0.165082f
C14761 DVSS.n6343 VSS 0.072078f
C14762 DVSS.n6344 VSS 0.105183f
C14763 DVSS.n6345 VSS 1.26652f
C14764 DVSS.n6346 VSS 1.2663f
C14765 DVSS.n6347 VSS 0.105306f
C14766 DVSS.n6348 VSS 0.165082f
C14767 DVSS.n6349 VSS 0.165082f
C14768 DVSS.n6350 VSS 0.165082f
C14769 DVSS.n6351 VSS 0.165082f
C14770 DVSS.n6352 VSS 0.165082f
C14771 DVSS.n6353 VSS 0.165082f
C14772 DVSS.n6354 VSS 0.165082f
C14773 DVSS.n6355 VSS 0.165082f
C14774 DVSS.n6356 VSS 0.165082f
C14775 DVSS.n6357 VSS 0.165082f
C14776 DVSS.n6358 VSS 0.165082f
C14777 DVSS.n6359 VSS 0.165082f
C14778 DVSS.n6360 VSS 0.165082f
C14779 DVSS.n6361 VSS 0.165082f
C14780 DVSS.n6362 VSS 0.165082f
C14781 DVSS.n6363 VSS 0.165082f
C14782 DVSS.n6364 VSS 0.165082f
C14783 DVSS.n6365 VSS 0.165082f
C14784 DVSS.n6366 VSS 0.165082f
C14785 DVSS.n6367 VSS 0.165082f
C14786 DVSS.n6368 VSS 0.165082f
C14787 DVSS.n6369 VSS 0.165082f
C14788 DVSS.n6370 VSS 0.165082f
C14789 DVSS.n6371 VSS 0.165082f
C14790 DVSS.n6372 VSS 0.165082f
C14791 DVSS.n6373 VSS 0.165082f
C14792 DVSS.n6374 VSS 0.165082f
C14793 DVSS.n6375 VSS 0.165082f
C14794 DVSS.n6376 VSS 0.165082f
C14795 DVSS.n6377 VSS 0.165082f
C14796 DVSS.n6378 VSS 0.165082f
C14797 DVSS.n6379 VSS 0.165082f
C14798 DVSS.n6380 VSS 0.165082f
C14799 DVSS.n6381 VSS 0.165082f
C14800 DVSS.n6382 VSS 0.165082f
C14801 DVSS.n6383 VSS 0.165082f
C14802 DVSS.n6384 VSS 0.165082f
C14803 DVSS.n6385 VSS 0.165082f
C14804 DVSS.n6386 VSS 0.165082f
C14805 DVSS.n6387 VSS 0.165082f
C14806 DVSS.n6388 VSS 0.165082f
C14807 DVSS.n6389 VSS 0.165082f
C14808 DVSS.n6390 VSS 0.165082f
C14809 DVSS.n6391 VSS 0.165082f
C14810 DVSS.n6392 VSS 0.165082f
C14811 DVSS.n6393 VSS 0.165082f
C14812 DVSS.n6394 VSS 0.165082f
C14813 DVSS.n6395 VSS 0.165082f
C14814 DVSS.n6396 VSS 0.165082f
C14815 DVSS.n6397 VSS 0.165082f
C14816 DVSS.n6398 VSS 0.165082f
C14817 DVSS.n6399 VSS 0.165082f
C14818 DVSS.n6400 VSS 0.165082f
C14819 DVSS.n6401 VSS 0.165082f
C14820 DVSS.n6402 VSS 0.165082f
C14821 DVSS.n6403 VSS 0.165082f
C14822 DVSS.n6404 VSS 0.165082f
C14823 DVSS.n6405 VSS 0.165082f
C14824 DVSS.n6406 VSS 0.165082f
C14825 DVSS.n6407 VSS 0.165082f
C14826 DVSS.n6408 VSS 0.165082f
C14827 DVSS.n6409 VSS 0.165082f
C14828 DVSS.n6410 VSS 0.165082f
C14829 DVSS.n6411 VSS 0.165082f
C14830 DVSS.n6412 VSS 0.165082f
C14831 DVSS.n6413 VSS 0.165082f
C14832 DVSS.n6414 VSS 0.165082f
C14833 DVSS.n6415 VSS 0.165082f
C14834 DVSS.n6416 VSS 0.165082f
C14835 DVSS.n6417 VSS 0.165082f
C14836 DVSS.n6418 VSS 0.165082f
C14837 DVSS.n6419 VSS 0.165082f
C14838 DVSS.n6420 VSS 0.165082f
C14839 DVSS.n6421 VSS 0.165082f
C14840 DVSS.n6422 VSS 0.165082f
C14841 DVSS.n6423 VSS 0.165082f
C14842 DVSS.n6424 VSS 0.165082f
C14843 DVSS.n6425 VSS 0.165082f
C14844 DVSS.n6426 VSS 0.165082f
C14845 DVSS.n6427 VSS 0.165082f
C14846 DVSS.n6428 VSS 0.165082f
C14847 DVSS.n6429 VSS 0.165082f
C14848 DVSS.n6430 VSS 0.165082f
C14849 DVSS.n6431 VSS 0.165082f
C14850 DVSS.n6432 VSS 0.165082f
C14851 DVSS.n6433 VSS 0.165082f
C14852 DVSS.n6434 VSS 0.165082f
C14853 DVSS.n6435 VSS 0.162757f
C14854 DVSS.n6436 VSS 0.341473f
C14855 DVSS.n6437 VSS 0.315112f
C14856 DVSS.n6438 VSS 0.616179f
C14857 DVSS.n6439 VSS 0.165082f
C14858 DVSS.n6440 VSS 0.165082f
C14859 DVSS.n6441 VSS 0.165082f
C14860 DVSS.n6442 VSS 0.098817f
C14861 DVSS.n6443 VSS 0.098817f
C14862 DVSS.n6444 VSS 0.084866f
C14863 DVSS.n6445 VSS 0.165082f
C14864 DVSS.n6446 VSS 0.148806f
C14865 DVSS.n6447 VSS 0.148806f
C14866 DVSS.n6448 VSS 0.165082f
C14867 DVSS.n6449 VSS 0.165082f
C14868 DVSS.n6450 VSS 0.165082f
C14869 DVSS.n6451 VSS 0.165082f
C14870 DVSS.n6452 VSS 0.165082f
C14871 DVSS.n6453 VSS 0.165082f
C14872 DVSS.n6454 VSS 0.165082f
C14873 DVSS.n6455 VSS 0.165082f
C14874 DVSS.n6456 VSS 0.165082f
C14875 DVSS.n6457 VSS 0.165082f
C14876 DVSS.n6458 VSS 0.165082f
C14877 DVSS.n6459 VSS 0.165082f
C14878 DVSS.n6460 VSS 0.165082f
C14879 DVSS.n6461 VSS 0.165082f
C14880 DVSS.n6462 VSS 0.165082f
C14881 DVSS.n6463 VSS 0.165082f
C14882 DVSS.n6464 VSS 0.165082f
C14883 DVSS.n6465 VSS 0.165082f
C14884 DVSS.n6466 VSS 0.165082f
C14885 DVSS.n6467 VSS 0.165082f
C14886 DVSS.n6468 VSS 0.165082f
C14887 DVSS.n6469 VSS 0.165082f
C14888 DVSS.n6470 VSS 0.165082f
C14889 DVSS.n6471 VSS 0.165082f
C14890 DVSS.n6472 VSS 0.165082f
C14891 DVSS.n6473 VSS 0.165082f
C14892 DVSS.n6474 VSS 0.165082f
C14893 DVSS.n6475 VSS 0.165082f
C14894 DVSS.n6476 VSS 0.165082f
C14895 DVSS.n6477 VSS 0.165082f
C14896 DVSS.n6478 VSS 0.165082f
C14897 DVSS.n6479 VSS 0.165082f
C14898 DVSS.n6480 VSS 0.165082f
C14899 DVSS.n6481 VSS 0.165082f
C14900 DVSS.n6482 VSS 0.165082f
C14901 DVSS.n6483 VSS 0.165082f
C14902 DVSS.n6484 VSS 0.165082f
C14903 DVSS.n6485 VSS 0.165082f
C14904 DVSS.n6486 VSS 0.165082f
C14905 DVSS.n6487 VSS 0.165082f
C14906 DVSS.n6488 VSS 0.165082f
C14907 DVSS.n6489 VSS 0.165082f
C14908 DVSS.n6490 VSS 0.165082f
C14909 DVSS.n6491 VSS 0.165082f
C14910 DVSS.n6492 VSS 0.165082f
C14911 DVSS.n6493 VSS 0.165082f
C14912 DVSS.n6494 VSS 0.165082f
C14913 DVSS.n6495 VSS 0.165082f
C14914 DVSS.n6496 VSS 0.165082f
C14915 DVSS.n6497 VSS 0.165082f
C14916 DVSS.n6498 VSS 0.165082f
C14917 DVSS.n6499 VSS 0.165082f
C14918 DVSS.n6500 VSS 0.165082f
C14919 DVSS.n6501 VSS 0.165082f
C14920 DVSS.n6502 VSS 0.165082f
C14921 DVSS.n6503 VSS 0.165082f
C14922 DVSS.n6504 VSS 0.165082f
C14923 DVSS.n6505 VSS 0.165082f
C14924 DVSS.n6506 VSS 0.165082f
C14925 DVSS.n6507 VSS 0.165082f
C14926 DVSS.n6508 VSS 0.165082f
C14927 DVSS.n6509 VSS 0.165082f
C14928 DVSS.n6510 VSS 0.165082f
C14929 DVSS.n6511 VSS 0.165082f
C14930 DVSS.n6512 VSS 0.165082f
C14931 DVSS.n6513 VSS 0.165082f
C14932 DVSS.n6514 VSS 0.165082f
C14933 DVSS.n6515 VSS 0.165082f
C14934 DVSS.n6516 VSS 0.165082f
C14935 DVSS.n6517 VSS 0.165082f
C14936 DVSS.n6518 VSS 0.165082f
C14937 DVSS.n6519 VSS 0.165082f
C14938 DVSS.n6520 VSS 0.165082f
C14939 DVSS.n6521 VSS 0.165082f
C14940 DVSS.n6522 VSS 0.165082f
C14941 DVSS.n6523 VSS 0.165082f
C14942 DVSS.n6524 VSS 0.165082f
C14943 DVSS.n6525 VSS 0.165082f
C14944 DVSS.n6526 VSS 0.165082f
C14945 DVSS.n6527 VSS 0.165082f
C14946 DVSS.n6528 VSS 0.165082f
C14947 DVSS.n6529 VSS 0.165082f
C14948 DVSS.n6530 VSS 0.165082f
C14949 DVSS.n6531 VSS 0.165082f
C14950 DVSS.n6532 VSS 0.165082f
C14951 DVSS.n6533 VSS 0.165082f
C14952 DVSS.n6534 VSS 0.165082f
C14953 DVSS.n6535 VSS 0.165082f
C14954 DVSS.n6536 VSS 0.165082f
C14955 DVSS.n6537 VSS 0.165082f
C14956 DVSS.n6538 VSS 0.165082f
C14957 DVSS.n6539 VSS 0.165082f
C14958 DVSS.n6540 VSS 0.165082f
C14959 DVSS.n6541 VSS 0.165082f
C14960 DVSS.n6542 VSS 0.165082f
C14961 DVSS.n6543 VSS 0.165082f
C14962 DVSS.n6544 VSS 0.165082f
C14963 DVSS.n6545 VSS 0.165082f
C14964 DVSS.n6546 VSS 0.165082f
C14965 DVSS.n6547 VSS 0.165082f
C14966 DVSS.n6548 VSS 0.165082f
C14967 DVSS.n6549 VSS 0.165082f
C14968 DVSS.n6550 VSS 0.165082f
C14969 DVSS.n6551 VSS 0.165082f
C14970 DVSS.n6552 VSS 0.165082f
C14971 DVSS.n6553 VSS 0.165082f
C14972 DVSS.n6554 VSS 0.165082f
C14973 DVSS.n6555 VSS 0.165082f
C14974 DVSS.n6556 VSS 0.165082f
C14975 DVSS.n6557 VSS 0.165082f
C14976 DVSS.n6558 VSS 0.165082f
C14977 DVSS.n6559 VSS 0.165082f
C14978 DVSS.n6560 VSS 0.165082f
C14979 DVSS.n6561 VSS 0.165082f
C14980 DVSS.n6562 VSS 0.165082f
C14981 DVSS.n6563 VSS 0.165082f
C14982 DVSS.n6564 VSS 0.165082f
C14983 DVSS.n6565 VSS 0.165082f
C14984 DVSS.n6566 VSS 0.165082f
C14985 DVSS.n6567 VSS 0.165082f
C14986 DVSS.n6568 VSS 0.165082f
C14987 DVSS.n6569 VSS 0.165082f
C14988 DVSS.n6570 VSS 0.165082f
C14989 DVSS.n6571 VSS 0.165082f
C14990 DVSS.n6572 VSS 0.165082f
C14991 DVSS.n6573 VSS 0.165082f
C14992 DVSS.n6574 VSS 0.165082f
C14993 DVSS.n6575 VSS 0.165082f
C14994 DVSS.n6576 VSS 0.165082f
C14995 DVSS.n6577 VSS 0.165082f
C14996 DVSS.n6578 VSS 0.165082f
C14997 DVSS.n6579 VSS 0.165082f
C14998 DVSS.n6580 VSS 0.165082f
C14999 DVSS.n6581 VSS 0.165082f
C15000 DVSS.n6582 VSS 0.165082f
C15001 DVSS.n6583 VSS 0.165082f
C15002 DVSS.n6584 VSS 0.165082f
C15003 DVSS.n6585 VSS 0.165082f
C15004 DVSS.n6586 VSS 0.165082f
C15005 DVSS.n6587 VSS 0.165082f
C15006 DVSS.n6588 VSS 0.165082f
C15007 DVSS.n6589 VSS 0.165082f
C15008 DVSS.n6590 VSS 0.165082f
C15009 DVSS.n6591 VSS 0.165082f
C15010 DVSS.n6592 VSS 0.165082f
C15011 DVSS.n6593 VSS 0.165082f
C15012 DVSS.n6594 VSS 0.165082f
C15013 DVSS.n6595 VSS 0.165082f
C15014 DVSS.n6596 VSS 0.165082f
C15015 DVSS.n6597 VSS 0.165082f
C15016 DVSS.n6598 VSS 0.165082f
C15017 DVSS.n6599 VSS 0.165082f
C15018 DVSS.n6600 VSS 0.165082f
C15019 DVSS.n6601 VSS 0.165082f
C15020 DVSS.n6602 VSS 0.165082f
C15021 DVSS.n6603 VSS 0.165082f
C15022 DVSS.n6604 VSS 0.165082f
C15023 DVSS.n6605 VSS 0.165082f
C15024 DVSS.n6606 VSS 0.165082f
C15025 DVSS.n6607 VSS 0.165082f
C15026 DVSS.n6608 VSS 0.165082f
C15027 DVSS.n6609 VSS 0.165082f
C15028 DVSS.n6610 VSS 0.165082f
C15029 DVSS.n6611 VSS 0.165082f
C15030 DVSS.n6612 VSS 0.165082f
C15031 DVSS.n6613 VSS 0.165082f
C15032 DVSS.n6614 VSS 0.165082f
C15033 DVSS.n6615 VSS 0.165082f
C15034 DVSS.n6616 VSS 0.165082f
C15035 DVSS.n6617 VSS 0.114511f
C15036 DVSS.n6618 VSS 0.165082f
C15037 DVSS.n6619 VSS 0.165082f
C15038 DVSS.n6620 VSS 0.165082f
C15039 DVSS.n6621 VSS 0.165082f
C15040 DVSS.n6622 VSS 0.165082f
C15041 DVSS.n6623 VSS 0.143575f
C15042 DVSS.n6624 VSS 0.165082f
C15043 DVSS.n6625 VSS 0.165082f
C15044 DVSS.n6626 VSS 0.165082f
C15045 DVSS.n6627 VSS 0.165082f
C15046 DVSS.n6628 VSS 0.165082f
C15047 DVSS.n6629 VSS 0.165082f
C15048 DVSS.n6630 VSS 0.165082f
C15049 DVSS.n6631 VSS 0.165082f
C15050 DVSS.n6632 VSS 0.165082f
C15051 DVSS.n6633 VSS 0.165082f
C15052 DVSS.n6634 VSS 0.165082f
C15053 DVSS.n6635 VSS 0.165082f
C15054 DVSS.n6636 VSS 0.165082f
C15055 DVSS.n6637 VSS 0.611712f
C15056 DVSS.n6638 VSS 0.165082f
C15057 DVSS.n6639 VSS 0.165082f
C15058 DVSS.n6640 VSS 0.165082f
C15059 DVSS.n6641 VSS 0.336866f
C15060 DVSS.n6642 VSS 1.22581f
C15061 DVSS.n6643 VSS 1.40516f
C15062 DVSS.n6644 VSS 0.064709f
C15063 DVSS.n6645 VSS 0.249392f
C15064 DVSS.n6646 VSS 0.038205f
C15065 DVSS.n6648 VSS 0.030471f
C15066 DVSS.n6650 VSS 0.74982f
C15067 DVSS.t25 VSS 0.330478f
C15068 DVSS.n6653 VSS 0.635269f
C15069 DVSS.n6655 VSS 0.74982f
C15070 DVSS.n6659 VSS 0.74982f
C15071 DVSS.n6662 VSS 0.116237f
C15072 DVSS.n6664 VSS 0.032106f
C15073 DVSS.n6665 VSS 0.032106f
C15074 DVSS.n6667 VSS 0.082541f
C15075 DVSS.n6668 VSS 0.082541f
C15076 DVSS.n6669 VSS 0.147063f
C15077 DVSS.n6670 VSS 0.052308f
C15078 DVSS.n6671 VSS 0.052308f
C15079 DVSS.n6672 VSS 0.052308f
C15080 DVSS.n6673 VSS 0.052308f
C15081 DVSS.n6674 VSS 0.052308f
C15082 DVSS.n6675 VSS 0.072078f
C15083 DVSS.n6677 VSS 0.052308f
C15084 DVSS.n6679 VSS 0.052308f
C15085 DVSS.n6681 VSS 0.052308f
C15086 DVSS.n6683 VSS 0.052308f
C15087 DVSS.n6689 VSS 0.082541f
C15088 DVSS.n6691 VSS 0.176874f
C15089 DVSS.n6692 VSS 0.176874f
C15090 DVSS.n6693 VSS 0.315134f
C15091 DVSS.n6694 VSS 0.052308f
C15092 DVSS.n6695 VSS 0.052308f
C15093 DVSS.n6696 VSS 0.052308f
C15094 DVSS.n6697 VSS 0.052308f
C15095 DVSS.n6698 VSS 0.052308f
C15096 DVSS.n6699 VSS 0.052308f
C15097 DVSS.n6700 VSS 0.052308f
C15098 DVSS.n6701 VSS 0.052308f
C15099 DVSS.n6702 VSS 0.052308f
C15100 DVSS.n6703 VSS 0.052308f
C15101 DVSS.n6704 VSS 0.154453f
C15102 DVSS.n6706 VSS 0.052308f
C15103 DVSS.n6708 VSS 0.052308f
C15104 DVSS.n6710 VSS 0.052308f
C15105 DVSS.n6712 VSS 0.052308f
C15106 DVSS.n6714 VSS 0.052308f
C15107 DVSS.n6716 VSS 0.052308f
C15108 DVSS.n6718 VSS 0.052308f
C15109 DVSS.n6720 VSS 0.052308f
C15110 DVSS.n6722 VSS 0.052308f
C15111 DVSS.n6724 VSS 0.052308f
C15112 DVSS.n6725 VSS 0.353747f
C15113 DVSS.n6726 VSS 0.154453f
C15114 DVSS.n6727 VSS 0.353747f
C15115 DVSS.n6728 VSS 0.353747f
C15116 DVSS.n6729 VSS 0.353747f
C15117 DVSS.n6730 VSS 0.282749f
C15118 DVSS.n6731 VSS 0.353747f
C15119 DVSS.n6732 VSS 1.31154f
C15120 DVSS.n6733 VSS 0.353747f
C15121 DVSS.n6734 VSS 0.176874f
C15122 DVSS.n6736 VSS 0.082541f
C15123 DVSS.n6737 VSS 0.082541f
C15124 DVSS.n6738 VSS 0.3147f
C15125 DVSS.n6739 VSS 0.052308f
C15126 DVSS.n6740 VSS 0.052308f
C15127 DVSS.n6741 VSS 0.052308f
C15128 DVSS.n6742 VSS 0.052308f
C15129 DVSS.n6743 VSS 0.052308f
C15130 DVSS.n6744 VSS 0.072078f
C15131 DVSS.n6745 VSS 0.045559f
C15132 DVSS.n6747 VSS 0.133296f
C15133 DVSS.t32 VSS 0.394423f
C15134 DVSS.n6749 VSS 0.233666f
C15135 DVSS.n6750 VSS 0.032106f
C15136 DVSS.n6752 VSS 0.027052f
C15137 DVSS.n6753 VSS 1.58569f
C15138 DVSS.n6755 VSS 1.58907f
C15139 DVSS.n6757 VSS 0.052308f
C15140 DVSS.n6759 VSS 0.052308f
C15141 DVSS.n6761 VSS 0.052308f
C15142 DVSS.n6762 VSS 0.072078f
C15143 DVSS.n6763 VSS 0.165082f
C15144 DVSS.n6764 VSS 0.165082f
C15145 DVSS.n6765 VSS 0.165082f
C15146 DVSS.n6766 VSS 0.165082f
C15147 DVSS.n6767 VSS 0.072078f
C15148 DVSS.n6768 VSS 0.165082f
C15149 DVSS.n6769 VSS 0.611712f
C15150 DVSS.n6770 VSS 0.165082f
C15151 DVSS.n6771 VSS 0.165082f
C15152 DVSS.n6772 VSS 0.165082f
C15153 DVSS.n6773 VSS 0.165082f
C15154 DVSS.n6774 VSS 0.165082f
C15155 DVSS.n6775 VSS 0.165082f
C15156 DVSS.n6776 VSS 0.165082f
C15157 DVSS.n6777 VSS 0.165082f
C15158 DVSS.n6778 VSS 0.165082f
C15159 DVSS.n6779 VSS 0.165082f
C15160 DVSS.n6780 VSS 0.072078f
C15161 DVSS.n6781 VSS 0.165082f
C15162 DVSS.n6782 VSS 0.165082f
C15163 DVSS.n6783 VSS 0.165082f
C15164 DVSS.n6784 VSS 0.165082f
C15165 DVSS.n6785 VSS 0.165082f
C15166 DVSS.n6786 VSS 0.165082f
C15167 DVSS.n6787 VSS 0.165082f
C15168 DVSS.n6788 VSS 0.165082f
C15169 DVSS.n6789 VSS 0.165082f
C15170 DVSS.n6790 VSS 0.165082f
C15171 DVSS.n6791 VSS 0.165082f
C15172 DVSS.n6792 VSS 0.165082f
C15173 DVSS.n6793 VSS 0.165082f
C15174 DVSS.n6794 VSS 0.165082f
C15175 DVSS.n6795 VSS 0.165082f
C15176 DVSS.n6796 VSS 0.165082f
C15177 DVSS.n6797 VSS 0.165082f
C15178 DVSS.n6798 VSS 0.165082f
C15179 DVSS.n6799 VSS 0.165082f
C15180 DVSS.n6800 VSS 0.165082f
C15181 DVSS.n6801 VSS 0.165082f
C15182 DVSS.n6802 VSS 0.165082f
C15183 DVSS.n6803 VSS 0.165082f
C15184 DVSS.n6804 VSS 0.165082f
C15185 DVSS.n6805 VSS 0.165082f
C15186 DVSS.n6806 VSS 0.165082f
C15187 DVSS.n6807 VSS 0.165082f
C15188 DVSS.n6808 VSS 0.165082f
C15189 DVSS.n6809 VSS 0.165082f
C15190 DVSS.n6810 VSS 0.165082f
C15191 DVSS.n6811 VSS 0.165082f
C15192 DVSS.n6812 VSS 0.165082f
C15193 DVSS.n6813 VSS 0.165082f
C15194 DVSS.n6814 VSS 0.165082f
C15195 DVSS.n6815 VSS 0.165082f
C15196 DVSS.n6816 VSS 0.165082f
C15197 DVSS.n6817 VSS 0.131949f
C15198 DVSS.n6818 VSS 0.165082f
C15199 DVSS.n6819 VSS 0.165082f
C15200 DVSS.n6820 VSS 0.165082f
C15201 DVSS.n6821 VSS 0.165082f
C15202 DVSS.n6822 VSS 0.072078f
C15203 DVSS.n6823 VSS 0.165082f
C15204 DVSS.n6824 VSS 0.165082f
C15205 DVSS.n6825 VSS 0.165082f
C15206 DVSS.n6826 VSS 0.165082f
C15207 DVSS.n6827 VSS 0.165082f
C15208 DVSS.n6828 VSS 0.165082f
C15209 DVSS.n6829 VSS 0.165082f
C15210 DVSS.n6830 VSS 0.165082f
C15211 DVSS.n6831 VSS 0.165082f
C15212 DVSS.n6832 VSS 0.131949f
C15213 DVSS.n6833 VSS 0.165082f
C15214 DVSS.n6834 VSS 0.072078f
C15215 DVSS.n6835 VSS 0.165082f
C15216 DVSS.n6836 VSS 0.072078f
C15217 DVSS.n6837 VSS 0.165082f
C15218 DVSS.n6838 VSS 0.165082f
C15219 DVSS.n6839 VSS 0.165082f
C15220 DVSS.n6840 VSS 0.165082f
C15221 DVSS.n6841 VSS 0.165082f
C15222 DVSS.n6842 VSS 0.165082f
C15223 DVSS.n6843 VSS 0.165082f
C15224 DVSS.n6844 VSS 0.165082f
C15225 DVSS.n6845 VSS 0.165082f
C15226 DVSS.n6846 VSS 0.165082f
C15227 DVSS.n6847 VSS 0.165082f
C15228 DVSS.n6848 VSS 0.165082f
C15229 DVSS.n6849 VSS 0.165082f
C15230 DVSS.n6850 VSS 0.131949f
C15231 DVSS.n6854 VSS 0.082541f
C15232 DVSS.n6857 VSS 0.052308f
C15233 DVSS.n6858 VSS 0.361112f
C15234 DVSS.n6859 VSS 0.438291f
C15235 DVSS.n6860 VSS 0.438291f
C15236 DVSS.n6861 VSS 0.052308f
C15237 DVSS.n6872 VSS 0.099554f
C15238 DVSS.n6874 VSS 0.672799f
C15239 DVSS.n6875 VSS 0.052308f
C15240 DVSS.n6876 VSS 0.052308f
C15241 DVSS.n6877 VSS 0.052308f
C15242 DVSS.n6878 VSS 0.052308f
C15243 DVSS.n6879 VSS 0.052308f
C15244 DVSS.n6880 VSS 0.052308f
C15245 DVSS.n6881 VSS 0.052308f
C15246 DVSS.n6882 VSS 0.052308f
C15247 DVSS.n6883 VSS 0.052308f
C15248 DVSS.n6884 VSS 0.052308f
C15249 DVSS.n6885 VSS 0.353747f
C15250 DVSS.n6886 VSS 0.154453f
C15251 DVSS.n6888 VSS 0.052308f
C15252 DVSS.n6889 VSS 0.052308f
C15253 DVSS.n6890 VSS 0.052308f
C15254 DVSS.n6891 VSS 0.052308f
C15255 DVSS.n6892 VSS 0.052308f
C15256 DVSS.n6893 VSS 0.052308f
C15257 DVSS.n6894 VSS 0.052308f
C15258 DVSS.n6895 VSS 0.052308f
C15259 DVSS.n6905 VSS 0.154453f
C15260 DVSS.n6906 VSS 0.176874f
C15261 DVSS.n6908 VSS 0.052308f
C15262 DVSS.n6909 VSS 0.052308f
C15263 DVSS.n6910 VSS 0.774638f
C15264 DVSS.n6911 VSS 0.052308f
C15265 DVSS.n6913 VSS 0.176874f
C15266 DVSS.n6914 VSS 0.154453f
C15267 DVSS.n6915 VSS 0.353747f
C15268 DVSS.n6916 VSS 0.353747f
C15269 DVSS.n6917 VSS 0.353747f
C15270 DVSS.n6918 VSS 0.353747f
C15271 DVSS.n6919 VSS 0.353747f
C15272 DVSS.n6920 VSS 0.353747f
C15273 DVSS.n6921 VSS 0.353747f
C15274 DVSS.n6922 VSS 0.353747f
C15275 DVSS.n6923 VSS 0.353747f
C15276 DVSS.n6924 VSS 0.353747f
C15277 DVSS.n6925 VSS 0.353747f
C15278 DVSS.n6926 VSS 0.353747f
C15279 DVSS.n6927 VSS 0.353747f
C15280 DVSS.n6928 VSS 0.353747f
C15281 DVSS.n6929 VSS 0.282749f
C15282 DVSS.n6930 VSS 0.353747f
C15283 DVSS.n6931 VSS 0.052308f
C15284 DVSS.n6932 VSS 0.052308f
C15285 DVSS.n6933 VSS 0.052308f
C15286 DVSS.n6934 VSS 0.052308f
C15287 DVSS.n6935 VSS 0.052308f
C15288 DVSS.n6936 VSS 0.052308f
C15289 DVSS.n6937 VSS 0.052308f
C15290 DVSS.n6938 VSS 0.052308f
C15291 DVSS.n6939 VSS 0.052308f
C15292 DVSS.n6940 VSS 0.052308f
C15293 DVSS.n6941 VSS 0.052308f
C15294 DVSS.n6942 VSS 0.031427f
C15295 DVSS.n6943 VSS 0.154453f
C15296 DVSS.n6944 VSS 0.052308f
C15297 DVSS.n6945 VSS 0.052308f
C15298 DVSS.n6946 VSS 0.052308f
C15299 DVSS.n6947 VSS 0.052308f
C15300 DVSS.n6948 VSS 0.052308f
C15301 DVSS.n6949 VSS 0.052308f
C15302 DVSS.n6950 VSS 0.052308f
C15303 DVSS.n6951 VSS 0.052308f
C15304 DVSS.n6952 VSS 0.052308f
C15305 DVSS.n6953 VSS 0.052308f
C15306 DVSS.n6954 VSS 0.052308f
C15307 DVSS.n6967 VSS 0.176874f
C15308 DVSS.n6968 VSS 0.154453f
C15309 DVSS.n6979 VSS 0.176874f
C15310 DVSS.n6980 VSS 0.353747f
C15311 DVSS.n6981 VSS 0.353747f
C15312 DVSS.n6982 VSS 0.293959f
C15313 DVSS.n6983 VSS 0.353747f
C15314 DVSS.n6984 VSS 0.353747f
C15315 DVSS.n6985 VSS 0.353747f
C15316 DVSS.n6986 VSS 0.353747f
C15317 DVSS.n6987 VSS 0.282749f
C15318 DVSS.n6988 VSS 0.353747f
C15319 DVSS.n6989 VSS 0.353747f
C15320 DVSS.n6990 VSS 0.353747f
C15321 DVSS.n6991 VSS 0.353747f
C15322 DVSS.n6992 VSS 0.353747f
C15323 DVSS.n6993 VSS 0.353747f
C15324 DVSS.n6994 VSS 0.353747f
C15325 DVSS.n6995 VSS 0.353747f
C15326 DVSS.n6996 VSS 0.353747f
C15327 DVSS.n6997 VSS 0.353747f
C15328 DVSS.n6998 VSS 0.353747f
C15329 DVSS.n6999 VSS 0.353747f
C15330 DVSS.n7000 VSS 0.353747f
C15331 DVSS.n7001 VSS 0.353747f
C15332 DVSS.n7002 VSS 0.353747f
C15333 DVSS.n7003 VSS 0.315134f
C15334 DVSS.n7004 VSS 0.353747f
C15335 DVSS.n7005 VSS 0.353747f
C15336 DVSS.n7006 VSS 0.353747f
C15337 DVSS.n7007 VSS 0.353747f
C15338 DVSS.n7008 VSS 0.353747f
C15339 DVSS.n7009 VSS 0.353747f
C15340 DVSS.n7010 VSS 0.353747f
C15341 DVSS.n7011 VSS 0.353747f
C15342 DVSS.n7012 VSS 0.353747f
C15343 DVSS.n7013 VSS 0.353747f
C15344 DVSS.n7014 VSS 0.353747f
C15345 DVSS.n7015 VSS 0.353747f
C15346 DVSS.n7016 VSS 0.353747f
C15347 DVSS.n7017 VSS 0.353747f
C15348 DVSS.n7018 VSS 0.353747f
C15349 DVSS.n7019 VSS 0.353747f
C15350 DVSS.n7020 VSS 0.353747f
C15351 DVSS.n7021 VSS 0.353747f
C15352 DVSS.n7022 VSS 0.353747f
C15353 DVSS.n7023 VSS 0.353747f
C15354 DVSS.n7024 VSS 0.353747f
C15355 DVSS.n7025 VSS 0.353747f
C15356 DVSS.n7026 VSS 0.154453f
C15357 DVSS.n7028 VSS 0.176874f
C15358 DVSS.n7029 VSS 0.099554f
C15359 DVSS.n7030 VSS 0.176874f
C15360 DVSS.n7031 VSS 0.255346f
C15361 DVSS.n7032 VSS 0.675109f
C15362 DVSS.n7033 VSS 0.425991f
C15363 DVSS.n7034 VSS 0.236662f
C15364 DVSS.n7035 VSS 0.353747f
C15365 DVSS.n7036 VSS 0.236662f
C15366 DVSS.n7037 VSS 0.353747f
C15367 DVSS.n7038 VSS 0.353747f
C15368 DVSS.n7039 VSS 0.353747f
C15369 DVSS.n7040 VSS 0.353747f
C15370 DVSS.n7041 VSS 0.353747f
C15371 DVSS.n7042 VSS 0.353747f
C15372 DVSS.n7043 VSS 0.353747f
C15373 DVSS.n7044 VSS 0.353747f
C15374 DVSS.n7045 VSS 0.154453f
C15375 DVSS.n7055 VSS 0.176874f
C15376 DVSS.n7058 VSS 0.052308f
C15377 DVSS.n7059 VSS 0.176874f
C15378 DVSS.n7060 VSS 0.438291f
C15379 DVSS.n7061 VSS 0.438291f
C15380 DVSS.n7062 VSS 0.082541f
C15381 DVSS.n7063 VSS 1.58907f
C15382 DVSS.n7064 VSS 1.58569f
C15383 DVSS.n7065 VSS 0.032106f
C15384 DVSS.n7066 VSS 0.045559f
C15385 DVSS.n7067 VSS 0.092157f
C15386 DVSS.n7068 VSS 0.044592f
C15387 DVSS.n7070 VSS 0.032106f
C15388 DVSS.n7071 VSS 0.032106f
C15389 DVSS.n7073 VSS 0.009955f
C15390 DVSS.n7074 VSS 0.019909f
C15391 DVSS.n7075 VSS 0.009955f
C15392 DVSS.n7077 VSS 0.180752f
C15393 DVSS.n7081 VSS 0.019909f
C15394 DVSS.n7082 VSS 0.019909f
C15395 DVSS.n7083 VSS 0.132478f
C15396 DVSS.n7084 VSS 0.017421f
C15397 DVSS.n7087 VSS 0.019909f
C15398 DVSS.n7091 VSS 0.019909f
C15399 DVSS.n7092 VSS 0.014932f
C15400 DVSS.n7093 VSS 0.017421f
C15401 DVSS.n7094 VSS 0.019909f
C15402 DVSS.n7095 VSS 0.132478f
C15403 DVSS.n7096 VSS 0.180752f
C15404 DVSS.n7097 VSS 0.35357f
C15405 DVSS.n7098 VSS 0.35357f
C15406 DVSS.n7100 VSS 0.019909f
C15407 DVSS.n7101 VSS 0.019909f
C15408 DVSS.n7102 VSS 0.134247f
C15409 DVSS.n7103 VSS 0.017421f
C15410 DVSS.n7104 VSS 0.014932f
C15411 DVSS.n7105 VSS 0.019909f
C15412 DVSS.n7106 VSS 0.180752f
C15413 DVSS.n7107 VSS 0.134247f
C15414 DVSS.n7108 VSS 0.017421f
C15415 DVSS.n7109 VSS 0.35357f
C15416 DVSS.n7110 VSS 0.35357f
C15417 DVSS.n7111 VSS 0.180752f
C15418 DVSS.n7112 VSS 0.180752f
C15419 DVSS.n7113 VSS 0.019909f
C15420 DVSS.n7114 VSS 0.019909f
C15421 DVSS.n7115 VSS 0.009955f
C15422 DVSS.n7116 VSS 0.009955f
C15423 DVSS.n7117 VSS 0.184214f
C15424 DVSS.n7118 VSS 0.421629f
C15425 DVSS.n7119 VSS 0.421629f
C15426 DVSS.n7120 VSS 0.019909f
C15427 DVSS.n7121 VSS 0.019909f
C15428 DVSS.n7122 VSS 0.009955f
C15429 DVSS.n7123 VSS 0.160088f
C15430 DVSS.n7124 VSS 0.179554f
C15431 DVSS.n7125 VSS 0.009955f
C15432 DVSS.n7126 VSS 0.019909f
C15433 DVSS.n7127 VSS 0.160088f
C15434 DVSS.n7128 VSS 0.179554f
C15435 DVSS.n7129 VSS 1.42561f
C15436 DVSS.n7130 VSS 1.42561f
C15437 DVSS.n7131 VSS 0.032106f
C15438 DVSS.n7132 VSS 0.045559f
C15439 DVSS.n7133 VSS 0.148938f
C15440 DVSS.n7134 VSS 0.548192f
C15441 DVSS.n7135 VSS 0.097211f
C15442 DVSS.n7137 VSS 0.032106f
C15443 DVSS.n7138 VSS 0.032106f
C15444 DVSS.n7140 VSS 0.009955f
C15445 DVSS.n7141 VSS 0.019909f
C15446 DVSS.n7142 VSS 0.019909f
C15447 DVSS.n7143 VSS 0.180752f
C15448 DVSS.n7144 VSS 0.009955f
C15449 DVSS.n7145 VSS 0.330782f
C15450 DVSS.n7146 VSS 0.211948f
C15451 DVSS.n7147 VSS 0.184214f
C15452 DVSS.n7148 VSS 0.157979f
C15453 DVSS.n7149 VSS 0.180752f
C15454 DVSS.n7150 VSS 0.297397f
C15455 DVSS.n7151 VSS 0.297397f
C15456 DVSS.n7152 VSS 0.032106f
C15457 DVSS.n7153 VSS 0.045559f
C15458 DVSS.n7154 VSS 0.096319f
C15459 DVSS.n7155 VSS 0.06562f
C15460 DVSS.n7156 VSS 0.061615f
C15461 DVSS.n7157 VSS 0.038205f
C15462 DVSS.n7158 VSS 0.035873f
C15463 DVSS.n7159 VSS 0.038205f
C15464 DVSS.n7160 VSS 0.035873f
C15465 DVSS.n7161 VSS 0.038205f
C15466 DVSS.n7162 VSS 0.035873f
C15467 DVSS.n7163 VSS 0.038205f
C15468 DVSS.n7164 VSS 0.035873f
C15469 DVSS.n7165 VSS 0.038205f
C15470 DVSS.n7166 VSS 0.035873f
C15471 DVSS.n7167 VSS 0.038205f
C15472 DVSS.n7168 VSS 0.038205f
C15473 DVSS.t9 VSS 0.330478f
C15474 DVSS.n7169 VSS 0.125906f
C15475 DVSS.n7170 VSS 0.038205f
C15476 DVSS.n7171 VSS 0.035873f
C15477 DVSS.n7172 VSS 0.038205f
C15478 DVSS.n7173 VSS 0.035873f
C15479 DVSS.n7174 VSS 0.038205f
C15480 DVSS.n7175 VSS 0.035873f
C15481 DVSS.n7176 VSS 0.038205f
C15482 DVSS.n7177 VSS 0.035873f
C15483 DVSS.n7178 VSS 0.038205f
C15484 DVSS.n7179 VSS 0.035873f
C15485 DVSS.n7180 VSS 0.038205f
C15486 DVSS.n7181 VSS 0.035873f
C15487 DVSS.n7182 VSS 0.066505f
C15488 DVSS.n7183 VSS 0.031887f
C15489 DVSS.n7184 VSS 0.066505f
C15490 DVSS.n7185 VSS 0.038205f
C15491 DVSS.n7186 VSS 0.035873f
C15492 DVSS.n7187 VSS 0.038205f
C15493 DVSS.n7188 VSS 0.038205f
C15494 DVSS.n7189 VSS 0.038205f
C15495 DVSS.n7190 VSS 0.035873f
C15496 DVSS.n7191 VSS 0.038205f
C15497 DVSS.n7192 VSS 0.038205f
C15498 DVSS.n7193 VSS 0.038205f
C15499 DVSS.n7194 VSS 0.035873f
C15500 DVSS.n7195 VSS 0.038205f
C15501 DVSS.n7196 VSS 0.038205f
C15502 DVSS.n7197 VSS 0.038205f
C15503 DVSS.n7198 VSS 0.035873f
C15504 DVSS.n7199 VSS 0.038205f
C15505 DVSS.n7200 VSS 0.038205f
C15506 DVSS.n7201 VSS 0.038205f
C15507 DVSS.n7202 VSS 0.035873f
C15508 DVSS.n7203 VSS 0.038205f
C15509 DVSS.n7204 VSS 0.038205f
C15510 DVSS.n7205 VSS 0.038205f
C15511 DVSS.n7206 VSS 0.035873f
C15512 DVSS.n7207 VSS 0.038205f
C15513 DVSS.n7208 VSS 0.038205f
C15514 DVSS.n7209 VSS 0.038205f
C15515 DVSS.n7210 VSS 0.026905f
C15516 DVSS.n7211 VSS 0.038205f
C15517 DVSS.n7212 VSS 0.038205f
C15518 DVSS.n7213 VSS 0.026905f
C15519 DVSS.n7214 VSS 0.020096f
C15520 DVSS.n7215 VSS 0.038205f
C15521 DVSS.n7216 VSS 0.038205f
C15522 DVSS.n7217 VSS 0.033714f
C15523 DVSS.n7218 VSS 0.038205f
C15524 DVSS.n7219 VSS 0.038205f
C15525 DVSS.n7220 VSS 0.038205f
C15526 DVSS.n7221 VSS 0.035873f
C15527 DVSS.n7222 VSS 0.038205f
C15528 DVSS.n7223 VSS 0.038205f
C15529 DVSS.n7224 VSS 0.038205f
C15530 DVSS.n7225 VSS 0.035873f
C15531 DVSS.n7226 VSS 0.038205f
C15532 DVSS.n7227 VSS 0.038205f
C15533 DVSS.n7228 VSS 0.038205f
C15534 DVSS.n7229 VSS 0.035873f
C15535 DVSS.n7230 VSS 0.038205f
C15536 DVSS.n7231 VSS 0.038205f
C15537 DVSS.n7232 VSS 0.038205f
C15538 DVSS.n7233 VSS 0.035873f
C15539 DVSS.n7234 VSS 0.038205f
C15540 DVSS.n7235 VSS 0.038205f
C15541 DVSS.n7236 VSS 0.038205f
C15542 DVSS.n7237 VSS 0.035873f
C15543 DVSS.n7238 VSS 0.038205f
C15544 DVSS.n7239 VSS 0.06562f
C15545 DVSS.n7240 VSS 0.030471f
C15546 DVSS.n7242 VSS 0.211218f
C15547 DVSS.n7244 VSS 0.038205f
C15548 DVSS.n7246 VSS 0.06562f
C15549 DVSS.n7247 VSS 0.061615f
C15550 DVSS.n7248 VSS 0.06562f
C15551 DVSS.n7250 VSS 0.211218f
C15552 DVSS.n7252 VSS 0.249392f
C15553 DVSS.n7253 VSS -0.427805f
C15554 DVSS.n7254 VSS 37.626503f
C15555 DVSS.n7255 VSS 14.8586f
C15556 DVSS.n7256 VSS 1.13994f
C15557 DVSS.n7257 VSS 9.96353f
C15558 DVSS.n7258 VSS 2.69552f
C15559 DVSS.n7259 VSS 9.972879f
C15560 DVSS.n7260 VSS 1.40512f
C15561 DVSS.n7261 VSS 2.56914f
C15562 DVSS.n7262 VSS 24.6928f
C15563 DVSS.n7263 VSS 25.8271f
C15564 DVSS.n7264 VSS 48.8624f
C15565 DVSS.n7265 VSS -0.427302f
C15566 DVSS.n7266 VSS 0.043865f
C15567 DVSS.n7269 VSS 0.043865f
C15568 DVSS.n7270 VSS 0.065379f
C15569 DVSS.n7271 VSS 0.069335f
C15570 DVSS.n7272 VSS 0.066505f
C15571 DVSS.n7273 VSS 0.038205f
C15572 DVSS.n7274 VSS 0.035873f
C15573 DVSS.n7275 VSS 0.038205f
C15574 DVSS.n7276 VSS 0.038205f
C15575 DVSS.n7277 VSS 0.038205f
C15576 DVSS.n7278 VSS 0.035873f
C15577 DVSS.n7279 VSS 0.038205f
C15578 DVSS.n7280 VSS 0.038205f
C15579 DVSS.n7281 VSS 0.038205f
C15580 DVSS.n7282 VSS 0.035873f
C15581 DVSS.n7283 VSS 0.038205f
C15582 DVSS.n7284 VSS 0.038205f
C15583 DVSS.n7285 VSS 0.038205f
C15584 DVSS.n7286 VSS 0.035873f
C15585 DVSS.n7287 VSS 0.038205f
C15586 DVSS.n7288 VSS 0.038205f
C15587 DVSS.n7289 VSS 0.038205f
C15588 DVSS.n7290 VSS 0.035873f
C15589 DVSS.n7291 VSS 0.038205f
C15590 DVSS.n7292 VSS 0.038205f
C15591 DVSS.n7293 VSS 0.038205f
C15592 DVSS.n7294 VSS 0.035873f
C15593 DVSS.n7295 VSS 0.038205f
C15594 DVSS.n7296 VSS 0.038205f
C15595 DVSS.n7297 VSS 0.038205f
C15596 DVSS.n7298 VSS 0.026905f
C15597 DVSS.n7299 VSS 0.038205f
C15598 DVSS.n7300 VSS 0.038205f
C15599 DVSS.n7301 VSS 0.038205f
C15600 DVSS.n7302 VSS 0.020096f
C15601 DVSS.n7303 VSS 0.038205f
C15602 DVSS.n7304 VSS 0.038205f
C15603 DVSS.n7305 VSS 0.038205f
C15604 DVSS.n7306 VSS 0.035873f
C15605 DVSS.n7307 VSS 0.038205f
C15606 DVSS.n7308 VSS 0.038205f
C15607 DVSS.n7309 VSS 0.038205f
C15608 DVSS.n7310 VSS 0.035873f
C15609 DVSS.n7311 VSS 0.038205f
C15610 DVSS.n7312 VSS 0.038205f
C15611 DVSS.n7313 VSS 0.038205f
C15612 DVSS.n7314 VSS 0.035873f
C15613 DVSS.n7315 VSS 0.038205f
C15614 DVSS.n7316 VSS 0.038205f
C15615 DVSS.n7317 VSS 0.038205f
C15616 DVSS.n7318 VSS 0.035873f
C15617 DVSS.n7319 VSS 0.038205f
C15618 DVSS.n7320 VSS 0.038205f
C15619 DVSS.n7321 VSS 0.038205f
C15620 DVSS.n7322 VSS 0.035873f
C15621 DVSS.n7323 VSS 0.038205f
C15622 DVSS.n7324 VSS 0.038205f
C15623 DVSS.n7326 VSS 0.069335f
C15624 DVSS.n7327 VSS 0.066505f
C15625 DVSS.n7328 VSS 0.049824f
C15626 DVSS.n7329 VSS 0.066505f
C15627 DVSS.n7330 VSS 0.069335f
C15628 DVSS.n7332 VSS 0.043865f
C15629 DVSS.n7333 VSS 0.396845f
C15630 DVSS.n7335 VSS 0.157135f
C15631 DVSS.n7337 VSS 0.066724f
C15632 DVSS.n7338 VSS 0.052308f
C15633 DVSS.n7339 VSS 0.186719f
C15634 DVSS.n7340 VSS 0.754249f
C15635 DVSS.n7342 VSS 0.242143f
C15636 DVSS.n7343 VSS 0.756156f
C15637 DVSS.n7345 VSS 0.157135f
C15638 DVSS.n7347 VSS 0.066724f
C15639 DVSS.n7348 VSS 0.052308f
C15640 DVSS.n7349 VSS 0.335771f
C15641 DVSS.n7350 VSS 0.754249f
C15642 DVSS.n7352 VSS 0.09309f
C15643 DVSS.n7354 VSS 0.157135f
C15644 DVSS.n7356 VSS 0.066724f
C15645 DVSS.n7357 VSS 0.052308f
C15646 DVSS.n7358 VSS 0.179185f
C15647 DVSS.n7359 VSS 0.754249f
C15648 DVSS.n7361 VSS 0.222771f
C15649 DVSS.n7362 VSS 0.331802f
C15650 DVSS.n7364 VSS 0.045559f
C15651 DVSS.n7365 VSS 0.058114f
C15652 DVSS.n7367 VSS 0.16051f
C15653 DVSS.n7368 VSS 0.048967f
C15654 DVSS.n7369 VSS 0.045559f
C15655 DVSS.n7371 VSS 0.764373f
C15656 DVSS.n7372 VSS 0.764373f
C15657 DVSS.n7373 VSS 0.048967f
C15658 DVSS.n7374 VSS 0.045559f
C15659 DVSS.n7376 VSS 0.048301f
C15660 DVSS.n7377 VSS 0.154453f
C15661 DVSS.n7378 VSS 0.774638f
C15662 DVSS.n7379 VSS 0.051675f
C15663 DVSS.n7380 VSS 0.176874f
C15664 DVSS.n7381 VSS 0.154453f
C15665 DVSS.n7382 VSS 0.353747f
C15666 DVSS.n7383 VSS 1.31154f
C15667 DVSS.n7384 VSS 0.353747f
C15668 DVSS.n7385 VSS 0.353747f
C15669 DVSS.n7386 VSS 0.353747f
C15670 DVSS.n7387 VSS 0.282749f
C15671 DVSS.n7388 VSS 0.353747f
C15672 DVSS.n7389 VSS 0.353747f
C15673 DVSS.n7390 VSS 0.353747f
C15674 DVSS.n7391 VSS 0.353747f
C15675 DVSS.n7392 VSS 0.353747f
C15676 DVSS.n7393 VSS 0.353747f
C15677 DVSS.n7394 VSS 0.353747f
C15678 DVSS.n7395 VSS 0.315134f
C15679 DVSS.n7396 VSS 0.154453f
C15680 DVSS.n7397 VSS 0.176874f
C15681 DVSS.n7398 VSS 0.044926f
C15682 DVSS.n7399 VSS 0.176874f
C15683 DVSS.n7400 VSS 0.154453f
C15684 DVSS.n7401 VSS 0.353747f
C15685 DVSS.n7402 VSS 0.353747f
C15686 DVSS.n7403 VSS 0.353747f
C15687 DVSS.n7404 VSS 0.353747f
C15688 DVSS.n7405 VSS 0.353747f
C15689 DVSS.n7406 VSS 0.282749f
C15690 DVSS.n7407 VSS 0.353747f
C15691 DVSS.n7408 VSS 0.353747f
C15692 DVSS.n7409 VSS 0.353747f
C15693 DVSS.n7410 VSS 0.353747f
C15694 DVSS.n7411 VSS 0.353747f
C15695 DVSS.n7412 VSS 0.353747f
C15696 DVSS.n7413 VSS 0.353747f
C15697 DVSS.n7414 VSS 0.315134f
C15698 DVSS.n7415 VSS 0.154453f
C15699 DVSS.n7417 VSS 0.176874f
C15700 DVSS.n7418 VSS 0.044926f
C15701 DVSS.n7419 VSS 0.176874f
C15702 DVSS.n7420 VSS 0.154453f
C15703 DVSS.n7421 VSS 0.353747f
C15704 DVSS.n7422 VSS 0.353747f
C15705 DVSS.n7423 VSS 0.353747f
C15706 DVSS.n7424 VSS 0.353747f
C15707 DVSS.n7425 VSS 0.353747f
C15708 DVSS.n7426 VSS 0.282749f
C15709 DVSS.n7427 VSS 0.353747f
C15710 DVSS.n7428 VSS 0.353747f
C15711 DVSS.n7429 VSS 0.353747f
C15712 DVSS.n7430 VSS 0.353747f
C15713 DVSS.n7431 VSS 0.353747f
C15714 DVSS.n7432 VSS 0.353747f
C15715 DVSS.n7433 VSS 0.353747f
C15716 DVSS.n7434 VSS 0.353747f
C15717 DVSS.n7435 VSS 0.353747f
C15718 DVSS.n7436 VSS 0.353747f
C15719 DVSS.n7437 VSS 0.353747f
C15720 DVSS.n7438 VSS 0.353747f
C15721 DVSS.n7439 VSS 0.353747f
C15722 DVSS.n7440 VSS 0.353747f
C15723 DVSS.n7441 VSS 0.353747f
C15724 DVSS.n7442 VSS 0.353747f
C15725 DVSS.n7443 VSS 0.353747f
C15726 DVSS.n7444 VSS 0.353747f
C15727 DVSS.n7445 VSS 0.353747f
C15728 DVSS.n7446 VSS 0.353747f
C15729 DVSS.n7447 VSS 0.353747f
C15730 DVSS.n7448 VSS 0.353747f
C15731 DVSS.n7449 VSS 0.353747f
C15732 DVSS.n7450 VSS 0.315134f
C15733 DVSS.n7451 VSS 0.154453f
C15734 DVSS.n7452 VSS 0.176874f
C15735 DVSS.n7453 VSS 0.044926f
C15736 DVSS.n7454 VSS 0.176874f
C15737 DVSS.n7455 VSS 0.154453f
C15738 DVSS.n7456 VSS 0.353747f
C15739 DVSS.n7457 VSS 0.353747f
C15740 DVSS.n7458 VSS 0.353747f
C15741 DVSS.n7459 VSS 0.353747f
C15742 DVSS.n7460 VSS 0.353747f
C15743 DVSS.n7461 VSS 0.282749f
C15744 DVSS.n7462 VSS 0.353747f
C15745 DVSS.n7463 VSS 0.353747f
C15746 DVSS.n7464 VSS 0.353747f
C15747 DVSS.n7465 VSS 0.353747f
C15748 DVSS.n7466 VSS 0.353747f
C15749 DVSS.n7467 VSS 0.353747f
C15750 DVSS.n7468 VSS 0.353747f
C15751 DVSS.n7469 VSS 0.353747f
C15752 DVSS.n7470 VSS 0.353747f
C15753 DVSS.n7471 VSS 0.353747f
C15754 DVSS.n7472 VSS 0.353747f
C15755 DVSS.n7473 VSS 0.353747f
C15756 DVSS.n7474 VSS 0.353747f
C15757 DVSS.n7475 VSS 0.353747f
C15758 DVSS.n7476 VSS 0.353747f
C15759 DVSS.n7477 VSS 0.353747f
C15760 DVSS.n7478 VSS 0.353747f
C15761 DVSS.n7479 VSS 0.353747f
C15762 DVSS.n7480 VSS 0.353747f
C15763 DVSS.n7481 VSS 0.353747f
C15764 DVSS.n7482 VSS 0.353747f
C15765 DVSS.n7483 VSS 0.353747f
C15766 DVSS.n7484 VSS 0.353747f
C15767 DVSS.n7485 VSS 0.341291f
C15768 DVSS.n7486 VSS 0.154453f
C15769 DVSS.n7487 VSS 0.176874f
C15770 DVSS.n7488 VSS 0.037674f
C15771 DVSS.n7489 VSS 0.176874f
C15772 DVSS.n7490 VSS 0.154453f
C15773 DVSS.n7491 VSS 0.353747f
C15774 DVSS.n7492 VSS 0.353747f
C15775 DVSS.n7493 VSS 0.353747f
C15776 DVSS.n7494 VSS 0.353747f
C15777 DVSS.n7495 VSS 0.353747f
C15778 DVSS.n7496 VSS 0.239153f
C15779 DVSS.n7497 VSS 0.154453f
C15780 DVSS.n7498 VSS 0.176874f
C15781 DVSS.n7499 VSS 0.037674f
C15782 DVSS.n7500 VSS 0.176874f
C15783 DVSS.n7501 VSS 0.154453f
C15784 DVSS.n7502 VSS 0.353747f
C15785 DVSS.n7503 VSS 0.353747f
C15786 DVSS.n7504 VSS 0.353747f
C15787 DVSS.n7505 VSS 0.353747f
C15788 DVSS.n7506 VSS 0.353747f
C15789 DVSS.n7507 VSS 0.353747f
C15790 DVSS.n7508 VSS 0.353747f
C15791 DVSS.n7509 VSS 0.353747f
C15792 DVSS.n7510 VSS 0.353747f
C15793 DVSS.n7511 VSS 0.353747f
C15794 DVSS.n7512 VSS 0.353747f
C15795 DVSS.n7513 VSS 0.353747f
C15796 DVSS.n7514 VSS 0.353747f
C15797 DVSS.n7515 VSS 0.353747f
C15798 DVSS.n7516 VSS 0.353747f
C15799 DVSS.n7517 VSS 0.353747f
C15800 DVSS.n7518 VSS 0.353747f
C15801 DVSS.n7519 VSS 0.353747f
C15802 DVSS.n7520 VSS 0.353747f
C15803 DVSS.n7521 VSS 0.353747f
C15804 DVSS.n7522 VSS 0.353747f
C15805 DVSS.n7523 VSS 0.353747f
C15806 DVSS.n7524 VSS 0.353747f
C15807 DVSS.n7525 VSS 0.353747f
C15808 DVSS.n7526 VSS 0.353747f
C15809 DVSS.n7527 VSS 0.353747f
C15810 DVSS.n7528 VSS 0.353747f
C15811 DVSS.n7529 VSS 0.353747f
C15812 DVSS.n7530 VSS 0.353747f
C15813 DVSS.n7531 VSS 0.154453f
C15814 DVSS.n7532 VSS 0.052308f
C15815 DVSS.n7533 VSS 0.052308f
C15816 DVSS.n7534 VSS 0.052308f
C15817 DVSS.n7535 VSS 0.052308f
C15818 DVSS.n7536 VSS 0.052308f
C15819 DVSS.n7537 VSS 0.052308f
C15820 DVSS.n7538 VSS 0.052308f
C15821 DVSS.n7539 VSS 0.052308f
C15822 DVSS.n7540 VSS 0.052308f
C15823 DVSS.n7541 VSS 0.052308f
C15824 DVSS.n7542 VSS 0.154453f
C15825 DVSS.n7553 VSS 0.176874f
C15826 DVSS.n7555 VSS 0.052308f
C15827 DVSS.n7556 VSS 0.176874f
C15828 DVSS.n7557 VSS 0.044926f
C15829 DVSS.n7558 VSS 0.176874f
C15830 DVSS.n7559 VSS 0.154453f
C15831 DVSS.n7560 VSS 0.353747f
C15832 DVSS.n7561 VSS 0.353747f
C15833 DVSS.n7562 VSS 0.353747f
C15834 DVSS.n7563 VSS 0.353747f
C15835 DVSS.n7564 VSS 0.353747f
C15836 DVSS.n7565 VSS 0.353747f
C15837 DVSS.n7566 VSS 0.353747f
C15838 DVSS.n7567 VSS 0.353747f
C15839 DVSS.n7568 VSS 0.353747f
C15840 DVSS.n7569 VSS 0.353747f
C15841 DVSS.n7570 VSS 0.353747f
C15842 DVSS.n7571 VSS 0.353747f
C15843 DVSS.n7572 VSS 0.353747f
C15844 DVSS.n7573 VSS 0.353747f
C15845 DVSS.n7574 VSS 0.353747f
C15846 DVSS.n7575 VSS 0.353747f
C15847 DVSS.n7576 VSS 0.353747f
C15848 DVSS.n7577 VSS 0.353747f
C15849 DVSS.n7578 VSS 0.353747f
C15850 DVSS.n7579 VSS 0.353747f
C15851 DVSS.n7580 VSS 0.353747f
C15852 DVSS.n7581 VSS 0.353747f
C15853 DVSS.n7582 VSS 0.353747f
C15854 DVSS.n7583 VSS 0.353747f
C15855 DVSS.n7584 VSS 0.353747f
C15856 DVSS.n7585 VSS 0.353747f
C15857 DVSS.n7586 VSS 0.353747f
C15858 DVSS.n7587 VSS 0.353747f
C15859 DVSS.n7588 VSS 0.353747f
C15860 DVSS.n7589 VSS 0.154453f
C15861 DVSS.n7590 VSS 0.052308f
C15862 DVSS.n7591 VSS 0.052308f
C15863 DVSS.n7592 VSS 0.052308f
C15864 DVSS.n7593 VSS 0.052308f
C15865 DVSS.n7594 VSS 0.052308f
C15866 DVSS.n7595 VSS 0.052308f
C15867 DVSS.n7596 VSS 0.052308f
C15868 DVSS.n7597 VSS 0.052308f
C15869 DVSS.n7598 VSS 0.052308f
C15870 DVSS.n7599 VSS 0.052308f
C15871 DVSS.n7600 VSS 0.154453f
C15872 DVSS.n7611 VSS 0.176874f
C15873 DVSS.n7613 VSS 0.052308f
C15874 DVSS.n7614 VSS 0.176874f
C15875 DVSS.n7615 VSS 0.044926f
C15876 DVSS.n7616 VSS 0.176874f
C15877 DVSS.n7617 VSS 0.154453f
C15878 DVSS.n7618 VSS 0.353747f
C15879 DVSS.n7619 VSS 0.353747f
C15880 DVSS.n7620 VSS 0.353747f
C15881 DVSS.n7621 VSS 0.353747f
C15882 DVSS.n7622 VSS 0.353747f
C15883 DVSS.n7623 VSS 0.353747f
C15884 DVSS.n7624 VSS 0.353747f
C15885 DVSS.n7625 VSS 0.353747f
C15886 DVSS.n7626 VSS 0.353747f
C15887 DVSS.n7627 VSS 0.353747f
C15888 DVSS.n7628 VSS 0.353747f
C15889 DVSS.n7629 VSS 0.353747f
C15890 DVSS.n7630 VSS 0.353747f
C15891 DVSS.n7631 VSS 0.154453f
C15892 DVSS.n7632 VSS 0.052308f
C15893 DVSS.n7633 VSS 0.052308f
C15894 DVSS.n7634 VSS 0.052308f
C15895 DVSS.n7635 VSS 0.052308f
C15896 DVSS.n7636 VSS 0.052308f
C15897 DVSS.n7637 VSS 0.052308f
C15898 DVSS.n7638 VSS 0.052308f
C15899 DVSS.n7639 VSS 0.052308f
C15900 DVSS.n7640 VSS 0.052308f
C15901 DVSS.n7641 VSS 0.052308f
C15902 DVSS.n7642 VSS 0.154453f
C15903 DVSS.n7653 VSS 0.176874f
C15904 DVSS.n7655 VSS 0.052308f
C15905 DVSS.n7656 VSS 0.176874f
C15906 DVSS.n7657 VSS 0.044926f
C15907 DVSS.n7658 VSS 0.176874f
C15908 DVSS.n7659 VSS 0.154453f
C15909 DVSS.n7660 VSS 0.353747f
C15910 DVSS.n7661 VSS 0.353747f
C15911 DVSS.n7662 VSS 0.353747f
C15912 DVSS.n7663 VSS 0.353747f
C15913 DVSS.n7664 VSS 0.353747f
C15914 DVSS.n7665 VSS 0.353747f
C15915 DVSS.n7666 VSS 0.353747f
C15916 DVSS.n7667 VSS 0.353747f
C15917 DVSS.n7668 VSS 0.318871f
C15918 DVSS.n7669 VSS 0.318871f
C15919 DVSS.n7670 VSS 0.21175f
C15920 DVSS.n7671 VSS 0.039859f
C15921 DVSS.n7672 VSS 0.348765f
C15922 DVSS.n7673 VSS 1.32112f
C15923 DVSS.n7674 VSS 0.682774f
C15924 DVSS.n7675 VSS 0.154453f
C15925 DVSS.n7676 VSS 0.353747f
C15926 DVSS.n7677 VSS 0.353747f
C15927 DVSS.n7678 VSS 0.154453f
C15928 DVSS.n7689 VSS 0.176874f
C15929 DVSS.n7692 VSS 0.052308f
C15930 DVSS.n7693 VSS 0.176874f
C15931 DVSS.n7694 VSS 0.051675f
C15932 DVSS.n7695 VSS 0.048301f
C15933 DVSS.n7696 VSS 0.048967f
C15934 DVSS.n7697 VSS 0.045559f
C15935 DVSS.n7698 VSS 0.041971f
C15936 DVSS.n7699 VSS 0.764373f
C15937 DVSS.n7700 VSS 0.058114f
C15938 DVSS.n7701 VSS 0.045559f
C15939 DVSS.n7702 VSS 0.045559f
C15940 DVSS.n7704 VSS 0.16051f
C15941 DVSS.n7705 VSS 0.041971f
C15942 DVSS.n7707 VSS 0.764373f
C15943 DVSS.n7708 VSS 0.048967f
C15944 DVSS.n7709 VSS 0.331802f
C15945 DVSS.n7711 VSS 0.157135f
C15946 DVSS.n7713 VSS 0.066724f
C15947 DVSS.n7714 VSS 0.052308f
C15948 DVSS.n7715 VSS 0.222771f
C15949 DVSS.n7716 VSS 0.754249f
C15950 DVSS.n7718 VSS 0.179185f
C15951 DVSS.n7720 VSS 0.066724f
C15952 DVSS.n7721 VSS 0.052308f
C15953 DVSS.n7722 VSS 0.09309f
C15954 DVSS.n7723 VSS 0.754249f
C15955 DVSS.n7725 VSS 0.335771f
C15956 DVSS.n7726 VSS 0.756156f
C15957 DVSS.n7729 VSS 0.082541f
C15958 DVSS.n7730 VSS 0.082541f
C15959 DVSS.n7731 VSS 0.134274f
C15960 DVSS.n7732 VSS 0.052308f
C15961 DVSS.n7733 VSS 0.052308f
C15962 DVSS.n7734 VSS 0.052308f
C15963 DVSS.n7735 VSS 0.052308f
C15964 DVSS.n7736 VSS 0.052308f
C15965 DVSS.n7737 VSS 0.072078f
C15966 DVSS.n7739 VSS 0.052308f
C15967 DVSS.n7741 VSS 0.052308f
C15968 DVSS.n7743 VSS 0.052308f
C15969 DVSS.n7745 VSS 0.052308f
C15970 DVSS.n7751 VSS 0.165082f
C15971 DVSS.n7752 VSS 0.072078f
C15972 DVSS.n7753 VSS 0.165082f
C15973 DVSS.n7754 VSS 0.165082f
C15974 DVSS.n7755 VSS 0.165082f
C15975 DVSS.n7756 VSS 0.165082f
C15976 DVSS.n7757 VSS 0.165082f
C15977 DVSS.n7758 VSS 0.165082f
C15978 DVSS.n7759 VSS 0.165082f
C15979 DVSS.n7760 VSS 0.165082f
C15980 DVSS.n7761 VSS 0.165082f
C15981 DVSS.n7762 VSS 0.165082f
C15982 DVSS.n7763 VSS 0.165082f
C15983 DVSS.n7764 VSS 0.156944f
C15984 DVSS.n7765 VSS 0.165082f
C15985 DVSS.n7766 VSS 0.165082f
C15986 DVSS.n7767 VSS 0.165082f
C15987 DVSS.n7768 VSS 0.165082f
C15988 DVSS.n7769 VSS 0.165082f
C15989 DVSS.n7770 VSS 0.072078f
C15990 DVSS.n7771 VSS 0.165082f
C15991 DVSS.n7772 VSS 0.165082f
C15992 DVSS.n7773 VSS 0.165082f
C15993 DVSS.n7774 VSS 0.165082f
C15994 DVSS.n7775 VSS 0.165082f
C15995 DVSS.n7776 VSS 0.165082f
C15996 DVSS.n7777 VSS 0.165082f
C15997 DVSS.n7778 VSS 0.165082f
C15998 DVSS.n7779 VSS 0.165082f
C15999 DVSS.n7780 VSS 0.165082f
C16000 DVSS.n7781 VSS 0.165082f
C16001 DVSS.n7782 VSS 0.165082f
C16002 DVSS.n7783 VSS 0.165082f
C16003 DVSS.n7784 VSS 0.165082f
C16004 DVSS.n7785 VSS 0.165082f
C16005 DVSS.n7786 VSS 0.165082f
C16006 DVSS.n7787 VSS 0.165082f
C16007 DVSS.n7788 VSS 0.165082f
C16008 DVSS.n7789 VSS 0.165082f
C16009 DVSS.n7790 VSS 0.165082f
C16010 DVSS.n7791 VSS 0.165082f
C16011 DVSS.n7792 VSS 0.165082f
C16012 DVSS.n7793 VSS 0.165082f
C16013 DVSS.n7794 VSS 0.165082f
C16014 DVSS.n7795 VSS 0.165082f
C16015 DVSS.n7796 VSS 0.165082f
C16016 DVSS.n7797 VSS 0.165082f
C16017 DVSS.n7798 VSS 0.165082f
C16018 DVSS.n7799 VSS 0.165082f
C16019 DVSS.n7800 VSS 0.165082f
C16020 DVSS.n7801 VSS 0.165082f
C16021 DVSS.n7802 VSS 0.165082f
C16022 DVSS.n7803 VSS 0.165082f
C16023 DVSS.n7804 VSS 0.165082f
C16024 DVSS.n7805 VSS 0.165082f
C16025 DVSS.n7806 VSS 0.165082f
C16026 DVSS.n7807 VSS 0.165082f
C16027 DVSS.n7808 VSS 0.165082f
C16028 DVSS.n7809 VSS 0.165082f
C16029 DVSS.n7810 VSS 0.165082f
C16030 DVSS.n7811 VSS 0.165082f
C16031 DVSS.n7812 VSS 0.165082f
C16032 DVSS.n7813 VSS 0.165082f
C16033 DVSS.n7814 VSS 0.165082f
C16034 DVSS.n7815 VSS 0.165082f
C16035 DVSS.n7816 VSS 0.165082f
C16036 DVSS.n7817 VSS 0.165082f
C16037 DVSS.n7818 VSS 0.165082f
C16038 DVSS.n7819 VSS 0.165082f
C16039 DVSS.n7820 VSS 0.165082f
C16040 DVSS.n7821 VSS 0.165082f
C16041 DVSS.n7822 VSS 0.165082f
C16042 DVSS.n7823 VSS 0.165082f
C16043 DVSS.n7824 VSS 0.165082f
C16044 DVSS.n7825 VSS 0.165082f
C16045 DVSS.n7826 VSS 0.165082f
C16046 DVSS.n7827 VSS 0.165082f
C16047 DVSS.n7828 VSS 0.165082f
C16048 DVSS.n7829 VSS 0.165082f
C16049 DVSS.n7830 VSS 0.165082f
C16050 DVSS.n7831 VSS 0.165082f
C16051 DVSS.n7832 VSS 0.165082f
C16052 DVSS.n7833 VSS 0.165082f
C16053 DVSS.n7834 VSS 0.165082f
C16054 DVSS.n7835 VSS 0.165082f
C16055 DVSS.n7836 VSS 0.165082f
C16056 DVSS.n7837 VSS 0.144737f
C16057 DVSS.n7838 VSS 0.165082f
C16058 DVSS.n7839 VSS 0.165082f
C16059 DVSS.n7840 VSS 0.165082f
C16060 DVSS.n7841 VSS 0.165082f
C16061 DVSS.n7842 VSS 0.165082f
C16062 DVSS.n7843 VSS 0.072078f
C16063 DVSS.n7844 VSS 0.082541f
C16064 DVSS.n7845 VSS 0.361727f
C16065 DVSS.n7846 VSS 0.082541f
C16066 DVSS.n7847 VSS 0.157135f
C16067 DVSS.n7848 VSS 0.157135f
C16068 DVSS.n7850 VSS 0.066724f
C16069 DVSS.n7851 VSS 0.052308f
C16070 DVSS.n7852 VSS 0.242143f
C16071 DVSS.n7853 VSS 0.754249f
C16072 DVSS.n7855 VSS 0.186719f
C16073 DVSS.n7856 VSS 0.043865f
C16074 DVSS.n7859 VSS 0.043865f
C16075 DVSS.n7860 VSS 0.396845f
C16076 DVSS.n7861 VSS 0.069335f
C16077 DVSS.n7862 VSS 0.066505f
C16078 DVSS.n7863 VSS 0.038205f
C16079 DVSS.n7864 VSS 0.038205f
C16080 DVSS.n7865 VSS 0.035873f
C16081 DVSS.n7866 VSS 0.038205f
C16082 DVSS.n7867 VSS 0.038205f
C16083 DVSS.n7868 VSS 0.024232f
C16084 DVSS.n7869 VSS 0.035873f
C16085 DVSS.n7870 VSS 0.021932f
C16086 DVSS.n7871 VSS 0.021932f
C16087 DVSS.n7872 VSS 0.035873f
C16088 DVSS.n7873 VSS 0.021932f
C16089 DVSS.n7874 VSS 0.021932f
C16090 DVSS.n7875 VSS 0.035873f
C16091 DVSS.n7876 VSS 0.021932f
C16092 DVSS.n7877 VSS 0.021932f
C16093 DVSS.n7878 VSS 0.035873f
C16094 DVSS.n7879 VSS 0.021932f
C16095 DVSS.n7880 VSS 0.021932f
C16096 DVSS.n7881 VSS 0.035873f
C16097 DVSS.n7882 VSS 0.035873f
C16098 DVSS.n7883 VSS 0.021755f
C16099 DVSS.n7884 VSS 0.019279f
C16100 DVSS.n7885 VSS 0.021755f
C16101 DVSS.n7886 VSS 0.019279f
C16102 DVSS.n7887 VSS 0.035873f
C16103 DVSS.n7888 VSS 0.021932f
C16104 DVSS.n7889 VSS 0.021932f
C16105 DVSS.n7890 VSS 0.035873f
C16106 DVSS.n7891 VSS 0.021932f
C16107 DVSS.n7892 VSS 0.021932f
C16108 DVSS.n7893 VSS 0.035873f
C16109 DVSS.n7894 VSS 0.021932f
C16110 DVSS.n7895 VSS 0.035873f
C16111 DVSS.t16 VSS 0.330478f
C16112 DVSS.n7896 VSS 0.125906f
C16113 DVSS.n7897 VSS 0.021932f
C16114 DVSS.n7898 VSS 0.026905f
C16115 DVSS.n7899 VSS 0.021932f
C16116 DVSS.n7900 VSS 0.019102f
C16117 DVSS.n7901 VSS 0.082541f
C16118 DVSS.n7902 VSS 0.019102f
C16119 DVSS.n7903 VSS 0.023878f
C16120 DVSS.n7904 VSS 0.038205f
C16121 DVSS.n7905 VSS 0.038205f
C16122 DVSS.n7906 VSS 0.035873f
C16123 DVSS.n7907 VSS 0.038205f
C16124 DVSS.n7908 VSS 0.038205f
C16125 DVSS.n7909 VSS 0.038205f
C16126 DVSS.n7910 VSS 0.038205f
C16127 DVSS.n7911 VSS 0.038205f
C16128 DVSS.n7912 VSS 0.035873f
C16129 DVSS.n7913 VSS 0.038205f
C16130 DVSS.n7914 VSS 0.038205f
C16131 DVSS.n7915 VSS 0.038205f
C16132 DVSS.n7916 VSS 0.038205f
C16133 DVSS.n7917 VSS 0.038205f
C16134 DVSS.n7918 VSS 0.038205f
C16135 DVSS.n7919 VSS 0.035873f
C16136 DVSS.n7920 VSS 0.035873f
C16137 DVSS.n7921 VSS 0.035873f
C16138 DVSS.n7922 VSS 0.038205f
C16139 DVSS.n7923 VSS 0.038205f
C16140 DVSS.n7924 VSS 0.038205f
C16141 DVSS.n7925 VSS 0.035873f
C16142 DVSS.n7926 VSS 0.035873f
C16143 DVSS.n7927 VSS 0.035873f
C16144 DVSS.n7928 VSS 0.038205f
C16145 DVSS.n7929 VSS 0.038205f
C16146 DVSS.n7930 VSS 0.038205f
C16147 DVSS.n7931 VSS 0.035873f
C16148 DVSS.n7932 VSS 0.033714f
C16149 DVSS.n7933 VSS 0.020096f
C16150 DVSS.n7934 VSS 0.023878f
C16151 DVSS.n7935 VSS 0.019102f
C16152 DVSS.n7936 VSS 0.082541f
C16153 DVSS.n7937 VSS 0.072078f
C16154 DVSS.n7938 VSS 0.165082f
C16155 DVSS.n7939 VSS 0.165082f
C16156 DVSS.n7940 VSS 0.165082f
C16157 DVSS.n7941 VSS 0.165082f
C16158 DVSS.n7942 VSS 0.165082f
C16159 DVSS.n7943 VSS 0.159269f
C16160 DVSS.n7944 VSS 0.165082f
C16161 DVSS.n7945 VSS 0.165082f
C16162 DVSS.n7946 VSS 0.165082f
C16163 DVSS.n7947 VSS 0.165082f
C16164 DVSS.n7948 VSS 0.165082f
C16165 DVSS.n7949 VSS 0.165082f
C16166 DVSS.n7950 VSS 0.165082f
C16167 DVSS.n7951 VSS 0.165082f
C16168 DVSS.n7952 VSS 0.165082f
C16169 DVSS.n7953 VSS 0.165082f
C16170 DVSS.n7954 VSS 0.165082f
C16171 DVSS.n7955 VSS 0.165082f
C16172 DVSS.n7956 VSS 0.165082f
C16173 DVSS.n7957 VSS 0.165082f
C16174 DVSS.n7958 VSS 0.165082f
C16175 DVSS.n7959 VSS 0.165082f
C16176 DVSS.n7960 VSS 0.165082f
C16177 DVSS.n7961 VSS 0.165082f
C16178 DVSS.n7962 VSS 0.165082f
C16179 DVSS.n7963 VSS 0.165082f
C16180 DVSS.n7964 VSS 0.165082f
C16181 DVSS.n7965 VSS 0.165082f
C16182 DVSS.n7966 VSS 0.165082f
C16183 DVSS.n7967 VSS 0.131949f
C16184 DVSS.n7972 VSS 0.082541f
C16185 DVSS.n7974 VSS 0.361727f
C16186 DVSS.n7975 VSS 0.082541f
C16187 DVSS.n7976 VSS 0.072078f
C16188 DVSS.n7977 VSS 0.165082f
C16189 DVSS.n7978 VSS 0.165082f
C16190 DVSS.n7979 VSS 0.165082f
C16191 DVSS.n7980 VSS 0.165082f
C16192 DVSS.n7981 VSS 0.165082f
C16193 DVSS.n7982 VSS 0.147063f
C16194 DVSS.n7983 VSS 0.165082f
C16195 DVSS.n7984 VSS 0.165082f
C16196 DVSS.n7985 VSS 0.165082f
C16197 DVSS.n7986 VSS 0.165082f
C16198 DVSS.n7987 VSS 0.165082f
C16199 DVSS.n7988 VSS 0.165082f
C16200 DVSS.n7989 VSS 0.165082f
C16201 DVSS.n7990 VSS 0.165082f
C16202 DVSS.n7991 VSS 0.165082f
C16203 DVSS.n7992 VSS 0.165082f
C16204 DVSS.n7993 VSS 0.165082f
C16205 DVSS.n7994 VSS 0.165082f
C16206 DVSS.n7995 VSS 0.165082f
C16207 DVSS.n7996 VSS 0.165082f
C16208 DVSS.n7997 VSS 0.165082f
C16209 DVSS.n7998 VSS 0.165082f
C16210 DVSS.n7999 VSS 0.165082f
C16211 DVSS.n8000 VSS 0.165082f
C16212 DVSS.n8001 VSS 0.165082f
C16213 DVSS.n8002 VSS 0.165082f
C16214 DVSS.n8003 VSS 0.165082f
C16215 DVSS.n8004 VSS 0.165082f
C16216 DVSS.n8005 VSS 0.165082f
C16217 DVSS.n8006 VSS 0.131949f
C16218 DVSS.n8011 VSS 0.082541f
C16219 DVSS.n8013 VSS 0.361727f
C16220 DVSS.n8014 VSS 0.082541f
C16221 DVSS.n8015 VSS 0.072078f
C16222 DVSS.n8016 VSS 0.165082f
C16223 DVSS.n8017 VSS 0.165082f
C16224 DVSS.n8018 VSS 0.165082f
C16225 DVSS.n8019 VSS 0.165082f
C16226 DVSS.n8020 VSS 0.165082f
C16227 DVSS.n8021 VSS 0.147063f
C16228 DVSS.n8022 VSS 0.165082f
C16229 DVSS.n8023 VSS 0.165082f
C16230 DVSS.n8024 VSS 0.165082f
C16231 DVSS.n8025 VSS 0.165082f
C16232 DVSS.n8026 VSS 0.165082f
C16233 DVSS.n8027 VSS 0.165082f
C16234 DVSS.n8028 VSS 0.165082f
C16235 DVSS.n8029 VSS 0.131949f
C16236 DVSS.n8034 VSS 0.082541f
C16237 DVSS.n8036 VSS 0.361727f
C16238 DVSS.n8037 VSS 0.082541f
C16239 DVSS.n8038 VSS 0.072078f
C16240 DVSS.n8039 VSS 0.165082f
C16241 DVSS.n8040 VSS 0.165082f
C16242 DVSS.n8041 VSS 0.165082f
C16243 DVSS.n8042 VSS 0.165082f
C16244 DVSS.n8043 VSS 0.165082f
C16245 DVSS.n8044 VSS 0.147063f
C16246 DVSS.n8045 VSS 0.165082f
C16247 DVSS.n8046 VSS 0.165082f
C16248 DVSS.n8047 VSS 0.165082f
C16249 DVSS.n8048 VSS 0.165082f
C16250 DVSS.n8049 VSS 0.165082f
C16251 DVSS.n8050 VSS 0.165082f
C16252 DVSS.n8051 VSS 0.165082f
C16253 DVSS.n8052 VSS 0.131949f
C16254 DVSS.n8056 VSS 0.082541f
C16255 DVSS.n8059 VSS 0.052308f
C16256 DVSS.n8060 VSS 0.361112f
C16257 DVSS.n8061 VSS 0.368477f
C16258 DVSS.n8062 VSS 0.365102f
C16259 DVSS.n8065 VSS 0.058114f
C16260 DVSS.n8067 VSS 0.041971f
C16261 DVSS.n8068 VSS 0.756569f
C16262 DVSS.n8069 VSS 0.048967f
C16263 DVSS.n8070 VSS 0.331802f
C16264 DVSS.n8072 VSS 0.222771f
C16265 DVSS.n8074 VSS 0.066724f
C16266 DVSS.n8075 VSS 0.052308f
C16267 DVSS.n8076 VSS 0.179185f
C16268 DVSS.n8078 VSS 0.09309f
C16269 DVSS.n8080 VSS 0.066724f
C16270 DVSS.n8081 VSS 0.052308f
C16271 DVSS.n8082 VSS 0.335771f
C16272 DVSS.n8083 VSS 0.756156f
C16273 DVSS.n8085 VSS 0.242143f
C16274 DVSS.n8087 VSS 0.066724f
C16275 DVSS.n8088 VSS 0.052308f
C16276 DVSS.n8089 VSS 0.186719f
C16277 DVSS.n8090 VSS 0.396845f
C16278 DVSS.n8092 VSS 0.043865f
C16279 DVSS.n8093 VSS 0.065379f
C16280 DVSS.n8095 VSS 0.069335f
C16281 DVSS.n8096 VSS 0.066505f
C16282 DVSS.n8097 VSS 0.049824f
C16283 DVSS.n8098 VSS 0.066505f
C16284 DVSS.n8099 VSS 0.069335f
C16285 DVSS.n8101 VSS 0.043865f
C16286 DVSS.n8102 VSS 0.065379f
C16287 DVSS.n8104 VSS 0.043865f
C16288 DVSS.n8105 VSS 0.396845f
C16289 DVSS.n8107 VSS 0.186719f
C16290 DVSS.n8109 VSS 0.066724f
C16291 DVSS.n8110 VSS 0.052308f
C16292 DVSS.n8111 VSS 0.242143f
C16293 DVSS.n8112 VSS 0.756156f
C16294 DVSS.n8114 VSS 0.335771f
C16295 DVSS.n8116 VSS 0.066724f
C16296 DVSS.n8117 VSS 0.052308f
C16297 DVSS.n8118 VSS 0.09309f
C16298 DVSS.n8119 VSS 0.361727f
C16299 DVSS.n8120 VSS 0.361727f
C16300 DVSS.n8121 VSS 0.082541f
C16301 DVSS.n8122 VSS 0.157135f
C16302 DVSS.n8123 VSS 0.082541f
C16303 DVSS.n8124 VSS 0.072078f
C16304 DVSS.n8125 VSS 0.165082f
C16305 DVSS.n8126 VSS 0.165082f
C16306 DVSS.n8127 VSS 0.165082f
C16307 DVSS.n8128 VSS 0.165082f
C16308 DVSS.n8129 VSS 0.165082f
C16309 DVSS.n8130 VSS 0.165082f
C16310 DVSS.n8131 VSS 0.165082f
C16311 DVSS.n8132 VSS 0.165082f
C16312 DVSS.n8133 VSS 0.165082f
C16313 DVSS.n8134 VSS 0.165082f
C16314 DVSS.n8135 VSS 0.165082f
C16315 DVSS.n8136 VSS 0.165082f
C16316 DVSS.n8137 VSS 0.165082f
C16317 DVSS.n8138 VSS 0.072078f
C16318 DVSS.n8139 VSS 0.052308f
C16319 DVSS.n8140 VSS 0.052308f
C16320 DVSS.n8144 VSS 0.072078f
C16321 DVSS.n8145 VSS 0.082541f
C16322 DVSS.n8147 VSS 0.052308f
C16323 DVSS.n8148 VSS 0.052308f
C16324 DVSS.n8149 VSS 0.082541f
C16325 DVSS.n8150 VSS 0.052308f
C16326 DVSS.n8152 VSS 0.082541f
C16327 DVSS.n8153 VSS 0.072078f
C16328 DVSS.n8154 VSS 0.165082f
C16329 DVSS.n8155 VSS 0.165082f
C16330 DVSS.n8156 VSS 0.165082f
C16331 DVSS.n8157 VSS 0.165082f
C16332 DVSS.n8158 VSS 0.165082f
C16333 DVSS.n8159 VSS 0.165082f
C16334 DVSS.n8160 VSS 0.165082f
C16335 DVSS.n8161 VSS 0.148806f
C16336 DVSS.n8162 VSS 0.148806f
C16337 DVSS.n8163 VSS 0.165082f
C16338 DVSS.n8164 VSS 0.084866f
C16339 DVSS.n8165 VSS 0.098817f
C16340 DVSS.n8166 VSS 0.165082f
C16341 DVSS.n8167 VSS 0.072078f
C16342 DVSS.n8168 VSS 0.165082f
C16343 DVSS.n8169 VSS 0.616179f
C16344 DVSS.n8170 VSS 0.319361f
C16345 DVSS.n8174 VSS 0.363609f
C16346 DVSS.n8177 VSS 0.052308f
C16347 DVSS.n8178 VSS 0.082541f
C16348 DVSS.n8179 VSS 0.368477f
C16349 DVSS.n8180 VSS 0.365102f
C16350 DVSS.n8181 VSS 0.048967f
C16351 DVSS.n8183 VSS 0.756569f
C16352 DVSS.n8184 VSS 0.041971f
C16353 DVSS.n8185 VSS 0.217854f
C16354 DVSS.n8186 VSS 0.133296f
C16355 DVSS.n8187 VSS 0.032106f
C16356 DVSS.n8189 VSS 0.045559f
C16357 DVSS.n8191 VSS 0.027052f
C16358 DVSS.n8192 VSS 0.233666f
C16359 DVSS.n8193 VSS 0.116237f
C16360 DVSS.n8194 VSS 0.74982f
C16361 DVSS.n8196 VSS 0.032106f
C16362 DVSS.n8197 VSS 0.032106f
C16363 DVSS.n8198 VSS 1.58569f
C16364 DVSS.n8199 VSS 0.092157f
C16365 DVSS.n8200 VSS 0.044592f
C16366 DVSS.n8201 VSS 0.74982f
C16367 DVSS.n8203 VSS 0.032106f
C16368 DVSS.n8204 VSS 0.032106f
C16369 DVSS.n8205 VSS 1.42561f
C16370 DVSS.n8206 VSS 0.148938f
C16371 DVSS.n8207 VSS 0.548192f
C16372 DVSS.n8208 VSS 0.097211f
C16373 DVSS.n8209 VSS 0.045559f
C16374 DVSS.n8210 VSS 0.096319f
C16375 DVSS.n8211 VSS 0.297397f
C16376 DVSS.n8212 VSS 0.297397f
C16377 DVSS.n8213 VSS 0.019909f
C16378 DVSS.n8214 VSS 0.019909f
C16379 DVSS.n8215 VSS 0.009955f
C16380 DVSS.n8216 VSS 0.157979f
C16381 DVSS.n8217 VSS 0.180752f
C16382 DVSS.n8218 VSS 0.180752f
C16383 DVSS.n8219 VSS 0.132478f
C16384 DVSS.n8220 VSS 0.017421f
C16385 DVSS.n8221 VSS 0.014932f
C16386 DVSS.n8222 VSS 0.017421f
C16387 DVSS.n8223 VSS 0.132478f
C16388 DVSS.n8224 VSS 0.132478f
C16389 DVSS.n8226 VSS 0.033721f
C16390 DVSS.n8228 VSS 0.033721f
C16391 DVSS.n8229 VSS 0.038205f
C16392 DVSS.n8231 VSS 0.306139f
C16393 DVSS.n8234 VSS 0.033721f
C16394 DVSS.n8235 VSS 0.033721f
C16395 DVSS.n8236 VSS 0.045559f
C16396 DVSS.n8237 VSS 0.306139f
C16397 DVSS.n8238 VSS 0.161143f
C16398 DVSS.n8239 VSS 0.161143f
C16399 DVSS.n8241 VSS 0.045559f
C16400 DVSS.n8243 VSS 0.267267f
C16401 DVSS.n8245 VSS 0.033721f
C16402 DVSS.n8246 VSS 0.033721f
C16403 DVSS.n8248 VSS 0.161143f
C16404 DVSS.n8249 VSS 0.306139f
C16405 DVSS.n8250 VSS 0.306139f
C16406 DVSS.n8252 VSS 0.033721f
C16407 DVSS.n8254 VSS 0.135131f
C16408 DVSS.n8255 VSS 0.029505f
C16409 DVSS.n8256 VSS 0.77032f
C16410 DVSS.n8257 VSS 1.41915f
C16411 DVSS.n8258 VSS 0.02529f
C16412 DVSS.n8259 VSS 0.029505f
C16413 DVSS.n8261 VSS 0.033721f
C16414 DVSS.n8263 VSS 0.045559f
C16415 DVSS.n8265 VSS 0.033721f
C16416 DVSS.n8266 VSS 0.033721f
C16417 DVSS.n8269 VSS 0.033721f
C16418 DVSS.n8270 VSS 0.328284f
C16419 DVSS.n8271 VSS 0.267267f
C16420 DVSS.n8272 VSS 0.161143f
C16421 DVSS.n8273 VSS 0.306139f
C16422 DVSS.n8274 VSS 0.306139f
C16423 DVSS.n8276 VSS 0.038205f
C16424 DVSS.n8278 VSS 0.033721f
C16425 DVSS.n8279 VSS 0.135131f
C16426 DVSS.n8280 VSS 0.135131f
C16427 DVSS.n8281 VSS 0.306139f
C16428 DVSS.n8282 VSS 0.038205f
C16429 DVSS.n8284 VSS 0.029505f
C16430 DVSS.n8285 VSS 1.41915f
C16431 DVSS.n8286 VSS 0.02529f
C16432 DVSS.n8287 VSS 0.029505f
C16433 DVSS.n8288 VSS 0.038205f
C16434 DVSS.n8290 VSS 0.306139f
C16435 DVSS.n8291 VSS 0.306139f
C16436 DVSS.n8292 VSS 0.157979f
C16437 DVSS.n8293 VSS 0.267267f
C16438 DVSS.n8294 VSS 0.330782f
C16439 DVSS.n8295 VSS 0.045718f
C16440 DVSS.n8296 VSS 0.04802f
C16441 DVSS.n8297 VSS 7.158741f
C16442 DVSS.n8298 VSS 0.04802f
C16443 DVSS.n8299 VSS 0.797916f
C16444 DVSS.n8300 VSS 1.41915f
C16445 DVSS.n8301 VSS 0.02529f
C16446 DVSS.n8302 VSS 0.029505f
C16447 DVSS.n8304 VSS 0.033721f
C16448 DVSS.n8306 VSS 0.135131f
C16449 DVSS.n8307 VSS 0.306139f
C16450 DVSS.n8308 VSS 0.306139f
C16451 DVSS.n8310 VSS 0.033721f
C16452 DVSS.n8311 VSS 0.033721f
C16453 DVSS.n8313 VSS 0.161143f
C16454 DVSS.n8314 VSS 0.267267f
C16455 DVSS.n8315 VSS 0.330782f
C16456 DVSS.n8316 VSS 0.211948f
C16457 DVSS.n8317 VSS 0.507231f
C16458 DVSS.n8318 VSS 7.158741f
C16459 DVSS.n8319 VSS 0.507231f
C16460 DVSS.n8320 VSS 0.211948f
C16461 DVSS.n8321 VSS 0.330782f
C16462 DVSS.n8324 VSS 0.033721f
C16463 DVSS.n8325 VSS 0.033721f
C16464 DVSS.n8326 VSS 0.045559f
C16465 DVSS.n8327 VSS 0.267267f
C16466 DVSS.n8328 VSS 0.157979f
C16467 DVSS.n8329 VSS 0.009955f
C16468 DVSS.n8330 VSS 0.009955f
C16469 DVSS.n8331 VSS 0.157979f
C16470 DVSS.n8333 VSS 0.421629f
C16471 DVSS.n8334 VSS 0.019909f
C16472 DVSS.n8335 VSS 0.019909f
C16473 DVSS.n8336 VSS 0.421629f
C16474 DVSS.n8337 VSS 0.009955f
C16475 DVSS.n8338 VSS 0.180752f
C16476 DVSS.n8339 VSS 0.160088f
C16477 DVSS.n8341 VSS 0.163463f
C16478 DVSS.n8344 VSS 0.052308f
C16479 DVSS.n8347 VSS 0.052308f
C16480 DVSS.n8348 VSS 0.082541f
C16481 DVSS.n8349 VSS 0.022779f
C16482 DVSS.n8350 VSS 0.026154f
C16483 DVSS.n8352 VSS 0.033721f
C16484 DVSS.n8353 VSS 0.025732f
C16485 DVSS.n8354 VSS 0.306139f
C16486 DVSS.n8355 VSS 0.306139f
C16487 DVSS.n8356 VSS 0.033721f
C16488 DVSS.n8358 VSS 0.021932f
C16489 DVSS.n8360 VSS 0.033721f
C16490 DVSS.n8362 VSS 0.026154f
C16491 DVSS.n8364 VSS 0.033721f
C16492 DVSS.n8366 VSS 0.033721f
C16493 DVSS.n8367 VSS 0.023201f
C16494 DVSS.n8368 VSS 0.033721f
C16495 DVSS.n8370 VSS 0.30411f
C16496 DVSS.n8371 VSS 0.025732f
C16497 DVSS.n8372 VSS 0.306139f
C16498 DVSS.n8373 VSS 0.019456f
C16499 DVSS.n8375 VSS 0.033721f
C16500 DVSS.n8376 VSS 0.306139f
C16501 DVSS.n8377 VSS 0.021579f
C16502 DVSS.n8378 VSS 0.029505f
C16503 DVSS.n8379 VSS 1.75989f
C16504 DVSS.n8380 VSS 0.02529f
C16505 DVSS.n8382 VSS 0.019456f
C16506 DVSS.n8384 VSS 0.033721f
C16507 DVSS.n8385 VSS 0.029505f
C16508 DVSS.n8386 VSS 0.021579f
C16509 DVSS.n8387 VSS 0.024409f
C16510 DVSS.n8388 VSS 0.082541f
C16511 DVSS.n8389 VSS 0.043865f
C16512 DVSS.n8391 VSS 0.025116f
C16513 DVSS.n8392 VSS 0.082541f
C16514 DVSS.n8393 VSS 0.072078f
C16515 DVSS.n8394 VSS 0.165082f
C16516 DVSS.n8395 VSS 0.165082f
C16517 DVSS.n8396 VSS 0.165082f
C16518 DVSS.n8397 VSS 0.165082f
C16519 DVSS.n8398 VSS 0.165082f
C16520 DVSS.n8399 VSS 0.10928f
C16521 DVSS.n8400 VSS 0.082541f
C16522 DVSS.n8402 VSS 0.141853f
C16523 DVSS.n8403 VSS 0.082541f
C16524 DVSS.n8404 VSS 0.159269f
C16525 DVSS.n8405 VSS 0.165082f
C16526 DVSS.n8406 VSS 0.165082f
C16527 DVSS.n8407 VSS 0.165082f
C16528 DVSS.n8408 VSS 0.165082f
C16529 DVSS.n8409 VSS 0.165082f
C16530 DVSS.n8410 VSS 0.165082f
C16531 DVSS.n8411 VSS 0.165082f
C16532 DVSS.n8412 VSS 0.165082f
C16533 DVSS.n8413 VSS 0.165082f
C16534 DVSS.n8414 VSS 0.165082f
C16535 DVSS.n8415 VSS 0.165082f
C16536 DVSS.n8416 VSS 0.165082f
C16537 DVSS.n8417 VSS 0.165082f
C16538 DVSS.n8418 VSS 0.165082f
C16539 DVSS.n8419 VSS 0.165082f
C16540 DVSS.n8420 VSS 0.165082f
C16541 DVSS.n8421 VSS 0.165082f
C16542 DVSS.n8422 VSS 0.165082f
C16543 DVSS.n8423 VSS 0.165082f
C16544 DVSS.n8424 VSS 0.165082f
C16545 DVSS.n8425 VSS 0.165082f
C16546 DVSS.n8426 VSS 0.165082f
C16547 DVSS.n8427 VSS 0.165082f
C16548 DVSS.n8428 VSS 0.131949f
C16549 DVSS.n8429 VSS 0.165082f
C16550 DVSS.n8430 VSS 0.165082f
C16551 DVSS.n8431 VSS 0.165082f
C16552 DVSS.n8432 VSS 0.165082f
C16553 DVSS.n8433 VSS 0.165082f
C16554 DVSS.n8434 VSS 0.072078f
C16555 DVSS.n8435 VSS 0.082541f
C16556 DVSS.n8438 VSS 0.052308f
C16557 DVSS.n8439 VSS 0.082541f
C16558 DVSS.n8440 VSS 0.169158f
C16559 DVSS.n8442 VSS 0.165783f
C16560 DVSS.n8444 VSS 0.045559f
C16561 DVSS.n8446 VSS 0.033721f
C16562 DVSS.n8447 VSS 0.246354f
C16563 DVSS.n8448 VSS 0.30411f
C16564 DVSS.n8449 VSS 0.30411f
C16565 DVSS.n8450 VSS 0.165783f
C16566 DVSS.n8451 VSS 0.169158f
C16567 DVSS.n8452 VSS 0.082541f
C16568 DVSS.n8453 VSS 0.022779f
C16569 DVSS.n8454 VSS 0.026154f
C16570 DVSS.n8456 VSS 0.033721f
C16571 DVSS.n8457 VSS 0.025732f
C16572 DVSS.n8458 VSS 0.07353f
C16573 DVSS.n8459 VSS 0.186081f
C16574 DVSS.n8460 VSS 0.136683f
C16575 DVSS.n8461 VSS 0.663966f
C16576 DVSS.n8462 VSS 13.1085f
C16577 DVSS.n8463 VSS 0.101916f
C16578 DVSS.n8464 VSS 0.994586f
C16579 DVSS.n8465 VSS 0.994586f
C16580 DVSS.n8466 VSS 1.75989f
C16581 DVSS.n8467 VSS 0.02529f
C16582 DVSS.n8468 VSS 0.029505f
C16583 DVSS.n8469 VSS 0.033721f
C16584 DVSS.n8470 VSS 0.206588f
C16585 DVSS.n8472 VSS 0.033721f
C16586 DVSS.n8474 VSS 0.139023f
C16587 DVSS.n8475 VSS 0.306139f
C16588 DVSS.n8476 VSS 0.306139f
C16589 DVSS.n8477 VSS 0.246354f
C16590 DVSS.n8478 VSS 0.033721f
C16591 DVSS.n8479 VSS 0.165783f
C16592 DVSS.n8480 VSS 0.30411f
C16593 DVSS.n8481 VSS 0.246354f
C16594 DVSS.n8482 VSS 0.30411f
C16595 DVSS.n8483 VSS 0.045559f
C16596 DVSS.n8484 VSS 0.094754f
C16597 DVSS.n8485 VSS 0.182276f
C16598 DVSS.n8486 VSS 0.07353f
C16599 DVSS.n8487 VSS 0.165783f
C16600 DVSS.n8488 VSS 0.169158f
C16601 DVSS.n8489 VSS 0.082541f
C16602 DVSS.n8490 VSS 0.022779f
C16603 DVSS.n8491 VSS 0.023201f
C16604 DVSS.n8492 VSS 0.033721f
C16605 DVSS.n8494 VSS 0.30411f
C16606 DVSS.n8495 VSS 0.025732f
C16607 DVSS.n8496 VSS 0.07353f
C16608 DVSS.n8497 VSS 0.186081f
C16609 DVSS.n8498 VSS 0.136683f
C16610 DVSS.n8499 VSS 0.663966f
C16611 DVSS.n8500 VSS 13.1085f
C16612 DVSS.n8501 VSS 0.663966f
C16613 DVSS.n8502 VSS 0.136683f
C16614 DVSS.n8503 VSS 0.102784f
C16615 DVSS.n8504 VSS 0.026154f
C16616 DVSS.n8505 VSS 0.019909f
C16617 DVSS.n8506 VSS 0.019909f
C16618 DVSS.n8507 VSS 0.026154f
C16619 DVSS.n8508 VSS 0.179554f
C16620 DVSS.n8509 VSS 0.179554f
C16621 DVSS.n8510 VSS 0.026154f
C16622 DVSS.n8511 VSS 0.019909f
C16623 DVSS.n8512 VSS 0.019909f
C16624 DVSS.n8513 VSS 0.026154f
C16625 DVSS.n8514 VSS 0.180752f
C16626 DVSS.n8515 VSS 0.180752f
C16627 DVSS.n8516 VSS 0.009955f
C16628 DVSS.n8517 VSS 0.019909f
C16629 DVSS.n8518 VSS 0.009955f
C16630 DVSS.n8519 VSS 0.017421f
C16631 DVSS.n8520 VSS 0.014932f
C16632 DVSS.n8521 VSS 0.017421f
C16633 DVSS.n8522 VSS 0.021932f
C16634 DVSS.n8523 VSS 0.009955f
C16635 DVSS.n8524 VSS 0.019909f
C16636 DVSS.n8525 VSS 0.021932f
C16637 DVSS.n8526 VSS 0.180752f
C16638 DVSS.n8527 VSS 0.180752f
C16639 DVSS.n8528 VSS 0.009955f
C16640 DVSS.n8529 VSS 0.019909f
C16641 DVSS.n8530 VSS 0.009955f
C16642 DVSS.n8531 VSS 0.019909f
C16643 DVSS.n8532 VSS 0.026154f
C16644 DVSS.n8534 VSS 0.176874f
C16645 DVSS.n8535 VSS 0.052308f
C16646 DVSS.n8536 VSS 0.052308f
C16647 DVSS.n8537 VSS 0.052308f
C16648 DVSS.n8538 VSS 0.030583f
C16649 DVSS.n8539 VSS 0.052308f
C16650 DVSS.n8540 VSS 0.052308f
C16651 DVSS.n8541 VSS 0.052308f
C16652 DVSS.n8542 VSS 0.154453f
C16653 DVSS.n8544 VSS 0.052308f
C16654 DVSS.n8546 VSS 0.052308f
C16655 DVSS.n8548 VSS 0.052308f
C16656 DVSS.n8550 VSS 0.052308f
C16657 DVSS.n8552 VSS 0.052308f
C16658 DVSS.n8554 VSS 0.052308f
C16659 DVSS.n8556 VSS 0.052308f
C16660 DVSS.n8558 VSS 0.052308f
C16661 DVSS.n8559 VSS 0.176874f
C16662 DVSS.n8560 VSS 0.022779f
C16663 DVSS.n8561 VSS 0.176874f
C16664 DVSS.n8562 VSS 0.282749f
C16665 DVSS.n8563 VSS 0.353747f
C16666 DVSS.n8564 VSS 0.353747f
C16667 DVSS.n8565 VSS 0.353747f
C16668 DVSS.n8566 VSS 0.353747f
C16669 DVSS.n8567 VSS 0.353747f
C16670 DVSS.n8568 VSS 0.353747f
C16671 DVSS.n8569 VSS 0.353747f
C16672 DVSS.n8570 VSS 0.353747f
C16673 DVSS.n8571 VSS 0.353747f
C16674 DVSS.n8572 VSS 0.353747f
C16675 DVSS.n8573 VSS 0.353747f
C16676 DVSS.n8574 VSS 0.353747f
C16677 DVSS.n8575 VSS 0.353747f
C16678 DVSS.n8576 VSS 0.353747f
C16679 DVSS.n8577 VSS 0.353747f
C16680 DVSS.n8578 VSS 0.353747f
C16681 DVSS.n8579 VSS 0.353747f
C16682 DVSS.n8580 VSS 0.353747f
C16683 DVSS.n8581 VSS 0.353747f
C16684 DVSS.n8582 VSS 0.353747f
C16685 DVSS.n8583 VSS 0.353747f
C16686 DVSS.n8584 VSS 0.353747f
C16687 DVSS.n8585 VSS 0.353747f
C16688 DVSS.n8586 VSS 0.353747f
C16689 DVSS.n8587 VSS 0.353747f
C16690 DVSS.n8588 VSS 0.353747f
C16691 DVSS.n8589 VSS 0.353747f
C16692 DVSS.n8590 VSS 0.353747f
C16693 DVSS.n8591 VSS 0.353747f
C16694 DVSS.n8592 VSS 0.353747f
C16695 DVSS.n8593 VSS 0.353747f
C16696 DVSS.n8594 VSS 0.353747f
C16697 DVSS.n8595 VSS 0.353747f
C16698 DVSS.n8596 VSS 0.353747f
C16699 DVSS.n8597 VSS 0.293959f
C16700 DVSS.n8598 VSS 0.293959f
C16701 DVSS.n8599 VSS 0.425991f
C16702 DVSS.n8600 VSS 0.675109f
C16703 DVSS.n8601 VSS 0.236662f
C16704 DVSS.n8602 VSS 0.236662f
C16705 DVSS.n8603 VSS 0.353747f
C16706 DVSS.n8604 VSS 0.353747f
C16707 DVSS.n8605 VSS 0.353747f
C16708 DVSS.n8606 VSS 0.353747f
C16709 DVSS.n8607 VSS 0.353747f
C16710 DVSS.n8608 VSS 0.353747f
C16711 DVSS.n8609 VSS 0.353747f
C16712 DVSS.n8610 VSS 0.353747f
C16713 DVSS.n8611 VSS 0.353747f
C16714 DVSS.n8612 VSS 0.353747f
C16715 DVSS.n8613 VSS 0.353747f
C16716 DVSS.n8614 VSS 0.353747f
C16717 DVSS.n8615 VSS 0.353747f
C16718 DVSS.n8616 VSS 0.353747f
C16719 DVSS.n8617 VSS 0.353747f
C16720 DVSS.n8618 VSS 0.353747f
C16721 DVSS.n8619 VSS 0.353747f
C16722 DVSS.n8620 VSS 0.353747f
C16723 DVSS.n8621 VSS 1.31155f
C16724 DVSS.n8622 VSS 0.353747f
C16725 DVSS.n8623 VSS 0.154453f
C16726 DVSS.n8634 VSS 0.176874f
C16727 DVSS.n8637 VSS 0.052308f
C16728 DVSS.n8638 VSS 0.776799f
C16729 DVSS.n8639 VSS 0.099554f
C16730 DVSS.n8640 VSS 0.099554f
C16731 DVSS.n8642 VSS 0.670635f
C16732 DVSS.n8643 VSS 0.052308f
C16733 DVSS.n8644 VSS 0.052308f
C16734 DVSS.n8645 VSS 0.052308f
C16735 DVSS.n8646 VSS 0.052308f
C16736 DVSS.n8647 VSS 0.052308f
C16737 DVSS.n8648 VSS 0.052308f
C16738 DVSS.n8649 VSS 0.052308f
C16739 DVSS.n8650 VSS 0.052308f
C16740 DVSS.n8651 VSS 0.052308f
C16741 DVSS.n8652 VSS 0.052308f
C16742 DVSS.n8653 VSS 0.052308f
C16743 DVSS.n8654 VSS 0.353747f
C16744 DVSS.n8655 VSS 0.154453f
C16745 DVSS.n8656 VSS 0.052308f
C16746 DVSS.n8657 VSS 0.052308f
C16747 DVSS.n8658 VSS 0.052308f
C16748 DVSS.n8659 VSS 0.052308f
C16749 DVSS.n8660 VSS 0.052308f
C16750 DVSS.n8661 VSS 0.052308f
C16751 DVSS.n8662 VSS 0.052308f
C16752 DVSS.n8663 VSS 0.052308f
C16753 DVSS.n8664 VSS 0.052308f
C16754 DVSS.n8665 VSS 0.052308f
C16755 DVSS.n8666 VSS 0.154453f
C16756 DVSS.n8677 VSS 0.176874f
C16757 DVSS.n8679 VSS 0.052308f
C16758 DVSS.n8680 VSS 0.776799f
C16759 DVSS.n8681 VSS 0.22484f
C16760 DVSS.n8682 VSS 0.176874f
C16761 DVSS.n8683 VSS 0.154453f
C16762 DVSS.n8684 VSS 0.353747f
C16763 DVSS.n8685 VSS 0.353747f
C16764 DVSS.n8686 VSS 0.353747f
C16765 DVSS.n8687 VSS 0.353747f
C16766 DVSS.n8688 VSS 0.353747f
C16767 DVSS.n8689 VSS 0.353747f
C16768 DVSS.n8690 VSS 0.353747f
C16769 DVSS.n8691 VSS 0.315134f
C16770 DVSS.n8692 VSS 0.353747f
C16771 DVSS.n8693 VSS 0.353747f
C16772 DVSS.n8694 VSS 0.353747f
C16773 DVSS.n8695 VSS 0.353747f
C16774 DVSS.n8696 VSS 0.353747f
C16775 DVSS.n8697 VSS 0.353747f
C16776 DVSS.n8698 VSS 0.154453f
C16777 DVSS.n8699 VSS 0.353747f
C16778 DVSS.n8700 VSS 0.353747f
C16779 DVSS.n8701 VSS 0.353747f
C16780 DVSS.n8702 VSS 0.353747f
C16781 DVSS.n8703 VSS 0.353747f
C16782 DVSS.n8704 VSS 0.353747f
C16783 DVSS.n8705 VSS 0.353747f
C16784 DVSS.n8706 VSS 0.353747f
C16785 DVSS.n8707 VSS 0.236662f
C16786 DVSS.n8708 VSS 0.236662f
C16787 DVSS.n8709 VSS 0.236662f
C16788 DVSS.n8710 VSS 0.425991f
C16789 DVSS.n8711 VSS 0.293959f
C16790 DVSS.n8712 VSS 0.293959f
C16791 DVSS.n8713 VSS 0.255346f
C16792 DVSS.n8714 VSS 0.154453f
C16793 DVSS.n8715 VSS 0.176874f
C16794 DVSS.n8716 VSS 0.052308f
C16795 DVSS.n8717 VSS 0.176874f
C16796 DVSS.n8718 VSS 0.154453f
C16797 DVSS.n8719 VSS 0.353747f
C16798 DVSS.n8720 VSS 0.353747f
C16799 DVSS.n8721 VSS 0.353747f
C16800 DVSS.n8722 VSS 0.353747f
C16801 DVSS.n8723 VSS 0.353747f
C16802 DVSS.n8724 VSS 0.282749f
C16803 DVSS.n8725 VSS 0.353747f
C16804 DVSS.n8726 VSS 0.353747f
C16805 DVSS.n8727 VSS 0.353747f
C16806 DVSS.n8728 VSS 0.353747f
C16807 DVSS.n8729 VSS 0.353747f
C16808 DVSS.n8730 VSS 0.353747f
C16809 DVSS.n8731 VSS 0.353747f
C16810 DVSS.n8732 VSS 0.353747f
C16811 DVSS.n8733 VSS 0.353747f
C16812 DVSS.n8734 VSS 0.353747f
C16813 DVSS.n8735 VSS 0.353747f
C16814 DVSS.n8736 VSS 0.353747f
C16815 DVSS.n8737 VSS 0.353747f
C16816 DVSS.n8738 VSS 0.353747f
C16817 DVSS.n8739 VSS 0.353747f
C16818 DVSS.n8740 VSS 0.353747f
C16819 DVSS.n8741 VSS 0.353747f
C16820 DVSS.n8742 VSS 0.353747f
C16821 DVSS.n8743 VSS 0.353747f
C16822 DVSS.n8744 VSS 0.353747f
C16823 DVSS.n8745 VSS 0.353747f
C16824 DVSS.n8746 VSS 0.353747f
C16825 DVSS.n8747 VSS 0.353747f
C16826 DVSS.n8748 VSS 0.315134f
C16827 DVSS.n8749 VSS 0.154453f
C16828 DVSS.n8750 VSS 0.176874f
C16829 DVSS.n8751 VSS 0.052308f
C16830 DVSS.n8752 VSS 0.176874f
C16831 DVSS.n8753 VSS 0.154453f
C16832 DVSS.n8754 VSS 0.353747f
C16833 DVSS.n8755 VSS 0.353747f
C16834 DVSS.n8756 VSS 0.353747f
C16835 DVSS.n8757 VSS 0.353747f
C16836 DVSS.n8758 VSS 0.353747f
C16837 DVSS.n8759 VSS 0.353747f
C16838 DVSS.n8760 VSS 0.282749f
C16839 DVSS.n8761 VSS 0.353747f
C16840 DVSS.n8762 VSS 0.353747f
C16841 DVSS.n8763 VSS 0.353747f
C16842 DVSS.n8764 VSS 0.226697f
C16843 DVSS.n8765 VSS 0.226697f
C16844 DVSS.n8766 VSS 0.425991f
C16845 DVSS.n8767 VSS 0.353747f
C16846 DVSS.n8768 VSS 0.353747f
C16847 DVSS.n8769 VSS 0.353747f
C16848 DVSS.n8770 VSS 0.353747f
C16849 DVSS.n8771 VSS 0.353747f
C16850 DVSS.n8772 VSS 0.353747f
C16851 DVSS.n8773 VSS 0.353747f
C16852 DVSS.n8774 VSS 0.353747f
C16853 DVSS.n8775 VSS 0.353747f
C16854 DVSS.n8776 VSS 0.353747f
C16855 DVSS.n8777 VSS 0.353747f
C16856 DVSS.n8788 VSS 0.176874f
C16857 DVSS.n8789 VSS 0.154453f
C16858 DVSS.n8790 VSS 0.239153f
C16859 DVSS.n8791 VSS 0.234171f
C16860 DVSS.n8792 VSS 0.353747f
C16861 DVSS.n8793 VSS 0.353747f
C16862 DVSS.n8794 VSS 0.353747f
C16863 DVSS.n8795 VSS 0.353747f
C16864 DVSS.n8796 VSS 0.353747f
C16865 DVSS.n8797 VSS 0.353747f
C16866 DVSS.n8798 VSS 0.353747f
C16867 DVSS.n8799 VSS 0.353747f
C16868 DVSS.n8800 VSS 0.353747f
C16869 DVSS.n8801 VSS 0.353747f
C16870 DVSS.n8802 VSS 0.353747f
C16871 DVSS.n8803 VSS 0.353747f
C16872 DVSS.n8804 VSS 0.353747f
C16873 DVSS.n8805 VSS 0.353747f
C16874 DVSS.n8806 VSS 0.353747f
C16875 DVSS.n8807 VSS 0.353747f
C16876 DVSS.n8808 VSS 0.303924f
C16877 DVSS.n8809 VSS 0.303924f
C16878 DVSS.n8810 VSS 0.303924f
C16879 DVSS.n8811 VSS 0.425991f
C16880 DVSS.n8812 VSS 0.425991f
C16881 DVSS.n8813 VSS 0.675109f
C16882 DVSS.n8814 VSS 0.226697f
C16883 DVSS.n8815 VSS 0.353747f
C16884 DVSS.n8816 VSS 0.226697f
C16885 DVSS.n8817 VSS 0.353747f
C16886 DVSS.n8818 VSS 0.353747f
C16887 DVSS.n8819 VSS 0.353747f
C16888 DVSS.n8820 VSS 0.353747f
C16889 DVSS.n8821 VSS 0.353747f
C16890 DVSS.n8822 VSS 0.353747f
C16891 DVSS.n8823 VSS 0.353747f
C16892 DVSS.n8824 VSS 0.353747f
C16893 DVSS.n8825 VSS 0.154453f
C16894 DVSS.n8826 VSS 0.052308f
C16895 DVSS.n8827 VSS 0.052308f
C16896 DVSS.n8828 VSS 0.052308f
C16897 DVSS.n8829 VSS 0.052308f
C16898 DVSS.n8830 VSS 0.052308f
C16899 DVSS.n8831 VSS 0.052308f
C16900 DVSS.n8832 VSS 0.052308f
C16901 DVSS.n8833 VSS 0.052308f
C16902 DVSS.n8834 VSS 0.052308f
C16903 DVSS.n8836 VSS 0.052308f
C16904 DVSS.n8838 VSS 0.052308f
C16905 DVSS.n8840 VSS 0.052308f
C16906 DVSS.n8842 VSS 0.052308f
C16907 DVSS.n8844 VSS 0.052308f
C16908 DVSS.n8846 VSS 0.052308f
C16909 DVSS.n8848 VSS 0.052308f
C16910 DVSS.n8850 VSS 0.052308f
C16911 DVSS.n8852 VSS 0.052308f
C16912 DVSS.n8854 VSS 0.052308f
C16913 DVSS.n8855 VSS 0.052308f
C16914 DVSS.n8856 VSS 0.176874f
C16915 DVSS.n8857 VSS 0.052308f
C16916 DVSS.n8859 VSS 0.176874f
C16917 DVSS.n8860 VSS 0.031427f
C16918 DVSS.n8861 VSS 0.031427f
C16919 DVSS.n8862 VSS 0.026354f
C16920 DVSS.n8865 VSS 0.048189f
C16921 DVSS.n8867 VSS 0.043865f
C16922 DVSS.n8869 VSS 0.397368f
C16923 DVSS.n8870 VSS 0.397368f
C16924 DVSS.n8871 VSS 0.052308f
C16925 DVSS.n8872 VSS 0.048189f
C16926 DVSS.n8873 VSS 0.026154f
C16927 DVSS.n8874 VSS 0.393287f
C16928 DVSS.n8875 VSS 0.393287f
C16929 DVSS.n8876 VSS 0.052308f
C16930 DVSS.n8877 VSS 0.048189f
C16931 DVSS.n8878 VSS 0.026154f
C16932 DVSS.n8879 VSS 0.173326f
C16933 DVSS.n8880 VSS 0.042395f
C16934 DVSS.n8882 VSS 0.045559f
C16935 DVSS.n8883 VSS 0.170217f
C16936 DVSS.n8884 VSS 0.026154f
C16937 DVSS.n8885 VSS 0.029924f
C16938 DVSS.n8886 VSS 0.029924f
C16939 DVSS.n8887 VSS 0.026154f
C16940 DVSS.n8888 VSS 0.029924f
C16941 DVSS.n8889 VSS 0.026154f
C16942 DVSS.n8890 VSS 0.041971f
C16943 DVSS.n8891 VSS 0.026154f
C16944 DVSS.n8892 VSS 0.041971f
C16945 DVSS.n8893 VSS 0.026154f
C16946 DVSS.n8894 VSS 0.041971f
C16947 DVSS.n8895 VSS 0.041971f
C16948 DVSS.n8896 VSS 0.023834f
C16949 DVSS.n8897 VSS 0.025099f
C16950 DVSS.n8898 VSS 0.041971f
C16951 DVSS.n8899 VSS 0.026154f
C16952 DVSS.n8900 VSS 0.041971f
C16953 DVSS.n8901 VSS 0.026154f
C16954 DVSS.n8902 VSS 0.041971f
C16955 DVSS.n8903 VSS 0.026154f
C16956 DVSS.n8904 VSS 0.041971f
C16957 DVSS.n8905 VSS 0.026154f
C16958 DVSS.n8906 VSS 0.041971f
C16959 DVSS.n8907 VSS 0.026154f
C16960 DVSS.n8908 VSS 0.041971f
C16961 DVSS.n8909 VSS 0.026154f
C16962 DVSS.n8910 VSS 0.041971f
C16963 DVSS.n8911 VSS 0.041971f
C16964 DVSS.n8912 VSS 0.02299f
C16965 DVSS.n8913 VSS 0.025943f
C16966 DVSS.n8914 VSS 0.041971f
C16967 DVSS.n8915 VSS 0.026154f
C16968 DVSS.n8916 VSS 0.041971f
C16969 DVSS.n8917 VSS 0.026154f
C16970 DVSS.n8918 VSS 0.041971f
C16971 DVSS.n8919 VSS 0.026154f
C16972 DVSS.n8920 VSS 0.041971f
C16973 DVSS.n8921 VSS 0.026154f
C16974 DVSS.n8922 VSS 0.041971f
C16975 DVSS.n8923 VSS 0.026154f
C16976 DVSS.n8924 VSS 0.041971f
C16977 DVSS.n8925 VSS 0.041971f
C16978 DVSS.n8926 VSS 0.025521f
C16979 DVSS.n8927 VSS 0.023412f
C16980 DVSS.n8928 VSS 0.041971f
C16981 DVSS.n8929 VSS 0.026154f
C16982 DVSS.n8930 VSS 0.041971f
C16983 DVSS.n8931 VSS 0.026154f
C16984 DVSS.n8932 VSS 0.041971f
C16985 DVSS.n8933 VSS 0.041971f
C16986 DVSS.n8934 VSS 0.026154f
C16987 DVSS.n8935 VSS 0.026154f
C16988 DVSS.n8936 VSS 0.022779f
C16989 DVSS.n8937 VSS 0.176874f
C16990 DVSS.n8938 VSS 0.022779f
C16991 DVSS.n8939 VSS 0.026154f
C16992 DVSS.n8940 VSS 0.041971f
C16993 DVSS.n8941 VSS 0.041971f
C16994 DVSS.n8942 VSS 0.031479f
C16995 DVSS.n8943 VSS 0.045559f
C16996 DVSS.n8944 VSS 0.045348f
C16997 DVSS.n8945 VSS 0.031479f
C16998 DVSS.n8946 VSS 0.041971f
C16999 DVSS.n8947 VSS 0.02299f
C17000 DVSS.n8948 VSS 0.025943f
C17001 DVSS.n8949 VSS 0.041971f
C17002 DVSS.n8950 VSS 0.026154f
C17003 DVSS.n8951 VSS 0.041971f
C17004 DVSS.n8952 VSS 0.026154f
C17005 DVSS.n8953 VSS 0.041971f
C17006 DVSS.n8954 VSS 0.026154f
C17007 DVSS.n8955 VSS 0.041971f
C17008 DVSS.n8956 VSS 0.026154f
C17009 DVSS.n8957 VSS 0.041971f
C17010 DVSS.n8958 VSS 0.026154f
C17011 DVSS.n8959 VSS 0.041971f
C17012 DVSS.n8960 VSS 0.041971f
C17013 DVSS.n8961 VSS 0.025521f
C17014 DVSS.n8962 VSS 0.023412f
C17015 DVSS.n8963 VSS 0.041971f
C17016 DVSS.n8964 VSS 0.026154f
C17017 DVSS.n8965 VSS 0.041971f
C17018 DVSS.n8966 VSS 0.026154f
C17019 DVSS.n8967 VSS 0.041971f
C17020 DVSS.n8968 VSS 0.026154f
C17021 DVSS.n8969 VSS 0.041971f
C17022 DVSS.n8970 VSS 0.026154f
C17023 DVSS.n8971 VSS 0.041971f
C17024 DVSS.n8972 VSS 0.026154f
C17025 DVSS.n8973 VSS 0.041971f
C17026 DVSS.n8974 VSS 0.026154f
C17027 DVSS.n8975 VSS 0.041971f
C17028 DVSS.n8976 VSS 0.041971f
C17029 DVSS.n8977 VSS 0.024678f
C17030 DVSS.n8978 VSS 0.024256f
C17031 DVSS.n8979 VSS 0.041971f
C17032 DVSS.n8980 VSS 0.026154f
C17033 DVSS.n8981 VSS 0.041971f
C17034 DVSS.n8982 VSS 0.026154f
C17035 DVSS.n8983 VSS 0.041971f
C17036 DVSS.n8984 VSS 0.026154f
C17037 DVSS.n8985 VSS 0.041971f
C17038 DVSS.n8986 VSS 0.026154f
C17039 DVSS.n8987 VSS 0.041971f
C17040 DVSS.n8988 VSS 0.026154f
C17041 DVSS.n8989 VSS 0.041971f
C17042 DVSS.n8990 VSS 0.026154f
C17043 DVSS.n8991 VSS 0.041971f
C17044 DVSS.n8992 VSS 0.041971f
C17045 DVSS.n8993 VSS 0.041971f
C17046 DVSS.n8994 VSS 0.025099f
C17047 DVSS.n8995 VSS 0.022779f
C17048 DVSS.n8996 VSS 0.176874f
C17049 DVSS.n8997 VSS 0.022779f
C17050 DVSS.n8998 VSS 0.026154f
C17051 DVSS.n8999 VSS 0.029924f
C17052 DVSS.n9000 VSS 0.029924f
C17053 DVSS.n9002 VSS 0.078891f
C17054 DVSS.n9003 VSS 0.036489f
C17055 DVSS.n9004 VSS 0.170217f
C17056 DVSS.n9006 VSS 0.173326f
C17057 DVSS.n9008 VSS 0.048189f
C17058 DVSS.n9009 VSS 0.036911f
C17059 DVSS.n9010 VSS 0.393287f
C17060 DVSS.n9012 VSS 0.393287f
C17061 DVSS.n9014 VSS 0.048189f
C17062 DVSS.n9015 VSS 0.036911f
C17063 DVSS.n9016 VSS 0.397368f
C17064 DVSS.n9017 VSS 0.038912f
C17065 DVSS.n9018 VSS 0.048189f
C17066 DVSS.n9019 VSS 0.043865f
C17067 DVSS.n9021 VSS 0.043865f
C17068 DVSS.n9023 VSS 0.397368f
C17069 DVSS.n9024 VSS 0.030953f
C17070 DVSS.n9025 VSS 0.030953f
C17071 DVSS.n9026 VSS 0.176874f
C17072 DVSS.n9027 VSS 0.083484f
C17073 DVSS.n9028 VSS 0.043865f
C17074 DVSS.n9029 VSS 0.043865f
C17075 DVSS.n9030 VSS 0.043865f
C17076 DVSS.n9031 VSS 0.043865f
C17077 DVSS.n9032 VSS 0.043865f
C17078 DVSS.n9033 VSS 0.043865f
C17079 DVSS.n9034 VSS 0.043865f
C17080 DVSS.n9035 VSS 0.043865f
C17081 DVSS.n9036 VSS 0.043865f
C17082 DVSS.n9037 VSS 0.043865f
C17083 DVSS.n9038 VSS 0.043865f
C17084 DVSS.n9039 VSS 0.154453f
C17085 DVSS.n9040 VSS 0.043865f
C17086 DVSS.n9041 VSS 0.043865f
C17087 DVSS.n9042 VSS 0.043865f
C17088 DVSS.n9043 VSS 0.043865f
C17089 DVSS.n9044 VSS 0.043865f
C17090 DVSS.n9045 VSS 0.043865f
C17091 DVSS.n9046 VSS 0.043865f
C17092 DVSS.n9047 VSS 0.043865f
C17093 DVSS.n9048 VSS 0.043865f
C17094 DVSS.n9049 VSS 0.043865f
C17095 DVSS.n9060 VSS 0.176874f
C17096 DVSS.n9062 VSS 0.043865f
C17097 DVSS.n9063 VSS 0.176874f
C17098 DVSS.n9064 VSS 0.083484f
C17099 DVSS.n9065 VSS 0.176874f
C17100 DVSS.n9066 VSS 0.234171f
C17101 DVSS.n9067 VSS 0.353747f
C17102 DVSS.n9068 VSS 0.353747f
C17103 DVSS.n9069 VSS 0.353747f
C17104 DVSS.n9070 VSS 0.353747f
C17105 DVSS.n9071 VSS 0.353747f
C17106 DVSS.n9072 VSS 0.353747f
C17107 DVSS.n9073 VSS 0.353747f
C17108 DVSS.n9074 VSS 0.353747f
C17109 DVSS.n9075 VSS 0.353747f
C17110 DVSS.n9076 VSS 0.353747f
C17111 DVSS.n9077 VSS 0.353747f
C17112 DVSS.n9078 VSS 0.353747f
C17113 DVSS.n9079 VSS 0.353747f
C17114 DVSS.n9080 VSS 0.353747f
C17115 DVSS.n9081 VSS 0.353747f
C17116 DVSS.n9082 VSS 0.353747f
C17117 DVSS.n9083 VSS 0.353747f
C17118 DVSS.n9084 VSS 0.353747f
C17119 DVSS.n9085 VSS 0.303924f
C17120 DVSS.n9086 VSS 0.303924f
C17121 DVSS.n9087 VSS 0.675109f
C17122 DVSS.n9088 VSS 0.425991f
C17123 DVSS.n9089 VSS 0.226697f
C17124 DVSS.n9090 VSS 0.226697f
C17125 DVSS.n9091 VSS 0.425991f
C17126 DVSS.n9092 VSS 0.303924f
C17127 DVSS.n9093 VSS 0.353747f
C17128 DVSS.n9094 VSS 0.353747f
C17129 DVSS.n9095 VSS 0.353747f
C17130 DVSS.n9096 VSS 0.353747f
C17131 DVSS.n9097 VSS 0.353747f
C17132 DVSS.n9098 VSS 0.353747f
C17133 DVSS.n9099 VSS 0.353747f
C17134 DVSS.n9100 VSS 0.353747f
C17135 DVSS.n9101 VSS 0.353747f
C17136 DVSS.n9102 VSS 0.353747f
C17137 DVSS.n9103 VSS 0.353747f
C17138 DVSS.n9104 VSS 0.353747f
C17139 DVSS.n9105 VSS 0.353747f
C17140 DVSS.n9106 VSS 0.353747f
C17141 DVSS.n9107 VSS 0.353747f
C17142 DVSS.n9108 VSS 0.353747f
C17143 DVSS.n9109 VSS 0.353747f
C17144 DVSS.n9110 VSS 0.353747f
C17145 DVSS.n9111 VSS 0.154453f
C17146 DVSS.n9113 VSS 0.043865f
C17147 DVSS.n9115 VSS 0.043865f
C17148 DVSS.n9117 VSS 0.043865f
C17149 DVSS.n9119 VSS 0.043865f
C17150 DVSS.n9121 VSS 0.043865f
C17151 DVSS.n9123 VSS 0.043865f
C17152 DVSS.n9125 VSS 0.043865f
C17153 DVSS.n9127 VSS 0.043865f
C17154 DVSS.n9128 VSS 0.176874f
C17155 DVSS.n9129 VSS 0.021932f
C17156 DVSS.n9130 VSS 0.176874f
C17157 DVSS.n9131 VSS 0.234171f
C17158 DVSS.n9132 VSS 0.353747f
C17159 DVSS.n9133 VSS 0.353747f
C17160 DVSS.n9134 VSS 0.353747f
C17161 DVSS.n9135 VSS 0.353747f
C17162 DVSS.n9136 VSS 0.353747f
C17163 DVSS.n9137 VSS 0.353747f
C17164 DVSS.n9138 VSS 0.154453f
C17165 DVSS.n9139 VSS 0.043865f
C17166 DVSS.n9140 VSS 0.043865f
C17167 DVSS.n9141 VSS 0.043865f
C17168 DVSS.n9142 VSS 0.043865f
C17169 DVSS.n9143 VSS 0.043865f
C17170 DVSS.n9144 VSS 0.043865f
C17171 DVSS.n9153 VSS 0.176874f
C17172 DVSS.n9155 VSS 0.043865f
C17173 DVSS.n9156 VSS 0.176874f
C17174 DVSS.n9157 VSS 0.043865f
C17175 DVSS.n9159 VSS 0.176874f
C17176 DVSS.n9160 VSS 0.336309f
C17177 DVSS.n9161 VSS 0.353747f
C17178 DVSS.n9162 VSS 0.353747f
C17179 DVSS.n9163 VSS 0.353747f
C17180 DVSS.n9164 VSS 0.353747f
C17181 DVSS.n9165 VSS 0.353747f
C17182 DVSS.n9166 VSS 0.353747f
C17183 DVSS.n9167 VSS 0.353747f
C17184 DVSS.n9168 VSS 0.353747f
C17185 DVSS.n9169 VSS 0.353747f
C17186 DVSS.n9170 VSS 0.353747f
C17187 DVSS.n9171 VSS 0.353747f
C17188 DVSS.n9172 VSS 0.353747f
C17189 DVSS.n9173 VSS 0.353747f
C17190 DVSS.n9174 VSS 0.353747f
C17191 DVSS.n9175 VSS 0.353747f
C17192 DVSS.n9176 VSS 0.425991f
C17193 DVSS.n9177 VSS 0.216732f
C17194 DVSS.n9178 VSS 0.216732f
C17195 DVSS.n9179 VSS 0.425991f
C17196 DVSS.n9180 VSS 0.675109f
C17197 DVSS.n9181 VSS 0.216732f
C17198 DVSS.n9182 VSS 0.216732f
C17199 DVSS.n9183 VSS 0.353747f
C17200 DVSS.n9184 VSS 0.353747f
C17201 DVSS.n9185 VSS 0.353747f
C17202 DVSS.n9186 VSS 0.353747f
C17203 DVSS.n9187 VSS 0.353747f
C17204 DVSS.n9188 VSS 0.353747f
C17205 DVSS.n9189 VSS 0.353747f
C17206 DVSS.n9190 VSS 0.353747f
C17207 DVSS.n9191 VSS 0.353747f
C17208 DVSS.n9192 VSS 0.353747f
C17209 DVSS.n9193 VSS 0.353747f
C17210 DVSS.n9194 VSS 0.353747f
C17211 DVSS.n9195 VSS 0.353747f
C17212 DVSS.n9196 VSS 0.353747f
C17213 DVSS.n9197 VSS 0.154453f
C17214 DVSS.n9208 VSS 0.176874f
C17215 DVSS.n9211 VSS 0.043865f
C17216 DVSS.n9212 VSS 0.176874f
C17217 DVSS.n9213 VSS 0.083484f
C17218 DVSS.n9214 VSS 0.083484f
C17219 DVSS.n9216 VSS 0.043865f
C17220 DVSS.n9218 VSS 0.043865f
C17221 DVSS.n9220 VSS 0.043865f
C17222 DVSS.n9222 VSS 0.043865f
C17223 DVSS.n9224 VSS 0.043865f
C17224 DVSS.n9226 VSS 0.043865f
C17225 DVSS.n9228 VSS 0.043865f
C17226 DVSS.n9230 VSS 0.043865f
C17227 DVSS.n9232 VSS 0.043865f
C17228 DVSS.n9234 VSS 0.043865f
C17229 DVSS.n9236 VSS 0.043865f
C17230 DVSS.n9238 VSS 0.043865f
C17231 DVSS.n9240 VSS 0.043865f
C17232 DVSS.n9242 VSS 0.043865f
C17233 DVSS.n9244 VSS 0.043865f
C17234 DVSS.n9246 VSS 0.043865f
C17235 DVSS.n9248 VSS 0.043865f
C17236 DVSS.n9250 VSS 0.043865f
C17237 DVSS.n9252 VSS 0.043865f
C17238 DVSS.n9254 VSS 0.043865f
C17239 DVSS.n9256 VSS 0.043865f
C17240 DVSS.n9258 VSS 0.043865f
C17241 DVSS.n9260 VSS 0.176874f
C17242 DVSS.n9261 VSS 0.154453f
C17243 DVSS.n9262 VSS 0.353747f
C17244 DVSS.n9263 VSS 0.353747f
C17245 DVSS.n9264 VSS 0.353747f
C17246 DVSS.n9265 VSS 0.353747f
C17247 DVSS.n9266 VSS 0.353747f
C17248 DVSS.n9267 VSS 0.336309f
C17249 DVSS.n9268 VSS 0.353747f
C17250 DVSS.n9269 VSS 0.353747f
C17251 DVSS.n9270 VSS 0.353747f
C17252 DVSS.n9271 VSS 0.353747f
C17253 DVSS.n9272 VSS 0.353747f
C17254 DVSS.n9273 VSS 0.353747f
C17255 DVSS.n9274 VSS 0.353747f
C17256 DVSS.n9275 VSS 0.353747f
C17257 DVSS.n9276 VSS 0.353747f
C17258 DVSS.n9277 VSS 0.353747f
C17259 DVSS.n9278 VSS 0.353747f
C17260 DVSS.n9279 VSS 0.353747f
C17261 DVSS.n9280 VSS 0.353747f
C17262 DVSS.n9281 VSS 0.353747f
C17263 DVSS.n9282 VSS 0.216732f
C17264 DVSS.n9283 VSS 0.216732f
C17265 DVSS.n9284 VSS 0.425991f
C17266 DVSS.n9285 VSS 0.353747f
C17267 DVSS.n9286 VSS 0.313888f
C17268 DVSS.n9287 VSS 0.313888f
C17269 DVSS.n9288 VSS 0.313888f
C17270 DVSS.n9289 VSS 0.353747f
C17271 DVSS.n9290 VSS 0.353747f
C17272 DVSS.n9291 VSS 0.353747f
C17273 DVSS.n9292 VSS 0.353747f
C17274 DVSS.n9293 VSS 0.353747f
C17275 DVSS.n9294 VSS 0.353747f
C17276 DVSS.n9295 VSS 0.353747f
C17277 DVSS.n9296 VSS 0.310152f
C17278 DVSS.n9297 VSS 0.353747f
C17279 DVSS.n9298 VSS 0.353747f
C17280 DVSS.n9299 VSS 0.353747f
C17281 DVSS.n9300 VSS 0.353747f
C17282 DVSS.n9301 VSS 0.353747f
C17283 DVSS.n9302 VSS 0.353747f
C17284 DVSS.n9303 VSS 0.353747f
C17285 DVSS.n9304 VSS 0.353747f
C17286 DVSS.n9305 VSS 0.353747f
C17287 DVSS.n9306 VSS 0.353747f
C17288 DVSS.n9307 VSS 0.353747f
C17289 DVSS.n9308 VSS 0.353747f
C17290 DVSS.n9309 VSS 0.353747f
C17291 DVSS.n9310 VSS 0.353747f
C17292 DVSS.n9311 VSS 0.353747f
C17293 DVSS.n9312 VSS 0.353747f
C17294 DVSS.n9313 VSS 0.353747f
C17295 DVSS.n9324 VSS 0.176874f
C17296 DVSS.n9325 VSS 0.154453f
C17297 DVSS.n9326 VSS 0.353747f
C17298 DVSS.n9327 VSS 0.353747f
C17299 DVSS.n9328 VSS 0.353747f
C17300 DVSS.n9329 VSS 0.353747f
C17301 DVSS.n9330 VSS 0.353747f
C17302 DVSS.n9331 VSS 0.353747f
C17303 DVSS.n9332 VSS 0.353747f
C17304 DVSS.n9333 VSS 0.353747f
C17305 DVSS.n9334 VSS 0.353747f
C17306 DVSS.n9335 VSS 0.353747f
C17307 DVSS.n9336 VSS 0.353747f
C17308 DVSS.n9337 VSS 0.353747f
C17309 DVSS.n9338 VSS 0.353747f
C17310 DVSS.n9339 VSS 0.353747f
C17311 DVSS.n9340 VSS 0.353747f
C17312 DVSS.n9341 VSS 0.353747f
C17313 DVSS.n9342 VSS 0.353747f
C17314 DVSS.n9343 VSS 0.353747f
C17315 DVSS.n9344 VSS 0.353747f
C17316 DVSS.n9345 VSS 0.353747f
C17317 DVSS.n9346 VSS 0.353747f
C17318 DVSS.n9347 VSS 0.353747f
C17319 DVSS.n9348 VSS 0.353747f
C17320 DVSS.n9349 VSS 0.353747f
C17321 DVSS.n9350 VSS 0.353747f
C17322 DVSS.n9351 VSS 0.353747f
C17323 DVSS.n9352 VSS 0.154453f
C17324 DVSS.n9363 VSS 0.176874f
C17325 DVSS.n9366 VSS 0.052308f
C17326 DVSS.n9367 VSS 0.176874f
C17327 DVSS.n9368 VSS 0.036911f
C17328 DVSS.n9370 VSS 0.048189f
C17329 DVSS.n9371 VSS 0.048189f
C17330 DVSS.n9372 VSS 0.052308f
C17331 DVSS.n9373 VSS 0.046402f
C17332 DVSS.n9375 VSS 0.052308f
C17333 DVSS.n9376 VSS 0.393287f
C17334 DVSS.n9377 VSS 0.036911f
C17335 DVSS.n9378 VSS 0.397368f
C17336 DVSS.n9380 VSS 0.043865f
C17337 DVSS.n9381 VSS 0.397368f
C17338 DVSS.n9382 VSS 0.030953f
C17339 DVSS.n9383 VSS 0.047218f
C17340 DVSS.n9384 VSS -2.20997f
C17341 DVSS.n9385 VSS 76.3007f
C17342 DVSS.n9386 VSS 16.4147f
C17343 DVSS.n9387 VSS 6.77029f
C17344 DVSS.n9388 VSS 1.8445f
C17345 DVSS.n9389 VSS -2.20997f
C17346 DVSS.n9390 VSS 0.035198f
C17347 DVSS.n9392 VSS 0.047218f
C17348 DVSS.n9394 VSS 0.021932f
C17349 DVSS.n9395 VSS 0.397368f
C17350 DVSS.n9397 VSS 0.397368f
C17351 DVSS.n9399 VSS 0.048189f
C17352 DVSS.n9402 VSS 0.048189f
C17353 DVSS.n9404 VSS 0.393287f
C17354 DVSS.n9406 VSS 0.393287f
C17355 DVSS.n9408 VSS 0.048189f
C17356 DVSS.n9411 VSS 0.048189f
C17357 DVSS.n9413 VSS 0.173326f
C17358 DVSS.n9415 VSS 0.170217f
C17359 DVSS.n9418 VSS 0.045559f
C17360 DVSS.n9419 VSS 0.078891f
C17361 DVSS.n9420 VSS 0.029924f
C17362 DVSS.n9421 VSS 0.026154f
C17363 DVSS.n9422 VSS 0.029924f
C17364 DVSS.n9423 VSS 0.026154f
C17365 DVSS.n9424 VSS 0.041971f
C17366 DVSS.n9425 VSS 0.026154f
C17367 DVSS.n9426 VSS 0.041971f
C17368 DVSS.n9427 VSS 0.026154f
C17369 DVSS.n9428 VSS 0.041971f
C17370 DVSS.n9429 VSS 0.041971f
C17371 DVSS.n9430 VSS 0.023834f
C17372 DVSS.n9431 VSS 0.025099f
C17373 DVSS.n9432 VSS 0.041971f
C17374 DVSS.n9433 VSS 0.026154f
C17375 DVSS.n9434 VSS 0.041971f
C17376 DVSS.n9435 VSS 0.026154f
C17377 DVSS.n9436 VSS 0.041971f
C17378 DVSS.n9437 VSS 0.026154f
C17379 DVSS.n9438 VSS 0.041971f
C17380 DVSS.n9439 VSS 0.026154f
C17381 DVSS.n9440 VSS 0.041971f
C17382 DVSS.n9441 VSS 0.026154f
C17383 DVSS.n9442 VSS 0.041971f
C17384 DVSS.n9443 VSS 0.026154f
C17385 DVSS.n9444 VSS 0.041971f
C17386 DVSS.n9445 VSS 0.041971f
C17387 DVSS.n9446 VSS 0.02299f
C17388 DVSS.n9447 VSS 0.025943f
C17389 DVSS.n9448 VSS 0.041971f
C17390 DVSS.n9449 VSS 0.026154f
C17391 DVSS.n9450 VSS 0.041971f
C17392 DVSS.n9451 VSS 0.026154f
C17393 DVSS.n9452 VSS 0.041971f
C17394 DVSS.n9453 VSS 0.026154f
C17395 DVSS.n9454 VSS 0.041971f
C17396 DVSS.n9455 VSS 0.026154f
C17397 DVSS.n9456 VSS 0.041971f
C17398 DVSS.n9457 VSS 0.026154f
C17399 DVSS.n9458 VSS 0.041971f
C17400 DVSS.n9459 VSS 0.041971f
C17401 DVSS.n9460 VSS 0.025521f
C17402 DVSS.n9461 VSS 0.023412f
C17403 DVSS.n9462 VSS 0.041971f
C17404 DVSS.n9463 VSS 0.026154f
C17405 DVSS.n9464 VSS 0.041971f
C17406 DVSS.n9465 VSS 0.026154f
C17407 DVSS.n9466 VSS 0.041971f
C17408 DVSS.n9467 VSS 0.041971f
C17409 DVSS.n9468 VSS 0.026154f
C17410 DVSS.n9469 VSS 0.026154f
C17411 DVSS.n9470 VSS 0.022779f
C17412 DVSS.n9471 VSS 0.176874f
C17413 DVSS.n9472 VSS 0.022779f
C17414 DVSS.n9473 VSS 0.026154f
C17415 DVSS.n9474 VSS 0.041971f
C17416 DVSS.n9475 VSS 0.041971f
C17417 DVSS.n9476 VSS 0.031479f
C17418 DVSS.n9477 VSS 0.045559f
C17419 DVSS.n9478 VSS 0.045348f
C17420 DVSS.n9479 VSS 0.031479f
C17421 DVSS.n9480 VSS 0.041971f
C17422 DVSS.n9481 VSS 0.02299f
C17423 DVSS.n9482 VSS 0.025943f
C17424 DVSS.n9483 VSS 0.041971f
C17425 DVSS.n9484 VSS 0.026154f
C17426 DVSS.n9485 VSS 0.041971f
C17427 DVSS.n9486 VSS 0.026154f
C17428 DVSS.n9487 VSS 0.041971f
C17429 DVSS.n9488 VSS 0.026154f
C17430 DVSS.n9489 VSS 0.041971f
C17431 DVSS.n9490 VSS 0.026154f
C17432 DVSS.n9491 VSS 0.041971f
C17433 DVSS.n9492 VSS 0.026154f
C17434 DVSS.n9493 VSS 0.041971f
C17435 DVSS.n9494 VSS 0.041971f
C17436 DVSS.n9495 VSS 0.025521f
C17437 DVSS.n9496 VSS 0.023412f
C17438 DVSS.n9497 VSS 0.041971f
C17439 DVSS.n9498 VSS 0.026154f
C17440 DVSS.n9499 VSS 0.041971f
C17441 DVSS.n9500 VSS 0.026154f
C17442 DVSS.n9501 VSS 0.041971f
C17443 DVSS.n9502 VSS 0.026154f
C17444 DVSS.n9503 VSS 0.041971f
C17445 DVSS.n9504 VSS 0.026154f
C17446 DVSS.n9505 VSS 0.041971f
C17447 DVSS.n9506 VSS 0.026154f
C17448 DVSS.n9507 VSS 0.041971f
C17449 DVSS.n9508 VSS 0.026154f
C17450 DVSS.n9509 VSS 0.041971f
C17451 DVSS.n9510 VSS 0.041971f
C17452 DVSS.n9511 VSS 0.024678f
C17453 DVSS.n9512 VSS 0.024256f
C17454 DVSS.n9513 VSS 0.041971f
C17455 DVSS.n9514 VSS 0.026154f
C17456 DVSS.n9515 VSS 0.041971f
C17457 DVSS.n9516 VSS 0.026154f
C17458 DVSS.n9517 VSS 0.041971f
C17459 DVSS.n9518 VSS 0.026154f
C17460 DVSS.n9519 VSS 0.041971f
C17461 DVSS.n9520 VSS 0.026154f
C17462 DVSS.n9521 VSS 0.041971f
C17463 DVSS.n9522 VSS 0.026154f
C17464 DVSS.n9523 VSS 0.041971f
C17465 DVSS.n9524 VSS 0.026154f
C17466 DVSS.n9525 VSS 0.041971f
C17467 DVSS.n9526 VSS 0.041971f
C17468 DVSS.n9527 VSS 0.023834f
C17469 DVSS.n9528 VSS 0.025099f
C17470 DVSS.n9529 VSS 0.041971f
C17471 DVSS.n9530 VSS 0.026154f
C17472 DVSS.n9531 VSS 0.041971f
C17473 DVSS.n9532 VSS 0.029924f
C17474 DVSS.n9533 VSS 0.029924f
C17475 DVSS.n9534 VSS 0.078891f
C17476 DVSS.n9535 VSS 0.045559f
C17477 DVSS.n9537 VSS 0.170217f
C17478 DVSS.n9540 VSS 0.052308f
C17479 DVSS.n9541 VSS 0.173326f
C17480 DVSS.n9542 VSS 0.036911f
C17481 DVSS.n9543 VSS 0.036911f
C17482 DVSS.n9544 VSS 0.176874f
C17483 DVSS.n9545 VSS 0.099554f
C17484 DVSS.n9546 VSS 0.099554f
C17485 DVSS.n9548 VSS 0.287731f
C17486 DVSS.n9549 VSS 0.052308f
C17487 DVSS.n9550 VSS 0.052308f
C17488 DVSS.n9551 VSS 0.052308f
C17489 DVSS.n9552 VSS 0.052308f
C17490 DVSS.n9553 VSS 0.052308f
C17491 DVSS.n9554 VSS 0.052308f
C17492 DVSS.n9555 VSS 0.052308f
C17493 DVSS.n9556 VSS 0.052308f
C17494 DVSS.n9557 VSS 0.052308f
C17495 DVSS.n9558 VSS 0.052308f
C17496 DVSS.n9559 VSS 0.052308f
C17497 DVSS.n9560 VSS 0.052308f
C17498 DVSS.n9561 VSS 0.052308f
C17499 DVSS.n9562 VSS 0.052308f
C17500 DVSS.n9563 VSS 0.052308f
C17501 DVSS.n9564 VSS 0.052308f
C17502 DVSS.n9565 VSS 0.052308f
C17503 DVSS.n9566 VSS 0.052308f
C17504 DVSS.n9576 VSS 0.176874f
C17505 DVSS.n9578 VSS 0.052308f
C17506 DVSS.n9579 VSS 0.052308f
C17507 DVSS.n9580 VSS 0.176874f
C17508 DVSS.n9581 VSS 0.052308f
C17509 DVSS.n9583 VSS 0.176874f
C17510 DVSS.n9584 VSS 0.154453f
C17511 DVSS.n9585 VSS 0.206768f
C17512 DVSS.n9586 VSS 0.353747f
C17513 DVSS.n9587 VSS 0.353747f
C17514 DVSS.n9588 VSS 0.353747f
C17515 DVSS.n9589 VSS 0.353747f
C17516 DVSS.n9590 VSS 0.353747f
C17517 DVSS.n9591 VSS 0.353747f
C17518 DVSS.n9592 VSS 0.353747f
C17519 DVSS.n9593 VSS 0.353747f
C17520 DVSS.n9594 VSS 0.353747f
C17521 DVSS.n9595 VSS 0.353747f
C17522 DVSS.n9596 VSS 0.353747f
C17523 DVSS.n9597 VSS 0.353747f
C17524 DVSS.n9598 VSS 0.353747f
C17525 DVSS.n9599 VSS 0.353747f
C17526 DVSS.n9600 VSS 0.353747f
C17527 DVSS.n9601 VSS 0.353747f
C17528 DVSS.n9602 VSS 0.353747f
C17529 DVSS.n9603 VSS 0.353747f
C17530 DVSS.n9604 VSS 0.353747f
C17531 DVSS.n9605 VSS 0.353747f
C17532 DVSS.n9606 VSS 0.353747f
C17533 DVSS.n9607 VSS 0.353747f
C17534 DVSS.n9608 VSS 0.353747f
C17535 DVSS.n9609 VSS 0.353747f
C17536 DVSS.n9610 VSS 0.353747f
C17537 DVSS.n9611 VSS 0.353747f
C17538 DVSS.n9612 VSS 0.353747f
C17539 DVSS.n9613 VSS 0.353747f
C17540 DVSS.n9614 VSS 0.353747f
C17541 DVSS.n9615 VSS 0.353747f
C17542 DVSS.n9616 VSS 0.353747f
C17543 DVSS.n9617 VSS 0.353747f
C17544 DVSS.n9618 VSS 0.353747f
C17545 DVSS.n9619 VSS 0.313888f
C17546 DVSS.n9620 VSS 0.313888f
C17547 DVSS.n9621 VSS 0.675109f
C17548 DVSS.n9622 VSS 0.425991f
C17549 DVSS.n9623 VSS 0.313888f
C17550 DVSS.n9624 VSS 0.353747f
C17551 DVSS.n9625 VSS 0.353747f
C17552 DVSS.n9626 VSS 0.353747f
C17553 DVSS.n9627 VSS 0.353747f
C17554 DVSS.n9628 VSS 0.287731f
C17555 DVSS.n9629 VSS 0.353747f
C17556 DVSS.n9630 VSS 0.353747f
C17557 DVSS.n9631 VSS 0.353747f
C17558 DVSS.n9632 VSS 0.353747f
C17559 DVSS.n9633 VSS 0.353747f
C17560 DVSS.n9634 VSS 0.154453f
C17561 DVSS.n9636 VSS 0.052308f
C17562 DVSS.n9638 VSS 0.052308f
C17563 DVSS.n9639 VSS 0.052308f
C17564 DVSS.n9641 VSS 0.052308f
C17565 DVSS.n9642 VSS 0.052308f
C17566 DVSS.n9644 VSS 0.052308f
C17567 DVSS.n9645 VSS 0.052308f
C17568 DVSS.n9647 VSS 0.052308f
C17569 DVSS.n9649 VSS 0.052308f
C17570 DVSS.n9650 VSS 0.052308f
C17571 DVSS.n9652 VSS 0.052308f
C17572 DVSS.n9653 VSS 0.052308f
C17573 DVSS.n9655 VSS 0.052308f
C17574 DVSS.n9656 VSS 0.052308f
C17575 DVSS.n9658 VSS 0.176874f
C17576 DVSS.n9659 VSS 0.026154f
C17577 DVSS.n9660 VSS 0.176874f
C17578 DVSS.n9661 VSS 0.310152f
C17579 DVSS.n9662 VSS 0.353747f
C17580 DVSS.n9663 VSS 0.353747f
C17581 DVSS.n9664 VSS 0.353747f
C17582 DVSS.n9665 VSS 0.353747f
C17583 DVSS.n9666 VSS 0.353747f
C17584 DVSS.n9667 VSS 0.353747f
C17585 DVSS.n9668 VSS 0.353747f
C17586 DVSS.n9669 VSS 0.353747f
C17587 DVSS.n9670 VSS 0.353747f
C17588 DVSS.n9671 VSS 0.353747f
C17589 DVSS.n9672 VSS 0.353747f
C17590 DVSS.n9673 VSS 0.353747f
C17591 DVSS.n9674 VSS 0.353747f
C17592 DVSS.n9675 VSS 0.353747f
C17593 DVSS.n9676 VSS 0.353747f
C17594 DVSS.n9677 VSS 0.353747f
C17595 DVSS.n9678 VSS 0.353747f
C17596 DVSS.n9679 VSS 0.353747f
C17597 DVSS.n9680 VSS 0.353747f
C17598 DVSS.n9681 VSS 0.353747f
C17599 DVSS.n9682 VSS 0.353747f
C17600 DVSS.n9683 VSS 0.353747f
C17601 DVSS.n9684 VSS 0.353747f
C17602 DVSS.n9685 VSS 0.287731f
C17603 DVSS.n9686 VSS 0.353747f
C17604 DVSS.n9687 VSS 0.353747f
C17605 DVSS.n9688 VSS 0.353747f
C17606 DVSS.n9689 VSS 0.353747f
C17607 DVSS.n9690 VSS 0.353747f
C17608 DVSS.n9691 VSS 0.154453f
C17609 DVSS.n9693 VSS 0.052308f
C17610 DVSS.n9695 VSS 0.052308f
C17611 DVSS.n9696 VSS 0.052308f
C17612 DVSS.n9698 VSS 0.052308f
C17613 DVSS.n9699 VSS 0.052308f
C17614 DVSS.n9701 VSS 0.052308f
C17615 DVSS.n9702 VSS 0.052308f
C17616 DVSS.n9704 VSS 0.052308f
C17617 DVSS.n9706 VSS 0.052308f
C17618 DVSS.n9707 VSS 0.052308f
C17619 DVSS.n9709 VSS 0.052308f
C17620 DVSS.n9710 VSS 0.052308f
C17621 DVSS.n9712 VSS 0.052308f
C17622 DVSS.n9713 VSS 0.052308f
C17623 DVSS.n9715 VSS 0.176874f
C17624 DVSS.n9716 VSS 0.026154f
C17625 DVSS.n9717 VSS 0.176874f
C17626 DVSS.n9718 VSS 0.163172f
C17627 DVSS.n9719 VSS 0.206768f
C17628 DVSS.n9720 VSS 0.206768f
C17629 DVSS.n9721 VSS 0.425991f
C17630 DVSS.n9722 VSS 0.323853f
C17631 DVSS.n9723 VSS 0.323853f
C17632 DVSS.n9724 VSS 0.323853f
C17633 DVSS.n9725 VSS 0.353747f
C17634 DVSS.n9726 VSS 0.287731f
C17635 DVSS.n9727 VSS 0.353747f
C17636 DVSS.n9728 VSS 0.353747f
C17637 DVSS.n9729 VSS 0.353747f
C17638 DVSS.n9730 VSS 0.353747f
C17639 DVSS.n9731 VSS 0.353747f
C17640 DVSS.n9732 VSS 0.353747f
C17641 DVSS.n9733 VSS 0.154453f
C17642 DVSS.n9734 VSS 0.049144f
C17643 DVSS.n9735 VSS 0.154453f
C17644 DVSS.n9736 VSS 0.052308f
C17645 DVSS.n9738 VSS 0.052308f
C17646 DVSS.n9739 VSS 0.052308f
C17647 DVSS.n9741 VSS 0.052308f
C17648 DVSS.n9742 VSS 0.052308f
C17649 DVSS.n9744 VSS 0.052308f
C17650 DVSS.n9745 VSS 0.052308f
C17651 DVSS.n9747 VSS 0.052308f
C17652 DVSS.n9748 VSS 0.052308f
C17653 DVSS.n9750 VSS 0.052308f
C17654 DVSS.n9751 VSS 0.052308f
C17655 DVSS.n9753 VSS 0.052308f
C17656 DVSS.n9754 VSS 0.052308f
C17657 DVSS.n9756 VSS 0.052308f
C17658 DVSS.n9757 VSS 0.052308f
C17659 DVSS.n9759 VSS 0.052308f
C17660 DVSS.n9760 VSS 0.052308f
C17661 DVSS.n9762 VSS 0.052308f
C17662 DVSS.n9763 VSS 0.052308f
C17663 DVSS.n9765 VSS 0.052308f
C17664 DVSS.n9766 VSS 0.052308f
C17665 DVSS.n9768 VSS 0.176874f
C17666 DVSS.n9769 VSS 0.022779f
C17667 DVSS.n9770 VSS 0.176874f
C17668 DVSS.n9771 VSS 0.154453f
C17669 DVSS.n9772 VSS 0.353747f
C17670 DVSS.n9773 VSS 0.353747f
C17671 DVSS.n9774 VSS 0.353747f
C17672 DVSS.n9775 VSS 0.353747f
C17673 DVSS.n9776 VSS 0.353747f
C17674 DVSS.n9777 VSS 0.353747f
C17675 DVSS.n9778 VSS 0.353747f
C17676 DVSS.n9779 VSS 0.353747f
C17677 DVSS.n9780 VSS 0.318871f
C17678 DVSS.n9781 VSS 0.318871f
C17679 DVSS.n9782 VSS 0.21175f
C17680 DVSS.n9783 VSS 0.181856f
C17681 DVSS.n9784 VSS 0.348765f
C17682 DVSS.n9785 VSS 0.682774f
C17683 DVSS.n9786 VSS 1.32112f
C17684 DVSS.n9787 VSS 0.353747f
C17685 DVSS.n9788 VSS 0.154453f
C17686 DVSS.n9799 VSS 0.176874f
C17687 DVSS.n9802 VSS 0.052308f
C17688 DVSS.n9803 VSS 0.176874f
C17689 DVSS.n9804 VSS 0.099554f
C17690 DVSS.n9805 VSS 0.099554f
C17691 DVSS.n9807 VSS 0.052308f
C17692 DVSS.n9809 VSS 0.052308f
C17693 DVSS.n9811 VSS 0.052308f
C17694 DVSS.n9813 VSS 0.052308f
C17695 DVSS.n9815 VSS 0.052308f
C17696 DVSS.n9817 VSS 0.052308f
C17697 DVSS.n9819 VSS 0.052308f
C17698 DVSS.n9821 VSS 0.052308f
C17699 DVSS.n9823 VSS 0.052308f
C17700 DVSS.n9825 VSS 0.052308f
C17701 DVSS.n9827 VSS 0.052308f
C17702 DVSS.n9839 VSS 0.176874f
C17703 DVSS.n9841 VSS 0.125804f
C17704 DVSS.n9842 VSS 0.099554f
C17705 DVSS.n9843 VSS 0.176874f
C17706 DVSS.n9844 VSS 0.154453f
C17707 DVSS.n9845 VSS 0.353747f
C17708 DVSS.n9846 VSS 0.682774f
C17709 DVSS.n9847 VSS 1.32112f
C17710 DVSS.n9848 VSS 0.262819f
C17711 DVSS.n9849 VSS 0.302678f
C17712 DVSS.n9850 VSS 0.227943f
C17713 DVSS.n9851 VSS 0.353747f
C17714 DVSS.n9852 VSS 0.353747f
C17715 DVSS.n9853 VSS 0.353747f
C17716 DVSS.n9854 VSS 0.353747f
C17717 DVSS.n9855 VSS 0.353747f
C17718 DVSS.n9856 VSS 0.353747f
C17719 DVSS.n9857 VSS 0.353747f
C17720 DVSS.n9858 VSS 0.353747f
C17721 DVSS.n9859 VSS 0.353747f
C17722 DVSS.n9860 VSS 0.353747f
C17723 DVSS.n9861 VSS 0.353747f
C17724 DVSS.n9862 VSS 0.353747f
C17725 DVSS.n9863 VSS 0.353747f
C17726 DVSS.n9864 VSS 0.353747f
C17727 DVSS.n9865 VSS 0.353747f
C17728 DVSS.n9866 VSS 0.323853f
C17729 DVSS.n9867 VSS 0.323853f
C17730 DVSS.n9868 VSS 0.675109f
C17731 DVSS.n9869 VSS 0.425991f
C17732 DVSS.n9870 VSS 0.206768f
C17733 DVSS.n9871 VSS 0.206768f
C17734 DVSS.n9872 VSS 0.425991f
C17735 DVSS.n9873 VSS 0.323853f
C17736 DVSS.n9874 VSS 0.353747f
C17737 DVSS.n9875 VSS 0.353747f
C17738 DVSS.n9876 VSS 0.353747f
C17739 DVSS.n9877 VSS 0.353747f
C17740 DVSS.n9878 VSS 0.287731f
C17741 DVSS.n9879 VSS 0.353747f
C17742 DVSS.n9880 VSS 0.353747f
C17743 DVSS.n9881 VSS 0.353747f
C17744 DVSS.n9882 VSS 0.353747f
C17745 DVSS.n9883 VSS 0.353747f
C17746 DVSS.n9884 VSS 0.353747f
C17747 DVSS.n9885 VSS 0.154453f
C17748 DVSS.n9886 VSS 0.176874f
C17749 DVSS.n9887 VSS 0.022779f
C17750 DVSS.n9888 VSS 0.176874f
C17751 DVSS.n9889 VSS 0.310152f
C17752 DVSS.n9890 VSS 0.353747f
C17753 DVSS.n9891 VSS 0.353747f
C17754 DVSS.n9892 VSS 0.353747f
C17755 DVSS.n9893 VSS 0.353747f
C17756 DVSS.n9894 VSS 0.346274f
C17757 DVSS.n9895 VSS 0.346274f
C17758 DVSS.n9896 VSS 0.346274f
C17759 DVSS.n9897 VSS 0.118331f
C17760 DVSS.n9898 VSS 0.052308f
C17761 DVSS.n9899 VSS 0.052308f
C17762 DVSS.n9900 VSS 0.052308f
C17763 DVSS.n9901 VSS 0.052308f
C17764 DVSS.n9902 VSS 0.052308f
C17765 DVSS.n9903 VSS 0.052308f
C17766 DVSS.n9904 VSS 0.052308f
C17767 DVSS.n9905 VSS 0.052308f
C17768 DVSS.n9906 VSS 0.052308f
C17769 DVSS.n9907 VSS 0.052308f
C17770 DVSS.n9908 VSS 0.052308f
C17771 DVSS.n9909 VSS 0.052308f
C17772 DVSS.n9910 VSS 0.052308f
C17773 DVSS.n9911 VSS 0.052308f
C17774 DVSS.n9912 VSS 0.052308f
C17775 DVSS.n9913 VSS 0.052308f
C17776 DVSS.n9914 VSS 0.052308f
C17777 DVSS.n9915 VSS 0.052308f
C17778 DVSS.n9916 VSS 0.052308f
C17779 DVSS.n9917 VSS 0.052308f
C17780 DVSS.n9918 VSS 0.052308f
C17781 DVSS.n9929 VSS 0.176874f
C17782 DVSS.n9931 VSS 0.052308f
C17783 DVSS.n9932 VSS 0.176874f
C17784 DVSS.n9933 VSS 0.22484f
C17785 DVSS.n9934 VSS 0.779994f
C17786 DVSS.n9935 VSS 0.682774f
C17787 DVSS.n9936 VSS 0.353747f
C17788 DVSS.n9937 VSS 0.353747f
C17789 DVSS.n9938 VSS 0.353747f
C17790 DVSS.n9939 VSS 0.321362f
C17791 DVDD.n0 VSS 0.189849f
C17792 DVDD.n1 VSS 0.210614f
C17793 DVDD.n2 VSS 0.210614f
C17794 DVDD.n3 VSS 0.091958f
C17795 DVDD.n4 VSS 0.013137f
C17796 DVDD.n5 VSS 0.013137f
C17797 DVDD.n6 VSS 0.013137f
C17798 DVDD.n7 VSS 0.013137f
C17799 DVDD.n8 VSS 0.013137f
C17800 DVDD.n9 VSS 0.013137f
C17801 DVDD.n10 VSS 0.013137f
C17802 DVDD.n11 VSS 0.013137f
C17803 DVDD.n12 VSS 0.013137f
C17804 DVDD.n13 VSS 0.013137f
C17805 DVDD.n14 VSS 0.013137f
C17806 DVDD.n15 VSS 0.013878f
C17807 DVDD.n16 VSS 0.210614f
C17808 DVDD.n17 VSS 0.210614f
C17809 DVDD.n18 VSS 0.210614f
C17810 DVDD.n19 VSS 0.210614f
C17811 DVDD.n20 VSS 0.105307f
C17812 DVDD.n21 VSS 0.210614f
C17813 DVDD.n22 VSS 0.210614f
C17814 DVDD.n23 VSS 0.210614f
C17815 DVDD.n24 VSS 0.105307f
C17816 DVDD.n25 VSS 0.066735f
C17817 DVDD.n26 VSS 0.066735f
C17818 DVDD.n27 VSS 0.066735f
C17819 DVDD.n28 VSS 0.066735f
C17820 DVDD.n29 VSS 0.066735f
C17821 DVDD.n30 VSS 0.091958f
C17822 DVDD.n32 VSS 1.85245f
C17823 DVDD.n35 VSS 0.066735f
C17824 DVDD.n38 VSS 0.066735f
C17825 DVDD.n41 VSS 0.066735f
C17826 DVDD.n44 VSS 0.066735f
C17827 DVDD.n46 VSS 0.560793f
C17828 DVDD.n47 VSS 0.210614f
C17829 DVDD.n48 VSS 0.210614f
C17830 DVDD.n49 VSS 0.210614f
C17831 DVDD.n50 VSS 0.210614f
C17832 DVDD.n51 VSS 0.210614f
C17833 DVDD.n52 VSS 0.210614f
C17834 DVDD.n53 VSS 0.210614f
C17835 DVDD.n54 VSS 0.210614f
C17836 DVDD.n55 VSS 0.105307f
C17837 DVDD.n56 VSS 0.210614f
C17838 DVDD.n57 VSS 0.210614f
C17839 DVDD.n58 VSS 0.210614f
C17840 DVDD.n59 VSS 0.105307f
C17841 DVDD.n60 VSS 0.029062f
C17842 DVDD.n61 VSS 0.029062f
C17843 DVDD.n62 VSS 0.029062f
C17844 DVDD.n63 VSS 0.029062f
C17845 DVDD.n64 VSS 0.029062f
C17846 DVDD.n65 VSS 0.091958f
C17847 DVDD.n66 VSS 0.029062f
C17848 DVDD.n67 VSS 0.029062f
C17849 DVDD.n68 VSS 0.029062f
C17850 DVDD.n69 VSS 0.029062f
C17851 DVDD.n70 VSS 0.029062f
C17852 DVDD.n71 VSS 0.033368f
C17853 DVDD.n72 VSS 0.091958f
C17854 DVDD.n73 VSS 0.105307f
C17855 DVDD.n74 VSS 0.058124f
C17856 DVDD.n75 VSS 0.114418f
C17857 DVDD.n76 VSS 0.114418f
C17858 DVDD.n77 VSS 0.058124f
C17859 DVDD.n78 VSS 0.15585f
C17860 DVDD.n79 VSS 0.05355f
C17861 DVDD.n80 VSS 0.114418f
C17862 DVDD.n81 VSS 0.029062f
C17863 DVDD.n82 VSS 0.029331f
C17864 DVDD.n83 VSS 0.027333f
C17865 DVDD.n84 VSS 0.197054f
C17866 DVDD.n85 VSS 0.217712f
C17867 DVDD.n86 VSS 0.013137f
C17868 DVDD.n87 VSS 0.066735f
C17869 DVDD.n88 VSS 0.197054f
C17870 DVDD.n89 VSS 0.197054f
C17871 DVDD.n90 VSS 0.013137f
C17872 DVDD.n91 VSS 0.033368f
C17873 DVDD.n92 VSS 0.033368f
C17874 DVDD.n93 VSS 0.026274f
C17875 DVDD.n94 VSS 0.030088f
C17876 DVDD.n95 VSS 0.060175f
C17877 DVDD.n96 VSS 0.059611f
C17878 DVDD.n97 VSS 0.026274f
C17879 DVDD.n98 VSS 0.060175f
C17880 DVDD.n99 VSS 0.057655f
C17881 DVDD.n100 VSS 0.170687f
C17882 DVDD.n101 VSS 0.060175f
C17883 DVDD.n102 VSS 0.045979f
C17884 DVDD.n103 VSS 1.62757f
C17885 DVDD.n104 VSS 0.557869f
C17886 DVDD.n105 VSS 0.556703f
C17887 DVDD.n106 VSS 0.197054f
C17888 DVDD.n107 VSS 0.033368f
C17889 DVDD.n108 VSS 0.197054f
C17890 DVDD.n109 VSS 0.026274f
C17891 DVDD.n110 VSS 0.026274f
C17892 DVDD.n111 VSS 0.272585f
C17893 DVDD.n112 VSS 0.029062f
C17894 DVDD.n113 VSS 0.066735f
C17895 DVDD.n114 VSS 0.029062f
C17896 DVDD.n115 VSS 0.013137f
C17897 DVDD.n116 VSS 0.197054f
C17898 DVDD.n117 VSS 0.197054f
C17899 DVDD.n118 VSS 0.026274f
C17900 DVDD.n119 VSS 0.611141f
C17901 DVDD.n120 VSS 0.197054f
C17902 DVDD.n121 VSS 0.197054f
C17903 DVDD.n122 VSS 0.271282f
C17904 DVDD.n123 VSS 0.197054f
C17905 DVDD.n124 VSS 0.197054f
C17906 DVDD.n125 VSS 0.029062f
C17907 DVDD.n126 VSS 0.029062f
C17908 DVDD.n127 VSS 0.066735f
C17909 DVDD.n128 VSS 0.066735f
C17910 DVDD.n129 VSS 0.197054f
C17911 DVDD.n130 VSS 0.033368f
C17912 DVDD.n131 VSS 0.033368f
C17913 DVDD.n132 VSS 0.030088f
C17914 DVDD.n133 VSS 0.029062f
C17915 DVDD.n134 VSS 0.114418f
C17916 DVDD.n135 VSS 0.114418f
C17917 DVDD.n136 VSS 0.033368f
C17918 DVDD.n137 VSS 0.225658f
C17919 DVDD.n138 VSS 0.026274f
C17920 DVDD.n139 VSS 0.02691f
C17921 DVDD.n140 VSS 0.060175f
C17922 DVDD.n141 VSS 0.173939f
C17923 DVDD.n142 VSS 0.033368f
C17924 DVDD.n143 VSS 0.048706f
C17925 DVDD.n144 VSS 0.029062f
C17926 DVDD.n145 VSS 0.201821f
C17927 DVDD.n146 VSS 0.548254f
C17928 DVDD.n147 VSS 0.033368f
C17929 DVDD.n148 VSS 0.066735f
C17930 DVDD.n149 VSS 0.066735f
C17931 DVDD.n150 VSS 0.066735f
C17932 DVDD.n151 VSS 0.548254f
C17933 DVDD.n152 VSS 0.201821f
C17934 DVDD.n153 VSS 0.033368f
C17935 DVDD.n154 VSS 0.048168f
C17936 DVDD.n155 VSS 0.060739f
C17937 DVDD.n156 VSS 0.029062f
C17938 DVDD.n157 VSS 0.114418f
C17939 DVDD.n158 VSS 0.114418f
C17940 DVDD.n159 VSS 0.114418f
C17941 DVDD.n160 VSS 0.058124f
C17942 DVDD.n161 VSS 0.114418f
C17943 DVDD.n162 VSS 0.114418f
C17944 DVDD.n163 VSS 0.114418f
C17945 DVDD.n164 VSS 0.030088f
C17946 DVDD.n165 VSS 0.030408f
C17947 DVDD.n166 VSS 0.197054f
C17948 DVDD.n167 VSS 0.197054f
C17949 DVDD.n168 VSS 0.033368f
C17950 DVDD.n169 VSS 0.066735f
C17951 DVDD.n170 VSS 0.197054f
C17952 DVDD.n171 VSS 0.033368f
C17953 DVDD.n172 VSS 0.032022f
C17954 DVDD.n173 VSS 0.033368f
C17955 DVDD.n174 VSS 0.026274f
C17956 DVDD.n175 VSS 0.030088f
C17957 DVDD.n176 VSS 0.060175f
C17958 DVDD.n177 VSS 0.044284f
C17959 DVDD.n178 VSS 0.02691f
C17960 DVDD.n179 VSS 0.026274f
C17961 DVDD.n180 VSS 0.060175f
C17962 DVDD.n181 VSS 0.061117f
C17963 DVDD.n182 VSS 0.173937f
C17964 DVDD.n183 VSS 0.556686f
C17965 DVDD.n184 VSS 0.554173f
C17966 DVDD.n185 VSS 0.344844f
C17967 DVDD.n186 VSS 0.332131f
C17968 DVDD.n187 VSS 0.27259f
C17969 DVDD.n188 VSS 0.271712f
C17970 DVDD.n189 VSS 0.045979f
C17971 DVDD.n190 VSS 0.332131f
C17972 DVDD.n191 VSS 0.344844f
C17973 DVDD.n192 VSS 0.611119f
C17974 DVDD.n193 VSS 0.06502f
C17975 DVDD.n194 VSS 0.044284f
C17976 DVDD.n195 VSS 0.344844f
C17977 DVDD.n196 VSS 0.332131f
C17978 DVDD.n197 VSS 0.045979f
C17979 DVDD.n198 VSS 0.332131f
C17980 DVDD.n199 VSS 0.451316f
C17981 DVDD.n200 VSS 1.65039f
C17982 DVDD.n201 VSS 0.197054f
C17983 DVDD.n202 VSS 0.197054f
C17984 DVDD.n203 VSS 0.197054f
C17985 DVDD.n204 VSS 0.451316f
C17986 DVDD.n205 VSS 0.724649f
C17987 DVDD.n206 VSS 0.535541f
C17988 DVDD.n207 VSS 0.535541f
C17989 DVDD.n208 VSS 0.197054f
C17990 DVDD.n209 VSS 0.451316f
C17991 DVDD.n210 VSS 0.344844f
C17992 DVDD.n211 VSS 0.197054f
C17993 DVDD.n212 VSS 0.197054f
C17994 DVDD.n213 VSS 0.611119f
C17995 DVDD.n214 VSS 0.045979f
C17996 DVDD.n215 VSS 0.332131f
C17997 DVDD.n216 VSS 0.344844f
C17998 DVDD.n217 VSS 0.044284f
C17999 DVDD.n218 VSS 0.332131f
C18000 DVDD.n219 VSS 0.344844f
C18001 DVDD.n220 VSS 0.271708f
C18002 DVDD.n221 VSS 0.344844f
C18003 DVDD.n222 VSS 0.332131f
C18004 DVDD.n223 VSS 0.272585f
C18005 DVDD.n224 VSS 0.044284f
C18006 DVDD.n225 VSS 0.045979f
C18007 DVDD.n226 VSS 0.332131f
C18008 DVDD.n227 VSS 0.557869f
C18009 DVDD.n228 VSS 3.32205f
C18010 DVDD.n229 VSS 0.565854f
C18011 DVDD.n230 VSS 0.045979f
C18012 DVDD.n231 VSS 0.332131f
C18013 DVDD.n232 VSS 0.344844f
C18014 DVDD.n233 VSS 0.044284f
C18015 DVDD.n234 VSS 0.332131f
C18016 DVDD.n235 VSS 0.344844f
C18017 DVDD.n236 VSS 0.045979f
C18018 DVDD.n237 VSS 0.332131f
C18019 DVDD.n238 VSS 0.044284f
C18020 DVDD.n239 VSS 0.344844f
C18021 DVDD.n240 VSS 1.30659f
C18022 DVDD.n241 VSS 0.451316f
C18023 DVDD.n242 VSS 0.197054f
C18024 DVDD.n243 VSS 0.225658f
C18025 DVDD.n244 VSS 0.197054f
C18026 DVDD.n245 VSS 0.033368f
C18027 DVDD.n246 VSS 0.032022f
C18028 DVDD.n247 VSS 0.114418f
C18029 DVDD.n248 VSS 0.114418f
C18030 DVDD.n249 VSS 0.029062f
C18031 DVDD.n250 VSS 0.033368f
C18032 DVDD.n251 VSS 0.225658f
C18033 DVDD.n252 VSS 0.197054f
C18034 DVDD.n253 VSS 0.451316f
C18035 DVDD.n254 VSS 0.455731f
C18036 DVDD.n255 VSS 0.058124f
C18037 DVDD.n256 VSS 0.114418f
C18038 DVDD.n257 VSS 0.058124f
C18039 DVDD.n258 VSS 0.114418f
C18040 DVDD.n259 VSS 0.058124f
C18041 DVDD.n260 VSS 0.114418f
C18042 DVDD.n261 VSS 0.058124f
C18043 DVDD.n262 VSS 0.114418f
C18044 DVDD.n263 VSS 0.058124f
C18045 DVDD.n264 VSS 0.114418f
C18046 DVDD.n265 VSS 0.277706f
C18047 DVDD.n266 VSS 0.114418f
C18048 DVDD.n267 VSS 0.066735f
C18049 DVDD.n268 VSS 0.225658f
C18050 DVDD.n269 VSS 0.451316f
C18051 DVDD.n270 VSS 0.724649f
C18052 DVDD.n271 VSS 0.724649f
C18053 DVDD.n272 VSS 0.225658f
C18054 DVDD.n273 VSS 0.197054f
C18055 DVDD.n274 VSS 0.217712f
C18056 DVDD.n275 VSS 0.033099f
C18057 DVDD.n276 VSS 0.197054f
C18058 DVDD.n277 VSS 0.535541f
C18059 DVDD.n278 VSS 0.451316f
C18060 DVDD.n279 VSS 0.451316f
C18061 DVDD.n280 VSS 0.451316f
C18062 DVDD.n281 VSS 0.225658f
C18063 DVDD.n282 VSS 0.204999f
C18064 DVDD.n283 VSS 0.033368f
C18065 DVDD.n284 VSS 0.029062f
C18066 DVDD.n285 VSS 0.114418f
C18067 DVDD.n286 VSS 0.114418f
C18068 DVDD.n287 VSS 0.277706f
C18069 DVDD.n288 VSS 0.033368f
C18070 DVDD.n289 VSS 0.429855f
C18071 DVDD.n290 VSS 0.204999f
C18072 DVDD.n291 VSS 1.28214f
C18073 DVDD.n292 VSS 0.451316f
C18074 DVDD.n293 VSS 0.217712f
C18075 DVDD.n294 VSS 0.197054f
C18076 DVDD.n295 VSS 0.033368f
C18077 DVDD.n296 VSS 0.225658f
C18078 DVDD.n297 VSS 0.029062f
C18079 DVDD.n298 VSS 0.114418f
C18080 DVDD.n299 VSS 0.114418f
C18081 DVDD.n300 VSS 0.029062f
C18082 DVDD.n301 VSS 0.029331f
C18083 DVDD.n302 VSS 0.029062f
C18084 DVDD.n303 VSS 0.033099f
C18085 DVDD.n304 VSS 0.114418f
C18086 DVDD.n305 VSS 0.114418f
C18087 DVDD.n306 VSS 0.114418f
C18088 DVDD.n307 VSS 0.033368f
C18089 DVDD.n308 VSS 0.225658f
C18090 DVDD.n309 VSS 0.332131f
C18091 DVDD.n310 VSS 0.451316f
C18092 DVDD.n311 VSS 0.451316f
C18093 DVDD.n312 VSS 0.451316f
C18094 DVDD.n313 VSS 0.197054f
C18095 DVDD.n314 VSS 0.029869f
C18096 DVDD.n315 VSS 0.029062f
C18097 DVDD.n316 VSS 0.029062f
C18098 DVDD.n317 VSS 0.032561f
C18099 DVDD.n318 VSS 0.114418f
C18100 DVDD.n319 VSS 0.114418f
C18101 DVDD.n320 VSS 0.114418f
C18102 DVDD.n321 VSS 0.048706f
C18103 DVDD.n322 VSS 0.201821f
C18104 DVDD.n323 VSS 0.548254f
C18105 DVDD.n324 VSS 0.451316f
C18106 DVDD.n325 VSS 0.750075f
C18107 DVDD.n326 VSS 0.750075f
C18108 DVDD.n327 VSS 0.451316f
C18109 DVDD.n328 VSS 0.451316f
C18110 DVDD.n329 VSS 0.201821f
C18111 DVDD.n330 VSS 0.197054f
C18112 DVDD.n331 VSS 0.033368f
C18113 DVDD.n332 VSS 0.032022f
C18114 DVDD.n333 VSS 0.114418f
C18115 DVDD.n334 VSS 0.114418f
C18116 DVDD.n335 VSS 0.058124f
C18117 DVDD.n336 VSS 0.048168f
C18118 DVDD.n337 VSS 0.220891f
C18119 DVDD.n338 VSS 0.029062f
C18120 DVDD.n339 VSS 0.029062f
C18121 DVDD.n340 VSS 0.033368f
C18122 DVDD.n341 VSS 0.114418f
C18123 DVDD.n342 VSS 0.114418f
C18124 DVDD.n343 VSS 0.114418f
C18125 DVDD.n344 VSS 0.029062f
C18126 DVDD.n345 VSS 0.033368f
C18127 DVDD.n346 VSS 0.225658f
C18128 DVDD.n347 VSS 0.197054f
C18129 DVDD.n348 VSS 0.026274f
C18130 DVDD.n349 VSS 0.197054f
C18131 DVDD.n350 VSS 0.013137f
C18132 DVDD.n351 VSS 0.066735f
C18133 DVDD.n352 VSS 0.197054f
C18134 DVDD.n353 VSS 0.46696f
C18135 DVDD.n354 VSS 0.06502f
C18136 DVDD.n355 VSS 0.06502f
C18137 DVDD.n356 VSS 0.029062f
C18138 DVDD.n357 VSS 0.026274f
C18139 DVDD.n358 VSS 0.197054f
C18140 DVDD.n359 VSS 0.066735f
C18141 DVDD.n360 VSS 0.344844f
C18142 DVDD.n361 VSS 0.197054f
C18143 DVDD.n362 VSS 0.197054f
C18144 DVDD.n363 VSS 0.225658f
C18145 DVDD.n364 VSS 0.029062f
C18146 DVDD.n365 VSS 0.029062f
C18147 DVDD.n366 VSS 0.033368f
C18148 DVDD.n367 VSS 0.114418f
C18149 DVDD.n368 VSS 0.114418f
C18150 DVDD.n369 VSS 0.033368f
C18151 DVDD.n370 VSS 0.029062f
C18152 DVDD.n371 VSS 0.197054f
C18153 DVDD.n372 VSS 0.029062f
C18154 DVDD.n373 VSS 0.197054f
C18155 DVDD.n374 VSS 0.026274f
C18156 DVDD.n375 VSS 0.029062f
C18157 DVDD.n376 VSS 0.026274f
C18158 DVDD.n377 VSS 0.033368f
C18159 DVDD.n378 VSS 0.033368f
C18160 DVDD.n379 VSS 0.131369f
C18161 DVDD.n380 VSS 0.131369f
C18162 DVDD.n381 VSS 0.033368f
C18163 DVDD.n382 VSS 0.029062f
C18164 DVDD.n383 VSS 0.066735f
C18165 DVDD.n384 VSS 0.066735f
C18166 DVDD.n385 VSS 0.204999f
C18167 DVDD.n386 VSS 0.033368f
C18168 DVDD.n387 VSS 0.033368f
C18169 DVDD.n388 VSS 0.029028f
C18170 DVDD.n389 VSS 0.029062f
C18171 DVDD.n390 VSS 0.114418f
C18172 DVDD.n391 VSS 0.15585f
C18173 DVDD.n392 VSS 0.130242f
C18174 DVDD.n393 VSS 0.197054f
C18175 DVDD.n394 VSS 0.225658f
C18176 DVDD.n395 VSS 0.027333f
C18177 DVDD.n396 VSS 0.026274f
C18178 DVDD.n397 VSS 0.060175f
C18179 DVDD.n398 VSS 0.060175f
C18180 DVDD.n399 VSS 0.045979f
C18181 DVDD.n400 VSS 0.060175f
C18182 DVDD.n401 VSS 0.033368f
C18183 DVDD.n402 VSS 0.114418f
C18184 DVDD.n403 VSS 0.114418f
C18185 DVDD.n404 VSS 0.131369f
C18186 DVDD.n405 VSS 0.131369f
C18187 DVDD.n406 VSS 0.033368f
C18188 DVDD.n407 VSS 0.131369f
C18189 DVDD.n408 VSS 0.033368f
C18190 DVDD.n409 VSS 0.197054f
C18191 DVDD.n410 VSS 0.033368f
C18192 DVDD.n411 VSS 0.033368f
C18193 DVDD.n412 VSS 0.030088f
C18194 DVDD.n413 VSS 0.060175f
C18195 DVDD.n414 VSS 0.045979f
C18196 DVDD.n415 VSS 0.170687f
C18197 DVDD.n416 VSS 0.451316f
C18198 DVDD.n417 VSS 0.344844f
C18199 DVDD.n418 VSS 0.344844f
C18200 DVDD.n419 VSS 0.332131f
C18201 DVDD.n420 VSS 0.344844f
C18202 DVDD.n421 VSS 0.044284f
C18203 DVDD.n422 VSS 0.565854f
C18204 DVDD.n423 VSS 0.332131f
C18205 DVDD.n424 VSS 0.344844f
C18206 DVDD.n425 VSS 0.332131f
C18207 DVDD.n426 VSS 0.451316f
C18208 DVDD.n427 VSS 0.451316f
C18209 DVDD.n428 VSS 0.197054f
C18210 DVDD.n429 VSS 0.033368f
C18211 DVDD.n430 VSS 0.197054f
C18212 DVDD.n431 VSS 0.029062f
C18213 DVDD.n432 VSS 0.560793f
C18214 DVDD.n433 VSS 0.066735f
C18215 DVDD.n434 VSS 0.217712f
C18216 DVDD.n435 VSS 0.033368f
C18217 DVDD.n436 VSS 0.033368f
C18218 DVDD.n437 VSS 0.029331f
C18219 DVDD.n438 VSS 0.059611f
C18220 DVDD.n439 VSS 0.057655f
C18221 DVDD.n440 VSS 0.060175f
C18222 DVDD.n441 VSS 0.026274f
C18223 DVDD.n442 VSS 0.026274f
C18224 DVDD.n443 VSS 0.033099f
C18225 DVDD.n444 VSS 0.029062f
C18226 DVDD.n445 VSS 0.15585f
C18227 DVDD.n446 VSS 0.058124f
C18228 DVDD.n447 VSS 0.114418f
C18229 DVDD.n448 VSS 0.124509f
C18230 DVDD.n449 VSS 0.124509f
C18231 DVDD.n450 VSS 0.114418f
C18232 DVDD.n451 VSS 0.277706f
C18233 DVDD.n452 VSS 0.058124f
C18234 DVDD.n453 VSS 0.114418f
C18235 DVDD.n454 VSS 0.058124f
C18236 DVDD.n455 VSS 0.114418f
C18237 DVDD.n456 VSS 0.105307f
C18238 DVDD.n457 VSS 0.105307f
C18239 DVDD.n458 VSS 0.033368f
C18240 DVDD.n459 VSS 0.105307f
C18241 DVDD.n460 VSS 0.187625f
C18242 DVDD.n461 VSS 0.029062f
C18243 DVDD.n462 VSS 0.029062f
C18244 DVDD.n463 VSS 0.029062f
C18245 DVDD.n464 VSS 0.029062f
C18246 DVDD.n465 VSS 0.210614f
C18247 DVDD.n466 VSS 0.091958f
C18248 DVDD.n467 VSS 0.210614f
C18249 DVDD.n468 VSS 0.210614f
C18250 DVDD.n469 VSS 0.210614f
C18251 DVDD.n470 VSS 0.210614f
C18252 DVDD.n471 VSS 0.210614f
C18253 DVDD.n472 VSS 0.210614f
C18254 DVDD.n473 VSS 0.210614f
C18255 DVDD.n474 VSS 0.210614f
C18256 DVDD.n475 VSS 0.210614f
C18257 DVDD.n476 VSS 0.210614f
C18258 DVDD.n477 VSS 0.210614f
C18259 DVDD.n478 VSS 0.210614f
C18260 DVDD.n479 VSS 0.210614f
C18261 DVDD.n480 VSS 0.210614f
C18262 DVDD.n481 VSS 0.210614f
C18263 DVDD.n482 VSS 0.210614f
C18264 DVDD.n483 VSS 0.210614f
C18265 DVDD.n484 VSS 0.029062f
C18266 DVDD.n485 VSS 0.029062f
C18267 DVDD.n486 VSS 0.029062f
C18268 DVDD.n487 VSS 0.029062f
C18269 DVDD.n488 VSS 0.029062f
C18270 DVDD.n489 VSS 0.091958f
C18271 DVDD.n490 VSS 0.029062f
C18272 DVDD.n491 VSS 0.029062f
C18273 DVDD.n492 VSS 0.029062f
C18274 DVDD.n493 VSS 0.029062f
C18275 DVDD.n494 VSS 0.029062f
C18276 DVDD.n495 VSS 0.033368f
C18277 DVDD.n496 VSS 0.105307f
C18278 DVDD.n497 VSS 0.050859f
C18279 DVDD.n498 VSS 0.105307f
C18280 DVDD.n499 VSS 0.091958f
C18281 DVDD.n500 VSS 0.210614f
C18282 DVDD.n501 VSS 0.210614f
C18283 DVDD.n502 VSS 0.210614f
C18284 DVDD.n503 VSS 0.091958f
C18285 DVDD.n504 VSS 0.210614f
C18286 DVDD.n505 VSS 0.210614f
C18287 DVDD.n506 VSS 0.210614f
C18288 DVDD.n507 VSS 0.210614f
C18289 DVDD.n508 VSS 0.210614f
C18290 DVDD.n509 VSS 0.210614f
C18291 DVDD.n510 VSS 0.210614f
C18292 DVDD.n511 VSS 0.210614f
C18293 DVDD.n512 VSS 0.210614f
C18294 DVDD.n513 VSS 0.210614f
C18295 DVDD.n514 VSS 0.210614f
C18296 DVDD.n515 VSS 0.210614f
C18297 DVDD.n516 VSS 0.210614f
C18298 DVDD.n517 VSS 0.210614f
C18299 DVDD.n518 VSS 0.210614f
C18300 DVDD.n519 VSS 0.210614f
C18301 DVDD.n520 VSS 0.210614f
C18302 DVDD.n521 VSS 0.029062f
C18303 DVDD.n522 VSS 0.029062f
C18304 DVDD.n523 VSS 0.029062f
C18305 DVDD.n524 VSS 0.029062f
C18306 DVDD.n525 VSS 0.029062f
C18307 DVDD.n526 VSS 0.091958f
C18308 DVDD.n527 VSS 0.029062f
C18309 DVDD.n528 VSS 0.029062f
C18310 DVDD.n529 VSS 0.029062f
C18311 DVDD.n530 VSS 0.029062f
C18312 DVDD.n531 VSS 0.029062f
C18313 DVDD.n532 VSS 0.033368f
C18314 DVDD.n533 VSS 0.105307f
C18315 DVDD.n534 VSS 0.105307f
C18316 DVDD.n535 VSS 0.032022f
C18317 DVDD.n536 VSS 0.114418f
C18318 DVDD.n537 VSS 0.114418f
C18319 DVDD.n538 VSS 0.058124f
C18320 DVDD.n539 VSS 0.114418f
C18321 DVDD.n540 VSS 0.277706f
C18322 DVDD.n541 VSS 0.114418f
C18323 DVDD.n542 VSS 0.058124f
C18324 DVDD.n543 VSS 0.114418f
C18325 DVDD.n544 VSS 0.114418f
C18326 DVDD.n545 VSS 0.058124f
C18327 DVDD.n546 VSS 0.114418f
C18328 DVDD.n547 VSS 0.38847f
C18329 DVDD.n548 VSS 0.105307f
C18330 DVDD.n549 VSS 0.105307f
C18331 DVDD.n550 VSS 0.033368f
C18332 DVDD.n551 VSS 0.105307f
C18333 DVDD.n552 VSS 0.171309f
C18334 DVDD.n553 VSS 0.029062f
C18335 DVDD.n554 VSS 0.029062f
C18336 DVDD.n555 VSS 0.029062f
C18337 DVDD.n556 VSS 0.029062f
C18338 DVDD.n557 VSS 0.029062f
C18339 DVDD.n558 VSS 0.210614f
C18340 DVDD.n559 VSS 0.091958f
C18341 DVDD.n560 VSS 0.210614f
C18342 DVDD.n561 VSS 0.210614f
C18343 DVDD.n562 VSS 0.210614f
C18344 DVDD.n563 VSS 0.210614f
C18345 DVDD.n564 VSS 0.210614f
C18346 DVDD.n565 VSS 0.210614f
C18347 DVDD.n566 VSS 0.210614f
C18348 DVDD.n567 VSS 0.210614f
C18349 DVDD.n568 VSS 0.210614f
C18350 DVDD.n569 VSS 0.210614f
C18351 DVDD.n570 VSS 0.210614f
C18352 DVDD.n571 VSS 0.210614f
C18353 DVDD.n572 VSS 0.210614f
C18354 DVDD.n573 VSS 0.210614f
C18355 DVDD.n574 VSS 0.210614f
C18356 DVDD.n575 VSS 0.210614f
C18357 DVDD.n576 VSS 0.210614f
C18358 DVDD.n577 VSS 0.029062f
C18359 DVDD.n578 VSS 0.029062f
C18360 DVDD.n579 VSS 0.754582f
C18361 DVDD.n580 VSS 0.029062f
C18362 DVDD.n581 VSS 0.029062f
C18363 DVDD.n582 VSS 0.091958f
C18364 DVDD.n583 VSS 0.029062f
C18365 DVDD.n584 VSS 0.029062f
C18366 DVDD.n585 VSS 0.029062f
C18367 DVDD.n586 VSS 0.029062f
C18368 DVDD.n587 VSS 0.029062f
C18369 DVDD.n588 VSS 0.033368f
C18370 DVDD.n589 VSS 0.105307f
C18371 DVDD.n590 VSS 0.049783f
C18372 DVDD.n591 VSS 0.105307f
C18373 DVDD.n592 VSS 0.091958f
C18374 DVDD.n593 VSS 0.210614f
C18375 DVDD.n594 VSS 0.210614f
C18376 DVDD.n595 VSS 0.210614f
C18377 DVDD.n596 VSS 0.091958f
C18378 DVDD.n597 VSS 0.210614f
C18379 DVDD.n598 VSS 0.210614f
C18380 DVDD.n599 VSS 0.210614f
C18381 DVDD.n600 VSS 0.210614f
C18382 DVDD.n601 VSS 0.210614f
C18383 DVDD.n602 VSS 0.210614f
C18384 DVDD.n603 VSS 0.210614f
C18385 DVDD.n604 VSS 0.210614f
C18386 DVDD.n605 VSS 0.210614f
C18387 DVDD.n606 VSS 0.105307f
C18388 DVDD.n607 VSS 0.210614f
C18389 DVDD.n608 VSS 0.210614f
C18390 DVDD.n609 VSS 0.210614f
C18391 DVDD.n610 VSS 0.091958f
C18392 DVDD.n611 VSS 0.105307f
C18393 DVDD.n612 VSS 0.066735f
C18394 DVDD.n613 VSS 0.066735f
C18395 DVDD.n614 VSS 0.066735f
C18396 DVDD.n615 VSS 0.066735f
C18397 DVDD.n616 VSS 0.066735f
C18398 DVDD.n617 VSS 0.091958f
C18399 DVDD.n619 VSS 0.871867f
C18400 DVDD.n621 VSS 0.066735f
C18401 DVDD.n623 VSS 0.066735f
C18402 DVDD.n625 VSS 0.066735f
C18403 DVDD.n627 VSS 0.066735f
C18404 DVDD.n633 VSS 0.210614f
C18405 DVDD.n634 VSS 0.210614f
C18406 DVDD.n635 VSS 0.210614f
C18407 DVDD.n636 VSS 0.210614f
C18408 DVDD.n637 VSS 0.105307f
C18409 DVDD.n638 VSS 0.210614f
C18410 DVDD.n639 VSS 0.210614f
C18411 DVDD.n640 VSS 0.189849f
C18412 DVDD.n641 VSS 0.091958f
C18413 DVDD.n642 VSS 0.105307f
C18414 DVDD.n643 VSS 0.029427f
C18415 DVDD.n644 VSS 0.029427f
C18416 DVDD.n645 VSS 0.029427f
C18417 DVDD.n646 VSS 0.029427f
C18418 DVDD.n647 VSS 0.029427f
C18419 DVDD.n648 VSS 0.091958f
C18420 DVDD.n649 VSS 0.256857f
C18421 DVDD.n650 VSS 0.029427f
C18422 DVDD.n651 VSS 0.029427f
C18423 DVDD.n652 VSS 0.029427f
C18424 DVDD.n653 VSS 0.029427f
C18425 DVDD.n654 VSS 0.029427f
C18426 DVDD.n655 VSS 0.042564f
C18427 DVDD.n656 VSS 0.131369f
C18428 DVDD.n657 VSS 0.131369f
C18429 DVDD.n658 VSS 0.042564f
C18430 DVDD.n659 VSS 0.124509f
C18431 DVDD.n660 VSS 0.026274f
C18432 DVDD.n661 VSS 0.131369f
C18433 DVDD.n662 VSS 0.026274f
C18434 DVDD.n663 VSS 0.131369f
C18435 DVDD.n664 VSS 0.026274f
C18436 DVDD.n665 VSS 0.131369f
C18437 DVDD.n666 VSS 0.026274f
C18438 DVDD.n667 VSS 0.131369f
C18439 DVDD.n668 VSS 0.026274f
C18440 DVDD.n669 VSS 0.131369f
C18441 DVDD.n670 VSS 0.026274f
C18442 DVDD.n671 VSS 0.131369f
C18443 DVDD.n672 VSS 0.102976f
C18444 DVDD.n673 VSS 0.114418f
C18445 DVDD.n674 VSS 0.058124f
C18446 DVDD.n675 VSS 0.114418f
C18447 DVDD.n676 VSS 0.058124f
C18448 DVDD.n677 VSS 0.114418f
C18449 DVDD.n678 VSS 0.058124f
C18450 DVDD.n679 VSS 0.114418f
C18451 DVDD.n680 VSS 0.058124f
C18452 DVDD.n681 VSS 0.114418f
C18453 DVDD.n682 VSS 0.058124f
C18454 DVDD.n683 VSS 0.114418f
C18455 DVDD.n684 VSS 0.058124f
C18456 DVDD.n685 VSS 0.114418f
C18457 DVDD.n686 VSS 0.058124f
C18458 DVDD.n687 VSS 0.058124f
C18459 DVDD.n688 VSS 0.114418f
C18460 DVDD.n689 VSS 0.114418f
C18461 DVDD.n690 VSS 0.058124f
C18462 DVDD.n691 VSS 0.114418f
C18463 DVDD.n692 VSS 0.058124f
C18464 DVDD.n693 VSS 0.058124f
C18465 DVDD.n694 VSS 0.114418f
C18466 DVDD.n695 VSS 0.114418f
C18467 DVDD.n696 VSS 0.114418f
C18468 DVDD.n697 VSS 0.058124f
C18469 DVDD.n698 VSS 0.058124f
C18470 DVDD.n699 VSS 0.058124f
C18471 DVDD.n700 VSS 0.114418f
C18472 DVDD.n701 VSS 0.114418f
C18473 DVDD.n702 VSS 0.114418f
C18474 DVDD.n703 VSS 0.114418f
C18475 DVDD.n704 VSS 0.033099f
C18476 DVDD.n705 VSS 0.029331f
C18477 DVDD.n706 VSS 0.114418f
C18478 DVDD.n707 VSS 0.033368f
C18479 DVDD.n708 VSS 0.114418f
C18480 DVDD.n709 VSS 0.033368f
C18481 DVDD.n710 VSS 0.114418f
C18482 DVDD.n711 VSS 0.033368f
C18483 DVDD.n712 VSS 0.114418f
C18484 DVDD.n713 VSS 0.033368f
C18485 DVDD.n714 VSS 0.114418f
C18486 DVDD.n715 VSS 0.033368f
C18487 DVDD.n716 VSS 0.114418f
C18488 DVDD.n717 VSS 0.033368f
C18489 DVDD.n718 VSS 0.114418f
C18490 DVDD.n719 VSS 0.114418f
C18491 DVDD.n720 VSS 0.032022f
C18492 DVDD.n721 VSS 0.030408f
C18493 DVDD.n722 VSS 0.114418f
C18494 DVDD.n723 VSS 0.033368f
C18495 DVDD.n724 VSS 0.38847f
C18496 DVDD.n725 VSS 0.747408f
C18497 DVDD.n726 VSS 0.029427f
C18498 DVDD.n727 VSS 0.131369f
C18499 DVDD.n728 VSS 0.029427f
C18500 DVDD.n729 VSS 0.131369f
C18501 DVDD.n730 VSS 0.029427f
C18502 DVDD.n731 VSS 0.131369f
C18503 DVDD.n732 VSS 0.029427f
C18504 DVDD.n733 VSS 0.131369f
C18505 DVDD.n734 VSS 0.029427f
C18506 DVDD.n735 VSS 0.131369f
C18507 DVDD.n736 VSS 0.029427f
C18508 DVDD.n737 VSS 0.131369f
C18509 DVDD.n738 VSS 0.029427f
C18510 DVDD.n739 VSS 0.131369f
C18511 DVDD.n740 VSS 0.029427f
C18512 DVDD.n741 VSS 0.131369f
C18513 DVDD.n742 VSS 0.029427f
C18514 DVDD.n743 VSS 0.425212f
C18515 DVDD.n744 VSS 0.809162f
C18516 DVDD.t9 VSS 5.27557f
C18517 DVDD.n745 VSS 0.15585f
C18518 DVDD.n746 VSS 0.277706f
C18519 DVDD.n747 VSS 0.277706f
C18520 DVDD.n748 VSS 0.15585f
C18521 DVDD.n749 VSS 0.114418f
C18522 DVDD.n750 VSS 0.114418f
C18523 DVDD.n751 VSS 0.058124f
C18524 DVDD.n752 VSS 0.058124f
C18525 DVDD.n753 VSS 0.058124f
C18526 DVDD.n754 VSS 0.114418f
C18527 DVDD.n755 VSS 0.114418f
C18528 DVDD.n756 VSS 0.114418f
C18529 DVDD.n757 VSS 0.058124f
C18530 DVDD.n758 VSS 0.058124f
C18531 DVDD.n759 VSS 0.058124f
C18532 DVDD.n760 VSS 0.114418f
C18533 DVDD.n761 VSS 0.114418f
C18534 DVDD.n762 VSS 0.114418f
C18535 DVDD.n763 VSS 0.058124f
C18536 DVDD.n764 VSS 0.058124f
C18537 DVDD.n765 VSS 0.058124f
C18538 DVDD.n766 VSS 0.114418f
C18539 DVDD.n767 VSS 0.114418f
C18540 DVDD.n768 VSS 0.114418f
C18541 DVDD.n769 VSS 0.058124f
C18542 DVDD.n770 VSS 0.058124f
C18543 DVDD.n771 VSS 0.058124f
C18544 DVDD.n772 VSS 0.114418f
C18545 DVDD.n773 VSS 0.114418f
C18546 DVDD.n774 VSS 0.114418f
C18547 DVDD.n775 VSS 0.058124f
C18548 DVDD.n776 VSS 0.058124f
C18549 DVDD.n777 VSS 0.058124f
C18550 DVDD.n778 VSS 0.114418f
C18551 DVDD.n779 VSS 0.114418f
C18552 DVDD.n780 VSS 0.114418f
C18553 DVDD.n781 VSS 0.058124f
C18554 DVDD.n782 VSS 0.058124f
C18555 DVDD.n783 VSS 0.058124f
C18556 DVDD.n784 VSS 0.114418f
C18557 DVDD.n785 VSS 0.114418f
C18558 DVDD.n786 VSS 0.114418f
C18559 DVDD.n787 VSS 0.058124f
C18560 DVDD.n788 VSS 0.058124f
C18561 DVDD.n789 VSS 0.058124f
C18562 DVDD.n790 VSS 0.124509f
C18563 DVDD.n791 VSS 0.131369f
C18564 DVDD.n792 VSS 0.026274f
C18565 DVDD.n793 VSS 0.131369f
C18566 DVDD.n794 VSS 0.131369f
C18567 DVDD.n795 VSS 0.026274f
C18568 DVDD.n796 VSS 0.131369f
C18569 DVDD.n797 VSS 0.102976f
C18570 DVDD.n798 VSS 0.131369f
C18571 DVDD.n799 VSS 0.026274f
C18572 DVDD.n800 VSS 0.026274f
C18573 DVDD.n801 VSS 0.026274f
C18574 DVDD.n802 VSS 0.131369f
C18575 DVDD.n803 VSS 0.131369f
C18576 DVDD.n804 VSS 0.131369f
C18577 DVDD.n805 VSS 0.026274f
C18578 DVDD.n806 VSS 0.026274f
C18579 DVDD.n807 VSS 0.025532f
C18580 DVDD.n808 VSS 0.131369f
C18581 DVDD.n809 VSS 0.013137f
C18582 DVDD.n810 VSS 0.131369f
C18583 DVDD.n811 VSS 0.013137f
C18584 DVDD.n812 VSS 0.131369f
C18585 DVDD.n813 VSS 0.013137f
C18586 DVDD.n814 VSS 0.131369f
C18587 DVDD.n815 VSS 0.013137f
C18588 DVDD.n816 VSS 0.131369f
C18589 DVDD.n817 VSS 0.013137f
C18590 DVDD.n818 VSS 0.131369f
C18591 DVDD.n819 VSS 0.013137f
C18592 DVDD.n820 VSS 0.131369f
C18593 DVDD.n821 VSS 0.013137f
C18594 DVDD.n822 VSS 0.131369f
C18595 DVDD.n823 VSS 0.013137f
C18596 DVDD.n824 VSS 0.131369f
C18597 DVDD.n825 VSS 0.013137f
C18598 DVDD.n826 VSS 0.131369f
C18599 DVDD.n827 VSS 0.131369f
C18600 DVDD.n828 VSS 0.131369f
C18601 DVDD.n829 VSS 0.131369f
C18602 DVDD.n830 VSS 0.026274f
C18603 DVDD.n831 VSS 0.026274f
C18604 DVDD.n832 VSS 0.026274f
C18605 DVDD.n833 VSS 0.131369f
C18606 DVDD.n834 VSS 0.131369f
C18607 DVDD.n835 VSS 0.131369f
C18608 DVDD.n836 VSS 0.026274f
C18609 DVDD.n837 VSS 0.026274f
C18610 DVDD.n838 VSS 0.025108f
C18611 DVDD.n839 VSS 0.131369f
C18612 DVDD.n840 VSS 0.013137f
C18613 DVDD.n841 VSS 0.029028f
C18614 DVDD.n842 VSS 0.029062f
C18615 DVDD.n843 VSS 0.033099f
C18616 DVDD.n844 VSS 0.114418f
C18617 DVDD.n845 VSS 0.114418f
C18618 DVDD.n846 VSS 0.114418f
C18619 DVDD.n847 VSS 0.114418f
C18620 DVDD.n848 VSS 0.033368f
C18621 DVDD.n849 VSS 0.030088f
C18622 DVDD.n850 VSS 0.197054f
C18623 DVDD.n851 VSS 0.013137f
C18624 DVDD.n852 VSS 0.066735f
C18625 DVDD.n853 VSS 0.197054f
C18626 DVDD.n854 VSS 0.013137f
C18627 DVDD.n855 VSS 0.032561f
C18628 DVDD.n856 VSS 0.026274f
C18629 DVDD.n857 VSS 0.030088f
C18630 DVDD.n858 VSS 0.044284f
C18631 DVDD.n859 VSS 0.060175f
C18632 DVDD.n860 VSS 0.060175f
C18633 DVDD.n861 VSS 0.173937f
C18634 DVDD.n862 VSS 0.061117f
C18635 DVDD.n863 VSS 0.060739f
C18636 DVDD.n864 VSS 0.033368f
C18637 DVDD.n865 VSS 0.033368f
C18638 DVDD.n866 VSS 0.197054f
C18639 DVDD.n867 VSS 0.220891f
C18640 DVDD.n868 VSS 0.013137f
C18641 DVDD.n869 VSS 0.066735f
C18642 DVDD.n870 VSS 0.548254f
C18643 DVDD.n871 VSS 0.201821f
C18644 DVDD.n872 VSS 0.013137f
C18645 DVDD.n873 VSS 0.048168f
C18646 DVDD.n874 VSS 0.033368f
C18647 DVDD.n875 VSS 0.061117f
C18648 DVDD.n876 VSS 0.026274f
C18649 DVDD.n877 VSS 0.029062f
C18650 DVDD.n878 VSS 0.114418f
C18651 DVDD.n879 VSS 0.114418f
C18652 DVDD.n880 VSS 0.033368f
C18653 DVDD.n881 VSS 0.030088f
C18654 DVDD.n882 VSS 0.197054f
C18655 DVDD.n883 VSS 0.197054f
C18656 DVDD.n884 VSS 0.013137f
C18657 DVDD.n885 VSS 0.066735f
C18658 DVDD.n886 VSS 0.013137f
C18659 DVDD.n887 VSS 0.114418f
C18660 DVDD.n888 VSS 0.114418f
C18661 DVDD.n889 VSS 0.033368f
C18662 DVDD.n890 VSS 0.030088f
C18663 DVDD.n891 VSS 0.197054f
C18664 DVDD.n892 VSS 0.013137f
C18665 DVDD.n893 VSS 0.066735f
C18666 DVDD.n894 VSS 0.197054f
C18667 DVDD.n895 VSS 0.013137f
C18668 DVDD.n896 VSS 0.033368f
C18669 DVDD.n897 VSS 0.026274f
C18670 DVDD.n898 VSS 0.029028f
C18671 DVDD.n899 VSS 0.045979f
C18672 DVDD.n900 VSS 0.060175f
C18673 DVDD.n901 VSS 0.060175f
C18674 DVDD.n902 VSS 0.060175f
C18675 DVDD.n903 VSS 0.026274f
C18676 DVDD.n904 VSS 0.033099f
C18677 DVDD.n905 VSS 0.130242f
C18678 DVDD.n906 VSS 0.197054f
C18679 DVDD.n907 VSS 0.535541f
C18680 DVDD.n908 VSS 0.013137f
C18681 DVDD.n909 VSS 0.066735f
C18682 DVDD.n910 VSS 0.066735f
C18683 DVDD.n911 VSS 0.535541f
C18684 DVDD.n912 VSS 0.197054f
C18685 DVDD.n913 VSS 0.131369f
C18686 DVDD.n914 VSS 0.114418f
C18687 DVDD.n915 VSS 0.114418f
C18688 DVDD.n916 VSS 0.033368f
C18689 DVDD.n917 VSS 0.027333f
C18690 DVDD.n918 VSS 0.029062f
C18691 DVDD.n919 VSS 0.217712f
C18692 DVDD.n920 VSS 0.013137f
C18693 DVDD.n921 VSS 0.131369f
C18694 DVDD.n922 VSS 0.131369f
C18695 DVDD.n923 VSS 0.013137f
C18696 DVDD.n924 VSS 0.013137f
C18697 DVDD.n925 VSS 0.131369f
C18698 DVDD.n926 VSS 0.013137f
C18699 DVDD.n927 VSS 0.131369f
C18700 DVDD.n928 VSS 0.131369f
C18701 DVDD.n929 VSS 0.013137f
C18702 DVDD.n930 VSS 0.114418f
C18703 DVDD.n931 VSS 0.114418f
C18704 DVDD.n932 VSS 0.114418f
C18705 DVDD.n933 VSS 0.029062f
C18706 DVDD.n934 VSS 0.058124f
C18707 DVDD.n935 VSS 0.048706f
C18708 DVDD.n936 VSS 0.114418f
C18709 DVDD.n937 VSS 0.114418f
C18710 DVDD.n938 VSS 0.114418f
C18711 DVDD.n939 VSS 0.114418f
C18712 DVDD.n940 VSS 0.029869f
C18713 DVDD.n941 VSS 0.029062f
C18714 DVDD.n942 VSS 0.225658f
C18715 DVDD.n943 VSS 0.013137f
C18716 DVDD.n944 VSS 0.013137f
C18717 DVDD.n945 VSS 0.131369f
C18718 DVDD.n946 VSS 0.013137f
C18719 DVDD.n947 VSS 0.131369f
C18720 DVDD.n948 VSS 0.131369f
C18721 DVDD.n949 VSS 0.014302f
C18722 DVDD.n950 VSS 0.026274f
C18723 DVDD.n951 VSS 0.023837f
C18724 DVDD.n952 VSS 0.131369f
C18725 DVDD.n953 VSS 0.131369f
C18726 DVDD.n954 VSS 0.013137f
C18727 DVDD.n955 VSS 0.013137f
C18728 DVDD.n956 VSS 0.013137f
C18729 DVDD.n957 VSS 0.750075f
C18730 DVDD.n958 VSS 0.451316f
C18731 DVDD.n959 VSS 0.332131f
C18732 DVDD.n960 VSS 0.451316f
C18733 DVDD.n961 VSS 0.451316f
C18734 DVDD.n962 VSS 0.451316f
C18735 DVDD.n963 VSS 0.451316f
C18736 DVDD.n964 VSS 0.451316f
C18737 DVDD.n965 VSS 0.548254f
C18738 DVDD.n966 VSS 0.750075f
C18739 DVDD.n967 VSS 0.750075f
C18740 DVDD.n968 VSS 0.750075f
C18741 DVDD.n969 VSS 0.451316f
C18742 DVDD.n970 VSS 0.451316f
C18743 DVDD.n971 VSS 0.451316f
C18744 DVDD.n972 VSS 0.332131f
C18745 DVDD.n973 VSS 0.451316f
C18746 DVDD.n974 VSS 0.451316f
C18747 DVDD.n975 VSS 0.451316f
C18748 DVDD.n976 VSS 0.197054f
C18749 DVDD.n977 VSS 0.225658f
C18750 DVDD.n978 VSS 0.013137f
C18751 DVDD.n979 VSS 0.013137f
C18752 DVDD.n980 VSS 0.131369f
C18753 DVDD.n981 VSS 0.013137f
C18754 DVDD.n982 VSS 0.131369f
C18755 DVDD.n983 VSS 0.013137f
C18756 DVDD.n984 VSS 0.131369f
C18757 DVDD.n985 VSS 0.013137f
C18758 DVDD.n986 VSS 0.131369f
C18759 DVDD.n987 VSS 0.013137f
C18760 DVDD.n988 VSS 0.131369f
C18761 DVDD.n989 VSS 0.013137f
C18762 DVDD.n990 VSS 0.131369f
C18763 DVDD.n991 VSS 0.131369f
C18764 DVDD.n992 VSS 0.013137f
C18765 DVDD.n993 VSS 0.013137f
C18766 DVDD.n994 VSS 0.013137f
C18767 DVDD.n995 VSS 0.204999f
C18768 DVDD.n996 VSS 0.029062f
C18769 DVDD.n997 VSS 0.029331f
C18770 DVDD.n998 VSS 0.114418f
C18771 DVDD.n999 VSS 0.15585f
C18772 DVDD.t4 VSS 5.27557f
C18773 DVDD.n1000 VSS 0.124509f
C18774 DVDD.n1001 VSS 0.038139f
C18775 DVDD.n1002 VSS 0.026274f
C18776 DVDD.n1003 VSS 0.217712f
C18777 DVDD.n1004 VSS 0.066735f
C18778 DVDD.n1005 VSS 0.026274f
C18779 DVDD.n1006 VSS 0.030088f
C18780 DVDD.n1007 VSS 0.060175f
C18781 DVDD.n1008 VSS 0.026274f
C18782 DVDD.n1009 VSS 0.066735f
C18783 DVDD.n1010 VSS 0.033368f
C18784 DVDD.n1011 VSS 0.197054f
C18785 DVDD.n1012 VSS 0.197054f
C18786 DVDD.n1013 VSS 0.014726f
C18787 DVDD.n1014 VSS 0.066735f
C18788 DVDD.n1015 VSS 0.451316f
C18789 DVDD.n1016 VSS 0.724649f
C18790 DVDD.n1017 VSS 0.451316f
C18791 DVDD.n1018 VSS 0.344844f
C18792 DVDD.n1019 VSS 0.451316f
C18793 DVDD.n1020 VSS 0.451316f
C18794 DVDD.n1021 VSS 0.451316f
C18795 DVDD.n1022 VSS 0.451316f
C18796 DVDD.n1023 VSS 0.451316f
C18797 DVDD.n1024 VSS 0.724649f
C18798 DVDD.n1025 VSS 0.724649f
C18799 DVDD.n1026 VSS 0.724649f
C18800 DVDD.n1027 VSS 0.451316f
C18801 DVDD.n1028 VSS 0.451316f
C18802 DVDD.n1029 VSS 0.451316f
C18803 DVDD.n1030 VSS 0.451316f
C18804 DVDD.n1031 VSS 0.451316f
C18805 DVDD.n1032 VSS 0.197054f
C18806 DVDD.n1033 VSS 0.026274f
C18807 DVDD.n1034 VSS 0.225658f
C18808 DVDD.n1035 VSS 0.066735f
C18809 DVDD.n1036 VSS 0.066735f
C18810 DVDD.n1037 VSS 0.197054f
C18811 DVDD.n1038 VSS 0.197054f
C18812 DVDD.n1039 VSS 0.013137f
C18813 DVDD.n1040 VSS 0.029062f
C18814 DVDD.n1041 VSS 0.033368f
C18815 DVDD.n1042 VSS 0.033368f
C18816 DVDD.n1043 VSS 0.026274f
C18817 DVDD.n1044 VSS 0.030088f
C18818 DVDD.n1045 VSS 0.060175f
C18819 DVDD.n1046 VSS 0.060739f
C18820 DVDD.n1047 VSS 0.026274f
C18821 DVDD.n1048 VSS 0.030088f
C18822 DVDD.n1049 VSS 0.033368f
C18823 DVDD.n1050 VSS 0.033368f
C18824 DVDD.n1051 VSS 0.197054f
C18825 DVDD.n1052 VSS 0.456124f
C18826 DVDD.n1053 VSS 0.013137f
C18827 DVDD.n1054 VSS 0.066735f
C18828 DVDD.n1056 VSS 0.225658f
C18829 DVDD.n1057 VSS 0.225658f
C18830 DVDD.n1058 VSS 0.216865f
C18831 DVDD.n1059 VSS 0.066735f
C18832 DVDD.n1060 VSS 0.066735f
C18833 DVDD.n1061 VSS 0.066735f
C18834 DVDD.n1062 VSS 0.066735f
C18835 DVDD.n1063 VSS 0.066735f
C18836 DVDD.n1064 VSS 0.066735f
C18837 DVDD.n1065 VSS 0.066735f
C18838 DVDD.n1066 VSS 0.066735f
C18839 DVDD.n1067 VSS 0.066735f
C18840 DVDD.n1068 VSS 0.066735f
C18841 DVDD.n1069 VSS 0.066735f
C18842 DVDD.n1070 VSS 0.197054f
C18843 DVDD.n1072 VSS 0.066735f
C18844 DVDD.n1074 VSS 0.066735f
C18845 DVDD.n1076 VSS 0.066735f
C18846 DVDD.n1078 VSS 0.066735f
C18847 DVDD.n1080 VSS 0.066735f
C18848 DVDD.n1082 VSS 0.066735f
C18849 DVDD.n1084 VSS 0.066735f
C18850 DVDD.n1086 VSS 0.066735f
C18851 DVDD.n1088 VSS 0.066735f
C18852 DVDD.n1090 VSS 0.066735f
C18853 DVDD.n1092 VSS 0.066735f
C18854 DVDD.n1095 VSS 0.120351f
C18855 DVDD.n1096 VSS 0.120351f
C18856 DVDD.n1097 VSS 0.066735f
C18857 DVDD.n1098 VSS 0.066735f
C18858 DVDD.n1099 VSS 0.066735f
C18859 DVDD.n1100 VSS 0.066735f
C18860 DVDD.n1101 VSS 0.066735f
C18861 DVDD.n1102 VSS 0.105095f
C18862 DVDD.n1104 VSS 0.066735f
C18863 DVDD.n1106 VSS 0.066735f
C18864 DVDD.n1108 VSS 0.066735f
C18865 DVDD.n1110 VSS 0.066735f
C18866 DVDD.n1116 VSS 0.120351f
C18867 DVDD.n1118 VSS 0.225658f
C18868 DVDD.n1119 VSS 0.225658f
C18869 DVDD.n1120 VSS 0.459262f
C18870 DVDD.n1121 VSS 0.066735f
C18871 DVDD.n1122 VSS 0.066735f
C18872 DVDD.n1123 VSS 0.066735f
C18873 DVDD.n1124 VSS 0.066735f
C18874 DVDD.n1125 VSS 0.066735f
C18875 DVDD.n1126 VSS 0.066735f
C18876 DVDD.n1127 VSS 0.066735f
C18877 DVDD.n1128 VSS 0.066735f
C18878 DVDD.n1129 VSS 0.066735f
C18879 DVDD.n1130 VSS 0.066735f
C18880 DVDD.n1131 VSS 0.066735f
C18881 DVDD.n1132 VSS 0.197054f
C18882 DVDD.n1134 VSS 0.066735f
C18883 DVDD.n1136 VSS 0.066735f
C18884 DVDD.n1138 VSS 0.066735f
C18885 DVDD.n1140 VSS 0.066735f
C18886 DVDD.n1142 VSS 0.066735f
C18887 DVDD.n1144 VSS 0.066735f
C18888 DVDD.n1146 VSS 0.066735f
C18889 DVDD.n1148 VSS 0.066735f
C18890 DVDD.n1150 VSS 0.066735f
C18891 DVDD.n1152 VSS 0.066735f
C18892 DVDD.n1154 VSS 0.066735f
C18893 DVDD.n1157 VSS 0.225658f
C18894 DVDD.n1158 VSS 0.225658f
C18895 DVDD.n1159 VSS 0.77709f
C18896 DVDD.n1160 VSS 0.066735f
C18897 DVDD.n1161 VSS 0.066735f
C18898 DVDD.n1162 VSS 0.066735f
C18899 DVDD.n1163 VSS 0.066735f
C18900 DVDD.n1164 VSS 0.066735f
C18901 DVDD.n1165 VSS 0.066735f
C18902 DVDD.n1166 VSS 0.066735f
C18903 DVDD.n1167 VSS 0.066735f
C18904 DVDD.n1168 VSS 0.066735f
C18905 DVDD.n1169 VSS 0.066735f
C18906 DVDD.n1170 VSS 0.066735f
C18907 DVDD.n1171 VSS 0.197054f
C18908 DVDD.n1173 VSS 0.066735f
C18909 DVDD.n1175 VSS 0.066735f
C18910 DVDD.n1177 VSS 0.066735f
C18911 DVDD.n1179 VSS 0.066735f
C18912 DVDD.n1181 VSS 0.066735f
C18913 DVDD.n1183 VSS 0.066735f
C18914 DVDD.n1185 VSS 0.066735f
C18915 DVDD.n1187 VSS 0.066735f
C18916 DVDD.n1189 VSS 0.066735f
C18917 DVDD.n1191 VSS 0.066735f
C18918 DVDD.n1193 VSS 0.066735f
C18919 DVDD.n1196 VSS 0.225658f
C18920 DVDD.n1197 VSS 0.225658f
C18921 DVDD.n1198 VSS 0.77709f
C18922 DVDD.n1199 VSS 0.066735f
C18923 DVDD.n1200 VSS 0.066735f
C18924 DVDD.n1201 VSS 0.066735f
C18925 DVDD.n1202 VSS 0.066735f
C18926 DVDD.n1203 VSS 0.066735f
C18927 DVDD.n1204 VSS 0.066735f
C18928 DVDD.n1205 VSS 0.066735f
C18929 DVDD.n1206 VSS 0.066735f
C18930 DVDD.n1207 VSS 0.066735f
C18931 DVDD.n1208 VSS 0.066735f
C18932 DVDD.n1209 VSS 0.066735f
C18933 DVDD.n1210 VSS 0.197054f
C18934 DVDD.n1212 VSS 0.066735f
C18935 DVDD.n1214 VSS 0.066735f
C18936 DVDD.n1216 VSS 0.066735f
C18937 DVDD.n1218 VSS 0.066735f
C18938 DVDD.n1220 VSS 0.066735f
C18939 DVDD.n1222 VSS 0.066735f
C18940 DVDD.n1224 VSS 0.066735f
C18941 DVDD.n1226 VSS 0.066735f
C18942 DVDD.n1228 VSS 0.066735f
C18943 DVDD.n1230 VSS 0.066735f
C18944 DVDD.n1232 VSS 0.066735f
C18945 DVDD.n1235 VSS 0.225658f
C18946 DVDD.n1236 VSS 0.225658f
C18947 DVDD.n1237 VSS 0.459262f
C18948 DVDD.n1238 VSS 0.066735f
C18949 DVDD.n1239 VSS 0.066735f
C18950 DVDD.n1240 VSS 0.05059f
C18951 DVDD.n1241 VSS 0.033368f
C18952 DVDD.n1242 VSS 0.049513f
C18953 DVDD.n1243 VSS 0.066735f
C18954 DVDD.n1244 VSS 0.066735f
C18955 DVDD.n1245 VSS 0.066735f
C18956 DVDD.n1246 VSS 0.066735f
C18957 DVDD.n1247 VSS 0.066735f
C18958 DVDD.n1248 VSS 0.066735f
C18959 DVDD.n1249 VSS 0.197054f
C18960 DVDD.n1251 VSS 0.066735f
C18961 DVDD.n1253 VSS 0.066735f
C18962 DVDD.n1255 VSS 0.066735f
C18963 DVDD.n1257 VSS 0.066735f
C18964 DVDD.n1259 VSS 0.066735f
C18965 DVDD.n1261 VSS 0.066735f
C18966 DVDD.n1263 VSS 0.066735f
C18967 DVDD.n1264 VSS 0.033368f
C18968 DVDD.n1265 VSS 0.033368f
C18969 DVDD.n1267 VSS 0.066735f
C18970 DVDD.n1269 VSS 0.066735f
C18971 DVDD.n1272 VSS 0.105307f
C18972 DVDD.n1273 VSS 0.105307f
C18973 DVDD.n1274 VSS 0.171309f
C18974 DVDD.n1275 VSS 0.066735f
C18975 DVDD.n1276 VSS 0.066735f
C18976 DVDD.n1277 VSS 0.066735f
C18977 DVDD.n1278 VSS 0.066735f
C18978 DVDD.n1279 VSS 0.066735f
C18979 DVDD.n1280 VSS 0.091958f
C18980 DVDD.n1282 VSS 0.066735f
C18981 DVDD.n1284 VSS 0.066735f
C18982 DVDD.n1286 VSS 0.066735f
C18983 DVDD.n1288 VSS 0.066735f
C18984 DVDD.n1294 VSS 0.105307f
C18985 DVDD.n1295 VSS 0.061481f
C18986 DVDD.n1296 VSS 0.360951f
C18987 DVDD.n1297 VSS 0.066735f
C18988 DVDD.n1299 VSS 0.061481f
C18989 DVDD.n1302 VSS 0.360856f
C18990 DVDD.n1303 VSS 0.970017f
C18991 DVDD.n1304 VSS 3.37246f
C18992 DVDD.n1305 VSS 4.58897f
C18993 DVDD.n1306 VSS 0.316328f
C18994 DVDD.n1309 VSS 0.638831f
C18995 DVDD.n1311 VSS 0.061481f
C18996 DVDD.n1312 VSS 0.061481f
C18997 DVDD.n1313 VSS 0.066735f
C18998 DVDD.n1314 VSS 0.352514f
C18999 DVDD.n1317 VSS 0.638831f
C19000 DVDD.n1319 VSS 0.061481f
C19001 DVDD.n1320 VSS 0.061481f
C19002 DVDD.n1321 VSS 0.066735f
C19003 DVDD.n1323 VSS 0.0127f
C19004 DVDD.n1324 VSS 0.025401f
C19005 DVDD.n1325 VSS 0.025401f
C19006 DVDD.n1326 VSS 0.176277f
C19007 DVDD.n1327 VSS 0.0127f
C19008 DVDD.n1328 VSS 0.342557f
C19009 DVDD.n1329 VSS 0.025401f
C19010 DVDD.n1330 VSS 0.348208f
C19011 DVDD.n1332 VSS 0.025401f
C19012 DVDD.n1333 VSS 0.0127f
C19013 DVDD.n1334 VSS 0.342557f
C19014 DVDD.n1335 VSS 0.144644f
C19015 DVDD.n1336 VSS 0.847098f
C19016 DVDD.t0 VSS 32.647602f
C19017 DVDD.n1337 VSS 1.30412f
C19018 DVDD.n1338 VSS 0.025401f
C19019 DVDD.n1339 VSS 0.130026f
C19020 DVDD.n1340 VSS 0.847098f
C19021 DVDD.n1341 VSS 1.30655f
C19022 DVDD.n1342 VSS 1.26891f
C19023 DVDD.n1343 VSS 1.30412f
C19024 DVDD.n1344 VSS 0.025401f
C19025 DVDD.n1345 VSS 0.025401f
C19026 DVDD.n1346 VSS 0.058124f
C19027 DVDD.n1347 VSS 0.058124f
C19028 DVDD.n1348 VSS 0.040796f
C19029 DVDD.n1349 VSS 0.029062f
C19030 DVDD.n1350 VSS 0.058124f
C19031 DVDD.n1351 VSS 0.058124f
C19032 DVDD.n1353 VSS 0.058124f
C19033 DVDD.n1354 VSS 0.348747f
C19034 DVDD.n1357 VSS 0.043021f
C19035 DVDD.n1358 VSS 0.043021f
C19036 DVDD.n1360 VSS 0.342557f
C19037 DVDD.n1362 VSS 0.058124f
C19038 DVDD.n1363 VSS 0.348747f
C19039 DVDD.n1366 VSS 0.043021f
C19040 DVDD.n1367 VSS 0.043021f
C19041 DVDD.n1369 VSS 0.342557f
C19042 DVDD.n1370 VSS 0.244982f
C19043 DVDD.n1371 VSS 0.130026f
C19044 DVDD.n1372 VSS 1.51198f
C19045 DVDD.n1373 VSS 0.063644f
C19046 DVDD.n1374 VSS 1.30655f
C19047 DVDD.n1375 VSS 1.30412f
C19048 DVDD.n1376 VSS 1.26891f
C19049 DVDD.n1377 VSS 0.025401f
C19050 DVDD.n1378 VSS 0.025401f
C19051 DVDD.n1379 VSS 0.058124f
C19052 DVDD.n1380 VSS 0.058124f
C19053 DVDD.n1381 VSS 0.040796f
C19054 DVDD.n1382 VSS 0.298559f
C19055 DVDD.n1383 VSS 0.034259f
C19056 DVDD.n1384 VSS 0.058124f
C19057 DVDD.n1385 VSS 0.025401f
C19058 DVDD.n1386 VSS 0.058124f
C19059 DVDD.n1387 VSS 0.025401f
C19060 DVDD.n1388 VSS 0.058124f
C19061 DVDD.n1389 VSS 0.022343f
C19062 DVDD.n1390 VSS 0.035652f
C19063 DVDD.n1391 VSS 0.029062f
C19064 DVDD.n1392 VSS 0.058124f
C19065 DVDD.n1393 VSS 0.307124f
C19066 DVDD.n1394 VSS 0.029062f
C19067 DVDD.n1395 VSS 0.058124f
C19068 DVDD.n1396 VSS 0.0127f
C19069 DVDD.n1398 VSS 0.0127f
C19070 DVDD.n1399 VSS 0.025401f
C19071 DVDD.n1400 VSS 0.025401f
C19072 DVDD.n1401 VSS 0.342557f
C19073 DVDD.n1402 VSS 0.0127f
C19074 DVDD.n1404 VSS 0.0127f
C19075 DVDD.n1405 VSS 0.025401f
C19076 DVDD.n1408 VSS 0.043021f
C19077 DVDD.n1409 VSS 0.387988f
C19078 DVDD.n1410 VSS 0.058124f
C19079 DVDD.n1411 VSS 0.043021f
C19080 DVDD.n1414 VSS 0.043021f
C19081 DVDD.n1415 VSS 0.387988f
C19082 DVDD.n1416 VSS 0.058124f
C19083 DVDD.n1417 VSS 0.043021f
C19084 DVDD.n1418 VSS 0.348747f
C19085 DVDD.n1419 VSS 0.043021f
C19086 DVDD.n1421 VSS 0.058124f
C19087 DVDD.n1423 VSS 0.043021f
C19088 DVDD.n1424 VSS 0.348747f
C19089 DVDD.n1426 VSS 0.043021f
C19090 DVDD.n1427 VSS 0.043021f
C19091 DVDD.n1429 VSS 0.058124f
C19092 DVDD.n1431 VSS 0.043021f
C19093 DVDD.n1432 VSS 0.348747f
C19094 DVDD.n1434 VSS 0.043021f
C19095 DVDD.n1435 VSS 0.043021f
C19096 DVDD.n1437 VSS 0.029062f
C19097 DVDD.n1438 VSS 0.040796f
C19098 DVDD.n1439 VSS 0.058124f
C19099 DVDD.n1440 VSS 0.058124f
C19100 DVDD.n1441 VSS 0.025401f
C19101 DVDD.n1442 VSS 0.058124f
C19102 DVDD.n1443 VSS 0.025401f
C19103 DVDD.n1444 VSS 0.058124f
C19104 DVDD.n1445 VSS 0.022343f
C19105 DVDD.n1449 VSS 0.043021f
C19106 DVDD.n1450 VSS 0.043021f
C19107 DVDD.n1454 VSS 0.043021f
C19108 DVDD.n1455 VSS 0.043021f
C19109 DVDD.n1457 VSS 0.058124f
C19110 DVDD.n1458 VSS 0.342557f
C19111 DVDD.n1461 VSS 0.058124f
C19112 DVDD.n1462 VSS 0.342557f
C19113 DVDD.n1465 VSS 0.043021f
C19114 DVDD.n1466 VSS 0.043021f
C19115 DVDD.n1470 VSS 0.043021f
C19116 DVDD.n1471 VSS 0.058124f
C19117 DVDD.n1472 VSS 0.043021f
C19118 DVDD.n1476 VSS 0.043021f
C19119 DVDD.n1477 VSS 0.058124f
C19120 DVDD.n1478 VSS 0.043021f
C19121 DVDD.n1481 VSS 0.342557f
C19122 DVDD.n1482 VSS 0.043021f
C19123 DVDD.n1483 VSS 0.348747f
C19124 DVDD.n1485 VSS 0.307124f
C19125 DVDD.n1486 VSS 0.348747f
C19126 DVDD.n1487 VSS 0.043021f
C19127 DVDD.n1488 VSS 0.348747f
C19128 DVDD.n1489 VSS 0.040796f
C19129 DVDD.n1490 VSS 0.058124f
C19130 DVDD.n1491 VSS 0.058124f
C19131 DVDD.n1492 VSS 0.025401f
C19132 DVDD.n1493 VSS 0.058124f
C19133 DVDD.n1494 VSS 0.025401f
C19134 DVDD.n1495 VSS 0.058124f
C19135 DVDD.n1496 VSS 1.62e-19
C19136 DVDD.n1497 VSS 0.181334f
C19137 DVDD.n1500 VSS -0.119061f
C19138 DVDD.n1501 VSS 0.066735f
C19139 DVDD.n1502 VSS 0.638831f
C19140 DVDD.n1506 VSS 0.348208f
C19141 DVDD.n1507 VSS 0.061481f
C19142 DVDD.n1508 VSS 0.501762f
C19143 DVDD.n1509 VSS 0.066735f
C19144 DVDD.n1512 VSS 0.105307f
C19145 DVDD.n1513 VSS 0.105307f
C19146 DVDD.n1514 VSS 0.187625f
C19147 DVDD.n1515 VSS 0.066735f
C19148 DVDD.n1516 VSS 0.066735f
C19149 DVDD.n1517 VSS 0.066735f
C19150 DVDD.n1518 VSS 0.066735f
C19151 DVDD.n1520 VSS 0.091958f
C19152 DVDD.n1522 VSS 0.066735f
C19153 DVDD.n1524 VSS 0.066735f
C19154 DVDD.n1526 VSS 0.066735f
C19155 DVDD.n1527 VSS 0.091958f
C19156 DVDD.n1529 VSS 0.225658f
C19157 DVDD.n1530 VSS 0.225658f
C19158 DVDD.n1531 VSS 0.402053f
C19159 DVDD.n1532 VSS 0.115442f
C19160 DVDD.n1533 VSS 0.066735f
C19161 DVDD.n1534 VSS 0.066735f
C19162 DVDD.n1535 VSS 0.05059f
C19163 DVDD.n1536 VSS 0.033368f
C19164 DVDD.n1537 VSS 0.049513f
C19165 DVDD.n1538 VSS 0.066735f
C19166 DVDD.n1539 VSS 0.048975f
C19167 DVDD.n1540 VSS 0.029062f
C19168 DVDD.n1541 VSS 0.066735f
C19169 DVDD.n1542 VSS 0.066735f
C19170 DVDD.n1543 VSS 0.049244f
C19171 DVDD.n1544 VSS 0.197054f
C19172 DVDD.n1546 VSS 0.066735f
C19173 DVDD.n1548 VSS 0.066735f
C19174 DVDD.n1549 VSS 0.059739f
C19175 DVDD.n1550 VSS 0.029062f
C19176 DVDD.n1552 VSS 0.066735f
C19177 DVDD.n1554 VSS 0.066735f
C19178 DVDD.n1555 VSS 0.033368f
C19179 DVDD.n1556 VSS 0.033368f
C19180 DVDD.n1558 VSS 0.066735f
C19181 DVDD.n1560 VSS 0.066735f
C19182 DVDD.n1561 VSS 0.036872f
C19183 DVDD.n1562 VSS 0.036905f
C19184 DVDD.n1563 VSS 0.451316f
C19185 DVDD.n1564 VSS 0.451316f
C19186 DVDD.n1565 VSS 0.451316f
C19187 DVDD.n1566 VSS 0.451316f
C19188 DVDD.n1567 VSS 0.451316f
C19189 DVDD.n1568 VSS 0.451316f
C19190 DVDD.n1569 VSS 0.451316f
C19191 DVDD.n1570 VSS 0.451316f
C19192 DVDD.n1571 VSS 0.451316f
C19193 DVDD.n1572 VSS 0.451316f
C19194 DVDD.n1573 VSS 0.451316f
C19195 DVDD.n1574 VSS 0.451316f
C19196 DVDD.n1575 VSS 0.451316f
C19197 DVDD.n1576 VSS 0.451316f
C19198 DVDD.n1577 VSS 0.451316f
C19199 DVDD.n1578 VSS 0.451316f
C19200 DVDD.n1579 VSS 0.451316f
C19201 DVDD.n1580 VSS 0.289224f
C19202 DVDD.n1581 VSS 0.451316f
C19203 DVDD.n1582 VSS 0.451316f
C19204 DVDD.n1583 VSS 0.289224f
C19205 DVDD.n1584 VSS 0.861315f
C19206 DVDD.n1585 VSS 0.387751f
C19207 DVDD.n1586 VSS 0.451316f
C19208 DVDD.n1587 VSS 0.543486f
C19209 DVDD.n1588 VSS 0.066735f
C19210 DVDD.n1589 VSS 0.066735f
C19211 DVDD.n1590 VSS 0.05059f
C19212 DVDD.n1591 VSS 0.033368f
C19213 DVDD.n1592 VSS 0.049513f
C19214 DVDD.n1593 VSS 0.066735f
C19215 DVDD.n1594 VSS 0.048975f
C19216 DVDD.n1595 VSS 0.029062f
C19217 DVDD.n1596 VSS 0.066735f
C19218 DVDD.n1597 VSS 0.066735f
C19219 DVDD.n1598 VSS 0.049244f
C19220 DVDD.n1599 VSS 0.115442f
C19221 DVDD.n1600 VSS 0.197054f
C19222 DVDD.n1601 VSS 0.029062f
C19223 DVDD.n1602 VSS 0.066735f
C19224 DVDD.n1603 VSS 0.066735f
C19225 DVDD.n1604 VSS 0.059739f
C19226 DVDD.n1605 VSS 0.029062f
C19227 DVDD.n1606 VSS 0.066735f
C19228 DVDD.n1607 VSS 0.066735f
C19229 DVDD.n1608 VSS 0.033368f
C19230 DVDD.n1609 VSS 0.033368f
C19231 DVDD.n1610 VSS 0.066735f
C19232 DVDD.n1611 VSS 0.066735f
C19233 DVDD.n1619 VSS 0.225658f
C19234 DVDD.n1620 VSS 0.559179f
C19235 DVDD.n1628 VSS 0.225658f
C19236 DVDD.n1629 VSS 0.197054f
C19237 DVDD.n1630 VSS 0.451316f
C19238 DVDD.n1631 VSS 0.451316f
C19239 DVDD.n1632 VSS 0.451316f
C19240 DVDD.n1633 VSS 0.451316f
C19241 DVDD.n1634 VSS 0.451316f
C19242 DVDD.n1635 VSS 0.451316f
C19243 DVDD.n1636 VSS 0.451316f
C19244 DVDD.n1637 VSS 0.451316f
C19245 DVDD.n1638 VSS 0.451316f
C19246 DVDD.n1639 VSS 0.451316f
C19247 DVDD.n1640 VSS 0.451316f
C19248 DVDD.n1641 VSS 0.451316f
C19249 DVDD.n1642 VSS 0.451316f
C19250 DVDD.n1643 VSS 0.451316f
C19251 DVDD.n1644 VSS 0.451316f
C19252 DVDD.n1645 VSS 0.451316f
C19253 DVDD.n1646 VSS 0.451316f
C19254 DVDD.n1647 VSS 0.451316f
C19255 DVDD.n1648 VSS 0.451316f
C19256 DVDD.n1649 VSS 0.451316f
C19257 DVDD.n1650 VSS 0.451316f
C19258 DVDD.n1651 VSS 0.451316f
C19259 DVDD.n1652 VSS 0.451316f
C19260 DVDD.n1653 VSS 0.451316f
C19261 DVDD.n1654 VSS 0.367092f
C19262 DVDD.n1655 VSS 0.451316f
C19263 DVDD.n1656 VSS 0.451316f
C19264 DVDD.n1657 VSS 0.451316f
C19265 DVDD.n1658 VSS 0.451316f
C19266 DVDD.n1659 VSS 0.451316f
C19267 DVDD.n1660 VSS 0.225658f
C19268 DVDD.n1661 VSS 0.115442f
C19269 DVDD.n1662 VSS 0.033368f
C19270 DVDD.n1663 VSS 0.049513f
C19271 DVDD.n1664 VSS 0.029062f
C19272 DVDD.n1665 VSS 0.197054f
C19273 DVDD.n1669 VSS 0.029062f
C19274 DVDD.n1672 VSS 0.033368f
C19275 DVDD.n1673 VSS 0.033368f
C19276 DVDD.n1677 VSS 0.033368f
C19277 DVDD.n1678 VSS 0.225658f
C19278 DVDD.n1679 VSS 0.033368f
C19279 DVDD.n1680 VSS 0.066735f
C19280 DVDD.n1681 VSS 0.066735f
C19281 DVDD.n1682 VSS 0.05059f
C19282 DVDD.n1683 VSS 0.066735f
C19283 DVDD.n1684 VSS 0.048975f
C19284 DVDD.n1685 VSS 0.066735f
C19285 DVDD.n1686 VSS 0.066735f
C19286 DVDD.n1687 VSS 0.049244f
C19287 DVDD.n1688 VSS 0.197054f
C19288 DVDD.n1690 VSS 0.066735f
C19289 DVDD.n1692 VSS 0.066735f
C19290 DVDD.n1693 VSS 0.059739f
C19291 DVDD.n1695 VSS 0.066735f
C19292 DVDD.n1697 VSS 0.066735f
C19293 DVDD.n1699 VSS 0.066735f
C19294 DVDD.n1701 VSS 0.066735f
C19295 DVDD.n1703 VSS 0.105307f
C19296 DVDD.n1704 VSS 0.105307f
C19297 DVDD.n1705 VSS 0.171309f
C19298 DVDD.n1707 VSS 0.066735f
C19299 DVDD.n1708 VSS 0.066735f
C19300 DVDD.n1709 VSS 0.066735f
C19301 DVDD.n1710 VSS 0.066735f
C19302 DVDD.n1711 VSS 0.066735f
C19303 DVDD.n1712 VSS 0.091958f
C19304 DVDD.n1714 VSS 0.066735f
C19305 DVDD.n1716 VSS 0.066735f
C19306 DVDD.n1718 VSS 0.066735f
C19307 DVDD.n1723 VSS 0.210614f
C19308 DVDD.n1724 VSS 0.091958f
C19309 DVDD.n1725 VSS 0.210614f
C19310 DVDD.n1726 VSS 0.210614f
C19311 DVDD.n1727 VSS 0.210614f
C19312 DVDD.n1728 VSS 0.210614f
C19313 DVDD.n1729 VSS 0.210614f
C19314 DVDD.n1730 VSS 0.210614f
C19315 DVDD.n1731 VSS 0.210614f
C19316 DVDD.n1732 VSS 0.210614f
C19317 DVDD.n1733 VSS 0.210614f
C19318 DVDD.n1734 VSS 0.210614f
C19319 DVDD.n1735 VSS 0.210614f
C19320 DVDD.n1736 VSS 0.210614f
C19321 DVDD.n1737 VSS 0.210614f
C19322 DVDD.n1738 VSS 0.210614f
C19323 DVDD.n1739 VSS 0.210614f
C19324 DVDD.n1740 VSS 0.210614f
C19325 DVDD.n1741 VSS 0.066735f
C19326 DVDD.n1742 VSS 0.066735f
C19327 DVDD.n1743 VSS 0.066735f
C19328 DVDD.n1744 VSS 0.066735f
C19329 DVDD.n1745 VSS 0.066735f
C19330 DVDD.n1746 VSS 0.091958f
C19331 DVDD.n1747 VSS 0.559179f
C19332 DVDD.n1748 VSS 0.066735f
C19333 DVDD.n1749 VSS 0.066735f
C19334 DVDD.n1750 VSS 0.066735f
C19335 DVDD.n1757 VSS 0.105307f
C19336 DVDD.n1758 VSS 0.091958f
C19337 DVDD.n1763 VSS 0.105307f
C19338 DVDD.n1764 VSS 0.210614f
C19339 DVDD.n1765 VSS 0.210614f
C19340 DVDD.n1766 VSS 0.210614f
C19341 DVDD.n1767 VSS 0.210614f
C19342 DVDD.n1768 VSS 0.210614f
C19343 DVDD.n1769 VSS 0.184658f
C19344 DVDD.n1770 VSS 0.210614f
C19345 DVDD.n1771 VSS 0.210614f
C19346 DVDD.n1772 VSS 0.210614f
C19347 DVDD.n1773 VSS 0.210614f
C19348 DVDD.n1774 VSS 0.210614f
C19349 DVDD.n1775 VSS 0.210614f
C19350 DVDD.n1776 VSS 0.210614f
C19351 DVDD.n1777 VSS 0.210614f
C19352 DVDD.n1778 VSS 0.210614f
C19353 DVDD.n1779 VSS 0.184658f
C19354 DVDD.n1780 VSS 0.171309f
C19355 DVDD.n1781 VSS 0.210614f
C19356 DVDD.n1782 VSS 0.210614f
C19357 DVDD.n1783 VSS 0.210614f
C19358 DVDD.n1784 VSS 0.105307f
C19359 DVDD.n1790 VSS 0.091958f
C19360 DVDD.n1792 VSS 0.062794f
C19361 DVDD.n1793 VSS 0.062794f
C19362 DVDD.n1794 VSS 0.062794f
C19363 DVDD.n1795 VSS 0.062794f
C19364 DVDD.n1796 VSS 0.062794f
C19365 DVDD.n1797 VSS 0.091958f
C19366 DVDD.n1799 VSS 0.181162f
C19367 DVDD.n1800 VSS 0.225658f
C19368 DVDD.n1801 VSS 0.367092f
C19369 DVDD.n1802 VSS 0.062794f
C19370 DVDD.n1803 VSS 0.062794f
C19371 DVDD.n1804 VSS 0.062794f
C19372 DVDD.n1805 VSS 0.062794f
C19373 DVDD.n1806 VSS 0.062794f
C19374 DVDD.n1807 VSS 0.062794f
C19375 DVDD.n1808 VSS 0.062794f
C19376 DVDD.n1809 VSS 0.062794f
C19377 DVDD.n1810 VSS 0.062794f
C19378 DVDD.n1811 VSS 0.062794f
C19379 DVDD.n1812 VSS 0.062794f
C19380 DVDD.n1813 VSS 0.079457f
C19381 DVDD.n1814 VSS 0.197054f
C19382 DVDD.n1816 VSS 0.062794f
C19383 DVDD.n1818 VSS 0.062794f
C19384 DVDD.n1820 VSS 0.062794f
C19385 DVDD.n1822 VSS 0.062794f
C19386 DVDD.n1824 VSS 0.062794f
C19387 DVDD.n1826 VSS 0.062794f
C19388 DVDD.n1828 VSS 0.062794f
C19389 DVDD.n1830 VSS 0.062794f
C19390 DVDD.n1832 VSS 0.062794f
C19391 DVDD.n1834 VSS 0.062794f
C19392 DVDD.n1835 VSS 0.451316f
C19393 DVDD.n1836 VSS 0.451316f
C19394 DVDD.n1837 VSS 0.451316f
C19395 DVDD.n1838 VSS 0.395696f
C19396 DVDD.n1839 VSS 0.451316f
C19397 DVDD.n1840 VSS 0.451316f
C19398 DVDD.n1841 VSS 0.543486f
C19399 DVDD.n1842 VSS 0.861315f
C19400 DVDD.n1843 VSS 0.451316f
C19401 DVDD.n1844 VSS 0.451316f
C19402 DVDD.n1845 VSS 0.451316f
C19403 DVDD.n1846 VSS 0.451316f
C19404 DVDD.n1847 VSS 0.451316f
C19405 DVDD.n1848 VSS 0.451316f
C19406 DVDD.n1849 VSS 0.451316f
C19407 DVDD.n1850 VSS 0.451316f
C19408 DVDD.n1851 VSS 0.451316f
C19409 DVDD.n1852 VSS 0.451316f
C19410 DVDD.n1853 VSS 0.197054f
C19411 DVDD.n1856 VSS 0.05059f
C19412 DVDD.n1857 VSS 0.033368f
C19413 DVDD.n1860 VSS 0.048975f
C19414 DVDD.n1861 VSS 0.029062f
C19415 DVDD.n1864 VSS 0.049244f
C19416 DVDD.n1865 VSS 0.115442f
C19417 DVDD.n1866 VSS 0.036898f
C19418 DVDD.n1867 VSS 0.011442f
C19419 DVDD.n1868 VSS 0.022884f
C19420 DVDD.n1869 VSS 0.022884f
C19421 DVDD.n1870 VSS 0.301797f
C19422 DVDD.n1871 VSS 0.033368f
C19423 DVDD.n1872 VSS 0.220876f
C19424 DVDD.n1873 VSS 0.011442f
C19425 DVDD.n1874 VSS 0.033368f
C19426 DVDD.n1875 VSS 0.13031f
C19427 DVDD.t25 VSS 1.69508f
C19428 DVDD.n1876 VSS 0.13031f
C19429 DVDD.n1878 VSS 0.022884f
C19430 DVDD.n1879 VSS 0.022884f
C19431 DVDD.n1880 VSS 0.011442f
C19432 DVDD.n1881 VSS 0.011442f
C19433 DVDD.n1882 VSS 0.220795f
C19434 DVDD.n1883 VSS 0.301873f
C19435 DVDD.n1884 VSS 0.036883f
C19436 DVDD.n1885 VSS 0.029062f
C19437 DVDD.n1886 VSS 0.059739f
C19438 DVDD.n1887 VSS 0.029062f
C19439 DVDD.n1888 VSS 0.033368f
C19440 DVDD.n1889 VSS 0.033368f
C19441 DVDD.n1891 VSS 0.225658f
C19442 DVDD.n1892 VSS 0.367092f
C19443 DVDD.n1893 VSS 0.066735f
C19444 DVDD.n1894 VSS 0.066735f
C19445 DVDD.n1895 VSS 0.049513f
C19446 DVDD.n1896 VSS 0.066735f
C19447 DVDD.n1897 VSS 0.066735f
C19448 DVDD.n1898 VSS 0.066735f
C19449 DVDD.n1899 VSS 0.197054f
C19450 DVDD.n1900 VSS 0.066735f
C19451 DVDD.n1901 VSS 0.066735f
C19452 DVDD.n1902 VSS 0.066735f
C19453 DVDD.n1903 VSS 0.066735f
C19454 DVDD.n1904 VSS 0.066735f
C19455 DVDD.n1905 VSS 0.451316f
C19456 DVDD.n1906 VSS 0.451316f
C19457 DVDD.n1907 VSS 0.451316f
C19458 DVDD.n1908 VSS 0.451316f
C19459 DVDD.n1909 VSS 0.451316f
C19460 DVDD.n1910 VSS 0.451316f
C19461 DVDD.n1911 VSS 0.451316f
C19462 DVDD.n1912 VSS 0.451316f
C19463 DVDD.n1913 VSS 0.451316f
C19464 DVDD.n1914 VSS 0.451316f
C19465 DVDD.n1915 VSS 0.451316f
C19466 DVDD.n1916 VSS 0.543486f
C19467 DVDD.n1917 VSS 0.543486f
C19468 DVDD.n1918 VSS 0.451316f
C19469 DVDD.n1919 VSS 0.451316f
C19470 DVDD.n1920 VSS 0.451316f
C19471 DVDD.n1921 VSS 0.220891f
C19472 DVDD.n1922 VSS 0.276511f
C19473 DVDD.n1923 VSS 0.276511f
C19474 DVDD.n1924 VSS 0.861315f
C19475 DVDD.n1925 VSS 0.276511f
C19476 DVDD.n1926 VSS 0.451316f
C19477 DVDD.n1927 VSS 0.861315f
C19478 DVDD.n1928 VSS 0.451316f
C19479 DVDD.n1929 VSS 0.861315f
C19480 DVDD.n1930 VSS 0.451316f
C19481 DVDD.n1931 VSS 0.451316f
C19482 DVDD.n1932 VSS 0.451316f
C19483 DVDD.n1933 VSS 0.451316f
C19484 DVDD.n1934 VSS 0.451316f
C19485 DVDD.n1935 VSS 0.451316f
C19486 DVDD.n1936 VSS 0.451316f
C19487 DVDD.n1937 VSS 0.451316f
C19488 DVDD.n1938 VSS 0.451316f
C19489 DVDD.n1939 VSS 0.451316f
C19490 DVDD.n1940 VSS 0.451316f
C19491 DVDD.n1941 VSS 0.367092f
C19492 DVDD.n1942 VSS 0.451316f
C19493 DVDD.n1943 VSS 0.451316f
C19494 DVDD.n1944 VSS 0.451316f
C19495 DVDD.n1945 VSS 0.451316f
C19496 DVDD.n1946 VSS 0.451316f
C19497 DVDD.n1947 VSS 0.225658f
C19498 DVDD.n1949 VSS 0.029062f
C19499 DVDD.n1953 VSS 0.029062f
C19500 DVDD.n1954 VSS 0.197054f
C19501 DVDD.n1958 VSS 0.029062f
C19502 DVDD.n1963 VSS 0.066735f
C19503 DVDD.n1964 VSS 0.066735f
C19504 DVDD.n1965 VSS 0.066735f
C19505 DVDD.n1966 VSS 0.057855f
C19506 DVDD.n1967 VSS 0.046553f
C19507 DVDD.n1968 VSS 0.066735f
C19508 DVDD.n1969 VSS 0.066735f
C19509 DVDD.n1970 VSS 0.066735f
C19510 DVDD.n1971 VSS 0.066735f
C19511 DVDD.n1972 VSS 0.063506f
C19512 DVDD.n1973 VSS 0.197054f
C19513 DVDD.n1974 VSS 0.066735f
C19514 DVDD.n1975 VSS 0.066735f
C19515 DVDD.n1976 VSS 0.045477f
C19516 DVDD.n1977 VSS 0.058932f
C19517 DVDD.n1978 VSS 0.066735f
C19518 DVDD.n1979 VSS 0.066735f
C19519 DVDD.n1980 VSS 0.066735f
C19520 DVDD.n1981 VSS 0.066735f
C19521 DVDD.n1982 VSS 0.04763f
C19522 DVDD.n1983 VSS 0.0369f
C19523 DVDD.n1988 VSS 0.451316f
C19524 DVDD.n1989 VSS 0.451316f
C19525 DVDD.n1990 VSS 0.451316f
C19526 DVDD.n1991 VSS 0.451316f
C19527 DVDD.n1992 VSS 0.451316f
C19528 DVDD.n1993 VSS 0.451316f
C19529 DVDD.n1994 VSS 0.451316f
C19530 DVDD.n1995 VSS 0.451316f
C19531 DVDD.n1996 VSS 0.451316f
C19532 DVDD.n1997 VSS 0.451316f
C19533 DVDD.n1998 VSS 0.451316f
C19534 DVDD.n1999 VSS 0.451316f
C19535 DVDD.n2000 VSS 0.451316f
C19536 DVDD.n2001 VSS 0.451316f
C19537 DVDD.n2002 VSS 0.451316f
C19538 DVDD.n2003 VSS 0.263798f
C19539 DVDD.n2004 VSS 0.861315f
C19540 DVDD.n2005 VSS 0.413177f
C19541 DVDD.n2006 VSS 0.451316f
C19542 DVDD.n2007 VSS 0.451316f
C19543 DVDD.n2008 VSS 0.451316f
C19544 DVDD.n2009 VSS 0.451316f
C19545 DVDD.n2010 VSS 0.451316f
C19546 DVDD.n2011 VSS 0.451316f
C19547 DVDD.n2012 VSS 0.451316f
C19548 DVDD.n2013 VSS 0.451316f
C19549 DVDD.n2014 VSS 0.451316f
C19550 DVDD.n2015 VSS 0.451316f
C19551 DVDD.n2016 VSS 0.062794f
C19552 DVDD.n2017 VSS 0.062794f
C19553 DVDD.n2018 VSS 0.062794f
C19554 DVDD.n2019 VSS 0.062794f
C19555 DVDD.n2020 VSS 0.062794f
C19556 DVDD.n2021 VSS 0.062794f
C19557 DVDD.n2022 VSS 0.062794f
C19558 DVDD.n2023 VSS 0.062794f
C19559 DVDD.n2024 VSS 0.062794f
C19560 DVDD.n2025 VSS 0.062794f
C19561 DVDD.n2026 VSS 0.062794f
C19562 DVDD.n2028 VSS 0.181162f
C19563 DVDD.n2029 VSS 0.225658f
C19564 DVDD.n2030 VSS 0.367092f
C19565 DVDD.n2031 VSS 0.062794f
C19566 DVDD.n2032 VSS 0.062794f
C19567 DVDD.n2033 VSS 0.062794f
C19568 DVDD.n2034 VSS 0.062794f
C19569 DVDD.n2035 VSS 0.031397f
C19570 DVDD.n2036 VSS 0.031397f
C19571 DVDD.n2037 VSS 0.031397f
C19572 DVDD.n2038 VSS 0.031397f
C19573 DVDD.n2039 VSS 0.031397f
C19574 DVDD.n2040 VSS 0.031397f
C19575 DVDD.n2041 VSS 0.031397f
C19576 DVDD.n2042 VSS 0.031836f
C19577 DVDD.n2043 VSS 0.197054f
C19578 DVDD.n2044 VSS 0.031397f
C19579 DVDD.n2045 VSS 0.031397f
C19580 DVDD.n2046 VSS 0.031397f
C19581 DVDD.n2047 VSS 0.031397f
C19582 DVDD.n2048 VSS 0.031397f
C19583 DVDD.n2049 VSS 0.031397f
C19584 DVDD.n2050 VSS 0.031397f
C19585 DVDD.n2052 VSS 0.044311f
C19586 DVDD.n2054 VSS 0.062794f
C19587 DVDD.n2056 VSS 0.062794f
C19588 DVDD.n2057 VSS 0.451316f
C19589 DVDD.n2058 VSS 0.451316f
C19590 DVDD.n2059 VSS 0.451316f
C19591 DVDD.n2060 VSS 0.395696f
C19592 DVDD.n2061 VSS 0.451316f
C19593 DVDD.n2062 VSS 0.451316f
C19594 DVDD.n2063 VSS 0.543486f
C19595 DVDD.n2064 VSS 0.451316f
C19596 DVDD.n2065 VSS 0.451316f
C19597 DVDD.n2066 VSS 0.451316f
C19598 DVDD.n2067 VSS 0.451316f
C19599 DVDD.n2068 VSS 0.451316f
C19600 DVDD.n2069 VSS 0.451316f
C19601 DVDD.n2070 VSS 0.451316f
C19602 DVDD.n2071 VSS 0.451316f
C19603 DVDD.n2072 VSS 0.451316f
C19604 DVDD.n2073 VSS 0.451316f
C19605 DVDD.n2074 VSS 0.197054f
C19606 DVDD.n2075 VSS 0.029062f
C19607 DVDD.n2076 VSS 0.029062f
C19608 DVDD.n2077 VSS 0.029062f
C19609 DVDD.n2078 VSS 0.029062f
C19610 DVDD.n2079 VSS 0.029062f
C19611 DVDD.n2080 VSS 0.029062f
C19612 DVDD.n2081 VSS 0.029062f
C19613 DVDD.n2082 VSS 0.029062f
C19614 DVDD.n2083 VSS 0.029062f
C19615 DVDD.n2084 VSS 0.029062f
C19616 DVDD.n2085 VSS 0.029062f
C19617 DVDD.n2086 VSS 0.029062f
C19618 DVDD.n2087 VSS 0.029062f
C19619 DVDD.n2088 VSS 0.029062f
C19620 DVDD.n2089 VSS 0.029062f
C19621 DVDD.n2090 VSS 0.057317f
C19622 DVDD.n2094 VSS 0.03875f
C19623 DVDD.n2096 VSS 0.225658f
C19624 DVDD.n2097 VSS 0.367092f
C19625 DVDD.n2098 VSS 0.066735f
C19626 DVDD.n2099 VSS 0.066735f
C19627 DVDD.n2100 VSS 0.066735f
C19628 DVDD.n2101 VSS 0.197054f
C19629 DVDD.n2102 VSS 0.066735f
C19630 DVDD.n2105 VSS 0.451316f
C19631 DVDD.n2106 VSS 0.451316f
C19632 DVDD.n2107 VSS 0.451316f
C19633 DVDD.n2108 VSS 0.451316f
C19634 DVDD.n2109 VSS 0.451316f
C19635 DVDD.n2110 VSS 0.451316f
C19636 DVDD.n2111 VSS 0.451316f
C19637 DVDD.n2112 VSS 0.451316f
C19638 DVDD.n2113 VSS 0.451316f
C19639 DVDD.n2114 VSS 0.451316f
C19640 DVDD.n2115 VSS 0.451316f
C19641 DVDD.n2116 VSS 0.861315f
C19642 DVDD.n2117 VSS 0.543486f
C19643 DVDD.n2118 VSS 0.451316f
C19644 DVDD.n2119 VSS 0.276511f
C19645 DVDD.n2120 VSS 0.197054f
C19646 DVDD.n2121 VSS 0.029062f
C19647 DVDD.n2122 VSS 0.029062f
C19648 DVDD.n2123 VSS 0.029062f
C19649 DVDD.n2124 VSS 0.029062f
C19650 DVDD.n2125 VSS 0.029062f
C19651 DVDD.n2126 VSS 0.029062f
C19652 DVDD.n2127 VSS 0.029062f
C19653 DVDD.n2128 VSS 0.029062f
C19654 DVDD.n2129 VSS 0.066735f
C19655 DVDD.n2130 VSS 0.066735f
C19656 DVDD.n2131 VSS 0.066735f
C19657 DVDD.n2132 VSS 0.066735f
C19658 DVDD.n2133 VSS 0.066735f
C19659 DVDD.n2134 VSS 0.066735f
C19660 DVDD.n2135 VSS 0.066735f
C19661 DVDD.n2136 VSS 0.057317f
C19662 DVDD.n2137 VSS 0.029062f
C19663 DVDD.n2138 VSS 0.029062f
C19664 DVDD.n2139 VSS 0.029062f
C19665 DVDD.n2140 VSS 0.029062f
C19666 DVDD.n2141 VSS 0.029062f
C19667 DVDD.n2142 VSS 0.029062f
C19668 DVDD.n2143 VSS 0.029062f
C19669 DVDD.n2149 VSS 0.225658f
C19670 DVDD.n2150 VSS 0.034444f
C19671 DVDD.n2151 VSS 0.197054f
C19672 DVDD.n2152 VSS 0.451316f
C19673 DVDD.n2153 VSS 0.451316f
C19674 DVDD.n2154 VSS 0.451316f
C19675 DVDD.n2155 VSS 0.451316f
C19676 DVDD.n2156 VSS 0.451316f
C19677 DVDD.n2157 VSS 0.451316f
C19678 DVDD.n2158 VSS 0.451316f
C19679 DVDD.n2159 VSS 0.451316f
C19680 DVDD.n2160 VSS 0.451316f
C19681 DVDD.n2161 VSS 0.451316f
C19682 DVDD.n2162 VSS 0.451316f
C19683 DVDD.n2163 VSS 0.451316f
C19684 DVDD.n2164 VSS 0.451316f
C19685 DVDD.n2165 VSS 0.451316f
C19686 DVDD.n2166 VSS 0.451316f
C19687 DVDD.n2167 VSS 0.360735f
C19688 DVDD.n2168 VSS 0.451316f
C19689 DVDD.n2169 VSS 0.451316f
C19690 DVDD.n2170 VSS 0.451316f
C19691 DVDD.n2171 VSS 0.225658f
C19692 DVDD.n2172 VSS 0.029062f
C19693 DVDD.n2173 VSS 0.029062f
C19694 DVDD.n2174 VSS 0.029062f
C19695 DVDD.n2175 VSS 0.029062f
C19696 DVDD.n2176 VSS 0.029062f
C19697 DVDD.n2177 VSS 0.029062f
C19698 DVDD.n2178 VSS 0.029062f
C19699 DVDD.n2179 VSS 0.029062f
C19700 DVDD.n2180 VSS 0.029062f
C19701 DVDD.n2181 VSS 0.029062f
C19702 DVDD.n2182 VSS 0.029062f
C19703 DVDD.n2183 VSS 0.029062f
C19704 DVDD.n2184 VSS 0.029062f
C19705 DVDD.n2185 VSS 0.029062f
C19706 DVDD.n2186 VSS 0.029062f
C19707 DVDD.n2187 VSS 0.057317f
C19708 DVDD.n2191 VSS 0.03875f
C19709 DVDD.n2193 VSS 0.338487f
C19710 DVDD.n2194 VSS 0.066735f
C19711 DVDD.n2195 VSS 0.066735f
C19712 DVDD.n2196 VSS 0.066735f
C19713 DVDD.n2197 VSS 0.387751f
C19714 DVDD.n2198 VSS 0.543486f
C19715 DVDD.n2199 VSS 0.543486f
C19716 DVDD.n2200 VSS 0.861315f
C19717 DVDD.n2201 VSS 0.451316f
C19718 DVDD.n2202 VSS 0.451316f
C19719 DVDD.n2203 VSS 0.861315f
C19720 DVDD.n2204 VSS 0.451316f
C19721 DVDD.n2205 VSS 0.543486f
C19722 DVDD.n2206 VSS 0.289224f
C19723 DVDD.n2207 VSS 0.225658f
C19724 DVDD.n2208 VSS 0.387751f
C19725 DVDD.n2209 VSS 0.451316f
C19726 DVDD.n2210 VSS 0.451316f
C19727 DVDD.n2212 VSS 0.029062f
C19728 DVDD.n2216 VSS 0.029062f
C19729 DVDD.n2217 VSS 0.197054f
C19730 DVDD.n2221 VSS 0.029062f
C19731 DVDD.n2226 VSS 0.066735f
C19732 DVDD.n2227 VSS 0.066735f
C19733 DVDD.n2228 VSS 0.066735f
C19734 DVDD.n2229 VSS 0.057855f
C19735 DVDD.n2230 VSS 0.046553f
C19736 DVDD.n2231 VSS 0.066735f
C19737 DVDD.n2232 VSS 0.066735f
C19738 DVDD.n2233 VSS 0.066735f
C19739 DVDD.n2234 VSS 0.066735f
C19740 DVDD.n2235 VSS 0.063506f
C19741 DVDD.n2236 VSS 0.197054f
C19742 DVDD.n2237 VSS 0.066735f
C19743 DVDD.n2238 VSS 0.066735f
C19744 DVDD.n2239 VSS 0.045477f
C19745 DVDD.n2240 VSS 0.058932f
C19746 DVDD.n2241 VSS 0.066735f
C19747 DVDD.n2242 VSS 0.066735f
C19748 DVDD.n2243 VSS 0.066735f
C19749 DVDD.n2244 VSS 0.066735f
C19750 DVDD.n2245 VSS 0.04763f
C19751 DVDD.n2246 VSS 0.033368f
C19752 DVDD.n2251 VSS 0.451316f
C19753 DVDD.n2252 VSS 0.451316f
C19754 DVDD.n2253 VSS 0.451316f
C19755 DVDD.n2254 VSS 0.451316f
C19756 DVDD.n2255 VSS 0.451316f
C19757 DVDD.n2256 VSS 0.451316f
C19758 DVDD.n2257 VSS 0.451316f
C19759 DVDD.n2258 VSS 0.451316f
C19760 DVDD.n2259 VSS 0.451316f
C19761 DVDD.n2260 VSS 0.451316f
C19762 DVDD.n2261 VSS 0.451316f
C19763 DVDD.n2262 VSS 0.451316f
C19764 DVDD.n2263 VSS 0.451316f
C19765 DVDD.n2264 VSS 0.451316f
C19766 DVDD.n2265 VSS 0.451316f
C19767 DVDD.n2266 VSS 0.451316f
C19768 DVDD.n2267 VSS 0.451316f
C19769 DVDD.n2268 VSS 0.451316f
C19770 DVDD.n2269 VSS 0.451316f
C19771 DVDD.n2270 VSS 0.451316f
C19772 DVDD.n2271 VSS 0.451316f
C19773 DVDD.n2272 VSS 0.451316f
C19774 DVDD.n2273 VSS 0.451316f
C19775 DVDD.n2274 VSS 0.451316f
C19776 DVDD.n2275 VSS 0.451316f
C19777 DVDD.n2276 VSS 0.451316f
C19778 DVDD.n2284 VSS 0.127013f
C19779 DVDD.n2285 VSS 0.197054f
C19780 DVDD.n2289 VSS 0.029062f
C19781 DVDD.n2290 VSS 0.029062f
C19782 DVDD.n2291 VSS 0.033368f
C19783 DVDD.n2292 VSS 0.225658f
C19784 DVDD.n2293 VSS 0.033368f
C19785 DVDD.n2294 VSS 0.225658f
C19786 DVDD.n2295 VSS 0.197054f
C19787 DVDD.n2296 VSS 0.04763f
C19788 DVDD.n2297 VSS 0.046553f
C19789 DVDD.n2298 VSS 0.045477f
C19790 DVDD.n2299 VSS 0.066735f
C19791 DVDD.n2300 VSS 0.066735f
C19792 DVDD.n2301 VSS 0.058932f
C19793 DVDD.n2302 VSS 0.066735f
C19794 DVDD.n2303 VSS 0.066735f
C19795 DVDD.n2304 VSS 0.066735f
C19796 DVDD.n2305 VSS 0.066735f
C19797 DVDD.n2306 VSS 0.056779f
C19798 DVDD.n2307 VSS 0.197054f
C19799 DVDD.n2308 VSS 0.451316f
C19800 DVDD.n2309 VSS 0.451316f
C19801 DVDD.n2310 VSS 0.451316f
C19802 DVDD.n2311 VSS 0.451316f
C19803 DVDD.n2312 VSS 0.451316f
C19804 DVDD.n2313 VSS 0.451316f
C19805 DVDD.n2314 VSS 0.451316f
C19806 DVDD.n2315 VSS 0.276511f
C19807 DVDD.n2316 VSS 0.220891f
C19808 DVDD.n2318 VSS 0.066735f
C19809 DVDD.n2320 VSS 0.066735f
C19810 DVDD.n2322 VSS 0.066735f
C19811 DVDD.n2323 VSS 0.057855f
C19812 DVDD.n2325 VSS 0.066735f
C19813 DVDD.n2327 VSS 0.066735f
C19814 DVDD.n2329 VSS 0.066735f
C19815 DVDD.n2331 VSS 0.066735f
C19816 DVDD.n2334 VSS 0.042106f
C19817 DVDD.n2335 VSS -1.46111f
C19818 DVDD.n2336 VSS 0.058124f
C19819 DVDD.n2340 VSS 0.042106f
C19820 DVDD.n2341 VSS 0.672082f
C19821 DVDD.n2342 VSS 2.21687f
C19822 DVDD.n2343 VSS 3.24347f
C19823 DVDD.n2345 VSS 0.033368f
C19824 DVDD.n2346 VSS 0.042106f
C19825 DVDD.n2348 VSS 0.042106f
C19826 DVDD.n2350 VSS 0.033368f
C19827 DVDD.n2351 VSS 0.042106f
C19828 DVDD.n2352 VSS 0.042106f
C19829 DVDD.n2353 VSS 0.058124f
C19830 DVDD.n2355 VSS 0.03875f
C19831 DVDD.n2358 VSS 0.042106f
C19832 DVDD.n2359 VSS 0.058124f
C19833 DVDD.n2363 VSS 0.042106f
C19834 DVDD.n2365 VSS 0.042106f
C19835 DVDD.n2366 VSS 0.042106f
C19836 DVDD.n2367 VSS 0.059201f
C19837 DVDD.n2368 VSS 0.23977f
C19838 DVDD.n2369 VSS 0.034444f
C19839 DVDD.n2370 VSS 0.379733f
C19840 DVDD.n2372 VSS 0.225658f
C19841 DVDD.n2374 VSS 0.225658f
C19842 DVDD.n2375 VSS 0.197054f
C19843 DVDD.n2376 VSS 0.04763f
C19844 DVDD.n2377 VSS 0.046553f
C19845 DVDD.n2378 VSS 0.045477f
C19846 DVDD.n2379 VSS 0.066735f
C19847 DVDD.n2380 VSS 0.066735f
C19848 DVDD.n2381 VSS 0.058932f
C19849 DVDD.n2382 VSS 0.066735f
C19850 DVDD.n2383 VSS 0.066735f
C19851 DVDD.n2384 VSS 0.066735f
C19852 DVDD.n2385 VSS 0.066735f
C19853 DVDD.n2386 VSS 0.056779f
C19854 DVDD.n2387 VSS 0.127013f
C19855 DVDD.n2388 VSS 0.360735f
C19856 DVDD.n2390 VSS 0.066735f
C19857 DVDD.n2392 VSS 0.066735f
C19858 DVDD.n2394 VSS 0.066735f
C19859 DVDD.n2395 VSS 0.057855f
C19860 DVDD.n2397 VSS 0.066735f
C19861 DVDD.n2399 VSS 0.066735f
C19862 DVDD.n2401 VSS 0.066735f
C19863 DVDD.n2403 VSS 0.066735f
C19864 DVDD.n2404 VSS 0.036872f
C19865 DVDD.n2405 VSS 0.011442f
C19866 DVDD.n2406 VSS 0.011442f
C19867 DVDD.n2407 VSS 0.011442f
C19868 DVDD.n2408 VSS 0.011442f
C19869 DVDD.n2409 VSS 0.0369f
C19870 DVDD.n2410 VSS 0.036871f
C19871 DVDD.n2411 VSS 0.301841f
C19872 DVDD.n2412 VSS 0.220837f
C19873 DVDD.n2413 VSS 0.033368f
C19874 DVDD.n2414 VSS 0.022884f
C19875 DVDD.n2415 VSS 0.022884f
C19876 DVDD.n2416 VSS 0.033368f
C19877 DVDD.n2417 VSS 0.13031f
C19878 DVDD.t31 VSS 1.69508f
C19879 DVDD.n2418 VSS 0.13031f
C19880 DVDD.n2419 VSS 0.033368f
C19881 DVDD.n2420 VSS 0.022884f
C19882 DVDD.n2421 VSS 0.022884f
C19883 DVDD.n2422 VSS 0.033368f
C19884 DVDD.n2423 VSS 0.220876f
C19885 DVDD.n2424 VSS 0.301797f
C19886 DVDD.n2425 VSS 0.036905f
C19887 DVDD.n2426 VSS 0.029062f
C19888 DVDD.n2427 VSS 0.036872f
C19889 DVDD.n2428 VSS 0.011442f
C19890 DVDD.n2429 VSS 0.011442f
C19891 DVDD.n2430 VSS 0.011442f
C19892 DVDD.n2431 VSS 0.011442f
C19893 DVDD.n2432 VSS 0.0369f
C19894 DVDD.n2433 VSS 0.036871f
C19895 DVDD.n2434 VSS 0.301841f
C19896 DVDD.n2435 VSS 0.220837f
C19897 DVDD.n2436 VSS 0.033368f
C19898 DVDD.n2437 VSS 0.022884f
C19899 DVDD.n2438 VSS 0.022884f
C19900 DVDD.n2439 VSS 0.033368f
C19901 DVDD.n2440 VSS 0.13031f
C19902 DVDD.t37 VSS 1.69508f
C19903 DVDD.n2441 VSS 0.13031f
C19904 DVDD.n2442 VSS 0.033368f
C19905 DVDD.n2443 VSS 0.022884f
C19906 DVDD.n2444 VSS 0.022884f
C19907 DVDD.n2445 VSS 0.033368f
C19908 DVDD.n2446 VSS 0.220876f
C19909 DVDD.n2447 VSS 0.301797f
C19910 DVDD.n2448 VSS 0.036905f
C19911 DVDD.n2449 VSS 0.029062f
C19912 DVDD.n2450 VSS 0.036872f
C19913 DVDD.n2451 VSS 0.402053f
C19914 DVDD.n2458 VSS 0.451316f
C19915 DVDD.n2459 VSS 0.451316f
C19916 DVDD.n2460 VSS 0.451316f
C19917 DVDD.n2461 VSS 0.451316f
C19918 DVDD.n2462 VSS 0.451316f
C19919 DVDD.n2463 VSS 0.451316f
C19920 DVDD.n2464 VSS 0.451316f
C19921 DVDD.n2465 VSS 0.360735f
C19922 DVDD.n2466 VSS 0.375037f
C19923 DVDD.n2467 VSS 0.861315f
C19924 DVDD.n2468 VSS 0.543486f
C19925 DVDD.n2469 VSS 0.451316f
C19926 DVDD.n2470 VSS 0.451316f
C19927 DVDD.n2471 VSS 0.861315f
C19928 DVDD.n2472 VSS 0.225658f
C19929 DVDD.n2473 VSS 0.726238f
C19930 DVDD.n2474 VSS 0.408409f
C19931 DVDD.n2486 VSS 0.127013f
C19932 DVDD.n2488 VSS 0.127013f
C19933 DVDD.n2489 VSS 0.402053f
C19934 DVDD.n2490 VSS 0.066735f
C19935 DVDD.n2491 VSS 0.066735f
C19936 DVDD.n2492 VSS 0.066735f
C19937 DVDD.n2493 VSS 0.066735f
C19938 DVDD.n2494 VSS 0.066735f
C19939 DVDD.n2495 VSS 0.066735f
C19940 DVDD.n2496 VSS 0.066735f
C19941 DVDD.n2497 VSS 0.066735f
C19942 DVDD.n2498 VSS 0.066735f
C19943 DVDD.n2499 VSS 0.066735f
C19944 DVDD.n2500 VSS 0.066735f
C19945 DVDD.n2501 VSS 0.451316f
C19946 DVDD.n2502 VSS 0.451316f
C19947 DVDD.n2503 VSS 0.451316f
C19948 DVDD.n2504 VSS 0.360735f
C19949 DVDD.n2505 VSS 0.451316f
C19950 DVDD.n2506 VSS 3.15709f
C19951 DVDD.n2507 VSS 0.451316f
C19952 DVDD.n2508 VSS 0.225658f
C19953 DVDD.n2521 VSS 0.225658f
C19954 DVDD.n2522 VSS 0.225658f
C19955 DVDD.n2523 VSS 2.66633f
C19956 DVDD.n2524 VSS 0.066735f
C19957 DVDD.n2525 VSS 0.066735f
C19958 DVDD.n2526 VSS 0.066735f
C19959 DVDD.n2527 VSS 0.066735f
C19960 DVDD.n2528 VSS 0.033368f
C19961 DVDD.n2529 VSS 0.033368f
C19962 DVDD.n2530 VSS 0.033368f
C19963 DVDD.n2531 VSS 0.033368f
C19964 DVDD.n2532 VSS 0.033368f
C19965 DVDD.n2533 VSS 0.033368f
C19966 DVDD.n2534 VSS 0.033368f
C19967 DVDD.n2535 VSS 0.033368f
C19968 DVDD.n2536 VSS 0.197054f
C19969 DVDD.n2537 VSS 0.033368f
C19970 DVDD.n2538 VSS 0.033368f
C19971 DVDD.n2539 VSS 0.033368f
C19972 DVDD.n2540 VSS 0.033368f
C19973 DVDD.n2541 VSS 0.033368f
C19974 DVDD.n2542 VSS 0.033368f
C19975 DVDD.n2543 VSS 0.033368f
C19976 DVDD.n2545 VSS 0.047092f
C19977 DVDD.n2547 VSS 0.066735f
C19978 DVDD.n2549 VSS 0.066735f
C19979 DVDD.n2550 VSS 0.930088f
C19980 DVDD.n2551 VSS 3.15709f
C19981 DVDD.n2552 VSS 0.451316f
C19982 DVDD.n2553 VSS 0.451316f
C19983 DVDD.n2554 VSS 0.451316f
C19984 DVDD.n2555 VSS 0.451316f
C19985 DVDD.n2556 VSS 0.451316f
C19986 DVDD.n2557 VSS 0.451316f
C19987 DVDD.n2558 VSS 0.451316f
C19988 DVDD.n2559 VSS 0.451316f
C19989 DVDD.n2560 VSS 0.451316f
C19990 DVDD.n2561 VSS 0.066735f
C19991 DVDD.n2562 VSS 0.066735f
C19992 DVDD.n2563 VSS 0.066735f
C19993 DVDD.n2564 VSS 0.066735f
C19994 DVDD.n2565 VSS 0.066735f
C19995 DVDD.n2566 VSS 0.066735f
C19996 DVDD.n2567 VSS 0.066735f
C19997 DVDD.n2568 VSS 0.066735f
C19998 DVDD.n2569 VSS 0.066735f
C19999 DVDD.n2570 VSS 0.066735f
C20000 DVDD.n2571 VSS 0.066735f
C20001 DVDD.n2572 VSS 0.127013f
C20002 DVDD.n2573 VSS 0.197054f
C20003 DVDD.n2574 VSS 0.066735f
C20004 DVDD.n2575 VSS 0.066735f
C20005 DVDD.n2576 VSS 0.066735f
C20006 DVDD.n2577 VSS 0.066735f
C20007 DVDD.n2578 VSS 0.066735f
C20008 DVDD.n2579 VSS 0.066735f
C20009 DVDD.n2580 VSS 0.066735f
C20010 DVDD.n2581 VSS 0.066735f
C20011 DVDD.n2582 VSS 0.066735f
C20012 DVDD.n2583 VSS 0.066735f
C20013 DVDD.n2584 VSS 0.066735f
C20014 DVDD.n2597 VSS 0.149379f
C20015 DVDD.n2609 VSS 0.225658f
C20016 DVDD.n2610 VSS 0.197054f
C20017 DVDD.n2611 VSS 0.451316f
C20018 DVDD.n2612 VSS 0.451316f
C20019 DVDD.n2613 VSS 0.451316f
C20020 DVDD.n2614 VSS 0.301937f
C20021 DVDD.n2615 VSS 0.543486f
C20022 DVDD.n2616 VSS 0.375037f
C20023 DVDD.n2617 VSS 0.451316f
C20024 DVDD.n2618 VSS 0.451316f
C20025 DVDD.n2619 VSS 0.451316f
C20026 DVDD.n2620 VSS 0.451316f
C20027 DVDD.n2621 VSS 0.451316f
C20028 DVDD.n2622 VSS 0.451316f
C20029 DVDD.n2623 VSS 0.451316f
C20030 DVDD.n2624 VSS 0.451316f
C20031 DVDD.n2625 VSS 0.451316f
C20032 DVDD.n2626 VSS 0.451316f
C20033 DVDD.n2627 VSS 0.451316f
C20034 DVDD.n2628 VSS 0.451316f
C20035 DVDD.n2629 VSS 0.451316f
C20036 DVDD.n2630 VSS 0.029062f
C20037 DVDD.n2631 VSS 0.029062f
C20038 DVDD.n2632 VSS 0.029062f
C20039 DVDD.n2633 VSS 0.029062f
C20040 DVDD.n2634 VSS 0.029062f
C20041 DVDD.n2635 VSS 0.029062f
C20042 DVDD.n2636 VSS 0.029062f
C20043 DVDD.n2637 VSS 0.029062f
C20044 DVDD.n2638 VSS 0.197054f
C20045 DVDD.n2642 VSS 0.057317f
C20046 DVDD.n2643 VSS 0.029062f
C20047 DVDD.n2644 VSS 0.029062f
C20048 DVDD.n2645 VSS 0.029062f
C20049 DVDD.n2646 VSS 0.029062f
C20050 DVDD.n2647 VSS 0.029062f
C20051 DVDD.n2648 VSS 0.029062f
C20052 DVDD.n2649 VSS 0.033368f
C20053 DVDD.n2650 VSS 0.114418f
C20054 DVDD.n2651 VSS 0.033368f
C20055 DVDD.n2652 VSS 0.124509f
C20056 DVDD.n2653 VSS 0.124509f
C20057 DVDD.n2654 VSS 0.114418f
C20058 DVDD.n2655 VSS 0.056779f
C20059 DVDD.n2656 VSS 0.225658f
C20060 DVDD.n2657 VSS 0.225658f
C20061 DVDD.n2658 VSS 0.033368f
C20062 DVDD.n2659 VSS 0.225658f
C20063 DVDD.n2660 VSS 0.197054f
C20064 DVDD.n2661 VSS 0.029062f
C20065 DVDD.n2662 VSS 0.029062f
C20066 DVDD.n2663 VSS 0.029062f
C20067 DVDD.n2664 VSS 0.029062f
C20068 DVDD.n2665 VSS 0.058393f
C20069 DVDD.n2666 VSS 0.066735f
C20070 DVDD.n2667 VSS 0.066735f
C20071 DVDD.n2668 VSS 0.029062f
C20072 DVDD.n2669 VSS 0.029062f
C20073 DVDD.n2670 VSS 0.029062f
C20074 DVDD.n2671 VSS 0.029062f
C20075 DVDD.n2672 VSS 0.360735f
C20076 DVDD.n2673 VSS 0.029062f
C20077 DVDD.n2674 VSS 0.029062f
C20078 DVDD.n2675 VSS 0.033368f
C20079 DVDD.n2676 VSS 0.114418f
C20080 DVDD.n2677 VSS 0.114418f
C20081 DVDD.n2678 VSS 0.033368f
C20082 DVDD.n2679 VSS 0.114418f
C20083 DVDD.n2680 VSS 0.033368f
C20084 DVDD.n2681 VSS 0.114418f
C20085 DVDD.n2682 VSS 0.114418f
C20086 DVDD.n2683 VSS 0.031484f
C20087 DVDD.n2684 VSS 0.030946f
C20088 DVDD.n2685 VSS 0.114418f
C20089 DVDD.n2686 VSS 0.033368f
C20090 DVDD.n2687 VSS 0.114418f
C20091 DVDD.n2688 VSS 0.033368f
C20092 DVDD.n2689 VSS 0.114418f
C20093 DVDD.n2690 VSS 0.033368f
C20094 DVDD.n2691 VSS 0.114418f
C20095 DVDD.n2692 VSS 0.033368f
C20096 DVDD.n2693 VSS 0.114418f
C20097 DVDD.n2694 VSS 0.033368f
C20098 DVDD.n2695 VSS 0.114418f
C20099 DVDD.n2696 VSS 0.033368f
C20100 DVDD.n2697 VSS 0.114418f
C20101 DVDD.n2698 VSS 0.114418f
C20102 DVDD.n2699 VSS 0.030408f
C20103 DVDD.n2700 VSS 0.032022f
C20104 DVDD.n2701 VSS 0.114418f
C20105 DVDD.n2702 VSS 0.033368f
C20106 DVDD.n2703 VSS 0.114418f
C20107 DVDD.n2704 VSS 0.033368f
C20108 DVDD.n2705 VSS 0.114418f
C20109 DVDD.n2706 VSS 0.114418f
C20110 DVDD.n2707 VSS 0.046553f
C20111 DVDD.n2708 VSS 0.058124f
C20112 DVDD.n2709 VSS 0.047092f
C20113 DVDD.n2710 VSS 0.114418f
C20114 DVDD.n2711 VSS 0.033368f
C20115 DVDD.n2712 VSS 0.114418f
C20116 DVDD.n2713 VSS 0.033368f
C20117 DVDD.n2714 VSS 0.114418f
C20118 DVDD.n2715 VSS 0.114418f
C20119 DVDD.n2716 VSS 0.031484f
C20120 DVDD.n2717 VSS 0.030946f
C20121 DVDD.n2718 VSS 0.114418f
C20122 DVDD.n2719 VSS 0.033368f
C20123 DVDD.n2720 VSS 0.114418f
C20124 DVDD.n2721 VSS 0.114418f
C20125 DVDD.n2722 VSS 0.033368f
C20126 DVDD.n2723 VSS 0.029062f
C20127 DVDD.n2726 VSS 0.066735f
C20128 DVDD.n2729 VSS 0.066735f
C20129 DVDD.n2732 VSS 0.066735f
C20130 DVDD.n2733 VSS 0.029062f
C20131 DVDD.n2734 VSS 0.029062f
C20132 DVDD.n2735 VSS 0.029062f
C20133 DVDD.n2736 VSS 0.029062f
C20134 DVDD.n2737 VSS 0.044401f
C20135 DVDD.n2738 VSS 0.114418f
C20136 DVDD.n2739 VSS 0.124509f
C20137 DVDD.n2740 VSS 0.124509f
C20138 DVDD.n2741 VSS 0.114418f
C20139 DVDD.n2742 VSS 0.054088f
C20140 DVDD.n2743 VSS 0.120351f
C20141 DVDD.n2744 VSS 0.058124f
C20142 DVDD.n2745 VSS 0.114418f
C20143 DVDD.n2746 VSS 0.058124f
C20144 DVDD.n2747 VSS 0.114418f
C20145 DVDD.n2748 VSS 0.058124f
C20146 DVDD.n2749 VSS 0.114418f
C20147 DVDD.n2750 VSS 0.058124f
C20148 DVDD.n2751 VSS 0.114418f
C20149 DVDD.n2752 VSS 0.058124f
C20150 DVDD.n2753 VSS 0.058124f
C20151 DVDD.n2754 VSS 0.114418f
C20152 DVDD.n2755 VSS 0.114418f
C20153 DVDD.n2756 VSS 0.114418f
C20154 DVDD.n2757 VSS 0.058124f
C20155 DVDD.n2758 VSS 0.058124f
C20156 DVDD.n2759 VSS 0.058124f
C20157 DVDD.n2760 VSS 0.114418f
C20158 DVDD.n2761 VSS 0.114418f
C20159 DVDD.n2762 VSS 0.114418f
C20160 DVDD.n2763 VSS 0.058124f
C20161 DVDD.n2764 VSS 0.058124f
C20162 DVDD.n2765 VSS 0.058124f
C20163 DVDD.n2766 VSS 0.114418f
C20164 DVDD.n2767 VSS 0.114418f
C20165 DVDD.n2768 VSS 0.114418f
C20166 DVDD.n2769 VSS 0.058124f
C20167 DVDD.n2770 VSS 0.058124f
C20168 DVDD.n2771 VSS 0.058124f
C20169 DVDD.n2772 VSS 0.114418f
C20170 DVDD.n2773 VSS 0.114418f
C20171 DVDD.n2774 VSS 0.114418f
C20172 DVDD.n2775 VSS 0.058124f
C20173 DVDD.n2776 VSS 0.045477f
C20174 DVDD.n2777 VSS 0.108485f
C20175 DVDD.n2778 VSS 0.026274f
C20176 DVDD.n2779 VSS 0.060175f
C20177 DVDD.n2780 VSS 0.060175f
C20178 DVDD.n2781 VSS 0.060175f
C20179 DVDD.n2782 VSS 0.030088f
C20180 DVDD.n2783 VSS 0.027333f
C20181 DVDD.n2785 VSS 0.093653f
C20182 DVDD.n2786 VSS 0.172475f
C20183 DVDD.n2787 VSS 0.154253f
C20184 DVDD.n2788 VSS 0.228836f
C20185 DVDD.n2789 VSS 0.060175f
C20186 DVDD.n2790 VSS 0.060175f
C20187 DVDD.n2791 VSS 0.026274f
C20188 DVDD.n2792 VSS 0.033368f
C20189 DVDD.n2793 VSS 0.030088f
C20190 DVDD.n2794 VSS 0.060175f
C20191 DVDD.n2795 VSS 0.026274f
C20192 DVDD.n2796 VSS 0.02691f
C20193 DVDD.n2797 VSS 0.043862f
C20194 DVDD.n2798 VSS 0.029062f
C20195 DVDD.n2799 VSS 0.114418f
C20196 DVDD.n2800 VSS 0.124509f
C20197 DVDD.n2801 VSS 0.124509f
C20198 DVDD.n2802 VSS 0.114418f
C20199 DVDD.n2803 VSS 0.054626f
C20200 DVDD.n2804 VSS 0.225658f
C20201 DVDD.n2805 VSS 0.225658f
C20202 DVDD.n2806 VSS 0.033368f
C20203 DVDD.n2807 VSS 0.225658f
C20204 DVDD.n2808 VSS 0.197054f
C20205 DVDD.n2809 VSS 0.066735f
C20206 DVDD.n2810 VSS 0.029062f
C20207 DVDD.n2811 VSS 0.029062f
C20208 DVDD.n2812 VSS 0.029062f
C20209 DVDD.n2813 VSS 0.029062f
C20210 DVDD.n2814 VSS 0.029062f
C20211 DVDD.n2815 VSS 0.029062f
C20212 DVDD.n2816 VSS 0.029062f
C20213 DVDD.n2817 VSS 0.029062f
C20214 DVDD.n2818 VSS 0.029062f
C20215 DVDD.n2819 VSS 0.029062f
C20216 DVDD.n2820 VSS 0.360735f
C20217 DVDD.n2821 VSS 0.029062f
C20218 DVDD.n2822 VSS 0.029062f
C20219 DVDD.n2823 VSS 0.029062f
C20220 DVDD.n2824 VSS 0.029062f
C20221 DVDD.n2825 VSS 0.029062f
C20222 DVDD.n2826 VSS 0.029062f
C20223 DVDD.n2827 VSS 0.029062f
C20224 DVDD.n2828 VSS 0.029062f
C20225 DVDD.n2829 VSS 0.033368f
C20226 DVDD.n2830 VSS 0.114418f
C20227 DVDD.n2831 VSS 0.114418f
C20228 DVDD.n2832 VSS 0.058124f
C20229 DVDD.n2833 VSS 0.051397f
C20230 DVDD.n2834 VSS 0.114418f
C20231 DVDD.n2835 VSS 0.033368f
C20232 DVDD.n2836 VSS 0.114418f
C20233 DVDD.n2837 VSS 0.114418f
C20234 DVDD.n2838 VSS 0.031484f
C20235 DVDD.n2839 VSS 0.030946f
C20236 DVDD.n2840 VSS 0.114418f
C20237 DVDD.n2841 VSS 0.033368f
C20238 DVDD.n2842 VSS 0.114418f
C20239 DVDD.n2843 VSS 0.033368f
C20240 DVDD.n2844 VSS 0.114418f
C20241 DVDD.n2845 VSS 0.033368f
C20242 DVDD.n2846 VSS 0.114418f
C20243 DVDD.n2847 VSS 0.033368f
C20244 DVDD.n2848 VSS 0.114418f
C20245 DVDD.n2849 VSS 0.033368f
C20246 DVDD.n2850 VSS 0.114418f
C20247 DVDD.n2851 VSS 0.033368f
C20248 DVDD.n2852 VSS 0.114418f
C20249 DVDD.n2853 VSS 0.114418f
C20250 DVDD.n2854 VSS 0.030408f
C20251 DVDD.n2855 VSS 0.032022f
C20252 DVDD.n2856 VSS 0.114418f
C20253 DVDD.n2857 VSS 0.033368f
C20254 DVDD.n2858 VSS 0.114418f
C20255 DVDD.n2859 VSS 0.033368f
C20256 DVDD.n2860 VSS 0.114418f
C20257 DVDD.n2861 VSS 0.033368f
C20258 DVDD.n2862 VSS 0.114418f
C20259 DVDD.n2863 VSS 0.033368f
C20260 DVDD.n2864 VSS 0.114418f
C20261 DVDD.n2865 VSS 0.033368f
C20262 DVDD.n2866 VSS 0.114418f
C20263 DVDD.n2867 VSS 0.033368f
C20264 DVDD.n2868 VSS 0.114418f
C20265 DVDD.n2869 VSS 0.114418f
C20266 DVDD.n2870 VSS 0.029331f
C20267 DVDD.n2871 VSS 0.033099f
C20268 DVDD.n2872 VSS 0.114418f
C20269 DVDD.n2873 VSS 0.114418f
C20270 DVDD.n2874 VSS 0.033368f
C20271 DVDD.n2875 VSS 0.029062f
C20272 DVDD.n2878 VSS 0.066735f
C20273 DVDD.n2879 VSS 0.058124f
C20274 DVDD.n2880 VSS 0.114418f
C20275 DVDD.n2881 VSS 0.124509f
C20276 DVDD.n2882 VSS 0.124509f
C20277 DVDD.n2883 VSS 0.114418f
C20278 DVDD.n2884 VSS 0.058124f
C20279 DVDD.n2885 VSS 0.114418f
C20280 DVDD.n2886 VSS 0.124509f
C20281 DVDD.n2887 VSS 0.124509f
C20282 DVDD.n2888 VSS 0.114418f
C20283 DVDD.n2889 VSS 0.04763f
C20284 DVDD.n2890 VSS 0.026274f
C20285 DVDD.n2891 VSS 0.030088f
C20286 DVDD.n2892 VSS 0.033368f
C20287 DVDD.n2893 VSS 0.197054f
C20288 DVDD.n2894 VSS 0.197054f
C20289 DVDD.n2895 VSS 0.033368f
C20290 DVDD.n2896 VSS 0.066735f
C20291 DVDD.n2897 VSS 0.066735f
C20292 DVDD.n2898 VSS 0.197054f
C20293 DVDD.n2899 VSS 0.033368f
C20294 DVDD.n2900 VSS 0.030088f
C20295 DVDD.n2901 VSS 0.032022f
C20296 DVDD.n2902 VSS 0.114418f
C20297 DVDD.n2903 VSS 0.114418f
C20298 DVDD.n2904 VSS 0.029062f
C20299 DVDD.n2905 VSS 0.033368f
C20300 DVDD.n2906 VSS 0.201821f
C20301 DVDD.n2907 VSS 0.026274f
C20302 DVDD.n2908 VSS 0.060175f
C20303 DVDD.n2909 VSS 0.060175f
C20304 DVDD.n2910 VSS 0.026274f
C20305 DVDD.n2911 VSS 0.060175f
C20306 DVDD.n2912 VSS 0.030088f
C20307 DVDD.n2913 VSS 0.026274f
C20308 DVDD.n2914 VSS 0.060175f
C20309 DVDD.n2915 VSS 0.173937f
C20310 DVDD.n2916 VSS 0.061117f
C20311 DVDD.n2917 VSS 0.058124f
C20312 DVDD.n2918 VSS 0.114418f
C20313 DVDD.n2919 VSS 0.058124f
C20314 DVDD.n2920 VSS 0.114418f
C20315 DVDD.n2921 VSS 0.058124f
C20316 DVDD.n2922 VSS 0.114418f
C20317 DVDD.n2923 VSS 0.058124f
C20318 DVDD.n2924 VSS 0.114418f
C20319 DVDD.n2925 VSS 0.058124f
C20320 DVDD.n2926 VSS 0.114418f
C20321 DVDD.n2927 VSS 0.058124f
C20322 DVDD.n2928 VSS 0.058124f
C20323 DVDD.n2929 VSS 0.114418f
C20324 DVDD.n2930 VSS 0.114418f
C20325 DVDD.n2931 VSS 0.114418f
C20326 DVDD.n2932 VSS 0.058124f
C20327 DVDD.n2933 VSS 0.058124f
C20328 DVDD.n2934 VSS 0.058124f
C20329 DVDD.n2935 VSS 0.114418f
C20330 DVDD.n2936 VSS 0.114418f
C20331 DVDD.n2937 VSS 0.114418f
C20332 DVDD.n2938 VSS 0.058124f
C20333 DVDD.n2939 VSS 0.058124f
C20334 DVDD.n2940 VSS 0.058124f
C20335 DVDD.n2941 VSS 0.114418f
C20336 DVDD.n2942 VSS 0.114418f
C20337 DVDD.n2943 VSS 0.114418f
C20338 DVDD.n2944 VSS 0.058124f
C20339 DVDD.n2945 VSS 0.058124f
C20340 DVDD.n2946 VSS 0.058124f
C20341 DVDD.n2947 VSS 0.114418f
C20342 DVDD.n2948 VSS 0.114418f
C20343 DVDD.n2949 VSS 0.114418f
C20344 DVDD.n2950 VSS 0.058124f
C20345 DVDD.n2951 VSS 0.058124f
C20346 DVDD.n2952 VSS 0.058124f
C20347 DVDD.n2953 VSS 0.114418f
C20348 DVDD.n2954 VSS 0.114418f
C20349 DVDD.n2955 VSS 0.114418f
C20350 DVDD.n2956 VSS 0.046553f
C20351 DVDD.n2957 VSS 0.455731f
C20352 DVDD.n2958 VSS 0.033368f
C20353 DVDD.n2959 VSS 0.066735f
C20354 DVDD.n2961 VSS 0.149379f
C20355 DVDD.n2962 VSS 0.225658f
C20356 DVDD.n2963 VSS 0.402053f
C20357 DVDD.n2964 VSS 0.066735f
C20358 DVDD.n2965 VSS 0.066735f
C20359 DVDD.n2966 VSS 0.066735f
C20360 DVDD.n2967 VSS 0.066735f
C20361 DVDD.n2968 VSS 0.066735f
C20362 DVDD.n2969 VSS 0.066735f
C20363 DVDD.n2970 VSS 0.066735f
C20364 DVDD.n2971 VSS 0.066735f
C20365 DVDD.n2972 VSS 0.066735f
C20366 DVDD.n2973 VSS 0.066735f
C20367 DVDD.n2974 VSS 0.066735f
C20368 DVDD.n2975 VSS 0.197054f
C20369 DVDD.n2977 VSS 0.066735f
C20370 DVDD.n2979 VSS 0.066735f
C20371 DVDD.n2981 VSS 0.066735f
C20372 DVDD.n2983 VSS 0.066735f
C20373 DVDD.n2985 VSS 0.066735f
C20374 DVDD.n2987 VSS 0.066735f
C20375 DVDD.n2989 VSS 0.066735f
C20376 DVDD.n2991 VSS 0.066735f
C20377 DVDD.n2993 VSS 0.066735f
C20378 DVDD.n2995 VSS 0.066735f
C20379 DVDD.n2997 VSS 0.066735f
C20380 DVDD.n3000 VSS 0.079669f
C20381 DVDD.n3001 VSS 0.120351f
C20382 DVDD.n3002 VSS 0.214428f
C20383 DVDD.n3003 VSS 0.066735f
C20384 DVDD.n3004 VSS 0.066735f
C20385 DVDD.n3005 VSS 0.066735f
C20386 DVDD.n3006 VSS 0.066735f
C20387 DVDD.n3007 VSS 0.066735f
C20388 DVDD.n3008 VSS 0.105095f
C20389 DVDD.n3010 VSS 0.066735f
C20390 DVDD.n3012 VSS 0.066735f
C20391 DVDD.n3014 VSS 0.066735f
C20392 DVDD.n3016 VSS 0.066735f
C20393 DVDD.n3022 VSS 0.120351f
C20394 DVDD.n3024 VSS 0.149379f
C20395 DVDD.n3025 VSS 0.225658f
C20396 DVDD.n3026 VSS 0.402053f
C20397 DVDD.n3027 VSS 0.066735f
C20398 DVDD.n3028 VSS 0.066735f
C20399 DVDD.n3029 VSS 0.066735f
C20400 DVDD.n3030 VSS 0.066735f
C20401 DVDD.n3031 VSS 0.066735f
C20402 DVDD.n3032 VSS 0.066735f
C20403 DVDD.n3033 VSS 0.066735f
C20404 DVDD.n3034 VSS 0.066735f
C20405 DVDD.n3035 VSS 0.066735f
C20406 DVDD.n3036 VSS 0.066735f
C20407 DVDD.n3037 VSS 0.066735f
C20408 DVDD.n3038 VSS 0.197054f
C20409 DVDD.n3040 VSS 0.066735f
C20410 DVDD.n3042 VSS 0.066735f
C20411 DVDD.n3044 VSS 0.066735f
C20412 DVDD.n3046 VSS 0.066735f
C20413 DVDD.n3048 VSS 0.066735f
C20414 DVDD.n3050 VSS 0.066735f
C20415 DVDD.n3052 VSS 0.066735f
C20416 DVDD.n3054 VSS 0.066735f
C20417 DVDD.n3056 VSS 0.066735f
C20418 DVDD.n3058 VSS 0.066735f
C20419 DVDD.n3060 VSS 0.066735f
C20420 DVDD.n3061 VSS 0.451316f
C20421 DVDD.n3062 VSS 0.451316f
C20422 DVDD.n3063 VSS 0.451316f
C20423 DVDD.n3064 VSS 0.451316f
C20424 DVDD.n3065 VSS 0.451316f
C20425 DVDD.n3066 VSS 0.451316f
C20426 DVDD.n3067 VSS 0.451316f
C20427 DVDD.n3068 VSS 0.451316f
C20428 DVDD.n3069 VSS 0.451316f
C20429 DVDD.n3070 VSS 0.451316f
C20430 DVDD.n3071 VSS 0.451316f
C20431 DVDD.n3072 VSS 0.451316f
C20432 DVDD.n3073 VSS 0.451316f
C20433 DVDD.n3074 VSS 0.451316f
C20434 DVDD.n3075 VSS 0.451316f
C20435 DVDD.n3076 VSS 0.451316f
C20436 DVDD.n3077 VSS 0.451316f
C20437 DVDD.n3078 VSS 0.451316f
C20438 DVDD.n3079 VSS 0.451316f
C20439 DVDD.n3080 VSS 0.451316f
C20440 DVDD.n3081 VSS 0.451316f
C20441 DVDD.n3082 VSS 0.451316f
C20442 DVDD.n3083 VSS 0.451316f
C20443 DVDD.n3084 VSS 0.451316f
C20444 DVDD.n3085 VSS 0.451316f
C20445 DVDD.n3086 VSS 0.451316f
C20446 DVDD.n3087 VSS 0.451316f
C20447 DVDD.n3088 VSS 0.451316f
C20448 DVDD.n3089 VSS 0.451316f
C20449 DVDD.n3090 VSS 0.451316f
C20450 DVDD.n3091 VSS 0.451316f
C20451 DVDD.n3092 VSS 0.451316f
C20452 DVDD.n3093 VSS 0.451316f
C20453 DVDD.n3094 VSS 0.289224f
C20454 DVDD.n3095 VSS 0.387751f
C20455 DVDD.n3096 VSS 0.451316f
C20456 DVDD.n3097 VSS 0.029062f
C20457 DVDD.n3098 VSS 0.029062f
C20458 DVDD.n3099 VSS 0.029062f
C20459 DVDD.n3100 VSS 0.029062f
C20460 DVDD.n3101 VSS 0.066735f
C20461 DVDD.n3102 VSS 0.066735f
C20462 DVDD.n3103 VSS 0.066735f
C20463 DVDD.n3104 VSS 0.029062f
C20464 DVDD.n3105 VSS 0.029062f
C20465 DVDD.n3106 VSS 0.029062f
C20466 DVDD.n3107 VSS 0.029062f
C20467 DVDD.n3108 VSS 0.029062f
C20468 DVDD.n3109 VSS 0.197054f
C20469 DVDD.n3110 VSS 0.029062f
C20470 DVDD.n3111 VSS 0.029062f
C20471 DVDD.n3112 VSS 0.029062f
C20472 DVDD.n3113 VSS 0.029062f
C20473 DVDD.n3114 VSS 0.058393f
C20474 DVDD.n3115 VSS 0.066735f
C20475 DVDD.n3116 VSS 0.066735f
C20476 DVDD.n3117 VSS 0.056779f
C20477 DVDD.n3118 VSS 0.029062f
C20478 DVDD.n3119 VSS 0.029062f
C20479 DVDD.n3120 VSS 0.029062f
C20480 DVDD.n3121 VSS 0.033368f
C20481 DVDD.n3122 VSS 0.225658f
C20482 DVDD.n3123 VSS 0.058124f
C20483 DVDD.n3124 VSS 0.114418f
C20484 DVDD.n3125 VSS 0.033368f
C20485 DVDD.n3126 VSS 0.114418f
C20486 DVDD.n3127 VSS 0.114418f
C20487 DVDD.n3128 VSS 0.031484f
C20488 DVDD.n3129 VSS 0.030946f
C20489 DVDD.n3130 VSS 0.114418f
C20490 DVDD.n3131 VSS 0.033368f
C20491 DVDD.n3132 VSS 0.114418f
C20492 DVDD.n3133 VSS 0.033368f
C20493 DVDD.n3134 VSS 0.114418f
C20494 DVDD.n3135 VSS 0.033368f
C20495 DVDD.n3136 VSS 0.114418f
C20496 DVDD.n3137 VSS 0.033368f
C20497 DVDD.n3138 VSS 0.114418f
C20498 DVDD.n3139 VSS 0.033368f
C20499 DVDD.n3140 VSS 0.15585f
C20500 DVDD.t13 VSS 5.27557f
C20501 DVDD.n3142 VSS 0.033368f
C20502 DVDD.n3143 VSS 0.15585f
C20503 DVDD.n3144 VSS 0.033368f
C20504 DVDD.n3145 VSS 0.114418f
C20505 DVDD.n3146 VSS 0.033368f
C20506 DVDD.n3147 VSS 0.114418f
C20507 DVDD.n3148 VSS 0.033368f
C20508 DVDD.n3149 VSS 0.114418f
C20509 DVDD.n3150 VSS 0.033368f
C20510 DVDD.n3151 VSS 0.114418f
C20511 DVDD.n3152 VSS 0.114418f
C20512 DVDD.n3153 VSS 0.031484f
C20513 DVDD.n3154 VSS 0.030946f
C20514 DVDD.n3155 VSS 0.114418f
C20515 DVDD.n3156 VSS 0.033368f
C20516 DVDD.n3157 VSS 0.114418f
C20517 DVDD.n3158 VSS 0.033368f
C20518 DVDD.n3159 VSS 0.114418f
C20519 DVDD.n3160 VSS 0.033368f
C20520 DVDD.n3161 VSS 0.114418f
C20521 DVDD.n3162 VSS 0.033368f
C20522 DVDD.n3163 VSS 0.114418f
C20523 DVDD.n3164 VSS 0.033368f
C20524 DVDD.n3165 VSS 0.114418f
C20525 DVDD.n3166 VSS 0.033368f
C20526 DVDD.n3167 VSS 0.114418f
C20527 DVDD.n3168 VSS 0.114418f
C20528 DVDD.n3169 VSS 0.030408f
C20529 DVDD.n3170 VSS 0.032022f
C20530 DVDD.n3171 VSS 0.114418f
C20531 DVDD.n3172 VSS 0.033368f
C20532 DVDD.n3173 VSS 0.114418f
C20533 DVDD.n3174 VSS 0.033368f
C20534 DVDD.n3175 VSS 0.114418f
C20535 DVDD.n3176 VSS 0.046553f
C20536 DVDD.n3177 VSS 0.114418f
C20537 DVDD.n3178 VSS 0.114418f
C20538 DVDD.n3179 VSS 0.114418f
C20539 DVDD.n3180 VSS 0.047092f
C20540 DVDD.n3184 VSS 0.225658f
C20541 DVDD.n3185 VSS 0.197054f
C20542 DVDD.n3186 VSS 0.451316f
C20543 DVDD.n3187 VSS 0.451316f
C20544 DVDD.n3188 VSS 0.451316f
C20545 DVDD.n3189 VSS 0.197054f
C20546 DVDD.n3190 VSS 0.451316f
C20547 DVDD.n3191 VSS 0.451316f
C20548 DVDD.n3192 VSS 0.451316f
C20549 DVDD.n3193 VSS 0.451316f
C20550 DVDD.n3194 VSS 0.451316f
C20551 DVDD.n3195 VSS 0.451316f
C20552 DVDD.n3196 VSS 0.451316f
C20553 DVDD.n3197 VSS 0.451316f
C20554 DVDD.n3198 VSS 0.451316f
C20555 DVDD.n3199 VSS 0.451316f
C20556 DVDD.n3200 VSS 0.451316f
C20557 DVDD.n3201 VSS 0.451316f
C20558 DVDD.n3202 VSS 0.451316f
C20559 DVDD.n3203 VSS 0.451316f
C20560 DVDD.n3204 VSS 0.451316f
C20561 DVDD.n3205 VSS 0.451316f
C20562 DVDD.n3206 VSS 0.451316f
C20563 DVDD.n3207 VSS 0.451316f
C20564 DVDD.n3208 VSS 0.451316f
C20565 DVDD.n3209 VSS 0.451316f
C20566 DVDD.n3210 VSS 0.451316f
C20567 DVDD.n3211 VSS 0.451316f
C20568 DVDD.n3212 VSS 0.451316f
C20569 DVDD.n3213 VSS 0.451316f
C20570 DVDD.n3214 VSS 0.451316f
C20571 DVDD.n3215 VSS 0.029062f
C20572 DVDD.n3216 VSS 0.029062f
C20573 DVDD.n3217 VSS 0.029062f
C20574 DVDD.n3218 VSS 0.029062f
C20575 DVDD.n3219 VSS 0.029062f
C20576 DVDD.n3220 VSS 0.029062f
C20577 DVDD.n3224 VSS 0.029062f
C20578 DVDD.n3225 VSS 0.029062f
C20579 DVDD.n3226 VSS 0.029062f
C20580 DVDD.n3227 VSS 0.197054f
C20581 DVDD.n3228 VSS 0.029062f
C20582 DVDD.n3229 VSS 0.029062f
C20583 DVDD.n3230 VSS 0.056779f
C20584 DVDD.n3231 VSS 0.029062f
C20585 DVDD.n3232 VSS 0.029062f
C20586 DVDD.n3233 VSS 0.029062f
C20587 DVDD.n3234 VSS 0.029062f
C20588 DVDD.n3235 VSS 0.029062f
C20589 DVDD.n3236 VSS 0.033368f
C20590 DVDD.n3237 VSS 0.225658f
C20591 DVDD.n3238 VSS 0.225658f
C20592 DVDD.n3239 VSS 0.031484f
C20593 DVDD.n3240 VSS 0.114418f
C20594 DVDD.n3241 VSS 0.114418f
C20595 DVDD.n3242 VSS 0.033368f
C20596 DVDD.n3243 VSS 0.114418f
C20597 DVDD.n3244 VSS 0.033368f
C20598 DVDD.n3245 VSS 0.114418f
C20599 DVDD.n3246 VSS 0.033368f
C20600 DVDD.n3247 VSS 0.114418f
C20601 DVDD.n3248 VSS 0.033368f
C20602 DVDD.n3249 VSS 0.15585f
C20603 DVDD.t30 VSS 5.27557f
C20604 DVDD.n3251 VSS 0.033368f
C20605 DVDD.n3252 VSS 0.15585f
C20606 DVDD.n3253 VSS 0.033368f
C20607 DVDD.n3254 VSS 0.114418f
C20608 DVDD.n3255 VSS 0.033368f
C20609 DVDD.n3256 VSS 0.114418f
C20610 DVDD.n3257 VSS 0.033368f
C20611 DVDD.n3258 VSS 0.114418f
C20612 DVDD.n3259 VSS 0.033368f
C20613 DVDD.n3260 VSS 0.114418f
C20614 DVDD.n3261 VSS 0.114418f
C20615 DVDD.n3262 VSS 0.031484f
C20616 DVDD.n3263 VSS 0.030946f
C20617 DVDD.n3264 VSS 0.114418f
C20618 DVDD.n3265 VSS 0.033368f
C20619 DVDD.n3266 VSS 0.114418f
C20620 DVDD.n3267 VSS 0.033368f
C20621 DVDD.n3268 VSS 0.114418f
C20622 DVDD.n3269 VSS 0.033368f
C20623 DVDD.n3270 VSS 0.114418f
C20624 DVDD.n3271 VSS 0.033368f
C20625 DVDD.n3272 VSS 0.114418f
C20626 DVDD.n3273 VSS 0.033368f
C20627 DVDD.n3274 VSS 0.114418f
C20628 DVDD.n3275 VSS 0.033368f
C20629 DVDD.n3276 VSS 0.114418f
C20630 DVDD.n3277 VSS 0.114418f
C20631 DVDD.n3278 VSS 0.030408f
C20632 DVDD.n3279 VSS 0.032022f
C20633 DVDD.n3280 VSS 0.114418f
C20634 DVDD.n3281 VSS 0.033368f
C20635 DVDD.n3282 VSS 0.114418f
C20636 DVDD.n3283 VSS 0.033368f
C20637 DVDD.n3284 VSS 0.114418f
C20638 DVDD.n3285 VSS 0.114418f
C20639 DVDD.n3286 VSS 0.046553f
C20640 DVDD.n3287 VSS 0.058124f
C20641 DVDD.n3288 VSS 0.047092f
C20642 DVDD.n3289 VSS 0.114418f
C20643 DVDD.n3290 VSS 0.033368f
C20644 DVDD.n3291 VSS 0.114418f
C20645 DVDD.n3292 VSS 0.033368f
C20646 DVDD.n3293 VSS 0.114418f
C20647 DVDD.n3294 VSS 0.114418f
C20648 DVDD.n3295 VSS 0.114418f
C20649 DVDD.n3296 VSS 0.030946f
C20650 DVDD.n3297 VSS 0.197054f
C20651 DVDD.n3298 VSS 0.058393f
C20652 DVDD.n3299 VSS 0.066735f
C20653 DVDD.n3300 VSS 0.066735f
C20654 DVDD.n3302 VSS 0.066735f
C20655 DVDD.n3303 VSS 0.066735f
C20656 DVDD.n3305 VSS 0.066735f
C20657 DVDD.n3307 VSS 0.451316f
C20658 DVDD.n3308 VSS 0.451316f
C20659 DVDD.n3309 VSS 0.451316f
C20660 DVDD.n3310 VSS 0.451316f
C20661 DVDD.n3311 VSS 0.451316f
C20662 DVDD.n3312 VSS 0.451316f
C20663 DVDD.n3313 VSS 0.276511f
C20664 DVDD.n3314 VSS 0.451316f
C20665 DVDD.n3315 VSS 0.543486f
C20666 DVDD.n3316 VSS 0.400464f
C20667 DVDD.n3317 VSS 0.451316f
C20668 DVDD.n3318 VSS 0.451316f
C20669 DVDD.n3319 VSS 0.451316f
C20670 DVDD.n3320 VSS 0.451316f
C20671 DVDD.n3321 VSS 0.451316f
C20672 DVDD.n3322 VSS 0.451316f
C20673 DVDD.n3323 VSS 0.451316f
C20674 DVDD.n3324 VSS 0.451316f
C20675 DVDD.n3325 VSS 0.451316f
C20676 DVDD.n3326 VSS 0.451316f
C20677 DVDD.n3327 VSS 0.451316f
C20678 DVDD.n3328 VSS 0.451316f
C20679 DVDD.n3329 VSS 0.451316f
C20680 DVDD.n3330 VSS 0.451316f
C20681 DVDD.n3331 VSS 0.451316f
C20682 DVDD.n3332 VSS 0.029062f
C20683 DVDD.n3333 VSS 0.029062f
C20684 DVDD.n3334 VSS 0.029062f
C20685 DVDD.n3335 VSS 0.029062f
C20686 DVDD.n3336 VSS 0.066735f
C20687 DVDD.n3337 VSS 0.066735f
C20688 DVDD.n3338 VSS 0.066735f
C20689 DVDD.n3339 VSS 0.029062f
C20690 DVDD.n3340 VSS 0.029062f
C20691 DVDD.n3341 VSS 0.029062f
C20692 DVDD.n3342 VSS 0.029062f
C20693 DVDD.n3343 VSS 0.029062f
C20694 DVDD.n3344 VSS 0.197054f
C20695 DVDD.n3345 VSS 0.029062f
C20696 DVDD.n3346 VSS 0.029062f
C20697 DVDD.n3347 VSS 0.029062f
C20698 DVDD.n3348 VSS 0.029062f
C20699 DVDD.n3349 VSS 0.058393f
C20700 DVDD.n3350 VSS 0.066735f
C20701 DVDD.n3351 VSS 0.066735f
C20702 DVDD.n3352 VSS 0.056779f
C20703 DVDD.n3353 VSS 0.029062f
C20704 DVDD.n3354 VSS 0.029062f
C20705 DVDD.n3355 VSS 0.029062f
C20706 DVDD.n3356 VSS 0.033368f
C20707 DVDD.n3357 VSS 0.225658f
C20708 DVDD.n3358 VSS 0.047092f
C20709 DVDD.n3362 VSS 0.225658f
C20710 DVDD.n3363 VSS 0.197054f
C20711 DVDD.n3364 VSS 0.451316f
C20712 DVDD.n3365 VSS 0.451316f
C20713 DVDD.n3366 VSS 0.451316f
C20714 DVDD.n3367 VSS 0.451316f
C20715 DVDD.n3368 VSS 0.451316f
C20716 DVDD.n3369 VSS 0.197054f
C20717 DVDD.n3370 VSS 0.451316f
C20718 DVDD.n3371 VSS 0.451316f
C20719 DVDD.n3372 VSS 0.451316f
C20720 DVDD.n3373 VSS 0.451316f
C20721 DVDD.n3374 VSS 0.451316f
C20722 DVDD.n3375 VSS 0.451316f
C20723 DVDD.n3376 VSS 0.451316f
C20724 DVDD.n3377 VSS 0.451316f
C20725 DVDD.n3378 VSS 0.451316f
C20726 DVDD.n3379 VSS 0.451316f
C20727 DVDD.n3380 VSS 0.451316f
C20728 DVDD.n3381 VSS 0.451316f
C20729 DVDD.n3382 VSS 0.451316f
C20730 DVDD.n3383 VSS 0.451316f
C20731 DVDD.n3384 VSS 0.263798f
C20732 DVDD.n3385 VSS 0.413177f
C20733 DVDD.n3386 VSS 0.451316f
C20734 DVDD.n3387 VSS 0.451316f
C20735 DVDD.n3388 VSS 0.451316f
C20736 DVDD.n3389 VSS 0.451316f
C20737 DVDD.n3390 VSS 0.451316f
C20738 DVDD.n3391 VSS 0.451316f
C20739 DVDD.n3392 VSS 0.451316f
C20740 DVDD.n3393 VSS 0.451316f
C20741 DVDD.n3394 VSS 0.451316f
C20742 DVDD.n3395 VSS 0.451316f
C20743 DVDD.n3396 VSS 0.031397f
C20744 DVDD.n3397 VSS 0.031397f
C20745 DVDD.n3398 VSS 0.031397f
C20746 DVDD.n3399 VSS 0.031397f
C20747 DVDD.n3400 VSS 0.062794f
C20748 DVDD.n3401 VSS 0.062794f
C20749 DVDD.n3402 VSS 0.062794f
C20750 DVDD.n3403 VSS 0.031397f
C20751 DVDD.n3404 VSS 0.031397f
C20752 DVDD.n3405 VSS 0.031397f
C20753 DVDD.n3406 VSS 0.031397f
C20754 DVDD.n3407 VSS 0.031837f
C20755 DVDD.n3408 VSS 0.197054f
C20756 DVDD.n3409 VSS 0.031397f
C20757 DVDD.n3410 VSS 0.031397f
C20758 DVDD.n3411 VSS 0.031397f
C20759 DVDD.n3412 VSS 0.031397f
C20760 DVDD.n3413 VSS 0.031397f
C20761 DVDD.n3414 VSS 0.131369f
C20762 DVDD.n3415 VSS 0.033368f
C20763 DVDD.n3416 VSS 0.15585f
C20764 DVDD.n3417 VSS 0.15585f
C20765 DVDD.n3418 VSS 0.131369f
C20766 DVDD.n3419 VSS 0.041272f
C20767 DVDD.n3420 VSS 0.120351f
C20768 DVDD.n3421 VSS 0.139516f
C20769 DVDD.n3422 VSS 0.048607f
C20770 DVDD.n3423 VSS 0.131369f
C20771 DVDD.n3424 VSS 0.048607f
C20772 DVDD.n3425 VSS 0.131369f
C20773 DVDD.n3426 VSS 0.048607f
C20774 DVDD.n3427 VSS 0.131369f
C20775 DVDD.n3428 VSS 0.048607f
C20776 DVDD.n3429 VSS 0.031397f
C20777 DVDD.n3430 VSS 0.131369f
C20778 DVDD.n3431 VSS 0.031397f
C20779 DVDD.n3432 VSS 0.131369f
C20780 DVDD.n3433 VSS 0.031397f
C20781 DVDD.n3434 VSS 0.131369f
C20782 DVDD.n3435 VSS 0.031397f
C20783 DVDD.n3436 VSS 0.131369f
C20784 DVDD.n3437 VSS 0.031397f
C20785 DVDD.n3438 VSS 0.131369f
C20786 DVDD.n3439 VSS 0.031397f
C20787 DVDD.n3440 VSS 0.131369f
C20788 DVDD.n3441 VSS 0.031397f
C20789 DVDD.n3442 VSS 0.131369f
C20790 DVDD.n3443 VSS 0.035844f
C20791 DVDD.n3444 VSS 0.131369f
C20792 DVDD.n3445 VSS 0.131369f
C20793 DVDD.n3446 VSS 0.131369f
C20794 DVDD.n3447 VSS 0.048607f
C20795 DVDD.n3448 VSS 0.048607f
C20796 DVDD.n3449 VSS 0.048607f
C20797 DVDD.n3450 VSS 0.131369f
C20798 DVDD.n3451 VSS 0.131369f
C20799 DVDD.n3452 VSS 0.131369f
C20800 DVDD.n3453 VSS 0.048607f
C20801 DVDD.n3454 VSS 0.048607f
C20802 DVDD.n3455 VSS 0.048607f
C20803 DVDD.n3456 VSS 0.131369f
C20804 DVDD.n3457 VSS 0.131369f
C20805 DVDD.n3458 VSS 0.131369f
C20806 DVDD.n3459 VSS 0.048607f
C20807 DVDD.n3460 VSS 0.048607f
C20808 DVDD.n3461 VSS 0.048607f
C20809 DVDD.n3462 VSS 0.131369f
C20810 DVDD.n3463 VSS 0.131369f
C20811 DVDD.n3464 VSS 0.131369f
C20812 DVDD.n3465 VSS 0.048607f
C20813 DVDD.n3466 VSS 0.033994f
C20814 DVDD.n3467 VSS 0.088144f
C20815 DVDD.n3468 VSS 0.195782f
C20816 DVDD.n3469 VSS 0.062794f
C20817 DVDD.n3470 VSS 0.062794f
C20818 DVDD.n3471 VSS 0.047855f
C20819 DVDD.n3472 VSS 0.031397f
C20820 DVDD.n3473 VSS 0.105095f
C20821 DVDD.n3474 VSS 0.031698f
C20822 DVDD.n3475 VSS 0.031397f
C20823 DVDD.n3478 VSS 0.062794f
C20824 DVDD.n3481 VSS 0.062794f
C20825 DVDD.n3483 VSS 0.061545f
C20826 DVDD.n3484 VSS 0.140961f
C20827 DVDD.n3485 VSS 0.10175f
C20828 DVDD.n3486 VSS 0.10175f
C20829 DVDD.n3487 VSS 0.070479f
C20830 DVDD.n3488 VSS 0.140961f
C20831 DVDD.n3489 VSS 0.127355f
C20832 DVDD.n3490 VSS 0.14195f
C20833 DVDD.n3491 VSS 0.140961f
C20834 DVDD.n3492 VSS 0.142138f
C20835 DVDD.n3493 VSS 0.063035f
C20836 DVDD.n3494 VSS 0.061545f
C20837 DVDD.n3495 VSS 0.070479f
C20838 DVDD.n3496 VSS 0.061545f
C20839 DVDD.n3497 VSS 0.070479f
C20840 DVDD.n3498 VSS 0.061545f
C20841 DVDD.n3499 VSS 0.140961f
C20842 DVDD.n3500 VSS 0.408805f
C20843 DVDD.n3501 VSS 0.140961f
C20844 DVDD.n3502 VSS 0.240702f
C20845 DVDD.n3503 VSS 0.240702f
C20846 DVDD.n3504 VSS 0.240702f
C20847 DVDD.n3505 VSS 0.240702f
C20848 DVDD.n3506 VSS 0.105095f
C20849 DVDD.n3507 VSS 0.240702f
C20850 DVDD.n3508 VSS 0.220361f
C20851 DVDD.n3509 VSS 0.140692f
C20852 DVDD.n3510 VSS 0.263798f
C20853 DVDD.n3511 VSS 0.413177f
C20854 DVDD.n3512 VSS 0.451316f
C20855 DVDD.n3513 VSS 0.451316f
C20856 DVDD.n3514 VSS 0.451316f
C20857 DVDD.n3515 VSS 0.451316f
C20858 DVDD.n3516 VSS 0.451316f
C20859 DVDD.n3517 VSS 0.451316f
C20860 DVDD.n3518 VSS 0.451316f
C20861 DVDD.n3519 VSS 0.451316f
C20862 DVDD.n3520 VSS 0.451316f
C20863 DVDD.n3521 VSS 0.451316f
C20864 DVDD.n3522 VSS 0.031397f
C20865 DVDD.n3523 VSS 0.031397f
C20866 DVDD.n3524 VSS 0.031397f
C20867 DVDD.n3525 VSS 0.031397f
C20868 DVDD.n3526 VSS 0.031397f
C20869 DVDD.n3527 VSS 0.031397f
C20870 DVDD.n3528 VSS 0.031397f
C20871 DVDD.n3529 VSS 0.031397f
C20872 DVDD.n3530 VSS 0.031397f
C20873 DVDD.n3531 VSS 0.031397f
C20874 DVDD.n3532 VSS 0.062794f
C20875 DVDD.n3533 VSS 0.08912f
C20876 DVDD.n3534 VSS 0.197054f
C20877 DVDD.n3535 VSS 0.062794f
C20878 DVDD.n3536 VSS 0.041779f
C20879 DVDD.n3537 VSS 0.031397f
C20880 DVDD.n3538 VSS 0.031397f
C20881 DVDD.n3539 VSS 0.031397f
C20882 DVDD.n3540 VSS 0.031397f
C20883 DVDD.n3541 VSS 0.031397f
C20884 DVDD.n3542 VSS 0.031397f
C20885 DVDD.n3543 VSS 0.031397f
C20886 DVDD.n3544 VSS 0.031397f
C20887 DVDD.n3545 VSS 0.031397f
C20888 DVDD.n3546 VSS 0.031397f
C20889 DVDD.n3549 VSS 0.225658f
C20890 DVDD.n3551 VSS 0.181162f
C20891 DVDD.n3552 VSS 0.048607f
C20892 DVDD.n3553 VSS 0.131369f
C20893 DVDD.n3554 VSS 0.15585f
C20894 DVDD.n3555 VSS 0.114418f
C20895 DVDD.n3556 VSS 0.054626f
C20896 DVDD.n3557 VSS 0.225658f
C20897 DVDD.n3558 VSS 0.225658f
C20898 DVDD.n3559 VSS 0.033368f
C20899 DVDD.n3560 VSS 0.225658f
C20900 DVDD.n3561 VSS 0.197054f
C20901 DVDD.n3562 VSS 0.029062f
C20902 DVDD.n3563 VSS 0.029062f
C20903 DVDD.n3564 VSS 0.029062f
C20904 DVDD.n3565 VSS 0.029062f
C20905 DVDD.n3566 VSS 0.029062f
C20906 DVDD.n3567 VSS 0.029062f
C20907 DVDD.n3568 VSS 0.029062f
C20908 DVDD.n3569 VSS 0.029062f
C20909 DVDD.n3570 VSS 0.029062f
C20910 DVDD.n3572 VSS 0.066735f
C20911 DVDD.n3574 VSS 0.058124f
C20912 DVDD.n3575 VSS 0.114418f
C20913 DVDD.n3576 VSS 0.124509f
C20914 DVDD.n3577 VSS 0.15585f
C20915 DVDD.n3578 VSS 0.131369f
C20916 DVDD.n3579 VSS 0.026274f
C20917 DVDD.n3580 VSS 0.131369f
C20918 DVDD.n3581 VSS 0.15585f
C20919 DVDD.n3582 VSS 0.15585f
C20920 DVDD.n3583 VSS 0.131369f
C20921 DVDD.n3584 VSS 0.013137f
C20922 DVDD.n3585 VSS 0.451316f
C20923 DVDD.n3586 VSS 0.451316f
C20924 DVDD.n3587 VSS 1.30659f
C20925 DVDD.n3588 VSS 0.455731f
C20926 DVDD.n3589 VSS 0.451316f
C20927 DVDD.n3590 VSS 0.451316f
C20928 DVDD.n3591 VSS 0.197054f
C20929 DVDD.n3592 VSS 0.131369f
C20930 DVDD.n3593 VSS 0.026274f
C20931 DVDD.n3594 VSS 0.131369f
C20932 DVDD.n3595 VSS 0.026274f
C20933 DVDD.n3596 VSS 0.131369f
C20934 DVDD.n3597 VSS 0.026274f
C20935 DVDD.n3598 VSS 0.131369f
C20936 DVDD.n3599 VSS 0.026274f
C20937 DVDD.n3600 VSS 0.131369f
C20938 DVDD.n3601 VSS 0.131369f
C20939 DVDD.n3602 VSS 0.026274f
C20940 DVDD.n3603 VSS 0.026274f
C20941 DVDD.n3604 VSS 0.026274f
C20942 DVDD.n3605 VSS 0.131369f
C20943 DVDD.n3606 VSS 0.131369f
C20944 DVDD.n3607 VSS 0.131369f
C20945 DVDD.n3608 VSS 0.026274f
C20946 DVDD.n3609 VSS 0.026274f
C20947 DVDD.n3610 VSS 0.026274f
C20948 DVDD.n3611 VSS 0.131369f
C20949 DVDD.n3612 VSS 0.131369f
C20950 DVDD.n3613 VSS 0.131369f
C20951 DVDD.n3614 VSS 0.026274f
C20952 DVDD.n3615 VSS 0.026274f
C20953 DVDD.n3616 VSS 0.026274f
C20954 DVDD.n3617 VSS 0.131369f
C20955 DVDD.n3618 VSS 0.131369f
C20956 DVDD.n3619 VSS 0.131369f
C20957 DVDD.n3620 VSS 0.026274f
C20958 DVDD.n3621 VSS 0.026274f
C20959 DVDD.n3622 VSS 0.026274f
C20960 DVDD.n3623 VSS 0.131369f
C20961 DVDD.n3624 VSS 0.131369f
C20962 DVDD.n3625 VSS 0.131369f
C20963 DVDD.n3626 VSS 0.026274f
C20964 DVDD.n3627 VSS 0.014726f
C20965 DVDD.n3628 VSS 0.013137f
C20966 DVDD.n3629 VSS 0.013137f
C20967 DVDD.n3630 VSS 0.131369f
C20968 DVDD.n3631 VSS 0.131369f
C20969 DVDD.n3632 VSS 0.013137f
C20970 DVDD.n3633 VSS 0.013137f
C20971 DVDD.n3634 VSS 0.225658f
C20972 DVDD.n3635 VSS 0.029062f
C20973 DVDD.n3636 VSS 0.032022f
C20974 DVDD.n3637 VSS 0.114418f
C20975 DVDD.n3638 VSS 0.114418f
C20976 DVDD.n3639 VSS 0.114418f
C20977 DVDD.n3640 VSS 0.029062f
C20978 DVDD.n3641 VSS 0.058124f
C20979 DVDD.n3642 VSS 0.114418f
C20980 DVDD.n3643 VSS 0.058124f
C20981 DVDD.n3644 VSS 0.114418f
C20982 DVDD.n3645 VSS 0.058124f
C20983 DVDD.n3646 VSS 0.114418f
C20984 DVDD.n3647 VSS 0.058124f
C20985 DVDD.n3648 VSS 0.114418f
C20986 DVDD.n3649 VSS 0.058124f
C20987 DVDD.n3650 VSS 0.058124f
C20988 DVDD.n3651 VSS 0.114418f
C20989 DVDD.n3652 VSS 0.058124f
C20990 DVDD.n3653 VSS 0.114418f
C20991 DVDD.n3654 VSS 0.058124f
C20992 DVDD.n3655 VSS 0.114418f
C20993 DVDD.n3656 VSS 0.058124f
C20994 DVDD.n3657 VSS 0.114418f
C20995 DVDD.n3658 VSS 0.058124f
C20996 DVDD.n3659 VSS 0.114418f
C20997 DVDD.n3660 VSS 0.058124f
C20998 DVDD.n3661 VSS 0.114418f
C20999 DVDD.n3662 VSS 0.058124f
C21000 DVDD.n3663 VSS 0.114418f
C21001 DVDD.n3664 VSS 0.114418f
C21002 DVDD.n3665 VSS 0.058124f
C21003 DVDD.n3666 VSS 0.058124f
C21004 DVDD.n3667 VSS 0.058124f
C21005 DVDD.n3668 VSS 0.114418f
C21006 DVDD.n3669 VSS 0.114418f
C21007 DVDD.n3670 VSS 0.114418f
C21008 DVDD.n3671 VSS 0.058124f
C21009 DVDD.n3672 VSS 0.058124f
C21010 DVDD.n3673 VSS 0.058124f
C21011 DVDD.n3674 VSS 0.114418f
C21012 DVDD.n3675 VSS 0.114418f
C21013 DVDD.n3676 VSS 0.114418f
C21014 DVDD.n3677 VSS 0.058124f
C21015 DVDD.n3678 VSS 0.058124f
C21016 DVDD.n3679 VSS 0.058124f
C21017 DVDD.n3680 VSS 0.114418f
C21018 DVDD.n3681 VSS 0.114418f
C21019 DVDD.n3682 VSS 0.114418f
C21020 DVDD.n3683 VSS 0.058124f
C21021 DVDD.n3684 VSS 0.058124f
C21022 DVDD.n3685 VSS 0.058124f
C21023 DVDD.n3686 VSS 0.114418f
C21024 DVDD.n3687 VSS 0.114418f
C21025 DVDD.n3688 VSS 0.114418f
C21026 DVDD.n3689 VSS 0.058124f
C21027 DVDD.n3690 VSS 0.058124f
C21028 DVDD.n3691 VSS 0.058124f
C21029 DVDD.n3692 VSS 0.114418f
C21030 DVDD.n3693 VSS 0.114418f
C21031 DVDD.n3694 VSS 0.114418f
C21032 DVDD.n3695 VSS 0.058124f
C21033 DVDD.n3696 VSS 0.058124f
C21034 DVDD.n3697 VSS 0.058124f
C21035 DVDD.n3698 VSS 0.114418f
C21036 DVDD.n3699 VSS 0.114418f
C21037 DVDD.n3700 VSS 0.114418f
C21038 DVDD.n3701 VSS 0.058124f
C21039 DVDD.n3702 VSS 0.277706f
C21040 DVDD.n3703 VSS 0.277706f
C21041 DVDD.n3704 VSS 0.058124f
C21042 DVDD.n3705 VSS 0.114418f
C21043 DVDD.n3706 VSS 0.114418f
C21044 DVDD.n3707 VSS 0.114418f
C21045 DVDD.n3708 VSS 0.058124f
C21046 DVDD.n3709 VSS 0.058124f
C21047 DVDD.n3710 VSS 0.058124f
C21048 DVDD.n3711 VSS 0.114418f
C21049 DVDD.n3712 VSS 0.114418f
C21050 DVDD.n3713 VSS 0.114418f
C21051 DVDD.n3714 VSS 0.058124f
C21052 DVDD.n3715 VSS 0.058124f
C21053 DVDD.n3716 VSS 0.058124f
C21054 DVDD.n3717 VSS 0.114418f
C21055 DVDD.n3718 VSS 0.114418f
C21056 DVDD.n3719 VSS 0.114418f
C21057 DVDD.n3720 VSS 0.058124f
C21058 DVDD.n3721 VSS 0.058124f
C21059 DVDD.n3722 VSS 0.058124f
C21060 DVDD.n3723 VSS 0.114418f
C21061 DVDD.n3724 VSS 0.114418f
C21062 DVDD.n3725 VSS 0.114418f
C21063 DVDD.n3726 VSS 0.058124f
C21064 DVDD.n3727 VSS 0.058124f
C21065 DVDD.n3728 VSS 0.058124f
C21066 DVDD.n3729 VSS 0.114418f
C21067 DVDD.n3730 VSS 0.114418f
C21068 DVDD.n3731 VSS 0.114418f
C21069 DVDD.n3732 VSS 0.058124f
C21070 DVDD.n3733 VSS 0.058124f
C21071 DVDD.n3734 VSS 0.046553f
C21072 DVDD.n3735 VSS 0.114418f
C21073 DVDD.n3736 VSS 0.114418f
C21074 DVDD.n3737 VSS 0.114418f
C21075 DVDD.n3738 VSS 0.114418f
C21076 DVDD.n3739 VSS 0.114418f
C21077 DVDD.n3740 VSS 0.030408f
C21078 DVDD.n3741 VSS 0.029062f
C21079 DVDD.n3742 VSS 0.225658f
C21080 DVDD.n3743 VSS 0.013137f
C21081 DVDD.n3744 VSS 0.013137f
C21082 DVDD.n3745 VSS 0.131369f
C21083 DVDD.n3746 VSS 0.131369f
C21084 DVDD.n3747 VSS 0.013137f
C21085 DVDD.n3748 VSS 0.013137f
C21086 DVDD.n3749 VSS 0.013137f
C21087 DVDD.n3750 VSS 0.124509f
C21088 DVDD.t19 VSS 5.27557f
C21089 DVDD.n3751 VSS 0.124509f
C21090 DVDD.n3752 VSS 0.101257f
C21091 DVDD.n3753 VSS 0.048607f
C21092 DVDD.n3754 VSS 0.131369f
C21093 DVDD.n3755 VSS 0.048607f
C21094 DVDD.n3756 VSS 0.131369f
C21095 DVDD.n3757 VSS 0.048607f
C21096 DVDD.n3758 VSS 0.131369f
C21097 DVDD.n3759 VSS 0.048607f
C21098 DVDD.n3760 VSS 0.131369f
C21099 DVDD.n3761 VSS 0.048607f
C21100 DVDD.n3762 VSS 0.131369f
C21101 DVDD.n3763 VSS 0.048607f
C21102 DVDD.n3764 VSS 0.076786f
C21103 DVDD.n3765 VSS 0.048607f
C21104 DVDD.n3766 VSS 0.131369f
C21105 DVDD.n3767 VSS 0.131369f
C21106 DVDD.n3768 VSS 0.131369f
C21107 DVDD.n3769 VSS 0.048607f
C21108 DVDD.n3770 VSS 0.048607f
C21109 DVDD.n3771 VSS 0.048607f
C21110 DVDD.n3772 VSS 0.131369f
C21111 DVDD.n3773 VSS 0.131369f
C21112 DVDD.n3774 VSS 0.131369f
C21113 DVDD.n3775 VSS 0.048607f
C21114 DVDD.n3776 VSS 0.048607f
C21115 DVDD.n3777 VSS 0.048607f
C21116 DVDD.n3778 VSS 0.131369f
C21117 DVDD.n3779 VSS 0.131369f
C21118 DVDD.n3780 VSS 0.131369f
C21119 DVDD.n3781 VSS 0.048607f
C21120 DVDD.n3782 VSS 0.048607f
C21121 DVDD.n3783 VSS 0.048607f
C21122 DVDD.n3784 VSS 0.131369f
C21123 DVDD.n3785 VSS 0.131369f
C21124 DVDD.n3786 VSS 0.131369f
C21125 DVDD.n3787 VSS 0.048607f
C21126 DVDD.n3788 VSS 0.048607f
C21127 DVDD.n3789 VSS 0.048607f
C21128 DVDD.n3790 VSS 0.131369f
C21129 DVDD.n3791 VSS 0.131369f
C21130 DVDD.n3792 VSS 0.131369f
C21131 DVDD.n3793 VSS 0.048607f
C21132 DVDD.n3794 VSS 0.048607f
C21133 DVDD.n3795 VSS 0.048607f
C21134 DVDD.n3796 VSS 0.131369f
C21135 DVDD.n3797 VSS 0.131369f
C21136 DVDD.n3798 VSS 0.131369f
C21137 DVDD.n3799 VSS 0.048607f
C21138 DVDD.n3800 VSS 0.048607f
C21139 DVDD.n3801 VSS 0.122706f
C21140 DVDD.n3802 VSS 0.124509f
C21141 DVDD.t11 VSS 5.27557f
C21142 DVDD.n3803 VSS 0.15585f
C21143 DVDD.n3804 VSS 0.156344f
C21144 DVDD.n3805 VSS 0.066735f
C21145 DVDD.n3807 VSS 0.16065f
C21146 DVDD.n3808 VSS 0.395696f
C21147 DVDD.n3809 VSS 0.029062f
C21148 DVDD.n3810 VSS 0.029062f
C21149 DVDD.n3811 VSS 0.029062f
C21150 DVDD.n3812 VSS 0.029062f
C21151 DVDD.n3813 VSS 0.029062f
C21152 DVDD.n3814 VSS 0.029062f
C21153 DVDD.n3815 VSS 0.029062f
C21154 DVDD.n3816 VSS 0.029062f
C21155 DVDD.n3817 VSS 0.029062f
C21156 DVDD.n3818 VSS 0.033368f
C21157 DVDD.n3819 VSS 0.058124f
C21158 DVDD.n3820 VSS 0.033368f
C21159 DVDD.n3821 VSS 0.114418f
C21160 DVDD.n3822 VSS 0.033368f
C21161 DVDD.n3823 VSS 0.114418f
C21162 DVDD.n3824 VSS 0.114418f
C21163 DVDD.n3825 VSS 0.033099f
C21164 DVDD.n3826 VSS 0.029331f
C21165 DVDD.n3827 VSS 0.114418f
C21166 DVDD.n3828 VSS 0.033368f
C21167 DVDD.n3829 VSS 0.114418f
C21168 DVDD.n3830 VSS 0.033368f
C21169 DVDD.n3831 VSS 0.114418f
C21170 DVDD.n3832 VSS 0.033368f
C21171 DVDD.n3833 VSS 0.114418f
C21172 DVDD.n3834 VSS 0.033368f
C21173 DVDD.n3835 VSS 0.114418f
C21174 DVDD.n3836 VSS 0.033368f
C21175 DVDD.n3837 VSS 0.114418f
C21176 DVDD.n3838 VSS 0.033368f
C21177 DVDD.n3839 VSS 0.114418f
C21178 DVDD.n3840 VSS 0.114418f
C21179 DVDD.n3841 VSS 0.032022f
C21180 DVDD.n3842 VSS 0.030408f
C21181 DVDD.n3843 VSS 0.114418f
C21182 DVDD.n3844 VSS 0.033368f
C21183 DVDD.n3845 VSS 0.114418f
C21184 DVDD.n3846 VSS 0.033368f
C21185 DVDD.n3847 VSS 0.114418f
C21186 DVDD.n3848 VSS 0.033368f
C21187 DVDD.n3849 VSS 0.114418f
C21188 DVDD.n3850 VSS 0.033368f
C21189 DVDD.n3851 VSS 0.114418f
C21190 DVDD.n3852 VSS 0.033368f
C21191 DVDD.n3853 VSS 0.114418f
C21192 DVDD.n3854 VSS 0.033368f
C21193 DVDD.n3855 VSS 0.114418f
C21194 DVDD.n3856 VSS 0.114418f
C21195 DVDD.n3857 VSS 0.030946f
C21196 DVDD.n3858 VSS 0.031484f
C21197 DVDD.n3859 VSS 0.114418f
C21198 DVDD.n3860 VSS 0.114418f
C21199 DVDD.n3861 VSS 0.114418f
C21200 DVDD.n3862 VSS 0.120351f
C21201 DVDD.n3863 VSS 0.033368f
C21202 DVDD.n3864 VSS 0.120351f
C21203 DVDD.n3865 VSS 0.061117f
C21204 DVDD.n3866 VSS 0.026274f
C21205 DVDD.n3867 VSS 0.033368f
C21206 DVDD.n3868 VSS 0.030088f
C21207 DVDD.n3869 VSS 0.060175f
C21208 DVDD.n3870 VSS 0.173937f
C21209 DVDD.n3871 VSS 0.060175f
C21210 DVDD.n3872 VSS 0.044284f
C21211 DVDD.n3873 VSS 0.026274f
C21212 DVDD.n3874 VSS 0.061085f
C21213 DVDD.n3876 VSS 0.172475f
C21214 DVDD.n3878 VSS 0.026274f
C21215 DVDD.n3879 VSS 0.030088f
C21216 DVDD.n3880 VSS 0.045979f
C21217 DVDD.n3881 VSS 0.044284f
C21218 DVDD.n3882 VSS 0.215276f
C21219 DVDD.n3883 VSS 0.240702f
C21220 DVDD.n3884 VSS 0.172475f
C21221 DVDD.n3885 VSS 0.092382f
C21222 DVDD.n3886 VSS 0.240702f
C21223 DVDD.n3887 VSS 0.211038f
C21224 DVDD.n3888 VSS 0.240702f
C21225 DVDD.n3889 VSS 0.240702f
C21226 DVDD.n3890 VSS 0.240702f
C21227 DVDD.n3891 VSS 0.240702f
C21228 DVDD.n3892 VSS 0.240702f
C21229 DVDD.n3893 VSS 0.451316f
C21230 DVDD.n3894 VSS 0.451316f
C21231 DVDD.n3895 VSS 0.451316f
C21232 DVDD.n3896 VSS 0.451316f
C21233 DVDD.n3897 VSS 0.451316f
C21234 DVDD.n3898 VSS 0.451316f
C21235 DVDD.n3899 VSS 0.451316f
C21236 DVDD.n3900 VSS 0.451316f
C21237 DVDD.n3901 VSS 0.451316f
C21238 DVDD.n3902 VSS 0.451316f
C21239 DVDD.n3903 VSS 0.451316f
C21240 DVDD.n3904 VSS 0.451316f
C21241 DVDD.n3905 VSS 0.451316f
C21242 DVDD.n3906 VSS 0.451316f
C21243 DVDD.n3907 VSS 0.451316f
C21244 DVDD.n3908 VSS 0.451316f
C21245 DVDD.n3909 VSS 0.451316f
C21246 DVDD.n3910 VSS 0.451316f
C21247 DVDD.n3911 VSS 0.451316f
C21248 DVDD.n3912 VSS 0.346009f
C21249 DVDD.n3913 VSS 0.346009f
C21250 DVDD.n3914 VSS 0.147472f
C21251 DVDD.n3915 VSS 0.240702f
C21252 DVDD.n3916 VSS 0.240702f
C21253 DVDD.n3917 VSS 0.240702f
C21254 DVDD.n3918 VSS 0.240702f
C21255 DVDD.n3919 VSS 0.240702f
C21256 DVDD.n3920 VSS 0.240702f
C21257 DVDD.n3921 VSS 0.240702f
C21258 DVDD.n3922 VSS 0.240702f
C21259 DVDD.n3923 VSS 0.215276f
C21260 DVDD.n3924 VSS 0.215276f
C21261 DVDD.n3925 VSS 0.240702f
C21262 DVDD.n3926 VSS 0.240702f
C21263 DVDD.n3927 VSS 0.240702f
C21264 DVDD.n3928 VSS 0.240702f
C21265 DVDD.n3929 VSS 0.240702f
C21266 DVDD.n3930 VSS 0.240702f
C21267 DVDD.n3931 VSS 0.240702f
C21268 DVDD.n3932 VSS 0.240702f
C21269 DVDD.n3933 VSS 0.240702f
C21270 DVDD.n3934 VSS 0.240702f
C21271 DVDD.n3935 VSS 0.240702f
C21272 DVDD.n3936 VSS 0.240702f
C21273 DVDD.n3937 VSS 0.240702f
C21274 DVDD.n3938 VSS 0.240702f
C21275 DVDD.n3939 VSS 0.240702f
C21276 DVDD.n3940 VSS 0.240702f
C21277 DVDD.n3941 VSS 0.213581f
C21278 DVDD.n3942 VSS 0.213581f
C21279 DVDD.n3943 VSS 0.213581f
C21280 DVDD.n3944 VSS 0.451316f
C21281 DVDD.n3945 VSS 0.451316f
C21282 DVDD.n3946 VSS 0.197054f
C21283 DVDD.n3947 VSS 0.066735f
C21284 DVDD.n3948 VSS 0.054626f
C21285 DVDD.n3949 VSS 0.029062f
C21286 DVDD.n3950 VSS 0.029062f
C21287 DVDD.n3951 VSS 0.029062f
C21288 DVDD.n3952 VSS 0.029062f
C21289 DVDD.n3953 VSS 0.029062f
C21290 DVDD.n3954 VSS 0.029062f
C21291 DVDD.n3955 VSS 0.029062f
C21292 DVDD.n3956 VSS 0.029062f
C21293 DVDD.n3957 VSS 0.029062f
C21294 DVDD.n3958 VSS 0.029062f
C21295 DVDD.n3959 VSS 0.029062f
C21296 DVDD.n3960 VSS 0.029062f
C21297 DVDD.n3961 VSS 0.029062f
C21298 DVDD.n3962 VSS 0.029062f
C21299 DVDD.n3963 VSS 0.029062f
C21300 DVDD.n3964 VSS 0.029062f
C21301 DVDD.n3965 VSS 0.029062f
C21302 DVDD.n3966 VSS 0.029062f
C21303 DVDD.n3967 VSS 0.029062f
C21304 DVDD.n3968 VSS 0.029062f
C21305 DVDD.n3969 VSS 0.066735f
C21306 DVDD.n3970 VSS 0.058124f
C21307 DVDD.n3971 VSS 0.114418f
C21308 DVDD.n3972 VSS 0.114418f
C21309 DVDD.n3973 VSS 0.058124f
C21310 DVDD.n3974 VSS 0.114418f
C21311 DVDD.n3975 VSS 0.114418f
C21312 DVDD.n3976 VSS 0.066735f
C21313 DVDD.n3977 VSS 0.225658f
C21314 DVDD.n3978 VSS 0.451316f
C21315 DVDD.n3979 VSS 0.724649f
C21316 DVDD.n3980 VSS 0.724649f
C21317 DVDD.n3981 VSS 0.225658f
C21318 DVDD.n3982 VSS 0.197054f
C21319 DVDD.n3983 VSS 0.217712f
C21320 DVDD.n3984 VSS 0.033099f
C21321 DVDD.n3985 VSS 0.197054f
C21322 DVDD.n3986 VSS 0.535541f
C21323 DVDD.n3987 VSS 0.451316f
C21324 DVDD.n3988 VSS 0.451316f
C21325 DVDD.n3989 VSS 0.344844f
C21326 DVDD.n3990 VSS 0.451316f
C21327 DVDD.n3991 VSS 0.225658f
C21328 DVDD.n3992 VSS 0.204999f
C21329 DVDD.n3993 VSS 0.033368f
C21330 DVDD.n3994 VSS 0.029062f
C21331 DVDD.n3995 VSS 0.114418f
C21332 DVDD.n3996 VSS 0.114418f
C21333 DVDD.n3997 VSS 0.033368f
C21334 DVDD.n3998 VSS 0.429855f
C21335 DVDD.n3999 VSS 0.204999f
C21336 DVDD.n4000 VSS 0.197054f
C21337 DVDD.n4001 VSS 0.225658f
C21338 DVDD.n4002 VSS 0.033368f
C21339 DVDD.n4003 VSS 0.114418f
C21340 DVDD.n4004 VSS 0.029062f
C21341 DVDD.n4005 VSS 0.114418f
C21342 DVDD.n4006 VSS 0.114418f
C21343 DVDD.n4007 VSS 0.029331f
C21344 DVDD.n4008 VSS 0.033099f
C21345 DVDD.n4009 VSS 0.217712f
C21346 DVDD.n4010 VSS 0.029062f
C21347 DVDD.n4011 VSS 0.029062f
C21348 DVDD.n4012 VSS 0.033368f
C21349 DVDD.n4013 VSS 0.114418f
C21350 DVDD.n4014 VSS 0.114418f
C21351 DVDD.n4015 VSS 0.114418f
C21352 DVDD.n4016 VSS 0.033368f
C21353 DVDD.n4017 VSS 0.225658f
C21354 DVDD.n4018 VSS 0.332131f
C21355 DVDD.n4019 VSS 0.451316f
C21356 DVDD.n4020 VSS 0.750075f
C21357 DVDD.n4021 VSS 0.197054f
C21358 DVDD.n4022 VSS 0.548254f
C21359 DVDD.n4023 VSS 0.548254f
C21360 DVDD.n4024 VSS 0.451316f
C21361 DVDD.n4025 VSS 0.451316f
C21362 DVDD.n4026 VSS 0.197054f
C21363 DVDD.n4027 VSS 0.225658f
C21364 DVDD.n4028 VSS 0.033368f
C21365 DVDD.n4029 VSS 0.114418f
C21366 DVDD.n4030 VSS 0.033368f
C21367 DVDD.n4031 VSS 0.220891f
C21368 DVDD.n4032 VSS 0.029062f
C21369 DVDD.n4033 VSS 0.114418f
C21370 DVDD.n4034 VSS 0.029062f
C21371 DVDD.n4035 VSS 0.114418f
C21372 DVDD.n4036 VSS 0.029062f
C21373 DVDD.n4037 VSS 0.032561f
C21374 DVDD.n4038 VSS 0.114418f
C21375 DVDD.n4039 VSS 0.114418f
C21376 DVDD.n4040 VSS 0.029869f
C21377 DVDD.n4041 VSS 0.197054f
C21378 DVDD.n4042 VSS 0.225658f
C21379 DVDD.n4043 VSS 0.029062f
C21380 DVDD.n4044 VSS 0.033368f
C21381 DVDD.n4045 VSS 0.220891f
C21382 DVDD.n4046 VSS 0.201821f
C21383 DVDD.n4047 VSS 0.029062f
C21384 DVDD.n4048 VSS 0.033368f
C21385 DVDD.n4049 VSS 0.114418f
C21386 DVDD.n4050 VSS 0.114418f
C21387 DVDD.n4051 VSS 0.048706f
C21388 DVDD.n4052 VSS 0.058124f
C21389 DVDD.n4053 VSS 0.048168f
C21390 DVDD.n4054 VSS 0.114418f
C21391 DVDD.n4055 VSS 0.114418f
C21392 DVDD.n4056 VSS 0.114418f
C21393 DVDD.n4057 VSS 0.033368f
C21394 DVDD.n4058 VSS 0.029062f
C21395 DVDD.n4059 VSS 0.201821f
C21396 DVDD.n4060 VSS 0.197054f
C21397 DVDD.n4061 VSS 0.225658f
C21398 DVDD.n4062 VSS 0.029062f
C21399 DVDD.n4063 VSS 0.030408f
C21400 DVDD.n4064 VSS 0.029062f
C21401 DVDD.n4065 VSS 0.032022f
C21402 DVDD.n4066 VSS 0.114418f
C21403 DVDD.n4067 VSS 0.114418f
C21404 DVDD.n4068 VSS 0.114418f
C21405 DVDD.n4069 VSS 0.029062f
C21406 DVDD.n4070 VSS 0.033368f
C21407 DVDD.n4071 VSS 0.197054f
C21408 DVDD.n4072 VSS 0.225658f
C21409 DVDD.n4073 VSS 0.029062f
C21410 DVDD.n4074 VSS 0.033368f
C21411 DVDD.n4075 VSS 0.114418f
C21412 DVDD.n4076 VSS 0.114418f
C21413 DVDD.n4077 VSS 0.033368f
C21414 DVDD.n4078 VSS 0.029062f
C21415 DVDD.n4079 VSS 0.225658f
C21416 DVDD.n4080 VSS 0.197054f
C21417 DVDD.n4081 VSS 0.332131f
C21418 DVDD.n4082 VSS 0.451316f
C21419 DVDD.n4083 VSS 0.451316f
C21420 DVDD.n4084 VSS 0.451316f
C21421 DVDD.n4085 VSS 0.451316f
C21422 DVDD.n4086 VSS 0.750075f
C21423 DVDD.n4087 VSS 0.750075f
C21424 DVDD.n4088 VSS 0.750075f
C21425 DVDD.n4089 VSS 0.451316f
C21426 DVDD.n4090 VSS 0.451316f
C21427 DVDD.n4091 VSS 0.451316f
C21428 DVDD.n4092 VSS 0.451316f
C21429 DVDD.n4093 VSS 0.451316f
C21430 DVDD.n4094 VSS 0.197054f
C21431 DVDD.n4095 VSS 0.225658f
C21432 DVDD.n4096 VSS 0.029062f
C21433 DVDD.n4097 VSS 0.033368f
C21434 DVDD.n4098 VSS 0.114418f
C21435 DVDD.n4099 VSS 0.114418f
C21436 DVDD.n4100 VSS 0.033368f
C21437 DVDD.n4101 VSS 0.029062f
C21438 DVDD.n4102 VSS 0.225658f
C21439 DVDD.n4103 VSS 0.197054f
C21440 DVDD.n4104 VSS 0.344844f
C21441 DVDD.n4105 VSS 0.451316f
C21442 DVDD.n4106 VSS 0.451316f
C21443 DVDD.n4107 VSS 1.28214f
C21444 DVDD.n4108 VSS 0.451316f
C21445 DVDD.n4109 VSS 0.451316f
C21446 DVDD.n4110 VSS 0.197054f
C21447 DVDD.n4111 VSS 0.447648f
C21448 DVDD.n4112 VSS 0.029062f
C21449 DVDD.n4113 VSS 0.05355f
C21450 DVDD.n4114 VSS 0.277706f
C21451 DVDD.n4115 VSS 0.15585f
C21452 DVDD.t24 VSS 5.27557f
C21453 DVDD.n4117 VSS 0.15585f
C21454 DVDD.n4118 VSS 0.029331f
C21455 DVDD.n4119 VSS 0.114418f
C21456 DVDD.n4120 VSS 0.114418f
C21457 DVDD.n4121 VSS 0.033368f
C21458 DVDD.n4122 VSS 0.029062f
C21459 DVDD.n4123 VSS 0.217712f
C21460 DVDD.n4124 VSS 0.197054f
C21461 DVDD.n4125 VSS 0.451316f
C21462 DVDD.n4126 VSS 0.451316f
C21463 DVDD.n4127 VSS 0.451316f
C21464 DVDD.n4128 VSS 0.724649f
C21465 DVDD.n4129 VSS 0.724649f
C21466 DVDD.n4130 VSS 0.535541f
C21467 DVDD.n4131 VSS 0.225658f
C21468 DVDD.n4132 VSS 0.10091f
C21469 DVDD.n4133 VSS 0.130242f
C21470 DVDD.n4134 VSS 0.066735f
C21471 DVDD.n4135 VSS 0.066735f
C21472 DVDD.n4136 VSS 0.204999f
C21473 DVDD.n4137 VSS 0.197054f
C21474 DVDD.n4138 VSS 0.451316f
C21475 DVDD.n4139 VSS 0.451316f
C21476 DVDD.n4140 VSS 0.451316f
C21477 DVDD.n4141 VSS 0.451316f
C21478 DVDD.n4142 VSS 0.451316f
C21479 DVDD.n4143 VSS 0.197054f
C21480 DVDD.n4144 VSS 0.197054f
C21481 DVDD.n4145 VSS 0.225658f
C21482 DVDD.n4146 VSS 0.04763f
C21483 DVDD.n4147 VSS 0.033368f
C21484 DVDD.n4148 VSS 0.197054f
C21485 DVDD.n4149 VSS 0.225658f
C21486 DVDD.n4150 VSS 0.451316f
C21487 DVDD.n4151 VSS 0.456124f
C21488 DVDD.n4152 VSS 0.197054f
C21489 DVDD.n4153 VSS 0.225658f
C21490 DVDD.n4154 VSS 0.033368f
C21491 DVDD.n4155 VSS 0.029062f
C21492 DVDD.n4156 VSS 0.114418f
C21493 DVDD.n4157 VSS 0.114418f
C21494 DVDD.n4158 VSS 0.029062f
C21495 DVDD.n4159 VSS 0.030408f
C21496 DVDD.n4160 VSS 0.029062f
C21497 DVDD.n4161 VSS 0.032022f
C21498 DVDD.n4162 VSS 0.114418f
C21499 DVDD.n4163 VSS 0.114418f
C21500 DVDD.n4164 VSS 0.114418f
C21501 DVDD.n4165 VSS 0.058124f
C21502 DVDD.n4166 VSS 0.114418f
C21503 DVDD.n4167 VSS 0.058124f
C21504 DVDD.n4168 VSS 0.114418f
C21505 DVDD.n4169 VSS 0.058124f
C21506 DVDD.n4170 VSS 0.114418f
C21507 DVDD.n4171 VSS 0.058124f
C21508 DVDD.n4172 VSS 0.114418f
C21509 DVDD.n4173 VSS 0.058124f
C21510 DVDD.n4174 VSS 0.114418f
C21511 DVDD.n4175 VSS 0.114418f
C21512 DVDD.n4176 VSS 0.058124f
C21513 DVDD.n4177 VSS 0.058124f
C21514 DVDD.n4178 VSS 0.058124f
C21515 DVDD.n4179 VSS 0.114418f
C21516 DVDD.n4180 VSS 0.114418f
C21517 DVDD.n4181 VSS 0.114418f
C21518 DVDD.n4182 VSS 0.058124f
C21519 DVDD.n4183 VSS 0.058124f
C21520 DVDD.n4184 VSS 0.058124f
C21521 DVDD.n4185 VSS 0.114418f
C21522 DVDD.n4186 VSS 0.114418f
C21523 DVDD.n4187 VSS 0.114418f
C21524 DVDD.n4188 VSS 0.058124f
C21525 DVDD.n4189 VSS 0.058124f
C21526 DVDD.n4190 VSS 0.058124f
C21527 DVDD.n4191 VSS 0.114418f
C21528 DVDD.n4192 VSS 0.114418f
C21529 DVDD.n4193 VSS 0.114418f
C21530 DVDD.n4194 VSS 0.058124f
C21531 DVDD.n4195 VSS 0.058124f
C21532 DVDD.n4196 VSS 0.058124f
C21533 DVDD.n4197 VSS 0.114418f
C21534 DVDD.n4198 VSS 0.114418f
C21535 DVDD.n4199 VSS 0.114418f
C21536 DVDD.n4200 VSS 0.058124f
C21537 DVDD.n4201 VSS 0.058124f
C21538 DVDD.n4202 VSS 0.046553f
C21539 DVDD.n4203 VSS 0.114418f
C21540 DVDD.n4204 VSS 0.114418f
C21541 DVDD.n4205 VSS 0.033368f
C21542 DVDD.n4206 VSS 0.029062f
C21543 DVDD.n4207 VSS 0.201821f
C21544 DVDD.n4208 VSS 0.197054f
C21545 DVDD.n4209 VSS 0.451316f
C21546 DVDD.n4210 VSS 0.455731f
C21547 DVDD.n4211 VSS 1.30659f
C21548 DVDD.n4212 VSS 0.451316f
C21549 DVDD.n4213 VSS 0.451316f
C21550 DVDD.n4214 VSS 0.197054f
C21551 DVDD.n4215 VSS 0.225658f
C21552 DVDD.n4216 VSS 0.029062f
C21553 DVDD.n4217 VSS 0.033368f
C21554 DVDD.n4218 VSS 0.029062f
C21555 DVDD.n4219 VSS 0.033368f
C21556 DVDD.n4220 VSS 0.15585f
C21557 DVDD.t34 VSS 5.27557f
C21558 DVDD.n4222 VSS 0.15585f
C21559 DVDD.n4223 VSS 0.277706f
C21560 DVDD.n4224 VSS 0.058124f
C21561 DVDD.n4225 VSS 0.114418f
C21562 DVDD.n4226 VSS 0.058124f
C21563 DVDD.n4227 VSS 0.114418f
C21564 DVDD.n4228 VSS 0.058124f
C21565 DVDD.n4229 VSS 0.114418f
C21566 DVDD.n4230 VSS 0.058124f
C21567 DVDD.n4231 VSS 0.114418f
C21568 DVDD.n4232 VSS 0.058124f
C21569 DVDD.n4233 VSS 0.114418f
C21570 DVDD.n4234 VSS 0.058124f
C21571 DVDD.n4235 VSS 0.114418f
C21572 DVDD.n4236 VSS 0.114418f
C21573 DVDD.n4237 VSS 0.058124f
C21574 DVDD.n4238 VSS 0.058124f
C21575 DVDD.n4239 VSS 0.058124f
C21576 DVDD.n4240 VSS 0.114418f
C21577 DVDD.n4241 VSS 0.114418f
C21578 DVDD.n4242 VSS 0.114418f
C21579 DVDD.n4243 VSS 0.058124f
C21580 DVDD.n4244 VSS 0.058124f
C21581 DVDD.n4245 VSS 0.058124f
C21582 DVDD.n4246 VSS 0.114418f
C21583 DVDD.n4247 VSS 0.114418f
C21584 DVDD.n4248 VSS 0.114418f
C21585 DVDD.n4249 VSS 0.058124f
C21586 DVDD.n4250 VSS 0.058124f
C21587 DVDD.n4251 VSS 0.058124f
C21588 DVDD.n4252 VSS 0.114418f
C21589 DVDD.n4253 VSS 0.114418f
C21590 DVDD.n4254 VSS 0.114418f
C21591 DVDD.n4255 VSS 0.058124f
C21592 DVDD.n4256 VSS 0.058124f
C21593 DVDD.n4257 VSS 0.058124f
C21594 DVDD.n4258 VSS 0.114418f
C21595 DVDD.n4259 VSS 0.114418f
C21596 DVDD.n4260 VSS 0.114418f
C21597 DVDD.n4261 VSS 0.058124f
C21598 DVDD.n4262 VSS 0.058124f
C21599 DVDD.n4263 VSS 0.058124f
C21600 DVDD.n4264 VSS 0.114418f
C21601 DVDD.n4265 VSS 0.114418f
C21602 DVDD.n4266 VSS 0.114418f
C21603 DVDD.n4267 VSS 0.058124f
C21604 DVDD.n4268 VSS 0.058124f
C21605 DVDD.n4269 VSS 0.058124f
C21606 DVDD.n4270 VSS 0.114418f
C21607 DVDD.n4271 VSS 0.114418f
C21608 DVDD.n4272 VSS 0.114418f
C21609 DVDD.n4273 VSS 0.058124f
C21610 DVDD.n4274 VSS 0.058124f
C21611 DVDD.n4275 VSS 0.277706f
C21612 DVDD.n4276 VSS 0.15585f
C21613 DVDD.t27 VSS 5.27557f
C21614 DVDD.n4278 VSS 0.15585f
C21615 DVDD.n4279 VSS 0.156344f
C21616 DVDD.n4282 VSS 0.225658f
C21617 DVDD.n4283 VSS 0.197054f
C21618 DVDD.n4285 VSS 0.225658f
C21619 DVDD.n4286 VSS 0.451316f
C21620 DVDD.n4287 VSS 0.451316f
C21621 DVDD.n4288 VSS 0.451316f
C21622 DVDD.n4289 VSS 0.451316f
C21623 DVDD.n4290 VSS 0.451316f
C21624 DVDD.n4291 VSS 0.451316f
C21625 DVDD.n4292 VSS 0.451316f
C21626 DVDD.n4293 VSS 0.451316f
C21627 DVDD.n4294 VSS 0.451316f
C21628 DVDD.n4295 VSS 0.451316f
C21629 DVDD.n4296 VSS 0.451316f
C21630 DVDD.n4297 VSS 0.451316f
C21631 DVDD.n4298 VSS 0.451316f
C21632 DVDD.n4299 VSS 0.451316f
C21633 DVDD.n4300 VSS 0.451316f
C21634 DVDD.n4301 VSS 0.360735f
C21635 DVDD.n4302 VSS 0.451316f
C21636 DVDD.n4303 VSS 0.451316f
C21637 DVDD.n4304 VSS 0.451316f
C21638 DVDD.n4305 VSS 0.225658f
C21639 DVDD.n4306 VSS 0.029062f
C21640 DVDD.n4307 VSS 0.029062f
C21641 DVDD.n4308 VSS 0.029062f
C21642 DVDD.n4309 VSS 0.029062f
C21643 DVDD.n4310 VSS 0.029062f
C21644 DVDD.n4311 VSS 0.029062f
C21645 DVDD.n4312 VSS 0.029062f
C21646 DVDD.n4313 VSS 0.029062f
C21647 DVDD.n4314 VSS 0.029062f
C21648 DVDD.n4315 VSS 0.029062f
C21649 DVDD.n4317 VSS 0.058124f
C21650 DVDD.n4318 VSS 0.114418f
C21651 DVDD.n4319 VSS 0.114418f
C21652 DVDD.n4320 VSS 0.058124f
C21653 DVDD.n4321 VSS 0.114418f
C21654 DVDD.n4322 VSS 0.058124f
C21655 DVDD.n4323 VSS 0.114418f
C21656 DVDD.n4324 VSS 0.058124f
C21657 DVDD.n4325 VSS 0.114418f
C21658 DVDD.n4326 VSS 0.058124f
C21659 DVDD.n4327 VSS 0.114418f
C21660 DVDD.n4328 VSS 0.058124f
C21661 DVDD.n4329 VSS 0.114418f
C21662 DVDD.n4330 VSS 0.058124f
C21663 DVDD.n4331 VSS 0.114418f
C21664 DVDD.n4332 VSS 0.114418f
C21665 DVDD.n4333 VSS 0.058124f
C21666 DVDD.n4334 VSS 0.058124f
C21667 DVDD.n4335 VSS 0.058124f
C21668 DVDD.n4336 VSS 0.114418f
C21669 DVDD.n4337 VSS 0.114418f
C21670 DVDD.n4338 VSS 0.114418f
C21671 DVDD.n4339 VSS 0.058124f
C21672 DVDD.n4340 VSS 0.058124f
C21673 DVDD.n4341 VSS 0.058124f
C21674 DVDD.n4342 VSS 0.114418f
C21675 DVDD.n4343 VSS 0.114418f
C21676 DVDD.n4344 VSS 0.114418f
C21677 DVDD.n4345 VSS 0.058124f
C21678 DVDD.n4346 VSS 0.058124f
C21679 DVDD.n4347 VSS 0.058124f
C21680 DVDD.n4348 VSS 0.114418f
C21681 DVDD.n4349 VSS 0.114418f
C21682 DVDD.n4350 VSS 0.114418f
C21683 DVDD.n4351 VSS 0.058124f
C21684 DVDD.n4352 VSS 0.058124f
C21685 DVDD.n4353 VSS 0.058124f
C21686 DVDD.n4354 VSS 0.114418f
C21687 DVDD.n4355 VSS 0.114418f
C21688 DVDD.n4356 VSS 0.114418f
C21689 DVDD.n4357 VSS 0.058124f
C21690 DVDD.n4358 VSS 0.058124f
C21691 DVDD.n4359 VSS 0.058124f
C21692 DVDD.n4360 VSS 0.114418f
C21693 DVDD.n4361 VSS 0.114418f
C21694 DVDD.n4362 VSS 0.114418f
C21695 DVDD.n4363 VSS 0.058124f
C21696 DVDD.n4364 VSS 0.058124f
C21697 DVDD.n4365 VSS 0.058124f
C21698 DVDD.n4366 VSS 0.114418f
C21699 DVDD.n4367 VSS 0.114418f
C21700 DVDD.n4368 VSS 0.114418f
C21701 DVDD.n4369 VSS 0.058124f
C21702 DVDD.n4370 VSS 0.058124f
C21703 DVDD.n4371 VSS 0.277706f
C21704 DVDD.n4372 VSS 0.15585f
C21705 DVDD.t8 VSS 5.27557f
C21706 DVDD.n4374 VSS 0.15585f
C21707 DVDD.n4375 VSS 0.156344f
C21708 DVDD.n4376 VSS 0.16065f
C21709 DVDD.n4377 VSS 0.054626f
C21710 DVDD.n4378 VSS 0.029062f
C21711 DVDD.n4379 VSS 0.029062f
C21712 DVDD.n4380 VSS 0.029062f
C21713 DVDD.n4381 VSS 0.029062f
C21714 DVDD.n4382 VSS 0.029062f
C21715 DVDD.n4383 VSS 0.029062f
C21716 DVDD.n4384 VSS 0.029062f
C21717 DVDD.n4385 VSS 0.029062f
C21718 DVDD.n4386 VSS 0.029062f
C21719 DVDD.n4387 VSS 0.033368f
C21720 DVDD.n4388 VSS 0.225658f
C21721 DVDD.n4389 VSS 0.051397f
C21722 DVDD.n4390 VSS 0.387751f
C21723 DVDD.n4391 VSS 0.289224f
C21724 DVDD.n4392 VSS 0.154253f
C21725 DVDD.n4393 VSS 0.240702f
C21726 DVDD.n4394 VSS 0.346009f
C21727 DVDD.n4395 VSS 0.240702f
C21728 DVDD.n4396 VSS 0.240702f
C21729 DVDD.n4397 VSS 0.240702f
C21730 DVDD.n4398 VSS 0.240702f
C21731 DVDD.n4399 VSS 0.240702f
C21732 DVDD.n4400 VSS 0.240702f
C21733 DVDD.n4401 VSS 0.240702f
C21734 DVDD.n4402 VSS 0.240702f
C21735 DVDD.n4403 VSS 0.240702f
C21736 DVDD.n4404 VSS 0.154253f
C21737 DVDD.n4405 VSS 0.154253f
C21738 DVDD.n4406 VSS 0.240702f
C21739 DVDD.n4407 VSS 0.240702f
C21740 DVDD.n4408 VSS 0.240702f
C21741 DVDD.n4409 VSS 0.240702f
C21742 DVDD.n4410 VSS 0.240702f
C21743 DVDD.n4411 VSS 0.240702f
C21744 DVDD.n4412 VSS 0.240702f
C21745 DVDD.n4413 VSS 0.240702f
C21746 DVDD.n4414 VSS 0.240702f
C21747 DVDD.n4415 VSS 0.240702f
C21748 DVDD.n4416 VSS 0.240702f
C21749 DVDD.n4417 VSS 0.240702f
C21750 DVDD.n4418 VSS 0.240702f
C21751 DVDD.n4419 VSS 0.240702f
C21752 DVDD.n4420 VSS 0.240702f
C21753 DVDD.n4421 VSS 0.240702f
C21754 DVDD.n4422 VSS 0.240702f
C21755 DVDD.n4423 VSS 0.240702f
C21756 DVDD.n4424 VSS 0.240702f
C21757 DVDD.n4425 VSS 0.154253f
C21758 DVDD.n4426 VSS 0.154253f
C21759 DVDD.n4427 VSS 0.451316f
C21760 DVDD.n4428 VSS 0.451316f
C21761 DVDD.n4429 VSS 0.451316f
C21762 DVDD.n4430 VSS 0.451316f
C21763 DVDD.n4431 VSS 0.451316f
C21764 DVDD.n4432 VSS 0.451316f
C21765 DVDD.n4433 VSS 0.451316f
C21766 DVDD.n4434 VSS 0.451316f
C21767 DVDD.n4435 VSS 0.451316f
C21768 DVDD.n4436 VSS 0.451316f
C21769 DVDD.n4437 VSS 0.451316f
C21770 DVDD.n4438 VSS 0.197054f
C21771 DVDD.n4439 VSS 0.451316f
C21772 DVDD.n4440 VSS 0.451316f
C21773 DVDD.n4441 VSS 0.451316f
C21774 DVDD.n4442 VSS 0.451316f
C21775 DVDD.n4443 VSS 0.451316f
C21776 DVDD.n4444 VSS 0.451316f
C21777 DVDD.n4445 VSS 0.451316f
C21778 DVDD.n4446 VSS 0.451316f
C21779 DVDD.n4447 VSS 0.451316f
C21780 DVDD.n4448 VSS 0.346009f
C21781 DVDD.n4449 VSS 0.301937f
C21782 DVDD.n4450 VSS 0.105095f
C21783 DVDD.n4451 VSS 0.240702f
C21784 DVDD.n4452 VSS 0.240702f
C21785 DVDD.n4453 VSS 0.240702f
C21786 DVDD.n4454 VSS 0.240702f
C21787 DVDD.n4455 VSS 0.192392f
C21788 DVDD.n4456 VSS 0.240702f
C21789 DVDD.n4457 VSS 0.240702f
C21790 DVDD.n4458 VSS 0.240702f
C21791 DVDD.n4459 VSS 0.120351f
C21792 DVDD.n4463 VSS 0.050859f
C21793 DVDD.n4464 VSS 0.033368f
C21794 DVDD.n4465 VSS 0.033368f
C21795 DVDD.n4466 VSS 0.131369f
C21796 DVDD.n4467 VSS 0.033368f
C21797 DVDD.n4468 VSS 0.131369f
C21798 DVDD.n4469 VSS 0.033368f
C21799 DVDD.n4470 VSS 0.225658f
C21800 DVDD.n4471 VSS 0.225658f
C21801 DVDD.n4472 VSS 0.225658f
C21802 DVDD.n4473 VSS 2.66633f
C21803 DVDD.n4474 VSS 0.033368f
C21804 DVDD.n4475 VSS 0.033368f
C21805 DVDD.n4476 VSS 0.033368f
C21806 DVDD.n4477 VSS 0.033368f
C21807 DVDD.n4478 VSS 0.033368f
C21808 DVDD.n4479 VSS 0.033368f
C21809 DVDD.n4480 VSS 0.033368f
C21810 DVDD.n4481 VSS 0.033368f
C21811 DVDD.n4482 VSS 0.033368f
C21812 DVDD.n4483 VSS 0.066735f
C21813 DVDD.n4484 VSS 0.066735f
C21814 DVDD.n4485 VSS 0.131369f
C21815 DVDD.n4486 VSS 0.066735f
C21816 DVDD.n4487 VSS 0.131369f
C21817 DVDD.n4488 VSS 0.066735f
C21818 DVDD.n4489 VSS 0.131369f
C21819 DVDD.n4490 VSS 0.066735f
C21820 DVDD.n4491 VSS 0.131369f
C21821 DVDD.n4492 VSS 0.066735f
C21822 DVDD.n4493 VSS 0.131369f
C21823 DVDD.n4494 VSS 0.066735f
C21824 DVDD.n4495 VSS 0.131369f
C21825 DVDD.n4496 VSS 0.066735f
C21826 DVDD.n4497 VSS 0.131369f
C21827 DVDD.n4498 VSS 0.066735f
C21828 DVDD.n4499 VSS 0.131369f
C21829 DVDD.n4500 VSS 0.066735f
C21830 DVDD.n4501 VSS 0.131369f
C21831 DVDD.n4502 VSS 0.066735f
C21832 DVDD.n4503 VSS 0.131369f
C21833 DVDD.n4504 VSS 0.066735f
C21834 DVDD.n4505 VSS 0.131369f
C21835 DVDD.n4506 VSS 0.066735f
C21836 DVDD.n4507 VSS 0.066735f
C21837 DVDD.n4508 VSS 0.197054f
C21838 DVDD.n4509 VSS 0.066735f
C21839 DVDD.n4510 VSS 0.026274f
C21840 DVDD.n4511 VSS 0.026274f
C21841 DVDD.n4512 VSS 0.030088f
C21842 DVDD.n4513 VSS 0.060175f
C21843 DVDD.n4514 VSS 0.059611f
C21844 DVDD.n4515 VSS 0.029028f
C21845 DVDD.n4516 VSS 0.217712f
C21846 DVDD.n4517 VSS 0.066735f
C21847 DVDD.n4518 VSS 0.066735f
C21848 DVDD.n4519 VSS 0.130242f
C21849 DVDD.n4520 VSS 0.033368f
C21850 DVDD.n4521 VSS 0.131369f
C21851 DVDD.n4522 VSS 0.033368f
C21852 DVDD.n4523 VSS 0.033368f
C21853 DVDD.n4524 VSS 0.033368f
C21854 DVDD.n4525 VSS 0.131369f
C21855 DVDD.n4526 VSS 0.131369f
C21856 DVDD.n4527 VSS 0.066735f
C21857 DVDD.n4528 VSS 0.225658f
C21858 DVDD.n4529 VSS 0.033368f
C21859 DVDD.n4530 VSS 0.033368f
C21860 DVDD.n4531 VSS 0.033368f
C21861 DVDD.n4532 VSS 0.033368f
C21862 DVDD.n4533 VSS 0.131369f
C21863 DVDD.n4534 VSS 0.033368f
C21864 DVDD.n4535 VSS 0.131369f
C21865 DVDD.n4536 VSS 0.131369f
C21866 DVDD.n4537 VSS 0.066735f
C21867 DVDD.n4538 VSS 0.131369f
C21868 DVDD.n4539 VSS 0.066735f
C21869 DVDD.n4540 VSS 0.131369f
C21870 DVDD.n4541 VSS 0.033368f
C21871 DVDD.n4542 VSS 0.105307f
C21872 DVDD.n4543 VSS 0.105307f
C21873 DVDD.n4544 VSS 0.105307f
C21874 DVDD.n4545 VSS 1.3091f
C21875 DVDD.n4546 VSS 0.033368f
C21876 DVDD.n4547 VSS 0.033368f
C21877 DVDD.n4548 VSS 0.033368f
C21878 DVDD.n4549 VSS 0.033368f
C21879 DVDD.n4550 VSS 0.033368f
C21880 DVDD.n4551 VSS 0.091958f
C21881 DVDD.n4552 VSS 0.033368f
C21882 DVDD.n4553 VSS 0.033368f
C21883 DVDD.n4554 VSS 0.033368f
C21884 DVDD.n4555 VSS 0.033368f
C21885 DVDD.n4556 VSS 0.033368f
C21886 DVDD.n4557 VSS 0.131369f
C21887 DVDD.n4558 VSS 0.066735f
C21888 DVDD.n4559 VSS 0.131369f
C21889 DVDD.n4560 VSS 0.066735f
C21890 DVDD.n4561 VSS 0.131369f
C21891 DVDD.n4562 VSS 0.15585f
C21892 DVDD.n4563 VSS 0.124509f
C21893 DVDD.n4564 VSS 0.114418f
C21894 DVDD.n4565 VSS 0.058124f
C21895 DVDD.n4566 VSS 0.114418f
C21896 DVDD.n4567 VSS 0.124509f
C21897 DVDD.n4568 VSS 0.925692f
C21898 DVDD.n4569 VSS 0.38847f
C21899 DVDD.n4570 VSS 0.105307f
C21900 DVDD.n4571 VSS 0.105307f
C21901 DVDD.n4572 VSS 0.033368f
C21902 DVDD.n4573 VSS 0.105307f
C21903 DVDD.n4574 VSS 0.187625f
C21904 DVDD.n4575 VSS 0.029062f
C21905 DVDD.n4576 VSS 0.029062f
C21906 DVDD.n4577 VSS 0.029062f
C21907 DVDD.n4578 VSS 0.029062f
C21908 DVDD.n4579 VSS 0.029062f
C21909 DVDD.n4580 VSS 0.210614f
C21910 DVDD.n4581 VSS 0.091958f
C21911 DVDD.n4582 VSS 0.210614f
C21912 DVDD.n4583 VSS 0.210614f
C21913 DVDD.n4584 VSS 0.210614f
C21914 DVDD.n4585 VSS 0.210614f
C21915 DVDD.n4586 VSS 0.210614f
C21916 DVDD.n4587 VSS 0.210614f
C21917 DVDD.n4588 VSS 0.210614f
C21918 DVDD.n4589 VSS 0.168343f
C21919 DVDD.n4590 VSS 0.210614f
C21920 DVDD.n4591 VSS 0.210614f
C21921 DVDD.n4592 VSS 0.210614f
C21922 DVDD.n4593 VSS 0.105307f
C21923 DVDD.n4600 VSS 0.187625f
C21924 DVDD.n4601 VSS 0.066735f
C21925 DVDD.n4602 VSS 0.066735f
C21926 DVDD.n4603 VSS 0.066735f
C21927 DVDD.n4604 VSS 0.066735f
C21928 DVDD.n4605 VSS 0.066735f
C21929 DVDD.n4606 VSS 0.210614f
C21930 DVDD.n4607 VSS 0.210614f
C21931 DVDD.n4608 VSS 0.210614f
C21932 DVDD.n4609 VSS 0.168343f
C21933 DVDD.n4610 VSS 0.210614f
C21934 DVDD.n4611 VSS 1.46014f
C21935 DVDD.n4612 VSS 0.210614f
C21936 DVDD.n4613 VSS 0.105307f
C21937 DVDD.n4614 VSS 0.65328f
C21938 DVDD.n4615 VSS 0.033368f
C21939 DVDD.n4616 VSS 0.033368f
C21940 DVDD.n4617 VSS 0.033368f
C21941 DVDD.n4618 VSS 0.033368f
C21942 DVDD.n4619 VSS 0.033368f
C21943 DVDD.n4620 VSS 0.033368f
C21944 DVDD.n4621 VSS 0.033368f
C21945 DVDD.n4622 VSS 0.033368f
C21946 DVDD.n4623 VSS 0.033368f
C21947 DVDD.n4624 VSS 0.033368f
C21948 DVDD.n4625 VSS 1.20359f
C21949 DVDD.n4626 VSS 0.066735f
C21950 DVDD.n4627 VSS 0.033368f
C21951 DVDD.n4628 VSS 0.431393f
C21952 DVDD.n4629 VSS 0.033368f
C21953 DVDD.n4630 VSS 0.131369f
C21954 DVDD.n4631 VSS 0.033368f
C21955 DVDD.n4632 VSS 0.131369f
C21956 DVDD.n4633 VSS 0.033368f
C21957 DVDD.n4634 VSS 0.131369f
C21958 DVDD.n4635 VSS 0.033368f
C21959 DVDD.n4636 VSS 0.131369f
C21960 DVDD.n4637 VSS 0.033368f
C21961 DVDD.n4638 VSS 0.131369f
C21962 DVDD.n4639 VSS 0.033368f
C21963 DVDD.n4640 VSS 0.131369f
C21964 DVDD.n4641 VSS 0.033368f
C21965 DVDD.n4642 VSS 0.131369f
C21966 DVDD.n4643 VSS 0.033368f
C21967 DVDD.n4644 VSS 0.131369f
C21968 DVDD.n4645 VSS 0.131369f
C21969 DVDD.n4646 VSS 0.131369f
C21970 DVDD.n4647 VSS 0.066735f
C21971 DVDD.n4648 VSS 0.066735f
C21972 DVDD.n4649 VSS 0.131369f
C21973 DVDD.n4650 VSS 0.066735f
C21974 DVDD.n4651 VSS 0.131369f
C21975 DVDD.n4652 VSS 0.066735f
C21976 DVDD.n4653 VSS 0.131369f
C21977 DVDD.n4654 VSS 0.066735f
C21978 DVDD.n4655 VSS 0.131369f
C21979 DVDD.n4656 VSS 0.066735f
C21980 DVDD.n4657 VSS 0.131369f
C21981 DVDD.n4658 VSS 0.066735f
C21982 DVDD.n4659 VSS 0.066735f
C21983 DVDD.n4660 VSS 0.131369f
C21984 DVDD.n4661 VSS 0.131369f
C21985 DVDD.n4662 VSS 0.131369f
C21986 DVDD.n4663 VSS 0.066735f
C21987 DVDD.n4664 VSS 0.066735f
C21988 DVDD.n4665 VSS 0.066735f
C21989 DVDD.n4666 VSS 0.131369f
C21990 DVDD.n4667 VSS 0.131369f
C21991 DVDD.n4668 VSS 0.131369f
C21992 DVDD.n4669 VSS 0.066735f
C21993 DVDD.n4670 VSS 0.066735f
C21994 DVDD.n4671 VSS 0.066735f
C21995 DVDD.n4672 VSS 0.131369f
C21996 DVDD.n4673 VSS 0.131369f
C21997 DVDD.n4674 VSS 0.131369f
C21998 DVDD.n4675 VSS 0.066735f
C21999 DVDD.n4676 VSS 0.066735f
C22000 DVDD.n4677 VSS 0.066735f
C22001 DVDD.n4678 VSS 0.131369f
C22002 DVDD.n4679 VSS 0.131369f
C22003 DVDD.n4680 VSS 0.131369f
C22004 DVDD.n4681 VSS 0.066735f
C22005 DVDD.n4682 VSS 0.066735f
C22006 DVDD.n4683 VSS 0.066735f
C22007 DVDD.n4684 VSS 0.131369f
C22008 DVDD.n4685 VSS 0.131369f
C22009 DVDD.n4686 VSS 0.131369f
C22010 DVDD.n4687 VSS 0.066735f
C22011 DVDD.n4688 VSS 0.066735f
C22012 DVDD.n4689 VSS 0.066735f
C22013 DVDD.n4690 VSS 0.131369f
C22014 DVDD.n4691 VSS 0.131369f
C22015 DVDD.n4692 VSS 0.131369f
C22016 DVDD.n4693 VSS 0.066735f
C22017 DVDD.n4694 VSS 0.26156f
C22018 DVDD.n4695 VSS 0.26156f
C22019 DVDD.n4696 VSS 0.066735f
C22020 DVDD.n4697 VSS 0.131369f
C22021 DVDD.n4698 VSS 0.131369f
C22022 DVDD.n4699 VSS 0.131369f
C22023 DVDD.n4700 VSS 0.066735f
C22024 DVDD.n4701 VSS 0.066735f
C22025 DVDD.n4702 VSS 0.066735f
C22026 DVDD.n4703 VSS 0.131369f
C22027 DVDD.n4704 VSS 0.131369f
C22028 DVDD.n4705 VSS 0.131369f
C22029 DVDD.n4706 VSS 0.063237f
C22030 DVDD.n4707 VSS 1.30905f
C22031 DVDD.n4708 VSS 0.407854f
C22032 DVDD.n4709 VSS 0.091958f
C22033 DVDD.n4710 VSS 0.091958f
C22034 DVDD.n4711 VSS 0.105307f
C22035 DVDD.n4712 VSS 0.033368f
C22036 DVDD.n4713 VSS 0.105307f
C22037 DVDD.n4714 VSS 0.091958f
C22038 DVDD.n4715 VSS 0.210614f
C22039 DVDD.n4716 VSS 0.210614f
C22040 DVDD.n4717 VSS 0.210614f
C22041 DVDD.n4718 VSS 0.210614f
C22042 DVDD.n4719 VSS 0.210614f
C22043 DVDD.n4720 VSS 0.210614f
C22044 DVDD.n4721 VSS 0.210614f
C22045 DVDD.n4722 VSS 0.210614f
C22046 DVDD.n4723 VSS 0.210614f
C22047 DVDD.n4724 VSS 0.210614f
C22048 DVDD.n4725 VSS 0.210614f
C22049 DVDD.n4726 VSS 0.210614f
C22050 DVDD.n4727 VSS 0.210614f
C22051 DVDD.n4728 VSS 0.091958f
C22052 DVDD.n4729 VSS 0.066735f
C22053 DVDD.n4730 VSS 0.066735f
C22054 DVDD.n4731 VSS 0.066735f
C22055 DVDD.n4732 VSS 0.066735f
C22056 DVDD.n4737 VSS 0.091958f
C22057 DVDD.n4738 VSS 0.105307f
C22058 DVDD.n4740 VSS 0.105307f
C22059 DVDD.n4741 VSS 0.105307f
C22060 DVDD.n4742 VSS 0.091958f
C22061 DVDD.n4747 VSS 0.066735f
C22062 DVDD.n4748 VSS 0.210614f
C22063 DVDD.n4749 VSS 0.210614f
C22064 DVDD.n4750 VSS 0.210614f
C22065 DVDD.n4751 VSS 0.210614f
C22066 DVDD.n4752 VSS 0.210614f
C22067 DVDD.n4753 VSS 0.210614f
C22068 DVDD.n4754 VSS 0.210614f
C22069 DVDD.n4755 VSS 0.210614f
C22070 DVDD.n4756 VSS 0.407854f
C22071 DVDD.n4757 VSS 0.091958f
C22072 DVDD.n4758 VSS 0.210614f
C22073 DVDD.n4759 VSS 0.091958f
C22074 DVDD.n4760 VSS 1.45939f
C22075 DVDD.n4761 VSS 0.210614f
C22076 DVDD.n4762 VSS 0.210614f
C22077 DVDD.n4763 VSS 0.210614f
C22078 DVDD.n4764 VSS 0.168343f
C22079 DVDD.n4765 VSS 0.210614f
C22080 DVDD.n4766 VSS 0.210614f
C22081 DVDD.n4767 VSS 0.210614f
C22082 DVDD.n4768 VSS 0.210614f
C22083 DVDD.n4769 VSS 0.210614f
C22084 DVDD.n4770 VSS 0.210614f
C22085 DVDD.n4771 VSS 0.210614f
C22086 DVDD.n4772 VSS 0.210614f
C22087 DVDD.n4773 VSS 0.187625f
C22088 DVDD.n4775 VSS 0.066735f
C22089 DVDD.n4776 VSS 0.066735f
C22090 DVDD.n4777 VSS 0.066735f
C22091 DVDD.n4778 VSS 0.066735f
C22092 DVDD.n4780 VSS 0.066735f
C22093 DVDD.n4782 VSS 0.066735f
C22094 DVDD.n4784 VSS 0.066735f
C22095 DVDD.n4786 VSS 0.066735f
C22096 DVDD.n4787 VSS 0.105307f
C22097 DVDD.n4788 VSS 0.091958f
C22098 DVDD.n4789 VSS 0.210614f
C22099 DVDD.n4790 VSS 0.091958f
C22100 DVDD.n4791 VSS 0.210614f
C22101 DVDD.n4792 VSS 0.210614f
C22102 DVDD.n4793 VSS 0.210614f
C22103 DVDD.n4794 VSS 0.210614f
C22104 DVDD.n4795 VSS 0.210614f
C22105 DVDD.n4796 VSS 0.210614f
C22106 DVDD.n4797 VSS 0.210614f
C22107 DVDD.n4798 VSS 0.210614f
C22108 DVDD.n4799 VSS 0.210614f
C22109 DVDD.n4800 VSS 0.210614f
C22110 DVDD.n4801 VSS 0.210614f
C22111 DVDD.n4802 VSS 0.210614f
C22112 DVDD.n4803 VSS 0.210614f
C22113 DVDD.n4804 VSS 0.210614f
C22114 DVDD.n4805 VSS 0.210614f
C22115 DVDD.n4806 VSS 0.210614f
C22116 DVDD.n4807 VSS 0.210614f
C22117 DVDD.n4808 VSS 0.210614f
C22118 DVDD.n4809 VSS 0.210614f
C22119 DVDD.n4810 VSS 0.210614f
C22120 DVDD.n4811 VSS 0.210614f
C22121 DVDD.n4812 VSS 0.210614f
C22122 DVDD.n4813 VSS 0.210614f
C22123 DVDD.n4814 VSS 0.210614f
C22124 DVDD.n4815 VSS 0.168343f
C22125 DVDD.n4816 VSS 0.105307f
C22126 DVDD.n4817 VSS 1.85245f
C22127 DVDD.n4818 VSS 1.85245f
C22128 DVDD.n4819 VSS 0.105307f
C22129 DVDD.n4820 VSS 0.871867f
C22130 DVDD.n4821 VSS 0.105307f
C22131 DVDD.n4822 VSS 0.091958f
C22132 DVDD.n4823 VSS 0.210614f
C22133 DVDD.n4824 VSS 0.210614f
C22134 DVDD.n4825 VSS 0.210614f
C22135 DVDD.n4826 VSS 0.210614f
C22136 DVDD.n4827 VSS 0.210614f
C22137 DVDD.n4828 VSS 0.210614f
C22138 DVDD.n4829 VSS 0.210614f
C22139 DVDD.n4830 VSS 0.210614f
C22140 DVDD.n4831 VSS 0.210614f
C22141 DVDD.n4832 VSS 0.210614f
C22142 DVDD.n4833 VSS 0.210614f
C22143 DVDD.n4834 VSS 0.210614f
C22144 DVDD.n4835 VSS 0.210614f
C22145 DVDD.n4836 VSS 0.210614f
C22146 DVDD.n4837 VSS 0.210614f
C22147 DVDD.n4838 VSS 0.210614f
C22148 DVDD.n4839 VSS 0.210614f
C22149 DVDD.n4840 VSS 0.210614f
C22150 DVDD.n4841 VSS 0.210614f
C22151 DVDD.n4842 VSS 0.210614f
C22152 DVDD.n4843 VSS 0.210614f
C22153 DVDD.n4844 VSS 0.210614f
C22154 DVDD.n4845 VSS 0.210614f
C22155 DVDD.n4846 VSS 0.210614f
C22156 DVDD.n4847 VSS 0.210614f
C22157 DVDD.n4848 VSS 0.210614f
C22158 DVDD.n4849 VSS 0.210614f
C22159 DVDD.n4850 VSS 0.210614f
C22160 DVDD.n4851 VSS 0.210614f
C22161 DVDD.n4852 VSS 0.210614f
C22162 DVDD.n4853 VSS 0.210614f
C22163 DVDD.n4854 VSS 0.210614f
C22164 DVDD.n4855 VSS 0.210614f
C22165 DVDD.n4856 VSS 0.210614f
C22166 DVDD.n4857 VSS 0.029062f
C22167 DVDD.n4858 VSS 0.029062f
C22168 DVDD.n4859 VSS 0.029062f
C22169 DVDD.n4860 VSS 0.029062f
C22170 DVDD.n4861 VSS 0.029062f
C22171 DVDD.n4862 VSS 0.091958f
C22172 DVDD.n4863 VSS 0.029062f
C22173 DVDD.n4864 VSS 0.029062f
C22174 DVDD.n4865 VSS 0.029062f
C22175 DVDD.n4866 VSS 0.029062f
C22176 DVDD.n4867 VSS 0.754582f
C22177 DVDD.n4868 VSS 0.032022f
C22178 DVDD.n4869 VSS 0.105307f
C22179 DVDD.n4870 VSS 0.114418f
C22180 DVDD.n4871 VSS 0.114418f
C22181 DVDD.n4872 VSS 0.058124f
C22182 DVDD.n4873 VSS 0.114418f
C22183 DVDD.n4874 VSS 0.058124f
C22184 DVDD.n4875 VSS 0.030408f
C22185 DVDD.n4876 VSS 0.114418f
C22186 DVDD.n4877 VSS 0.033368f
C22187 DVDD.n4878 VSS 0.38847f
C22188 DVDD.n4879 VSS 0.747408f
C22189 DVDD.t10 VSS 5.27557f
C22190 DVDD.n4881 VSS 0.058124f
C22191 DVDD.n4882 VSS 0.114418f
C22192 DVDD.n4883 VSS 0.058124f
C22193 DVDD.n4884 VSS 0.114418f
C22194 DVDD.n4885 VSS 0.058124f
C22195 DVDD.n4886 VSS 0.114418f
C22196 DVDD.n4887 VSS 0.058124f
C22197 DVDD.n4888 VSS 0.114418f
C22198 DVDD.n4889 VSS 0.058124f
C22199 DVDD.n4890 VSS 0.114418f
C22200 DVDD.n4891 VSS 0.058124f
C22201 DVDD.n4892 VSS 0.114418f
C22202 DVDD.n4893 VSS 0.058124f
C22203 DVDD.n4894 VSS 0.114418f
C22204 DVDD.n4895 VSS 0.058124f
C22205 DVDD.n4896 VSS 0.114418f
C22206 DVDD.n4897 VSS 0.058124f
C22207 DVDD.n4898 VSS 0.114418f
C22208 DVDD.n4899 VSS 0.114418f
C22209 DVDD.n4900 VSS 0.058124f
C22210 DVDD.t39 VSS 5.27557f
C22211 DVDD.n4902 VSS 0.15585f
C22212 DVDD.n4903 VSS 0.114418f
C22213 DVDD.n4904 VSS 0.058124f
C22214 DVDD.n4905 VSS 0.058124f
C22215 DVDD.n4906 VSS 0.114418f
C22216 DVDD.n4907 VSS 0.114418f
C22217 DVDD.n4908 VSS 0.114418f
C22218 DVDD.n4909 VSS 0.058124f
C22219 DVDD.n4910 VSS 0.058124f
C22220 DVDD.n4911 VSS 0.058124f
C22221 DVDD.n4912 VSS 0.114418f
C22222 DVDD.n4913 VSS 0.114418f
C22223 DVDD.n4914 VSS 0.114418f
C22224 DVDD.n4915 VSS 0.114418f
C22225 DVDD.n4916 VSS 0.032022f
C22226 DVDD.n4917 VSS 0.030408f
C22227 DVDD.n4918 VSS 0.114418f
C22228 DVDD.n4919 VSS 0.033368f
C22229 DVDD.n4920 VSS 0.114418f
C22230 DVDD.n4921 VSS 0.033368f
C22231 DVDD.n4922 VSS 0.114418f
C22232 DVDD.n4923 VSS 0.033368f
C22233 DVDD.n4924 VSS 0.114418f
C22234 DVDD.n4925 VSS 0.033368f
C22235 DVDD.n4926 VSS 0.114418f
C22236 DVDD.n4927 VSS 0.033368f
C22237 DVDD.n4928 VSS 0.114418f
C22238 DVDD.n4929 VSS 0.033368f
C22239 DVDD.n4930 VSS 0.114418f
C22240 DVDD.n4931 VSS 0.114418f
C22241 DVDD.n4932 VSS 0.030946f
C22242 DVDD.n4933 VSS 0.031484f
C22243 DVDD.n4934 VSS 0.114418f
C22244 DVDD.n4935 VSS 0.033368f
C22245 DVDD.n4936 VSS 0.114418f
C22246 DVDD.n4937 VSS 0.114418f
C22247 DVDD.n4938 VSS 0.051397f
C22248 DVDD.n4939 VSS 0.058124f
C22249 DVDD.n4940 VSS 0.058124f
C22250 DVDD.n4941 VSS 0.114418f
C22251 DVDD.n4942 VSS 0.114418f
C22252 DVDD.n4943 VSS 0.114418f
C22253 DVDD.n4944 VSS 0.058124f
C22254 DVDD.n4945 VSS 0.058124f
C22255 DVDD.n4946 VSS 0.058124f
C22256 DVDD.n4947 VSS 0.114418f
C22257 DVDD.n4948 VSS 0.114418f
C22258 DVDD.n4949 VSS 0.15585f
C22259 DVDD.n4950 VSS 0.277706f
C22260 DVDD.t15 VSS 5.27557f
C22261 DVDD.n4952 VSS 0.15585f
C22262 DVDD.n4953 VSS 0.277706f
C22263 DVDD.n4954 VSS 0.058124f
C22264 DVDD.n4955 VSS 0.058124f
C22265 DVDD.n4956 VSS 0.114418f
C22266 DVDD.n4957 VSS 0.114418f
C22267 DVDD.n4958 VSS 0.114418f
C22268 DVDD.n4959 VSS 0.058124f
C22269 DVDD.n4960 VSS 0.058124f
C22270 DVDD.n4961 VSS 0.058124f
C22271 DVDD.n4962 VSS 0.114418f
C22272 DVDD.n4963 VSS 0.114418f
C22273 DVDD.n4964 VSS 0.114418f
C22274 DVDD.n4965 VSS 0.058124f
C22275 DVDD.n4966 VSS 0.058124f
C22276 DVDD.n4967 VSS 0.058124f
C22277 DVDD.n4968 VSS 0.114418f
C22278 DVDD.n4969 VSS 0.114418f
C22279 DVDD.n4970 VSS 0.114418f
C22280 DVDD.n4971 VSS 0.058124f
C22281 DVDD.n4972 VSS 0.058124f
C22282 DVDD.n4973 VSS 0.058124f
C22283 DVDD.n4974 VSS 0.114418f
C22284 DVDD.n4975 VSS 0.114418f
C22285 DVDD.n4976 VSS 0.114418f
C22286 DVDD.n4977 VSS 0.058124f
C22287 DVDD.n4978 VSS 0.058124f
C22288 DVDD.n4979 VSS 0.058124f
C22289 DVDD.n4980 VSS 0.114418f
C22290 DVDD.n4981 VSS 0.114418f
C22291 DVDD.n4982 VSS 0.114418f
C22292 DVDD.n4983 VSS 0.058124f
C22293 DVDD.n4984 VSS 0.058124f
C22294 DVDD.n4985 VSS 0.058124f
C22295 DVDD.n4986 VSS 0.114418f
C22296 DVDD.n4987 VSS 0.114418f
C22297 DVDD.n4988 VSS 0.114418f
C22298 DVDD.n4989 VSS 0.058124f
C22299 DVDD.n4990 VSS 0.058124f
C22300 DVDD.n4991 VSS 0.058124f
C22301 DVDD.n4992 VSS 0.114418f
C22302 DVDD.n4993 VSS 0.114418f
C22303 DVDD.n4994 VSS 0.15585f
C22304 DVDD.n4995 VSS 0.277706f
C22305 DVDD.n4996 VSS 0.277706f
C22306 DVDD.n4997 VSS 0.15585f
C22307 DVDD.n4998 VSS 0.114418f
C22308 DVDD.n4999 VSS 0.114418f
C22309 DVDD.n5000 VSS 0.058124f
C22310 DVDD.n5001 VSS 0.058124f
C22311 DVDD.n5002 VSS 0.058124f
C22312 DVDD.n5003 VSS 0.114418f
C22313 DVDD.n5004 VSS 0.114418f
C22314 DVDD.n5005 VSS 0.114418f
C22315 DVDD.n5006 VSS 0.058124f
C22316 DVDD.n5007 VSS 0.058124f
C22317 DVDD.n5008 VSS 0.049783f
C22318 DVDD.n5009 VSS 0.114418f
C22319 DVDD.n5010 VSS 0.033368f
C22320 DVDD.n5011 VSS 0.114418f
C22321 DVDD.n5012 VSS 0.114418f
C22322 DVDD.n5013 VSS 0.033099f
C22323 DVDD.n5014 VSS 0.029331f
C22324 DVDD.n5015 VSS 0.114418f
C22325 DVDD.n5016 VSS 0.033368f
C22326 DVDD.n5017 VSS 0.114418f
C22327 DVDD.n5018 VSS 0.033368f
C22328 DVDD.n5019 VSS 0.114418f
C22329 DVDD.n5020 VSS 0.033368f
C22330 DVDD.n5021 VSS 0.114418f
C22331 DVDD.n5022 VSS 0.033368f
C22332 DVDD.n5023 VSS 0.114418f
C22333 DVDD.n5024 VSS 0.033368f
C22334 DVDD.n5025 VSS 0.114418f
C22335 DVDD.n5026 VSS 0.114418f
C22336 DVDD.n5027 VSS 0.033368f
C22337 DVDD.n5028 VSS 0.105307f
C22338 DVDD.n5029 VSS 0.091958f
C22339 DVDD.n5030 VSS 0.210614f
C22340 DVDD.n5031 VSS 0.210614f
C22341 DVDD.n5032 VSS 0.210614f
C22342 DVDD.n5033 VSS 0.091958f
C22343 DVDD.n5034 VSS 0.210614f
C22344 DVDD.n5035 VSS 0.210614f
C22345 DVDD.n5036 VSS 0.210614f
C22346 DVDD.n5037 VSS 0.210614f
C22347 DVDD.n5038 VSS 0.210614f
C22348 DVDD.n5039 VSS 0.210614f
C22349 DVDD.n5040 VSS 0.210614f
C22350 DVDD.n5041 VSS 0.210614f
C22351 DVDD.n5042 VSS 0.210614f
C22352 DVDD.n5043 VSS 0.210614f
C22353 DVDD.n5044 VSS 0.210614f
C22354 DVDD.n5045 VSS 0.210614f
C22355 DVDD.n5046 VSS 0.210614f
C22356 DVDD.n5047 VSS 0.210614f
C22357 DVDD.n5048 VSS 0.210614f
C22358 DVDD.n5049 VSS 0.210614f
C22359 DVDD.n5050 VSS 0.210614f
C22360 DVDD.n5051 VSS 0.210614f
C22361 DVDD.n5052 VSS 0.210614f
C22362 DVDD.n5053 VSS 0.210614f
C22363 DVDD.n5054 VSS 0.210614f
C22364 DVDD.n5055 VSS 0.210614f
C22365 DVDD.n5056 VSS 0.210614f
C22366 DVDD.n5057 VSS 0.210614f
C22367 DVDD.n5058 VSS 0.210614f
C22368 DVDD.n5059 VSS 0.210614f
C22369 DVDD.n5060 VSS 0.210614f
C22370 DVDD.n5061 VSS 0.210614f
C22371 DVDD.n5062 VSS 0.210614f
C22372 DVDD.n5063 VSS 0.210614f
C22373 DVDD.n5064 VSS 0.210614f
C22374 DVDD.n5065 VSS 0.210614f
C22375 DVDD.n5066 VSS 0.210614f
C22376 DVDD.n5067 VSS 0.210614f
C22377 DVDD.n5068 VSS 0.210614f
C22378 DVDD.n5069 VSS 0.210614f
C22379 DVDD.n5070 VSS 0.210614f
C22380 DVDD.n5071 VSS 0.210614f
C22381 DVDD.n5072 VSS 0.210614f
C22382 DVDD.n5073 VSS 0.210614f
C22383 DVDD.n5074 VSS 0.210614f
C22384 DVDD.n5075 VSS 0.210614f
C22385 DVDD.n5076 VSS 0.210614f
C22386 DVDD.n5077 VSS 0.210614f
C22387 DVDD.n5078 VSS 0.210614f
C22388 DVDD.n5079 VSS 0.168343f
C22389 DVDD.n5080 VSS 0.105307f
C22390 DVDD.n5081 VSS 0.029062f
C22391 DVDD.n5082 VSS 0.105307f
C22392 DVDD.n5083 VSS 0.187625f
C22393 DVDD.n5084 VSS 0.210614f
C22394 DVDD.n5085 VSS 0.210614f
C22395 DVDD.n5086 VSS 0.210614f
C22396 DVDD.n5087 VSS 0.210614f
C22397 DVDD.n5088 VSS 0.210614f
C22398 DVDD.n5089 VSS 0.210614f
C22399 DVDD.n5090 VSS 0.210614f
C22400 DVDD.n5091 VSS 0.210614f
C22401 DVDD.n5092 VSS 0.210614f
C22402 DVDD.n5093 VSS 0.210614f
C22403 DVDD.n5094 VSS 0.210614f
C22404 DVDD.n5095 VSS 0.210614f
C22405 DVDD.n5096 VSS 0.210614f
C22406 DVDD.n5097 VSS 0.210614f
C22407 DVDD.n5098 VSS 0.210614f
C22408 DVDD.n5099 VSS 0.210614f
C22409 DVDD.n5100 VSS 0.210614f
C22410 DVDD.n5101 VSS 0.210614f
C22411 DVDD.n5102 VSS 0.210614f
C22412 DVDD.n5103 VSS 0.210614f
C22413 DVDD.n5104 VSS 0.210614f
C22414 DVDD.n5105 VSS 0.210614f
C22415 DVDD.n5106 VSS 0.210614f
C22416 DVDD.n5107 VSS 0.168343f
C22417 DVDD.n5108 VSS 0.210614f
C22418 DVDD.n5109 VSS 0.091958f
C22419 DVDD.n5110 VSS 0.210614f
C22420 DVDD.n5111 VSS 0.210614f
C22421 DVDD.n5112 VSS 0.210614f
C22422 DVDD.n5113 VSS 0.210614f
C22423 DVDD.n5114 VSS 0.210614f
C22424 DVDD.n5115 VSS 0.091958f
C22425 DVDD.n5116 VSS 0.029062f
C22426 DVDD.n5117 VSS 0.029062f
C22427 DVDD.n5118 VSS 0.029062f
C22428 DVDD.n5119 VSS 0.029062f
C22429 DVDD.n5120 VSS 0.033368f
C22430 DVDD.n5121 VSS 0.114418f
C22431 DVDD.n5122 VSS 0.030408f
C22432 DVDD.n5123 VSS 0.032022f
C22433 DVDD.n5124 VSS 0.114418f
C22434 DVDD.n5125 VSS 0.033368f
C22435 DVDD.n5126 VSS 0.114418f
C22436 DVDD.n5127 VSS 0.033368f
C22437 DVDD.n5128 VSS 0.114418f
C22438 DVDD.n5129 VSS 0.033368f
C22439 DVDD.n5130 VSS 0.114418f
C22440 DVDD.n5131 VSS 0.033368f
C22441 DVDD.n5132 VSS 0.114418f
C22442 DVDD.n5133 VSS 0.114418f
C22443 DVDD.n5134 VSS 0.114418f
C22444 DVDD.n5135 VSS 0.058124f
C22445 DVDD.n5136 VSS 0.114418f
C22446 DVDD.n5137 VSS 0.114418f
C22447 DVDD.n5138 VSS 0.058124f
C22448 DVDD.n5139 VSS 0.058124f
C22449 DVDD.n5140 VSS 0.058124f
C22450 DVDD.n5141 VSS 0.114418f
C22451 DVDD.n5142 VSS 0.114418f
C22452 DVDD.n5143 VSS 0.114418f
C22453 DVDD.n5144 VSS 0.058124f
C22454 DVDD.n5145 VSS 0.058124f
C22455 DVDD.n5146 VSS 0.049783f
C22456 DVDD.n5147 VSS 0.114418f
C22457 DVDD.n5148 VSS 0.033368f
C22458 DVDD.n5149 VSS 0.114418f
C22459 DVDD.n5150 VSS 0.114418f
C22460 DVDD.n5151 VSS 0.033099f
C22461 DVDD.n5152 VSS 0.029331f
C22462 DVDD.n5153 VSS 0.114418f
C22463 DVDD.n5154 VSS 0.114418f
C22464 DVDD.n5155 VSS 0.033368f
C22465 DVDD.n5156 VSS 0.029062f
C22466 DVDD.n5157 VSS 0.105307f
C22467 DVDD.n5158 VSS 0.754582f
C22468 DVDD.n5159 VSS 0.747408f
C22469 DVDD.t1 VSS 5.27557f
C22470 DVDD.n5160 VSS 0.15585f
C22471 DVDD.n5161 VSS 0.277706f
C22472 DVDD.n5162 VSS 0.058124f
C22473 DVDD.n5163 VSS 0.114418f
C22474 DVDD.n5164 VSS 0.058124f
C22475 DVDD.n5165 VSS 0.114418f
C22476 DVDD.n5166 VSS 0.058124f
C22477 DVDD.n5167 VSS 0.114418f
C22478 DVDD.n5168 VSS 0.058124f
C22479 DVDD.n5169 VSS 0.114418f
C22480 DVDD.n5170 VSS 0.058124f
C22481 DVDD.n5171 VSS 0.114418f
C22482 DVDD.n5172 VSS 0.058124f
C22483 DVDD.n5173 VSS 0.114418f
C22484 DVDD.n5174 VSS 0.058124f
C22485 DVDD.n5175 VSS 0.114418f
C22486 DVDD.n5176 VSS 0.114418f
C22487 DVDD.n5177 VSS 0.058124f
C22488 DVDD.n5178 VSS 0.058124f
C22489 DVDD.n5179 VSS 0.058124f
C22490 DVDD.n5180 VSS 0.114418f
C22491 DVDD.n5181 VSS 0.114418f
C22492 DVDD.n5182 VSS 0.114418f
C22493 DVDD.n5183 VSS 0.058124f
C22494 DVDD.n5184 VSS 0.058124f
C22495 DVDD.n5185 VSS 0.058124f
C22496 DVDD.n5186 VSS 0.114418f
C22497 DVDD.n5187 VSS 0.114418f
C22498 DVDD.n5188 VSS 0.114418f
C22499 DVDD.n5189 VSS 0.058124f
C22500 DVDD.n5190 VSS 0.058124f
C22501 DVDD.n5191 VSS 0.058124f
C22502 DVDD.n5192 VSS 0.114418f
C22503 DVDD.n5193 VSS 0.114418f
C22504 DVDD.n5194 VSS 0.114418f
C22505 DVDD.n5195 VSS 0.058124f
C22506 DVDD.n5196 VSS 0.058124f
C22507 DVDD.n5197 VSS 0.058124f
C22508 DVDD.n5198 VSS 0.114418f
C22509 DVDD.n5199 VSS 0.114418f
C22510 DVDD.n5200 VSS 0.114418f
C22511 DVDD.n5201 VSS 0.058124f
C22512 DVDD.n5202 VSS 0.058124f
C22513 DVDD.n5203 VSS 0.058124f
C22514 DVDD.n5204 VSS 0.114418f
C22515 DVDD.n5205 VSS 0.114418f
C22516 DVDD.n5206 VSS 0.114418f
C22517 DVDD.n5207 VSS 0.058124f
C22518 DVDD.n5208 VSS 0.058124f
C22519 DVDD.n5209 VSS 0.058124f
C22520 DVDD.n5210 VSS 0.114418f
C22521 DVDD.n5211 VSS 0.114418f
C22522 DVDD.n5212 VSS 0.114418f
C22523 DVDD.n5213 VSS 0.058124f
C22524 DVDD.n5214 VSS 0.058124f
C22525 DVDD.n5215 VSS 0.277706f
C22526 DVDD.n5216 VSS 0.15585f
C22527 DVDD.t7 VSS 5.27557f
C22528 DVDD.n5217 VSS 0.124509f
C22529 DVDD.n5218 VSS 0.26156f
C22530 DVDD.n5219 VSS 0.26156f
C22531 DVDD.n5220 VSS 0.131369f
C22532 DVDD.n5221 VSS 0.066735f
C22533 DVDD.n5222 VSS 0.066735f
C22534 DVDD.n5223 VSS 0.066735f
C22535 DVDD.n5224 VSS 0.131369f
C22536 DVDD.n5225 VSS 0.131369f
C22537 DVDD.n5226 VSS 0.131369f
C22538 DVDD.n5227 VSS 0.066735f
C22539 DVDD.n5228 VSS 0.066735f
C22540 DVDD.n5229 VSS 0.064852f
C22541 DVDD.n5230 VSS 0.131369f
C22542 DVDD.n5231 VSS 0.033368f
C22543 DVDD.n5232 VSS 0.131369f
C22544 DVDD.n5233 VSS 0.033368f
C22545 DVDD.n5234 VSS 0.131369f
C22546 DVDD.n5235 VSS 0.033368f
C22547 DVDD.n5236 VSS 0.131369f
C22548 DVDD.n5237 VSS 0.033368f
C22549 DVDD.n5238 VSS 0.131369f
C22550 DVDD.n5239 VSS 0.033368f
C22551 DVDD.n5240 VSS 0.131369f
C22552 DVDD.n5241 VSS 0.033368f
C22553 DVDD.n5242 VSS 0.131369f
C22554 DVDD.n5243 VSS 0.033368f
C22555 DVDD.n5244 VSS 0.131369f
C22556 DVDD.n5245 VSS 0.131369f
C22557 DVDD.n5246 VSS 0.131369f
C22558 DVDD.n5247 VSS 0.033368f
C22559 DVDD.n5248 VSS 0.033368f
C22560 DVDD.n5249 VSS 1.20429f
C22561 DVDD.n5250 VSS 0.033368f
C22562 DVDD.n5251 VSS 0.035251f
C22563 DVDD.n5252 VSS 0.131369f
C22564 DVDD.n5253 VSS 0.131369f
C22565 DVDD.n5254 VSS 0.131369f
C22566 DVDD.n5255 VSS 0.066735f
C22567 DVDD.n5256 VSS 0.066735f
C22568 DVDD.n5257 VSS 0.066735f
C22569 DVDD.n5258 VSS 0.131369f
C22570 DVDD.n5259 VSS 0.131369f
C22571 DVDD.n5260 VSS 0.131369f
C22572 DVDD.n5261 VSS 0.066735f
C22573 DVDD.n5262 VSS 0.26156f
C22574 DVDD.n5263 VSS 0.063775f
C22575 DVDD.n5264 VSS 0.26156f
C22576 DVDD.n5265 VSS 0.124509f
C22577 DVDD.t33 VSS 5.27557f
C22578 DVDD.n5266 VSS 0.124509f
C22579 DVDD.n5267 VSS 0.096874f
C22580 DVDD.n5268 VSS 0.124053f
C22581 DVDD.n5269 VSS 0.225658f
C22582 DVDD.n5270 VSS 0.130242f
C22583 DVDD.n5271 VSS 0.066735f
C22584 DVDD.n5272 VSS 0.204999f
C22585 DVDD.n5273 VSS 0.066735f
C22586 DVDD.n5274 VSS 0.027333f
C22587 DVDD.n5275 VSS 0.026274f
C22588 DVDD.n5276 VSS 0.060175f
C22589 DVDD.n5277 VSS 0.057655f
C22590 DVDD.n5278 VSS 0.170687f
C22591 DVDD.n5279 VSS 0.060175f
C22592 DVDD.n5280 VSS 0.060175f
C22593 DVDD.n5281 VSS 0.026274f
C22594 DVDD.n5282 VSS 0.030088f
C22595 DVDD.n5283 VSS 0.066735f
C22596 DVDD.n5284 VSS 0.225658f
C22597 DVDD.n5285 VSS 0.066735f
C22598 DVDD.n5286 VSS 0.066735f
C22599 DVDD.n5287 VSS 0.225658f
C22600 DVDD.n5288 VSS 0.037404f
C22601 DVDD.n5289 VSS 0.033368f
C22602 DVDD.n5290 VSS 0.033368f
C22603 DVDD.n5291 VSS 0.033368f
C22604 DVDD.n5292 VSS 0.131369f
C22605 DVDD.n5293 VSS 0.033368f
C22606 DVDD.n5294 VSS 0.131369f
C22607 DVDD.n5295 VSS 0.131369f
C22608 DVDD.n5296 VSS 0.033368f
C22609 DVDD.n5297 VSS 0.451316f
C22610 DVDD.n5298 VSS 0.451316f
C22611 DVDD.n5299 VSS 1.30659f
C22612 DVDD.n5300 VSS 0.451316f
C22613 DVDD.n5301 VSS 0.451316f
C22614 DVDD.n5302 VSS 0.197054f
C22615 DVDD.n5303 VSS 0.225658f
C22616 DVDD.n5304 VSS 0.033368f
C22617 DVDD.n5305 VSS 0.033368f
C22618 DVDD.n5306 VSS 0.033368f
C22619 DVDD.n5307 VSS 0.033368f
C22620 DVDD.n5308 VSS 0.131369f
C22621 DVDD.n5309 VSS 0.037404f
C22622 DVDD.n5310 VSS 0.131369f
C22623 DVDD.n5311 VSS 0.131369f
C22624 DVDD.n5312 VSS 0.131369f
C22625 DVDD.n5313 VSS 0.066735f
C22626 DVDD.n5314 VSS 0.066735f
C22627 DVDD.n5315 VSS 0.066735f
C22628 DVDD.n5316 VSS 0.131369f
C22629 DVDD.n5317 VSS 0.131369f
C22630 DVDD.n5318 VSS 0.131369f
C22631 DVDD.n5319 VSS 0.066735f
C22632 DVDD.n5320 VSS 0.066735f
C22633 DVDD.n5321 VSS 0.066735f
C22634 DVDD.n5322 VSS 0.131369f
C22635 DVDD.n5323 VSS 0.131369f
C22636 DVDD.n5324 VSS 0.131369f
C22637 DVDD.n5325 VSS 0.066735f
C22638 DVDD.n5326 VSS 0.066735f
C22639 DVDD.n5327 VSS 0.066735f
C22640 DVDD.n5328 VSS 0.131369f
C22641 DVDD.n5329 VSS 0.131369f
C22642 DVDD.n5330 VSS 0.131369f
C22643 DVDD.n5331 VSS 0.066735f
C22644 DVDD.n5332 VSS 0.066735f
C22645 DVDD.n5333 VSS 0.066735f
C22646 DVDD.n5334 VSS 0.131369f
C22647 DVDD.n5335 VSS 0.131369f
C22648 DVDD.n5336 VSS 0.131369f
C22649 DVDD.n5337 VSS 0.066735f
C22650 DVDD.n5338 VSS 0.26156f
C22651 DVDD.n5339 VSS 0.26156f
C22652 DVDD.n5340 VSS 0.066735f
C22653 DVDD.n5341 VSS 0.066735f
C22654 DVDD.n5342 VSS 0.131369f
C22655 DVDD.n5343 VSS 0.131369f
C22656 DVDD.n5344 VSS 0.131369f
C22657 DVDD.n5345 VSS 0.066735f
C22658 DVDD.n5346 VSS 0.066735f
C22659 DVDD.n5347 VSS 0.066735f
C22660 DVDD.n5348 VSS 0.131369f
C22661 DVDD.n5349 VSS 0.131369f
C22662 DVDD.n5350 VSS 0.131369f
C22663 DVDD.n5351 VSS 0.066735f
C22664 DVDD.n5352 VSS 0.066735f
C22665 DVDD.n5353 VSS 0.066735f
C22666 DVDD.n5354 VSS 0.131369f
C22667 DVDD.n5355 VSS 0.131369f
C22668 DVDD.n5356 VSS 0.131369f
C22669 DVDD.n5357 VSS 0.066735f
C22670 DVDD.n5358 VSS 0.066735f
C22671 DVDD.n5359 VSS 0.066735f
C22672 DVDD.n5360 VSS 0.131369f
C22673 DVDD.n5361 VSS 0.131369f
C22674 DVDD.n5362 VSS 0.131369f
C22675 DVDD.n5363 VSS 0.066735f
C22676 DVDD.n5364 VSS 0.066735f
C22677 DVDD.n5365 VSS 0.066735f
C22678 DVDD.n5366 VSS 0.131369f
C22679 DVDD.n5367 VSS 0.131369f
C22680 DVDD.n5368 VSS 0.131369f
C22681 DVDD.n5369 VSS 0.066735f
C22682 DVDD.n5370 VSS 0.066735f
C22683 DVDD.n5371 VSS 0.066735f
C22684 DVDD.n5372 VSS 0.131369f
C22685 DVDD.n5373 VSS 0.131369f
C22686 DVDD.n5374 VSS 0.131369f
C22687 DVDD.n5375 VSS 0.066735f
C22688 DVDD.n5376 VSS 0.150424f
C22689 DVDD.n5377 VSS 0.150424f
C22690 DVDD.n5378 VSS 3.15709f
C22691 DVDD.n5379 VSS 0.451316f
C22692 DVDD.n5380 VSS 0.451316f
C22693 DVDD.n5381 VSS 0.451316f
C22694 DVDD.n5382 VSS 0.451316f
C22695 DVDD.n5383 VSS 0.451316f
C22696 DVDD.n5384 VSS 0.451316f
C22697 DVDD.n5385 VSS 0.451316f
C22698 DVDD.n5386 VSS 0.451316f
C22699 DVDD.n5387 VSS 0.451316f
C22700 DVDD.n5388 VSS 0.301937f
C22701 DVDD.n5389 VSS 0.451316f
C22702 DVDD.n5400 VSS 0.225658f
C22703 DVDD.n5401 VSS 0.197054f
C22704 DVDD.n5402 VSS 0.451316f
C22705 DVDD.n5403 VSS 0.451316f
C22706 DVDD.n5404 VSS 0.451316f
C22707 DVDD.n5405 VSS 0.451316f
C22708 DVDD.n5406 VSS 0.451316f
C22709 DVDD.n5407 VSS 0.451316f
C22710 DVDD.n5408 VSS 0.451316f
C22711 DVDD.n5409 VSS 0.360735f
C22712 DVDD.n5410 VSS 0.451316f
C22713 DVDD.n5411 VSS 0.197054f
C22714 DVDD.n5412 VSS 0.451316f
C22715 DVDD.n5413 VSS 0.197054f
C22716 DVDD.n5414 VSS 0.451316f
C22717 DVDD.n5415 VSS 0.930088f
C22718 DVDD.n5416 VSS 0.197054f
C22719 DVDD.n5419 VSS 0.066735f
C22720 DVDD.n5421 VSS 0.033368f
C22721 DVDD.n5422 VSS 0.044401f
C22722 DVDD.n5423 VSS 0.033368f
C22723 DVDD.n5424 VSS 0.033368f
C22724 DVDD.n5425 VSS 0.033368f
C22725 DVDD.n5426 VSS 0.033368f
C22726 DVDD.n5427 VSS 0.033368f
C22727 DVDD.n5428 VSS 0.033368f
C22728 DVDD.n5429 VSS 0.033368f
C22729 DVDD.n5430 VSS 0.033368f
C22730 DVDD.n5431 VSS 0.033368f
C22731 DVDD.n5432 VSS 0.131369f
C22732 DVDD.n5433 VSS 0.033368f
C22733 DVDD.n5434 VSS 0.131369f
C22734 DVDD.n5435 VSS 0.033368f
C22735 DVDD.n5436 VSS 0.131369f
C22736 DVDD.n5437 VSS 0.033368f
C22737 DVDD.n5438 VSS 0.131369f
C22738 DVDD.n5439 VSS 0.033368f
C22739 DVDD.n5440 VSS 0.131369f
C22740 DVDD.n5441 VSS 0.033368f
C22741 DVDD.n5442 VSS 0.131369f
C22742 DVDD.n5443 VSS 0.033368f
C22743 DVDD.n5444 VSS 0.131369f
C22744 DVDD.n5445 VSS 0.033368f
C22745 DVDD.n5446 VSS 0.131369f
C22746 DVDD.n5447 VSS 0.033368f
C22747 DVDD.n5448 VSS 0.131369f
C22748 DVDD.n5449 VSS 0.033368f
C22749 DVDD.n5450 VSS 0.131369f
C22750 DVDD.n5451 VSS 0.033368f
C22751 DVDD.n5452 VSS 0.131369f
C22752 DVDD.n5453 VSS 0.033368f
C22753 DVDD.n5454 VSS 0.131369f
C22754 DVDD.n5455 VSS 0.033368f
C22755 DVDD.n5456 VSS 0.131369f
C22756 DVDD.n5457 VSS 0.033368f
C22757 DVDD.n5458 VSS 0.131369f
C22758 DVDD.n5459 VSS 0.033368f
C22759 DVDD.n5460 VSS 0.131369f
C22760 DVDD.n5461 VSS 0.033368f
C22761 DVDD.n5462 VSS 0.131369f
C22762 DVDD.n5463 VSS 0.131369f
C22763 DVDD.n5464 VSS 0.033368f
C22764 DVDD.n5465 VSS 0.033368f
C22765 DVDD.n5466 VSS 2.63355f
C22766 DVDD.n5467 VSS 0.033368f
C22767 DVDD.n5468 VSS 0.033368f
C22768 DVDD.n5469 VSS 0.131369f
C22769 DVDD.n5470 VSS 0.131369f
C22770 DVDD.n5471 VSS 0.044401f
C22771 DVDD.n5472 VSS 0.066735f
C22772 DVDD.n5473 VSS 0.050859f
C22773 DVDD.n5474 VSS 0.131369f
C22774 DVDD.n5475 VSS 0.033368f
C22775 DVDD.n5476 VSS 0.131369f
C22776 DVDD.n5477 VSS 0.131369f
C22777 DVDD.n5478 VSS 0.033368f
C22778 DVDD.n5479 VSS 0.033368f
C22779 DVDD.n5480 VSS 0.033368f
C22780 DVDD.n5481 VSS 0.033368f
C22781 DVDD.n5482 VSS 0.105095f
C22782 DVDD.n5483 VSS 0.120351f
C22783 DVDD.n5484 VSS 0.066735f
C22784 DVDD.n5485 VSS 0.131369f
C22785 DVDD.n5486 VSS 0.066735f
C22786 DVDD.n5487 VSS 0.131369f
C22787 DVDD.n5488 VSS 0.066735f
C22788 DVDD.n5489 VSS 0.131369f
C22789 DVDD.n5490 VSS 0.066735f
C22790 DVDD.n5491 VSS 0.131369f
C22791 DVDD.n5492 VSS 0.225658f
C22792 DVDD.n5493 VSS 0.225658f
C22793 DVDD.n5494 VSS 0.033368f
C22794 DVDD.n5495 VSS 0.225658f
C22795 DVDD.n5496 VSS 2.66633f
C22796 DVDD.n5497 VSS 0.033368f
C22797 DVDD.n5498 VSS 0.033368f
C22798 DVDD.n5499 VSS 0.033368f
C22799 DVDD.n5500 VSS 0.033368f
C22800 DVDD.n5501 VSS 0.066735f
C22801 DVDD.n5502 VSS 0.066735f
C22802 DVDD.n5503 VSS 0.066735f
C22803 DVDD.n5504 VSS 0.033368f
C22804 DVDD.n5505 VSS 0.033368f
C22805 DVDD.n5506 VSS 0.033368f
C22806 DVDD.n5507 VSS 0.033368f
C22807 DVDD.n5508 VSS 3.15709f
C22808 DVDD.n5509 VSS 0.451316f
C22809 DVDD.n5510 VSS 0.451316f
C22810 DVDD.n5511 VSS 0.451316f
C22811 DVDD.n5512 VSS 0.451316f
C22812 DVDD.n5513 VSS 0.451316f
C22813 DVDD.n5514 VSS 0.451316f
C22814 DVDD.n5515 VSS 0.451316f
C22815 DVDD.n5516 VSS 0.451316f
C22816 DVDD.n5517 VSS 0.451316f
C22817 DVDD.n5518 VSS 0.451316f
C22818 DVDD.n5519 VSS 0.451316f
C22819 DVDD.n5520 VSS 0.451316f
C22820 DVDD.n5521 VSS 0.451316f
C22821 DVDD.n5522 VSS 0.451316f
C22822 DVDD.n5523 VSS 0.360735f
C22823 DVDD.n5524 VSS 0.451316f
C22824 DVDD.n5525 VSS 0.197054f
C22825 DVDD.n5526 VSS 0.451316f
C22826 DVDD.n5527 VSS 0.197054f
C22827 DVDD.n5528 VSS 0.451316f
C22828 DVDD.n5529 VSS 0.930088f
C22829 DVDD.n5530 VSS 0.197054f
C22830 DVDD.n5531 VSS 0.033368f
C22831 DVDD.n5532 VSS 0.033368f
C22832 DVDD.n5533 VSS 0.033368f
C22833 DVDD.n5534 VSS 0.033368f
C22834 DVDD.n5535 VSS 0.131369f
C22835 DVDD.n5536 VSS 0.033368f
C22836 DVDD.n5537 VSS 0.131369f
C22837 DVDD.n5538 VSS 0.033368f
C22838 DVDD.n5539 VSS 0.131369f
C22839 DVDD.n5540 VSS 0.033368f
C22840 DVDD.n5541 VSS 0.131369f
C22841 DVDD.n5542 VSS 0.033368f
C22842 DVDD.n5543 VSS 0.131369f
C22843 DVDD.n5544 VSS 0.033368f
C22844 DVDD.n5545 VSS 0.131369f
C22845 DVDD.n5546 VSS 0.131369f
C22846 DVDD.n5547 VSS 0.131369f
C22847 DVDD.n5548 VSS 0.033368f
C22848 DVDD.n5549 VSS 0.033368f
C22849 DVDD.n5550 VSS 0.033368f
C22850 DVDD.n5552 VSS 0.048168f
C22851 DVDD.n5555 VSS 0.066735f
C22852 DVDD.n5558 VSS 0.066735f
C22853 DVDD.n5560 VSS 0.033368f
C22854 DVDD.n5561 VSS 0.046553f
C22855 DVDD.n5562 VSS 0.033368f
C22856 DVDD.n5563 VSS 0.033368f
C22857 DVDD.n5564 VSS 0.033368f
C22858 DVDD.n5565 VSS 0.033368f
C22859 DVDD.n5566 VSS 0.066735f
C22860 DVDD.n5567 VSS 0.033368f
C22861 DVDD.n5568 VSS 0.131369f
C22862 DVDD.n5569 VSS 0.033368f
C22863 DVDD.n5570 VSS 0.131369f
C22864 DVDD.n5571 VSS 0.033368f
C22865 DVDD.n5572 VSS 0.131369f
C22866 DVDD.n5573 VSS 0.033368f
C22867 DVDD.n5574 VSS 0.131369f
C22868 DVDD.n5575 VSS 0.033368f
C22869 DVDD.n5576 VSS 0.131369f
C22870 DVDD.n5577 VSS 0.033368f
C22871 DVDD.n5578 VSS 0.131369f
C22872 DVDD.n5579 VSS 0.131369f
C22873 DVDD.n5580 VSS 0.033368f
C22874 DVDD.n5581 VSS 0.131369f
C22875 DVDD.n5582 VSS 0.033368f
C22876 DVDD.n5583 VSS 0.131369f
C22877 DVDD.n5584 VSS 0.033368f
C22878 DVDD.n5585 VSS 0.131369f
C22879 DVDD.n5586 VSS 0.033368f
C22880 DVDD.n5587 VSS 0.131369f
C22881 DVDD.n5588 VSS 0.033368f
C22882 DVDD.n5589 VSS 0.131369f
C22883 DVDD.n5590 VSS 0.033368f
C22884 DVDD.n5591 VSS 0.131369f
C22885 DVDD.n5592 VSS 0.033368f
C22886 DVDD.n5593 VSS 0.131369f
C22887 DVDD.n5594 VSS 0.033368f
C22888 DVDD.n5595 VSS 0.131369f
C22889 DVDD.n5596 VSS 0.033368f
C22890 DVDD.n5597 VSS 0.131369f
C22891 DVDD.n5598 VSS 0.033368f
C22892 DVDD.n5599 VSS 0.131369f
C22893 DVDD.n5600 VSS 0.033368f
C22894 DVDD.n5601 VSS 0.131369f
C22895 DVDD.n5602 VSS 0.033368f
C22896 DVDD.n5603 VSS 0.131369f
C22897 DVDD.n5604 VSS 0.033368f
C22898 DVDD.n5605 VSS 0.131369f
C22899 DVDD.n5606 VSS 0.033368f
C22900 DVDD.n5607 VSS 0.131369f
C22901 DVDD.n5608 VSS 0.047092f
C22902 DVDD.n5609 VSS 0.131369f
C22903 DVDD.n5610 VSS 0.131369f
C22904 DVDD.n5611 VSS 0.131369f
C22905 DVDD.n5612 VSS 0.046553f
C22906 DVDD.n5613 VSS 0.033368f
C22907 DVDD.n5614 VSS 2.63355f
C22908 DVDD.n5615 VSS 0.033368f
C22909 DVDD.n5616 VSS 0.048168f
C22910 DVDD.n5617 VSS 0.066735f
C22911 DVDD.n5618 VSS 0.131369f
C22912 DVDD.n5619 VSS 0.131369f
C22913 DVDD.n5620 VSS 0.131369f
C22914 DVDD.n5621 VSS 0.066735f
C22915 DVDD.n5622 VSS 0.066735f
C22916 DVDD.n5623 VSS 0.066735f
C22917 DVDD.n5624 VSS 0.131369f
C22918 DVDD.n5625 VSS 0.131369f
C22919 DVDD.n5626 VSS 0.131369f
C22920 DVDD.n5627 VSS 0.066735f
C22921 DVDD.n5628 VSS 0.066735f
C22922 DVDD.n5629 VSS 0.066735f
C22923 DVDD.n5630 VSS 0.131369f
C22924 DVDD.n5631 VSS 0.131369f
C22925 DVDD.n5632 VSS 0.131369f
C22926 DVDD.n5633 VSS 0.066735f
C22927 DVDD.n5634 VSS 0.066735f
C22928 DVDD.n5635 VSS 0.066735f
C22929 DVDD.n5636 VSS 0.131369f
C22930 DVDD.n5637 VSS 0.131369f
C22931 DVDD.n5638 VSS 0.131369f
C22932 DVDD.n5639 VSS 0.043862f
C22933 DVDD.n5640 VSS 1.17574f
C22934 DVDD.n5641 VSS 0.043862f
C22935 DVDD.n5642 VSS 0.066735f
C22936 DVDD.n5643 VSS 0.066735f
C22937 DVDD.n5644 VSS 0.353796f
C22938 DVDD.n5645 VSS 0.556696f
C22939 DVDD.n5646 VSS 0.557897f
C22940 DVDD.n5647 VSS 1.25096f
C22941 DVDD.n5648 VSS 0.147472f
C22942 DVDD.n5649 VSS 0.147472f
C22943 DVDD.n5650 VSS 0.105095f
C22944 DVDD.n5652 VSS 0.066735f
C22945 DVDD.n5654 VSS 0.066735f
C22946 DVDD.n5656 VSS 0.066735f
C22947 DVDD.n5657 VSS 0.027121f
C22948 DVDD.n5658 VSS 0.033368f
C22949 DVDD.n5659 VSS 0.120351f
C22950 DVDD.n5660 VSS 0.105095f
C22951 DVDD.n5661 VSS 0.240702f
C22952 DVDD.n5662 VSS 0.240702f
C22953 DVDD.n5663 VSS 0.240702f
C22954 DVDD.n5664 VSS 0.240702f
C22955 DVDD.n5665 VSS 0.240702f
C22956 DVDD.n5666 VSS 0.240702f
C22957 DVDD.n5667 VSS 0.240702f
C22958 DVDD.n5668 VSS 0.240702f
C22959 DVDD.n5669 VSS 0.240702f
C22960 DVDD.n5670 VSS 0.240702f
C22961 DVDD.n5671 VSS 0.240702f
C22962 DVDD.n5672 VSS 0.240702f
C22963 DVDD.n5673 VSS 0.240702f
C22964 DVDD.n5674 VSS 0.240702f
C22965 DVDD.n5675 VSS 0.161033f
C22966 DVDD.n5676 VSS 0.182751f
C22967 DVDD.n5677 VSS 0.138891f
C22968 DVDD.n5678 VSS 0.097467f
C22969 DVDD.n5679 VSS 0.161033f
C22970 DVDD.n5680 VSS 0.240702f
C22971 DVDD.n5681 VSS 0.20002f
C22972 DVDD.n5682 VSS 0.240702f
C22973 DVDD.n5683 VSS 0.240702f
C22974 DVDD.n5684 VSS 0.240702f
C22975 DVDD.n5685 VSS 0.240702f
C22976 DVDD.n5686 VSS 0.240702f
C22977 DVDD.n5687 VSS 0.240702f
C22978 DVDD.n5688 VSS 0.240702f
C22979 DVDD.n5689 VSS 0.105095f
C22980 DVDD.n5690 VSS 0.228836f
C22981 DVDD.n5691 VSS 0.214428f
C22982 DVDD.n5692 VSS 0.240702f
C22983 DVDD.n5693 VSS 0.240702f
C22984 DVDD.n5694 VSS 0.240702f
C22985 DVDD.n5695 VSS 0.240702f
C22986 DVDD.n5696 VSS 0.240702f
C22987 DVDD.n5697 VSS 0.240702f
C22988 DVDD.n5698 VSS 0.240702f
C22989 DVDD.n5699 VSS 0.240702f
C22990 DVDD.n5700 VSS 0.240702f
C22991 DVDD.n5701 VSS 0.240702f
C22992 DVDD.n5702 VSS 0.240702f
C22993 DVDD.n5703 VSS 0.240702f
C22994 DVDD.n5704 VSS 0.240702f
C22995 DVDD.n5705 VSS 0.240702f
C22996 DVDD.n5706 VSS 0.240702f
C22997 DVDD.n5707 VSS 0.192392f
C22998 DVDD.n5708 VSS 0.20002f
C22999 DVDD.n5709 VSS 0.346009f
C23000 DVDD.n5710 VSS 0.360735f
C23001 DVDD.n5711 VSS 0.375037f
C23002 DVDD.n5712 VSS 0.375037f
C23003 DVDD.n5713 VSS 0.451316f
C23004 DVDD.n5714 VSS 0.451316f
C23005 DVDD.n5715 VSS 0.451316f
C23006 DVDD.n5716 VSS 0.451316f
C23007 DVDD.n5717 VSS 0.451316f
C23008 DVDD.n5718 VSS 0.451316f
C23009 DVDD.n5719 VSS 0.451316f
C23010 DVDD.n5720 VSS 0.451316f
C23011 DVDD.n5721 VSS 0.451316f
C23012 DVDD.n5722 VSS 0.451316f
C23013 DVDD.n5723 VSS 0.451316f
C23014 DVDD.n5724 VSS 0.451316f
C23015 DVDD.n5725 VSS 0.451316f
C23016 DVDD.n5726 VSS 0.402053f
C23017 DVDD.n5727 VSS 0.451316f
C23018 DVDD.n5728 VSS 0.451316f
C23019 DVDD.n5729 VSS 0.451316f
C23020 DVDD.n5730 VSS 0.451316f
C23021 DVDD.n5731 VSS 0.197054f
C23022 DVDD.n5732 VSS 0.451316f
C23023 DVDD.n5733 VSS 0.451316f
C23024 DVDD.n5734 VSS 0.451316f
C23025 DVDD.n5735 VSS 0.451316f
C23026 DVDD.n5736 VSS 0.451316f
C23027 DVDD.n5737 VSS 0.451316f
C23028 DVDD.n5738 VSS 0.451316f
C23029 DVDD.n5739 VSS 0.451316f
C23030 DVDD.n5740 VSS 0.451316f
C23031 DVDD.n5741 VSS 0.451316f
C23032 DVDD.n5742 VSS 0.451316f
C23033 DVDD.n5743 VSS 0.451316f
C23034 DVDD.n5744 VSS 0.451316f
C23035 DVDD.n5745 VSS 0.451316f
C23036 DVDD.n5746 VSS 0.451316f
C23037 DVDD.n5747 VSS 0.451316f
C23038 DVDD.n5748 VSS 0.451316f
C23039 DVDD.n5749 VSS 0.451316f
C23040 DVDD.n5750 VSS 0.451316f
C23041 DVDD.n5751 VSS 0.451316f
C23042 DVDD.n5752 VSS 0.451316f
C23043 DVDD.n5753 VSS 0.451316f
C23044 DVDD.n5754 VSS 0.451316f
C23045 DVDD.n5755 VSS 0.451316f
C23046 DVDD.n5756 VSS 0.289224f
C23047 DVDD.n5757 VSS 0.289224f
C23048 DVDD.n5758 VSS 0.338487f
C23049 DVDD.n5759 VSS 0.346009f
C23050 DVDD.n5760 VSS 0.054088f
C23051 DVDD.n5761 VSS 0.066735f
C23052 DVDD.n5762 VSS 0.066735f
C23053 DVDD.n5763 VSS 0.061085f
C23054 DVDD.n5764 VSS 0.029062f
C23055 DVDD.n5765 VSS 0.105095f
C23056 DVDD.n5766 VSS 0.029062f
C23057 DVDD.n5767 VSS 0.033368f
C23058 DVDD.n5768 VSS 0.114418f
C23059 DVDD.n5769 VSS 0.033368f
C23060 DVDD.n5770 VSS 0.114418f
C23061 DVDD.n5771 VSS 0.114418f
C23062 DVDD.n5772 VSS 0.043862f
C23063 DVDD.n5773 VSS 0.058124f
C23064 DVDD.n5774 VSS 0.114418f
C23065 DVDD.n5775 VSS 0.114418f
C23066 DVDD.n5776 VSS 0.114418f
C23067 DVDD.n5777 VSS 0.114418f
C23068 DVDD.n5778 VSS 0.031484f
C23069 DVDD.n5779 VSS 0.030946f
C23070 DVDD.n5780 VSS 0.114418f
C23071 DVDD.n5781 VSS 0.033368f
C23072 DVDD.n5782 VSS 0.114418f
C23073 DVDD.n5783 VSS 0.033368f
C23074 DVDD.n5784 VSS 0.114418f
C23075 DVDD.n5785 VSS 0.033368f
C23076 DVDD.n5786 VSS 0.114418f
C23077 DVDD.n5787 VSS 0.033368f
C23078 DVDD.n5788 VSS 0.114418f
C23079 DVDD.n5789 VSS 0.033368f
C23080 DVDD.n5790 VSS 0.114418f
C23081 DVDD.n5791 VSS 0.033368f
C23082 DVDD.n5792 VSS 0.114418f
C23083 DVDD.n5793 VSS 0.114418f
C23084 DVDD.n5794 VSS 0.030408f
C23085 DVDD.n5795 VSS 0.032022f
C23086 DVDD.n5796 VSS 0.114418f
C23087 DVDD.n5797 VSS 0.033368f
C23088 DVDD.n5798 VSS 0.114418f
C23089 DVDD.n5799 VSS 0.033368f
C23090 DVDD.n5800 VSS 0.114418f
C23091 DVDD.n5801 VSS 0.033368f
C23092 DVDD.n5802 VSS 0.114418f
C23093 DVDD.n5803 VSS 0.033368f
C23094 DVDD.n5804 VSS 0.114418f
C23095 DVDD.n5805 VSS 0.033368f
C23096 DVDD.n5806 VSS 0.114418f
C23097 DVDD.n5807 VSS 0.033368f
C23098 DVDD.n5808 VSS 0.114418f
C23099 DVDD.n5809 VSS 0.114418f
C23100 DVDD.n5810 VSS 0.029331f
C23101 DVDD.n5811 VSS 0.033099f
C23102 DVDD.n5812 VSS 0.114418f
C23103 DVDD.n5813 VSS 0.033368f
C23104 DVDD.n5814 VSS 0.114418f
C23105 DVDD.n5815 VSS 0.033368f
C23106 DVDD.n5816 VSS 0.114418f
C23107 DVDD.n5817 VSS 0.033368f
C23108 DVDD.n5818 VSS 0.114418f
C23109 DVDD.n5819 VSS 0.033368f
C23110 DVDD.n5820 VSS 0.15585f
C23111 DVDD.t21 VSS 5.27557f
C23112 DVDD.n5822 VSS 0.15585f
C23113 DVDD.n5823 VSS 0.033368f
C23114 DVDD.n5824 VSS 0.029062f
C23115 DVDD.n5825 VSS 0.066735f
C23116 DVDD.n5826 VSS 0.066735f
C23117 DVDD.n5827 VSS 0.066735f
C23118 DVDD.n5828 VSS 0.033368f
C23119 DVDD.n5829 VSS 0.120351f
C23120 DVDD.n5830 VSS 0.058124f
C23121 DVDD.n5831 VSS 0.15585f
C23122 DVDD.n5832 VSS 0.114418f
C23123 DVDD.n5833 VSS 0.058124f
C23124 DVDD.n5834 VSS 0.114418f
C23125 DVDD.n5835 VSS 0.058124f
C23126 DVDD.n5836 VSS 0.114418f
C23127 DVDD.n5837 VSS 0.058124f
C23128 DVDD.n5838 VSS 0.114418f
C23129 DVDD.n5839 VSS 0.044401f
C23130 DVDD.t36 VSS 5.27557f
C23131 DVDD.n5841 VSS 0.033368f
C23132 DVDD.n5842 VSS 0.15585f
C23133 DVDD.n5843 VSS 0.033368f
C23134 DVDD.n5844 VSS 0.114418f
C23135 DVDD.n5845 VSS 0.033368f
C23136 DVDD.n5846 VSS 0.114418f
C23137 DVDD.n5847 VSS 0.033368f
C23138 DVDD.n5848 VSS 0.114418f
C23139 DVDD.n5849 VSS 0.033368f
C23140 DVDD.n5850 VSS 0.114418f
C23141 DVDD.n5851 VSS 0.114418f
C23142 DVDD.n5852 VSS 0.032561f
C23143 DVDD.n5853 VSS 0.029869f
C23144 DVDD.n5854 VSS 0.114418f
C23145 DVDD.n5855 VSS 0.033368f
C23146 DVDD.n5856 VSS 0.114418f
C23147 DVDD.n5857 VSS 0.033368f
C23148 DVDD.n5858 VSS 0.114418f
C23149 DVDD.n5859 VSS 0.033368f
C23150 DVDD.n5860 VSS 0.114418f
C23151 DVDD.n5861 VSS 0.114418f
C23152 DVDD.n5862 VSS 0.114418f
C23153 DVDD.n5863 VSS 0.058124f
C23154 DVDD.n5864 VSS 0.058124f
C23155 DVDD.n5865 VSS 0.058124f
C23156 DVDD.n5866 VSS 0.114418f
C23157 DVDD.n5867 VSS 0.114418f
C23158 DVDD.n5868 VSS 0.114418f
C23159 DVDD.n5869 VSS 0.058124f
C23160 DVDD.n5870 VSS 0.058124f
C23161 DVDD.n5871 VSS 0.058124f
C23162 DVDD.n5872 VSS 0.114418f
C23163 DVDD.n5873 VSS 0.114418f
C23164 DVDD.n5874 VSS 0.114418f
C23165 DVDD.n5875 VSS 0.058124f
C23166 DVDD.n5876 VSS 0.058124f
C23167 DVDD.n5877 VSS 0.058124f
C23168 DVDD.n5878 VSS 0.114418f
C23169 DVDD.n5879 VSS 0.114418f
C23170 DVDD.n5880 VSS 0.114418f
C23171 DVDD.n5881 VSS 0.058124f
C23172 DVDD.n5882 VSS 0.058124f
C23173 DVDD.n5883 VSS 0.058124f
C23174 DVDD.n5884 VSS 0.114418f
C23175 DVDD.n5885 VSS 0.114418f
C23176 DVDD.n5886 VSS 0.114418f
C23177 DVDD.n5887 VSS 0.045477f
C23178 DVDD.n5891 VSS 0.120351f
C23179 DVDD.n5892 VSS 0.105095f
C23180 DVDD.n5896 VSS 0.240702f
C23181 DVDD.n5897 VSS 0.240702f
C23182 DVDD.n5898 VSS 0.240702f
C23183 DVDD.n5899 VSS 0.105095f
C23184 DVDD.n5900 VSS 0.240702f
C23185 DVDD.n5901 VSS 0.240702f
C23186 DVDD.n5902 VSS 0.240702f
C23187 DVDD.n5903 VSS 0.240702f
C23188 DVDD.n5904 VSS 0.240702f
C23189 DVDD.n5905 VSS 0.222056f
C23190 DVDD.n5906 VSS 0.222056f
C23191 DVDD.n5907 VSS 0.271712f
C23192 DVDD.n5908 VSS 0.27258f
C23193 DVDD.n5909 VSS 0.240702f
C23194 DVDD.n5910 VSS 0.287049f
C23195 DVDD.n5911 VSS 0.240702f
C23196 DVDD.n5912 VSS 0.674186f
C23197 DVDD.n5913 VSS 0.240702f
C23198 DVDD.n5914 VSS 0.240702f
C23199 DVDD.n5915 VSS 0.240702f
C23200 DVDD.n5916 VSS 0.240702f
C23201 DVDD.n5917 VSS 0.120351f
C23202 DVDD.n5918 VSS 0.240702f
C23203 DVDD.n5919 VSS 0.240702f
C23204 DVDD.n5920 VSS 0.240702f
C23205 DVDD.n5921 VSS 0.105095f
C23206 DVDD.n5922 VSS 0.120351f
C23207 DVDD.n5923 VSS 0.029062f
C23208 DVDD.n5924 VSS 0.061085f
C23209 DVDD.n5928 VSS 0.105095f
C23210 DVDD.n5929 VSS 0.029062f
C23211 DVDD.n5930 VSS 0.029062f
C23212 DVDD.n5931 VSS 0.043862f
C23213 DVDD.n5932 VSS 0.066735f
C23214 DVDD.n5933 VSS 0.066735f
C23215 DVDD.n5934 VSS 0.114418f
C23216 DVDD.n5935 VSS 0.058124f
C23217 DVDD.n5936 VSS 0.114418f
C23218 DVDD.n5937 VSS 0.058124f
C23219 DVDD.n5938 VSS 0.114418f
C23220 DVDD.n5939 VSS 0.058124f
C23221 DVDD.n5940 VSS 0.114418f
C23222 DVDD.n5941 VSS 0.058124f
C23223 DVDD.t22 VSS 5.27557f
C23224 DVDD.n5943 VSS 0.033368f
C23225 DVDD.n5944 VSS 0.15585f
C23226 DVDD.n5945 VSS 0.033368f
C23227 DVDD.n5946 VSS 0.114418f
C23228 DVDD.n5947 VSS 0.033368f
C23229 DVDD.n5948 VSS 0.114418f
C23230 DVDD.n5949 VSS 0.033368f
C23231 DVDD.n5950 VSS 0.114418f
C23232 DVDD.n5951 VSS 0.033368f
C23233 DVDD.n5952 VSS 0.114418f
C23234 DVDD.n5953 VSS 0.114418f
C23235 DVDD.n5954 VSS 0.032561f
C23236 DVDD.n5955 VSS 0.029869f
C23237 DVDD.n5956 VSS 0.114418f
C23238 DVDD.n5957 VSS 0.033368f
C23239 DVDD.n5958 VSS 0.114418f
C23240 DVDD.n5959 VSS 0.033368f
C23241 DVDD.n5960 VSS 0.114418f
C23242 DVDD.n5961 VSS 0.033368f
C23243 DVDD.n5962 VSS 0.114418f
C23244 DVDD.n5963 VSS 0.114418f
C23245 DVDD.n5964 VSS 0.044401f
C23246 DVDD.n5965 VSS 0.058124f
C23247 DVDD.n5966 VSS 0.114418f
C23248 DVDD.n5967 VSS 0.114418f
C23249 DVDD.n5968 VSS 0.114418f
C23250 DVDD.n5969 VSS 0.058124f
C23251 DVDD.n5970 VSS 0.058124f
C23252 DVDD.n5971 VSS 0.058124f
C23253 DVDD.n5972 VSS 0.114418f
C23254 DVDD.n5973 VSS 0.114418f
C23255 DVDD.n5974 VSS 0.114418f
C23256 DVDD.n5975 VSS 0.058124f
C23257 DVDD.n5976 VSS 0.058124f
C23258 DVDD.n5977 VSS 0.058124f
C23259 DVDD.n5978 VSS 0.114418f
C23260 DVDD.n5979 VSS 0.114418f
C23261 DVDD.n5980 VSS 0.114418f
C23262 DVDD.n5981 VSS 0.058124f
C23263 DVDD.n5982 VSS 0.058124f
C23264 DVDD.n5983 VSS 0.058124f
C23265 DVDD.n5984 VSS 0.114418f
C23266 DVDD.n5985 VSS 0.114418f
C23267 DVDD.n5986 VSS 0.114418f
C23268 DVDD.n5987 VSS 0.058124f
C23269 DVDD.n5988 VSS 0.058124f
C23270 DVDD.n5989 VSS 0.045477f
C23271 DVDD.n5990 VSS 0.114418f
C23272 DVDD.n5991 VSS 0.15585f
C23273 DVDD.n5992 VSS 0.033368f
C23274 DVDD.n5993 VSS 0.054088f
C23275 DVDD.n5994 VSS 0.147472f
C23276 DVDD.n5995 VSS 0.117808f
C23277 DVDD.n5997 VSS 0.066735f
C23278 DVDD.n5999 VSS 0.066735f
C23279 DVDD.n6001 VSS 0.066735f
C23280 DVDD.n6002 VSS 0.120351f
C23281 DVDD.n6003 VSS 0.114418f
C23282 DVDD.n6004 VSS 0.114418f
C23283 DVDD.n6005 VSS 0.058124f
C23284 DVDD.n6006 VSS 0.051397f
C23285 DVDD.n6007 VSS 0.114418f
C23286 DVDD.n6008 VSS 0.033368f
C23287 DVDD.n6009 VSS 0.114418f
C23288 DVDD.n6010 VSS 0.114418f
C23289 DVDD.n6011 VSS 0.031484f
C23290 DVDD.n6012 VSS 0.030946f
C23291 DVDD.n6013 VSS 0.114418f
C23292 DVDD.n6014 VSS 0.033368f
C23293 DVDD.n6015 VSS 0.114418f
C23294 DVDD.n6016 VSS 0.033368f
C23295 DVDD.n6017 VSS 0.114418f
C23296 DVDD.n6018 VSS 0.033368f
C23297 DVDD.n6019 VSS 0.114418f
C23298 DVDD.n6020 VSS 0.033368f
C23299 DVDD.n6021 VSS 0.114418f
C23300 DVDD.n6022 VSS 0.033368f
C23301 DVDD.n6023 VSS 0.114418f
C23302 DVDD.n6024 VSS 0.033368f
C23303 DVDD.n6025 VSS 0.114418f
C23304 DVDD.n6026 VSS 0.114418f
C23305 DVDD.n6027 VSS 0.030408f
C23306 DVDD.n6028 VSS 0.032022f
C23307 DVDD.n6029 VSS 0.114418f
C23308 DVDD.n6030 VSS 0.033368f
C23309 DVDD.n6031 VSS 0.114418f
C23310 DVDD.n6032 VSS 0.033368f
C23311 DVDD.n6033 VSS 0.114418f
C23312 DVDD.n6034 VSS 0.033368f
C23313 DVDD.n6035 VSS 0.114418f
C23314 DVDD.n6036 VSS 0.033368f
C23315 DVDD.n6037 VSS 0.114418f
C23316 DVDD.n6038 VSS 0.033368f
C23317 DVDD.n6039 VSS 0.114418f
C23318 DVDD.n6040 VSS 0.033368f
C23319 DVDD.n6041 VSS 0.114418f
C23320 DVDD.n6042 VSS 0.114418f
C23321 DVDD.n6043 VSS 0.029331f
C23322 DVDD.n6044 VSS 0.033099f
C23323 DVDD.n6045 VSS 0.114418f
C23324 DVDD.n6046 VSS 0.033368f
C23325 DVDD.n6047 VSS 0.114418f
C23326 DVDD.n6048 VSS 0.033368f
C23327 DVDD.n6049 VSS 0.114418f
C23328 DVDD.n6050 VSS 0.033368f
C23329 DVDD.n6051 VSS 0.114418f
C23330 DVDD.n6052 VSS 0.033368f
C23331 DVDD.n6053 VSS 0.15585f
C23332 DVDD.t3 VSS 5.27557f
C23333 DVDD.n6055 VSS 0.033368f
C23334 DVDD.n6056 VSS 0.15585f
C23335 DVDD.n6057 VSS 0.033368f
C23336 DVDD.n6058 VSS 0.114418f
C23337 DVDD.n6059 VSS 0.114418f
C23338 DVDD.n6060 VSS 0.033368f
C23339 DVDD.n6061 VSS 0.029062f
C23340 DVDD.n6062 VSS 0.120351f
C23341 DVDD.n6063 VSS 0.105095f
C23342 DVDD.n6064 VSS 0.240702f
C23343 DVDD.n6065 VSS 0.240702f
C23344 DVDD.n6066 VSS 0.240702f
C23345 DVDD.n6067 VSS 0.240702f
C23346 DVDD.n6068 VSS 0.240702f
C23347 DVDD.n6069 VSS 0.195782f
C23348 DVDD.n6070 VSS 0.240702f
C23349 DVDD.n6071 VSS 0.240702f
C23350 DVDD.n6072 VSS 0.240702f
C23351 DVDD.n6073 VSS 0.240702f
C23352 DVDD.n6074 VSS 0.240702f
C23353 DVDD.n6075 VSS 0.240702f
C23354 DVDD.n6076 VSS 0.240702f
C23355 DVDD.n6077 VSS 0.240702f
C23356 DVDD.n6078 VSS 0.240702f
C23357 DVDD.n6079 VSS 0.161033f
C23358 DVDD.n6080 VSS 0.161033f
C23359 DVDD.n6081 VSS 0.161033f
C23360 DVDD.n6082 VSS 0.701473f
C23361 DVDD.n6083 VSS 0.222056f
C23362 DVDD.n6084 VSS 0.240702f
C23363 DVDD.n6085 VSS 0.240702f
C23364 DVDD.n6086 VSS 0.240702f
C23365 DVDD.n6087 VSS 0.240702f
C23366 DVDD.n6088 VSS 0.240702f
C23367 DVDD.n6089 VSS 0.240702f
C23368 DVDD.n6090 VSS 0.240702f
C23369 DVDD.n6091 VSS 0.240702f
C23370 DVDD.n6092 VSS 0.240702f
C23371 DVDD.n6093 VSS 0.240702f
C23372 DVDD.n6094 VSS 0.192392f
C23373 DVDD.n6095 VSS 0.120351f
C23374 DVDD.n6096 VSS 0.029062f
C23375 DVDD.n6097 VSS 0.120351f
C23376 DVDD.n6098 VSS 0.180526f
C23377 DVDD.n6099 VSS 0.2068f
C23378 DVDD.n6100 VSS 0.2068f
C23379 DVDD.n6101 VSS 0.346009f
C23380 DVDD.n6102 VSS 0.387751f
C23381 DVDD.n6103 VSS 0.451316f
C23382 DVDD.n6104 VSS 0.451316f
C23383 DVDD.n6105 VSS 0.197054f
C23384 DVDD.n6106 VSS 0.197054f
C23385 DVDD.n6107 VSS 0.066735f
C23386 DVDD.n6109 VSS 0.066735f
C23387 DVDD.n6111 VSS 0.225658f
C23388 DVDD.n6112 VSS 0.029062f
C23389 DVDD.n6113 VSS 0.225658f
C23390 DVDD.n6114 VSS 0.197054f
C23391 DVDD.n6115 VSS 0.451316f
C23392 DVDD.n6116 VSS 0.451316f
C23393 DVDD.n6117 VSS 0.451316f
C23394 DVDD.n6118 VSS 0.451316f
C23395 DVDD.n6119 VSS 0.451316f
C23396 DVDD.n6120 VSS 0.451316f
C23397 DVDD.n6121 VSS 0.451316f
C23398 DVDD.n6122 VSS 0.451316f
C23399 DVDD.n6123 VSS 0.451316f
C23400 DVDD.n6124 VSS 0.451316f
C23401 DVDD.n6125 VSS 0.451316f
C23402 DVDD.n6126 VSS 0.451316f
C23403 DVDD.n6127 VSS 0.451316f
C23404 DVDD.n6128 VSS 0.451316f
C23405 DVDD.n6129 VSS 0.451316f
C23406 DVDD.n6130 VSS 0.451316f
C23407 DVDD.n6131 VSS 0.451316f
C23408 DVDD.n6132 VSS 0.451316f
C23409 DVDD.n6133 VSS 0.451316f
C23410 DVDD.n6134 VSS 0.451316f
C23411 DVDD.n6135 VSS 0.451316f
C23412 DVDD.n6136 VSS 0.451316f
C23413 DVDD.n6137 VSS 0.451316f
C23414 DVDD.n6138 VSS 0.451316f
C23415 DVDD.n6139 VSS 0.451316f
C23416 DVDD.n6140 VSS 0.451316f
C23417 DVDD.n6141 VSS 0.451316f
C23418 DVDD.n6142 VSS 0.451316f
C23419 DVDD.n6143 VSS 0.451316f
C23420 DVDD.n6144 VSS 0.451316f
C23421 DVDD.n6145 VSS 0.451316f
C23422 DVDD.n6146 VSS 0.367092f
C23423 DVDD.n6147 VSS 0.451316f
C23424 DVDD.n6148 VSS 0.451316f
C23425 DVDD.n6149 VSS 0.451316f
C23426 DVDD.n6150 VSS 0.451316f
C23427 DVDD.n6151 VSS 0.451316f
C23428 DVDD.n6152 VSS 0.197054f
C23429 DVDD.n6153 VSS 0.225658f
C23430 DVDD.n6154 VSS 0.16065f
C23431 DVDD.n6155 VSS 0.225658f
C23432 DVDD.n6156 VSS 0.220891f
C23433 DVDD.n6157 VSS 0.276511f
C23434 DVDD.n6158 VSS 0.276511f
C23435 DVDD.n6159 VSS 0.346009f
C23436 DVDD.n6160 VSS 0.400464f
C23437 DVDD.n6161 VSS 0.400464f
C23438 DVDD.n6162 VSS 0.400464f
C23439 DVDD.n6163 VSS 0.451316f
C23440 DVDD.n6164 VSS 0.451316f
C23441 DVDD.n6165 VSS 0.451316f
C23442 DVDD.n6166 VSS 0.451316f
C23443 DVDD.n6167 VSS 0.451316f
C23444 DVDD.n6168 VSS 0.451316f
C23445 DVDD.n6169 VSS 0.451316f
C23446 DVDD.n6170 VSS 0.451316f
C23447 DVDD.n6171 VSS 0.451316f
C23448 DVDD.n6172 VSS 0.451316f
C23449 DVDD.n6173 VSS 0.451316f
C23450 DVDD.n6174 VSS 0.451316f
C23451 DVDD.n6175 VSS 0.451316f
C23452 DVDD.n6176 VSS 0.451316f
C23453 DVDD.n6177 VSS 0.451316f
C23454 DVDD.n6178 VSS 0.451316f
C23455 DVDD.n6179 VSS 0.451316f
C23456 DVDD.n6180 VSS 0.367092f
C23457 DVDD.n6181 VSS 0.451316f
C23458 DVDD.n6182 VSS 0.451316f
C23459 DVDD.n6183 VSS 0.451316f
C23460 DVDD.n6184 VSS 0.451316f
C23461 DVDD.n6185 VSS 0.451316f
C23462 DVDD.n6186 VSS 0.197054f
C23463 DVDD.n6187 VSS 0.451316f
C23464 DVDD.n6188 VSS 0.197054f
C23465 DVDD.n6189 VSS 0.451316f
C23466 DVDD.n6190 VSS 0.451316f
C23467 DVDD.n6191 VSS 0.451316f
C23468 DVDD.n6192 VSS 0.451316f
C23469 DVDD.n6193 VSS 0.451316f
C23470 DVDD.n6194 VSS 0.451316f
C23471 DVDD.n6195 VSS 0.451316f
C23472 DVDD.n6196 VSS 0.451316f
C23473 DVDD.n6197 VSS 0.451316f
C23474 DVDD.n6198 VSS 0.451316f
C23475 DVDD.n6199 VSS 0.451316f
C23476 DVDD.n6200 VSS 0.451316f
C23477 DVDD.n6201 VSS 0.451316f
C23478 DVDD.n6202 VSS 0.451316f
C23479 DVDD.n6203 VSS 0.451316f
C23480 DVDD.n6204 VSS 0.451316f
C23481 DVDD.n6205 VSS 0.263798f
C23482 DVDD.n6206 VSS 0.451316f
C23483 DVDD.n6207 VSS 0.451316f
C23484 DVDD.n6208 VSS 0.451316f
C23485 DVDD.n6209 VSS 0.263798f
C23486 DVDD.n6210 VSS 0.346009f
C23487 DVDD.n6211 VSS 0.140692f
C23488 DVDD.n6212 VSS 0.240702f
C23489 DVDD.n6213 VSS 0.240702f
C23490 DVDD.n6214 VSS 0.140692f
C23491 DVDD.n6215 VSS 0.240702f
C23492 DVDD.n6216 VSS 0.240702f
C23493 DVDD.n6217 VSS 0.240702f
C23494 DVDD.n6218 VSS 0.240702f
C23495 DVDD.n6219 VSS 0.240702f
C23496 DVDD.n6220 VSS 0.240702f
C23497 DVDD.n6221 VSS 0.240702f
C23498 DVDD.n6222 VSS 0.240702f
C23499 DVDD.n6223 VSS 0.240702f
C23500 DVDD.n6224 VSS 0.240702f
C23501 DVDD.n6225 VSS 0.240702f
C23502 DVDD.n6226 VSS 0.240702f
C23503 DVDD.n6227 VSS 0.240702f
C23504 DVDD.n6228 VSS 0.240702f
C23505 DVDD.n6229 VSS 0.240702f
C23506 DVDD.n6230 VSS 0.105095f
C23507 DVDD.n6231 VSS 0.240702f
C23508 DVDD.n6232 VSS 0.167813f
C23509 DVDD.n6233 VSS 0.167813f
C23510 DVDD.n6234 VSS 0.172475f
C23511 DVDD.n6235 VSS 0.045979f
C23512 DVDD.n6236 VSS 0.060175f
C23513 DVDD.n6237 VSS 0.170687f
C23514 DVDD.n6238 VSS 0.060175f
C23515 DVDD.n6239 VSS 0.027333f
C23516 DVDD.n6240 VSS 0.066735f
C23517 DVDD.n6242 VSS 0.026274f
C23518 DVDD.n6243 VSS 0.057655f
C23519 DVDD.n6244 VSS 0.059611f
C23520 DVDD.n6245 VSS 0.058124f
C23521 DVDD.n6246 VSS 0.114418f
C23522 DVDD.n6247 VSS 0.058124f
C23523 DVDD.n6248 VSS 0.114418f
C23524 DVDD.n6249 VSS 0.058124f
C23525 DVDD.n6250 VSS 0.114418f
C23526 DVDD.n6251 VSS 0.058124f
C23527 DVDD.n6252 VSS 0.114418f
C23528 DVDD.n6253 VSS 0.044401f
C23529 DVDD.n6254 VSS 0.033368f
C23530 DVDD.n6255 VSS 0.114418f
C23531 DVDD.n6256 VSS 0.033368f
C23532 DVDD.n6257 VSS 0.114418f
C23533 DVDD.n6258 VSS 0.033368f
C23534 DVDD.n6259 VSS 0.114418f
C23535 DVDD.n6260 VSS 0.033368f
C23536 DVDD.n6261 VSS 0.114418f
C23537 DVDD.n6262 VSS 0.114418f
C23538 DVDD.n6263 VSS 0.032561f
C23539 DVDD.n6264 VSS 0.029869f
C23540 DVDD.n6265 VSS 0.114418f
C23541 DVDD.n6266 VSS 0.033368f
C23542 DVDD.n6267 VSS 0.114418f
C23543 DVDD.n6268 VSS 0.033368f
C23544 DVDD.n6269 VSS 0.114418f
C23545 DVDD.n6270 VSS 0.033368f
C23546 DVDD.n6271 VSS 0.114418f
C23547 DVDD.n6272 VSS 0.114418f
C23548 DVDD.n6273 VSS 0.114418f
C23549 DVDD.n6274 VSS 0.058124f
C23550 DVDD.n6275 VSS 0.058124f
C23551 DVDD.n6276 VSS 0.058124f
C23552 DVDD.n6277 VSS 0.114418f
C23553 DVDD.n6278 VSS 0.114418f
C23554 DVDD.n6279 VSS 0.114418f
C23555 DVDD.n6280 VSS 0.058124f
C23556 DVDD.n6281 VSS 0.058124f
C23557 DVDD.n6282 VSS 0.058124f
C23558 DVDD.n6283 VSS 0.114418f
C23559 DVDD.n6284 VSS 0.114418f
C23560 DVDD.n6285 VSS 0.114418f
C23561 DVDD.n6286 VSS 0.058124f
C23562 DVDD.n6287 VSS 0.058124f
C23563 DVDD.n6288 VSS 0.058124f
C23564 DVDD.n6289 VSS 0.114418f
C23565 DVDD.n6290 VSS 0.114418f
C23566 DVDD.n6291 VSS 0.114418f
C23567 DVDD.n6292 VSS 0.058124f
C23568 DVDD.n6293 VSS 0.058124f
C23569 DVDD.n6294 VSS 0.058124f
C23570 DVDD.n6295 VSS 0.114418f
C23571 DVDD.n6296 VSS 0.114418f
C23572 DVDD.n6297 VSS 0.114418f
C23573 DVDD.n6298 VSS 0.045477f
C23574 DVDD.n6299 VSS 0.029062f
C23575 DVDD.n6300 VSS 0.033368f
C23576 DVDD.n6301 VSS 0.054088f
C23577 DVDD.n6303 VSS 0.066735f
C23578 DVDD.n6304 VSS 0.029028f
C23579 DVDD.n6305 VSS 0.026274f
C23580 DVDD.n6306 VSS 0.060175f
C23581 DVDD.n6307 VSS 0.060175f
C23582 DVDD.n6308 VSS 0.026274f
C23583 DVDD.n6309 VSS 0.030088f
C23584 DVDD.n6310 VSS 0.066735f
C23585 DVDD.n6312 VSS 0.066735f
C23586 DVDD.n6314 VSS 0.066735f
C23587 DVDD.n6315 VSS 0.030088f
C23588 DVDD.n6316 VSS 0.026274f
C23589 DVDD.n6317 VSS 0.060175f
C23590 DVDD.n6318 VSS 0.060175f
C23591 DVDD.n6319 VSS 0.026274f
C23592 DVDD.n6320 VSS 0.030088f
C23593 DVDD.n6321 VSS 0.029062f
C23594 DVDD.n6322 VSS 0.114418f
C23595 DVDD.n6323 VSS 0.033368f
C23596 DVDD.n6324 VSS 0.029062f
C23597 DVDD.n6325 VSS 0.02691f
C23598 DVDD.n6326 VSS 0.060739f
C23599 DVDD.n6327 VSS 0.029062f
C23600 DVDD.n6328 VSS 0.043862f
C23601 DVDD.n6329 VSS 0.114418f
C23602 DVDD.n6330 VSS 0.114418f
C23603 DVDD.n6331 VSS 0.114418f
C23604 DVDD.n6332 VSS 0.051397f
C23605 DVDD.n6333 VSS 0.029062f
C23606 DVDD.n6334 VSS 0.225658f
C23607 DVDD.n6335 VSS 0.029062f
C23608 DVDD.n6336 VSS 0.033368f
C23609 DVDD.n6337 VSS 0.15585f
C23610 DVDD.n6338 VSS 0.031397f
C23611 DVDD.n6339 VSS 0.131369f
C23612 DVDD.n6340 VSS 0.031397f
C23613 DVDD.n6341 VSS 0.131369f
C23614 DVDD.n6342 VSS 0.031397f
C23615 DVDD.n6343 VSS 0.131369f
C23616 DVDD.n6344 VSS 0.031397f
C23617 DVDD.n6345 VSS 0.131369f
C23618 DVDD.n6346 VSS 0.031397f
C23619 DVDD.n6347 VSS 0.131369f
C23620 DVDD.n6348 VSS 0.031397f
C23621 DVDD.n6349 VSS 0.131369f
C23622 DVDD.n6350 VSS 0.031397f
C23623 DVDD.n6351 VSS 0.131369f
C23624 DVDD.n6352 VSS 0.031397f
C23625 DVDD.n6353 VSS 0.131369f
C23626 DVDD.n6354 VSS 0.031397f
C23627 DVDD.n6355 VSS 0.131369f
C23628 DVDD.n6356 VSS 0.031397f
C23629 DVDD.n6357 VSS 0.131369f
C23630 DVDD.n6358 VSS 0.031397f
C23631 DVDD.n6359 VSS 0.131369f
C23632 DVDD.n6360 VSS 0.031397f
C23633 DVDD.n6361 VSS 0.131369f
C23634 DVDD.n6362 VSS 0.031397f
C23635 DVDD.n6363 VSS 0.131369f
C23636 DVDD.n6364 VSS 0.031397f
C23637 DVDD.n6365 VSS 0.131369f
C23638 DVDD.n6366 VSS 0.031397f
C23639 DVDD.n6367 VSS 0.131369f
C23640 DVDD.n6368 VSS 0.031397f
C23641 DVDD.n6369 VSS 0.131369f
C23642 DVDD.n6370 VSS 0.031397f
C23643 DVDD.n6371 VSS 0.131369f
C23644 DVDD.n6372 VSS 0.031397f
C23645 DVDD.n6373 VSS 0.131369f
C23646 DVDD.n6374 VSS 0.031397f
C23647 DVDD.n6375 VSS 0.124509f
C23648 DVDD.t20 VSS 5.27557f
C23649 DVDD.n6376 VSS 0.031397f
C23650 DVDD.n6377 VSS 0.124509f
C23651 DVDD.n6378 VSS 0.031397f
C23652 DVDD.n6379 VSS 0.131369f
C23653 DVDD.n6380 VSS 0.031397f
C23654 DVDD.n6381 VSS 0.131369f
C23655 DVDD.n6382 VSS 0.037371f
C23656 DVDD.n6383 VSS 0.131369f
C23657 DVDD.n6384 VSS 0.131369f
C23658 DVDD.n6385 VSS 0.131369f
C23659 DVDD.n6386 VSS 0.034156f
C23660 DVDD.n6387 VSS 0.197054f
C23661 DVDD.n6388 VSS 0.451316f
C23662 DVDD.n6389 VSS 0.451316f
C23663 DVDD.n6390 VSS 0.451316f
C23664 DVDD.n6391 VSS 0.40682f
C23665 DVDD.n6392 VSS 0.050852f
C23666 DVDD.n6393 VSS 2.07943f
C23667 DVDD.n6394 VSS 0.6412f
C23668 DVDD.n6395 VSS 0.40682f
C23669 DVDD.n6396 VSS 0.197054f
C23670 DVDD.n6397 VSS 0.225658f
C23671 DVDD.n6398 VSS 0.031583f
C23672 DVDD.n6399 VSS 0.225658f
C23673 DVDD.n6400 VSS 0.367092f
C23674 DVDD.n6401 VSS 0.451316f
C23675 DVDD.n6402 VSS 0.451316f
C23676 DVDD.n6403 VSS 0.451316f
C23677 DVDD.n6404 VSS 0.451316f
C23678 DVDD.n6405 VSS 0.451316f
C23679 DVDD.n6406 VSS 0.395696f
C23680 DVDD.n6407 VSS 0.451316f
C23681 DVDD.n6408 VSS 0.197054f
C23682 DVDD.n6409 VSS 0.451316f
C23683 DVDD.n6420 VSS 0.225658f
C23684 DVDD.n6421 VSS 0.197054f
C23685 DVDD.n6422 VSS 0.451316f
C23686 DVDD.n6423 VSS 0.413177f
C23687 DVDD.n6424 VSS 0.346009f
C23688 DVDD.n6425 VSS 0.220361f
C23689 DVDD.n6426 VSS 0.105095f
C23690 DVDD.n6427 VSS 0.240702f
C23691 DVDD.n6428 VSS 0.240702f
C23692 DVDD.n6429 VSS 0.240702f
C23693 DVDD.n6430 VSS 0.240702f
C23694 DVDD.n6431 VSS 0.240702f
C23695 DVDD.n6432 VSS 0.211038f
C23696 DVDD.n6433 VSS 0.240702f
C23697 DVDD.n6434 VSS 0.240702f
C23698 DVDD.n6435 VSS 0.240702f
C23699 DVDD.n6436 VSS 0.240702f
C23700 DVDD.n6437 VSS 0.240702f
C23701 DVDD.n6438 VSS 0.240702f
C23702 DVDD.n6439 VSS 0.240702f
C23703 DVDD.n6440 VSS 0.240702f
C23704 DVDD.n6441 VSS 0.240702f
C23705 DVDD.n6442 VSS 0.105095f
C23706 DVDD.n6443 VSS 0.208495f
C23707 DVDD.n6444 VSS 0.208495f
C23708 DVDD.n6445 VSS 0.127355f
C23709 DVDD.n6446 VSS 0.103735f
C23710 DVDD.n6447 VSS 0.103735f
C23711 DVDD.n6448 VSS 0.061545f
C23712 DVDD.n6449 VSS 0.082435f
C23713 DVDD.n6450 VSS 0.055589f
C23714 DVDD.n6451 VSS 0.070479f
C23715 DVDD.n6452 VSS 0.070479f
C23716 DVDD.n6453 VSS 0.061545f
C23717 DVDD.n6454 VSS 0.140961f
C23718 DVDD.n6455 VSS 0.140961f
C23719 DVDD.n6456 VSS 0.401144f
C23720 DVDD.n6457 VSS 0.133867f
C23721 DVDD.n6458 VSS 0.140961f
C23722 DVDD.n6459 VSS 0.061545f
C23723 DVDD.n6460 VSS 0.064028f
C23724 DVDD.n6461 VSS 0.067998f
C23725 DVDD.n6463 VSS 0.062794f
C23726 DVDD.n6464 VSS 0.120351f
C23727 DVDD.n6465 VSS 0.031467f
C23728 DVDD.n6466 VSS 0.031397f
C23729 DVDD.n6467 VSS 0.124509f
C23730 DVDD.t35 VSS 5.27557f
C23731 DVDD.n6468 VSS 0.124509f
C23732 DVDD.n6469 VSS 0.031397f
C23733 DVDD.n6470 VSS 0.045323f
C23734 DVDD.n6471 VSS 0.062794f
C23735 DVDD.n6472 VSS 0.062794f
C23736 DVDD.n6473 VSS 0.043804f
C23737 DVDD.n6474 VSS 0.031397f
C23738 DVDD.n6475 VSS 0.031397f
C23739 DVDD.n6476 VSS 0.031397f
C23740 DVDD.n6477 VSS 0.031397f
C23741 DVDD.n6481 VSS 0.225658f
C23742 DVDD.n6485 VSS 0.181162f
C23743 DVDD.n6486 VSS 0.048607f
C23744 DVDD.n6487 VSS 0.131369f
C23745 DVDD.n6488 VSS 0.033368f
C23746 DVDD.n6489 VSS 0.15585f
C23747 DVDD.n6490 VSS 0.033368f
C23748 DVDD.n6491 VSS 0.114418f
C23749 DVDD.n6492 VSS 0.033368f
C23750 DVDD.n6493 VSS 0.114418f
C23751 DVDD.n6494 VSS 0.033368f
C23752 DVDD.n6495 VSS 0.114418f
C23753 DVDD.n6496 VSS 0.033368f
C23754 DVDD.n6497 VSS 0.114418f
C23755 DVDD.n6498 VSS 0.114418f
C23756 DVDD.n6499 VSS 0.031484f
C23757 DVDD.n6500 VSS 0.030946f
C23758 DVDD.n6501 VSS 0.114418f
C23759 DVDD.n6502 VSS 0.033368f
C23760 DVDD.n6503 VSS 0.114418f
C23761 DVDD.n6504 VSS 0.033368f
C23762 DVDD.n6505 VSS 0.114418f
C23763 DVDD.n6506 VSS 0.033368f
C23764 DVDD.n6507 VSS 0.114418f
C23765 DVDD.n6508 VSS 0.033368f
C23766 DVDD.n6509 VSS 0.114418f
C23767 DVDD.n6510 VSS 0.033368f
C23768 DVDD.n6511 VSS 0.114418f
C23769 DVDD.n6512 VSS 0.033368f
C23770 DVDD.n6513 VSS 0.114418f
C23771 DVDD.n6514 VSS 0.114418f
C23772 DVDD.n6515 VSS 0.030408f
C23773 DVDD.n6516 VSS 0.032022f
C23774 DVDD.n6517 VSS 0.114418f
C23775 DVDD.n6518 VSS 0.033368f
C23776 DVDD.n6519 VSS 0.114418f
C23777 DVDD.n6520 VSS 0.033368f
C23778 DVDD.n6521 VSS 0.114418f
C23779 DVDD.n6522 VSS 0.114418f
C23780 DVDD.n6523 VSS 0.046553f
C23781 DVDD.n6524 VSS 0.058124f
C23782 DVDD.n6525 VSS 0.114418f
C23783 DVDD.n6526 VSS 0.114418f
C23784 DVDD.n6527 VSS 0.114418f
C23785 DVDD.n6528 VSS 0.033368f
C23786 DVDD.n6529 VSS 0.114418f
C23787 DVDD.n6530 VSS 0.114418f
C23788 DVDD.n6531 VSS 0.031484f
C23789 DVDD.n6532 VSS 0.030946f
C23790 DVDD.n6533 VSS 0.114418f
C23791 DVDD.n6534 VSS 0.033368f
C23792 DVDD.n6535 VSS 0.114418f
C23793 DVDD.n6536 VSS 0.033368f
C23794 DVDD.n6537 VSS 0.114418f
C23795 DVDD.n6538 VSS 0.033368f
C23796 DVDD.n6539 VSS 0.114418f
C23797 DVDD.n6540 VSS 0.033368f
C23798 DVDD.n6541 VSS 0.114418f
C23799 DVDD.n6542 VSS 0.033368f
C23800 DVDD.n6543 VSS 0.15585f
C23801 DVDD.n6544 VSS 0.031397f
C23802 DVDD.n6545 VSS 0.131369f
C23803 DVDD.n6546 VSS 0.031397f
C23804 DVDD.n6547 VSS 0.131369f
C23805 DVDD.n6548 VSS 0.031397f
C23806 DVDD.n6549 VSS 0.131369f
C23807 DVDD.n6550 VSS 0.031397f
C23808 DVDD.n6551 VSS 0.131369f
C23809 DVDD.n6552 VSS 0.031397f
C23810 DVDD.n6553 VSS 0.131369f
C23811 DVDD.n6554 VSS 0.031397f
C23812 DVDD.n6555 VSS 0.131369f
C23813 DVDD.n6556 VSS 0.031397f
C23814 DVDD.n6557 VSS 0.124509f
C23815 DVDD.t16 VSS 5.27557f
C23816 DVDD.n6558 VSS 0.031397f
C23817 DVDD.n6559 VSS 0.124509f
C23818 DVDD.n6560 VSS 0.031397f
C23819 DVDD.n6561 VSS 0.131369f
C23820 DVDD.n6562 VSS 0.031397f
C23821 DVDD.n6563 VSS 0.131369f
C23822 DVDD.n6564 VSS 0.031397f
C23823 DVDD.n6565 VSS 0.131369f
C23824 DVDD.n6566 VSS 0.031397f
C23825 DVDD.n6567 VSS 0.131369f
C23826 DVDD.n6568 VSS 0.031397f
C23827 DVDD.n6569 VSS 0.131369f
C23828 DVDD.n6570 VSS 0.031397f
C23829 DVDD.n6571 VSS 0.131369f
C23830 DVDD.n6572 VSS 0.031397f
C23831 DVDD.n6573 VSS 0.131369f
C23832 DVDD.n6574 VSS 0.031397f
C23833 DVDD.n6575 VSS 0.131369f
C23834 DVDD.n6576 VSS 0.031397f
C23835 DVDD.n6577 VSS 0.131369f
C23836 DVDD.n6578 VSS 0.031397f
C23837 DVDD.n6579 VSS 0.131369f
C23838 DVDD.n6580 VSS 0.031397f
C23839 DVDD.n6581 VSS 0.131369f
C23840 DVDD.n6582 VSS 0.031397f
C23841 DVDD.n6583 VSS 0.131369f
C23842 DVDD.n6584 VSS 0.031397f
C23843 DVDD.n6585 VSS 0.131369f
C23844 DVDD.n6586 VSS 0.031397f
C23845 DVDD.n6587 VSS 0.131369f
C23846 DVDD.n6588 VSS 0.035291f
C23847 DVDD.n6589 VSS 0.131369f
C23848 DVDD.n6590 VSS 0.131369f
C23849 DVDD.n6591 VSS 0.131369f
C23850 DVDD.n6592 VSS 0.035031f
C23851 DVDD.n6593 VSS 0.197054f
C23852 DVDD.n6594 VSS 0.451316f
C23853 DVDD.n6595 VSS 0.451316f
C23854 DVDD.n6596 VSS 0.451316f
C23855 DVDD.n6597 VSS 0.40682f
C23856 DVDD.n6598 VSS 0.050852f
C23857 DVDD.n6599 VSS 2.07943f
C23858 DVDD.n6600 VSS 0.6412f
C23859 DVDD.n6601 VSS 0.40682f
C23860 DVDD.n6602 VSS 0.197054f
C23861 DVDD.n6603 VSS 0.225658f
C23862 DVDD.n6604 VSS 0.031818f
C23863 DVDD.n6605 VSS 0.225658f
C23864 DVDD.n6606 VSS 0.367092f
C23865 DVDD.n6607 VSS 0.451316f
C23866 DVDD.n6608 VSS 0.451316f
C23867 DVDD.n6609 VSS 0.451316f
C23868 DVDD.n6610 VSS 0.451316f
C23869 DVDD.n6611 VSS 0.451316f
C23870 DVDD.n6612 VSS 0.395696f
C23871 DVDD.n6613 VSS 0.451316f
C23872 DVDD.n6614 VSS 0.197054f
C23873 DVDD.n6615 VSS 0.451316f
C23874 DVDD.n6626 VSS 0.225658f
C23875 DVDD.n6627 VSS 0.197054f
C23876 DVDD.n6628 VSS 0.451316f
C23877 DVDD.n6629 VSS 0.413177f
C23878 DVDD.n6630 VSS 0.543486f
C23879 DVDD.n6631 VSS 0.263798f
C23880 DVDD.n6632 VSS 0.263798f
C23881 DVDD.n6633 VSS 0.451316f
C23882 DVDD.n6634 VSS 0.451316f
C23883 DVDD.n6635 VSS 0.451316f
C23884 DVDD.n6636 VSS 0.451316f
C23885 DVDD.n6637 VSS 0.451316f
C23886 DVDD.n6638 VSS 0.451316f
C23887 DVDD.n6639 VSS 0.451316f
C23888 DVDD.n6640 VSS 0.451316f
C23889 DVDD.n6641 VSS 0.451316f
C23890 DVDD.n6642 VSS 0.451316f
C23891 DVDD.n6643 VSS 0.451316f
C23892 DVDD.n6644 VSS 0.395696f
C23893 DVDD.n6648 VSS 0.225658f
C23894 DVDD.n6649 VSS 0.029062f
C23895 DVDD.n6650 VSS 0.225658f
C23896 DVDD.n6651 VSS 0.367092f
C23897 DVDD.n6652 VSS 0.451316f
C23898 DVDD.n6653 VSS 0.451316f
C23899 DVDD.n6654 VSS 0.451316f
C23900 DVDD.n6655 VSS 0.451316f
C23901 DVDD.n6656 VSS 0.451316f
C23902 DVDD.n6657 VSS 0.451316f
C23903 DVDD.n6658 VSS 0.451316f
C23904 DVDD.n6659 VSS 0.451316f
C23905 DVDD.n6660 VSS 0.451316f
C23906 DVDD.n6661 VSS 0.451316f
C23907 DVDD.n6662 VSS 0.451316f
C23908 DVDD.n6663 VSS 0.451316f
C23909 DVDD.n6664 VSS 0.451316f
C23910 DVDD.n6665 VSS 0.451316f
C23911 DVDD.n6666 VSS 0.451316f
C23912 DVDD.n6667 VSS 0.400464f
C23913 DVDD.n6668 VSS 0.400464f
C23914 DVDD.n6669 VSS 0.543486f
C23915 DVDD.n6670 VSS 0.220891f
C23916 DVDD.n6671 VSS 0.276511f
C23917 DVDD.n6672 VSS 0.451316f
C23918 DVDD.n6673 VSS 0.197054f
C23919 DVDD.n6674 VSS 0.225658f
C23920 DVDD.n6675 VSS 0.029062f
C23921 DVDD.n6676 VSS 0.225658f
C23922 DVDD.n6677 VSS 0.367092f
C23923 DVDD.n6678 VSS 0.451316f
C23924 DVDD.n6679 VSS 0.451316f
C23925 DVDD.n6680 VSS 0.451316f
C23926 DVDD.n6681 VSS 0.451316f
C23927 DVDD.n6682 VSS 0.451316f
C23928 DVDD.n6683 VSS 0.451316f
C23929 DVDD.n6684 VSS 0.451316f
C23930 DVDD.n6685 VSS 0.451316f
C23931 DVDD.n6686 VSS 0.451316f
C23932 DVDD.n6687 VSS 0.451316f
C23933 DVDD.n6688 VSS 0.451316f
C23934 DVDD.n6689 VSS 0.451316f
C23935 DVDD.n6690 VSS 0.451316f
C23936 DVDD.n6691 VSS 0.451316f
C23937 DVDD.n6692 VSS 0.451316f
C23938 DVDD.n6693 VSS 0.451316f
C23939 DVDD.n6694 VSS 0.451316f
C23940 DVDD.n6695 VSS 0.451316f
C23941 DVDD.n6696 VSS 0.451316f
C23942 DVDD.n6697 VSS 0.451316f
C23943 DVDD.n6698 VSS 0.451316f
C23944 DVDD.n6699 VSS 0.451316f
C23945 DVDD.n6700 VSS 0.360735f
C23946 DVDD.n6704 VSS 0.225658f
C23947 DVDD.n6705 VSS 0.029062f
C23948 DVDD.n6706 VSS 0.225658f
C23949 DVDD.n6707 VSS 0.338487f
C23950 DVDD.n6708 VSS 0.387751f
C23951 DVDD.n6709 VSS 0.543486f
C23952 DVDD.n6710 VSS 0.289224f
C23953 DVDD.n6711 VSS 0.289224f
C23954 DVDD.n6712 VSS 0.451316f
C23955 DVDD.n6713 VSS 0.451316f
C23956 DVDD.n6714 VSS 0.451316f
C23957 DVDD.n6715 VSS 0.451316f
C23958 DVDD.n6716 VSS 0.451316f
C23959 DVDD.n6717 VSS 0.451316f
C23960 DVDD.n6718 VSS 0.451316f
C23961 DVDD.n6719 VSS 0.451316f
C23962 DVDD.n6720 VSS 0.451316f
C23963 DVDD.n6721 VSS 0.451316f
C23964 DVDD.n6722 VSS 0.451316f
C23965 DVDD.n6723 VSS 0.451316f
C23966 DVDD.n6724 VSS 0.451316f
C23967 DVDD.n6725 VSS 0.451316f
C23968 DVDD.n6726 VSS 0.451316f
C23969 DVDD.n6727 VSS 0.451316f
C23970 DVDD.n6728 VSS 0.451316f
C23971 DVDD.n6729 VSS 0.197054f
C23972 DVDD.n6730 VSS 0.451316f
C23973 DVDD.n6731 VSS 0.197054f
C23974 DVDD.n6732 VSS 0.451316f
C23975 DVDD.n6733 VSS 0.402053f
C23976 DVDD.n6734 VSS 0.451316f
C23977 DVDD.n6735 VSS 0.451316f
C23978 DVDD.n6736 VSS 0.451316f
C23979 DVDD.n6737 VSS 0.451316f
C23980 DVDD.n6738 VSS 0.451316f
C23981 DVDD.n6739 VSS 0.451316f
C23982 DVDD.n6740 VSS 0.451316f
C23983 DVDD.n6741 VSS 0.451316f
C23984 DVDD.n6742 VSS 0.451316f
C23985 DVDD.n6743 VSS 0.451316f
C23986 DVDD.n6744 VSS 0.451316f
C23987 DVDD.n6745 VSS 0.360735f
C23988 DVDD.n6746 VSS 0.375037f
C23989 DVDD.n6747 VSS 0.375037f
C23990 DVDD.n6748 VSS 0.543486f
C23991 DVDD.n6749 VSS 0.301937f
C23992 DVDD.n6750 VSS 0.408409f
C23993 DVDD.n6751 VSS 0.182751f
C23994 DVDD.n6752 VSS 0.301937f
C23995 DVDD.n6753 VSS 0.451316f
C23996 DVDD.n6754 VSS 0.197054f
C23997 DVDD.n6765 VSS 0.225658f
C23998 DVDD.n6767 VSS 0.127013f
C23999 DVDD.n6768 VSS 0.225658f
C24000 DVDD.n6769 VSS 0.559179f
C24001 DVDD.n6770 VSS 0.559179f
C24002 DVDD.n6771 VSS 0.120351f
C24003 DVDD.n6772 VSS 0.128627f
C24004 DVDD.n6773 VSS 0.128627f
C24005 DVDD.n6774 VSS 0.225658f
C24006 DVDD.n6775 VSS 1.85083f
C24007 DVDD.n6776 VSS 1.85083f
C24008 DVDD.n6777 VSS 0.456124f
C24009 DVDD.n6778 VSS 0.029062f
C24010 DVDD.n6779 VSS 0.060739f
C24011 DVDD.n6780 VSS 0.02691f
C24012 DVDD.n6781 VSS 0.029062f
C24013 DVDD.n6782 VSS 0.033368f
C24014 DVDD.n6783 VSS 0.114418f
C24015 DVDD.n6784 VSS 0.114418f
C24016 DVDD.n6785 VSS 0.114418f
C24017 DVDD.n6786 VSS 0.030408f
C24018 DVDD.n6787 VSS 0.029062f
C24019 DVDD.n6788 VSS 0.225658f
C24020 DVDD.n6789 VSS 0.066735f
C24021 DVDD.n6790 VSS 0.066735f
C24022 DVDD.n6791 VSS 0.225658f
C24023 DVDD.n6792 VSS 0.029062f
C24024 DVDD.n6793 VSS 0.033368f
C24025 DVDD.n6794 VSS 0.029062f
C24026 DVDD.n6795 VSS 0.033368f
C24027 DVDD.n6796 VSS 0.15585f
C24028 DVDD.t12 VSS 5.27557f
C24029 DVDD.n6797 VSS 0.15585f
C24030 DVDD.n6798 VSS 0.277706f
C24031 DVDD.n6799 VSS 0.058124f
C24032 DVDD.n6800 VSS 0.114418f
C24033 DVDD.n6801 VSS 0.058124f
C24034 DVDD.n6802 VSS 0.114418f
C24035 DVDD.n6803 VSS 0.058124f
C24036 DVDD.n6804 VSS 0.114418f
C24037 DVDD.n6805 VSS 0.058124f
C24038 DVDD.n6806 VSS 0.114418f
C24039 DVDD.n6807 VSS 0.058124f
C24040 DVDD.n6808 VSS 0.114418f
C24041 DVDD.n6809 VSS 0.058124f
C24042 DVDD.n6810 VSS 0.114418f
C24043 DVDD.n6811 VSS 0.114418f
C24044 DVDD.n6812 VSS 0.058124f
C24045 DVDD.n6813 VSS 0.058124f
C24046 DVDD.n6814 VSS 0.058124f
C24047 DVDD.n6815 VSS 0.114418f
C24048 DVDD.n6816 VSS 0.114418f
C24049 DVDD.n6817 VSS 0.114418f
C24050 DVDD.n6818 VSS 0.058124f
C24051 DVDD.n6819 VSS 0.058124f
C24052 DVDD.n6820 VSS 0.058124f
C24053 DVDD.n6821 VSS 0.114418f
C24054 DVDD.n6822 VSS 0.114418f
C24055 DVDD.n6823 VSS 0.114418f
C24056 DVDD.n6824 VSS 0.058124f
C24057 DVDD.n6825 VSS 0.058124f
C24058 DVDD.n6826 VSS 0.058124f
C24059 DVDD.n6827 VSS 0.114418f
C24060 DVDD.n6828 VSS 0.114418f
C24061 DVDD.n6829 VSS 0.114418f
C24062 DVDD.n6830 VSS 0.058124f
C24063 DVDD.n6831 VSS 0.058124f
C24064 DVDD.n6832 VSS 0.058124f
C24065 DVDD.n6833 VSS 0.114418f
C24066 DVDD.n6834 VSS 0.114418f
C24067 DVDD.n6835 VSS 0.114418f
C24068 DVDD.n6836 VSS 0.058124f
C24069 DVDD.n6837 VSS 0.058124f
C24070 DVDD.n6838 VSS 0.058124f
C24071 DVDD.n6839 VSS 0.114418f
C24072 DVDD.n6840 VSS 0.114418f
C24073 DVDD.n6841 VSS 0.114418f
C24074 DVDD.n6842 VSS 0.058124f
C24075 DVDD.n6843 VSS 0.058124f
C24076 DVDD.n6844 VSS 0.058124f
C24077 DVDD.n6845 VSS 0.114418f
C24078 DVDD.n6846 VSS 0.114418f
C24079 DVDD.n6847 VSS 0.114418f
C24080 DVDD.n6848 VSS 0.058124f
C24081 DVDD.n6849 VSS 0.058124f
C24082 DVDD.n6850 VSS 0.277706f
C24083 DVDD.n6851 VSS 0.15585f
C24084 DVDD.t40 VSS 5.27557f
C24085 DVDD.n6852 VSS 0.15585f
C24086 DVDD.n6853 VSS 0.156344f
C24087 DVDD.n6855 VSS 0.16065f
C24088 DVDD.n6856 VSS 0.225658f
C24089 DVDD.n6857 VSS 0.029062f
C24090 DVDD.n6858 VSS 0.033368f
C24091 DVDD.n6859 VSS 0.15585f
C24092 DVDD.t18 VSS 5.27557f
C24093 DVDD.n6860 VSS 0.15585f
C24094 DVDD.n6861 VSS 0.029062f
C24095 DVDD.n6862 VSS 0.033368f
C24096 DVDD.n6863 VSS 0.114418f
C24097 DVDD.n6864 VSS 0.114418f
C24098 DVDD.n6865 VSS 0.033368f
C24099 DVDD.n6866 VSS 0.029062f
C24100 DVDD.n6867 VSS 0.060739f
C24101 DVDD.n6868 VSS 0.061117f
C24102 DVDD.n6869 VSS 0.173937f
C24103 DVDD.n6870 VSS 0.060175f
C24104 DVDD.n6871 VSS 0.026274f
C24105 DVDD.n6872 VSS 0.030088f
C24106 DVDD.n6873 VSS 0.061085f
C24107 DVDD.n6875 VSS 0.066735f
C24108 DVDD.n6877 VSS 0.066735f
C24109 DVDD.n6878 VSS 0.030088f
C24110 DVDD.n6879 VSS 0.026274f
C24111 DVDD.n6880 VSS 0.044284f
C24112 DVDD.n6881 VSS 0.044284f
C24113 DVDD.n6882 VSS 0.172475f
C24114 DVDD.n6883 VSS 0.045979f
C24115 DVDD.n6884 VSS 0.045979f
C24116 DVDD.n6885 VSS 0.026274f
C24117 DVDD.n6886 VSS 0.026274f
C24118 DVDD.n6887 VSS 0.030088f
C24119 DVDD.n6888 VSS 0.066735f
C24120 DVDD.n6890 VSS 0.066735f
C24121 DVDD.n6893 VSS 0.066735f
C24122 DVDD.n6894 VSS 0.029028f
C24123 DVDD.n6895 VSS 0.026274f
C24124 DVDD.n6896 VSS 0.060175f
C24125 DVDD.n6897 VSS 0.170687f
C24126 DVDD.n6898 VSS 0.057655f
C24127 DVDD.n6899 VSS 0.059611f
C24128 DVDD.n6900 VSS 0.029062f
C24129 DVDD.n6901 VSS 0.033368f
C24130 DVDD.n6902 VSS 0.15585f
C24131 DVDD.t28 VSS 5.27557f
C24132 DVDD.n6903 VSS 0.033368f
C24133 DVDD.n6904 VSS 0.15585f
C24134 DVDD.n6905 VSS 0.033368f
C24135 DVDD.n6906 VSS 0.114418f
C24136 DVDD.n6907 VSS 0.033368f
C24137 DVDD.n6908 VSS 0.114418f
C24138 DVDD.n6909 VSS 0.033368f
C24139 DVDD.n6910 VSS 0.114418f
C24140 DVDD.n6911 VSS 0.033368f
C24141 DVDD.n6912 VSS 0.114418f
C24142 DVDD.n6913 VSS 0.114418f
C24143 DVDD.n6914 VSS 0.032561f
C24144 DVDD.n6915 VSS 0.029869f
C24145 DVDD.n6916 VSS 0.114418f
C24146 DVDD.n6917 VSS 0.033368f
C24147 DVDD.n6918 VSS 0.114418f
C24148 DVDD.n6919 VSS 0.033368f
C24149 DVDD.n6920 VSS 0.114418f
C24150 DVDD.n6921 VSS 0.114418f
C24151 DVDD.n6922 VSS 0.033368f
C24152 DVDD.n6923 VSS 0.029062f
C24153 DVDD.n6924 VSS 0.225658f
C24154 DVDD.n6925 VSS 0.029062f
C24155 DVDD.n6926 VSS 0.033368f
C24156 DVDD.n6927 VSS 0.15585f
C24157 DVDD.t5 VSS 5.27557f
C24158 DVDD.n6928 VSS 0.033368f
C24159 DVDD.n6929 VSS 0.15585f
C24160 DVDD.n6930 VSS 0.114418f
C24161 DVDD.n6931 VSS 0.033368f
C24162 DVDD.n6932 VSS 0.029062f
C24163 DVDD.n6934 VSS 0.225658f
C24164 DVDD.n6935 VSS 0.197054f
C24165 DVDD.n6936 VSS 0.066735f
C24166 DVDD.n6937 VSS 0.066735f
C24167 DVDD.n6938 VSS 0.066735f
C24168 DVDD.n6939 VSS 0.360735f
C24169 DVDD.n6940 VSS 0.066735f
C24170 DVDD.n6941 VSS 0.066735f
C24171 DVDD.n6942 VSS 0.451316f
C24172 DVDD.n6943 VSS 0.451316f
C24173 DVDD.n6944 VSS 0.451316f
C24174 DVDD.n6945 VSS 0.451316f
C24175 DVDD.n6946 VSS 0.451316f
C24176 DVDD.n6947 VSS 0.451316f
C24177 DVDD.n6948 VSS 0.451316f
C24178 DVDD.n6949 VSS 0.451316f
C24179 DVDD.n6950 VSS 0.451316f
C24180 DVDD.n6951 VSS 0.451316f
C24181 DVDD.n6952 VSS 0.451316f
C24182 DVDD.n6953 VSS 0.451316f
C24183 DVDD.n6954 VSS 0.451316f
C24184 DVDD.n6955 VSS 0.451316f
C24185 DVDD.n6956 VSS 0.451316f
C24186 DVDD.n6957 VSS 0.451316f
C24187 DVDD.n6958 VSS 0.451316f
C24188 DVDD.n6959 VSS 0.451316f
C24189 DVDD.n6960 VSS 0.451316f
C24190 DVDD.n6961 VSS 0.451316f
C24191 DVDD.n6962 VSS 0.451316f
C24192 DVDD.n6963 VSS 0.451316f
C24193 DVDD.n6964 VSS 0.451316f
C24194 DVDD.n6965 VSS 0.451316f
C24195 DVDD.n6966 VSS 0.451316f
C24196 DVDD.n6967 VSS 0.451316f
C24197 DVDD.n6968 VSS 0.451316f
C24198 DVDD.n6969 VSS 0.451316f
C24199 DVDD.n6970 VSS 0.451316f
C24200 DVDD.n6971 VSS 0.451316f
C24201 DVDD.n6972 VSS 0.451316f
C24202 DVDD.n6973 VSS 0.451316f
C24203 DVDD.n6974 VSS 0.451316f
C24204 DVDD.n6975 VSS 0.451316f
C24205 DVDD.n6976 VSS 0.197054f
C24206 DVDD.n6979 VSS 0.225658f
C24207 DVDD.n6981 VSS 0.066735f
C24208 DVDD.n6982 VSS 0.225658f
C24209 DVDD.n6983 VSS 0.066735f
C24210 DVDD.n6985 VSS 0.225658f
C24211 DVDD.n6986 VSS 0.402053f
C24212 DVDD.n6987 VSS 0.451316f
C24213 DVDD.n6988 VSS 0.451316f
C24214 DVDD.n6989 VSS 0.451316f
C24215 DVDD.n6990 VSS 0.451316f
C24216 DVDD.n6991 VSS 0.451316f
C24217 DVDD.n6992 VSS 0.451316f
C24218 DVDD.n6993 VSS 0.451316f
C24219 DVDD.n6994 VSS 0.451316f
C24220 DVDD.n6995 VSS 0.451316f
C24221 DVDD.n6996 VSS 0.451316f
C24222 DVDD.n6997 VSS 0.451316f
C24223 DVDD.n6998 VSS 0.360735f
C24224 DVDD.n6999 VSS 0.375037f
C24225 DVDD.n7000 VSS 0.861315f
C24226 DVDD.n7001 VSS 0.301937f
C24227 DVDD.n7002 VSS 0.182751f
C24228 DVDD.n7003 VSS 0.225658f
C24229 DVDD.n7004 VSS 0.127013f
C24230 DVDD.n7005 VSS 0.225658f
C24231 DVDD.n7006 VSS 0.402053f
C24232 DVDD.n7007 VSS 0.451316f
C24233 DVDD.n7008 VSS 0.451316f
C24234 DVDD.n7009 VSS 0.451316f
C24235 DVDD.n7010 VSS 0.451316f
C24236 DVDD.n7011 VSS 0.451316f
C24237 DVDD.n7012 VSS 0.360735f
C24238 DVDD.n7013 VSS 0.451316f
C24239 DVDD.n7014 VSS 0.197054f
C24240 DVDD.n7015 VSS 0.451316f
C24241 DVDD.n7016 VSS 0.451316f
C24242 DVDD.n7017 VSS 0.197054f
C24243 DVDD.n7020 VSS 0.225658f
C24244 DVDD.n7023 VSS 0.066735f
C24245 DVDD.n7024 VSS 2.63355f
C24246 DVDD.n7025 VSS 0.127013f
C24247 DVDD.n7026 VSS 0.127013f
C24248 DVDD.n7029 VSS 0.225658f
C24249 DVDD.n7030 VSS 0.225658f
C24250 DVDD.n7031 VSS 2.66323f
C24251 DVDD.n7032 VSS 0.066735f
C24252 DVDD.n7033 VSS 0.066735f
C24253 DVDD.n7034 VSS 0.066735f
C24254 DVDD.n7035 VSS 0.066735f
C24255 DVDD.n7036 VSS 0.066735f
C24256 DVDD.n7037 VSS 0.066735f
C24257 DVDD.n7038 VSS 0.066735f
C24258 DVDD.n7039 VSS 0.066735f
C24259 DVDD.n7040 VSS 0.066735f
C24260 DVDD.n7041 VSS 0.066735f
C24261 DVDD.n7042 VSS 0.066735f
C24262 DVDD.n7043 VSS 0.197054f
C24263 DVDD.n7045 VSS 0.066735f
C24264 DVDD.n7047 VSS 0.066735f
C24265 DVDD.n7049 VSS 0.066735f
C24266 DVDD.n7051 VSS 0.066735f
C24267 DVDD.n7053 VSS 0.066735f
C24268 DVDD.n7055 VSS 0.066735f
C24269 DVDD.n7057 VSS 0.066735f
C24270 DVDD.n7059 VSS 0.066735f
C24271 DVDD.n7061 VSS 0.066735f
C24272 DVDD.n7063 VSS 0.066735f
C24273 DVDD.n7065 VSS 0.066735f
C24274 DVDD.n7068 VSS 0.105307f
C24275 DVDD.n7069 VSS 0.105307f
C24276 DVDD.n7070 VSS 1.28462f
C24277 DVDD.n7071 VSS 0.066735f
C24278 DVDD.n7072 VSS 0.066735f
C24279 DVDD.n7073 VSS 0.066735f
C24280 DVDD.n7074 VSS 0.066735f
C24281 DVDD.n7075 VSS 0.066735f
C24282 DVDD.n7076 VSS 0.091958f
C24283 DVDD.n7078 VSS 0.066735f
C24284 DVDD.n7080 VSS 0.066735f
C24285 DVDD.n7082 VSS 0.066735f
C24286 DVDD.n7084 VSS 0.066735f
C24287 DVDD.n7090 VSS 0.420368f
C24288 DVDD.n7091 VSS 0.091958f
C24289 DVDD.n7092 VSS 0.210614f
C24290 DVDD.n7093 VSS 0.210614f
C24291 DVDD.n7094 VSS 0.210614f
C24292 DVDD.n7095 VSS 0.210614f
C24293 DVDD.n7096 VSS 0.210614f
C24294 DVDD.n7097 VSS 0.210614f
C24295 DVDD.n7098 VSS 0.210614f
C24296 DVDD.n7099 VSS 0.066735f
C24297 DVDD.n7100 VSS 0.066735f
C24298 DVDD.n7101 VSS 0.066735f
C24299 DVDD.n7102 VSS 0.066735f
C24300 DVDD.n7103 VSS 0.066735f
C24301 DVDD.n7104 VSS 0.091958f
C24302 DVDD.n7106 VSS 0.149379f
C24303 DVDD.n7107 VSS 0.225658f
C24304 DVDD.n7108 VSS 0.402053f
C24305 DVDD.n7109 VSS 0.066735f
C24306 DVDD.n7110 VSS 0.066735f
C24307 DVDD.n7111 VSS 0.05059f
C24308 DVDD.n7112 VSS 0.033368f
C24309 DVDD.n7113 VSS 0.049513f
C24310 DVDD.n7114 VSS 0.066735f
C24311 DVDD.n7115 VSS 0.066735f
C24312 DVDD.n7116 VSS 0.066735f
C24313 DVDD.n7117 VSS 0.066735f
C24314 DVDD.n7118 VSS 0.066735f
C24315 DVDD.n7119 VSS 0.066735f
C24316 DVDD.n7120 VSS 0.197054f
C24317 DVDD.n7122 VSS 0.066735f
C24318 DVDD.n7124 VSS 0.066735f
C24319 DVDD.n7126 VSS 0.066735f
C24320 DVDD.n7128 VSS 0.066735f
C24321 DVDD.n7130 VSS 0.066735f
C24322 DVDD.n7132 VSS 0.066735f
C24323 DVDD.n7134 VSS 0.066735f
C24324 DVDD.n7135 VSS 0.033368f
C24325 DVDD.n7136 VSS 0.033368f
C24326 DVDD.n7137 VSS 0.033368f
C24327 DVDD.n7138 VSS 0.033368f
C24328 DVDD.n7140 VSS 0.061481f
C24329 DVDD.n7142 VSS 0.061481f
C24330 DVDD.n7143 VSS 0.033368f
C24331 DVDD.n7145 VSS 0.033368f
C24332 DVDD.n7146 VSS 0.061481f
C24333 DVDD.n7148 VSS 0.061481f
C24334 DVDD.n7149 VSS 0.033368f
C24335 DVDD.n7151 VSS 0.033368f
C24336 DVDD.n7152 VSS 0.033368f
C24337 DVDD.n7154 VSS 0.061481f
C24338 DVDD.n7156 VSS 0.061481f
C24339 DVDD.n7157 VSS 0.033368f
C24340 DVDD.n7158 VSS 0.033368f
C24341 DVDD.n7160 VSS 0.061481f
C24342 DVDD.n7162 VSS 0.061481f
C24343 DVDD.n7164 VSS 0.033368f
C24344 DVDD.n7165 VSS 0.033368f
C24345 DVDD.n7166 VSS 0.033368f
C24346 DVDD.n7168 VSS 0.061481f
C24347 DVDD.n7170 VSS 0.061481f
C24348 DVDD.n7171 VSS 0.033368f
C24349 DVDD.n7172 VSS 0.360951f
C24350 DVDD.n7173 VSS 0.033368f
C24351 DVDD.n7175 VSS 0.360951f
C24352 DVDD.n7176 VSS 0.033368f
C24353 DVDD.n7177 VSS 0.501762f
C24354 DVDD.n7178 VSS 0.033368f
C24355 DVDD.n7180 VSS 0.501762f
C24356 DVDD.n7181 VSS 0.033368f
C24357 DVDD.n7182 VSS 0.316328f
C24358 DVDD.n7183 VSS -2.30734f
C24359 DVDD.n7184 VSS 0.316328f
C24360 DVDD.n7185 VSS 0.033368f
C24361 DVDD.n7186 VSS 0.501762f
C24362 DVDD.n7187 VSS 0.033368f
C24363 DVDD.n7189 VSS 0.501762f
C24364 DVDD.n7190 VSS 0.033368f
C24365 DVDD.n7191 VSS 0.360951f
C24366 DVDD.n7192 VSS 0.360951f
C24367 DVDD.n7194 VSS 0.033368f
C24368 DVDD.n7195 VSS 0.061481f
C24369 DVDD.n7197 VSS 0.033368f
C24370 DVDD.n7198 VSS 0.061481f
C24371 DVDD.n7200 VSS 0.970017f
C24372 DVDD.n7201 VSS 0.033368f
C24373 DVDD.n7202 VSS 0.033368f
C24374 DVDD.n7204 VSS 0.066735f
C24375 DVDD.n7205 VSS 0.451316f
C24376 DVDD.n7206 VSS 0.451316f
C24377 DVDD.n7207 VSS 0.451316f
C24378 DVDD.n7208 VSS 0.360735f
C24379 DVDD.n7209 VSS 0.451316f
C24380 DVDD.n7210 VSS 3.1729f
C24381 DVDD.n7211 VSS 0.929942f
C24382 DVDD.n7222 VSS 0.225658f
C24383 DVDD.n7223 VSS 0.197054f
C24384 DVDD.n7224 VSS 0.451316f
C24385 DVDD.n7225 VSS 0.197054f
C24386 DVDD.n7226 VSS 0.451316f
C24387 DVDD.n7227 VSS 0.451316f
C24388 DVDD.n7228 VSS 0.451316f
C24389 DVDD.n7229 VSS 0.451316f
C24390 DVDD.n7230 VSS 0.451316f
C24391 DVDD.n7231 VSS 0.451316f
C24392 DVDD.n7232 VSS 0.451316f
C24393 DVDD.n7233 VSS 0.451316f
C24394 DVDD.n7234 VSS 0.451316f
C24395 DVDD.n7235 VSS 0.451316f
C24396 DVDD.n7236 VSS 0.451316f
C24397 DVDD.n7237 VSS 0.451316f
C24398 DVDD.n7238 VSS 0.451316f
C24399 DVDD.n7239 VSS 0.451316f
C24400 DVDD.n7240 VSS 0.301937f
C24401 DVDD.n7241 VSS 0.375037f
C24402 DVDD.n7242 VSS 0.451316f
C24403 DVDD.n7243 VSS 0.451316f
C24404 DVDD.n7244 VSS 0.451316f
C24405 DVDD.n7245 VSS 0.451316f
C24406 DVDD.n7246 VSS 0.451316f
C24407 DVDD.n7247 VSS 0.451316f
C24408 DVDD.n7248 VSS 0.451316f
C24409 DVDD.n7249 VSS 0.451316f
C24410 DVDD.n7250 VSS 0.451316f
C24411 DVDD.n7251 VSS 0.451316f
C24412 DVDD.n7252 VSS 0.451316f
C24413 DVDD.n7253 VSS 0.451316f
C24414 DVDD.n7254 VSS 0.451316f
C24415 DVDD.n7255 VSS 0.451316f
C24416 DVDD.n7256 VSS 0.451316f
C24417 DVDD.n7257 VSS 0.451316f
C24418 DVDD.n7258 VSS 0.451316f
C24419 DVDD.n7259 VSS 0.451316f
C24420 DVDD.n7260 VSS 0.451316f
C24421 DVDD.n7261 VSS 0.451316f
C24422 DVDD.n7262 VSS 0.451316f
C24423 DVDD.n7263 VSS 0.451316f
C24424 DVDD.n7264 VSS 0.451316f
C24425 DVDD.n7265 VSS 0.451316f
C24426 DVDD.n7266 VSS 0.360735f
C24427 DVDD.n7267 VSS 0.375037f
C24428 DVDD.n7268 VSS 0.543486f
C24429 DVDD.n7269 VSS 0.182751f
C24430 DVDD.n7270 VSS 0.301937f
C24431 DVDD.n7271 VSS 0.451316f
C24432 DVDD.n7272 VSS 0.197054f
C24433 DVDD.n7281 VSS 0.225658f
C24434 DVDD.n7284 VSS 0.066735f
C24435 DVDD.n7285 VSS 0.225658f
C24436 DVDD.n7286 VSS 0.559179f
C24437 DVDD.n7287 VSS 0.559179f
C24438 DVDD.n7288 VSS 0.066735f
C24439 DVDD.n7289 VSS 0.066735f
C24440 DVDD.n7290 VSS 0.066735f
C24441 DVDD.n7291 VSS 0.066735f
C24442 DVDD.n7298 VSS 0.105307f
C24443 DVDD.n7299 VSS 0.091958f
C24444 DVDD.n7304 VSS 0.105307f
C24445 DVDD.n7305 VSS 0.210614f
C24446 DVDD.n7306 VSS 0.210614f
C24447 DVDD.n7307 VSS 0.210614f
C24448 DVDD.n7308 VSS 0.210614f
C24449 DVDD.n7309 VSS 0.210614f
C24450 DVDD.n7310 VSS 0.168343f
C24451 DVDD.n7311 VSS 0.210614f
C24452 DVDD.n7312 VSS 0.210614f
C24453 DVDD.n7313 VSS 0.210614f
C24454 DVDD.n7314 VSS 0.210614f
C24455 DVDD.n7315 VSS 0.210614f
C24456 DVDD.n7316 VSS 0.210614f
C24457 DVDD.n7317 VSS 0.210614f
C24458 DVDD.n7318 VSS 0.210614f
C24459 DVDD.n7319 VSS 0.210614f
C24460 DVDD.n7320 VSS 0.168343f
C24461 DVDD.n7321 VSS 0.210614f
C24462 DVDD.n7322 VSS 0.210614f
C24463 DVDD.n7323 VSS 0.210614f
C24464 DVDD.n7324 VSS 0.210614f
C24465 DVDD.n7325 VSS 0.210614f
C24466 DVDD.n7326 VSS 0.210614f
C24467 DVDD.n7327 VSS 0.210614f
C24468 DVDD.n7328 VSS 0.210614f
C24469 DVDD.n7329 VSS 0.187625f
C24470 DVDD.n7330 VSS 0.210614f
C24471 DVDD.n7331 VSS 0.210614f
C24472 DVDD.n7332 VSS 0.210614f
C24473 DVDD.n7333 VSS 0.105307f
C24474 DVDD.n7339 VSS 0.091958f
C24475 DVDD.n7342 VSS 0.066735f
C24476 DVDD.n7344 VSS 0.061481f
C24477 DVDD.n7347 VSS 0.0127f
C24478 DVDD.n7348 VSS 0.0127f
C24479 DVDD.n7349 VSS 0.025401f
C24480 DVDD.n7351 VSS 0.025401f
C24481 DVDD.n7352 VSS 0.229078f
C24482 DVDD.n7353 VSS 0.229078f
C24483 DVDD.n7354 VSS 0.0127f
C24484 DVDD.n7355 VSS 0.025401f
C24485 DVDD.n7356 VSS 0.0127f
C24486 DVDD.n7357 VSS 0.025401f
C24487 DVDD.n7358 VSS 0.348208f
C24488 DVDD.n7359 VSS 0.352514f
C24489 DVDD.n7361 VSS 0.066735f
C24490 DVDD.n7362 VSS 0.061481f
C24491 DVDD.n7363 VSS 0.638831f
C24492 DVDD.n7364 VSS 0.066735f
C24493 DVDD.n7365 VSS 0.066735f
C24494 DVDD.n7366 VSS 0.066735f
C24495 DVDD.n7367 VSS 0.066735f
C24496 DVDD.n7368 VSS 0.066735f
C24497 DVDD.n7369 VSS 0.091958f
C24498 DVDD.n7370 VSS 0.066735f
C24499 DVDD.n7371 VSS 0.066735f
C24500 DVDD.n7372 VSS 0.066735f
C24501 DVDD.n7373 VSS 0.210614f
C24502 DVDD.n7374 VSS 0.210614f
C24503 DVDD.n7375 VSS 0.210614f
C24504 DVDD.n7376 VSS 0.210614f
C24505 DVDD.n7377 VSS 0.210614f
C24506 DVDD.n7378 VSS 0.210614f
C24507 DVDD.n7379 VSS 0.210614f
C24508 DVDD.n7380 VSS 0.210614f
C24509 DVDD.n7381 VSS 0.210614f
C24510 DVDD.n7382 VSS 0.210614f
C24511 DVDD.n7383 VSS 0.210614f
C24512 DVDD.n7384 VSS 0.210614f
C24513 DVDD.n7385 VSS 0.210614f
C24514 DVDD.n7386 VSS 0.210614f
C24515 DVDD.n7387 VSS 0.210614f
C24516 DVDD.n7388 VSS 0.210614f
C24517 DVDD.n7389 VSS 0.210614f
C24518 DVDD.n7390 VSS 0.210614f
C24519 DVDD.n7391 VSS 0.210614f
C24520 DVDD.n7392 VSS 0.210614f
C24521 DVDD.n7393 VSS 0.210614f
C24522 DVDD.n7394 VSS 0.210614f
C24523 DVDD.n7395 VSS 0.210614f
C24524 DVDD.n7396 VSS 0.210614f
C24525 DVDD.n7397 VSS 0.210614f
C24526 DVDD.n7398 VSS 0.210614f
C24527 DVDD.n7399 VSS 0.210614f
C24528 DVDD.n7400 VSS 0.210614f
C24529 DVDD.n7401 VSS 0.210614f
C24530 DVDD.n7402 VSS 0.210614f
C24531 DVDD.n7403 VSS 0.210614f
C24532 DVDD.n7404 VSS 0.210614f
C24533 DVDD.n7405 VSS 0.210614f
C24534 DVDD.n7406 VSS 0.210614f
C24535 DVDD.n7407 VSS 0.210614f
C24536 DVDD.n7408 VSS 0.210614f
C24537 DVDD.n7409 VSS 0.210614f
C24538 DVDD.n7410 VSS 0.210614f
C24539 DVDD.n7411 VSS 0.210614f
C24540 DVDD.n7412 VSS 0.210614f
C24541 DVDD.n7413 VSS 0.210614f
C24542 DVDD.n7414 VSS 0.210614f
C24543 DVDD.n7415 VSS 0.210614f
C24544 DVDD.n7416 VSS 0.210614f
C24545 DVDD.n7417 VSS 0.210614f
C24546 DVDD.n7418 VSS 0.210614f
C24547 DVDD.n7419 VSS 0.210614f
C24548 DVDD.n7420 VSS 0.210614f
C24549 DVDD.n7421 VSS 0.168343f
C24550 DVDD.n7425 VSS 0.105307f
C24551 DVDD.n7427 VSS 0.066735f
C24552 DVDD.n7428 VSS 0.105307f
C24553 DVDD.n7429 VSS 0.638831f
C24554 DVDD.n7430 VSS 0.105307f
C24555 DVDD.n7431 VSS 0.091958f
C24556 DVDD.n7432 VSS 0.210614f
C24557 DVDD.n7433 VSS 0.210614f
C24558 DVDD.n7434 VSS 0.210614f
C24559 DVDD.n7435 VSS 0.210614f
C24560 DVDD.n7436 VSS 0.210614f
C24561 DVDD.n7437 VSS 0.210614f
C24562 DVDD.n7438 VSS 0.210614f
C24563 DVDD.n7439 VSS 0.210614f
C24564 DVDD.n7440 VSS 0.210614f
C24565 DVDD.n7441 VSS 0.210614f
C24566 DVDD.n7442 VSS 0.210614f
C24567 DVDD.n7443 VSS 0.210614f
C24568 DVDD.n7444 VSS 0.210614f
C24569 DVDD.n7445 VSS 0.210614f
C24570 DVDD.n7446 VSS 0.210614f
C24571 DVDD.n7447 VSS 0.210614f
C24572 DVDD.n7448 VSS 0.210614f
C24573 DVDD.n7449 VSS 0.210614f
C24574 DVDD.n7450 VSS 0.210614f
C24575 DVDD.n7451 VSS 0.210614f
C24576 DVDD.n7452 VSS 0.210614f
C24577 DVDD.n7453 VSS 0.210614f
C24578 DVDD.n7454 VSS 0.210614f
C24579 DVDD.n7455 VSS 0.210614f
C24580 DVDD.n7456 VSS 0.210614f
C24581 DVDD.n7457 VSS 0.210614f
C24582 DVDD.n7458 VSS 0.210614f
C24583 DVDD.n7459 VSS 0.210614f
C24584 DVDD.n7460 VSS 0.091958f
C24585 DVDD.n7461 VSS 0.210614f
C24586 DVDD.n7462 VSS 0.210614f
C24587 DVDD.n7463 VSS 0.210614f
C24588 DVDD.n7464 VSS 0.210614f
C24589 DVDD.n7465 VSS 0.210614f
C24590 DVDD.n7466 VSS 0.210614f
C24591 DVDD.n7467 VSS 0.210614f
C24592 DVDD.n7468 VSS 0.210614f
C24593 DVDD.n7469 VSS 0.210614f
C24594 DVDD.n7470 VSS 0.210614f
C24595 DVDD.n7471 VSS 0.210614f
C24596 DVDD.n7472 VSS 0.210614f
C24597 DVDD.n7473 VSS 0.210614f
C24598 DVDD.n7474 VSS 0.210614f
C24599 DVDD.n7475 VSS 0.210614f
C24600 DVDD.n7476 VSS 0.210614f
C24601 DVDD.n7477 VSS 0.210614f
C24602 DVDD.n7478 VSS 0.210614f
C24603 DVDD.n7479 VSS 0.210614f
C24604 DVDD.n7480 VSS 0.210614f
C24605 DVDD.n7481 VSS 0.210614f
C24606 DVDD.n7482 VSS 0.210614f
C24607 DVDD.n7483 VSS 0.210614f
C24608 DVDD.n7484 VSS 0.091958f
C24609 DVDD.n7485 VSS 0.105307f
C24610 DVDD.n7486 VSS 0.638831f
C24611 DVDD.n7487 VSS 0.105307f
C24612 DVDD.n7488 VSS 0.187625f
C24613 DVDD.n7489 VSS 0.210614f
C24614 DVDD.n7490 VSS 0.210614f
C24615 DVDD.n7491 VSS 0.210614f
C24616 DVDD.n7492 VSS 0.210614f
C24617 DVDD.n7493 VSS 0.210614f
C24618 DVDD.n7494 VSS 0.210614f
C24619 DVDD.n7495 VSS 0.210614f
C24620 DVDD.n7496 VSS 0.168343f
C24621 DVDD.n7497 VSS 0.210614f
C24622 DVDD.n7498 VSS 0.210614f
C24623 DVDD.n7499 VSS 0.210614f
C24624 DVDD.n7500 VSS 1.46996f
C24625 DVDD.n7501 VSS 0.210614f
C24626 DVDD.n7502 VSS 0.091958f
C24627 DVDD.n7503 VSS 0.105307f
C24628 DVDD.n7504 VSS 5.4567f
C24629 DVDD.n7505 VSS 1.20568f
C24630 DVDD.n7506 VSS 0.559179f
C24631 DVDD.n7507 VSS 0.559179f
C24632 DVDD.n7508 VSS 2.62099f
C24633 DVDD.n7509 VSS 0.127013f
C24634 DVDD.n7510 VSS 2.66633f
C24635 DVDD.n7511 VSS 0.066735f
C24636 DVDD.n7512 VSS 0.066735f
C24637 DVDD.n7513 VSS 0.066735f
C24638 DVDD.n7514 VSS 0.066735f
C24639 DVDD.n7515 VSS 0.066735f
C24640 DVDD.n7516 VSS 0.066735f
C24641 DVDD.n7517 VSS 0.066735f
C24642 DVDD.n7518 VSS 0.066735f
C24643 DVDD.n7519 VSS 0.066735f
C24644 DVDD.n7520 VSS 0.066735f
C24645 DVDD.n7521 VSS 0.066735f
C24646 DVDD.n7522 VSS 0.930088f
C24647 DVDD.n7523 VSS 0.197054f
C24648 DVDD.n7524 VSS 0.066735f
C24649 DVDD.n7525 VSS 0.066735f
C24650 DVDD.n7526 VSS 0.066735f
C24651 DVDD.n7527 VSS 0.066735f
C24652 DVDD.n7528 VSS 0.066735f
C24653 DVDD.n7529 VSS 0.066735f
C24654 DVDD.n7530 VSS 0.066735f
C24655 DVDD.n7531 VSS 0.066735f
C24656 DVDD.n7532 VSS 0.066735f
C24657 DVDD.n7533 VSS 0.066735f
C24658 DVDD.n7534 VSS 0.197054f
C24659 DVDD.n7545 VSS 0.225658f
C24660 DVDD.n7547 VSS 0.066735f
C24661 DVDD.n7548 VSS 2.63355f
C24662 DVDD.n7549 VSS 0.127013f
C24663 DVDD.n7550 VSS 0.225658f
C24664 DVDD.n7551 VSS 0.197054f
C24665 DVDD.n7552 VSS 0.451316f
C24666 DVDD.n7553 VSS 0.451316f
C24667 DVDD.n7554 VSS 0.451316f
C24668 DVDD.n7555 VSS 0.451316f
C24669 DVDD.n7556 VSS 0.451316f
C24670 DVDD.n7557 VSS 0.451316f
C24671 DVDD.n7558 VSS 0.451316f
C24672 DVDD.n7559 VSS 0.451316f
C24673 DVDD.n7560 VSS 0.451316f
C24674 DVDD.n7561 VSS 0.451316f
C24675 DVDD.n7562 VSS 0.451316f
C24676 DVDD.n7563 VSS 0.451316f
C24677 DVDD.n7564 VSS 0.451316f
C24678 DVDD.n7565 VSS 0.197054f
C24679 DVDD.n7566 VSS 0.066735f
C24680 DVDD.n7567 VSS 0.066735f
C24681 DVDD.n7568 VSS 0.066735f
C24682 DVDD.n7569 VSS 0.066735f
C24683 DVDD.n7570 VSS 0.066735f
C24684 DVDD.n7571 VSS 0.066735f
C24685 DVDD.n7572 VSS 0.066735f
C24686 DVDD.n7573 VSS 0.066735f
C24687 DVDD.n7574 VSS 0.066735f
C24688 DVDD.n7575 VSS 0.066735f
C24689 DVDD.n7576 VSS 0.197054f
C24690 DVDD.n7587 VSS 0.225658f
C24691 DVDD.n7589 VSS 0.066735f
C24692 DVDD.n7590 VSS 0.225658f
C24693 DVDD.n7591 VSS 0.127013f
C24694 DVDD.n7592 VSS 0.149379f
C24695 DVDD.n7593 VSS 0.726238f
C24696 DVDD.n7594 VSS 0.182751f
C24697 DVDD.n7595 VSS 0.301937f
C24698 DVDD.n7596 VSS 0.301937f
C24699 DVDD.n7597 VSS 0.861315f
C24700 DVDD.n7598 VSS 0.375037f
C24701 DVDD.n7599 VSS 0.451316f
C24702 DVDD.n7600 VSS 0.451316f
C24703 DVDD.n7601 VSS 0.451316f
C24704 DVDD.n7602 VSS 0.451316f
C24705 DVDD.n7603 VSS 0.451316f
C24706 DVDD.n7604 VSS 0.451316f
C24707 DVDD.n7605 VSS 0.451316f
C24708 DVDD.n7606 VSS 0.451316f
C24709 DVDD.n7607 VSS 0.451316f
C24710 DVDD.n7608 VSS 0.451316f
C24711 DVDD.n7609 VSS 0.451316f
C24712 DVDD.n7610 VSS 0.451316f
C24713 DVDD.n7611 VSS 0.451316f
C24714 DVDD.n7612 VSS 0.451316f
C24715 DVDD.n7613 VSS 0.451316f
C24716 DVDD.n7614 VSS 0.451316f
C24717 DVDD.n7615 VSS 0.451316f
C24718 DVDD.n7616 VSS 0.451316f
C24719 DVDD.n7617 VSS 0.451316f
C24720 DVDD.n7618 VSS 0.451316f
C24721 DVDD.n7619 VSS 0.451316f
C24722 DVDD.n7620 VSS 0.451316f
C24723 DVDD.n7621 VSS 0.451316f
C24724 DVDD.n7622 VSS 0.451316f
C24725 DVDD.n7623 VSS 0.451316f
C24726 DVDD.n7624 VSS 0.451316f
C24727 DVDD.n7625 VSS 0.451316f
C24728 DVDD.n7626 VSS 0.451316f
C24729 DVDD.n7627 VSS 0.451316f
C24730 DVDD.n7628 VSS 0.451316f
C24731 DVDD.n7629 VSS 0.451316f
C24732 DVDD.n7630 VSS 0.451316f
C24733 DVDD.n7631 VSS 0.451316f
C24734 DVDD.n7632 VSS 0.451316f
C24735 DVDD.n7633 VSS 0.289224f
C24736 DVDD.n7634 VSS 0.289224f
C24737 DVDD.n7635 VSS 0.451316f
C24738 DVDD.n7636 VSS 0.451316f
C24739 DVDD.n7637 VSS 0.451316f
C24740 DVDD.n7638 VSS 0.451316f
C24741 DVDD.n7639 VSS 0.451316f
C24742 DVDD.n7640 VSS 0.451316f
C24743 DVDD.n7641 VSS 0.451316f
C24744 DVDD.n7642 VSS 0.451316f
C24745 DVDD.n7643 VSS 0.451316f
C24746 DVDD.n7644 VSS 0.451316f
C24747 DVDD.n7645 VSS 0.451316f
C24748 DVDD.n7646 VSS 0.451316f
C24749 DVDD.n7647 VSS 0.451316f
C24750 DVDD.n7648 VSS 0.451316f
C24751 DVDD.n7649 VSS 0.451316f
C24752 DVDD.n7650 VSS 0.451316f
C24753 DVDD.n7651 VSS 0.451316f
C24754 DVDD.n7652 VSS 0.451316f
C24755 DVDD.n7653 VSS 0.197054f
C24756 DVDD.n7654 VSS 0.451316f
C24757 DVDD.n7655 VSS 0.451316f
C24758 DVDD.n7656 VSS 0.197054f
C24759 DVDD.n7660 VSS 0.225658f
C24760 DVDD.n7661 VSS 0.022884f
C24761 DVDD.n7662 VSS 0.022884f
C24762 DVDD.n7663 VSS 0.011442f
C24763 DVDD.n7664 VSS 0.036871f
C24764 DVDD.n7665 VSS 0.301841f
C24765 DVDD.n7666 VSS 0.220837f
C24766 DVDD.n7667 VSS 0.011442f
C24767 DVDD.n7668 VSS 0.022884f
C24768 DVDD.n7669 VSS 0.022884f
C24769 DVDD.n7670 VSS 0.011442f
C24770 DVDD.n7671 VSS 0.13031f
C24771 DVDD.t6 VSS 1.69508f
C24772 DVDD.n7672 VSS 0.13031f
C24773 DVDD.n7673 VSS 0.033368f
C24774 DVDD.n7674 VSS 0.011442f
C24775 DVDD.n7675 VSS 0.220876f
C24776 DVDD.n7676 VSS 0.301797f
C24777 DVDD.n7677 VSS 0.036905f
C24778 DVDD.n7678 VSS 0.029062f
C24779 DVDD.n7679 VSS 0.225658f
C24780 DVDD.n7680 VSS 0.063506f
C24781 DVDD.n7681 VSS 0.042106f
C24782 DVDD.n7682 VSS 0.042106f
C24783 DVDD.n7683 VSS 0.059201f
C24784 DVDD.n7684 VSS 0.379733f
C24785 DVDD.n7685 VSS 0.034444f
C24786 DVDD.n7686 VSS 0.672082f
C24787 DVDD.n7687 VSS 0.243708f
C24788 DVDD.n7689 VSS 0.672082f
C24789 DVDD.n7690 VSS 0.033368f
C24790 DVDD.n7693 VSS 0.042106f
C24791 DVDD.n7694 VSS 0.033368f
C24792 DVDD.n7695 VSS 0.379733f
C24793 DVDD.n7696 VSS 0.379733f
C24794 DVDD.n7697 VSS 0.033368f
C24795 DVDD.n7700 VSS 0.042106f
C24796 DVDD.n7701 VSS 0.033368f
C24797 DVDD.n7702 VSS 0.23977f
C24798 DVDD.n7703 VSS 0.033368f
C24799 DVDD.n7705 VSS 0.042106f
C24800 DVDD.n7706 VSS 0.042106f
C24801 DVDD.n7708 VSS 0.042106f
C24802 DVDD.n7710 VSS 0.033368f
C24803 DVDD.n7713 VSS 0.042106f
C24804 DVDD.n7714 VSS 0.042106f
C24805 DVDD.n7716 VSS 0.033368f
C24806 DVDD.n7718 VSS 0.042106f
C24807 DVDD.n7719 VSS 0.033368f
C24808 DVDD.n7720 VSS 0.379733f
C24809 DVDD.n7722 VSS 0.033368f
C24810 DVDD.n7723 VSS 0.379733f
C24811 DVDD.n7724 VSS 0.033368f
C24812 DVDD.n7725 VSS 0.23977f
C24813 DVDD.n7726 VSS -1.46111f
C24814 DVDD.n7727 VSS 2.21687f
C24815 DVDD.n7728 VSS 3.24347f
C24816 DVDD.n7729 VSS 0.243708f
C24817 DVDD.n7731 VSS 0.042106f
C24818 DVDD.n7732 VSS 0.042106f
C24819 DVDD.n7733 VSS 0.059201f
C24820 DVDD.n7734 VSS 0.672082f
C24821 DVDD.n7735 VSS 0.034444f
C24822 DVDD.n7736 VSS 0.379733f
C24823 DVDD.n7737 VSS 0.379733f
C24824 DVDD.n7738 VSS 0.042106f
C24825 DVDD.n7740 VSS 0.042106f
C24826 DVDD.n7742 VSS 0.058124f
C24827 DVDD.n7743 VSS 0.23977f
C24828 DVDD.n7745 VSS 0.059201f
C24829 DVDD.n7746 VSS 0.063506f
C24830 DVDD.n7747 VSS 0.225658f
C24831 DVDD.n7748 VSS 0.029062f
C24832 DVDD.n7749 VSS 0.225658f
C24833 DVDD.n7750 VSS 0.367092f
C24834 DVDD.n7751 VSS 0.451316f
C24835 DVDD.n7752 VSS 0.451316f
C24836 DVDD.n7753 VSS 0.451316f
C24837 DVDD.n7754 VSS 0.451316f
C24838 DVDD.n7755 VSS 0.451316f
C24839 DVDD.n7756 VSS 0.451316f
C24840 DVDD.n7757 VSS 0.451316f
C24841 DVDD.n7758 VSS 0.451316f
C24842 DVDD.n7759 VSS 0.451316f
C24843 DVDD.n7760 VSS 0.451316f
C24844 DVDD.n7761 VSS 0.451316f
C24845 DVDD.n7762 VSS 0.451316f
C24846 DVDD.n7763 VSS 0.451316f
C24847 DVDD.n7764 VSS 0.451316f
C24848 DVDD.n7765 VSS 0.451316f
C24849 DVDD.n7766 VSS 0.451316f
C24850 DVDD.n7767 VSS 0.451316f
C24851 DVDD.n7768 VSS 0.451316f
C24852 DVDD.n7769 VSS 0.451316f
C24853 DVDD.n7770 VSS 0.451316f
C24854 DVDD.n7771 VSS 0.451316f
C24855 DVDD.n7772 VSS 0.451316f
C24856 DVDD.n7773 VSS 0.360735f
C24857 DVDD.n7776 VSS 0.225658f
C24858 DVDD.n7777 VSS 0.056779f
C24859 DVDD.n7778 VSS 0.225658f
C24860 DVDD.n7779 VSS 0.127013f
C24861 DVDD.n7780 VSS 0.225658f
C24862 DVDD.n7781 VSS 0.197054f
C24863 DVDD.n7782 VSS 0.451316f
C24864 DVDD.n7783 VSS 0.387751f
C24865 DVDD.n7784 VSS 0.338487f
C24866 DVDD.n7785 VSS 0.861315f
C24867 DVDD.n7786 VSS 0.861315f
C24868 DVDD.n7787 VSS 0.289224f
C24869 DVDD.n7788 VSS 0.289224f
C24870 DVDD.n7789 VSS 0.289224f
C24871 DVDD.n7790 VSS 0.861315f
C24872 DVDD.n7791 VSS 0.387751f
C24873 DVDD.n7792 VSS 0.451316f
C24874 DVDD.n7793 VSS 0.451316f
C24875 DVDD.n7794 VSS 0.197054f
C24876 DVDD.n7795 VSS 0.066735f
C24877 DVDD.n7798 VSS 0.197054f
C24878 DVDD.n7799 VSS 0.225658f
C24879 DVDD.n7801 VSS 0.066735f
C24880 DVDD.n7802 VSS 0.066735f
C24881 DVDD.n7803 VSS 0.225658f
C24882 DVDD.n7804 VSS 0.066735f
C24883 DVDD.n7806 VSS 0.225658f
C24884 DVDD.n7807 VSS 0.197054f
C24885 DVDD.n7808 VSS 0.451316f
C24886 DVDD.n7809 VSS 0.451316f
C24887 DVDD.n7810 VSS 0.451316f
C24888 DVDD.n7811 VSS 0.451316f
C24889 DVDD.n7812 VSS 0.451316f
C24890 DVDD.n7813 VSS 0.451316f
C24891 DVDD.n7814 VSS 0.451316f
C24892 DVDD.n7815 VSS 0.451316f
C24893 DVDD.n7816 VSS 0.451316f
C24894 DVDD.n7817 VSS 0.451316f
C24895 DVDD.n7818 VSS 0.451316f
C24896 DVDD.n7819 VSS 0.451316f
C24897 DVDD.n7820 VSS 0.451316f
C24898 DVDD.n7821 VSS 0.451316f
C24899 DVDD.n7822 VSS 0.451316f
C24900 DVDD.n7823 VSS 0.451316f
C24901 DVDD.n7824 VSS 0.451316f
C24902 DVDD.n7825 VSS 0.451316f
C24903 DVDD.n7826 VSS 0.451316f
C24904 DVDD.n7827 VSS 0.451316f
C24905 DVDD.n7828 VSS 0.451316f
C24906 DVDD.n7829 VSS 0.451316f
C24907 DVDD.n7830 VSS 0.451316f
C24908 DVDD.n7831 VSS 0.451316f
C24909 DVDD.n7832 VSS 0.451316f
C24910 DVDD.n7833 VSS 0.451316f
C24911 DVDD.n7834 VSS 0.451316f
C24912 DVDD.n7835 VSS 0.451316f
C24913 DVDD.n7836 VSS 0.451316f
C24914 DVDD.n7837 VSS 0.451316f
C24915 DVDD.n7838 VSS 0.451316f
C24916 DVDD.n7842 VSS 0.225658f
C24917 DVDD.n7843 VSS 0.367092f
C24918 DVDD.n7844 VSS 0.451316f
C24919 DVDD.n7845 VSS 0.451316f
C24920 DVDD.n7846 VSS 0.451316f
C24921 DVDD.n7847 VSS 0.451316f
C24922 DVDD.n7848 VSS 0.451316f
C24923 DVDD.n7849 VSS 0.451316f
C24924 DVDD.n7850 VSS 0.197054f
C24925 DVDD.n7851 VSS 0.225658f
C24926 DVDD.n7852 VSS 0.03875f
C24927 DVDD.n7853 VSS 0.225658f
C24928 DVDD.n7854 VSS 0.220891f
C24929 DVDD.n7855 VSS 0.276511f
C24930 DVDD.n7856 VSS 0.861315f
C24931 DVDD.n7857 VSS 0.400464f
C24932 DVDD.n7858 VSS 0.400464f
C24933 DVDD.n7859 VSS 0.400464f
C24934 DVDD.n7860 VSS 0.451316f
C24935 DVDD.n7861 VSS 0.451316f
C24936 DVDD.n7862 VSS 0.451316f
C24937 DVDD.n7863 VSS 0.451316f
C24938 DVDD.n7864 VSS 0.451316f
C24939 DVDD.n7865 VSS 0.451316f
C24940 DVDD.n7866 VSS 0.451316f
C24941 DVDD.n7867 VSS 0.451316f
C24942 DVDD.n7868 VSS 0.451316f
C24943 DVDD.n7869 VSS 0.451316f
C24944 DVDD.n7870 VSS 0.451316f
C24945 DVDD.n7871 VSS 0.451316f
C24946 DVDD.n7872 VSS 0.451316f
C24947 DVDD.n7873 VSS 0.451316f
C24948 DVDD.n7874 VSS 0.451316f
C24949 DVDD.n7875 VSS 0.451316f
C24950 DVDD.n7876 VSS 0.451316f
C24951 DVDD.n7877 VSS 0.451316f
C24952 DVDD.n7878 VSS 0.451316f
C24953 DVDD.n7879 VSS 0.451316f
C24954 DVDD.n7880 VSS 0.451316f
C24955 DVDD.n7881 VSS 0.451316f
C24956 DVDD.n7882 VSS 0.451316f
C24957 DVDD.n7883 VSS 0.451316f
C24958 DVDD.n7884 VSS 0.451316f
C24959 DVDD.n7885 VSS 0.197054f
C24960 DVDD.n7886 VSS 0.225658f
C24961 DVDD.n7888 VSS 0.066735f
C24962 DVDD.n7889 VSS 0.066735f
C24963 DVDD.n7890 VSS 0.225658f
C24964 DVDD.n7891 VSS 0.066735f
C24965 DVDD.n7893 VSS 0.225658f
C24966 DVDD.n7894 VSS 0.395696f
C24967 DVDD.n7895 VSS 0.451316f
C24968 DVDD.n7896 VSS 0.451316f
C24969 DVDD.n7897 VSS 0.451316f
C24970 DVDD.n7898 VSS 0.451316f
C24971 DVDD.n7899 VSS 0.451316f
C24972 DVDD.n7900 VSS 0.451316f
C24973 DVDD.n7901 VSS 0.451316f
C24974 DVDD.n7902 VSS 0.451316f
C24975 DVDD.n7903 VSS 0.451316f
C24976 DVDD.n7904 VSS 0.451316f
C24977 DVDD.n7905 VSS 0.451316f
C24978 DVDD.n7906 VSS 0.451316f
C24979 DVDD.n7907 VSS 0.451316f
C24980 DVDD.n7908 VSS 0.451316f
C24981 DVDD.n7909 VSS 0.451316f
C24982 DVDD.n7910 VSS 0.263798f
C24983 DVDD.n7911 VSS 0.263798f
C24984 DVDD.n7912 VSS 0.263798f
C24985 DVDD.n7913 VSS 0.861315f
C24986 DVDD.n7914 VSS 0.413177f
C24987 DVDD.n7915 VSS 0.413177f
C24988 DVDD.n7926 VSS 0.225658f
C24989 DVDD.n7927 VSS 0.197054f
C24990 DVDD.n7928 VSS 0.451316f
C24991 DVDD.n7929 VSS 0.197054f
C24992 DVDD.n7930 VSS 0.451316f
C24993 DVDD.n7931 VSS 0.451316f
C24994 DVDD.n7932 VSS 0.451316f
C24995 DVDD.n7933 VSS 0.451316f
C24996 DVDD.n7934 VSS 0.451316f
C24997 DVDD.n7935 VSS 0.451316f
C24998 DVDD.n7936 VSS 0.451316f
C24999 DVDD.n7937 VSS 0.451316f
C25000 DVDD.n7938 VSS 0.451316f
C25001 DVDD.n7939 VSS 0.451316f
C25002 DVDD.n7940 VSS 0.451316f
C25003 DVDD.n7941 VSS 0.451316f
C25004 DVDD.n7942 VSS 0.451316f
C25005 DVDD.n7943 VSS 0.451316f
C25006 DVDD.n7944 VSS 0.451316f
C25007 DVDD.n7945 VSS 0.232015f
C25008 DVDD.n7946 VSS 2.07943f
C25009 DVDD.n7947 VSS 0.6412f
C25010 DVDD.n7948 VSS 0.197054f
C25011 DVDD.n7949 VSS 0.40682f
C25012 DVDD.n7950 VSS 0.451316f
C25013 DVDD.n7951 VSS 0.197054f
C25014 DVDD.n7954 VSS 0.225658f
C25015 DVDD.n7957 VSS 0.062794f
C25016 DVDD.n7958 VSS 0.225658f
C25017 DVDD.n7959 VSS 0.079457f
C25018 DVDD.n7960 VSS 0.079457f
C25019 DVDD.n7961 VSS 0.197054f
C25020 DVDD.n7962 VSS 0.062794f
C25021 DVDD.n7963 VSS 0.062794f
C25022 DVDD.n7964 VSS 0.062794f
C25023 DVDD.n7965 VSS 0.062794f
C25024 DVDD.n7966 VSS 0.062794f
C25025 DVDD.n7967 VSS 0.062794f
C25026 DVDD.n7968 VSS 0.062794f
C25027 DVDD.n7969 VSS 0.062794f
C25028 DVDD.n7970 VSS 0.062794f
C25029 DVDD.n7971 VSS 0.062794f
C25030 DVDD.n7972 VSS 0.062794f
C25031 DVDD.n7985 VSS 0.181162f
C25032 DVDD.n7997 VSS 0.225658f
C25033 DVDD.n7998 VSS 0.197054f
C25034 DVDD.n7999 VSS 0.451316f
C25035 DVDD.n8000 VSS 0.451316f
C25036 DVDD.n8001 VSS 0.451316f
C25037 DVDD.n8002 VSS 0.40682f
C25038 DVDD.n8003 VSS 0.050852f
C25039 DVDD.n8004 VSS 2.07943f
C25040 DVDD.n8005 VSS 0.6412f
C25041 DVDD.n8006 VSS 0.40682f
C25042 DVDD.n8007 VSS 0.197054f
C25043 DVDD.n8008 VSS 0.225658f
C25044 DVDD.n8009 VSS 0.079457f
C25045 DVDD.n8010 VSS 0.225658f
C25046 DVDD.n8011 VSS 0.367092f
C25047 DVDD.n8012 VSS 0.451316f
C25048 DVDD.n8013 VSS 0.451316f
C25049 DVDD.n8014 VSS 0.451316f
C25050 DVDD.n8015 VSS 0.451316f
C25051 DVDD.n8016 VSS 0.451316f
C25052 DVDD.n8017 VSS 0.395696f
C25053 DVDD.n8018 VSS 0.451316f
C25054 DVDD.n8019 VSS 0.197054f
C25055 DVDD.n8020 VSS 0.451316f
C25056 DVDD.n8031 VSS 0.225658f
C25057 DVDD.n8032 VSS 0.197054f
C25058 DVDD.n8033 VSS 0.451316f
C25059 DVDD.n8034 VSS 0.413177f
C25060 DVDD.n8035 VSS 0.861315f
C25061 DVDD.n8036 VSS 0.263798f
C25062 DVDD.n8037 VSS 0.263798f
C25063 DVDD.n8038 VSS 0.451316f
C25064 DVDD.n8039 VSS 0.451316f
C25065 DVDD.n8040 VSS 0.451316f
C25066 DVDD.n8041 VSS 0.451316f
C25067 DVDD.n8042 VSS 0.451316f
C25068 DVDD.n8043 VSS 0.451316f
C25069 DVDD.n8044 VSS 0.451316f
C25070 DVDD.n8045 VSS 0.451316f
C25071 DVDD.n8046 VSS 0.451316f
C25072 DVDD.n8047 VSS 0.451316f
C25073 DVDD.n8048 VSS 0.451316f
C25074 DVDD.n8049 VSS 0.395696f
C25075 DVDD.n8052 VSS 0.225658f
C25076 DVDD.n8053 VSS 0.056779f
C25077 DVDD.n8054 VSS 0.225658f
C25078 DVDD.n8055 VSS 0.127013f
C25079 DVDD.n8056 VSS 0.225658f
C25080 DVDD.n8057 VSS 0.197054f
C25081 DVDD.n8058 VSS 0.451316f
C25082 DVDD.n8059 VSS 0.451316f
C25083 DVDD.n8060 VSS 0.451316f
C25084 DVDD.n8061 VSS 0.451316f
C25085 DVDD.n8062 VSS 0.451316f
C25086 DVDD.n8063 VSS 0.451316f
C25087 DVDD.n8064 VSS 0.451316f
C25088 DVDD.n8065 VSS 0.451316f
C25089 DVDD.n8066 VSS 0.451316f
C25090 DVDD.n8067 VSS 0.451316f
C25091 DVDD.n8068 VSS 0.451316f
C25092 DVDD.n8069 VSS 0.451316f
C25093 DVDD.n8070 VSS 0.451316f
C25094 DVDD.n8071 VSS 0.451316f
C25095 DVDD.n8072 VSS 0.451316f
C25096 DVDD.n8073 VSS 0.451316f
C25097 DVDD.n8074 VSS 0.451316f
C25098 DVDD.n8075 VSS 0.400464f
C25099 DVDD.n8076 VSS 0.400464f
C25100 DVDD.n8077 VSS 0.400464f
C25101 DVDD.n8078 VSS 0.861315f
C25102 DVDD.n8079 VSS 0.543486f
C25103 DVDD.n8080 VSS 0.400464f
C25104 DVDD.n8081 VSS 0.400464f
C25105 DVDD.n8082 VSS 0.400464f
C25106 DVDD.n8083 VSS 0.451316f
C25107 DVDD.n8084 VSS 0.451316f
C25108 DVDD.n8085 VSS 0.451316f
C25109 DVDD.n8086 VSS 0.451316f
C25110 DVDD.n8087 VSS 0.451316f
C25111 DVDD.n8088 VSS 0.451316f
C25112 DVDD.n8089 VSS 0.451316f
C25113 DVDD.n8090 VSS 0.451316f
C25114 DVDD.n8091 VSS 0.451316f
C25115 DVDD.n8092 VSS 0.451316f
C25116 DVDD.n8093 VSS 0.451316f
C25117 DVDD.n8094 VSS 0.451316f
C25118 DVDD.n8095 VSS 0.451316f
C25119 DVDD.n8096 VSS 0.451316f
C25120 DVDD.n8097 VSS 0.451316f
C25121 DVDD.n8098 VSS 0.451316f
C25122 DVDD.n8099 VSS 0.451316f
C25123 DVDD.n8100 VSS 0.451316f
C25124 DVDD.n8101 VSS 0.451316f
C25125 DVDD.n8102 VSS 0.451316f
C25126 DVDD.n8103 VSS 0.451316f
C25127 DVDD.n8104 VSS 0.451316f
C25128 DVDD.n8105 VSS 0.451316f
C25129 DVDD.n8106 VSS 0.451316f
C25130 DVDD.n8107 VSS 0.451316f
C25131 DVDD.n8108 VSS 0.197054f
C25132 DVDD.n8115 VSS 0.225658f
C25133 DVDD.n8117 VSS 0.066735f
C25134 DVDD.n8118 VSS 0.225658f
C25135 DVDD.n8119 VSS 0.559179f
C25136 DVDD.n8120 VSS 0.225658f
C25137 DVDD.n8121 VSS 0.395696f
C25138 DVDD.n8122 VSS 0.451316f
C25139 DVDD.n8123 VSS 0.451316f
C25140 DVDD.n8124 VSS 0.451316f
C25141 DVDD.n8125 VSS 0.451316f
C25142 DVDD.n8126 VSS 0.451316f
C25143 DVDD.n8127 VSS 0.451316f
C25144 DVDD.n8128 VSS 0.451316f
C25145 DVDD.n8129 VSS 0.451316f
C25146 DVDD.n8130 VSS 0.451316f
C25147 DVDD.n8131 VSS 0.451316f
C25148 DVDD.n8132 VSS 0.451316f
C25149 DVDD.n8133 VSS 0.451316f
C25150 DVDD.n8134 VSS 0.451316f
C25151 DVDD.n8135 VSS 0.451316f
C25152 DVDD.n8136 VSS 0.451316f
C25153 DVDD.n8137 VSS 0.263798f
C25154 DVDD.n8138 VSS 0.263798f
C25155 DVDD.n8139 VSS 0.263798f
C25156 DVDD.n8140 VSS 0.543486f
C25157 DVDD.n8141 VSS 0.413177f
C25158 DVDD.n8142 VSS 0.413177f
C25159 DVDD.n8151 VSS 0.225658f
C25160 DVDD.n8152 VSS 0.197054f
C25161 DVDD.n8153 VSS 0.451316f
C25162 DVDD.n8154 VSS 0.197054f
C25163 DVDD.n8155 VSS 0.451316f
C25164 DVDD.n8156 VSS 0.451316f
C25165 DVDD.n8157 VSS 0.451316f
C25166 DVDD.n8158 VSS 0.451316f
C25167 DVDD.n8159 VSS 0.451316f
C25168 DVDD.n8160 VSS 0.451316f
C25169 DVDD.n8161 VSS 0.451316f
C25170 DVDD.n8162 VSS 0.451316f
C25171 DVDD.n8163 VSS 0.451316f
C25172 DVDD.n8164 VSS 0.451316f
C25173 DVDD.n8165 VSS 0.451316f
C25174 DVDD.n8166 VSS 0.451316f
C25175 DVDD.n8167 VSS 0.451316f
C25176 DVDD.n8168 VSS 0.451316f
C25177 DVDD.n8169 VSS 0.40682f
C25178 DVDD.n8170 VSS 0.050852f
C25179 DVDD.n8171 VSS 2.07943f
C25180 DVDD.n8172 VSS 0.6412f
C25181 DVDD.n8173 VSS 0.197054f
C25182 DVDD.n8174 VSS 0.40682f
C25183 DVDD.n8175 VSS 0.451316f
C25184 DVDD.n8176 VSS 0.197054f
C25185 DVDD.n8187 VSS 0.225658f
C25186 DVDD.n8190 VSS 0.062794f
C25187 DVDD.n8191 VSS 0.225658f
C25188 DVDD.n8192 VSS 0.249601f
C25189 DVDD.n8193 VSS 0.249601f
C25190 DVDD.n8194 VSS 0.062794f
C25191 DVDD.n8195 VSS 0.062794f
C25192 DVDD.n8196 VSS 0.062794f
C25193 DVDD.n8200 VSS 0.189849f
C25194 DVDD.n8201 VSS 0.189849f
C25195 DVDD.n8202 VSS 0.023731f
C25196 DVDD.n8203 VSS 0.277232f
C25197 DVDD.n8204 VSS 1.01509f
C25198 DVDD.n8205 VSS 0.084542f
C25199 DVDD.n8207 VSS 0.062794f
C25200 DVDD.n8208 VSS 0.105307f
C25201 DVDD.n8209 VSS -2.07648f
C25202 DVDD.n8210 VSS 0.105307f
C25203 DVDD.n8211 VSS 0.091958f
C25204 DVDD.n8212 VSS 0.210614f
C25205 DVDD.n8213 VSS 0.210614f
C25206 DVDD.n8214 VSS 0.210614f
C25207 DVDD.n8215 VSS 0.210614f
C25208 DVDD.n8216 VSS 0.210614f
C25209 DVDD.n8217 VSS 0.210614f
C25210 DVDD.n8218 VSS 0.210614f
C25211 DVDD.n8219 VSS 0.210614f
C25212 DVDD.n8220 VSS 0.210614f
C25213 DVDD.n8221 VSS 0.210614f
C25214 DVDD.n8222 VSS 0.210614f
C25215 DVDD.n8223 VSS 0.210614f
C25216 DVDD.n8224 VSS 0.091958f
C25217 DVDD.n8225 VSS 0.210614f
C25218 DVDD.n8226 VSS 0.091958f
C25219 DVDD.n8227 VSS 0.210614f
C25220 DVDD.n8228 VSS 0.210614f
C25221 DVDD.n8229 VSS 0.210614f
C25222 DVDD.n8230 VSS 0.210614f
C25223 DVDD.n8231 VSS 0.210614f
C25224 DVDD.n8232 VSS 0.210614f
C25225 DVDD.n8233 VSS 0.210614f
C25226 DVDD.n8234 VSS 0.210614f
C25227 DVDD.n8235 VSS 0.210614f
C25228 DVDD.n8236 VSS 0.210614f
C25229 DVDD.n8237 VSS 0.210614f
C25230 DVDD.n8238 VSS 0.210614f
C25231 DVDD.n8239 VSS 0.210614f
C25232 DVDD.n8240 VSS 0.210614f
C25233 DVDD.n8241 VSS 0.210614f
C25234 DVDD.n8242 VSS 0.210614f
C25235 DVDD.n8243 VSS 0.210614f
C25236 DVDD.n8244 VSS 0.210614f
C25237 DVDD.n8245 VSS 0.210614f
C25238 DVDD.n8246 VSS 0.210614f
C25239 DVDD.n8247 VSS 0.210614f
C25240 DVDD.n8248 VSS 0.210614f
C25241 DVDD.n8249 VSS 0.091958f
C25242 DVDD.n8250 VSS 0.105307f
C25243 DVDD.n8251 VSS 0.066735f
C25244 DVDD.n8252 VSS 0.105307f
C25245 DVDD.n8253 VSS 0.171309f
C25246 DVDD.n8254 VSS 0.210614f
C25247 DVDD.n8255 VSS 0.210614f
C25248 DVDD.n8256 VSS 0.210614f
C25249 DVDD.n8257 VSS 0.210614f
C25250 DVDD.n8258 VSS 0.210614f
C25251 DVDD.n8259 VSS 0.210614f
C25252 DVDD.n8260 VSS 0.210614f
C25253 DVDD.n8261 VSS 0.210614f
C25254 DVDD.n8262 VSS 0.210614f
C25255 DVDD.n8263 VSS 0.210614f
C25256 DVDD.n8264 VSS 0.210614f
C25257 DVDD.n8265 VSS 0.210614f
C25258 DVDD.n8266 VSS 0.210614f
C25259 DVDD.n8267 VSS 0.210614f
C25260 DVDD.n8268 VSS 0.210614f
C25261 DVDD.n8269 VSS 0.210614f
C25262 DVDD.n8270 VSS 0.210614f
C25263 DVDD.n8271 VSS 0.210614f
C25264 DVDD.n8272 VSS 0.210614f
C25265 DVDD.n8273 VSS 0.210614f
C25266 DVDD.n8274 VSS 0.210614f
C25267 DVDD.n8275 VSS 0.210614f
C25268 DVDD.n8276 VSS 0.210614f
C25269 DVDD.n8277 VSS 0.184658f
C25270 DVDD.n8278 VSS 0.210614f
C25271 DVDD.n8279 VSS 0.210614f
C25272 DVDD.n8280 VSS 0.210614f
C25273 DVDD.n8281 VSS 0.210614f
C25274 DVDD.n8282 VSS 0.210614f
C25275 DVDD.n8283 VSS 0.091958f
C25276 DVDD.n8284 VSS 0.105307f
C25277 DVDD.n8286 VSS 0.066735f
C25278 DVDD.n8287 VSS 0.105307f
C25279 DVDD.n8288 VSS 0.559179f
C25280 DVDD.n8289 VSS 0.559179f
C25281 DVDD.n8290 VSS 0.225658f
C25282 DVDD.n8291 VSS 0.029062f
C25283 DVDD.n8292 VSS 0.225658f
C25284 DVDD.n8293 VSS 0.197054f
C25285 DVDD.n8294 VSS 0.451316f
C25286 DVDD.n8295 VSS 0.451316f
C25287 DVDD.n8296 VSS 0.451316f
C25288 DVDD.n8297 VSS 0.451316f
C25289 DVDD.n8298 VSS 0.451316f
C25290 DVDD.n8299 VSS 0.451316f
C25291 DVDD.n8300 VSS 0.451316f
C25292 DVDD.n8301 VSS 0.451316f
C25293 DVDD.n8302 VSS 0.451316f
C25294 DVDD.n8303 VSS 0.451316f
C25295 DVDD.n8304 VSS 0.451316f
C25296 DVDD.n8305 VSS 0.451316f
C25297 DVDD.n8306 VSS 0.451316f
C25298 DVDD.n8307 VSS 0.451316f
C25299 DVDD.n8308 VSS 0.451316f
C25300 DVDD.n8309 VSS 0.451316f
C25301 DVDD.n8310 VSS 0.451316f
C25302 DVDD.n8311 VSS 0.451316f
C25303 DVDD.n8312 VSS 0.451316f
C25304 DVDD.n8313 VSS 0.451316f
C25305 DVDD.n8314 VSS 0.451316f
C25306 DVDD.n8315 VSS 0.451316f
C25307 DVDD.n8316 VSS 0.451316f
C25308 DVDD.n8317 VSS 0.360735f
C25309 DVDD.n8318 VSS 0.451316f
C25310 DVDD.n8319 VSS 0.451316f
C25311 DVDD.n8320 VSS 0.197054f
C25312 DVDD.n8321 VSS 0.225658f
C25313 DVDD.n8322 VSS 0.559179f
C25314 DVDD.n8323 VSS 0.225658f
C25315 DVDD.n8324 VSS 0.338487f
C25316 DVDD.n8325 VSS 0.387751f
C25317 DVDD.n8326 VSS 0.543486f
C25318 DVDD.n8327 VSS 0.289224f
C25319 DVDD.n8328 VSS 0.451316f
C25320 DVDD.n8329 VSS 0.451316f
C25321 DVDD.n8330 VSS 0.451316f
C25322 DVDD.n8331 VSS 0.451316f
C25323 DVDD.n8332 VSS 0.451316f
C25324 DVDD.n8333 VSS 0.451316f
C25325 DVDD.n8334 VSS 0.451316f
C25326 DVDD.n8335 VSS 0.451316f
C25327 DVDD.n8336 VSS 0.451316f
C25328 DVDD.n8337 VSS 0.451316f
C25329 DVDD.n8338 VSS 0.451316f
C25330 DVDD.n8339 VSS 0.451316f
C25331 DVDD.n8340 VSS 0.451316f
C25332 DVDD.n8341 VSS 0.451316f
C25333 DVDD.n8342 VSS 0.451316f
C25334 DVDD.n8343 VSS 0.360735f
C25335 DVDD.n8344 VSS 0.451316f
C25336 DVDD.n8345 VSS 0.197054f
C25337 DVDD.n8346 VSS 0.451316f
C25338 DVDD.n8347 VSS 0.451316f
C25339 DVDD.n8348 VSS 0.197054f
C25340 DVDD.n8356 VSS 0.225658f
C25341 DVDD.n8357 VSS 0.029062f
C25342 DVDD.n8358 VSS 0.225658f
C25343 DVDD.n8359 VSS 0.559179f
C25344 DVDD.n8360 VSS 0.559179f
C25345 DVDD.n8361 VSS 0.066735f
C25346 DVDD.n8365 VSS 0.105307f
C25347 DVDD.n8368 VSS 0.066735f
C25348 DVDD.n8369 VSS 0.105307f
C25349 DVDD.n8370 VSS 0.638831f
C25350 DVDD.n8371 VSS 0.638831f
C25351 DVDD.n8372 VSS 0.066735f
C25352 DVDD.n8374 VSS 0.061481f
C25353 DVDD.n8376 VSS 0.501762f
C25354 DVDD.n8377 VSS 0.352514f
C25355 DVDD.n8378 VSS 0.360951f
C25356 DVDD.n8379 VSS 0.360951f
C25357 DVDD.n8380 VSS 0.061481f
C25358 DVDD.n8382 VSS 0.066735f
C25359 DVDD.n8383 VSS 0.061481f
C25360 DVDD.n8385 VSS 0.970017f
C25361 DVDD.n8386 VSS 0.360856f
C25362 DVDD.n8387 VSS 0.35655f
C25363 DVDD.n8388 VSS 0.176277f
C25364 DVDD.n8389 VSS 0.043231f
C25365 DVDD.n8390 VSS 0.022343f
C25366 DVDD.n8391 VSS 0.058124f
C25367 DVDD.n8392 VSS 0.058124f
C25368 DVDD.n8393 VSS 0.058124f
C25369 DVDD.n8394 VSS 0.025401f
C25370 DVDD.n8395 VSS 0.025401f
C25371 DVDD.n8396 VSS 0.025401f
C25372 DVDD.n8397 VSS 0.058124f
C25373 DVDD.n8398 VSS 0.058124f
C25374 DVDD.n8399 VSS 0.058124f
C25375 DVDD.n8400 VSS 0.025401f
C25376 DVDD.n8401 VSS 0.025401f
C25377 DVDD.n8402 VSS 0.022343f
C25378 DVDD.n8403 VSS 0.058124f
C25379 DVDD.n8404 VSS 0.058124f
C25380 DVDD.n8405 VSS 0.029062f
C25381 DVDD.n8406 VSS 0.035652f
C25382 DVDD.n8407 VSS 0.029062f
C25383 DVDD.n8408 VSS 0.058124f
C25384 DVDD.n8409 VSS 0.058124f
C25385 DVDD.n8410 VSS 0.025401f
C25386 DVDD.n8411 VSS 0.025401f
C25387 DVDD.n8412 VSS 0.022343f
C25388 DVDD.n8413 VSS 0.058124f
C25389 DVDD.n8414 VSS 0.058124f
C25390 DVDD.n8415 VSS 0.298559f
C25391 DVDD.n8416 VSS 0.307124f
C25392 DVDD.n8417 VSS 0.348747f
C25393 DVDD.n8418 VSS 0.043021f
C25394 DVDD.n8419 VSS 0.342557f
C25395 DVDD.n8420 VSS 0.387988f
C25396 DVDD.n8421 VSS 0.387988f
C25397 DVDD.n8424 VSS 0.043021f
C25398 DVDD.n8425 VSS 0.043021f
C25399 DVDD.n8426 VSS 0.043021f
C25400 DVDD.n8427 VSS 0.342557f
C25401 DVDD.n8428 VSS 0.244982f
C25402 DVDD.n8429 VSS 2.2453f
C25403 DVDD.n8430 VSS 0.446943f
C25404 DVDD.n8431 VSS 0.043021f
C25405 DVDD.n8433 VSS 0.244982f
C25406 DVDD.n8434 VSS 0.058124f
C25407 DVDD.n8435 VSS 0.387988f
C25408 DVDD.n8436 VSS 0.043021f
C25409 DVDD.n8438 VSS 0.387988f
C25410 DVDD.n8439 VSS 0.058124f
C25411 DVDD.n8440 VSS 0.307124f
C25412 DVDD.n8441 VSS 0.298559f
C25413 DVDD.n8442 VSS 0.029062f
C25414 DVDD.n8443 VSS 0.058124f
C25415 DVDD.n8444 VSS 0.058124f
C25416 DVDD.n8445 VSS 0.058124f
C25417 DVDD.n8446 VSS 0.022343f
C25418 DVDD.n8448 VSS 0.022343f
C25419 DVDD.n8449 VSS 0.35655f
C25420 DVDD.n8450 VSS 0.02105f
C25421 DVDD.n8451 VSS 0.058124f
C25422 DVDD.n8452 VSS 0.058124f
C25423 DVDD.n8453 VSS 0.058124f
C25424 DVDD.n8454 VSS 0.025401f
C25425 DVDD.n8455 VSS 0.025401f
C25426 DVDD.n8456 VSS 0.025401f
C25427 DVDD.n8457 VSS 0.058124f
C25428 DVDD.n8458 VSS 0.058124f
C25429 DVDD.n8459 VSS 0.058124f
C25430 DVDD.n8460 VSS 0.025401f
C25431 DVDD.n8461 VSS 0.025401f
C25432 DVDD.n8462 VSS 0.025401f
C25433 DVDD.n8463 VSS 0.058124f
C25434 DVDD.n8464 VSS 0.058124f
C25435 DVDD.n8465 VSS 0.029062f
C25436 DVDD.n8466 VSS 0.058124f
C25437 DVDD.n8467 VSS 0.035652f
C25438 DVDD.n8468 VSS 0.040796f
C25439 DVDD.n8469 VSS 0.022343f
C25440 DVDD.n8470 VSS 0.058124f
C25441 DVDD.n8471 VSS 0.058124f
C25442 DVDD.n8472 VSS 0.058124f
C25443 DVDD.n8473 VSS 0.025401f
C25444 DVDD.n8474 VSS 0.025401f
C25445 DVDD.n8475 VSS 0.025401f
C25446 DVDD.n8476 VSS 0.058124f
C25447 DVDD.n8477 VSS 0.058124f
C25448 DVDD.n8478 VSS 0.058124f
C25449 DVDD.n8479 VSS 0.025401f
C25450 DVDD.n8480 VSS 0.025401f
C25451 DVDD.n8481 VSS 0.022343f
C25452 DVDD.n8482 VSS 0.058124f
C25453 DVDD.n8483 VSS 0.058124f
C25454 DVDD.n8484 VSS 0.058124f
C25455 DVDD.n8485 VSS 0.025401f
C25456 DVDD.n8486 VSS 0.025401f
C25457 DVDD.n8487 VSS 0.022343f
C25458 DVDD.n8488 VSS 0.058124f
C25459 DVDD.n8489 VSS 0.058124f
C25460 DVDD.n8490 VSS 0.034259f
C25461 DVDD.n8491 VSS 0.058124f
C25462 DVDD.n8492 VSS 0.029062f
C25463 DVDD.n8493 VSS 0.298559f
C25464 DVDD.n8494 VSS 0.307124f
C25465 DVDD.n8495 VSS 0.348747f
C25466 DVDD.n8497 VSS 0.387988f
C25467 DVDD.n8498 VSS 0.387988f
C25468 DVDD.n8499 VSS 0.348747f
C25469 DVDD.n8501 VSS 0.244982f
C25470 DVDD.n8502 VSS 2.2453f
C25471 DVDD.n8503 VSS 0.446943f
C25472 DVDD.n8504 VSS 0.244982f
C25473 DVDD.n8505 VSS 0.348747f
C25474 DVDD.n8507 VSS 0.387988f
C25475 DVDD.n8508 VSS 0.348747f
C25476 DVDD.n8509 VSS 0.043021f
C25477 DVDD.n8511 VSS 0.348747f
C25478 DVDD.n8513 VSS 0.387988f
C25479 DVDD.n8514 VSS 0.342557f
C25480 DVDD.n8515 VSS 0.025401f
C25481 DVDD.n8516 VSS 0.342557f
C25482 DVDD.n8517 VSS 0.0127f
C25483 DVDD.n8519 VSS 0.0127f
C25484 DVDD.n8520 VSS 0.025401f
C25485 DVDD.n8521 VSS 0.025401f
C25486 DVDD.n8522 VSS 0.405257f
C25487 DVDD.n8523 VSS 0.063648f
C25488 DVDD.n8524 VSS 0.058124f
C25489 DVDD.n8525 VSS 0.022343f
C25490 DVDD.n8526 VSS 0.058124f
C25491 DVDD.n8527 VSS 0.025401f
C25492 DVDD.n8528 VSS 0.025401f
C25493 DVDD.n8529 VSS 0.025401f
C25494 DVDD.n8530 VSS 0.689855f
C25495 DVDD.n8531 VSS 0.374234f
C25496 DVDD.n8532 VSS 0.226026f
C25497 DVDD.n8534 VSS 0.025401f
C25498 DVDD.n8535 VSS 0.025401f
C25499 DVDD.n8536 VSS 0.0127f
C25500 DVDD.n8537 VSS 0.0127f
C25501 DVDD.n8538 VSS 0.229078f
C25502 DVDD.n8539 VSS 0.229078f
C25503 DVDD.n8540 VSS 0.405257f
C25504 DVDD.n8541 VSS 0.144644f
C25505 DVDD.n8542 VSS 0.263887f
C25506 DVDD.n8543 VSS 0.144644f
C25507 DVDD.n8544 VSS 0.405257f
C25508 DVDD.n8545 VSS 0.229078f
C25509 DVDD.n8546 VSS 0.229078f
C25510 DVDD.n8547 VSS 0.405257f
C25511 DVDD.n8548 VSS 0.226029f
C25512 DVDD.n8549 VSS 0.374234f
C25513 DVDD.n8550 VSS 0.689855f
C25514 DVDD.n8551 VSS 0.025401f
C25515 DVDD.n8552 VSS 0.025401f
C25516 DVDD.n8553 VSS 0.025401f
C25517 DVDD.n8554 VSS 0.058124f
C25518 DVDD.n8555 VSS 0.058124f
C25519 DVDD.n8556 VSS 0.058124f
C25520 DVDD.n8557 VSS 0.298559f
C25521 DVDD.n8558 VSS 0.040796f
C25522 DVDD.n8559 VSS 0.022343f
C25523 DVDD.n8560 VSS 0.058124f
C25524 DVDD.n8561 VSS 0.058124f
C25525 DVDD.n8562 VSS 0.058124f
C25526 DVDD.n8563 VSS 0.025401f
C25527 DVDD.n8564 VSS 0.025401f
C25528 DVDD.n8565 VSS 0.025401f
C25529 DVDD.n8566 VSS 0.058124f
C25530 DVDD.n8567 VSS 0.058124f
C25531 DVDD.n8568 VSS 0.058124f
C25532 DVDD.n8569 VSS 0.025401f
C25533 DVDD.n8570 VSS 0.025401f
C25534 DVDD.n8571 VSS 0.022343f
C25535 DVDD.n8572 VSS 0.058124f
C25536 DVDD.n8573 VSS 0.058124f
C25537 DVDD.n8574 VSS 0.029062f
C25538 DVDD.n8575 VSS 0.058124f
C25539 DVDD.n8576 VSS 0.029062f
C25540 DVDD.n8577 VSS 0.058124f
C25541 DVDD.n8578 VSS 0.058124f
C25542 DVDD.n8579 VSS 0.022343f
C25543 DVDD.n8580 VSS 0.025401f
C25544 DVDD.n8581 VSS 0.025401f
C25545 DVDD.n8582 VSS 0.058124f
C25546 DVDD.n8583 VSS 0.058124f
C25547 DVDD.n8584 VSS 0.058124f
C25548 DVDD.n8585 VSS 0.025401f
C25549 DVDD.n8586 VSS 0.130026f
C25550 DVDD.n8587 VSS 16.8082f
C25551 DVDD.n8588 VSS 0.847098f
C25552 DVDD.n8589 VSS 1.30412f
C25553 DVDD.n8590 VSS 2.2453f
C25554 DVDD.n8591 VSS 0.446943f
C25555 DVDD.n8592 VSS 0.244982f
C25556 DVDD.n8593 VSS 0.342557f
C25557 DVDD.n8594 VSS 0.043021f
C25558 DVDD.n8595 VSS 0.348747f
C25559 DVDD.n8596 VSS 0.387988f
C25560 DVDD.n8597 VSS 0.387988f
C25561 DVDD.n8598 VSS 0.342557f
C25562 DVDD.n8599 VSS 0.043021f
C25563 DVDD.n8600 VSS 0.348747f
C25564 DVDD.n8601 VSS 0.307124f
C25565 DVDD.n8602 VSS 0.298559f
C25566 DVDD.n8603 VSS 0.029062f
C25567 DVDD.n8604 VSS 0.058124f
C25568 DVDD.n8605 VSS 0.035652f
C25569 DVDD.n8606 VSS 0.058124f
C25570 DVDD.n8607 VSS 0.058124f
C25571 DVDD.n8608 VSS 0.022343f
C25572 DVDD.n8609 VSS 0.025401f
C25573 DVDD.n8610 VSS 0.025401f
C25574 DVDD.n8611 VSS 0.058124f
C25575 DVDD.n8612 VSS 0.058124f
C25576 DVDD.n8613 VSS 0.058124f
C25577 DVDD.n8614 VSS 0.025401f
C25578 DVDD.n8615 VSS 0.130026f
C25579 DVDD.n8616 VSS 16.8082f
C25580 DVDD.n8617 VSS 0.847098f
C25581 DVDD.n8618 VSS 1.51198f
C25582 DVDD.n8619 VSS 0.263887f
C25583 DVDD.n8620 VSS 0.0127f
C25584 DVDD.n8621 VSS 0.144644f
C25585 DVDD.n8622 VSS 0.342557f
C25586 DVDD.n8623 VSS 0.229078f
C25587 DVDD.n8624 VSS 0.229078f
C25588 DVDD.n8625 VSS 0.342557f
C25589 DVDD.n8626 VSS 0.181334f
C25590 DVDD.n8627 VSS 0.348208f
C25591 DVDD.n8628 VSS 0.352514f
C25592 DVDD.n8630 VSS 0.066735f
C25593 DVDD.n8631 VSS 0.360951f
C25594 DVDD.n8632 VSS 0.638831f
C25595 DVDD.n8633 VSS 0.501762f
C25596 DVDD.n8635 VSS 0.066735f
C25597 DVDD.n8636 VSS 0.501762f
C25598 DVDD.n8637 VSS 0.638831f
C25599 DVDD.n8638 VSS 0.316328f
C25600 DVDD.n8639 VSS -2.30734f
C25601 DVDD.n8640 VSS 3.37246f
C25602 DVDD.n8641 VSS 4.58897f
C25603 DVDD.n8642 VSS -0.119061f
C25604 DVDD.n8644 VSS 0.066735f
C25605 DVDD.n8645 VSS 0.970017f
C25606 DVDD.n8646 VSS 0.638831f
C25607 DVDD.n8647 VSS 0.638831f
C25608 DVDD.n8648 VSS 0.105307f
C25609 DVDD.n8649 VSS 0.559179f
C25610 DVDD.n8650 VSS 0.559179f
C25611 DVDD.n8651 VSS 0.187519f
C25612 DVDD.n8652 VSS 0.127013f
C25613 DVDD.n8653 VSS 0.127013f
C25614 DVDD.n8654 VSS 0.187519f
C25615 DVDD.n8655 VSS 0.127013f
C25616 DVDD.n8656 VSS 0.127013f
C25617 DVDD.n8657 VSS 0.187519f
C25618 DVDD.n8658 VSS 0.127013f
C25619 DVDD.n8659 VSS 0.127013f
C25620 DVDD.n8660 VSS 0.187519f
C25621 DVDD.n8661 VSS 0.559179f
C25622 DVDD.n8662 VSS 0.559179f
C25623 DVDD.n8663 VSS 0.10001f
C25624 DVDD.n8664 VSS 0.128627f
C25625 DVDD.n8665 VSS 0.128627f
C25626 DVDD.n8666 VSS 0.187519f
C25627 DVDD.n8667 VSS 1.85083f
C25628 DVDD.n8668 VSS 1.85083f
C25629 DVDD.n8669 VSS 0.066735f
C25630 DVDD.n8670 VSS 0.201821f
C25631 DVDD.n8671 VSS 0.029062f
C25632 DVDD.n8672 VSS 0.02691f
C25633 DVDD.n8673 VSS 0.026274f
C25634 DVDD.n8674 VSS 0.060175f
C25635 DVDD.n8675 VSS 0.061117f
C25636 DVDD.n8676 VSS 0.173937f
C25637 DVDD.n8677 VSS 0.060175f
C25638 DVDD.n8678 VSS 0.060175f
C25639 DVDD.n8679 VSS 0.026274f
C25640 DVDD.n8680 VSS 0.030088f
C25641 DVDD.n8681 VSS 0.029062f
C25642 DVDD.n8682 VSS 0.225658f
C25643 DVDD.n8683 VSS 0.066735f
C25644 DVDD.n8684 VSS 0.066735f
C25645 DVDD.n8685 VSS 0.066735f
C25646 DVDD.n8686 VSS 0.225658f
C25647 DVDD.n8687 VSS 0.04763f
C25648 DVDD.n8688 VSS 0.030088f
C25649 DVDD.n8689 VSS 0.026274f
C25650 DVDD.n8690 VSS 0.060175f
C25651 DVDD.n8691 VSS 0.059611f
C25652 DVDD.n8692 VSS 0.057655f
C25653 DVDD.n8693 VSS 0.060175f
C25654 DVDD.n8694 VSS 0.170687f
C25655 DVDD.n8695 VSS 0.060175f
C25656 DVDD.n8696 VSS 0.026274f
C25657 DVDD.n8697 VSS 0.029028f
C25658 DVDD.n8698 VSS 0.027333f
C25659 DVDD.n8699 VSS 0.066735f
C25660 DVDD.n8700 VSS 0.204999f
C25661 DVDD.n8701 VSS 0.026274f
C25662 DVDD.n8702 VSS 0.04884f
C25663 DVDD.n8703 VSS 0.225658f
C25664 DVDD.n8704 VSS 0.130242f
C25665 DVDD.n8705 VSS 0.130242f
C25666 DVDD.n8706 VSS 0.225658f
C25667 DVDD.n8707 VSS 0.10091f
C25668 DVDD.n8708 VSS 0.059656f
C25669 DVDD.n8709 VSS 0.057608f
C25670 DVDD.n8710 VSS 0.170688f
C25671 DVDD.n8711 VSS 0.060175f
C25672 DVDD.n8712 VSS 0.026274f
C25673 DVDD.n8713 VSS 0.030088f
C25674 DVDD.n8714 VSS 0.029062f
C25675 DVDD.n8715 VSS 0.225658f
C25676 DVDD.n8716 VSS 0.066735f
C25677 DVDD.n8717 VSS 0.066735f
C25678 DVDD.n8718 VSS 0.225658f
C25679 DVDD.n8719 VSS 0.029062f
C25680 DVDD.n8720 VSS 0.033368f
C25681 DVDD.n8721 VSS 0.114418f
C25682 DVDD.n8722 VSS 0.114418f
C25683 DVDD.n8723 VSS 0.033368f
C25684 DVDD.n8724 VSS 0.060175f
C25685 DVDD.n8725 VSS 0.030088f
C25686 DVDD.n8726 VSS 0.026274f
C25687 DVDD.n8727 VSS 0.060175f
C25688 DVDD.n8728 VSS 0.044284f
C25689 DVDD.n8729 VSS 0.173937f
C25690 DVDD.n8730 VSS 0.060175f
C25691 DVDD.n8731 VSS 0.060175f
C25692 DVDD.n8732 VSS 0.026274f
C25693 DVDD.n8733 VSS 0.030088f
C25694 DVDD.n8734 VSS 0.029062f
C25695 DVDD.n8735 VSS 0.225658f
C25696 DVDD.n8736 VSS 0.066735f
C25697 DVDD.n8737 VSS 0.066735f
C25698 DVDD.n8738 VSS 0.225658f
C25699 DVDD.n8739 VSS 0.029062f
C25700 DVDD.n8740 VSS 0.032022f
C25701 DVDD.n8741 VSS 0.030408f
C25702 DVDD.n8742 VSS 0.114418f
C25703 DVDD.n8743 VSS 0.114418f
C25704 DVDD.n8744 VSS 0.033368f
C25705 DVDD.n8745 VSS 0.029062f
C25706 DVDD.n8746 VSS 0.02691f
C25707 DVDD.n8747 VSS 0.060739f
C25708 DVDD.n8748 VSS 0.029062f
C25709 DVDD.n8749 VSS 0.220891f
C25710 DVDD.n8750 VSS 0.130242f
C25711 DVDD.n8751 VSS 0.130242f
C25712 DVDD.n8752 VSS 0.066735f
C25713 DVDD.n8753 VSS 0.201821f
C25714 DVDD.n8754 VSS 0.029062f
C25715 DVDD.n8755 VSS 0.02691f
C25716 DVDD.n8756 VSS 0.026274f
C25717 DVDD.n8757 VSS 0.060175f
C25718 DVDD.n8758 VSS 0.060175f
C25719 DVDD.n8759 VSS 0.026274f
C25720 DVDD.n8760 VSS 0.030088f
C25721 DVDD.n8761 VSS 0.029062f
C25722 DVDD.n8762 VSS 0.225658f
C25723 DVDD.n8763 VSS 0.066735f
C25724 DVDD.n8764 VSS 0.066735f
C25725 DVDD.n8765 VSS 0.225658f
C25726 DVDD.n8766 VSS 0.029062f
C25727 DVDD.n8767 VSS 0.033368f
C25728 DVDD.n8768 VSS 0.114418f
C25729 DVDD.n8769 VSS 0.114418f
C25730 DVDD.n8770 VSS 0.033368f
C25731 DVDD.n8771 VSS 0.029062f
C25732 DVDD.n8772 VSS 0.225658f
C25733 DVDD.n8773 VSS 0.013137f
C25734 DVDD.n8774 VSS 0.013137f
C25735 DVDD.n8775 VSS 0.131369f
C25736 DVDD.n8776 VSS 0.131369f
C25737 DVDD.n8777 VSS 0.013137f
C25738 DVDD.n8778 VSS 0.013137f
C25739 DVDD.n8779 VSS 0.013137f
C25740 DVDD.n8780 VSS 0.131369f
C25741 DVDD.n8781 VSS 0.451316f
C25742 DVDD.n8782 VSS 0.451316f
C25743 DVDD.n8783 VSS 0.344844f
C25744 DVDD.n8784 VSS 0.451316f
C25745 DVDD.n8785 VSS 0.451316f
C25746 DVDD.n8786 VSS 1.28214f
C25747 DVDD.n8787 VSS 0.429855f
C25748 DVDD.n8788 VSS 0.447648f
C25749 DVDD.n8789 VSS 0.013137f
C25750 DVDD.n8790 VSS 0.013137f
C25751 DVDD.n8791 VSS 0.131369f
C25752 DVDD.n8792 VSS 0.131369f
C25753 DVDD.n8793 VSS 0.124509f
C25754 DVDD.n8794 VSS 0.102976f
C25755 DVDD.n8795 VSS 0.102976f
C25756 DVDD.n8796 VSS 0.124509f
C25757 DVDD.t38 VSS 5.27557f
C25758 DVDD.n8797 VSS 0.114418f
C25759 DVDD.n8798 VSS 0.058124f
C25760 DVDD.n8799 VSS 0.114418f
C25761 DVDD.n8800 VSS 0.114418f
C25762 DVDD.n8801 VSS 0.032022f
C25763 DVDD.n8802 VSS 0.030408f
C25764 DVDD.n8803 VSS 0.114418f
C25765 DVDD.n8804 VSS 0.033368f
C25766 DVDD.n8805 VSS 0.114418f
C25767 DVDD.n8806 VSS 0.033368f
C25768 DVDD.n8807 VSS 0.114418f
C25769 DVDD.n8808 VSS 0.033368f
C25770 DVDD.n8809 VSS 0.114418f
C25771 DVDD.n8810 VSS 0.033368f
C25772 DVDD.n8811 VSS 0.114418f
C25773 DVDD.n8812 VSS 0.033368f
C25774 DVDD.n8813 VSS 0.114418f
C25775 DVDD.n8814 VSS 0.033368f
C25776 DVDD.n8815 VSS 0.114418f
C25777 DVDD.n8816 VSS 0.114418f
C25778 DVDD.n8817 VSS 0.030946f
C25779 DVDD.n8818 VSS 0.031484f
C25780 DVDD.n8819 VSS 0.114418f
C25781 DVDD.n8820 VSS 0.033368f
C25782 DVDD.n8821 VSS 0.114418f
C25783 DVDD.n8822 VSS 0.114418f
C25784 DVDD.n8823 VSS 0.051397f
C25785 DVDD.n8824 VSS 0.058124f
C25786 DVDD.n8825 VSS 0.058124f
C25787 DVDD.n8826 VSS 0.114418f
C25788 DVDD.n8827 VSS 0.114418f
C25789 DVDD.n8828 VSS 0.114418f
C25790 DVDD.n8829 VSS 0.058124f
C25791 DVDD.n8830 VSS 0.058124f
C25792 DVDD.n8831 VSS 0.058124f
C25793 DVDD.n8832 VSS 0.114418f
C25794 DVDD.n8833 VSS 0.114418f
C25795 DVDD.n8834 VSS 0.15585f
C25796 DVDD.n8835 VSS 0.277706f
C25797 DVDD.n8836 VSS 0.277706f
C25798 DVDD.n8837 VSS 0.15585f
C25799 DVDD.t14 VSS 5.27557f
C25800 DVDD.n8838 VSS 0.124509f
C25801 DVDD.n8839 VSS 0.131369f
C25802 DVDD.n8840 VSS 0.026274f
C25803 DVDD.n8841 VSS 0.026274f
C25804 DVDD.n8842 VSS 0.026274f
C25805 DVDD.n8843 VSS 0.131369f
C25806 DVDD.n8844 VSS 0.131369f
C25807 DVDD.n8845 VSS 0.131369f
C25808 DVDD.n8846 VSS 0.026274f
C25809 DVDD.n8847 VSS 0.026274f
C25810 DVDD.n8848 VSS 0.026274f
C25811 DVDD.n8849 VSS 0.131369f
C25812 DVDD.n8850 VSS 0.131369f
C25813 DVDD.n8851 VSS 0.131369f
C25814 DVDD.n8852 VSS 0.026274f
C25815 DVDD.n8853 VSS 0.026274f
C25816 DVDD.n8854 VSS 0.026274f
C25817 DVDD.n8855 VSS 0.131369f
C25818 DVDD.n8856 VSS 0.131369f
C25819 DVDD.n8857 VSS 0.131369f
C25820 DVDD.n8858 VSS 0.026274f
C25821 DVDD.n8859 VSS 0.026274f
C25822 DVDD.n8860 VSS 0.026274f
C25823 DVDD.n8861 VSS 0.131369f
C25824 DVDD.n8862 VSS 0.131369f
C25825 DVDD.n8863 VSS 0.131369f
C25826 DVDD.n8864 VSS 0.026274f
C25827 DVDD.n8865 VSS 0.026274f
C25828 DVDD.n8866 VSS 0.026274f
C25829 DVDD.n8867 VSS 0.131369f
C25830 DVDD.n8868 VSS 0.131369f
C25831 DVDD.n8869 VSS 0.131369f
C25832 DVDD.n8870 VSS 0.026274f
C25833 DVDD.n8871 VSS 0.026274f
C25834 DVDD.n8872 VSS 0.026274f
C25835 DVDD.n8873 VSS 0.131369f
C25836 DVDD.n8874 VSS 0.131369f
C25837 DVDD.n8875 VSS 0.124509f
C25838 DVDD.n8876 VSS 0.101549f
C25839 DVDD.n8877 VSS 0.11754f
C25840 DVDD.n8878 VSS 0.042564f
C25841 DVDD.n8879 VSS 0.131369f
C25842 DVDD.n8880 VSS 0.131369f
C25843 DVDD.n8881 VSS 0.131369f
C25844 DVDD.n8882 VSS 0.042564f
C25845 DVDD.n8883 VSS 0.042564f
C25846 DVDD.n8884 VSS 0.042564f
C25847 DVDD.n8885 VSS 0.131369f
C25848 DVDD.n8886 VSS 0.131369f
C25849 DVDD.n8887 VSS 0.131369f
C25850 DVDD.n8888 VSS 0.039704f
C25851 DVDD.n8889 VSS 0.277232f
C25852 DVDD.n8890 VSS 0.108274f
C25853 DVDD.n8891 VSS 1.01509f
C25854 DVDD.n8892 VSS 0.084542f
C25855 DVDD.n8893 VSS 0.027756f
C25856 DVDD.n8894 VSS 0.105307f
C25857 DVDD.n8895 VSS 0.091958f
C25858 DVDD.n8896 VSS 0.210614f
C25859 DVDD.n8897 VSS 0.210614f
C25860 DVDD.n8898 VSS 0.210614f
C25861 DVDD.n8899 VSS 0.210614f
C25862 DVDD.n8900 VSS 0.210614f
C25863 DVDD.n8901 VSS 0.171309f
C25864 DVDD.n8902 VSS 0.210614f
C25865 DVDD.n8903 VSS 0.210614f
C25866 DVDD.n8904 VSS 0.210614f
C25867 DVDD.n8905 VSS 0.210614f
C25868 DVDD.n8906 VSS 0.210614f
C25869 DVDD.n8907 VSS 0.210614f
C25870 DVDD.n8908 VSS 0.210614f
C25871 DVDD.n8909 VSS 0.184658f
C25872 DVDD.n8910 VSS 0.105307f
C25873 DVDD.n8911 VSS 1.85245f
C25874 DVDD.n8912 VSS 0.105307f
C25875 DVDD.n8913 VSS 0.091958f
C25876 DVDD.n8914 VSS 0.210614f
C25877 DVDD.n8915 VSS 0.210614f
C25878 DVDD.n8916 VSS 0.210614f
C25879 DVDD.n8917 VSS 0.210614f
C25880 DVDD.n8918 VSS 0.210614f
C25881 DVDD.n8919 VSS 0.171309f
C25882 DVDD.n8920 VSS 0.210614f
C25883 DVDD.n8921 VSS 0.210614f
C25884 DVDD.n8922 VSS 0.210614f
C25885 DVDD.n8923 VSS 0.210614f
C25886 DVDD.n8924 VSS 0.210614f
C25887 DVDD.n8925 VSS 0.210614f
C25888 DVDD.n8926 VSS 0.210614f
C25889 DVDD.n8927 VSS 0.210614f
C25890 DVDD.n8928 VSS 0.210614f
C25891 DVDD.n8929 VSS 0.210614f
C25892 DVDD.n8930 VSS 0.210614f
C25893 DVDD.n8931 VSS 0.210614f
C25894 DVDD.n8932 VSS 0.210614f
C25895 DVDD.n8933 VSS 0.210614f
C25896 DVDD.n8934 VSS 0.210614f
C25897 DVDD.n8935 VSS 0.184658f
C25898 DVDD.n8936 VSS 0.105307f
C25899 DVDD.n8937 VSS 0.029062f
C25900 DVDD.n8938 VSS 0.105307f
C25901 DVDD.n8939 VSS 0.171309f
C25902 DVDD.n8940 VSS 0.210614f
C25903 DVDD.n8941 VSS 0.210614f
C25904 DVDD.n8942 VSS 0.210614f
C25905 DVDD.n8943 VSS 0.210614f
C25906 DVDD.n8944 VSS 0.210614f
C25907 DVDD.n8945 VSS 0.210614f
C25908 DVDD.n8946 VSS 0.210614f
C25909 DVDD.n8947 VSS 0.210614f
C25910 DVDD.n8948 VSS 0.210614f
C25911 DVDD.n8949 VSS 0.210614f
C25912 DVDD.n8950 VSS 0.210614f
C25913 DVDD.n8951 VSS 0.210614f
C25914 DVDD.n8952 VSS 0.210614f
C25915 DVDD.n8953 VSS 0.210614f
C25916 DVDD.n8954 VSS 0.210614f
C25917 DVDD.n8955 VSS 0.210614f
C25918 DVDD.n8956 VSS 0.210614f
C25919 DVDD.n8957 VSS 0.210614f
C25920 DVDD.n8958 VSS 0.210614f
C25921 DVDD.n8959 VSS 0.210614f
C25922 DVDD.n8960 VSS 0.210614f
C25923 DVDD.n8961 VSS 0.210614f
C25924 DVDD.n8962 VSS 0.210614f
C25925 DVDD.n8963 VSS 0.184658f
C25926 DVDD.n8964 VSS 0.210614f
C25927 DVDD.n8965 VSS 0.091958f
C25928 DVDD.n8966 VSS 0.210614f
C25929 DVDD.n8967 VSS 0.210614f
C25930 DVDD.n8968 VSS 0.210614f
C25931 DVDD.n8969 VSS 0.210614f
C25932 DVDD.n8970 VSS 0.210614f
C25933 DVDD.n8971 VSS 0.091958f
C25934 DVDD.n8972 VSS 0.029062f
C25935 DVDD.n8973 VSS 0.029062f
C25936 DVDD.n8974 VSS 0.029062f
C25937 DVDD.n8975 VSS 0.029062f
C25938 DVDD.n8976 VSS 0.033368f
C25939 DVDD.n8977 VSS 0.114418f
C25940 DVDD.n8978 VSS 0.030408f
C25941 DVDD.n8979 VSS 0.032022f
C25942 DVDD.n8980 VSS 0.114418f
C25943 DVDD.n8981 VSS 0.033368f
C25944 DVDD.n8982 VSS 0.114418f
C25945 DVDD.n8983 VSS 0.033368f
C25946 DVDD.n8984 VSS 0.114418f
C25947 DVDD.n8985 VSS 0.033368f
C25948 DVDD.n8986 VSS 0.114418f
C25949 DVDD.n8987 VSS 0.033368f
C25950 DVDD.n8988 VSS 0.114418f
C25951 DVDD.n8989 VSS 0.114418f
C25952 DVDD.n8990 VSS 0.114418f
C25953 DVDD.n8991 VSS 0.058124f
C25954 DVDD.n8992 VSS 0.114418f
C25955 DVDD.n8993 VSS 0.114418f
C25956 DVDD.n8994 VSS 0.058124f
C25957 DVDD.n8995 VSS 0.058124f
C25958 DVDD.n8996 VSS 0.058124f
C25959 DVDD.n8997 VSS 0.114418f
C25960 DVDD.n8998 VSS 0.114418f
C25961 DVDD.n8999 VSS 0.114418f
C25962 DVDD.n9000 VSS 0.058124f
C25963 DVDD.n9001 VSS 0.058124f
C25964 DVDD.n9002 VSS 0.049783f
C25965 DVDD.n9003 VSS 0.114418f
C25966 DVDD.n9004 VSS 0.033368f
C25967 DVDD.n9005 VSS 0.114418f
C25968 DVDD.n9006 VSS 0.114418f
C25969 DVDD.n9007 VSS 0.033099f
C25970 DVDD.n9008 VSS 0.029331f
C25971 DVDD.n9009 VSS 0.114418f
C25972 DVDD.n9010 VSS 0.114418f
C25973 DVDD.n9011 VSS 0.033368f
C25974 DVDD.n9012 VSS 0.029062f
C25975 DVDD.n9013 VSS 0.105307f
C25976 DVDD.n9014 VSS 0.754582f
C25977 DVDD.n9015 VSS 0.747408f
C25978 DVDD.t26 VSS 5.27557f
C25979 DVDD.n9017 VSS 0.15585f
C25980 DVDD.n9018 VSS 0.277706f
C25981 DVDD.n9019 VSS 0.058124f
C25982 DVDD.n9020 VSS 0.114418f
C25983 DVDD.n9021 VSS 0.058124f
C25984 DVDD.n9022 VSS 0.114418f
C25985 DVDD.n9023 VSS 0.058124f
C25986 DVDD.n9024 VSS 0.114418f
C25987 DVDD.n9025 VSS 0.058124f
C25988 DVDD.n9026 VSS 0.114418f
C25989 DVDD.n9027 VSS 0.058124f
C25990 DVDD.n9028 VSS 0.114418f
C25991 DVDD.n9029 VSS 0.058124f
C25992 DVDD.n9030 VSS 0.114418f
C25993 DVDD.n9031 VSS 0.114418f
C25994 DVDD.n9032 VSS 0.058124f
C25995 DVDD.n9033 VSS 0.058124f
C25996 DVDD.n9034 VSS 0.058124f
C25997 DVDD.n9035 VSS 0.114418f
C25998 DVDD.n9036 VSS 0.114418f
C25999 DVDD.n9037 VSS 0.114418f
C26000 DVDD.n9038 VSS 0.058124f
C26001 DVDD.n9039 VSS 0.058124f
C26002 DVDD.n9040 VSS 0.058124f
C26003 DVDD.n9041 VSS 0.114418f
C26004 DVDD.n9042 VSS 0.114418f
C26005 DVDD.n9043 VSS 0.114418f
C26006 DVDD.n9044 VSS 0.058124f
C26007 DVDD.n9045 VSS 0.058124f
C26008 DVDD.n9046 VSS 0.058124f
C26009 DVDD.n9047 VSS 0.114418f
C26010 DVDD.n9048 VSS 0.114418f
C26011 DVDD.n9049 VSS 0.114418f
C26012 DVDD.n9050 VSS 0.058124f
C26013 DVDD.n9051 VSS 0.058124f
C26014 DVDD.n9052 VSS 0.058124f
C26015 DVDD.n9053 VSS 0.114418f
C26016 DVDD.n9054 VSS 0.114418f
C26017 DVDD.n9055 VSS 0.114418f
C26018 DVDD.n9056 VSS 0.058124f
C26019 DVDD.n9057 VSS 0.058124f
C26020 DVDD.n9058 VSS 0.058124f
C26021 DVDD.n9059 VSS 0.114418f
C26022 DVDD.n9060 VSS 0.114418f
C26023 DVDD.n9061 VSS 0.114418f
C26024 DVDD.n9062 VSS 0.058124f
C26025 DVDD.n9063 VSS 0.058124f
C26026 DVDD.n9064 VSS 0.058124f
C26027 DVDD.n9065 VSS 0.114418f
C26028 DVDD.n9066 VSS 0.114418f
C26029 DVDD.n9067 VSS 0.114418f
C26030 DVDD.n9068 VSS 0.058124f
C26031 DVDD.n9069 VSS 0.058124f
C26032 DVDD.n9070 VSS 0.277706f
C26033 DVDD.n9071 VSS 0.15585f
C26034 DVDD.t29 VSS 5.27557f
C26035 DVDD.n9073 VSS 0.15585f
C26036 DVDD.n9074 VSS 0.277706f
C26037 DVDD.n9075 VSS 0.058124f
C26038 DVDD.n9076 VSS 0.114418f
C26039 DVDD.n9077 VSS 0.058124f
C26040 DVDD.n9078 VSS 0.033368f
C26041 DVDD.n9079 VSS 0.114418f
C26042 DVDD.n9080 VSS 0.033368f
C26043 DVDD.n9081 VSS 0.114418f
C26044 DVDD.n9082 VSS 0.033368f
C26045 DVDD.n9083 VSS 0.114418f
C26046 DVDD.n9084 VSS 0.033368f
C26047 DVDD.n9085 VSS 0.114418f
C26048 DVDD.n9086 VSS 0.033368f
C26049 DVDD.n9087 VSS 0.114418f
C26050 DVDD.n9088 VSS 0.114418f
C26051 DVDD.n9089 VSS 0.030946f
C26052 DVDD.n9090 VSS 0.031484f
C26053 DVDD.n9091 VSS 0.114418f
C26054 DVDD.n9092 VSS 0.033368f
C26055 DVDD.n9093 VSS 0.114418f
C26056 DVDD.n9094 VSS 0.051397f
C26057 DVDD.n9095 VSS 0.114418f
C26058 DVDD.n9096 VSS 0.114418f
C26059 DVDD.n9097 VSS 0.114418f
C26060 DVDD.n9098 VSS 0.058124f
C26061 DVDD.n9099 VSS 0.058124f
C26062 DVDD.n9100 VSS 0.058124f
C26063 DVDD.n9101 VSS 0.114418f
C26064 DVDD.n9102 VSS 0.114418f
C26065 DVDD.n9103 VSS 0.114418f
C26066 DVDD.n9104 VSS 0.058124f
C26067 DVDD.n9105 VSS 0.058124f
C26068 DVDD.n9106 VSS 0.277706f
C26069 DVDD.n9107 VSS 0.15585f
C26070 DVDD.t23 VSS 5.27557f
C26071 DVDD.n9109 VSS 0.15585f
C26072 DVDD.n9110 VSS 0.114418f
C26073 DVDD.n9111 VSS 0.058124f
C26074 DVDD.n9112 VSS 0.058124f
C26075 DVDD.n9113 VSS 0.058124f
C26076 DVDD.n9114 VSS 0.114418f
C26077 DVDD.n9115 VSS 0.114418f
C26078 DVDD.n9116 VSS 0.114418f
C26079 DVDD.n9117 VSS 0.058124f
C26080 DVDD.n9118 VSS 0.058124f
C26081 DVDD.n9119 VSS 0.050859f
C26082 DVDD.n9120 VSS 0.114418f
C26083 DVDD.n9121 VSS 0.033368f
C26084 DVDD.n9122 VSS 0.114418f
C26085 DVDD.n9123 VSS 0.114418f
C26086 DVDD.n9124 VSS 0.114418f
C26087 DVDD.n9125 VSS 0.030408f
C26088 DVDD.n9126 VSS 0.091958f
C26089 DVDD.n9127 VSS 0.210614f
C26090 DVDD.n9128 VSS 0.210614f
C26091 DVDD.n9129 VSS 0.210614f
C26092 DVDD.n9130 VSS 0.210614f
C26093 DVDD.n9131 VSS 0.210614f
C26094 DVDD.n9132 VSS 0.210614f
C26095 DVDD.n9133 VSS 0.210614f
C26096 DVDD.n9134 VSS 0.184658f
C26097 DVDD.n9135 VSS 0.210614f
C26098 DVDD.n9136 VSS 0.210614f
C26099 DVDD.n9137 VSS 0.210614f
C26100 DVDD.n9138 VSS 0.210614f
C26101 DVDD.n9139 VSS 0.210614f
C26102 DVDD.n9140 VSS 0.210614f
C26103 DVDD.n9141 VSS 0.210614f
C26104 DVDD.n9142 VSS 0.210614f
C26105 DVDD.n9143 VSS 0.171309f
C26106 DVDD.n9144 VSS 0.210614f
C26107 DVDD.n9145 VSS 0.210614f
C26108 DVDD.n9146 VSS 0.210614f
C26109 DVDD.n9147 VSS 0.210614f
C26110 DVDD.n9148 VSS 0.210614f
C26111 DVDD.n9149 VSS 0.210614f
C26112 DVDD.n9150 VSS 0.210614f
C26113 DVDD.n9151 VSS 0.210614f
C26114 DVDD.n9152 VSS 0.210614f
C26115 DVDD.n9153 VSS 0.210614f
C26116 DVDD.n9154 VSS 0.210614f
C26117 DVDD.n9155 VSS 0.210614f
C26118 DVDD.n9156 VSS 0.210614f
C26119 DVDD.n9157 VSS 0.210614f
C26120 DVDD.n9158 VSS 0.210614f
C26121 DVDD.n9159 VSS 0.210614f
C26122 DVDD.n9160 VSS 0.210614f
C26123 DVDD.n9161 VSS 0.210614f
C26124 DVDD.n9162 VSS 0.210614f
C26125 DVDD.n9163 VSS 0.210614f
C26126 DVDD.n9164 VSS 0.210614f
C26127 DVDD.n9165 VSS 0.210614f
C26128 DVDD.n9166 VSS 0.210614f
C26129 DVDD.n9167 VSS 0.210614f
C26130 DVDD.n9168 VSS 0.210614f
C26131 DVDD.n9169 VSS 0.210614f
C26132 DVDD.n9170 VSS 0.210614f
C26133 DVDD.n9171 VSS 0.210614f
C26134 DVDD.n9172 VSS 0.091958f
C26135 DVDD.n9173 VSS 0.105307f
C26136 DVDD.n9174 VSS 0.029062f
C26137 DVDD.n9175 VSS 0.105307f
C26138 DVDD.n9176 VSS 0.171309f
C26139 DVDD.n9177 VSS 0.210614f
C26140 DVDD.n9178 VSS 0.210614f
C26141 DVDD.n9179 VSS 0.210614f
C26142 DVDD.n9180 VSS 0.210614f
C26143 DVDD.n9181 VSS 0.210614f
C26144 DVDD.n9182 VSS 0.210614f
C26145 DVDD.n9183 VSS 0.210614f
C26146 DVDD.n9184 VSS 0.210614f
C26147 DVDD.n9185 VSS 0.210614f
C26148 DVDD.n9186 VSS 0.210614f
C26149 DVDD.n9187 VSS 0.210614f
C26150 DVDD.n9188 VSS 0.210614f
C26151 DVDD.n9189 VSS 0.210614f
C26152 DVDD.n9190 VSS 0.210614f
C26153 DVDD.n9191 VSS 0.210614f
C26154 DVDD.n9192 VSS 0.210614f
C26155 DVDD.n9193 VSS 0.210614f
C26156 DVDD.n9194 VSS 0.210614f
C26157 DVDD.n9195 VSS 0.210614f
C26158 DVDD.n9196 VSS 0.210614f
C26159 DVDD.n9197 VSS 0.210614f
C26160 DVDD.n9198 VSS 0.210614f
C26161 DVDD.n9199 VSS 0.210614f
C26162 DVDD.n9200 VSS 0.210614f
C26163 DVDD.n9201 VSS 0.210614f
C26164 DVDD.n9202 VSS 0.210614f
C26165 DVDD.n9203 VSS 0.210614f
C26166 DVDD.n9204 VSS 0.210614f
C26167 DVDD.n9205 VSS 0.210614f
C26168 DVDD.n9206 VSS 0.210614f
C26169 DVDD.n9207 VSS 0.168343f
C26170 DVDD.n9208 VSS 0.105307f
C26171 DVDD.n9209 VSS 0.029062f
C26172 DVDD.n9210 VSS 0.105307f
C26173 DVDD.n9211 VSS 0.187625f
C26174 DVDD.n9212 VSS 0.210614f
C26175 DVDD.n9213 VSS 0.210614f
C26176 DVDD.n9214 VSS 0.210614f
C26177 DVDD.n9215 VSS 0.210614f
C26178 DVDD.n9216 VSS 0.210614f
C26179 DVDD.n9217 VSS 0.210614f
C26180 DVDD.n9218 VSS 0.210614f
C26181 DVDD.n9219 VSS 0.210614f
C26182 DVDD.n9220 VSS 0.210614f
C26183 DVDD.n9221 VSS 0.210614f
C26184 DVDD.n9222 VSS 0.210614f
C26185 DVDD.n9223 VSS 0.210614f
C26186 DVDD.n9224 VSS 0.210614f
C26187 DVDD.n9225 VSS 0.210614f
C26188 DVDD.n9226 VSS 0.210614f
C26189 DVDD.n9227 VSS 0.210614f
C26190 DVDD.n9228 VSS 0.210614f
C26191 DVDD.n9229 VSS 0.210614f
C26192 DVDD.n9230 VSS 0.210614f
C26193 DVDD.n9231 VSS 0.210614f
C26194 DVDD.n9232 VSS 0.210614f
C26195 DVDD.n9233 VSS 0.210614f
C26196 DVDD.n9234 VSS 0.210614f
C26197 DVDD.n9235 VSS 0.168343f
C26198 DVDD.n9236 VSS 0.210614f
C26199 DVDD.n9237 VSS 0.091958f
C26200 DVDD.n9238 VSS 0.210614f
C26201 DVDD.n9239 VSS 0.210614f
C26202 DVDD.n9240 VSS 0.210614f
C26203 DVDD.n9241 VSS 0.210614f
C26204 DVDD.n9242 VSS 0.210614f
C26205 DVDD.n9243 VSS 0.091958f
C26206 DVDD.n9244 VSS 0.029062f
C26207 DVDD.n9245 VSS 0.029062f
C26208 DVDD.n9246 VSS 0.029062f
C26209 DVDD.n9247 VSS 0.029062f
C26210 DVDD.n9248 VSS 0.029062f
C26211 DVDD.n9249 VSS 0.033368f
C26212 DVDD.n9250 VSS 0.032022f
C26213 DVDD.n9251 VSS 0.114418f
C26214 DVDD.n9252 VSS 0.031484f
C26215 DVDD.n9253 VSS 0.030946f
C26216 DVDD.n9254 VSS 0.114418f
C26217 DVDD.n9255 VSS 0.033368f
C26218 DVDD.n9256 VSS 0.114418f
C26219 DVDD.n9257 VSS 0.033368f
C26220 DVDD.n9258 VSS 0.114418f
C26221 DVDD.n9259 VSS 0.033368f
C26222 DVDD.n9260 VSS 0.114418f
C26223 DVDD.n9261 VSS 0.033368f
C26224 DVDD.n9262 VSS 0.114418f
C26225 DVDD.n9263 VSS 0.033368f
C26226 DVDD.n9264 VSS 0.114418f
C26227 DVDD.n9265 VSS 0.114418f
C26228 DVDD.n9266 VSS 0.114418f
C26229 DVDD.n9267 VSS 0.058124f
C26230 DVDD.n9268 VSS 0.114418f
C26231 DVDD.n9269 VSS 0.058124f
C26232 DVDD.n9270 VSS 0.058124f
C26233 DVDD.n9271 VSS 0.114418f
C26234 DVDD.n9272 VSS 0.114418f
C26235 DVDD.n9273 VSS 0.114418f
C26236 DVDD.n9274 VSS 0.058124f
C26237 DVDD.n9275 VSS 0.058124f
C26238 DVDD.n9276 VSS 0.050859f
C26239 DVDD.n9277 VSS 0.114418f
C26240 DVDD.n9278 VSS 0.033368f
C26241 DVDD.n9279 VSS 0.114418f
C26242 DVDD.n9280 VSS 0.114418f
C26243 DVDD.n9281 VSS 0.114418f
C26244 DVDD.n9282 VSS 0.030408f
C26245 DVDD.n9283 VSS 0.029062f
C26246 DVDD.n9284 VSS 0.105307f
C26247 DVDD.n9285 VSS 0.029062f
C26248 DVDD.n9286 VSS 0.051397f
C26249 DVDD.n9287 VSS 0.114418f
C26250 DVDD.n9288 VSS 0.114418f
C26251 DVDD.n9289 VSS 0.114418f
C26252 DVDD.n9290 VSS 0.058124f
C26253 DVDD.n9291 VSS 0.058124f
C26254 DVDD.n9292 VSS 0.058124f
C26255 DVDD.n9293 VSS 0.114418f
C26256 DVDD.n9294 VSS 0.114418f
C26257 DVDD.n9295 VSS 0.114418f
C26258 DVDD.n9296 VSS 0.058124f
C26259 DVDD.n9297 VSS 0.058124f
C26260 DVDD.n9298 VSS 0.277706f
C26261 DVDD.n9299 VSS 0.15585f
C26262 DVDD.t32 VSS 5.27557f
C26263 DVDD.n9300 VSS 0.15585f
C26264 DVDD.n9301 VSS 0.277706f
C26265 DVDD.n9302 VSS 0.277706f
C26266 DVDD.n9303 VSS 0.05355f
C26267 DVDD.n9304 VSS 0.114418f
C26268 DVDD.n9305 VSS 0.114418f
C26269 DVDD.n9306 VSS 0.114418f
C26270 DVDD.n9307 VSS 0.114418f
C26271 DVDD.n9308 VSS 0.114418f
C26272 DVDD.n9309 VSS 0.114418f
C26273 DVDD.n9310 VSS 0.114418f
C26274 DVDD.n9311 VSS 0.033368f
C26275 DVDD.n9312 VSS 0.029062f
C26276 DVDD.n9313 VSS 0.029028f
C26277 DVDD.n9314 VSS 0.027333f
C26278 DVDD.n9315 VSS 0.029062f
C26279 DVDD.n9316 VSS 0.204999f
C26280 DVDD.n9317 VSS 0.066735f
C26281 DVDD.n9318 VSS 0.560793f
C26282 DVDD.n9319 VSS 0.447648f
C26283 DVDD.n9320 VSS 0.429855f
C26284 DVDD.n9321 VSS 1.28214f
C26285 DVDD.n9322 VSS 0.451316f
C26286 DVDD.n9323 VSS 0.451316f
C26287 DVDD.n9324 VSS 0.344844f
C26288 DVDD.n9325 VSS 0.344844f
C26289 DVDD.n9326 VSS 0.451316f
C26290 DVDD.n9327 VSS 0.225658f
C26291 DVDD.n9328 VSS 0.197054f
C26292 DVDD.n9329 VSS 0.197054f
C26293 DVDD.n9330 VSS 0.451316f
C26294 DVDD.n9331 VSS 0.750075f
C26295 DVDD.n9332 VSS 0.451316f
C26296 DVDD.n9333 VSS 0.332131f
C26297 DVDD.n9334 VSS 0.451316f
C26298 DVDD.n9335 VSS 0.451316f
C26299 DVDD.n9336 VSS 0.451316f
C26300 DVDD.n9337 VSS 0.451316f
C26301 DVDD.n9338 VSS 0.451316f
C26302 DVDD.n9339 VSS 0.750075f
C26303 DVDD.n9340 VSS 0.750075f
C26304 DVDD.n9341 VSS 0.750075f
C26305 DVDD.n9342 VSS 0.451316f
C26306 DVDD.n9343 VSS 0.451316f
C26307 DVDD.n9344 VSS 0.451316f
C26308 DVDD.n9345 VSS 0.451316f
C26309 DVDD.n9346 VSS 0.332131f
C26310 DVDD.n9347 VSS 0.332131f
C26311 DVDD.n9348 VSS 0.060175f
C26312 DVDD.n9349 VSS 0.030088f
C26313 DVDD.n9350 VSS 0.026274f
C26314 DVDD.n9351 VSS 0.060175f
C26315 DVDD.n9352 VSS 0.044284f
C26316 DVDD.n9353 VSS 0.044284f
C26317 DVDD.n9354 VSS 3.42659f
C26318 DVDD.n9355 VSS 0.045979f
C26319 DVDD.n9356 VSS 0.060175f
C26320 DVDD.n9357 VSS 0.060175f
C26321 DVDD.n9358 VSS 0.026274f
C26322 DVDD.n9359 VSS 0.030088f
C26323 DVDD.n9360 VSS 0.029062f
C26324 DVDD.n9361 VSS 0.225658f
C26325 DVDD.n9362 VSS 0.033368f
C26326 DVDD.n9363 VSS 0.033368f
C26327 DVDD.n9364 VSS 0.131369f
C26328 DVDD.n9365 VSS 0.033368f
C26329 DVDD.n9366 VSS 0.131369f
C26330 DVDD.n9367 VSS 0.033368f
C26331 DVDD.n9368 VSS 0.131369f
C26332 DVDD.n9369 VSS 0.131369f
C26333 DVDD.n9370 VSS 0.033368f
C26334 DVDD.n9371 VSS 0.033368f
C26335 DVDD.n9372 VSS 0.033368f
C26336 DVDD.n9373 VSS 0.033368f
C26337 DVDD.n9374 VSS 0.033368f
C26338 DVDD.n9375 VSS 0.131369f
C26339 DVDD.n9376 VSS 0.131369f
C26340 DVDD.n9377 VSS 0.036328f
C26341 DVDD.n9378 VSS 0.066735f
C26342 DVDD.n9379 VSS 0.060546f
C26343 DVDD.n9380 VSS 0.131369f
C26344 DVDD.n9381 VSS 0.131369f
C26345 DVDD.n9382 VSS 0.033368f
C26346 DVDD.n9383 VSS 0.033368f
C26347 DVDD.n9384 VSS 0.033368f
C26348 DVDD.n9385 VSS 0.131369f
C26349 DVDD.n9386 VSS 0.033368f
C26350 DVDD.n9387 VSS 0.131369f
C26351 DVDD.n9388 VSS 0.131369f
C26352 DVDD.n9389 VSS 0.033368f
C26353 DVDD.n9390 VSS 0.033368f
C26354 DVDD.n9391 VSS 0.225658f
C26355 DVDD.n9392 VSS 0.029062f
C26356 DVDD.n9393 VSS 0.033368f
C26357 DVDD.n9394 VSS 0.114418f
C26358 DVDD.n9395 VSS 0.114418f
C26359 DVDD.n9396 VSS 0.114418f
C26360 DVDD.n9397 VSS 0.033368f
C26361 DVDD.n9398 VSS 0.225658f
C26362 DVDD.n9399 VSS 0.029062f
C26363 DVDD.n9400 VSS 0.030088f
C26364 DVDD.n9401 VSS 0.026274f
C26365 DVDD.n9402 VSS 0.030088f
C26366 DVDD.n9403 VSS 0.026274f
C26367 DVDD.n9404 VSS 0.060175f
C26368 DVDD.n9405 VSS 0.170688f
C26369 DVDD.n9406 VSS 0.057608f
C26370 DVDD.n9407 VSS 0.059656f
C26371 DVDD.n9408 VSS 0.10091f
C26372 DVDD.n9409 VSS 0.033099f
C26373 DVDD.n9410 VSS 0.029331f
C26374 DVDD.n9411 VSS 0.114418f
C26375 DVDD.n9412 VSS 0.114418f
C26376 DVDD.n9413 VSS 0.033368f
C26377 DVDD.n9414 VSS 0.029062f
C26378 DVDD.n9415 VSS 0.217712f
C26379 DVDD.n9416 VSS 0.066735f
C26380 DVDD.n9417 VSS 0.066735f
C26381 DVDD.n9418 VSS 0.225658f
C26382 DVDD.n9419 VSS 0.033368f
C26383 DVDD.n9420 VSS 0.033368f
C26384 DVDD.n9421 VSS 0.131369f
C26385 DVDD.n9422 VSS 0.131369f
C26386 DVDD.n9423 VSS 0.033368f
C26387 DVDD.n9424 VSS 0.033368f
C26388 DVDD.n9425 VSS 3.34178f
C26389 DVDD.n9426 VSS 0.451316f
C26390 DVDD.n9427 VSS 0.451316f
C26391 DVDD.n9428 VSS 0.451316f
C26392 DVDD.n9429 VSS 0.332131f
C26393 DVDD.n9430 VSS 0.197054f
C26394 DVDD.n9431 VSS 0.225658f
C26395 DVDD.n9432 VSS 0.029062f
C26396 DVDD.n9433 VSS 0.033368f
C26397 DVDD.n9434 VSS 0.114418f
C26398 DVDD.n9435 VSS 0.114418f
C26399 DVDD.n9436 VSS 0.114418f
C26400 DVDD.n9437 VSS 0.030408f
C26401 DVDD.n9438 VSS 0.029062f
C26402 DVDD.n9439 VSS 0.225658f
C26403 DVDD.n9440 VSS 0.197054f
C26404 DVDD.n9441 VSS 0.451316f
C26405 DVDD.n9442 VSS 0.750075f
C26406 DVDD.n9443 VSS 0.750075f
C26407 DVDD.n9444 VSS 0.548254f
C26408 DVDD.n9445 VSS 0.220891f
C26409 DVDD.n9446 VSS 0.029062f
C26410 DVDD.n9447 VSS 0.033368f
C26411 DVDD.n9448 VSS 0.114418f
C26412 DVDD.n9449 VSS 0.114418f
C26413 DVDD.n9450 VSS 0.033368f
C26414 DVDD.n9451 VSS 0.029062f
C26415 DVDD.n9452 VSS 0.225658f
C26416 DVDD.n9453 VSS 0.197054f
C26417 DVDD.n9454 VSS 0.451316f
C26418 DVDD.n9455 VSS 0.451316f
C26419 DVDD.n9456 VSS 0.197054f
C26420 DVDD.n9457 VSS 0.225658f
C26421 DVDD.n9458 VSS 0.029062f
C26422 DVDD.n9459 VSS 0.033368f
C26423 DVDD.n9460 VSS 0.114418f
C26424 DVDD.n9461 VSS 0.033368f
C26425 DVDD.n9462 VSS 0.114418f
C26426 DVDD.n9463 VSS 0.114418f
C26427 DVDD.n9464 VSS 0.033368f
C26428 DVDD.n9465 VSS 0.029062f
C26429 DVDD.n9466 VSS 0.225658f
C26430 DVDD.n9467 VSS 0.197054f
C26431 DVDD.n9468 VSS 0.451316f
C26432 DVDD.n9469 VSS 0.451316f
C26433 DVDD.n9470 VSS 0.197054f
C26434 DVDD.n9471 VSS 0.447648f
C26435 DVDD.n9472 VSS 0.029062f
C26436 DVDD.n9473 VSS 0.05355f
C26437 DVDD.n9474 VSS 0.277706f
C26438 DVDD.n9475 VSS 0.15585f
C26439 DVDD.t2 VSS 5.27557f
C26440 DVDD.n9477 VSS 0.15585f
C26441 DVDD.n9478 VSS 0.029331f
C26442 DVDD.n9479 VSS 0.114418f
C26443 DVDD.n9480 VSS 0.114418f
C26444 DVDD.n9481 VSS 0.033368f
C26445 DVDD.n9482 VSS 0.029062f
C26446 DVDD.n9483 VSS 0.217712f
C26447 DVDD.n9484 VSS 0.197054f
C26448 DVDD.n9485 VSS 0.451316f
C26449 DVDD.n9486 VSS 0.451316f
C26450 DVDD.n9487 VSS 0.451316f
C26451 DVDD.n9488 VSS 0.724649f
C26452 DVDD.n9489 VSS 0.724649f
C26453 DVDD.n9490 VSS 0.535541f
C26454 DVDD.n9491 VSS 0.225658f
C26455 DVDD.n9492 VSS 0.10091f
C26456 DVDD.n9493 VSS 0.130242f
C26457 DVDD.n9494 VSS 0.066735f
C26458 DVDD.n9495 VSS 0.066735f
C26459 DVDD.n9496 VSS 0.204999f
C26460 DVDD.n9497 VSS 0.197054f
C26461 DVDD.n9498 VSS 0.451316f
C26462 DVDD.n9499 VSS 0.451316f
C26463 DVDD.n9500 VSS 0.451316f
C26464 DVDD.n9501 VSS 0.451316f
C26465 DVDD.n9502 VSS 0.451316f
C26466 DVDD.n9503 VSS 0.197054f
C26467 DVDD.n9504 VSS 0.197054f
C26468 DVDD.n9505 VSS 0.225658f
C26469 DVDD.n9506 VSS 0.04763f
C26470 DVDD.n9507 VSS 0.029062f
C26471 DVDD.n9508 VSS 0.033368f
C26472 DVDD.n9509 VSS 0.029062f
C26473 DVDD.n9510 VSS 0.033368f
C26474 DVDD.n9511 VSS 0.15585f
C26475 DVDD.t17 VSS 5.27557f
C26476 DVDD.n9513 VSS 0.15585f
C26477 DVDD.n9514 VSS 0.114418f
C26478 DVDD.n9515 VSS 0.058124f
C26479 DVDD.n9516 VSS 0.058124f
C26480 DVDD.n9517 VSS 0.058124f
C26481 DVDD.n9518 VSS 0.114418f
C26482 DVDD.n9519 VSS 0.114418f
C26483 DVDD.n9520 VSS 0.114418f
C26484 DVDD.n9521 VSS 0.058124f
C26485 DVDD.n9522 VSS 0.058124f
C26486 DVDD.n9523 VSS 0.058124f
C26487 DVDD.n9524 VSS 0.114418f
C26488 DVDD.n9525 VSS 0.114418f
C26489 DVDD.n9526 VSS 0.114418f
C26490 DVDD.n9527 VSS 0.058124f
C26491 DVDD.n9528 VSS 0.058124f
C26492 DVDD.n9529 VSS 0.058124f
C26493 DVDD.n9530 VSS 0.114418f
C26494 DVDD.n9531 VSS 0.114418f
C26495 DVDD.n9532 VSS 0.114418f
C26496 DVDD.n9533 VSS 0.058124f
C26497 DVDD.n9534 VSS 0.058124f
C26498 DVDD.n9535 VSS 0.058124f
C26499 DVDD.n9536 VSS 0.114418f
C26500 DVDD.n9537 VSS 0.114418f
C26501 DVDD.n9538 VSS 0.114418f
C26502 DVDD.n9539 VSS 0.058124f
C26503 DVDD.n9540 VSS 0.058124f
C26504 DVDD.n9541 VSS 0.058124f
C26505 DVDD.n9542 VSS 0.114418f
C26506 DVDD.n9543 VSS 0.114418f
C26507 DVDD.n9544 VSS 0.114418f
C26508 DVDD.n9545 VSS 0.046553f
C26509 DVDD.n9546 VSS 0.029062f
C26510 DVDD.n9547 VSS 0.456124f
C26511 DVDD.n9548 VSS 0.201821f
C26512 DVDD.n9549 VSS 0.029062f
C26513 DVDD.n9550 VSS 0.033368f
C26514 DVDD.n9551 VSS 0.114418f
C26515 DVDD.n9552 VSS 0.114418f
C26516 DVDD.n9553 VSS 0.114418f
C26517 DVDD.n9554 VSS 0.030408f
C26518 DVDD.n9555 VSS 0.029062f
C26519 DVDD.n9556 VSS 0.225658f
C26520 DVDD.n9557 VSS 0.197054f
C26521 DVDD.n9558 VSS 0.451316f
C26522 DVDD.n9559 VSS 0.451316f
C26523 DVDD.n9560 VSS 0.332131f
C26524 DVDD.n9561 VSS 3.4242f
C26525 DVDD.n9562 VSS 0.556669f
C26526 DVDD.n9563 VSS 1.62732f
C26527 DVDD.n9564 VSS 0.344844f
C26528 DVDD.n9565 VSS 0.451316f
C26529 DVDD.n9566 VSS 0.451316f
C26530 DVDD.n9567 VSS 0.451316f
C26531 DVDD.n9568 VSS 0.451316f
C26532 DVDD.n9569 VSS 0.451316f
C26533 DVDD.n9570 VSS 0.724649f
C26534 DVDD.n9571 VSS 0.724649f
C26535 DVDD.n9572 VSS 0.724649f
C26536 DVDD.n9573 VSS 0.451316f
C26537 DVDD.n9574 VSS 0.451316f
C26538 DVDD.n9575 VSS 0.451316f
C26539 DVDD.n9576 VSS 0.451316f
C26540 DVDD.n9577 VSS 0.344844f
C26541 DVDD.n9578 VSS 0.344844f
C26542 DVDD.n9579 VSS 3.44612f
C26543 DVDD.n9580 VSS 0.044284f
C26544 DVDD.n9581 VSS 0.060175f
C26545 DVDD.n9582 VSS 0.060175f
C26546 DVDD.n9583 VSS 0.026274f
C26547 DVDD.n9584 VSS 0.030088f
C26548 DVDD.n9585 VSS 0.029062f
C26549 DVDD.n9586 VSS 0.225658f
C26550 DVDD.n9587 VSS 0.066735f
C26551 DVDD.n9588 VSS 0.066735f
C26552 DVDD.n9589 VSS 0.225658f
C26553 DVDD.n9590 VSS 0.029062f
C26554 DVDD.n9591 VSS 0.033368f
C26555 DVDD.n9592 VSS 0.114418f
C26556 DVDD.n9593 VSS 0.114418f
C26557 DVDD.n9594 VSS 0.033368f
C26558 DVDD.n9595 VSS 0.029062f
C26559 DVDD.n9596 VSS 0.220891f
C26560 DVDD.n9597 VSS 0.130242f
C26561 DVDD.n9598 VSS 0.130242f
C26562 DVDD.n9599 VSS 0.220891f
C26563 DVDD.n9600 VSS 0.029062f
C26564 DVDD.n9601 VSS 0.060786f
C26565 DVDD.n9602 VSS 0.061067f
C26566 DVDD.n9603 VSS 0.060175f
C26567 DVDD.n9604 VSS 0.026274f
C26568 DVDD.n9605 VSS 0.030088f
C26569 DVDD.n9606 VSS 0.029062f
C26570 DVDD.n9607 VSS 0.029869f
C26571 DVDD.n9608 VSS 0.032561f
C26572 DVDD.n9609 VSS 0.114418f
C26573 DVDD.n9610 VSS 0.114418f
C26574 DVDD.n9611 VSS 0.033368f
C26575 DVDD.n9612 VSS 0.029062f
C26576 DVDD.n9613 VSS 0.225658f
C26577 DVDD.n9614 VSS 0.066735f
C26578 DVDD.n9615 VSS 0.066735f
C26579 DVDD.n9616 VSS 3.31978f
C26580 DVDD.n9617 VSS 0.026274f
C26581 DVDD.n9618 VSS 0.045979f
C26582 DVDD.n9619 VSS 0.060175f
C26583 DVDD.n9620 VSS 0.026274f
C26584 DVDD.n9621 VSS 0.030088f
C26585 DVDD.n9622 VSS 0.029062f
C26586 DVDD.n9623 VSS 0.225658f
C26587 DVDD.n9624 VSS 0.066735f
C26588 DVDD.n9625 VSS 0.066735f
C26589 DVDD.n9626 VSS 0.066735f
C26590 DVDD.n9627 VSS 0.204999f
C26591 DVDD.n9628 VSS 0.029062f
C26592 DVDD.n9629 VSS 0.033368f
C26593 DVDD.n9630 VSS 0.114418f
C26594 DVDD.n9631 VSS 0.114418f
C26595 DVDD.n9632 VSS 0.15585f
C26596 DVDD.n9633 VSS 0.277706f
C26597 DVDD.n9634 VSS 0.277706f
C26598 DVDD.n9635 VSS 0.058124f
C26599 DVDD.n9636 VSS 0.114418f
C26600 DVDD.n9637 VSS 0.114418f
C26601 DVDD.n9638 VSS 0.114418f
C26602 DVDD.n9639 VSS 0.058124f
C26603 DVDD.n9640 VSS 0.058124f
C26604 DVDD.n9641 VSS 0.058124f
C26605 DVDD.n9642 VSS 0.114418f
C26606 DVDD.n9643 VSS 0.114418f
C26607 DVDD.n9644 VSS 0.114418f
C26608 DVDD.n9645 VSS 0.050859f
C26609 DVDD.n9646 VSS 0.029062f
C26610 DVDD.n9647 VSS 0.105307f
C26611 DVDD.n9648 VSS 0.091958f
C26612 DVDD.n9649 VSS 0.210614f
C26613 DVDD.n9650 VSS 0.210614f
C26614 DVDD.n9651 VSS 0.210614f
C26615 DVDD.n9652 VSS 0.210614f
C26616 DVDD.n9653 VSS 0.210614f
C26617 DVDD.n9654 VSS 0.184658f
C26618 DVDD.n9655 VSS 0.210614f
C26619 DVDD.n9656 VSS 0.210614f
C26620 DVDD.n9657 VSS 0.210614f
C26621 DVDD.n9658 VSS 0.210614f
C26622 DVDD.n9659 VSS 0.210614f
C26623 DVDD.n9660 VSS 0.210614f
C26624 DVDD.n9661 VSS 0.210614f
C26625 DVDD.n9662 VSS 0.210614f
C26626 DVDD.n9663 VSS 0.210614f
C26627 DVDD.n9664 VSS 0.210614f
C26628 DVDD.n9665 VSS 0.210614f
C26629 DVDD.n9666 VSS 0.210614f
C26630 DVDD.n9667 VSS 0.210614f
C26631 DVDD.n9668 VSS 0.210614f
C26632 DVDD.n9669 VSS 0.210614f
C26633 DVDD.n9670 VSS 0.171309f
C26634 DVDD.n9671 VSS 0.091958f
C26635 DVDD.n9672 VSS 0.105307f
C26636 DVDD.n9673 VSS 0.560793f
C26637 DVDD.n9674 VSS 0.105307f
C26638 DVDD.n9675 VSS 0.091958f
C26639 DVDD.n9676 VSS 0.210614f
C26640 DVDD.n9677 VSS 0.210614f
C26641 DVDD.n9678 VSS 0.210614f
C26642 DVDD.n9679 VSS 0.210614f
C26643 DVDD.n9680 VSS 0.210614f
C26644 DVDD.n9681 VSS 0.184658f
C26645 DVDD.n9682 VSS 0.210614f
C26646 DVDD.n9683 VSS 0.210614f
C26647 DVDD.n9684 VSS 0.210614f
C26648 DVDD.n9685 VSS 0.210614f
C26649 DVDD.n9686 VSS 0.210614f
C26650 DVDD.n9687 VSS 0.210614f
C26651 DVDD.n9688 VSS 0.210614f
C26652 DVDD.n9689 VSS 0.210614f
C26653 DVDD.n9690 VSS 0.149061f
C26654 DVDD.n9691 VSS 0.105307f
C26655 DVDD.n9692 VSS 0.013137f
C26656 DVDD.n9693 VSS 0.105307f
C26657 DVDD.n9694 VSS 0.180209f
C26658 DVDD.n9695 VSS 0.210614f
C26659 DVDD.n9696 VSS 0.189849f
C26660 DVDD.n9697 VSS 0.210614f
C26661 DVDD.n9698 VSS 0.108274f
C26662 DVDD.n9699 VSS 0.27725f
C26663 DVDD.n9700 VSS 1.01479f
.ends

