* NGSPICE file created from gf180mcu_fd_io__bi_t_pex.ext - technology: gf180mcuD

.subckt gf180mcu_fd_io__bi_t_pex DVSS DVDD PAD SL A Y PDRV1 PDRV0 PD CS OE IE PU VDD
+ VSS
X0 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t1 SL.t0 VSS.t23 VSS.t22 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
D0 CS.t0 VDD.t12 diode_pd2nw_06v0 pj=4u area=1p
X1 DVSS.t174 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t2 DVSS.t173 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t1 DVDD.t58 DVDD.t57 pfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t1 VSS.t8 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS.t0 DVDD.t26 ppolyf_u r_width=0.8u r_length=35.7u
X5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t3 VDD.t5 VDD.t4 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X6 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t2 GF_NI_BI_T_BASE_0.ndrive_x_<0>.t0 DVDD.t25 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X7 DVDD.t194 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB.t0 DVDD.t193 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X8 GF_NI_BI_T_BASE_0.ndrive_x_<0>.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t3 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t0 DVDD.t22 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X9 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t2 DVDD.t63 DVDD.t62 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X10 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS PAD.t3 w_4468_53342# ppolyf_u r_width=2.5u r_length=2.8u
X11 PAD GF_NI_BI_T_BASE_0.pdrive_y_<0>.t4 DVDD DVDD.t195 pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X12 GF_NI_BI_T_BASE_0.pdrive_y_<1>.t0 DVDD.t205 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t0 DVSS.t32 nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X13 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t3 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t4 DVSS.t5 nfet_06v0 ad=0.689p pd=3.17u as=0.689p ps=3.17u w=2.65u l=0.7u
X14 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t4 DVSS.t206 GF_NI_BI_T_BASE_0.ndrive_x_<0>.t2 DVDD.t186 pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X15 PAD GF_NI_BI_T_BASE_0.ndrive_x_<1>.t3 DVSS DVSS.t117 nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.14364n pd=83.56u as=10.639999p ps=76.56u w=38u l=1.15u
X16 DVSS.t102 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t2 DVSS.t101 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X17 DVDD.t206 DVSS.t33 cap_nmos_06v0 c_width=5u c_length=1.5u
X18 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t2 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t2 DVSS.t37 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X19 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t2 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t8 DVSS.t62 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X20 PU.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t0 VSS.t15 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X21 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t1 DVDD.t188 DVDD.t187 pfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X22 VDD.t9 PU.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t0 VDD.t8 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X23 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS PAD.t5 w_4468_53342# ppolyf_u r_width=2.5u r_length=2.8u
X24 DVSS.t127 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t0 DVSS.t126 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X25 PAD GF_NI_BI_T_BASE_0.pdrive_x_<2>.t4 DVDD DVDD.t100 pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X26 GF_NI_BI_T_BASE_0.ndrive_x_<3>.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t2 DVSS.t131 DVSS.t130 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X27 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t2 DVDD.t203 DVDD.t202 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X28 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t3 DVDD.t192 DVDD.t191 pfet_06v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X29 Y.t11 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t2 VSS.t28 VSS.t27 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
D1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS DVDD diode_pd2nw_06v0 pj=42u area=20p
X30 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t1 PDRV0.t1 VDD.t7 VDD.t6 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X31 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t3 DVDD.t157 DVDD.t156 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X32 DVSS.t203 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t3 GF_NI_BI_T_BASE_0.pdrive_y_<3>.t2 DVSS.t202 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X33 a_5575_63014.t5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t3 DVSS.t59 DVDD.t18 pfet_06v0 ad=0.836p pd=4.68u as=0.494p ps=2.42u w=1.9u l=0.7u
X34 PAD GF_NI_BI_T_BASE_0.ndrive_x_<0>.t3 DVSS DVSS.t53 nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.14364n pd=83.56u as=10.639999p ps=76.56u w=38u l=1.15u
X35 DVSS.t160 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t3 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t2 DVSS.t159 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X36 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t0 VDD.t14 VDD.t13 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X37 DVSS.t58 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t4 a_5575_63014.t4 DVDD.t17 pfet_06v0 ad=0.494p pd=2.42u as=0.836p ps=4.68u w=1.9u l=0.7u
X38 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS.t1 DVDD.t26 ppolyf_u r_width=0.8u r_length=35.7u
X39 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t4 DVDD.t16 DVDD.t15 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X40 DVDD.t120 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t0 DVDD.t119 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X41 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t2 DVDD.t147 DVDD.t146 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X42 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t2 DVDD.t163 DVDD.t162 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X43 DVSS.t77 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t2 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t3 DVSS.t76 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X44 DVDD.t56 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB.t0 DVDD.t55 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X45 DVDD.t167 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t0 DVDD.t166 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X46 PAD GF_NI_BI_T_BASE_0.pdrive_x_<3>.t4 DVDD DVDD.t176 pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X47 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t0 IE.t0 VSS.t37 VSS.t36 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X48 VDD.t27 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t3 Y.t5 VDD.t26 pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X49 Y.t4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t4 VDD.t29 VDD.t28 pfet_06v0 ad=0.91p pd=4.02u as=1.54p ps=7.88u w=3.5u l=0.7u
X50 DVDD.t207 DVSS.t34 cap_nmos_06v0 c_width=5u c_length=1.5u
X51 DVSS.t133 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t1 DVSS.t132 nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
D2 DVSS.t19 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS diode_nd2ps_06v0 pj=42u area=20p
X52 GF_NI_BI_T_BASE_0.pdrive_y_<1>.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t3 DVSS.t151 DVSS.t150 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X53 DVDD.t171 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t3 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t1 DVDD.t170 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X54 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t3 DVSS.t147 DVSS.t146 nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X55 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t2 DVDD.t110 DVDD.t109 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X56 DVDD.t42 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t3 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t0 DVDD.t41 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X57 DVSS.t158 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t1 DVSS.t157 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X58 DVSS.t166 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t0 DVSS.t165 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X59 DVSS.t189 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t4 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t3 DVSS.t188 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X60 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t5 DVSS.t191 DVSS.t190 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X61 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t3 DVDD.t128 DVDD.t127 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X62 DVDD.t112 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB.t0 DVDD.t111 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X63 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t0 DVSS.t8 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X64 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.MINUS.t0 DVDD.t26 ppolyf_u r_width=0.8u r_length=35.7u
X65 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t0 DVSS.t80 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X66 DVDD.t143 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t4 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t1 DVDD.t142 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X67 DVDD.t136 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t4 GF_NI_BI_T_BASE_0.pdrive_y_<1>.t3 DVDD.t135 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X68 VDD.t64 CS.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t0 VDD.t63 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X69 DVSS.t180 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t1 DVSS.t179 nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X70 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t6 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t2 DVDD.t182 DVSS.t196 nfet_06v0 ad=0.572p pd=3.48u as=0.572p ps=3.48u w=1.3u l=0.7u
X71 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t5 GF_NI_BI_T_BASE_0.ndrive_x_<3>.t1 DVDD.t21 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
D3 IE.t1 VDD.t36 diode_pd2nw_06v0 pj=4u area=1p
X72 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t4 DVDD.t114 DVDD.t113 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X73 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t0 OE.t3 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S.t0 VSS.t41 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X74 PAD GF_NI_BI_T_BASE_0.pdrive_y_<2>.t4 DVDD DVDD.t199 pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X75 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t3 GF_NI_BI_T_BASE_0.pdrive_y_<3>.t3 DVSS.t95 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X76 DVDD.t208 DVSS.t35 cap_nmos_06v0 c_width=5u c_length=1.5u
X77 GF_NI_BI_T_BASE_0.ndrive_x_<3>.t2 DVSS.t207 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t4 DVDD.t185 pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X78 GF_NI_BI_T_BASE_0.pdrive_y_<3>.t3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t4 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t2 DVSS.t40 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X79 DVDD.t209 DVSS.t36 cap_nmos_06v0 c_width=5u c_length=1.5u
X80 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t4 DVSS.t116 DVSS.t115 nfet_06v0 ad=1.408p pd=7.28u as=0.832p ps=3.72u w=3.2u l=0.7u
X81 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S.t1 VDD.t65 VSS.t1 VSS.t0 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X82 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t6 GF_NI_BI_T_BASE_0.ndrive_x_<2>.t0 DVDD.t19 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X83 VDD.t59 PDRV1.t1 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t0 VDD.t58 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X84 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t3 VDD.t32 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X85 DVSS.t137 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t4 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t1 DVSS.t136 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X86 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t6 DVDD.t70 DVDD.t69 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X87 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t0 OE.t4 VDD.t53 VDD.t52 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X88 VDD.t55 OE.t5 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t0 VDD.t54 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X89 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t0 A.t0 VDD.t48 VDD.t47 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X90 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t0 DVDD.t210 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t0 DVSS.t37 nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X91 DVDD.t211 DVSS.t38 cap_nmos_06v0 c_width=5u c_length=1.5u
X92 VSS.t12 PU.t3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D.t0 VSS.t11 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X93 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t0 SL.t1 VDD.t21 VDD.t20 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X94 DVSS GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t5 PAD DVSS.t50 nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.639999p pd=76.56u as=0.14364n ps=83.56u w=38u l=1.15u
X95 VDD.t11 PU.t4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t0 VDD.t10 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X96 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t3 DVSS.t110 DVSS.t109 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X97 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t3 VDD.t42 VDD.t41 pfet_06v0 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.7u
X98 DVDD GF_NI_BI_T_BASE_0.pdrive_y_<3>.t4 PAD DVDD.t64 pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X99 DVDD.t28 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t4 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t1 DVDD.t27 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X100 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t13 DVSS.t104 DVSS.t103 nfet_06v0 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.7u
X101 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.MINUS.t1 DVDD.t26 ppolyf_u r_width=0.8u r_length=35.7u
X102 DVSS.t84 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t0 DVSS.t83 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X103 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB.t3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t1 DVDD.t93 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X104 GF_NI_BI_T_BASE_0.pdrive_y_<1>.t3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t5 DVDD.t138 DVDD.t137 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X105 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t5 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t6 DVSS.t16 nfet_06v0 ad=1.166p pd=6.18u as=0.689p ps=3.17u w=2.65u l=0.7u
X106 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t7 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t1 DVSS.t18 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X107 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t5 DVDD.t30 DVDD.t29 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X108 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t0 OE.t6 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S.t0 VSS.t24 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X109 DVSS GF_NI_BI_T_BASE_0.ndrive_y_<0>.t5 PAD DVSS.t20 nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.639999p pd=76.56u as=0.14364n ps=83.56u w=38u l=1.15u
X110 DVDD.t212 DVSS.t39 cap_nmos_06v0 c_width=5u c_length=1.5u
X111 DVSS.t198 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t0 DVSS.t197 nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X112 VDD.t44 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t0 VDD.t43 pfet_06v0 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.7u
D4 VSS.t50 OE.t2 diode_pd2nw_06v0 pj=1.92u area=0.2304p
X113 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t2 DVDD.t198 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X114 DVSS.t69 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t4 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t1 DVSS.t68 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X115 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t3 DVSS.t73 DVSS.t72 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X116 DVDD.t60 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVDD.t59 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X117 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t5 DVSS.t67 DVSS.t66 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X118 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t0 DVSS.t138 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X119 DVDD.t54 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t1 DVDD.t53 pfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X120 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t11 DVDD.t141 pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X121 DVSS.t178 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t1 DVSS.t177 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X122 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t5 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t4 DVSS.t17 nfet_06v0 ad=0.689p pd=3.17u as=1.166p ps=6.18u w=2.65u l=0.7u
X123 VDD.t31 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t5 Y.t3 VDD.t30 pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X124 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_2.PLUS.t1 DVDD.t26 ppolyf_u r_width=0.8u r_length=35.7u
X125 VSS.t14 PU.t5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t1 VSS.t13 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X126 DVSS.t182 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN DVSS.t181 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X127 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t5 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t2 DVSS.t98 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X128 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<1>.t4 PAD DVDD.t85 pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X129 GF_NI_BI_T_BASE_0.ndrive_x_<1>.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t7 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t1 DVDD.t20 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X130 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t5 DVSS.t7 DVSS.t6 nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X131 VSS.t26 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t6 Y.t10 VSS.t25 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X132 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t3 DVSS.t135 DVSS.t134 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X133 Y.t9 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t7 VSS.t19 VSS.t18 nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X134 DVDD.t149 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t1 DVDD.t148 pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X135 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S DVSS.t199 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X136 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t4 DVSS.t172 DVSS.t171 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X137 GF_NI_BI_T_BASE_0.pdrive_y_<3>.t0 DVDD.t213 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t0 DVSS.t40 nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X138 DVSS.t153 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t6 GF_NI_BI_T_BASE_0.pdrive_y_<1>.t2 DVSS.t152 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X139 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t6 DVDD.t40 DVDD.t39 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X140 DVDD.t214 DVSS.t41 cap_nmos_06v0 c_width=3u c_length=3u
X141 DVSS.t57 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t8 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t1 DVSS.t56 nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X142 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t4 DVSS.t129 DVSS.t128 nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X143 VDD.t16 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t8 Y.t2 VDD.t15 pfet_06v0 ad=1.54p pd=7.88u as=0.91p ps=4.02u w=3.5u l=0.7u
X144 PAD GF_NI_BI_T_BASE_0.ndrive_x_<2>.t3 DVSS DVSS.t141 nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.14364n pd=83.56u as=10.639999p ps=76.56u w=38u l=1.15u
X145 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t6 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t3 DVSS.t44 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X146 DVDD.t130 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t0 DVDD.t129 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X147 DVDD.t13 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t1 DVDD.t12 pfet_06v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X148 a_5575_63014.t1 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t6 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t10 DVDD.t2 pfet_06v0 ad=0.946p pd=5.18u as=0.559p ps=2.67u w=2.15u l=0.7u
X149 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t4 DVDD.t134 DVDD.t133 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
D5 VSS.t51 VDD.t60 diode_pd2nw_06v0 pj=1.92u area=0.2304p
X150 GF_NI_BI_T_BASE_0.ndrive_x_<2>.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t9 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t0 DVDD.t14 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X151 VSS.t5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t1 VSS.t4 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
D6 VSS.t52 OE.t1 diode_pd2nw_06v0 pj=1.92u area=0.2304p
X152 DVDD.t140 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t6 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t0 DVDD.t139 pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X153 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t4 DVSS.t208 GF_NI_BI_T_BASE_0.ndrive_x_<2>.t2 DVDD.t184 pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X154 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_2.PLUS.t0 DVDD.t61 ppolyf_u r_width=0.8u r_length=22.999998u
X155 DVDD.t68 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t0 DVDD.t67 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X156 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t7 DVDD.t72 DVDD.t71 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X157 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t1 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t3 DVSS.t82 DVSS.t81 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X158 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t1 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t3 DVSS.t176 DVSS.t175 nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X159 DVSS.t140 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t2 GF_NI_BI_T_BASE_0.ndrive_x_<0>.t1 DVSS.t139 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X160 Y.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t9 VDD.t18 VDD.t17 pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X161 DVDD.t215 DVSS.t42 cap_nmos_06v0 c_width=3u c_length=3u
X162 DVDD.t155 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t1 DVDD.t154 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X163 DVSS.t30 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t6 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t1 DVSS.t29 nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X164 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t0 PD.t0 VDD.t57 VDD.t56 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X165 GF_NI_BI_T_BASE_0.pdrive_y_<3>.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t6 DVSS.t65 DVSS.t64 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
D7 A.t1 VDD.t19 diode_pd2nw_06v0 pj=4u area=1p
X166 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t7 GF_NI_BI_T_BASE_0.pdrive_y_<1>.t1 DVSS.t99 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X167 DVDD.t38 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t7 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t0 DVDD.t37 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X168 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t7 DVSS.t28 DVSS.t27 nfet_06v0 ad=0.832p pd=3.72u as=1.408p ps=7.28u w=3.2u l=0.7u
X169 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t3 DVSS.t201 DVSS.t200 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X170 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<0>.t4 PAD DVDD.t79 pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X171 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t1 IE.t2 VDD.t46 VDD.t45 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X172 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_4.PLUS.t1 DVDD.t26 ppolyf_u r_width=0.8u r_length=35.7u
X173 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t0 PD.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t2 VSS.t42 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X174 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t3 DVDD.t190 DVDD.t189 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X175 DVDD.t32 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t7 GF_NI_BI_T_BASE_0.pdrive_y_<3>.t1 DVDD.t31 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X176 VDD.t23 OE.t7 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t1 VDD.t22 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X177 PAD GF_NI_BI_T_BASE_0.pdrive_x_<1>.t5 DVDD DVDD.t88 pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X178 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t1 VDD.t49 VDD.t51 VDD.t50 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X179 DVSS.t162 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t5 GF_NI_BI_T_BASE_0.ndrive_x_<3>.t0 DVSS.t161 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X180 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t6 DVSS.t10 DVSS.t9 nfet_06v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X181 DVSS GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t5 PAD DVSS.t92 nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.639999p pd=76.56u as=0.14364n ps=83.56u w=38u l=1.15u
X182 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t2 DVSS.t97 DVSS.t96 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
D8 VSS.t53 OE.t0 diode_pd2nw_06v0 pj=1.92u area=0.2304p
X183 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t3 DVDD.t126 DVDD.t125 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X184 DVDD.t169 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVDD.t168 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X185 DVSS.t195 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t2 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t1 DVSS.t194 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X186 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t7 DVDD.t52 DVDD.t51 pfet_06v0 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.7u
D9 SL.t2 VDD.t19 diode_pd2nw_06v0 pj=4u area=1p
X187 DVDD.t216 DVSS.t43 cap_nmos_06v0 c_width=3u c_length=3u
X188 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t1 VSS.t17 VSS.t16 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X189 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t8 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t4 DVSS.t15 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X190 DVSS.t106 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t14 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t1 DVSS.t105 nfet_06v0 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.7u
X191 DVDD.t165 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t0 DVDD.t164 pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X192 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t1 DVDD.t217 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t2 DVSS.t44 nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X193 DVDD.t122 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t7 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t3 DVDD.t121 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X194 DVDD.t218 DVSS.t45 cap_nmos_06v0 c_width=5u c_length=1.5u
X195 a_5575_63014.t3 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t7 DVDD.t11 DVDD.t10 pfet_06v0 ad=0.836p pd=4.68u as=0.494p ps=2.42u w=1.9u l=0.7u
X196 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S.t1 PDRV0.t2 VSS.t10 VSS.t9 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X197 VSS.t21 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t10 Y.t8 VSS.t20 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X198 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t5 VDD.t38 VDD.t37 pfet_06v0 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.7u
X199 DVSS GF_NI_BI_T_BASE_0.ndrive_y_<2>.t5 PAD DVSS.t87 nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.639999p pd=76.56u as=0.14364n ps=83.56u w=38u l=1.15u
X200 DVDD GF_NI_BI_T_BASE_0.pdrive_y_<1>.t4 PAD DVDD.t106 pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X201 GF_NI_BI_T_BASE_0.ndrive_x_<1>.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t4 DVSS.t112 DVSS.t111 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X202 DVDD.t24 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t8 a_5575_63014.t2 DVDD.t23 pfet_06v0 ad=0.494p pd=2.42u as=0.836p ps=4.68u w=1.9u l=0.7u
X203 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t6 DVSS.t164 DVSS.t163 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X204 DVSS.t114 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t5 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t3 DVSS.t113 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X205 VDD.t40 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t6 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t0 VDD.t39 pfet_06v0 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.7u
X206 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t2 DVSS.t145 DVSS.t144 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X207 DVDD.t161 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t0 DVDD.t160 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X208 GF_NI_BI_T_BASE_0.pdrive_y_<3>.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t8 DVDD.t34 DVDD.t33 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
D10 PU.t6 VDD.t12 diode_pd2nw_06v0 pj=4u area=1p
X209 VSS.t7 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D.t1 VSS.t6 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X210 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t9 DVDD.t50 DVDD.t49 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X211 DVSS.t61 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t8 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB.t1 DVSS.t60 nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X212 PU.t0 PD.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t1 VDD.t33 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X213 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t7 DVDD.t97 DVDD.t96 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X214 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t9 DVSS.t24 DVSS.t23 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X215 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t5 DVDD.t173 DVDD.t172 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X216 GF_NI_BI_T_BASE_0.ndrive_x_<0>.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t4 DVSS.t149 DVSS.t148 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X217 DVSS.t75 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t4 GF_NI_BI_T_BASE_0.ndrive_x_<2>.t1 DVSS.t74 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X218 VSS.t31 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t11 Y.t7 VSS.t30 nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X219 VDD.t3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.Z VDD.t2 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X220 VDD.t25 OE.t8 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t1 VDD.t24 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X221 DVDD.t219 DVSS.t46 cap_nmos_06v0 c_width=5u c_length=1.5u
X222 DVDD.t220 DVSS.t47 cap_nmos_06v0 c_width=3u c_length=3u
X223 VSS.t3 CS.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t1 VSS.t2 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X224 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS PAD.t4 w_4468_53342# ppolyf_u r_width=2.5u r_length=2.8u
X225 DVDD.t5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t10 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t0 DVDD.t4 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X226 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t5 DVDD.t78 DVDD.t77 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X227 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t3 DVSS.t86 DVSS.t85 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X228 VSS.t35 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t7 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t1 VSS.t34 nfet_06v0 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.7u
X229 PAD GF_NI_BI_T_BASE_0.ndrive_x_<3>.t3 DVSS DVSS.t185 nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.14364n pd=83.56u as=10.639999p ps=76.56u w=38u l=1.15u
X230 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<3>.t5 PAD DVDD.t179 pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X231 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t8 VSS.t47 VSS.t46 nfet_06v0 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.7u
X232 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t4 DVDD.t118 DVDD.t117 pfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X233 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t7 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S DVSS.t156 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X234 DVDD.t74 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t8 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t1 DVDD.t73 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X235 DVSS.t170 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t6 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t1 DVSS.t169 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X236 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t1 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t9 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t6 DVSS.t63 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X237 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_4.PLUS.t0 DVDD.t26 ppolyf_u r_width=0.8u r_length=35.7u
X238 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t11 DVSS.t2 DVSS.t1 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X239 DVDD.t99 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t6 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t0 DVDD.t98 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X240 DVDD.t221 DVSS.t48 cap_nmos_06v0 c_width=5u c_length=1.5u
X241 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t5 DVSS.t184 DVSS.t183 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X242 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t5 DVSS.t79 DVSS.t78 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X243 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t5 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t10 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t0 DVSS.t31 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
D11 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS DVDD diode_pd2nw_06v0 pj=42u area=20p
X244 GF_NI_BI_T_BASE_0.ndrive_x_<3>.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t12 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t3 DVDD.t0 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X245 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t8 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t2 DVSS.t100 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X246 DVDD.t222 DVSS.t49 cap_nmos_06v0 c_width=5u c_length=1.5u
X247 Y.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t12 VDD.t35 VDD.t34 pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X248 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t4 DVSS.t91 DVSS.t90 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X249 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t13 GF_NI_BI_T_BASE_0.ndrive_x_<1>.t1 DVDD.t1 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X250 DVSS.t14 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t10 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB.t1 DVSS.t13 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X251 DVSS.t155 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t1 DVSS.t154 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X252 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t10 DVDD.t9 DVDD.t8 pfet_06v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X253 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t9 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t11 a_5575_63014.t0 DVDD.t3 pfet_06v0 ad=0.559p pd=2.67u as=0.946p ps=5.18u w=2.15u l=0.7u
X254 Y.t6 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t13 VSS.t33 VSS.t32 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X255 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t1 DVDD.t75 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X256 GF_NI_BI_T_BASE_0.pdrive_y_<1>.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t9 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t2 DVSS.t32 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X257 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t7 DVSS.t168 DVSS.t167 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X258 GF_NI_BI_T_BASE_0.ndrive_x_<1>.t2 DVSS.t209 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t4 DVDD.t183 pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X259 VSS.t44 PDRV1.t2 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S.t0 VSS.t43 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X260 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t0 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t5 DVDD.t159 DVDD.t158 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X261 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t5 DVDD.t46 DVDD.t45 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X262 DVDD.t116 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t5 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t3 DVDD.t115 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X263 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D.t0 PD.t3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.Z VSS.t29 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X264 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S.t1 OE.t9 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t1 VSS.t38 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X265 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t15 DVDD.t95 DVDD.t94 pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X266 VSS.t40 OE.t10 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S.t1 VSS.t39 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
D12 DVSS.t19 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS diode_nd2ps_06v0 pj=42u area=20p
X267 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S.t0 A.t2 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t1 VSS.t45 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X268 GF_NI_BI_T_BASE_0.ndrive_x_<2>.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t6 DVSS.t71 DVSS.t70 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X269 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.Z PD.t4 VDD.t62 VDD.t61 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X270 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<2>.t5 PAD DVDD.t103 pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X271 DVSS.t123 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB.t1 DVSS.t122 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
D13 VSS.t54 PDRV1.t0 diode_pd2nw_06v0 pj=1.92u area=0.2304p
X272 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t0 PD.t5 VSS.t49 VSS.t48 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X273 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS PAD.t21 w_4468_53342# ppolyf_u r_width=2.5u r_length=2.8u
X274 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t1 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t3 DVDD.t92 DVDD.t91 pfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X275 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t8 DVDD.t153 DVDD.t152 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X276 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t6 DVSS.t125 DVSS.t124 nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X277 DVDD.t175 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t3 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t0 DVDD.t174 pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X278 DVDD.t145 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t0 DVDD.t144 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X279 DVSS.t12 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t11 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t1 DVSS.t11 nfet_06v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X280 PAD GF_NI_BI_T_BASE_0.pdrive_x_<0>.t5 DVDD DVDD.t82 pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X281 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t8 DVDD.t36 DVDD.t35 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X282 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t12 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t2 DVDD.t204 pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X283 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t2 DVSS.t108 DVSS.t107 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X284 DVSS.t121 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t6 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t2 DVSS.t120 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X285 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t3 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t12 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t3 DVSS.t0 nfet_06v0 ad=0.689p pd=3.17u as=0.689p ps=3.17u w=2.65u l=0.7u
X286 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t7 DVSS.t193 DVSS.t192 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X287 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t1 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t0 DVDD.t76 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X288 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t8 DVDD.t124 DVDD.t123 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
D14 PD.t6 VDD.t36 diode_pd2nw_06v0 pj=4u area=1p
X289 VDD.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t0 VDD.t0 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X290 DVDD.t151 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t9 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t0 DVDD.t150 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X291 DVSS.t26 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t11 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t0 DVSS.t25 nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X292 DVDD.t48 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t12 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t0 DVDD.t47 pfet_06v0 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.7u
X293 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t12 DVSS.t4 DVSS.t3 nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
D15 VSS.t55 PDRV0.t0 diode_pd2nw_06v0 pj=1.92u area=0.2304p
X294 DVDD.t44 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t7 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t2 DVDD.t43 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X295 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t1 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t3 DVDD.t132 DVDD.t131 pfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X296 DVSS.t205 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t7 GF_NI_BI_T_BASE_0.ndrive_x_<1>.t0 DVSS.t204 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
R0 SL.n2 SL.t1 43.0184
R1 SL.n2 SL.t0 30.9212
R2 SL.n1 SL 27.184
R3 SL SL.n1 4.56015
R4 SL SL.n2 4.00158
R5 SL.n1 SL.n0 3.59134
R6 SL SL.t2 2.6293
R7 SL.n0 SL.t2 2.60635
R8 SL.n0 SL 0.02345
R9 VSS.n2636 VSS.n2617 196056
R10 VSS.n5290 VSS.n5289 37210.9
R11 VSS.n5711 VSS.n11 32548.6
R12 VSS.n5449 VSS.n5448 32385.4
R13 VSS.n2635 VSS.n2203 30893.3
R14 VSS.n5691 VSS.n5690 27088.7
R15 VSS.n5454 VSS.n1290 25861.7
R16 VSS.n4204 VSS.n2617 21519.5
R17 VSS.n5690 VSS.n5689 20471.6
R18 VSS.n5294 VSS.n2200 19823.1
R19 VSS.n5455 VSS.n5454 19552.7
R20 VSS.n5304 VSS.n5303 17654
R21 VSS.n5710 VSS.n12 16516.8
R22 VSS.n2080 VSS.n1292 16516.8
R23 VSS.n5304 VSS.n2187 16432
R24 VSS.n4326 VSS.n2203 16400
R25 VSS.n4327 VSS.n4325 16252.3
R26 VSS.n5691 VSS.n12 16242.7
R27 VSS.n1292 VSS.n1290 16242.7
R28 VSS.n5317 VSS.n2187 16230.9
R29 VSS.n5291 VSS.n2202 16230.9
R30 VSS.n5305 VSS.n5304 16230.9
R31 VSS.n5303 VSS.n2099 16230.9
R32 VSS.n5435 VSS.n2091 16230.9
R33 VSS.n4199 VSS.n2635 15030.2
R34 VSS.n4199 VSS.n2634 14984.7
R35 VSS.n4327 VSS.n4326 14824
R36 VSS.n5294 VSS.n5293 14824
R37 VSS.n5692 VSS.n5691 14769.2
R38 VSS.n1290 VSS.n1172 14767.1
R39 VSS.n5289 VSS.n2203 13915.8
R40 VSS.n4868 VSS.n4866 12369.1
R41 VSS.n3620 VSS.n2410 12369.1
R42 VSS.n3246 VSS.n2704 12369.1
R43 VSS.n3248 VSS.n3247 12369.1
R44 VSS.n5293 VSS.n5292 11473.2
R45 VSS.n5292 VSS.n5291 10835.5
R46 VSS.n5290 VSS.n2178 9379.2
R47 VSS.n4867 VSS.n2237 8636.96
R48 VSS.n5291 VSS.n5290 8547.5
R49 VSS.n3602 VSS.n2635 7940.47
R50 VSS.n5448 VSS.n2081 7811.82
R51 VSS.n4204 VSS.n4203 7328.63
R52 VSS.n5177 VSS.n2223 6939.76
R53 VSS.n4325 VSS.n4324 6651.3
R54 VSS.n5302 VSS.n5301 6538.35
R55 VSS.n3247 VSS.n3246 6519.88
R56 VSS.n4869 VSS.n4868 6104.43
R57 VSS.n5289 VSS.n5288 5387.7
R58 VSS.n5318 VSS.n2186 4902.86
R59 VSS.n5346 VSS.n2177 4902.86
R60 VSS.n2193 VSS.n2105 4902.86
R61 VSS.n5302 VSS.n2091 4526.71
R62 VSS.n2797 VSS.n2634 4493.06
R63 VSS.n5266 VSS.n2237 3620.98
R64 VSS.n4325 VSS.n2617 3491.91
R65 VSS.n5293 VSS.n2201 3437.85
R66 VSS.n4326 VSS.n2201 3435.27
R67 VSS.n4127 VSS.n3777 3354.59
R68 VSS.n4127 VSS.n3779 3354.59
R69 VSS.n5303 VSS.n5302 3311.99
R70 VSS.n4205 VSS.n4204 3307.91
R71 VSS.n3247 VSS.n2797 3136.7
R72 VSS.n4324 VSS.n2200 3086.59
R73 VSS.n5345 VSS.n2178 2875.76
R74 VSS.n4670 VSS.n2510 2717.55
R75 VSS.n4670 VSS.n2511 2717.55
R76 VSS.n5332 VSS.n5331 2717.55
R77 VSS.n5331 VSS.n2185 2717.55
R78 VSS.n4868 VSS.n4867 2581.97
R79 VSS.n5712 VSS.n9 2402.48
R80 VSS.n5712 VSS.n10 2401.2
R81 VSS.n5450 VSS.n9 2400.01
R82 VSS.n5450 VSS.n10 2398.73
R83 VSS.n3246 VSS.n3245 2395.26
R84 VSS.n1744 VSS.n13 2286.22
R85 VSS.n1742 VSS.n1729 2282.35
R86 VSS.n1743 VSS.n1742 2282.35
R87 VSS.n1729 VSS.n1293 2278.48
R88 VSS.n1744 VSS.n1743 2277.19
R89 VSS.n4208 VSS.n2091 2219.8
R90 VSS.n5709 VSS.n13 2185.59
R91 VSS.n2079 VSS.n1293 2179.14
R92 VSS.n5292 VSS.n2187 2099.5
R93 VSS.n5344 VSS.n11 1924.39
R94 VSS.n4325 VSS.n4323 1819.86
R95 VSS.n909 VSS.n220 1814.99
R96 VSS.n910 VSS.n909 1813.28
R97 VSS.n3245 VSS.n2410 1508.72
R98 VSS.n5328 VSS.n5327 1449.32
R99 VSS.n5406 VSS.n2111 1375
R100 VSS.n5327 VSS.n5319 1235.04
R101 VSS.n5327 VSS.n5320 1235.04
R102 VSS.n4198 VSS.n4194 1219.32
R103 VSS.n4203 VSS.t13 1116.18
R104 VSS.n5178 VSS.n2274 1105.19
R105 VSS.n5416 VSS.n2104 1089.54
R106 VSS.t48 VSS.n4198 1038.26
R107 VSS.n5178 VSS.n5177 1024.12
R108 VSS.n2080 VSS.n2079 967.646
R109 VSS.n5710 VSS.n5709 967.646
R110 VSS.t15 VSS.t13 953.457
R111 VSS.t0 VSS.n2111 882.342
R112 VSS.t43 VSS.n2111 882.342
R113 VSS.n4205 VSS.n2630 835.686
R114 VSS.n4867 VSS.n2274 826.212
R115 VSS.n5331 VSS.n2186 815.005
R116 VSS.n5407 VSS.n5406 800.532
R117 VSS.t41 VSS.n5306 798.532
R118 VSS.n5316 VSS.t38 798.532
R119 VSS.n4843 VSS.t24 797.183
R120 VSS.n4199 VSS.t48 744.888
R121 VSS.n5405 VSS.n2112 709.234
R122 VSS.n5347 VSS.n2176 709.234
R123 VSS.n5306 VSS.n5305 693.769
R124 VSS.n5317 VSS.n5316 693.769
R125 VSS.n4843 VSS.n2202 693.769
R126 VSS.n5407 VSS.n2105 676.944
R127 VSS.n3622 VSS.n3621 675.573
R128 VSS.n3622 VSS.n2239 675.573
R129 VSS.n5262 VSS.n2240 675.573
R130 VSS.n5416 VSS.n5415 651.337
R131 VSS.n4850 VSS.t9 640.203
R132 VSS.n5331 VSS.n5328 626.841
R133 VSS.n5328 VSS.n2176 614.595
R134 VSS.n4194 VSS.n2636 614.245
R135 VSS.n5449 VSS.n2080 608.972
R136 VSS.n5711 VSS.n5710 608.972
R137 VSS.n5345 VSS.n5344 588.939
R138 VSS.n4871 VSS.n2408 586.833
R139 VSS.n5346 VSS.n5345 578.966
R140 VSS.n3256 VSS.n2634 562.811
R141 VSS.n5319 VSS.n5318 549.35
R142 VSS.n5320 VSS.n2177 549.35
R143 VSS.n2193 VSS.n2104 547.1
R144 VSS.n3244 VSS.n2408 517.379
R145 VSS.n4200 VSS.t42 515.692
R146 VSS.n2510 VSS.n2093 488.243
R147 VSS.n2511 VSS.n2097 488.243
R148 VSS.n5332 VSS.n2182 488.243
R149 VSS.n2185 VSS.n2179 488.243
R150 VSS.n3244 VSS.n2273 478.878
R151 VSS.n3521 VSS.n2725 472.197
R152 VSS.n4871 VSS.n2409 447.923
R153 VSS.n4200 VSS.t15 437.764
R154 VSS.n2186 VSS.n2112 426.43
R155 VSS.n3520 VSS.n2707 396.685
R156 VSS.n5447 VSS.n2082 393.92
R157 VSS.n2090 VSS.n2089 388.551
R158 VSS.t8 VSS.n2627 363.911
R159 VSS.n2627 VSS.t6 363.911
R160 VSS.n5263 VSS.n5262 360.44
R161 VSS.n5423 VSS.n5422 355.668
R162 VSS.n3619 VSS.n2697 344.332
R163 VSS.n4865 VSS.n2411 344.332
R164 VSS.n3255 VSS.t4 343.325
R165 VSS.n3612 VSS.t16 343.325
R166 VSS.n3612 VSS.t2 343.325
R167 VSS.n4858 VSS.t36 343.325
R168 VSS.n5406 VSS.n5405 341.812
R169 VSS.n2730 VSS.t34 334.264
R170 VSS.t18 VSS.n2730 330.236
R171 VSS.n5307 VSS.t41 325.932
R172 VSS.n5312 VSS.t38 325.932
R173 VSS.n5425 VSS.n2100 325.471
R174 VSS.n5263 VSS.n2239 315.134
R175 VSS.n5422 VSS.n2102 302.654
R176 VSS.n3608 VSS.n2704 300.031
R177 VSS.n3620 VSS.n3619 300.031
R178 VSS.n3621 VSS.n3620 300.031
R179 VSS.n4866 VSS.n2240 300.031
R180 VSS.n4866 VSS.n4865 300.031
R181 VSS.n5440 VSS.n2090 299.969
R182 VSS.n5265 VSS.n5264 290.733
R183 VSS.n3601 VSS.n2707 278.889
R184 VSS.n4208 VSS.n2081 271
R185 VSS.n4870 VSS.n2410 266.361
R186 VSS.n4206 VSS.n4205 255.427
R187 VSS.t27 VSS.t30 245.663
R188 VSS.t34 VSS.t46 245.663
R189 VSS.n5307 VSS.t0 242.12
R190 VSS.n5312 VSS.t43 242.12
R191 VSS.n4849 VSS.t24 236.487
R192 VSS.n3840 VSS.n3777 233.749
R193 VSS.n4069 VSS.n3779 233.749
R194 VSS.t22 VSS.n2092 229.507
R195 VSS.n2520 VSS.t22 229.507
R196 VSS.n3607 VSS.n2703 227.541
R197 VSS.n2200 VSS.n2195 224.798
R198 VSS.n5267 VSS.n5266 219.064
R199 VSS.t45 VSS.n2509 212.731
R200 VSS.t42 VSS.n4199 208.569
R201 VSS.n3249 VSS.t20 208.411
R202 VSS.n3521 VSS.n3520 203.377
R203 VSS.n5439 VSS.n5435 199.98
R204 VSS.n2509 VSS.n2099 199.98
R205 VSS.n3603 VSS.n3602 197.337
R206 VSS.n2797 VSS.n2408 187.429
R207 VSS.n4850 VSS.n2178 185.811
R208 VSS.n5440 VSS.n5439 181.861
R209 VSS.t9 VSS.n4849 175.677
R210 VSS.n2637 VSS.n2636 170.571
R211 VSS.t11 VSS.n4214 162.298
R212 VSS.n5434 VSS.n2092 154.346
R213 VSS.n3248 VSS.t32 154.043
R214 VSS.n5450 VSS.n5449 152.252
R215 VSS.n5712 VSS.n5711 152.252
R216 VSS.n4308 VSS.t29 150.202
R217 VSS.n4870 VSS.n4869 149.083
R218 VSS.t25 VSS.n3531 149.01
R219 VSS.n5305 VSS.n2193 146.669
R220 VSS.n5318 VSS.n5317 146.669
R221 VSS.n2202 VSS.n2177 146.669
R222 VSS.n3532 VSS.t32 145.988
R223 VSS.n4214 VSS.n2081 137.097
R224 VSS.n4670 VSS.n2520 134.886
R225 VSS.n5415 VSS.n2105 131.381
R226 VSS.n5433 VSS.n2083 129.345
R227 VSS.n5342 VSS.n5339 129.345
R228 VSS.n5427 VSS.n2098 129.345
R229 VSS.n5408 VSS.n2110 129.345
R230 VSS.n5446 VSS.n2083 128.957
R231 VSS.n5343 VSS.n5342 128.957
R232 VSS.n4215 VSS.t11 122.984
R233 VSS.n4215 VSS.t8 122.984
R234 VSS.t29 VSS.n4306 122.984
R235 VSS.n5347 VSS.n5346 118.02
R236 VSS.n4308 VSS.n4307 114.919
R237 VSS.n4315 VSS.n4314 114.919
R238 VSS.n4316 VSS.n4315 114.919
R239 VSS.n4316 VSS.n2618 114.919
R240 VSS.n4322 VSS.n2618 114.919
R241 VSS.n5300 VSS.n2195 114.919
R242 VSS.n5301 VSS.n2194 112.903
R243 VSS.n4323 VSS.n4322 111.895
R244 VSS.n5179 VSS.n2273 110.056
R245 VSS.t6 VSS.n2625 108.871
R246 VSS.n5268 VSS.n5267 102.416
R247 VSS.n4669 VSS.n2523 102.356
R248 VSS.n5330 VSS.n2183 102.356
R249 VSS.n5426 VSS.n5425 102.004
R250 VSS.n5693 VSS.n15 99.728
R251 VSS.n1294 VSS.n1171 99.7229
R252 VSS.n3532 VSS.t25 99.6752
R253 VSS.n4307 VSS.n2622 98.7908
R254 VSS.n5426 VSS.n2099 97.977
R255 VSS.n3531 VSS.t18 96.6548
R256 VSS.t46 VSS.n2725 95.648
R257 VSS.n2089 VSS.n2082 93.2795
R258 VSS.t20 VSS.n3248 91.6207
R259 VSS.n3608 VSS.n3607 90.6139
R260 VSS.n910 VSS.n219 86.0408
R261 VSS.n4671 VSS.t39 83.8845
R262 VSS.n3603 VSS.n2704 82.5594
R263 VSS.n4858 VSS.n2237 81.5525
R264 VSS.n220 VSS.n219 80.8661
R265 VSS.n4671 VSS.t45 79.858
R266 VSS.t39 VSS.n4670 73.8184
R267 VSS.n4128 VSS.n3775 73.4718
R268 VSS.n4128 VSS.n3776 73.4718
R269 VSS.n3884 VSS.n3778 73.2997
R270 VSS.n3785 VSS.n3778 73.2997
R271 VSS.n5414 VSS.n2106 72.4894
R272 VSS.n2078 VSS.n1294 69.3341
R273 VSS.n5708 VSS.n15 69.3341
R274 VSS.n2630 VSS.n2081 64.5166
R275 VSS.t30 VSS.n2796 61.4162
R276 VSS.n5333 VSS.n2183 61.1338
R277 VSS.n2184 VSS.n2183 61.1338
R278 VSS.n2523 VSS.n2521 61.1338
R279 VSS.n2523 VSS.n2522 61.1338
R280 VSS.n2519 VSS.n2512 59.6561
R281 VSS.n4859 VSS.n2412 59.6561
R282 VSS.n3254 VSS.n2795 59.6561
R283 VSS.n908 VSS.n219 58.4662
R284 VSS.n2106 VSS.n2098 56.4672
R285 VSS.n5408 VSS.n2106 56.4672
R286 VSS.n4864 VSS.n2412 56.0005
R287 VSS.n3618 VSS.n2698 56.0005
R288 VSS.n3250 VSS.n2795 56.0005
R289 VSS.n4192 VSS.n2637 55.8444
R290 VSS.n5417 VSS.n2102 53.0152
R291 VSS.n5435 VSS.n5434 45.6334
R292 VSS.n5417 VSS.n5416 41.6069
R293 VSS.n5433 VSS.n2093 40.8338
R294 VSS.n5339 VSS.n2179 40.8338
R295 VSS.n2182 VSS.n2110 40.8338
R296 VSS.n5427 VSS.n2097 40.8338
R297 VSS.n4126 VSS.n3780 40.2769
R298 VSS.n4126 VSS.n3781 40.2769
R299 VSS.n5267 VSS.n2224 39.6013
R300 VSS.n2409 VSS.n2273 38.5005
R301 VSS.n3256 VSS.n3255 37.2527
R302 VSS.n3249 VSS.t27 37.2527
R303 VSS.n3613 VSS.n2702 33.0561
R304 VSS.n5423 VSS.n2100 30.1987
R305 VSS.n5457 VSS.n5456 29.2479
R306 VSS.n5457 VSS.n1285 29.2479
R307 VSS.n5463 VSS.n1285 29.2479
R308 VSS.n5464 VSS.n5463 29.2479
R309 VSS.n5465 VSS.n5464 29.2479
R310 VSS.n5465 VSS.n1281 29.2479
R311 VSS.n5471 VSS.n1281 29.2479
R312 VSS.n5472 VSS.n5471 29.2479
R313 VSS.n5473 VSS.n5472 29.2479
R314 VSS.n5473 VSS.n1277 29.2479
R315 VSS.n5479 VSS.n1277 29.2479
R316 VSS.n5480 VSS.n5479 29.2479
R317 VSS.n5481 VSS.n5480 29.2479
R318 VSS.n5481 VSS.n1273 29.2479
R319 VSS.n5487 VSS.n1273 29.2479
R320 VSS.n5488 VSS.n5487 29.2479
R321 VSS.n5489 VSS.n5488 29.2479
R322 VSS.n5489 VSS.n1269 29.2479
R323 VSS.n5495 VSS.n1269 29.2479
R324 VSS.n5496 VSS.n5495 29.2479
R325 VSS.n5497 VSS.n5496 29.2479
R326 VSS.n5497 VSS.n1265 29.2479
R327 VSS.n5503 VSS.n1265 29.2479
R328 VSS.n5504 VSS.n5503 29.2479
R329 VSS.n5505 VSS.n5504 29.2479
R330 VSS.n5505 VSS.n1261 29.2479
R331 VSS.n5511 VSS.n1261 29.2479
R332 VSS.n5512 VSS.n5511 29.2479
R333 VSS.n5513 VSS.n5512 29.2479
R334 VSS.n5513 VSS.n1257 29.2479
R335 VSS.n5519 VSS.n1257 29.2479
R336 VSS.n5520 VSS.n5519 29.2479
R337 VSS.n5521 VSS.n5520 29.2479
R338 VSS.n5521 VSS.n1253 29.2479
R339 VSS.n5527 VSS.n1253 29.2479
R340 VSS.n5528 VSS.n5527 29.2479
R341 VSS.n5529 VSS.n5528 29.2479
R342 VSS.n5529 VSS.n1249 29.2479
R343 VSS.n5535 VSS.n1249 29.2479
R344 VSS.n5536 VSS.n5535 29.2479
R345 VSS.n5537 VSS.n5536 29.2479
R346 VSS.n5537 VSS.n1245 29.2479
R347 VSS.n5543 VSS.n1245 29.2479
R348 VSS.n5544 VSS.n5543 29.2479
R349 VSS.n5545 VSS.n5544 29.2479
R350 VSS.n5545 VSS.n1241 29.2479
R351 VSS.n5551 VSS.n1241 29.2479
R352 VSS.n5552 VSS.n5551 29.2479
R353 VSS.n5553 VSS.n5552 29.2479
R354 VSS.n5553 VSS.n1237 29.2479
R355 VSS.n5559 VSS.n1237 29.2479
R356 VSS.n5560 VSS.n5559 29.2479
R357 VSS.n5561 VSS.n5560 29.2479
R358 VSS.n5561 VSS.n1233 29.2479
R359 VSS.n5568 VSS.n1233 29.2479
R360 VSS.n5569 VSS.n5568 29.2479
R361 VSS.n5571 VSS.n1229 29.2479
R362 VSS.n5577 VSS.n1229 29.2479
R363 VSS.n5578 VSS.n5577 29.2479
R364 VSS.n5579 VSS.n5578 29.2479
R365 VSS.n5579 VSS.n1225 29.2479
R366 VSS.n5585 VSS.n1225 29.2479
R367 VSS.n5586 VSS.n5585 29.2479
R368 VSS.n5587 VSS.n5586 29.2479
R369 VSS.n5587 VSS.n1221 29.2479
R370 VSS.n5593 VSS.n1221 29.2479
R371 VSS.n5594 VSS.n5593 29.2479
R372 VSS.n5595 VSS.n5594 29.2479
R373 VSS.n5595 VSS.n1217 29.2479
R374 VSS.n5601 VSS.n1217 29.2479
R375 VSS.n5602 VSS.n5601 29.2479
R376 VSS.n5603 VSS.n5602 29.2479
R377 VSS.n5603 VSS.n1213 29.2479
R378 VSS.n5609 VSS.n1213 29.2479
R379 VSS.n5610 VSS.n5609 29.2479
R380 VSS.n5611 VSS.n5610 29.2479
R381 VSS.n5611 VSS.n1209 29.2479
R382 VSS.n5617 VSS.n1209 29.2479
R383 VSS.n5618 VSS.n5617 29.2479
R384 VSS.n5619 VSS.n5618 29.2479
R385 VSS.n5619 VSS.n1205 29.2479
R386 VSS.n5625 VSS.n1205 29.2479
R387 VSS.n5626 VSS.n5625 29.2479
R388 VSS.n5627 VSS.n5626 29.2479
R389 VSS.n5627 VSS.n1201 29.2479
R390 VSS.n5633 VSS.n1201 29.2479
R391 VSS.n5634 VSS.n5633 29.2479
R392 VSS.n5635 VSS.n5634 29.2479
R393 VSS.n5635 VSS.n1197 29.2479
R394 VSS.n5641 VSS.n1197 29.2479
R395 VSS.n5642 VSS.n5641 29.2479
R396 VSS.n5643 VSS.n5642 29.2479
R397 VSS.n5643 VSS.n1193 29.2479
R398 VSS.n5649 VSS.n1193 29.2479
R399 VSS.n5650 VSS.n5649 29.2479
R400 VSS.n5651 VSS.n5650 29.2479
R401 VSS.n5651 VSS.n1189 29.2479
R402 VSS.n5657 VSS.n1189 29.2479
R403 VSS.n5658 VSS.n5657 29.2479
R404 VSS.n5659 VSS.n5658 29.2479
R405 VSS.n5659 VSS.n1185 29.2479
R406 VSS.n5665 VSS.n1185 29.2479
R407 VSS.n5666 VSS.n5665 29.2479
R408 VSS.n5667 VSS.n5666 29.2479
R409 VSS.n5667 VSS.n1181 29.2479
R410 VSS.n5673 VSS.n1181 29.2479
R411 VSS.n5674 VSS.n5673 29.2479
R412 VSS.n5675 VSS.n5674 29.2479
R413 VSS.n5675 VSS.n1177 29.2479
R414 VSS.n5681 VSS.n1177 29.2479
R415 VSS.n5682 VSS.n5681 29.2479
R416 VSS.n5683 VSS.n5682 29.2479
R417 VSS.n5683 VSS.n1173 29.2479
R418 VSS.n3610 VSS.n2702 26.6005
R419 VSS.n2702 VSS.n2698 26.6005
R420 VSS.n3611 VSS.n2703 26.1777
R421 VSS.n5456 VSS.n5455 21.9361
R422 VSS.n5448 VSS.n5447 21.4748
R423 VSS.n3602 VSS.n3601 20.1368
R424 VSS.n5689 VSS.n5688 19.8187
R425 VSS.n4314 VSS.n2622 16.1295
R426 VSS.n2086 VSS.n2085 15.9461
R427 VSS.n5341 VSS.n5340 15.9461
R428 VSS.n5409 VSS.n2109 15.9461
R429 VSS.n2525 VSS.n2524 15.9461
R430 VSS.n5713 VSS.n8 14.9684
R431 VSS.n5571 VSS.n5570 14.8601
R432 VSS.n5453 VSS.n5451 14.6638
R433 VSS.n5570 VSS.n5569 14.3883
R434 VSS.n2705 DVSS 14.1351
R435 VSS.n4306 VSS.n2625 14.1134
R436 VSS.n4530 VSS.n4528 12.4433
R437 VSS.n5689 VSS.n1173 12.0297
R438 VSS.n5314 VSS 10.8266
R439 VSS.n2191 VSS 10.8266
R440 VSS.n4844 VSS 10.8266
R441 VSS.n5714 VSS.n7 10.6065
R442 VSS.n2765 VSS.n1291 10.6065
R443 VSS.n5455 VSS.n1289 9.91235
R444 VSS.n2764 VSS.n7 8.06976
R445 VSS.n2765 VSS.n2764 8.03441
R446 VSS.n3884 VSS.n3781 7.77509
R447 VSS.n3785 VSS.n3780 7.77509
R448 VSS.n1745 VSS.n14 7.61966
R449 VSS.n1741 VSS.n1735 7.60677
R450 VSS.n1741 VSS.n1728 7.60677
R451 VSS.n3780 VSS.n3775 7.60296
R452 VSS.n3781 VSS.n3776 7.60296
R453 VSS.n1735 VSS.n1295 7.59387
R454 VSS.n1745 VSS.n1728 7.58957
R455 VSS.n5708 VSS.n14 7.28428
R456 VSS.n2078 VSS.n1295 7.26279
R457 VSS.n3251 VSS.n2701 6.95655
R458 VSS.n3523 VSS.t47 6.33948
R459 VSS.n3525 VSS.t35 6.33948
R460 VSS.n4196 VSS.n4195 6.3005
R461 VSS.n3528 VSS.n3527 6.3005
R462 VSS.n2732 VSS.n2731 6.3005
R463 VSS.n2792 VSS.n2791 6.3005
R464 VSS.n2794 VSS.n2793 6.3005
R465 VSS.n2632 VSS.n2631 6.3005
R466 VSS.n5714 VSS.n5713 6.19648
R467 VSS.n5451 VSS.n1291 6.19648
R468 VSS.n4862 VSS.n2414 5.57932
R469 VSS.n5702 VSS.n5701 5.42247
R470 VSS VSS.t54 5.2005
R471 VSS VSS.t52 5.2005
R472 VSS VSS.t51 5.2005
R473 VSS VSS.t53 5.2005
R474 VSS VSS.t55 5.2005
R475 VSS VSS.t50 5.2005
R476 VSS.n5270 VSS.n2223 5.2005
R477 VSS.n5287 VSS.n2223 5.2005
R478 VSS.n5270 VSS.n2224 5.2005
R479 VSS.n2224 VSS.n2210 5.2005
R480 VSS.n2224 VSS.n2208 5.2005
R481 VSS.n2224 VSS.n2211 5.2005
R482 VSS.n2224 VSS.n2207 5.2005
R483 VSS.n2224 VSS.n2212 5.2005
R484 VSS.n2224 VSS.n2206 5.2005
R485 VSS.n2224 VSS.n2213 5.2005
R486 VSS.n2224 VSS.n2205 5.2005
R487 VSS.n2224 VSS.n2214 5.2005
R488 VSS.n5284 VSS.n2224 5.2005
R489 VSS.n5287 VSS.n2224 5.2005
R490 VSS.n5270 VSS.n2217 5.2005
R491 VSS.n2217 VSS.n2210 5.2005
R492 VSS.n2217 VSS.n2208 5.2005
R493 VSS.n2217 VSS.n2211 5.2005
R494 VSS.n2217 VSS.n2207 5.2005
R495 VSS.n2217 VSS.n2212 5.2005
R496 VSS.n2217 VSS.n2206 5.2005
R497 VSS.n2217 VSS.n2213 5.2005
R498 VSS.n2217 VSS.n2205 5.2005
R499 VSS.n2217 VSS.n2214 5.2005
R500 VSS.n5287 VSS.n2217 5.2005
R501 VSS.n5270 VSS.n2225 5.2005
R502 VSS.n2225 VSS.n2210 5.2005
R503 VSS.n2225 VSS.n2208 5.2005
R504 VSS.n2225 VSS.n2211 5.2005
R505 VSS.n2225 VSS.n2207 5.2005
R506 VSS.n2225 VSS.n2212 5.2005
R507 VSS.n2225 VSS.n2206 5.2005
R508 VSS.n2225 VSS.n2213 5.2005
R509 VSS.n2225 VSS.n2205 5.2005
R510 VSS.n2225 VSS.n2214 5.2005
R511 VSS.n5287 VSS.n2225 5.2005
R512 VSS.n5270 VSS.n2216 5.2005
R513 VSS.n2216 VSS.n2210 5.2005
R514 VSS.n2216 VSS.n2208 5.2005
R515 VSS.n2216 VSS.n2211 5.2005
R516 VSS.n2216 VSS.n2207 5.2005
R517 VSS.n2216 VSS.n2212 5.2005
R518 VSS.n2216 VSS.n2206 5.2005
R519 VSS.n2216 VSS.n2213 5.2005
R520 VSS.n2216 VSS.n2205 5.2005
R521 VSS.n2216 VSS.n2214 5.2005
R522 VSS.n5287 VSS.n2216 5.2005
R523 VSS.n5270 VSS.n2226 5.2005
R524 VSS.n2226 VSS.n2210 5.2005
R525 VSS.n2226 VSS.n2208 5.2005
R526 VSS.n2226 VSS.n2211 5.2005
R527 VSS.n2226 VSS.n2207 5.2005
R528 VSS.n2226 VSS.n2212 5.2005
R529 VSS.n2226 VSS.n2206 5.2005
R530 VSS.n2226 VSS.n2213 5.2005
R531 VSS.n2226 VSS.n2205 5.2005
R532 VSS.n2226 VSS.n2214 5.2005
R533 VSS.n5287 VSS.n2226 5.2005
R534 VSS.n5270 VSS.n2215 5.2005
R535 VSS.n2215 VSS.n2210 5.2005
R536 VSS.n2215 VSS.n2208 5.2005
R537 VSS.n2215 VSS.n2211 5.2005
R538 VSS.n2215 VSS.n2207 5.2005
R539 VSS.n2215 VSS.n2212 5.2005
R540 VSS.n2215 VSS.n2206 5.2005
R541 VSS.n2215 VSS.n2213 5.2005
R542 VSS.n2215 VSS.n2205 5.2005
R543 VSS.n2215 VSS.n2214 5.2005
R544 VSS.n5287 VSS.n2215 5.2005
R545 VSS.n5288 VSS.n2210 5.2005
R546 VSS.n5288 VSS.n2208 5.2005
R547 VSS.n5288 VSS.n2211 5.2005
R548 VSS.n5288 VSS.n2207 5.2005
R549 VSS.n5288 VSS.n2212 5.2005
R550 VSS.n5288 VSS.n2206 5.2005
R551 VSS.n5288 VSS.n2213 5.2005
R552 VSS.n5288 VSS.n2205 5.2005
R553 VSS.n5288 VSS.n2214 5.2005
R554 VSS.n5288 VSS.n5287 5.2005
R555 VSS.n4528 VSS.n2546 5.08553
R556 VSS.n5268 VSS.n2232 4.84618
R557 VSS.n2230 VSS.n2217 4.84618
R558 VSS.n5282 VSS.n2225 4.84618
R559 VSS.n2229 VSS.n2216 4.84618
R560 VSS.n5283 VSS.n2226 4.84618
R561 VSS.n2228 VSS.n2215 4.84618
R562 VSS.n5288 VSS.n2204 4.84618
R563 VSS.n2232 VSS.n2223 4.84618
R564 VSS.n2230 VSS.n2224 4.84618
R565 VSS.n5282 VSS.n2217 4.84618
R566 VSS.n2229 VSS.n2225 4.84618
R567 VSS.n5283 VSS.n2216 4.84618
R568 VSS.n2228 VSS.n2226 4.84618
R569 VSS.n2215 VSS.n2204 4.84618
R570 VSS.n4303 VSS.n4302 4.82802
R571 VSS.n4285 VSS.n4284 4.66866
R572 VSS.n4686 VSS.n4685 4.66866
R573 VSS.n5314 VSS 4.5005
R574 VSS.n2191 VSS 4.5005
R575 VSS.n4844 VSS 4.5005
R576 VSS.n4437 VSS.n2608 4.5005
R577 VSS.n2614 VSS.n2608 4.5005
R578 VSS.n4439 VSS.n2608 4.5005
R579 VSS.n4437 VSS.n2610 4.5005
R580 VSS.n2614 VSS.n2610 4.5005
R581 VSS.n4439 VSS.n2610 4.5005
R582 VSS.n4439 VSS.n2607 4.5005
R583 VSS.n2614 VSS.n2607 4.5005
R584 VSS.n4437 VSS.n2607 4.5005
R585 VSS.n4439 VSS.n2611 4.5005
R586 VSS.n2614 VSS.n2611 4.5005
R587 VSS.n4437 VSS.n2611 4.5005
R588 VSS.n4437 VSS.n2606 4.5005
R589 VSS.n2614 VSS.n2606 4.5005
R590 VSS.n4439 VSS.n2606 4.5005
R591 VSS.n4439 VSS.n2612 4.5005
R592 VSS.n2614 VSS.n2612 4.5005
R593 VSS.n4437 VSS.n2612 4.5005
R594 VSS.n4437 VSS.n2605 4.5005
R595 VSS.n2614 VSS.n2605 4.5005
R596 VSS.n4439 VSS.n2605 4.5005
R597 VSS.n4439 VSS.n4438 4.5005
R598 VSS.n4438 VSS.n2614 4.5005
R599 VSS.n4438 VSS.n4437 4.5005
R600 VSS.n2074 VSS.n2073 4.5005
R601 VSS.n2073 VSS.n2071 4.5005
R602 VSS.n2073 VSS.n2067 4.5005
R603 VSS.n2072 VSS.n1594 4.5005
R604 VSS.n2073 VSS.n2072 4.5005
R605 VSS.n1597 VSS.n1595 4.5005
R606 VSS.n2062 VSS.n1595 4.5005
R607 VSS.n2065 VSS.n1595 4.5005
R608 VSS.n2066 VSS.n1597 4.5005
R609 VSS.n2066 VSS.n2065 4.5005
R610 VSS.n2065 VSS.n1602 4.5005
R611 VSS.n2065 VSS.n1605 4.5005
R612 VSS.n2065 VSS.n1601 4.5005
R613 VSS.n2065 VSS.n1607 4.5005
R614 VSS.n2065 VSS.n1600 4.5005
R615 VSS.n2065 VSS.n1609 4.5005
R616 VSS.n2065 VSS.n1599 4.5005
R617 VSS.n2064 VSS.n2062 4.5005
R618 VSS.n2065 VSS.n2064 4.5005
R619 VSS.n1854 VSS.n1797 4.5005
R620 VSS.n1857 VSS.n1797 4.5005
R621 VSS.n1797 VSS.n1792 4.5005
R622 VSS.n1854 VSS.n1820 4.5005
R623 VSS.n1820 VSS.n1792 4.5005
R624 VSS.n1807 VSS.n1792 4.5005
R625 VSS.n1806 VSS.n1792 4.5005
R626 VSS.n1804 VSS.n1792 4.5005
R627 VSS.n1803 VSS.n1792 4.5005
R628 VSS.n1801 VSS.n1792 4.5005
R629 VSS.n1800 VSS.n1792 4.5005
R630 VSS.n1799 VSS.n1792 4.5005
R631 VSS.n1857 VSS.n1856 4.5005
R632 VSS.n1856 VSS.n1792 4.5005
R633 VSS.n1819 VSS.n1818 4.5005
R634 VSS.n1818 VSS.n1810 4.5005
R635 VSS.n1810 VSS.n16 4.5005
R636 VSS.n1813 VSS.n16 4.5005
R637 VSS.n1815 VSS.n16 4.5005
R638 VSS.n1818 VSS.n1817 4.5005
R639 VSS.n1817 VSS.n16 4.5005
R640 VSS.n1144 VSS.n34 4.5005
R641 VSS.n1142 VSS.n1141 4.5005
R642 VSS.n1140 VSS.n1139 4.5005
R643 VSS.n1078 VSS.n77 4.5005
R644 VSS.n5701 VSS.n32 4.5005
R645 VSS.n1145 VSS.n33 4.5005
R646 VSS.n5703 VSS.n27 4.5005
R647 VSS.n27 VSS.n19 4.5005
R648 VSS.n27 VSS.n20 4.5005
R649 VSS.n27 VSS.n22 4.5005
R650 VSS.n24 VSS.n20 4.5005
R651 VSS.n24 VSS.n22 4.5005
R652 VSS.n5703 VSS.n28 4.5005
R653 VSS.n28 VSS.n19 4.5005
R654 VSS.n28 VSS.n20 4.5005
R655 VSS.n28 VSS.n22 4.5005
R656 VSS.n5703 VSS.n26 4.5005
R657 VSS.n26 VSS.n19 4.5005
R658 VSS.n26 VSS.n20 4.5005
R659 VSS.n26 VSS.n22 4.5005
R660 VSS.n30 VSS.n20 4.5005
R661 VSS.n30 VSS.n22 4.5005
R662 VSS.n25 VSS.n20 4.5005
R663 VSS.n25 VSS.n22 4.5005
R664 VSS.n5703 VSS.n29 4.5005
R665 VSS.n29 VSS.n19 4.5005
R666 VSS.n29 VSS.n20 4.5005
R667 VSS.n29 VSS.n22 4.5005
R668 VSS.n5704 VSS.n20 4.5005
R669 VSS.n5704 VSS.n22 4.5005
R670 VSS.n20 VSS.n18 4.5005
R671 VSS.n22 VSS.n18 4.5005
R672 VSS.n19 VSS.n18 4.5005
R673 VSS.n5703 VSS.n18 4.5005
R674 VSS.n5704 VSS.n19 4.5005
R675 VSS.n5704 VSS.n5703 4.5005
R676 VSS.n25 VSS.n19 4.5005
R677 VSS.n5703 VSS.n25 4.5005
R678 VSS.n30 VSS.n19 4.5005
R679 VSS.n5703 VSS.n30 4.5005
R680 VSS.n24 VSS.n19 4.5005
R681 VSS.n5703 VSS.n24 4.5005
R682 VSS.n5702 VSS.n22 4.5005
R683 VSS.n5702 VSS.n20 4.5005
R684 VSS.n5702 VSS.n19 4.5005
R685 VSS.n5703 VSS.n5702 4.5005
R686 VSS.n4135 VSS.n3768 4.5005
R687 VSS.n3771 VSS.n3768 4.5005
R688 VSS.n4134 VSS.n3771 4.5005
R689 VSS.n4135 VSS.n4134 4.5005
R690 VSS.n3918 VSS.n3769 4.5005
R691 VSS.n3784 VSS.n3769 4.5005
R692 VSS.n4145 VSS.n3759 4.5005
R693 VSS.n4145 VSS.n4144 4.5005
R694 VSS.n4144 VSS.n4143 4.5005
R695 VSS.n4143 VSS.n3759 4.5005
R696 VSS.n3879 VSS.n3760 4.5005
R697 VSS.n3880 VSS.n3879 4.5005
R698 VSS.n4163 VSS.n3731 4.5005
R699 VSS.n4163 VSS.n3733 4.5005
R700 VSS.n4163 VSS.n3730 4.5005
R701 VSS.n4163 VSS.n4162 4.5005
R702 VSS.n4162 VSS.n4161 4.5005
R703 VSS.n4161 VSS.n3730 4.5005
R704 VSS.n4161 VSS.n3733 4.5005
R705 VSS.n4161 VSS.n3731 4.5005
R706 VSS.n3788 VSS.n3732 4.5005
R707 VSS.n3818 VSS.n3732 4.5005
R708 VSS.n3818 VSS.n3817 4.5005
R709 VSS.n3818 VSS.n3789 4.5005
R710 VSS.n3819 VSS.n3788 4.5005
R711 VSS.n3819 VSS.n3818 4.5005
R712 VSS.n3948 VSS.n3888 4.5005
R713 VSS.n3948 VSS.n3892 4.5005
R714 VSS.n3948 VSS.n3893 4.5005
R715 VSS.n3948 VSS.n3900 4.5005
R716 VSS.n3905 VSS.n3900 4.5005
R717 VSS.n3905 VSS.n3893 4.5005
R718 VSS.n3905 VSS.n3892 4.5005
R719 VSS.n3905 VSS.n3888 4.5005
R720 VSS.n3890 VSS.n3887 4.5005
R721 VSS.n4118 VSS.n3890 4.5005
R722 VSS.n4118 VSS.n4117 4.5005
R723 VSS.n4118 VSS.n3889 4.5005
R724 VSS.n4119 VSS.n3887 4.5005
R725 VSS.n4119 VSS.n4118 4.5005
R726 VSS.n4066 VSS.n4057 4.5005
R727 VSS.n4066 VSS.n3964 4.5005
R728 VSS.n4072 VSS.n4057 4.5005
R729 VSS.n4072 VSS.n3964 4.5005
R730 VSS.n4079 VSS.n3964 4.5005
R731 VSS.n4079 VSS.n4057 4.5005
R732 VSS.n4088 VSS.n3965 4.5005
R733 VSS.n4090 VSS.n3965 4.5005
R734 VSS.n4090 VSS.n4089 4.5005
R735 VSS.n4089 VSS.n4088 4.5005
R736 VSS.n4077 VSS.n3964 4.5005
R737 VSS.n4077 VSS.n4057 4.5005
R738 VSS.n4072 VSS.n4070 4.5005
R739 VSS.n4072 VSS.n4071 4.5005
R740 VSS.n4084 VSS.n4058 4.5005
R741 VSS.n4085 VSS.n4084 4.5005
R742 VSS.n3726 VSS.n3724 4.5005
R743 VSS.n3746 VSS.n3726 4.5005
R744 VSS.n3951 VSS.n3907 4.5005
R745 VSS.n3952 VSS.n3951 4.5005
R746 VSS.n4086 VSS.n4058 4.5005
R747 VSS.n4086 VSS.n4085 4.5005
R748 VSS.n4131 VSS.n3774 4.5005
R749 VSS.n4131 VSS.n4130 4.5005
R750 VSS.n4146 VSS.n3758 4.5005
R751 VSS.n4146 VSS.n3755 4.5005
R752 VSS.n3719 VSS.n2654 4.5005
R753 VSS.n3719 VSS.n3718 4.5005
R754 VSS.n3718 VSS.n2663 4.5005
R755 VSS.n3718 VSS.n2660 4.5005
R756 VSS.n3718 VSS.n2665 4.5005
R757 VSS.n3718 VSS.n2659 4.5005
R758 VSS.n3718 VSS.n2667 4.5005
R759 VSS.n3718 VSS.n2658 4.5005
R760 VSS.n3718 VSS.n2669 4.5005
R761 VSS.n3718 VSS.n2657 4.5005
R762 VSS.n3717 VSS.n2654 4.5005
R763 VSS.n3718 VSS.n3717 4.5005
R764 VSS.n4170 VSS.n4169 4.5005
R765 VSS.n4169 VSS.n4168 4.5005
R766 VSS.n3805 VSS.n3804 4.5005
R767 VSS.n3805 VSS.n3796 4.5005
R768 VSS.n3806 VSS.n3805 4.5005
R769 VSS.n3806 VSS.n3720 4.5005
R770 VSS.n3796 VSS.n3720 4.5005
R771 VSS.n3804 VSS.n3720 4.5005
R772 VSS.n3866 VSS.n3841 4.5005
R773 VSS.n3821 VSS.n2648 4.5005
R774 VSS.n3835 VSS.n2644 4.5005
R775 VSS.n3835 VSS.n2648 4.5005
R776 VSS.n3823 VSS.n2644 4.5005
R777 VSS.n3823 VSS.n2648 4.5005
R778 VSS.n3821 VSS.n2644 4.5005
R779 VSS.n3866 VSS.n2644 4.5005
R780 VSS.n3866 VSS.n2648 4.5005
R781 VSS.n3867 VSS.n3866 4.5005
R782 VSS.n2561 VSS.n2556 4.5005
R783 VSS.n4514 VSS.n2561 4.5005
R784 VSS.n4512 VSS.n2561 4.5005
R785 VSS.n2563 VSS.n2556 4.5005
R786 VSS.n4514 VSS.n2563 4.5005
R787 VSS.n4512 VSS.n2563 4.5005
R788 VSS.n4512 VSS.n2560 4.5005
R789 VSS.n4514 VSS.n2560 4.5005
R790 VSS.n2560 VSS.n2556 4.5005
R791 VSS.n2564 VSS.n2556 4.5005
R792 VSS.n4514 VSS.n2564 4.5005
R793 VSS.n4512 VSS.n2564 4.5005
R794 VSS.n2559 VSS.n2556 4.5005
R795 VSS.n4514 VSS.n2559 4.5005
R796 VSS.n4512 VSS.n2559 4.5005
R797 VSS.n4512 VSS.n2565 4.5005
R798 VSS.n4514 VSS.n2565 4.5005
R799 VSS.n2565 VSS.n2556 4.5005
R800 VSS.n4512 VSS.n2558 4.5005
R801 VSS.n4514 VSS.n2558 4.5005
R802 VSS.n2558 VSS.n2556 4.5005
R803 VSS.n2566 VSS.n2556 4.5005
R804 VSS.n4514 VSS.n2566 4.5005
R805 VSS.n4512 VSS.n2566 4.5005
R806 VSS.n4512 VSS.n2557 4.5005
R807 VSS.n4514 VSS.n2557 4.5005
R808 VSS.n2557 VSS.n2556 4.5005
R809 VSS.n4513 VSS.n4512 4.5005
R810 VSS.n4514 VSS.n4513 4.5005
R811 VSS.n4513 VSS.n2556 4.5005
R812 VSS.n3864 VSS.n3863 4.5005
R813 VSS.n3860 VSS.n2616 4.5005
R814 VSS.n3865 VSS.n3864 4.5005
R815 VSS.n3865 VSS.n3859 4.5005
R816 VSS.n3865 VSS.n2616 4.5005
R817 VSS.n4856 VSS.n2416 4.5005
R818 VSS.n4856 VSS.n4855 4.5005
R819 VSS.n4855 VSS.n2424 4.5005
R820 VSS.n4855 VSS.n2421 4.5005
R821 VSS.n4855 VSS.n2426 4.5005
R822 VSS.n4855 VSS.n2420 4.5005
R823 VSS.n4855 VSS.n2428 4.5005
R824 VSS.n4855 VSS.n2419 4.5005
R825 VSS.n4855 VSS.n2430 4.5005
R826 VSS.n4855 VSS.n2418 4.5005
R827 VSS.n4854 VSS.n2416 4.5005
R828 VSS.n4855 VSS.n4854 4.5005
R829 VSS.n4685 VSS.n4684 4.5005
R830 VSS.n2502 VSS.n2501 4.5005
R831 VSS.n4676 VSS.n4675 4.5005
R832 VSS.n2508 VSS.n2506 4.5005
R833 VSS.n4279 VSS.n4277 4.5005
R834 VSS.n4284 VSS.n4283 4.5005
R835 VSS.n4853 VSS.n0 4.5005
R836 VSS.n4853 VSS.n4825 4.5005
R837 VSS.n4842 VSS.n0 4.5005
R838 VSS.n4836 VSS.n1 4.5005
R839 VSS.n4838 VSS.n1 4.5005
R840 VSS.n4840 VSS.n1 4.5005
R841 VSS.n4842 VSS.n1 4.5005
R842 VSS.n4853 VSS.n1 4.5005
R843 VSS.n4834 VSS.n4825 4.5005
R844 VSS.n4832 VSS.n4825 4.5005
R845 VSS.n4830 VSS.n4825 4.5005
R846 VSS.n4828 VSS.n4825 4.5005
R847 VSS.n4826 VSS.n1 4.5005
R848 VSS.n4826 VSS.n4825 4.5005
R849 VSS.n4861 VSS.n4856 4.24863
R850 VSS.n1289 VSS.n1288 4.05657
R851 VSS.n5458 VSS.n1288 4.05657
R852 VSS.n5458 VSS.n1286 4.05657
R853 VSS.n5462 VSS.n1286 4.05657
R854 VSS.n5462 VSS.n1284 4.05657
R855 VSS.n5466 VSS.n1284 4.05657
R856 VSS.n5466 VSS.n1282 4.05657
R857 VSS.n5470 VSS.n1282 4.05657
R858 VSS.n5470 VSS.n1280 4.05657
R859 VSS.n5474 VSS.n1280 4.05657
R860 VSS.n5474 VSS.n1278 4.05657
R861 VSS.n5478 VSS.n1278 4.05657
R862 VSS.n5478 VSS.n1276 4.05657
R863 VSS.n5482 VSS.n1276 4.05657
R864 VSS.n5482 VSS.n1274 4.05657
R865 VSS.n5486 VSS.n1274 4.05657
R866 VSS.n5486 VSS.n1272 4.05657
R867 VSS.n5490 VSS.n1272 4.05657
R868 VSS.n5490 VSS.n1270 4.05657
R869 VSS.n5494 VSS.n1270 4.05657
R870 VSS.n5494 VSS.n1268 4.05657
R871 VSS.n5498 VSS.n1268 4.05657
R872 VSS.n5498 VSS.n1266 4.05657
R873 VSS.n5502 VSS.n1266 4.05657
R874 VSS.n5502 VSS.n1264 4.05657
R875 VSS.n5506 VSS.n1264 4.05657
R876 VSS.n5506 VSS.n1262 4.05657
R877 VSS.n5510 VSS.n1262 4.05657
R878 VSS.n5510 VSS.n1260 4.05657
R879 VSS.n5514 VSS.n1260 4.05657
R880 VSS.n5514 VSS.n1258 4.05657
R881 VSS.n5518 VSS.n1258 4.05657
R882 VSS.n5518 VSS.n1256 4.05657
R883 VSS.n5522 VSS.n1256 4.05657
R884 VSS.n5522 VSS.n1254 4.05657
R885 VSS.n5526 VSS.n1254 4.05657
R886 VSS.n5526 VSS.n1252 4.05657
R887 VSS.n5530 VSS.n1252 4.05657
R888 VSS.n5530 VSS.n1250 4.05657
R889 VSS.n5534 VSS.n1250 4.05657
R890 VSS.n5534 VSS.n1248 4.05657
R891 VSS.n5538 VSS.n1248 4.05657
R892 VSS.n5538 VSS.n1246 4.05657
R893 VSS.n5542 VSS.n1246 4.05657
R894 VSS.n5542 VSS.n1244 4.05657
R895 VSS.n5546 VSS.n1244 4.05657
R896 VSS.n5546 VSS.n1242 4.05657
R897 VSS.n5550 VSS.n1242 4.05657
R898 VSS.n5550 VSS.n1240 4.05657
R899 VSS.n5554 VSS.n1240 4.05657
R900 VSS.n5554 VSS.n1238 4.05657
R901 VSS.n5558 VSS.n1238 4.05657
R902 VSS.n5558 VSS.n1236 4.05657
R903 VSS.n5562 VSS.n1236 4.05657
R904 VSS.n5562 VSS.n1234 4.05657
R905 VSS.n5567 VSS.n1234 4.05657
R906 VSS.n5567 VSS.n1232 4.05657
R907 VSS.n5572 VSS.n1232 4.05657
R908 VSS.n5572 VSS.n1230 4.05657
R909 VSS.n5576 VSS.n1230 4.05657
R910 VSS.n5576 VSS.n1228 4.05657
R911 VSS.n5580 VSS.n1228 4.05657
R912 VSS.n5580 VSS.n1226 4.05657
R913 VSS.n5584 VSS.n1226 4.05657
R914 VSS.n5584 VSS.n1224 4.05657
R915 VSS.n5588 VSS.n1224 4.05657
R916 VSS.n5588 VSS.n1222 4.05657
R917 VSS.n5592 VSS.n1222 4.05657
R918 VSS.n5592 VSS.n1220 4.05657
R919 VSS.n5596 VSS.n1220 4.05657
R920 VSS.n5596 VSS.n1218 4.05657
R921 VSS.n5600 VSS.n1218 4.05657
R922 VSS.n5600 VSS.n1216 4.05657
R923 VSS.n5604 VSS.n1216 4.05657
R924 VSS.n5604 VSS.n1214 4.05657
R925 VSS.n5608 VSS.n1214 4.05657
R926 VSS.n5608 VSS.n1212 4.05657
R927 VSS.n5612 VSS.n1212 4.05657
R928 VSS.n5612 VSS.n1210 4.05657
R929 VSS.n5616 VSS.n1210 4.05657
R930 VSS.n5616 VSS.n1208 4.05657
R931 VSS.n5620 VSS.n1208 4.05657
R932 VSS.n5620 VSS.n1206 4.05657
R933 VSS.n5624 VSS.n1206 4.05657
R934 VSS.n5624 VSS.n1204 4.05657
R935 VSS.n5628 VSS.n1204 4.05657
R936 VSS.n5628 VSS.n1202 4.05657
R937 VSS.n5632 VSS.n1202 4.05657
R938 VSS.n5632 VSS.n1200 4.05657
R939 VSS.n5636 VSS.n1200 4.05657
R940 VSS.n5636 VSS.n1198 4.05657
R941 VSS.n5640 VSS.n1198 4.05657
R942 VSS.n5640 VSS.n1196 4.05657
R943 VSS.n5644 VSS.n1196 4.05657
R944 VSS.n5644 VSS.n1194 4.05657
R945 VSS.n5648 VSS.n1194 4.05657
R946 VSS.n5648 VSS.n1192 4.05657
R947 VSS.n5652 VSS.n1192 4.05657
R948 VSS.n5652 VSS.n1190 4.05657
R949 VSS.n5656 VSS.n1190 4.05657
R950 VSS.n5656 VSS.n1188 4.05657
R951 VSS.n5660 VSS.n1188 4.05657
R952 VSS.n5660 VSS.n1186 4.05657
R953 VSS.n5664 VSS.n1186 4.05657
R954 VSS.n5664 VSS.n1184 4.05657
R955 VSS.n5668 VSS.n1184 4.05657
R956 VSS.n5668 VSS.n1182 4.05657
R957 VSS.n5672 VSS.n1182 4.05657
R958 VSS.n5672 VSS.n1180 4.05657
R959 VSS.n5676 VSS.n1180 4.05657
R960 VSS.n5676 VSS.n1178 4.05657
R961 VSS.n5680 VSS.n1178 4.05657
R962 VSS.n5680 VSS.n1176 4.05657
R963 VSS.n5684 VSS.n1176 4.05657
R964 VSS.n5684 VSS.n1174 4.05657
R965 VSS.n5688 VSS.n1174 4.05657
R966 VSS.n3260 VSS.n2633 3.8345
R967 VSS.n4861 VSS.n4860 3.7805
R968 VSS.n4862 VSS.n4861 3.77031
R969 VSS.n5326 VSS.n5322 3.68022
R970 VSS.n3681 VSS.n2694 3.37368
R971 VSS.n4195 VSS 3.18489
R972 VSS.n3527 VSS 3.18489
R973 VSS.n2731 VSS 3.18489
R974 VSS.n2791 VSS 3.18489
R975 VSS.n2793 VSS 3.18489
R976 VSS.n2631 VSS 3.18489
R977 VSS.n2513 VSS.t23 3.17811
R978 VSS.n3253 VSS.t5 3.17811
R979 VSS.n4857 VSS.t37 3.17811
R980 VSS.n2700 VSS.t17 3.17811
R981 VSS.n2699 VSS.t3 3.17811
R982 VSS.n4323 VSS.n2194 3.02469
R983 VSS.n4854 VSS.n4853 2.95295
R984 VSS.n5421 VSS.n2103 2.90887
R985 VSS.n5315 VSS.n5314 2.81187
R986 VSS.n2192 VSS.n2191 2.81187
R987 VSS.n4845 VSS.n4844 2.81187
R988 VSS.n5183 VSS.n5182 2.75988
R989 VSS.n5688 VSS.n5687 2.6005
R990 VSS.n5686 VSS.n1174 2.6005
R991 VSS.n1174 VSS.n1173 2.6005
R992 VSS.n5685 VSS.n5684 2.6005
R993 VSS.n5684 VSS.n5683 2.6005
R994 VSS.n1176 VSS.n1175 2.6005
R995 VSS.n5682 VSS.n1176 2.6005
R996 VSS.n5680 VSS.n5679 2.6005
R997 VSS.n5681 VSS.n5680 2.6005
R998 VSS.n5678 VSS.n1178 2.6005
R999 VSS.n1178 VSS.n1177 2.6005
R1000 VSS.n5677 VSS.n5676 2.6005
R1001 VSS.n5676 VSS.n5675 2.6005
R1002 VSS.n1180 VSS.n1179 2.6005
R1003 VSS.n5674 VSS.n1180 2.6005
R1004 VSS.n5672 VSS.n5671 2.6005
R1005 VSS.n5673 VSS.n5672 2.6005
R1006 VSS.n5670 VSS.n1182 2.6005
R1007 VSS.n1182 VSS.n1181 2.6005
R1008 VSS.n5669 VSS.n5668 2.6005
R1009 VSS.n5668 VSS.n5667 2.6005
R1010 VSS.n1184 VSS.n1183 2.6005
R1011 VSS.n5666 VSS.n1184 2.6005
R1012 VSS.n5664 VSS.n5663 2.6005
R1013 VSS.n5665 VSS.n5664 2.6005
R1014 VSS.n5662 VSS.n1186 2.6005
R1015 VSS.n1186 VSS.n1185 2.6005
R1016 VSS.n5661 VSS.n5660 2.6005
R1017 VSS.n5660 VSS.n5659 2.6005
R1018 VSS.n1188 VSS.n1187 2.6005
R1019 VSS.n5658 VSS.n1188 2.6005
R1020 VSS.n5656 VSS.n5655 2.6005
R1021 VSS.n5657 VSS.n5656 2.6005
R1022 VSS.n5654 VSS.n1190 2.6005
R1023 VSS.n1190 VSS.n1189 2.6005
R1024 VSS.n5653 VSS.n5652 2.6005
R1025 VSS.n5652 VSS.n5651 2.6005
R1026 VSS.n1192 VSS.n1191 2.6005
R1027 VSS.n5650 VSS.n1192 2.6005
R1028 VSS.n5648 VSS.n5647 2.6005
R1029 VSS.n5649 VSS.n5648 2.6005
R1030 VSS.n5646 VSS.n1194 2.6005
R1031 VSS.n1194 VSS.n1193 2.6005
R1032 VSS.n5645 VSS.n5644 2.6005
R1033 VSS.n5644 VSS.n5643 2.6005
R1034 VSS.n1196 VSS.n1195 2.6005
R1035 VSS.n5642 VSS.n1196 2.6005
R1036 VSS.n5640 VSS.n5639 2.6005
R1037 VSS.n5641 VSS.n5640 2.6005
R1038 VSS.n5638 VSS.n1198 2.6005
R1039 VSS.n1198 VSS.n1197 2.6005
R1040 VSS.n5637 VSS.n5636 2.6005
R1041 VSS.n5636 VSS.n5635 2.6005
R1042 VSS.n1200 VSS.n1199 2.6005
R1043 VSS.n5634 VSS.n1200 2.6005
R1044 VSS.n5632 VSS.n5631 2.6005
R1045 VSS.n5633 VSS.n5632 2.6005
R1046 VSS.n5630 VSS.n1202 2.6005
R1047 VSS.n1202 VSS.n1201 2.6005
R1048 VSS.n5629 VSS.n5628 2.6005
R1049 VSS.n5628 VSS.n5627 2.6005
R1050 VSS.n1204 VSS.n1203 2.6005
R1051 VSS.n5626 VSS.n1204 2.6005
R1052 VSS.n5624 VSS.n5623 2.6005
R1053 VSS.n5625 VSS.n5624 2.6005
R1054 VSS.n5622 VSS.n1206 2.6005
R1055 VSS.n1206 VSS.n1205 2.6005
R1056 VSS.n5621 VSS.n5620 2.6005
R1057 VSS.n5620 VSS.n5619 2.6005
R1058 VSS.n1208 VSS.n1207 2.6005
R1059 VSS.n5618 VSS.n1208 2.6005
R1060 VSS.n5616 VSS.n5615 2.6005
R1061 VSS.n5617 VSS.n5616 2.6005
R1062 VSS.n5614 VSS.n1210 2.6005
R1063 VSS.n1210 VSS.n1209 2.6005
R1064 VSS.n5613 VSS.n5612 2.6005
R1065 VSS.n5612 VSS.n5611 2.6005
R1066 VSS.n1212 VSS.n1211 2.6005
R1067 VSS.n5610 VSS.n1212 2.6005
R1068 VSS.n5608 VSS.n5607 2.6005
R1069 VSS.n5609 VSS.n5608 2.6005
R1070 VSS.n5606 VSS.n1214 2.6005
R1071 VSS.n1214 VSS.n1213 2.6005
R1072 VSS.n5605 VSS.n5604 2.6005
R1073 VSS.n5604 VSS.n5603 2.6005
R1074 VSS.n1216 VSS.n1215 2.6005
R1075 VSS.n5602 VSS.n1216 2.6005
R1076 VSS.n5600 VSS.n5599 2.6005
R1077 VSS.n5601 VSS.n5600 2.6005
R1078 VSS.n5598 VSS.n1218 2.6005
R1079 VSS.n1218 VSS.n1217 2.6005
R1080 VSS.n5597 VSS.n5596 2.6005
R1081 VSS.n5596 VSS.n5595 2.6005
R1082 VSS.n1220 VSS.n1219 2.6005
R1083 VSS.n5594 VSS.n1220 2.6005
R1084 VSS.n5592 VSS.n5591 2.6005
R1085 VSS.n5593 VSS.n5592 2.6005
R1086 VSS.n5590 VSS.n1222 2.6005
R1087 VSS.n1222 VSS.n1221 2.6005
R1088 VSS.n5589 VSS.n5588 2.6005
R1089 VSS.n5588 VSS.n5587 2.6005
R1090 VSS.n1224 VSS.n1223 2.6005
R1091 VSS.n5586 VSS.n1224 2.6005
R1092 VSS.n5584 VSS.n5583 2.6005
R1093 VSS.n5585 VSS.n5584 2.6005
R1094 VSS.n5582 VSS.n1226 2.6005
R1095 VSS.n1226 VSS.n1225 2.6005
R1096 VSS.n5581 VSS.n5580 2.6005
R1097 VSS.n5580 VSS.n5579 2.6005
R1098 VSS.n1228 VSS.n1227 2.6005
R1099 VSS.n5578 VSS.n1228 2.6005
R1100 VSS.n5576 VSS.n5575 2.6005
R1101 VSS.n5577 VSS.n5576 2.6005
R1102 VSS.n5574 VSS.n1230 2.6005
R1103 VSS.n1230 VSS.n1229 2.6005
R1104 VSS.n5573 VSS.n5572 2.6005
R1105 VSS.n5572 VSS.n5571 2.6005
R1106 VSS.n5565 VSS.n1232 2.6005
R1107 VSS.n5569 VSS.n1232 2.6005
R1108 VSS.n5567 VSS.n5566 2.6005
R1109 VSS.n5568 VSS.n5567 2.6005
R1110 VSS.n5564 VSS.n1234 2.6005
R1111 VSS.n1234 VSS.n1233 2.6005
R1112 VSS.n5563 VSS.n5562 2.6005
R1113 VSS.n5562 VSS.n5561 2.6005
R1114 VSS.n1236 VSS.n1235 2.6005
R1115 VSS.n5560 VSS.n1236 2.6005
R1116 VSS.n5558 VSS.n5557 2.6005
R1117 VSS.n5559 VSS.n5558 2.6005
R1118 VSS.n5556 VSS.n1238 2.6005
R1119 VSS.n1238 VSS.n1237 2.6005
R1120 VSS.n5555 VSS.n5554 2.6005
R1121 VSS.n5554 VSS.n5553 2.6005
R1122 VSS.n1240 VSS.n1239 2.6005
R1123 VSS.n5552 VSS.n1240 2.6005
R1124 VSS.n5550 VSS.n5549 2.6005
R1125 VSS.n5551 VSS.n5550 2.6005
R1126 VSS.n5548 VSS.n1242 2.6005
R1127 VSS.n1242 VSS.n1241 2.6005
R1128 VSS.n5547 VSS.n5546 2.6005
R1129 VSS.n5546 VSS.n5545 2.6005
R1130 VSS.n1244 VSS.n1243 2.6005
R1131 VSS.n5544 VSS.n1244 2.6005
R1132 VSS.n5542 VSS.n5541 2.6005
R1133 VSS.n5543 VSS.n5542 2.6005
R1134 VSS.n5540 VSS.n1246 2.6005
R1135 VSS.n1246 VSS.n1245 2.6005
R1136 VSS.n5539 VSS.n5538 2.6005
R1137 VSS.n5538 VSS.n5537 2.6005
R1138 VSS.n1248 VSS.n1247 2.6005
R1139 VSS.n5536 VSS.n1248 2.6005
R1140 VSS.n5534 VSS.n5533 2.6005
R1141 VSS.n5535 VSS.n5534 2.6005
R1142 VSS.n5532 VSS.n1250 2.6005
R1143 VSS.n1250 VSS.n1249 2.6005
R1144 VSS.n5531 VSS.n5530 2.6005
R1145 VSS.n5530 VSS.n5529 2.6005
R1146 VSS.n1252 VSS.n1251 2.6005
R1147 VSS.n5528 VSS.n1252 2.6005
R1148 VSS.n5526 VSS.n5525 2.6005
R1149 VSS.n5527 VSS.n5526 2.6005
R1150 VSS.n5524 VSS.n1254 2.6005
R1151 VSS.n1254 VSS.n1253 2.6005
R1152 VSS.n5523 VSS.n5522 2.6005
R1153 VSS.n5522 VSS.n5521 2.6005
R1154 VSS.n1256 VSS.n1255 2.6005
R1155 VSS.n5520 VSS.n1256 2.6005
R1156 VSS.n5518 VSS.n5517 2.6005
R1157 VSS.n5519 VSS.n5518 2.6005
R1158 VSS.n5516 VSS.n1258 2.6005
R1159 VSS.n1258 VSS.n1257 2.6005
R1160 VSS.n5515 VSS.n5514 2.6005
R1161 VSS.n5514 VSS.n5513 2.6005
R1162 VSS.n1260 VSS.n1259 2.6005
R1163 VSS.n5512 VSS.n1260 2.6005
R1164 VSS.n5510 VSS.n5509 2.6005
R1165 VSS.n5511 VSS.n5510 2.6005
R1166 VSS.n5508 VSS.n1262 2.6005
R1167 VSS.n1262 VSS.n1261 2.6005
R1168 VSS.n5507 VSS.n5506 2.6005
R1169 VSS.n5506 VSS.n5505 2.6005
R1170 VSS.n1264 VSS.n1263 2.6005
R1171 VSS.n5504 VSS.n1264 2.6005
R1172 VSS.n5502 VSS.n5501 2.6005
R1173 VSS.n5503 VSS.n5502 2.6005
R1174 VSS.n5500 VSS.n1266 2.6005
R1175 VSS.n1266 VSS.n1265 2.6005
R1176 VSS.n5499 VSS.n5498 2.6005
R1177 VSS.n5498 VSS.n5497 2.6005
R1178 VSS.n1268 VSS.n1267 2.6005
R1179 VSS.n5496 VSS.n1268 2.6005
R1180 VSS.n5494 VSS.n5493 2.6005
R1181 VSS.n5495 VSS.n5494 2.6005
R1182 VSS.n5492 VSS.n1270 2.6005
R1183 VSS.n1270 VSS.n1269 2.6005
R1184 VSS.n5491 VSS.n5490 2.6005
R1185 VSS.n5490 VSS.n5489 2.6005
R1186 VSS.n1272 VSS.n1271 2.6005
R1187 VSS.n5488 VSS.n1272 2.6005
R1188 VSS.n5486 VSS.n5485 2.6005
R1189 VSS.n5487 VSS.n5486 2.6005
R1190 VSS.n5484 VSS.n1274 2.6005
R1191 VSS.n1274 VSS.n1273 2.6005
R1192 VSS.n5483 VSS.n5482 2.6005
R1193 VSS.n5482 VSS.n5481 2.6005
R1194 VSS.n1276 VSS.n1275 2.6005
R1195 VSS.n5480 VSS.n1276 2.6005
R1196 VSS.n5478 VSS.n5477 2.6005
R1197 VSS.n5479 VSS.n5478 2.6005
R1198 VSS.n5476 VSS.n1278 2.6005
R1199 VSS.n1278 VSS.n1277 2.6005
R1200 VSS.n5475 VSS.n5474 2.6005
R1201 VSS.n5474 VSS.n5473 2.6005
R1202 VSS.n1280 VSS.n1279 2.6005
R1203 VSS.n5472 VSS.n1280 2.6005
R1204 VSS.n5470 VSS.n5469 2.6005
R1205 VSS.n5471 VSS.n5470 2.6005
R1206 VSS.n5468 VSS.n1282 2.6005
R1207 VSS.n1282 VSS.n1281 2.6005
R1208 VSS.n5467 VSS.n5466 2.6005
R1209 VSS.n5466 VSS.n5465 2.6005
R1210 VSS.n1284 VSS.n1283 2.6005
R1211 VSS.n5464 VSS.n1284 2.6005
R1212 VSS.n5462 VSS.n5461 2.6005
R1213 VSS.n5463 VSS.n5462 2.6005
R1214 VSS.n5460 VSS.n1286 2.6005
R1215 VSS.n1286 VSS.n1285 2.6005
R1216 VSS.n5459 VSS.n5458 2.6005
R1217 VSS.n5458 VSS.n5457 2.6005
R1218 VSS.n1288 VSS.n1287 2.6005
R1219 VSS.n5456 VSS.n1288 2.6005
R1220 VSS.n5452 VSS.n1289 2.6005
R1221 VSS.n5251 DVSS 2.57245
R1222 VSS.n5252 VSS.n5251 2.57069
R1223 VSS.n2167 VSS.n18 2.43717
R1224 VSS.n2223 VSS.n2222 2.41753
R1225 VSS.n2223 VSS.n2221 2.41753
R1226 VSS.n2223 VSS.n2220 2.41753
R1227 VSS.n2223 VSS.n2219 2.41753
R1228 VSS.n5281 VSS.n2223 2.41753
R1229 VSS.n5269 VSS.n5268 2.41753
R1230 VSS.n5268 VSS.n2236 2.41753
R1231 VSS.n5268 VSS.n2235 2.41753
R1232 VSS.n5268 VSS.n2234 2.41753
R1233 VSS.n5268 VSS.n2233 2.41753
R1234 VSS.n5268 VSS.n2218 2.41753
R1235 VSS.n5288 VSS.n2209 2.41753
R1236 VSS.n5336 VSS.n5335 2.41274
R1237 VSS.n5337 VSS.n5336 2.41274
R1238 VSS.n5431 VSS.n5430 2.41274
R1239 VSS.n5430 VSS.n5429 2.41274
R1240 VSS.n5251 DVSS 2.32795
R1241 VSS.n3260 VSS.n3259 2.311
R1242 VSS.n3605 VSS.n2694 2.28324
R1243 VSS.n3828 VSS.n3825 2.2728
R1244 VSS.n5425 VSS.n5424 2.25682
R1245 VSS.n5418 VSS.n2104 2.25682
R1246 VSS.n2528 VSS.n2103 2.25392
R1247 VSS.n653 VSS.n358 2.2505
R1248 VSS.n652 VSS.n651 2.2505
R1249 VSS.n650 VSS.n359 2.2505
R1250 VSS.n649 VSS.n648 2.2505
R1251 VSS.n647 VSS.n360 2.2505
R1252 VSS.n646 VSS.n645 2.2505
R1253 VSS.n644 VSS.n361 2.2505
R1254 VSS.n643 VSS.n642 2.2505
R1255 VSS.n641 VSS.n362 2.2505
R1256 VSS.n640 VSS.n639 2.2505
R1257 VSS.n638 VSS.n363 2.2505
R1258 VSS.n637 VSS.n636 2.2505
R1259 VSS.n634 VSS.n364 2.2505
R1260 VSS.n633 VSS.n632 2.2505
R1261 VSS.n537 VSS.n536 2.2505
R1262 VSS.n538 VSS.n534 2.2505
R1263 VSS.n540 VSS.n539 2.2505
R1264 VSS.n541 VSS.n533 2.2505
R1265 VSS.n543 VSS.n542 2.2505
R1266 VSS.n544 VSS.n532 2.2505
R1267 VSS.n546 VSS.n545 2.2505
R1268 VSS.n547 VSS.n531 2.2505
R1269 VSS.n549 VSS.n548 2.2505
R1270 VSS.n550 VSS.n530 2.2505
R1271 VSS.n552 VSS.n551 2.2505
R1272 VSS.n553 VSS.n529 2.2505
R1273 VSS.n555 VSS.n554 2.2505
R1274 VSS.n556 VSS.n528 2.2505
R1275 VSS.n558 VSS.n557 2.2505
R1276 VSS.n559 VSS.n527 2.2505
R1277 VSS.n561 VSS.n560 2.2505
R1278 VSS.n562 VSS.n526 2.2505
R1279 VSS.n564 VSS.n563 2.2505
R1280 VSS.n565 VSS.n525 2.2505
R1281 VSS.n567 VSS.n566 2.2505
R1282 VSS.n568 VSS.n524 2.2505
R1283 VSS.n570 VSS.n569 2.2505
R1284 VSS.n666 VSS.n354 2.2505
R1285 VSS.n668 VSS.n667 2.2505
R1286 VSS.n665 VSS.n353 2.2505
R1287 VSS.n664 VSS.n663 2.2505
R1288 VSS.n662 VSS.n355 2.2505
R1289 VSS.n661 VSS.n660 2.2505
R1290 VSS.n659 VSS.n356 2.2505
R1291 VSS.n658 VSS.n657 2.2505
R1292 VSS.n656 VSS.n357 2.2505
R1293 VSS.n655 VSS.n654 2.2505
R1294 VSS.n105 VSS.n104 2.2505
R1295 VSS.n184 VSS.n183 2.2505
R1296 VSS.n185 VSS.n182 2.2505
R1297 VSS.n187 VSS.n186 2.2505
R1298 VSS.n188 VSS.n181 2.2505
R1299 VSS.n190 VSS.n189 2.2505
R1300 VSS.n191 VSS.n180 2.2505
R1301 VSS.n193 VSS.n192 2.2505
R1302 VSS.n196 VSS.n195 2.2505
R1303 VSS.n197 VSS.n178 2.2505
R1304 VSS.n199 VSS.n198 2.2505
R1305 VSS.n200 VSS.n177 2.2505
R1306 VSS.n202 VSS.n201 2.2505
R1307 VSS.n203 VSS.n176 2.2505
R1308 VSS.n205 VSS.n204 2.2505
R1309 VSS.n206 VSS.n175 2.2505
R1310 VSS.n208 VSS.n207 2.2505
R1311 VSS.n209 VSS.n174 2.2505
R1312 VSS.n211 VSS.n210 2.2505
R1313 VSS.n212 VSS.n173 2.2505
R1314 VSS.n214 VSS.n213 2.2505
R1315 VSS.n215 VSS.n172 2.2505
R1316 VSS.n914 VSS.n913 2.2505
R1317 VSS.n912 VSS.n171 2.2505
R1318 VSS.n233 VSS.n218 2.2505
R1319 VSS.n235 VSS.n234 2.2505
R1320 VSS.n236 VSS.n232 2.2505
R1321 VSS.n238 VSS.n237 2.2505
R1322 VSS.n239 VSS.n231 2.2505
R1323 VSS.n241 VSS.n240 2.2505
R1324 VSS.n242 VSS.n230 2.2505
R1325 VSS.n244 VSS.n243 2.2505
R1326 VSS.n245 VSS.n229 2.2505
R1327 VSS.n247 VSS.n246 2.2505
R1328 VSS.n248 VSS.n228 2.2505
R1329 VSS.n250 VSS.n249 2.2505
R1330 VSS.n251 VSS.n227 2.2505
R1331 VSS.n253 VSS.n252 2.2505
R1332 VSS.n254 VSS.n226 2.2505
R1333 VSS.n256 VSS.n255 2.2505
R1334 VSS.n257 VSS.n225 2.2505
R1335 VSS.n259 VSS.n258 2.2505
R1336 VSS.n260 VSS.n224 2.2505
R1337 VSS.n262 VSS.n261 2.2505
R1338 VSS.n903 VSS.n223 2.2505
R1339 VSS.n905 VSS.n904 2.2505
R1340 VSS.n194 VSS.n179 2.2505
R1341 VSS.n3912 VSS.n3908 2.2505
R1342 VSS.n3941 VSS.n3940 2.2505
R1343 VSS.n3931 VSS.n3930 2.2505
R1344 VSS.n3925 VSS.n3924 2.2505
R1345 VSS.n3872 VSS.n3745 2.2505
R1346 VSS.n4153 VSS.n4152 2.2505
R1347 VSS.n3751 VSS.n3742 2.2505
R1348 VSS.n3749 VSS.n3735 2.2505
R1349 VSS.n4059 VSS.n3958 2.2505
R1350 VSS.n4099 VSS.n4098 2.2505
R1351 VSS.n3956 VSS.n3903 2.2505
R1352 VSS.n4106 VSS.n4105 2.2505
R1353 VSS.n4082 VSS.n4064 2.2505
R1354 VSS.n4074 VSS.n4073 2.2505
R1355 VSS.n4076 VSS.n4075 2.2505
R1356 VSS.n4078 VSS.n4065 2.2505
R1357 VSS.n4081 VSS.n4080 2.2505
R1358 VSS.n4062 VSS.n4061 2.2505
R1359 VSS.n4060 VSS.n3955 2.2505
R1360 VSS.n4100 VSS.n3954 2.2505
R1361 VSS.n4102 VSS.n4101 2.2505
R1362 VSS.n4104 VSS.n4103 2.2505
R1363 VSS.n3953 VSS.n3902 2.2505
R1364 VSS.n3946 VSS.n3945 2.2505
R1365 VSS.n3944 VSS.n3943 2.2505
R1366 VSS.n3942 VSS.n3909 2.2505
R1367 VSS.n3927 VSS.n3910 2.2505
R1368 VSS.n3929 VSS.n3928 2.2505
R1369 VSS.n3926 VSS.n3773 2.2505
R1370 VSS.n4149 VSS.n4148 2.2505
R1371 VSS.n4151 VSS.n4150 2.2505
R1372 VSS.n3754 VSS.n3744 2.2505
R1373 VSS.n3753 VSS.n3752 2.2505
R1374 VSS.n3750 VSS.n3748 2.2505
R1375 VSS.n3747 VSS.n3725 2.2505
R1376 VSS.n4167 VSS.n4166 2.2505
R1377 VSS.n2652 VSS.n2650 2.2505
R1378 VSS.n4172 VSS.n4171 2.2505
R1379 VSS.n3797 VSS.n2651 2.2505
R1380 VSS.n4174 VSS.n4173 2.2505
R1381 VSS.n3828 VSS.n3827 2.2505
R1382 VSS.n3839 VSS.n3838 2.2505
R1383 VSS.n3837 VSS.n3836 2.2505
R1384 VSS.n3834 VSS.n3833 2.2505
R1385 VSS.n3832 VSS.n3831 2.2505
R1386 VSS.n3830 VSS.n3824 2.2505
R1387 VSS.n3261 VSS.n3260 2.2505
R1388 VSS.n2075 VSS.n2074 2.24683
R1389 VSS.n2069 VSS.n2068 2.24683
R1390 VSS.n1819 VSS.n1809 2.24683
R1391 VSS.n5699 VSS.n32 2.24648
R1392 VSS.n5697 VSS.n32 2.24648
R1393 VSS.n1148 VSS.n32 2.24648
R1394 VSS.n1146 VSS.n32 2.24648
R1395 VSS.n1147 VSS.n33 2.24648
R1396 VSS.n1149 VSS.n33 2.24648
R1397 VSS.n5698 VSS.n33 2.24648
R1398 VSS.n5700 VSS.n33 2.24648
R1399 VSS.n3863 VSS.n3862 2.24442
R1400 VSS.n3861 VSS.n3860 2.24442
R1401 VSS.n2076 VSS.n1593 2.24405
R1402 VSS.n2070 VSS.n1594 2.24405
R1403 VSS.n2076 VSS.n1592 2.24405
R1404 VSS.n1812 VSS.n1811 2.24405
R1405 VSS.n1818 VSS.n1814 2.24405
R1406 VSS.n1816 VSS.n1811 2.24405
R1407 VSS.n3816 VSS.n3788 2.24386
R1408 VSS.n3815 VSS.n3814 2.24386
R1409 VSS.n3814 VSS.n3787 2.24386
R1410 VSS.n4116 VSS.n3887 2.24386
R1411 VSS.n4115 VSS.n4114 2.24386
R1412 VSS.n4114 VSS.n3886 2.24386
R1413 VSS.n1604 VSS.n1597 2.24304
R1414 VSS.n2062 VSS.n1596 2.24304
R1415 VSS.n1606 VSS.n1597 2.24304
R1416 VSS.n2062 VSS.n1612 2.24304
R1417 VSS.n1608 VSS.n1597 2.24304
R1418 VSS.n2062 VSS.n1611 2.24304
R1419 VSS.n2063 VSS.n1597 2.24304
R1420 VSS.n2062 VSS.n1610 2.24304
R1421 VSS.n1857 VSS.n1796 2.24304
R1422 VSS.n1854 VSS.n1808 2.24304
R1423 VSS.n1857 VSS.n1795 2.24304
R1424 VSS.n1854 VSS.n1805 2.24304
R1425 VSS.n1857 VSS.n1794 2.24304
R1426 VSS.n1854 VSS.n1802 2.24304
R1427 VSS.n1857 VSS.n1793 2.24304
R1428 VSS.n1855 VSS.n1854 2.24304
R1429 VSS.n3715 VSS.n2655 2.24304
R1430 VSS.n2662 VSS.n2654 2.24304
R1431 VSS.n3715 VSS.n2673 2.24304
R1432 VSS.n2664 VSS.n2654 2.24304
R1433 VSS.n3715 VSS.n2672 2.24304
R1434 VSS.n2666 VSS.n2654 2.24304
R1435 VSS.n3715 VSS.n2671 2.24304
R1436 VSS.n2668 VSS.n2654 2.24304
R1437 VSS.n3716 VSS.n3715 2.24304
R1438 VSS.n2423 VSS.n2416 2.24304
R1439 VSS.n3372 VSS.n2415 2.24304
R1440 VSS.n2425 VSS.n2416 2.24304
R1441 VSS.n3372 VSS.n3369 2.24304
R1442 VSS.n2427 VSS.n2416 2.24304
R1443 VSS.n3372 VSS.n3370 2.24304
R1444 VSS.n2429 VSS.n2416 2.24304
R1445 VSS.n3372 VSS.n3371 2.24304
R1446 VSS.n3372 VSS.n2431 2.24304
R1447 VSS.n4841 VSS.n4825 2.24304
R1448 VSS.n4839 VSS.n0 2.24304
R1449 VSS.n4835 VSS.n0 2.24304
R1450 VSS.n4837 VSS.n4825 2.24304
R1451 VSS.n4833 VSS.n1 2.24304
R1452 VSS.n4829 VSS.n1 2.24304
R1453 VSS.n4831 VSS.n0 2.24304
R1454 VSS.n4827 VSS.n0 2.24304
R1455 VSS.n3949 VSS.n3904 2.24011
R1456 VSS.n3949 VSS.n3947 2.24011
R1457 VSS.n4164 VSS.n3729 2.24011
R1458 VSS.n4164 VSS.n3727 2.24011
R1459 VSS.n3795 VSS.n3723 2.24011
R1460 VSS.n3795 VSS.n2653 2.24011
R1461 VSS.n3728 VSS.n3726 2.24011
R1462 VSS.n3757 VSS.n3756 2.24011
R1463 VSS.n4133 VSS.n3772 2.24011
R1464 VSS.n3951 VSS.n3906 2.24011
R1465 VSS.n4169 VSS.n3721 2.24011
R1466 VSS.n3922 VSS.n3919 2.23777
R1467 VSS.n3920 VSS.n3769 2.23777
R1468 VSS.n3922 VSS.n3921 2.23777
R1469 VSS.n3877 VSS.n3876 2.23777
R1470 VSS.n3879 VSS.n3878 2.23777
R1471 VSS.n3876 VSS.n3871 2.23777
R1472 VSS.n1143 VSS.n1142 2.23644
R1473 VSS.n35 VSS.n34 2.23644
R1474 VSS.n1142 VSS.n38 2.23644
R1475 VSS.n39 VSS.n34 2.23644
R1476 VSS.n1142 VSS.n40 2.23644
R1477 VSS.n41 VSS.n34 2.23644
R1478 VSS.n1142 VSS.n42 2.23644
R1479 VSS.n43 VSS.n34 2.23644
R1480 VSS.n1142 VSS.n44 2.23644
R1481 VSS.n45 VSS.n34 2.23644
R1482 VSS.n1142 VSS.n46 2.23644
R1483 VSS.n47 VSS.n34 2.23644
R1484 VSS.n1142 VSS.n48 2.23644
R1485 VSS.n49 VSS.n34 2.23644
R1486 VSS.n1142 VSS.n50 2.23644
R1487 VSS.n51 VSS.n34 2.23644
R1488 VSS.n1142 VSS.n52 2.23644
R1489 VSS.n53 VSS.n34 2.23644
R1490 VSS.n1142 VSS.n54 2.23644
R1491 VSS.n55 VSS.n34 2.23644
R1492 VSS.n77 VSS.n56 2.23644
R1493 VSS.n1139 VSS.n67 2.23644
R1494 VSS.n77 VSS.n76 2.23644
R1495 VSS.n1139 VSS.n66 2.23644
R1496 VSS.n77 VSS.n75 2.23644
R1497 VSS.n1139 VSS.n65 2.23644
R1498 VSS.n77 VSS.n74 2.23644
R1499 VSS.n1139 VSS.n64 2.23644
R1500 VSS.n77 VSS.n73 2.23644
R1501 VSS.n1139 VSS.n63 2.23644
R1502 VSS.n77 VSS.n72 2.23644
R1503 VSS.n1139 VSS.n62 2.23644
R1504 VSS.n77 VSS.n71 2.23644
R1505 VSS.n1139 VSS.n61 2.23644
R1506 VSS.n77 VSS.n70 2.23644
R1507 VSS.n1139 VSS.n60 2.23644
R1508 VSS.n77 VSS.n69 2.23644
R1509 VSS.n1139 VSS.n59 2.23644
R1510 VSS.n77 VSS.n68 2.23644
R1511 VSS.n1139 VSS.n58 2.23644
R1512 VSS.n4305 VSS.n2622 2.16228
R1513 VSS.n5692 VSS.n1172 2.15282
R1514 VSS.n3522 VSS.n3517 2.12226
R1515 VSS.n3640 VSS.n3639 2.10421
R1516 VSS.n2707 VSS.n2706 2.10097
R1517 VSS.n4672 VSS.n2509 2.07167
R1518 VSS.n5301 VSS.n5300 2.01663
R1519 VSS.n5258 VSS.n5257 1.96906
R1520 VSS.n2514 VSS.n2092 1.94426
R1521 VSS.n3609 VSS.n3608 1.94426
R1522 VSS.n4194 VSS.n4193 1.91475
R1523 VSS.n4198 VSS.n4197 1.91081
R1524 VSS.n3257 VSS.n3256 1.89625
R1525 VSS.n5174 VSS.n2271 1.87995
R1526 VSS.n5334 VSS.n5333 1.81109
R1527 VSS.n2521 VSS.n2094 1.81109
R1528 VSS.n2184 VSS.n2180 1.81109
R1529 VSS.n2522 VSS.n2096 1.81109
R1530 VSS.n5439 VSS.n5438 1.80682
R1531 VSS.n2630 VSS 1.7864
R1532 VSS.n4203 VSS 1.7864
R1533 VSS.n5342 VSS.n5341 1.73383
R1534 VSS.n5342 VSS.n11 1.73383
R1535 VSS.n5409 VSS.n5408 1.73383
R1536 VSS.n5408 VSS.n5407 1.73383
R1537 VSS.n2525 VSS.n2098 1.73383
R1538 VSS.n2102 VSS.n2098 1.73383
R1539 VSS.n2086 VSS.n2083 1.73383
R1540 VSS.n2089 VSS.n2083 1.73383
R1541 VSS.n5687 VSS.n8 1.69455
R1542 VSS.n907 VSS.n906 1.66284
R1543 VSS.n5446 VSS.n5445 1.66212
R1544 VSS.n907 VSS.n221 1.64846
R1545 VSS.n5316 VSS.n5315 1.61108
R1546 VSS.n5306 VSS.n2192 1.61108
R1547 VSS.n4845 VSS.n4843 1.61108
R1548 VSS.n3562 VSS.n3561 1.59033
R1549 VSS.n3553 VSS.n2729 1.59033
R1550 VSS.n2728 VSS.n2723 1.59033
R1551 VSS.n2726 VSS.n2719 1.59033
R1552 VSS.n3518 VSS.n2715 1.59033
R1553 VSS.n3587 VSS.n3586 1.59033
R1554 VSS.n3650 VSS.n3623 1.59033
R1555 VSS.n3674 VSS.n3673 1.59033
R1556 VSS.n3664 VSS.n2241 1.59033
R1557 VSS.n2516 VSS.t40 1.57022
R1558 VSS.n2626 VSS.t7 1.57022
R1559 VSS.n2628 VSS.t12 1.57022
R1560 VSS.n2188 VSS.t44 1.57022
R1561 VSS.n2190 VSS.t1 1.57022
R1562 VSS.n4846 VSS.t10 1.57022
R1563 VSS.n3617 VSS.n2414 1.56129
R1564 VSS.n4217 VSS.n2627 1.52301
R1565 VSS.n3605 VSS.n2703 1.51243
R1566 VSS.n5432 DVSS 1.50997
R1567 VSS.n5428 DVSS 1.50997
R1568 VSS.n2181 DVSS 1.50997
R1569 VSS.n5338 DVSS 1.50997
R1570 VSS.n1772 VSS.n1762 1.50734
R1571 VSS.n1787 VSS.n1786 1.50734
R1572 VSS.n1726 VSS.n1724 1.50734
R1573 VSS.n1904 VSS.n1903 1.50734
R1574 VSS.n1702 VSS.n1700 1.50734
R1575 VSS.n1942 VSS.n1941 1.50734
R1576 VSS.n1989 VSS.n1988 1.50734
R1577 VSS.n1974 VSS.n1973 1.50734
R1578 VSS.n2021 VSS.n2020 1.50734
R1579 VSS.n2006 VSS.n2005 1.50734
R1580 VSS.n1628 VSS.n1618 1.50734
R1581 VSS.n1643 VSS.n1642 1.50734
R1582 VSS.n2937 VSS.n2925 1.5055
R1583 VSS.n5171 VSS.n5170 1.5055
R1584 VSS.n2937 VSS.n2936 1.5055
R1585 VSS.n5170 VSS.n2278 1.5055
R1586 VSS.n5329 VSS.n2113 1.50326
R1587 VSS.n4668 VSS.n4667 1.50326
R1588 VSS.n4513 VSS.n2568 1.50157
R1589 VSS.n4333 VSS.n4332 1.5005
R1590 VSS.n4335 VSS.n4334 1.5005
R1591 VSS.n4337 VSS.n4336 1.5005
R1592 VSS.n4339 VSS.n4338 1.5005
R1593 VSS.n4341 VSS.n4340 1.5005
R1594 VSS.n4343 VSS.n4342 1.5005
R1595 VSS.n4345 VSS.n4344 1.5005
R1596 VSS.n4347 VSS.n4346 1.5005
R1597 VSS.n4330 VSS.n2613 1.5005
R1598 VSS.n1641 VSS.n1634 1.5005
R1599 VSS.n2039 VSS.n2038 1.5005
R1600 VSS.n1632 VSS.n1626 1.5005
R1601 VSS.n2046 VSS.n2045 1.5005
R1602 VSS.n1627 VSS.n1623 1.5005
R1603 VSS.n1663 VSS.n1661 1.5005
R1604 VSS.n2010 VSS.n2009 1.5005
R1605 VSS.n1731 VSS.n1658 1.5005
R1606 VSS.n1730 VSS.n1651 1.5005
R1607 VSS.n2019 VSS.n2018 1.5005
R1608 VSS.n1688 VSS.n1686 1.5005
R1609 VSS.n1978 VSS.n1977 1.5005
R1610 VSS.n1737 VSS.n1683 1.5005
R1611 VSS.n1736 VSS.n1678 1.5005
R1612 VSS.n1987 VSS.n1986 1.5005
R1613 VSS.n1936 VSS.n1715 1.5005
R1614 VSS.n1938 VSS.n1708 1.5005
R1615 VSS.n1951 VSS.n1950 1.5005
R1616 VSS.n1706 VSS.n1703 1.5005
R1617 VSS.n1957 VSS.n1956 1.5005
R1618 VSS.n1898 VSS.n1757 1.5005
R1619 VSS.n1900 VSS.n1750 1.5005
R1620 VSS.n1913 VSS.n1912 1.5005
R1621 VSS.n1748 VSS.n1727 1.5005
R1622 VSS.n1919 VSS.n1918 1.5005
R1623 VSS.n1785 VSS.n1778 1.5005
R1624 VSS.n1874 VSS.n1873 1.5005
R1625 VSS.n1776 VSS.n1770 1.5005
R1626 VSS.n1881 VSS.n1880 1.5005
R1627 VSS.n1771 VSS.n1767 1.5005
R1628 VSS.n5706 VSS.n5705 1.5005
R1629 VSS.n21 VSS.n17 1.5005
R1630 VSS.n1151 VSS.n1150 1.5005
R1631 VSS.n1153 VSS.n1152 1.5005
R1632 VSS.n1155 VSS.n1154 1.5005
R1633 VSS.n1157 VSS.n1156 1.5005
R1634 VSS.n1159 VSS.n1158 1.5005
R1635 VSS.n1161 VSS.n1160 1.5005
R1636 VSS.n1163 VSS.n1162 1.5005
R1637 VSS.n1165 VSS.n1164 1.5005
R1638 VSS.n1167 VSS.n1166 1.5005
R1639 VSS.n1168 VSS.n31 1.5005
R1640 VSS.n5112 VSS.n5111 1.5005
R1641 VSS.n5110 VSS.n2275 1.5005
R1642 VSS.n5172 VSS.n5171 1.5005
R1643 VSS.n5114 VSS.n5113 1.5005
R1644 VSS.n5109 VSS.n2289 1.5005
R1645 VSS.n5108 VSS.n5107 1.5005
R1646 VSS.n5096 VSS.n2291 1.5005
R1647 VSS.n5095 VSS.n5094 1.5005
R1648 VSS.n5093 VSS.n5092 1.5005
R1649 VSS.n5091 VSS.n2301 1.5005
R1650 VSS.n5070 VSS.n2302 1.5005
R1651 VSS.n5072 VSS.n5071 1.5005
R1652 VSS.n5068 VSS.n5067 1.5005
R1653 VSS.n2313 VSS.n2312 1.5005
R1654 VSS.n5045 VSS.n5044 1.5005
R1655 VSS.n5043 VSS.n5042 1.5005
R1656 VSS.n2322 VSS.n2321 1.5005
R1657 VSS.n5026 VSS.n5025 1.5005
R1658 VSS.n5024 VSS.n2332 1.5005
R1659 VSS.n5023 VSS.n5022 1.5005
R1660 VSS.n2334 VSS.n2333 1.5005
R1661 VSS.n5002 VSS.n5001 1.5005
R1662 VSS.n5000 VSS.n4999 1.5005
R1663 VSS.n2343 VSS.n2342 1.5005
R1664 VSS.n4983 VSS.n4982 1.5005
R1665 VSS.n2354 VSS.n2353 1.5005
R1666 VSS.n4964 VSS.n4963 1.5005
R1667 VSS.n4966 VSS.n4965 1.5005
R1668 VSS.n4961 VSS.n2361 1.5005
R1669 VSS.n4960 VSS.n4959 1.5005
R1670 VSS.n4948 VSS.n2365 1.5005
R1671 VSS.n4947 VSS.n4946 1.5005
R1672 VSS.n4945 VSS.n4944 1.5005
R1673 VSS.n4943 VSS.n2375 1.5005
R1674 VSS.n4919 VSS.n2376 1.5005
R1675 VSS.n4921 VSS.n4920 1.5005
R1676 VSS.n4917 VSS.n4916 1.5005
R1677 VSS.n2387 VSS.n2386 1.5005
R1678 VSS.n4893 VSS.n4892 1.5005
R1679 VSS.n4891 VSS.n4890 1.5005
R1680 VSS.n2396 VSS.n2395 1.5005
R1681 VSS.n4874 VSS.n4873 1.5005
R1682 VSS.n2407 VSS.n2406 1.5005
R1683 VSS.n3224 VSS.n3223 1.5005
R1684 VSS.n3222 VSS.n3220 1.5005
R1685 VSS.n2808 VSS.n2807 1.5005
R1686 VSS.n3234 VSS.n3233 1.5005
R1687 VSS.n3236 VSS.n3235 1.5005
R1688 VSS.n2806 VSS.n2804 1.5005
R1689 VSS.n3188 VSS.n3187 1.5005
R1690 VSS.n3185 VSS.n2818 1.5005
R1691 VSS.n3184 VSS.n3183 1.5005
R1692 VSS.n2820 VSS.n2819 1.5005
R1693 VSS.n3167 VSS.n3166 1.5005
R1694 VSS.n3165 VSS.n3164 1.5005
R1695 VSS.n2829 VSS.n2828 1.5005
R1696 VSS.n3147 VSS.n3146 1.5005
R1697 VSS.n3145 VSS.n2839 1.5005
R1698 VSS.n3144 VSS.n3143 1.5005
R1699 VSS.n2841 VSS.n2840 1.5005
R1700 VSS.n3123 VSS.n3122 1.5005
R1701 VSS.n3120 VSS.n3119 1.5005
R1702 VSS.n2850 VSS.n2849 1.5005
R1703 VSS.n3103 VSS.n3102 1.5005
R1704 VSS.n3101 VSS.n3100 1.5005
R1705 VSS.n3099 VSS.n3098 1.5005
R1706 VSS.n3097 VSS.n3096 1.5005
R1707 VSS.n2862 VSS.n2861 1.5005
R1708 VSS.n3084 VSS.n3083 1.5005
R1709 VSS.n3082 VSS.n3081 1.5005
R1710 VSS.n2874 VSS.n2873 1.5005
R1711 VSS.n3050 VSS.n3049 1.5005
R1712 VSS.n3048 VSS.n3047 1.5005
R1713 VSS.n3046 VSS.n3045 1.5005
R1714 VSS.n3044 VSS.n3043 1.5005
R1715 VSS.n2885 VSS.n2884 1.5005
R1716 VSS.n3023 VSS.n3022 1.5005
R1717 VSS.n3021 VSS.n3020 1.5005
R1718 VSS.n2896 VSS.n2895 1.5005
R1719 VSS.n2996 VSS.n2995 1.5005
R1720 VSS.n2994 VSS.n2903 1.5005
R1721 VSS.n2993 VSS.n2992 1.5005
R1722 VSS.n2905 VSS.n2904 1.5005
R1723 VSS.n2976 VSS.n2975 1.5005
R1724 VSS.n2974 VSS.n2973 1.5005
R1725 VSS.n2951 VSS.n2916 1.5005
R1726 VSS.n2953 VSS.n2952 1.5005
R1727 VSS.n2950 VSS.n2949 1.5005
R1728 VSS.n2948 VSS.n2924 1.5005
R1729 VSS.n2930 VSS.n2925 1.5005
R1730 VSS.n5124 VSS.n5123 1.5005
R1731 VSS.n5122 VSS.n2278 1.5005
R1732 VSS.n2936 VSS.n2935 1.5005
R1733 VSS.n2934 VSS.n2933 1.5005
R1734 VSS.n2932 VSS.n2920 1.5005
R1735 VSS.n2958 VSS.n2957 1.5005
R1736 VSS.n2959 VSS.n2918 1.5005
R1737 VSS.n2968 VSS.n2967 1.5005
R1738 VSS.n2966 VSS.n2965 1.5005
R1739 VSS.n2964 VSS.n2963 1.5005
R1740 VSS.n2962 VSS.n2961 1.5005
R1741 VSS.n2901 VSS.n2900 1.5005
R1742 VSS.n3001 VSS.n3000 1.5005
R1743 VSS.n3002 VSS.n2898 1.5005
R1744 VSS.n3015 VSS.n3014 1.5005
R1745 VSS.n3013 VSS.n3012 1.5005
R1746 VSS.n3011 VSS.n3010 1.5005
R1747 VSS.n3009 VSS.n3008 1.5005
R1748 VSS.n3006 VSS.n3004 1.5005
R1749 VSS.n3005 VSS.n2878 1.5005
R1750 VSS.n3055 VSS.n3054 1.5005
R1751 VSS.n3056 VSS.n2876 1.5005
R1752 VSS.n3076 VSS.n3075 1.5005
R1753 VSS.n3074 VSS.n3073 1.5005
R1754 VSS.n3072 VSS.n3071 1.5005
R1755 VSS.n3070 VSS.n3069 1.5005
R1756 VSS.n3067 VSS.n3057 1.5005
R1757 VSS.n3066 VSS.n3065 1.5005
R1758 VSS.n3064 VSS.n3063 1.5005
R1759 VSS.n3062 VSS.n3061 1.5005
R1760 VSS.n3060 VSS.n3059 1.5005
R1761 VSS.n3128 VSS.n3127 1.5005
R1762 VSS.n3129 VSS.n2843 1.5005
R1763 VSS.n3137 VSS.n3136 1.5005
R1764 VSS.n3135 VSS.n3134 1.5005
R1765 VSS.n3133 VSS.n3132 1.5005
R1766 VSS.n3131 VSS.n3130 1.5005
R1767 VSS.n2831 VSS.n2824 1.5005
R1768 VSS.n3172 VSS.n3171 1.5005
R1769 VSS.n3173 VSS.n2822 1.5005
R1770 VSS.n3177 VSS.n3176 1.5005
R1771 VSS.n3175 VSS.n3174 1.5005
R1772 VSS.n2800 VSS.n2798 1.5005
R1773 VSS.n3241 VSS.n3240 1.5005
R1774 VSS.n2801 VSS.n2799 1.5005
R1775 VSS.n3204 VSS.n3203 1.5005
R1776 VSS.n3207 VSS.n3206 1.5005
R1777 VSS.n3208 VSS.n3199 1.5005
R1778 VSS.n3216 VSS.n3215 1.5005
R1779 VSS.n3214 VSS.n3213 1.5005
R1780 VSS.n3212 VSS.n3211 1.5005
R1781 VSS.n3210 VSS.n3209 1.5005
R1782 VSS.n2398 VSS.n2391 1.5005
R1783 VSS.n4898 VSS.n4897 1.5005
R1784 VSS.n4899 VSS.n2389 1.5005
R1785 VSS.n4911 VSS.n4910 1.5005
R1786 VSS.n4908 VSS.n4907 1.5005
R1787 VSS.n4906 VSS.n4905 1.5005
R1788 VSS.n4904 VSS.n4903 1.5005
R1789 VSS.n4902 VSS.n4900 1.5005
R1790 VSS.n2370 VSS.n2369 1.5005
R1791 VSS.n4953 VSS.n4952 1.5005
R1792 VSS.n4955 VSS.n4954 1.5005
R1793 VSS.n2358 VSS.n2357 1.5005
R1794 VSS.n4971 VSS.n4970 1.5005
R1795 VSS.n4973 VSS.n4972 1.5005
R1796 VSS.n4975 VSS.n2355 1.5005
R1797 VSS.n4977 VSS.n4976 1.5005
R1798 VSS.n4979 VSS.n4978 1.5005
R1799 VSS.n2345 VSS.n2338 1.5005
R1800 VSS.n5007 VSS.n5006 1.5005
R1801 VSS.n5008 VSS.n2336 1.5005
R1802 VSS.n5016 VSS.n5015 1.5005
R1803 VSS.n5014 VSS.n5013 1.5005
R1804 VSS.n5012 VSS.n5011 1.5005
R1805 VSS.n5010 VSS.n5009 1.5005
R1806 VSS.n2324 VSS.n2317 1.5005
R1807 VSS.n5050 VSS.n5049 1.5005
R1808 VSS.n5051 VSS.n2315 1.5005
R1809 VSS.n5062 VSS.n5061 1.5005
R1810 VSS.n5059 VSS.n5058 1.5005
R1811 VSS.n5057 VSS.n5056 1.5005
R1812 VSS.n5055 VSS.n2304 1.5005
R1813 VSS.n5054 VSS.n5053 1.5005
R1814 VSS.n2296 VSS.n2295 1.5005
R1815 VSS.n5101 VSS.n5100 1.5005
R1816 VSS.n5103 VSS.n5102 1.5005
R1817 VSS.n2286 VSS.n2285 1.5005
R1818 VSS.n5120 VSS.n5119 1.5005
R1819 VSS.n5121 VSS.n2284 1.5005
R1820 VSS.n5126 VSS.n5125 1.5005
R1821 VSS.n5118 VSS.n2283 1.5005
R1822 VSS.n5117 VSS.n5116 1.5005
R1823 VSS.n5105 VSS.n5104 1.5005
R1824 VSS.n2298 VSS.n2294 1.5005
R1825 VSS.n5099 VSS.n5098 1.5005
R1826 VSS.n5052 VSS.n2305 1.5005
R1827 VSS.n5090 VSS.n2304 1.5005
R1828 VSS.n5074 VSS.n2310 1.5005
R1829 VSS.n2316 VSS.n2309 1.5005
R1830 VSS.n5065 VSS.n5063 1.5005
R1831 VSS.n5048 VSS.n5047 1.5005
R1832 VSS.n2326 VSS.n2318 1.5005
R1833 VSS.n5040 VSS.n2325 1.5005
R1834 VSS.n5028 VSS.n2331 1.5005
R1835 VSS.n2337 VSS.n2330 1.5005
R1836 VSS.n5019 VSS.n5017 1.5005
R1837 VSS.n5005 VSS.n5004 1.5005
R1838 VSS.n2347 VSS.n2339 1.5005
R1839 VSS.n4997 VSS.n2346 1.5005
R1840 VSS.n4985 VSS.n2352 1.5005
R1841 VSS.n4974 VSS.n2351 1.5005
R1842 VSS.n2363 VSS.n2356 1.5005
R1843 VSS.n4969 VSS.n4968 1.5005
R1844 VSS.n4957 VSS.n4956 1.5005
R1845 VSS.n2372 VSS.n2368 1.5005
R1846 VSS.n4951 VSS.n4950 1.5005
R1847 VSS.n4901 VSS.n2379 1.5005
R1848 VSS.n4941 VSS.n2378 1.5005
R1849 VSS.n4923 VSS.n2384 1.5005
R1850 VSS.n2390 VSS.n2383 1.5005
R1851 VSS.n4914 VSS.n4912 1.5005
R1852 VSS.n4896 VSS.n4895 1.5005
R1853 VSS.n2400 VSS.n2392 1.5005
R1854 VSS.n4888 VSS.n2399 1.5005
R1855 VSS.n4876 VSS.n2405 1.5005
R1856 VSS.n3200 VSS.n2404 1.5005
R1857 VSS.n3226 VSS.n3217 1.5005
R1858 VSS.n3205 VSS.n2811 1.5005
R1859 VSS.n3231 VSS.n2810 1.5005
R1860 VSS.n3202 VSS.n3201 1.5005
R1861 VSS.n3239 VSS.n3238 1.5005
R1862 VSS.n3190 VSS.n2817 1.5005
R1863 VSS.n2823 VSS.n2816 1.5005
R1864 VSS.n3180 VSS.n3178 1.5005
R1865 VSS.n3170 VSS.n3169 1.5005
R1866 VSS.n2833 VSS.n2825 1.5005
R1867 VSS.n3162 VSS.n2832 1.5005
R1868 VSS.n3149 VSS.n2838 1.5005
R1869 VSS.n2844 VSS.n2837 1.5005
R1870 VSS.n3140 VSS.n3138 1.5005
R1871 VSS.n3126 VSS.n3125 1.5005
R1872 VSS.n2853 VSS.n2846 1.5005
R1873 VSS.n3117 VSS.n2852 1.5005
R1874 VSS.n3105 VSS.n2858 1.5005
R1875 VSS.n3058 VSS.n2857 1.5005
R1876 VSS.n3068 VSS.n2866 1.5005
R1877 VSS.n3094 VSS.n2864 1.5005
R1878 VSS.n3086 VSS.n2871 1.5005
R1879 VSS.n2877 VSS.n2870 1.5005
R1880 VSS.n3079 VSS.n3077 1.5005
R1881 VSS.n3053 VSS.n3052 1.5005
R1882 VSS.n3036 VSS.n2879 1.5005
R1883 VSS.n3007 VSS.n2888 1.5005
R1884 VSS.n3041 VSS.n2887 1.5005
R1885 VSS.n3025 VSS.n2893 1.5005
R1886 VSS.n2899 VSS.n2892 1.5005
R1887 VSS.n3018 VSS.n3016 1.5005
R1888 VSS.n2999 VSS.n2998 1.5005
R1889 VSS.n2908 VSS.n2901 1.5005
R1890 VSS.n2990 VSS.n2907 1.5005
R1891 VSS.n2978 VSS.n2913 1.5005
R1892 VSS.n2919 VSS.n2912 1.5005
R1893 VSS.n2971 VSS.n2969 1.5005
R1894 VSS.n2956 VSS.n2955 1.5005
R1895 VSS.n2928 VSS.n2921 1.5005
R1896 VSS.n2946 VSS.n2927 1.5005
R1897 VSS.n5126 VSS.n2276 1.5005
R1898 VSS.n2290 VSS.n2283 1.5005
R1899 VSS.n5116 VSS.n5115 1.5005
R1900 VSS.n5106 VSS.n5105 1.5005
R1901 VSS.n2298 VSS.n2292 1.5005
R1902 VSS.n5098 VSS.n5097 1.5005
R1903 VSS.n2305 VSS.n2300 1.5005
R1904 VSS.n5091 VSS.n5090 1.5005
R1905 VSS.n5074 VSS.n5073 1.5005
R1906 VSS.n2311 VSS.n2309 1.5005
R1907 VSS.n5066 VSS.n5065 1.5005
R1908 VSS.n5047 VSS.n5046 1.5005
R1909 VSS.n2326 VSS.n2320 1.5005
R1910 VSS.n5041 VSS.n5040 1.5005
R1911 VSS.n5028 VSS.n5027 1.5005
R1912 VSS.n5021 VSS.n2330 1.5005
R1913 VSS.n5020 VSS.n5019 1.5005
R1914 VSS.n5004 VSS.n5003 1.5005
R1915 VSS.n2347 VSS.n2341 1.5005
R1916 VSS.n4998 VSS.n4997 1.5005
R1917 VSS.n4985 VSS.n4984 1.5005
R1918 VSS.n4962 VSS.n2351 1.5005
R1919 VSS.n2364 VSS.n2363 1.5005
R1920 VSS.n4968 VSS.n4967 1.5005
R1921 VSS.n4958 VSS.n4957 1.5005
R1922 VSS.n2372 VSS.n2366 1.5005
R1923 VSS.n4950 VSS.n4949 1.5005
R1924 VSS.n2379 VSS.n2374 1.5005
R1925 VSS.n4942 VSS.n4941 1.5005
R1926 VSS.n4923 VSS.n4922 1.5005
R1927 VSS.n2385 VSS.n2383 1.5005
R1928 VSS.n4915 VSS.n4914 1.5005
R1929 VSS.n4895 VSS.n4894 1.5005
R1930 VSS.n2400 VSS.n2394 1.5005
R1931 VSS.n4889 VSS.n4888 1.5005
R1932 VSS.n4876 VSS.n4875 1.5005
R1933 VSS.n3221 VSS.n2404 1.5005
R1934 VSS.n3226 VSS.n3225 1.5005
R1935 VSS.n3219 VSS.n2811 1.5005
R1936 VSS.n3232 VSS.n3231 1.5005
R1937 VSS.n3201 VSS.n2805 1.5005
R1938 VSS.n3238 VSS.n3237 1.5005
R1939 VSS.n3190 VSS.n3189 1.5005
R1940 VSS.n3182 VSS.n2816 1.5005
R1941 VSS.n3181 VSS.n3180 1.5005
R1942 VSS.n3169 VSS.n3168 1.5005
R1943 VSS.n2833 VSS.n2827 1.5005
R1944 VSS.n3163 VSS.n3162 1.5005
R1945 VSS.n3149 VSS.n3148 1.5005
R1946 VSS.n3142 VSS.n2837 1.5005
R1947 VSS.n3141 VSS.n3140 1.5005
R1948 VSS.n3125 VSS.n3124 1.5005
R1949 VSS.n2853 VSS.n2848 1.5005
R1950 VSS.n3118 VSS.n3117 1.5005
R1951 VSS.n3105 VSS.n3104 1.5005
R1952 VSS.n2859 VSS.n2857 1.5005
R1953 VSS.n2866 VSS.n2860 1.5005
R1954 VSS.n3095 VSS.n3094 1.5005
R1955 VSS.n3086 VSS.n3085 1.5005
R1956 VSS.n2872 VSS.n2870 1.5005
R1957 VSS.n3080 VSS.n3079 1.5005
R1958 VSS.n3052 VSS.n3051 1.5005
R1959 VSS.n3036 VSS.n2881 1.5005
R1960 VSS.n2888 VSS.n2883 1.5005
R1961 VSS.n3042 VSS.n3041 1.5005
R1962 VSS.n3025 VSS.n3024 1.5005
R1963 VSS.n2894 VSS.n2892 1.5005
R1964 VSS.n3019 VSS.n3018 1.5005
R1965 VSS.n2998 VSS.n2997 1.5005
R1966 VSS.n2908 VSS.n2903 1.5005
R1967 VSS.n2991 VSS.n2990 1.5005
R1968 VSS.n2978 VSS.n2977 1.5005
R1969 VSS.n2914 VSS.n2912 1.5005
R1970 VSS.n2972 VSS.n2971 1.5005
R1971 VSS.n2955 VSS.n2954 1.5005
R1972 VSS.n2928 VSS.n2923 1.5005
R1973 VSS.n2947 VSS.n2946 1.5005
R1974 VSS.n5182 VSS.n5181 1.5005
R1975 VSS.n3842 VSS.n2567 1.5005
R1976 VSS.n3844 VSS.n3843 1.5005
R1977 VSS.n3846 VSS.n3845 1.5005
R1978 VSS.n3848 VSS.n3847 1.5005
R1979 VSS.n3850 VSS.n3849 1.5005
R1980 VSS.n3852 VSS.n3851 1.5005
R1981 VSS.n3854 VSS.n3853 1.5005
R1982 VSS.n3856 VSS.n3855 1.5005
R1983 VSS.n3858 VSS.n3857 1.5005
R1984 VSS.n4329 VSS.n2615 1.49818
R1985 VSS.n3607 VSS.n3606 1.49138
R1986 VSS.n4672 VSS.n4671 1.48621
R1987 VSS.n4123 VSS.n4122 1.44688
R1988 VSS.n3882 VSS.n3881 1.44688
R1989 VSS.n5414 VSS.n5413 1.39741
R1990 VSS.n5453 VSS.n5452 1.38664
R1991 VSS.n3840 VSS.n3780 1.35477
R1992 VSS.n4069 VSS.n3781 1.35477
R1993 VSS.n5255 DVSS 1.35085
R1994 VSS.n3614 VSS.n2701 1.328
R1995 VSS.n3538 VSS.n3533 1.31286
R1996 VSS.n3600 VSS.n3599 1.31286
R1997 VSS.n2695 VSS.n2688 1.31286
R1998 VSS.n2244 VSS.n2242 1.31286
R1999 VSS.n2185 VSS.n2184 1.3005
R2000 VSS.n5333 VSS.n5332 1.3005
R2001 VSS.n2522 VSS.n2511 1.3005
R2002 VSS.n2521 VSS.n2510 1.3005
R2003 VSS.n4849 VSS.n4848 1.3005
R2004 VSS.n5308 VSS.n5307 1.3005
R2005 VSS.n5313 VSS.n5312 1.3005
R2006 VSS.n4216 VSS.n4215 1.3005
R2007 VSS.n4306 VSS.n4305 1.3005
R2008 VSS.n3254 VSS 1.28985
R2009 VSS.n5351 VSS.n2173 1.26649
R2010 VSS.n3568 VSS.n3567 1.25594
R2011 VSS.n3651 VSS.n3624 1.25594
R2012 DVSS VSS.n4206 1.23516
R2013 VSS.n4206 DVSS 1.23404
R2014 VSS.n2087 VSS.n2086 1.23176
R2015 VSS.n5341 VSS.n2174 1.23176
R2016 VSS.n5410 VSS.n5409 1.23176
R2017 VSS.n2526 VSS.n2525 1.23176
R2018 VSS.n4750 VSS.n2189 1.19925
R2019 VSS.n5257 VSS.n5256 1.16402
R2020 VSS.n2084 VSS.n2082 1.15745
R2021 VSS.n3604 VSS.n3603 1.15606
R2022 VSS.n5424 VSS.n5423 1.15606
R2023 VSS.n5418 VSS.n5417 1.15606
R2024 VSS.n4192 VSS.n4191 1.13009
R2025 VSS.n3639 VSS.n2238 1.10843
R2026 VSS.n3621 VSS.n2695 1.10563
R2027 VSS.n2242 VSS.n2240 1.10563
R2028 VSS.n3533 VSS.n3532 1.10563
R2029 VSS.n3601 VSS.n3600 1.10563
R2030 VSS.n4195 VSS.t49 1.0925
R2031 VSS.n3527 VSS.t19 1.0925
R2032 VSS.n2731 VSS.t33 1.0925
R2033 VSS.n2731 VSS.t26 1.0925
R2034 VSS.n2791 VSS.t28 1.0925
R2035 VSS.n2791 VSS.t21 1.0925
R2036 VSS.n2793 VSS.t31 1.0925
R2037 VSS.n2631 VSS.t14 1.0925
R2038 VSS.n2175 VSS.n2113 1.08844
R2039 VSS.n5403 VSS.n2113 1.08844
R2040 VSS.n4667 VSS.n4666 1.08844
R2041 VSS.n4667 VSS.n2088 1.08844
R2042 VSS.n5441 VSS.n2088 1.0805
R2043 VSS.n5348 VSS.n2175 1.0805
R2044 VSS.n5404 VSS.n5403 1.0805
R2045 VSS.n4666 VSS.n2530 1.0805
R2046 VSS.n5257 VSS.n2238 1.07932
R2047 VSS.n2077 VSS.n1591 1.07349
R2048 VSS.n4193 VSS.n2637 1.07241
R2049 VSS.n3720 VSS.n3719 1.05604
R2050 VSS.n2519 VSS.n2518 1.05029
R2051 VSS.n3252 VSS.n2795 1.0405
R2052 VSS.n2796 VSS.n2795 1.0405
R2053 VSS.n3611 VSS.n3610 1.0405
R2054 VSS.n3616 VSS.n2698 1.0405
R2055 VSS.n2698 VSS.n2697 1.0405
R2056 VSS.n2413 VSS.n2412 1.0405
R2057 VSS.n2412 VSS.n2411 1.0405
R2058 VSS.n5339 VSS.n5338 1.0405
R2059 VSS.n5339 VSS.n2176 1.0405
R2060 VSS.n2181 VSS.n2110 1.0405
R2061 VSS.n2112 VSS.n2110 1.0405
R2062 VSS.n5428 VSS.n5427 1.0405
R2063 VSS.n5427 VSS.n5426 1.0405
R2064 VSS.n5433 VSS.n5432 1.0405
R2065 VSS.n5434 VSS.n5433 1.0405
R2066 VSS.n2512 VSS.t22 1.0405
R2067 VSS.n2796 VSS.t4 1.00732
R2068 VSS.t16 VSS.n3611 1.00732
R2069 VSS.t2 VSS.n2697 1.00732
R2070 VSS.t36 VSS.n2411 1.00732
R2071 VSS.n3624 VSS.n2239 1.00517
R2072 VSS.n3567 VSS.n2725 1.00517
R2073 VSS VSS.n3522 1.00241
R2074 VSS.n3610 VSS.n3609 0.996088
R2075 VSS.n2514 VSS.n2512 0.996088
R2076 VSS.n5256 VSS.n5252 0.992621
R2077 VSS.n5442 DVSS 0.972907
R2078 VSS.n5349 DVSS 0.972907
R2079 VSS.n2108 DVSS 0.972907
R2080 VSS.n5443 VSS.n2087 0.971611
R2081 VSS.n5350 VSS.n2174 0.971611
R2082 VSS.n5411 VSS.n5410 0.971611
R2083 VSS.n2527 VSS.n2526 0.971611
R2084 VSS.n3522 VSS.n3521 0.945955
R2085 VSS.n4851 VSS.n4850 0.945955
R2086 VSS.n2189 VSS.n2111 0.945955
R2087 VSS.n5327 VSS.n5326 0.945955
R2088 VSS.n5422 VSS.n5421 0.945955
R2089 VSS.n2529 DVSS 0.92317
R2090 VSS.n3361 VSS.n7 0.922809
R2091 VSS.n5715 VSS.n5714 0.922714
R2092 VSS.n2766 VSS.n2765 0.922457
R2093 VSS.n4237 VSS.n1291 0.922457
R2094 VSS.n4202 VSS.n4201 0.910322
R2095 VSS.n1587 VSS.n1296 0.902282
R2096 VSS.n1588 VSS.n1587 0.902198
R2097 VSS.n1588 VSS.n1297 0.902161
R2098 VSS.n1297 VSS.n1296 0.901878
R2099 VSS.n5182 VSS.n2271 0.882658
R2100 VSS.n1591 VSS.n1590 0.879171
R2101 VSS.n5695 VSS.n1169 0.879171
R2102 VSS.n5353 VSS.n5352 0.875955
R2103 VSS.n5402 VSS.n5401 0.875955
R2104 VSS.n4665 VSS.n4664 0.875955
R2105 VSS.n3681 VSS.n3680 0.875366
R2106 VSS.n3640 VSS.n2696 0.875366
R2107 VSS.n5259 VSS.n5258 0.875366
R2108 VSS.n4197 VSS.n2633 0.873402
R2109 VSS.n1169 VSS.n1168 0.870066
R2110 VSS.n3564 VSS.n2730 0.867167
R2111 VSS.n3520 VSS.n3519 0.867167
R2112 VSS.n3678 VSS.n3622 0.867167
R2113 VSS.n5262 VSS.n5261 0.867167
R2114 VSS.n4863 VSS.n2413 0.843937
R2115 VSS.n3617 VSS.n3616 0.843937
R2116 VSS.n3252 VSS.n3251 0.843937
R2117 VSS.n3639 VSS.n2694 0.827218
R2118 VSS.n1145 VSS.n1144 0.820816
R2119 VSS.n2701 VSS.n2414 0.815237
R2120 VSS.n4529 VSS.n2088 0.803519
R2121 VSS.n5321 VSS.n2175 0.803519
R2122 VSS.n5403 VSS.n5402 0.803519
R2123 VSS.n4666 VSS.n4665 0.803519
R2124 VSS.n5352 DVSS 0.801151
R2125 VSS.n5437 VSS.n2090 0.8005
R2126 VSS.n4309 VSS.n2623 0.796907
R2127 VSS.n4313 VSS.n2623 0.796907
R2128 VSS.n4313 VSS.n2621 0.796907
R2129 VSS.n4317 VSS.n2621 0.796907
R2130 VSS.n4317 VSS.n2619 0.796907
R2131 VSS.n4321 VSS.n2619 0.796907
R2132 VSS.n4321 VSS.n2196 0.796907
R2133 VSS.n5299 VSS.n2196 0.796907
R2134 VSS.n5299 VSS.n2197 0.796907
R2135 VSS.n4851 VSS 0.78605
R2136 VSS.n5253 DVSS 0.783069
R2137 VSS.n5254 DVSS 0.783069
R2138 VSS.n3866 VSS.n3865 0.778288
R2139 VSS.n4574 VSS.n2103 0.774059
R2140 VSS.n2173 VSS.n2172 0.752663
R2141 VSS.n4860 VSS 0.751638
R2142 VSS.n3881 VSS.n3782 0.7505
R2143 VSS.n4124 VSS.n4123 0.7505
R2144 DVSS VSS.n4192 0.746344
R2145 VSS.n282 VSS.n122 0.745113
R2146 VSS.n824 VSS.n305 0.745113
R2147 VSS.n751 VSS.n330 0.745113
R2148 VSS.n3786 VSS.n3785 0.743357
R2149 VSS.n3785 VSS.n3777 0.743357
R2150 VSS.n4067 VSS.n3776 0.743357
R2151 VSS.n3779 VSS.n3776 0.743357
R2152 VSS.n3885 VSS.n3884 0.743357
R2153 VSS.n3884 VSS.n3779 0.743357
R2154 VSS.n3822 VSS.n3775 0.743357
R2155 VSS.n3777 VSS.n3775 0.743357
R2156 VSS.n283 VSS.n282 0.736857
R2157 VSS.n825 VSS.n824 0.736857
R2158 VSS.n751 VSS.n750 0.736857
R2159 VSS.n3870 VSS.n3869 0.735937
R2160 VSS.n4121 VSS.n4120 0.735937
R2161 VSS.n5444 VSS.n2084 0.7304
R2162 VSS.n3682 VSS.n3681 0.71546
R2163 VSS.n3641 VSS.n3640 0.71546
R2164 VSS.n5258 VSS.n5250 0.71546
R2165 VSS.n2530 VSS.n2529 0.707265
R2166 VSS.n5334 VSS.n2182 0.693432
R2167 VSS.n2180 VSS.n2179 0.693432
R2168 VSS.n2097 VSS.n2096 0.693432
R2169 VSS.n2094 VSS.n2093 0.693432
R2170 VSS.n5429 VSS.n2096 0.682241
R2171 VSS.n5335 VSS.n5334 0.682241
R2172 VSS.n5337 VSS.n2180 0.682241
R2173 VSS.n5431 VSS.n2094 0.682241
R2174 VSS.n4329 VSS.n4328 0.666308
R2175 VSS.n5296 VSS.n5295 0.66242
R2176 VSS.n5442 VSS.n5441 0.662265
R2177 VSS.n5349 VSS.n5348 0.662265
R2178 VSS.n5404 VSS.n2108 0.662265
R2179 VSS.n4328 VSS.n2616 0.64762
R2180 VSS.n5254 VSS.n5253 0.646382
R2181 VSS.n1773 VSS.n1769 0.643357
R2182 VSS.n1879 VSS.n1878 0.643357
R2183 VSS.n1876 VSS.n1875 0.643357
R2184 VSS.n1775 VSS.n1774 0.643357
R2185 VSS.n1917 VSS.n1916 0.643357
R2186 VSS.n1915 VSS.n1914 0.643357
R2187 VSS.n1899 VSS.n1747 0.643357
R2188 VSS.n1902 VSS.n1901 0.643357
R2189 VSS.n1955 VSS.n1954 0.643357
R2190 VSS.n1953 VSS.n1952 0.643357
R2191 VSS.n1937 VSS.n1705 0.643357
R2192 VSS.n1940 VSS.n1939 0.643357
R2193 VSS.n1677 VSS.n1676 0.643357
R2194 VSS.n1739 VSS.n1738 0.643357
R2195 VSS.n1687 VSS.n1685 0.643357
R2196 VSS.n1976 VSS.n1975 0.643357
R2197 VSS.n1650 VSS.n1649 0.643357
R2198 VSS.n1733 VSS.n1732 0.643357
R2199 VSS.n1662 VSS.n1660 0.643357
R2200 VSS.n2008 VSS.n2007 0.643357
R2201 VSS.n1629 VSS.n1625 0.643357
R2202 VSS.n2044 VSS.n2043 0.643357
R2203 VSS.n2041 VSS.n2040 0.643357
R2204 VSS.n1631 VSS.n1630 0.643357
R2205 VSS.n4217 VSS.n4216 0.634889
R2206 VSS.n2101 DVSS 0.621687
R2207 VSS.n5419 DVSS 0.621687
R2208 VSS.n5324 DVSS 0.621687
R2209 VSS.n5323 DVSS 0.621687
R2210 VSS.n5255 VSS.n5254 0.618588
R2211 VSS.n5177 VSS.n5176 0.612265
R2212 VSS.n5295 DVSS 0.600908
R2213 VSS.n5271 VSS.n2231 0.588678
R2214 VSS.n4864 VSS.n4863 0.585632
R2215 VSS.n3618 VSS.n3617 0.585632
R2216 VSS.n3251 VSS.n3250 0.585632
R2217 VSS.n3679 VSS.n2695 0.584525
R2218 VSS.n5260 VSS.n2242 0.584525
R2219 VSS.n3563 VSS.n3533 0.584525
R2220 VSS.n3600 VSS.n2708 0.584525
R2221 VSS.n2931 VSS.n2408 0.578278
R2222 VSS.n2409 DVSS 0.578278
R2223 VSS.n2409 VSS.n2274 0.578278
R2224 VSS.n5271 VSS.n5270 0.578278
R2225 VSS.n5272 VSS.n2210 0.578278
R2226 VSS.n5273 VSS.n2208 0.578278
R2227 VSS.n5274 VSS.n2211 0.578278
R2228 VSS.n5275 VSS.n2207 0.578278
R2229 VSS.n5276 VSS.n2212 0.578278
R2230 VSS.n5277 VSS.n2206 0.578278
R2231 VSS.n5278 VSS.n2213 0.578278
R2232 VSS.n5279 VSS.n2205 0.578278
R2233 VSS.n5280 VSS.n2214 0.578278
R2234 VSS.n5285 VSS.n5284 0.578278
R2235 VSS.n5287 VSS.n5286 0.578278
R2236 VSS.n5297 VSS.n2197 0.578278
R2237 VSS.n2197 VSS.n2195 0.578278
R2238 VSS.n5300 VSS.n5299 0.578278
R2239 VSS.n2196 VSS.n2194 0.578278
R2240 VSS.n4322 VSS.n4321 0.578278
R2241 VSS.n2619 VSS.n2618 0.578278
R2242 VSS.n4317 VSS.n4316 0.578278
R2243 VSS.n4315 VSS.n2621 0.578278
R2244 VSS.n4314 VSS.n4313 0.578278
R2245 VSS.n4307 VSS.n2623 0.578278
R2246 VSS.n4309 VSS.n4308 0.578278
R2247 VSS.n5299 VSS.n5298 0.578278
R2248 VSS.n2198 VSS.n2196 0.578278
R2249 VSS.n4321 VSS.n4320 0.578278
R2250 VSS.n4319 VSS.n2619 0.578278
R2251 VSS.n4318 VSS.n4317 0.578278
R2252 VSS.n2621 VSS.n2620 0.578278
R2253 VSS.n4313 VSS.n4312 0.578278
R2254 VSS.n4311 VSS.n2623 0.578278
R2255 VSS.n4310 VSS.n4309 0.578278
R2256 VSS.n4863 VSS.n4862 0.563
R2257 VSS.n5310 VSS.n2189 0.557079
R2258 VSS.n3615 VSS.n3614 0.557079
R2259 VSS.n5421 VSS.n5420 0.557079
R2260 VSS.n5326 VSS.n5325 0.557079
R2261 VSS.n3606 VSS.n3604 0.557079
R2262 VSS.n5315 VSS.n5313 0.553108
R2263 VSS.n5308 VSS.n2192 0.553108
R2264 VSS.n4848 VSS.n4845 0.553108
R2265 VSS.n2706 VSS.n2705 0.549281
R2266 VSS.n3526 VSS.n3524 0.545794
R2267 VSS.n5438 VSS.n5437 0.545794
R2268 VSS.n5443 VSS.n5442 0.545794
R2269 VSS.n5351 VSS.n5350 0.545794
R2270 VSS.n5350 VSS.n5349 0.545794
R2271 VSS.n5411 VSS.n2108 0.545794
R2272 VSS.n5412 VSS.n5411 0.545794
R2273 VSS.n2527 VSS.n2107 0.545794
R2274 VSS.n3679 VSS.n3678 0.545794
R2275 VSS.n5261 VSS.n5260 0.545794
R2276 VSS.n3519 VSS.n2708 0.545794
R2277 VSS.n3564 VSS.n3563 0.545794
R2278 VSS.n5438 DVSS 0.544093
R2279 VSS.n5436 DVSS 0.544093
R2280 VSS.n5437 DVSS 0.544018
R2281 VSS.n3258 VSS.n3257 0.543147
R2282 VSS.n5322 VSS.n5321 0.533549
R2283 VSS.n3870 VSS.n3786 0.5255
R2284 VSS.n4121 VSS.n3885 0.5255
R2285 VSS.n3250 VSS.n3249 0.5205
R2286 VSS.n3619 VSS.n3618 0.5205
R2287 VSS.n4865 VSS.n4864 0.5205
R2288 VSS.n4304 VSS.n2626 0.519124
R2289 VSS.n2629 VSS.n2628 0.519124
R2290 VSS.n5311 VSS.n2188 0.519124
R2291 VSS.n5309 VSS.n2190 0.519124
R2292 VSS.n4847 VSS.n4846 0.519124
R2293 VSS.n2944 VSS.n2939 0.5005
R2294 VSS.n2943 VSS.n2940 0.5005
R2295 VSS.n2942 VSS.n2941 0.5005
R2296 VSS.n2911 VSS.n2910 0.5005
R2297 VSS.n2981 VSS.n2980 0.5005
R2298 VSS.n2982 VSS.n2909 0.5005
R2299 VSS.n2988 VSS.n2983 0.5005
R2300 VSS.n2987 VSS.n2984 0.5005
R2301 VSS.n2986 VSS.n2985 0.5005
R2302 VSS.n2891 VSS.n2890 0.5005
R2303 VSS.n3028 VSS.n3027 0.5005
R2304 VSS.n3029 VSS.n2889 0.5005
R2305 VSS.n3039 VSS.n3030 0.5005
R2306 VSS.n3038 VSS.n3031 0.5005
R2307 VSS.n3035 VSS.n3032 0.5005
R2308 VSS.n3034 VSS.n3033 0.5005
R2309 VSS.n2869 VSS.n2868 0.5005
R2310 VSS.n3089 VSS.n3088 0.5005
R2311 VSS.n3090 VSS.n2867 0.5005
R2312 VSS.n3092 VSS.n3091 0.5005
R2313 VSS.n2856 VSS.n2855 0.5005
R2314 VSS.n3108 VSS.n3107 0.5005
R2315 VSS.n3109 VSS.n2854 0.5005
R2316 VSS.n3115 VSS.n3110 0.5005
R2317 VSS.n3114 VSS.n3111 0.5005
R2318 VSS.n3113 VSS.n3112 0.5005
R2319 VSS.n2836 VSS.n2835 0.5005
R2320 VSS.n3152 VSS.n3151 0.5005
R2321 VSS.n3153 VSS.n2834 0.5005
R2322 VSS.n3160 VSS.n3154 0.5005
R2323 VSS.n3159 VSS.n3155 0.5005
R2324 VSS.n3158 VSS.n3157 0.5005
R2325 VSS.n3156 VSS.n2814 0.5005
R2326 VSS.n3192 VSS.n2815 0.5005
R2327 VSS.n3193 VSS.n2813 0.5005
R2328 VSS.n3195 VSS.n3194 0.5005
R2329 VSS.n3196 VSS.n2812 0.5005
R2330 VSS.n3229 VSS.n3197 0.5005
R2331 VSS.n3228 VSS.n3198 0.5005
R2332 VSS.n2403 VSS.n2402 0.5005
R2333 VSS.n4879 VSS.n4878 0.5005
R2334 VSS.n4880 VSS.n2401 0.5005
R2335 VSS.n4886 VSS.n4881 0.5005
R2336 VSS.n4885 VSS.n4882 0.5005
R2337 VSS.n4884 VSS.n4883 0.5005
R2338 VSS.n2382 VSS.n2381 0.5005
R2339 VSS.n4926 VSS.n4925 0.5005
R2340 VSS.n4927 VSS.n2380 0.5005
R2341 VSS.n4939 VSS.n4928 0.5005
R2342 VSS.n4938 VSS.n4929 0.5005
R2343 VSS.n4937 VSS.n4930 0.5005
R2344 VSS.n4936 VSS.n4931 0.5005
R2345 VSS.n4935 VSS.n4932 0.5005
R2346 VSS.n4934 VSS.n4933 0.5005
R2347 VSS.n2350 VSS.n2349 0.5005
R2348 VSS.n4988 VSS.n4987 0.5005
R2349 VSS.n4989 VSS.n2348 0.5005
R2350 VSS.n4995 VSS.n4990 0.5005
R2351 VSS.n4994 VSS.n4991 0.5005
R2352 VSS.n4993 VSS.n4992 0.5005
R2353 VSS.n2329 VSS.n2328 0.5005
R2354 VSS.n5031 VSS.n5030 0.5005
R2355 VSS.n5032 VSS.n2327 0.5005
R2356 VSS.n5038 VSS.n5033 0.5005
R2357 VSS.n5037 VSS.n5034 0.5005
R2358 VSS.n5036 VSS.n5035 0.5005
R2359 VSS.n2308 VSS.n2307 0.5005
R2360 VSS.n5077 VSS.n5076 0.5005
R2361 VSS.n5078 VSS.n2306 0.5005
R2362 VSS.n5088 VSS.n5079 0.5005
R2363 VSS.n5087 VSS.n5080 0.5005
R2364 VSS.n5086 VSS.n5081 0.5005
R2365 VSS.n5085 VSS.n5082 0.5005
R2366 VSS.n5084 VSS.n5083 0.5005
R2367 VSS.n2282 VSS.n2281 0.5005
R2368 VSS.n5129 VSS.n5128 0.5005
R2369 VSS.n5130 VSS.n2280 0.5005
R2370 VSS.n5168 VSS.n5131 0.5005
R2371 VSS.n5167 VSS.n5132 0.5005
R2372 VSS.n5166 VSS.n5133 0.5005
R2373 VSS.n5136 VSS.n5134 0.5005
R2374 VSS.n5162 VSS.n5137 0.5005
R2375 VSS.n5161 VSS.n5138 0.5005
R2376 VSS.n5141 VSS.n5139 0.5005
R2377 VSS.n5157 VSS.n5142 0.5005
R2378 VSS.n5156 VSS.n5143 0.5005
R2379 VSS.n5155 VSS.n5144 0.5005
R2380 VSS.n5146 VSS.n5145 0.5005
R2381 VSS.n5151 VSS.n5147 0.5005
R2382 VSS.n5150 VSS.n5148 0.5005
R2383 VSS.n5163 VSS.n5162 0.5005
R2384 VSS.n5164 VSS.n5134 0.5005
R2385 VSS.n5166 VSS.n5165 0.5005
R2386 VSS.n5167 VSS.n2279 0.5005
R2387 VSS.n5169 VSS.n5168 0.5005
R2388 VSS.n2280 VSS.n2277 0.5005
R2389 VSS.n5128 VSS.n5127 0.5005
R2390 VSS.n2288 VSS.n2282 0.5005
R2391 VSS.n5084 VSS.n2287 0.5005
R2392 VSS.n5085 VSS.n2293 0.5005
R2393 VSS.n5086 VSS.n2299 0.5005
R2394 VSS.n5087 VSS.n2297 0.5005
R2395 VSS.n5089 VSS.n5088 0.5005
R2396 VSS.n2306 VSS.n2303 0.5005
R2397 VSS.n5076 VSS.n5075 0.5005
R2398 VSS.n5064 VSS.n2308 0.5005
R2399 VSS.n5036 VSS.n2314 0.5005
R2400 VSS.n5037 VSS.n2319 0.5005
R2401 VSS.n5039 VSS.n5038 0.5005
R2402 VSS.n2327 VSS.n2323 0.5005
R2403 VSS.n5030 VSS.n5029 0.5005
R2404 VSS.n5018 VSS.n2329 0.5005
R2405 VSS.n4993 VSS.n2335 0.5005
R2406 VSS.n4994 VSS.n2340 0.5005
R2407 VSS.n4996 VSS.n4995 0.5005
R2408 VSS.n2348 VSS.n2344 0.5005
R2409 VSS.n4987 VSS.n4986 0.5005
R2410 VSS.n2362 VSS.n2350 0.5005
R2411 VSS.n4934 VSS.n2360 0.5005
R2412 VSS.n4935 VSS.n2359 0.5005
R2413 VSS.n4936 VSS.n2367 0.5005
R2414 VSS.n4937 VSS.n2373 0.5005
R2415 VSS.n4938 VSS.n2371 0.5005
R2416 VSS.n4940 VSS.n4939 0.5005
R2417 VSS.n2380 VSS.n2377 0.5005
R2418 VSS.n4925 VSS.n4924 0.5005
R2419 VSS.n4913 VSS.n2382 0.5005
R2420 VSS.n4884 VSS.n2388 0.5005
R2421 VSS.n4885 VSS.n2393 0.5005
R2422 VSS.n4887 VSS.n4886 0.5005
R2423 VSS.n2401 VSS.n2397 0.5005
R2424 VSS.n4878 VSS.n4877 0.5005
R2425 VSS.n3218 VSS.n2403 0.5005
R2426 VSS.n3228 VSS.n3227 0.5005
R2427 VSS.n3230 VSS.n3229 0.5005
R2428 VSS.n2812 VSS.n2809 0.5005
R2429 VSS.n3194 VSS.n2803 0.5005
R2430 VSS.n3193 VSS.n2802 0.5005
R2431 VSS.n3192 VSS.n3191 0.5005
R2432 VSS.n3179 VSS.n2814 0.5005
R2433 VSS.n3158 VSS.n2821 0.5005
R2434 VSS.n3159 VSS.n2826 0.5005
R2435 VSS.n3161 VSS.n3160 0.5005
R2436 VSS.n2834 VSS.n2830 0.5005
R2437 VSS.n3151 VSS.n3150 0.5005
R2438 VSS.n3139 VSS.n2836 0.5005
R2439 VSS.n3113 VSS.n2842 0.5005
R2440 VSS.n3114 VSS.n2847 0.5005
R2441 VSS.n3116 VSS.n3115 0.5005
R2442 VSS.n2854 VSS.n2851 0.5005
R2443 VSS.n3107 VSS.n3106 0.5005
R2444 VSS.n2865 VSS.n2856 0.5005
R2445 VSS.n3093 VSS.n3092 0.5005
R2446 VSS.n2867 VSS.n2863 0.5005
R2447 VSS.n3088 VSS.n3087 0.5005
R2448 VSS.n3078 VSS.n2869 0.5005
R2449 VSS.n3034 VSS.n2875 0.5005
R2450 VSS.n3035 VSS.n2880 0.5005
R2451 VSS.n3038 VSS.n3037 0.5005
R2452 VSS.n3040 VSS.n3039 0.5005
R2453 VSS.n2889 VSS.n2886 0.5005
R2454 VSS.n3027 VSS.n3026 0.5005
R2455 VSS.n3017 VSS.n2891 0.5005
R2456 VSS.n2986 VSS.n2897 0.5005
R2457 VSS.n2987 VSS.n2902 0.5005
R2458 VSS.n2989 VSS.n2988 0.5005
R2459 VSS.n2909 VSS.n2906 0.5005
R2460 VSS.n2980 VSS.n2979 0.5005
R2461 VSS.n2970 VSS.n2911 0.5005
R2462 VSS.n2942 VSS.n2917 0.5005
R2463 VSS.n2943 VSS.n2922 0.5005
R2464 VSS.n2945 VSS.n2944 0.5005
R2465 VSS.n2929 VSS.n2926 0.5005
R2466 VSS.n5161 VSS.n5160 0.5005
R2467 VSS.n5159 VSS.n5139 0.5005
R2468 VSS.n5158 VSS.n5157 0.5005
R2469 VSS.n5156 VSS.n5140 0.5005
R2470 VSS.n5155 VSS.n5154 0.5005
R2471 VSS.n5153 VSS.n5145 0.5005
R2472 VSS.n5152 VSS.n5151 0.5005
R2473 VSS VSS.n4857 0.497977
R2474 VSS VSS.n2700 0.497977
R2475 VSS VSS.n2699 0.497977
R2476 VSS VSS.n3253 0.497977
R2477 VSS.n3676 VSS.n3624 0.497868
R2478 VSS.n3567 VSS.n3566 0.497868
R2479 VSS.n4201 VSS.n4200 0.495738
R2480 VSS.n1079 VSS.n1078 0.490418
R2481 VSS.n2517 VSS.n2516 0.478861
R2482 VSS.n5265 VSS.n2227 0.477527
R2483 VSS.n5266 VSS.n5265 0.473227
R2484 VSS.n3255 VSS.n3254 0.473227
R2485 VSS.n3614 VSS.n3613 0.473227
R2486 VSS.n3613 VSS.n3612 0.473227
R2487 VSS.n4860 VSS.n4859 0.473227
R2488 VSS.n4859 VSS.n4858 0.473227
R2489 VSS.n2520 VSS.n2519 0.473227
R2490 VSS.n5437 DVSS 0.469029
R2491 VSS.n2931 DVSS 0.467804
R2492 DVSS VSS.n2931 0.467804
R2493 VSS.n2528 VSS.n2527 0.465755
R2494 VSS.n4238 VSS.n4237 0.461183
R2495 VSS.n2515 VSS.n2513 0.457714
R2496 VSS.n2766 VSS.n2762 0.455549
R2497 VSS.n3363 VSS.n3361 0.455549
R2498 VSS.n1832 VSS.n1830 0.455549
R2499 VSS.n5715 VSS.n4 0.455549
R2500 VSS.n4302 VSS.n4301 0.452884
R2501 VSS.n4852 VSS.n4851 0.452868
R2502 VSS.n4302 VSS.n4218 0.452744
R2503 VSS.n3362 VSS.n3359 0.4505
R2504 VSS.n3368 VSS.n3360 0.4505
R2505 VSS.n3374 VSS.n3358 0.4505
R2506 VSS.n3376 VSS.n3375 0.4505
R2507 VSS.n3377 VSS.n3357 0.4505
R2508 VSS.n3379 VSS.n3378 0.4505
R2509 VSS.n3356 VSS.n3355 0.4505
R2510 VSS.n3384 VSS.n3383 0.4505
R2511 VSS.n3385 VSS.n3354 0.4505
R2512 VSS.n3387 VSS.n3386 0.4505
R2513 VSS.n3352 VSS.n3351 0.4505
R2514 VSS.n3392 VSS.n3391 0.4505
R2515 VSS.n3393 VSS.n3350 0.4505
R2516 VSS.n3395 VSS.n3394 0.4505
R2517 VSS.n3348 VSS.n3347 0.4505
R2518 VSS.n3400 VSS.n3399 0.4505
R2519 VSS.n3401 VSS.n3346 0.4505
R2520 VSS.n3403 VSS.n3402 0.4505
R2521 VSS.n3344 VSS.n3343 0.4505
R2522 VSS.n3408 VSS.n3407 0.4505
R2523 VSS.n3409 VSS.n3342 0.4505
R2524 VSS.n3411 VSS.n3410 0.4505
R2525 VSS.n3340 VSS.n3339 0.4505
R2526 VSS.n3416 VSS.n3415 0.4505
R2527 VSS.n3417 VSS.n3338 0.4505
R2528 VSS.n3419 VSS.n3418 0.4505
R2529 VSS.n3336 VSS.n3335 0.4505
R2530 VSS.n3424 VSS.n3423 0.4505
R2531 VSS.n3425 VSS.n3334 0.4505
R2532 VSS.n3427 VSS.n3426 0.4505
R2533 VSS.n3332 VSS.n3331 0.4505
R2534 VSS.n3432 VSS.n3431 0.4505
R2535 VSS.n3433 VSS.n3330 0.4505
R2536 VSS.n3435 VSS.n3434 0.4505
R2537 VSS.n3328 VSS.n3327 0.4505
R2538 VSS.n3440 VSS.n3439 0.4505
R2539 VSS.n3441 VSS.n3326 0.4505
R2540 VSS.n3443 VSS.n3442 0.4505
R2541 VSS.n3324 VSS.n3323 0.4505
R2542 VSS.n3448 VSS.n3447 0.4505
R2543 VSS.n3449 VSS.n3322 0.4505
R2544 VSS.n3451 VSS.n3450 0.4505
R2545 VSS.n3320 VSS.n3319 0.4505
R2546 VSS.n3456 VSS.n3455 0.4505
R2547 VSS.n3457 VSS.n3318 0.4505
R2548 VSS.n3459 VSS.n3458 0.4505
R2549 VSS.n3316 VSS.n3315 0.4505
R2550 VSS.n3464 VSS.n3463 0.4505
R2551 VSS.n3465 VSS.n3314 0.4505
R2552 VSS.n3467 VSS.n3466 0.4505
R2553 VSS.n3312 VSS.n3311 0.4505
R2554 VSS.n3472 VSS.n3471 0.4505
R2555 VSS.n3473 VSS.n3310 0.4505
R2556 VSS.n3475 VSS.n3474 0.4505
R2557 VSS.n3308 VSS.n3307 0.4505
R2558 VSS.n3480 VSS.n3479 0.4505
R2559 VSS.n3481 VSS.n3306 0.4505
R2560 VSS.n3483 VSS.n3482 0.4505
R2561 VSS.n3304 VSS.n3303 0.4505
R2562 VSS.n3488 VSS.n3487 0.4505
R2563 VSS.n3489 VSS.n3302 0.4505
R2564 VSS.n3491 VSS.n3490 0.4505
R2565 VSS.n3300 VSS.n3299 0.4505
R2566 VSS.n3496 VSS.n3495 0.4505
R2567 VSS.n3497 VSS.n3298 0.4505
R2568 VSS.n3499 VSS.n3498 0.4505
R2569 VSS.n3296 VSS.n3295 0.4505
R2570 VSS.n3504 VSS.n3503 0.4505
R2571 VSS.n3505 VSS.n3294 0.4505
R2572 VSS.n3507 VSS.n3506 0.4505
R2573 VSS.n3292 VSS.n3291 0.4505
R2574 VSS.n3512 VSS.n3511 0.4505
R2575 VSS.n3513 VSS.n2737 0.4505
R2576 VSS.n2770 VSS.n2769 0.4505
R2577 VSS.n2771 VSS.n2761 0.4505
R2578 VSS.n2773 VSS.n2772 0.4505
R2579 VSS.n2759 VSS.n2758 0.4505
R2580 VSS.n2778 VSS.n2777 0.4505
R2581 VSS.n2779 VSS.n2757 0.4505
R2582 VSS.n2781 VSS.n2780 0.4505
R2583 VSS.n2755 VSS.n2754 0.4505
R2584 VSS.n2786 VSS.n2785 0.4505
R2585 VSS.n2787 VSS.n2753 0.4505
R2586 VSS.n2789 VSS.n2788 0.4505
R2587 VSS.n2751 VSS.n2750 0.4505
R2588 VSS.n3265 VSS.n3264 0.4505
R2589 VSS.n3266 VSS.n2749 0.4505
R2590 VSS.n3268 VSS.n3267 0.4505
R2591 VSS.n2747 VSS.n2746 0.4505
R2592 VSS.n3273 VSS.n3272 0.4505
R2593 VSS.n3274 VSS.n2745 0.4505
R2594 VSS.n3276 VSS.n3275 0.4505
R2595 VSS.n2743 VSS.n2742 0.4505
R2596 VSS.n3281 VSS.n3280 0.4505
R2597 VSS.n3282 VSS.n2741 0.4505
R2598 VSS.n3284 VSS.n3283 0.4505
R2599 VSS.n2739 VSS.n2738 0.4505
R2600 VSS.n3289 VSS.n3288 0.4505
R2601 VSS.n3290 VSS.n2736 0.4505
R2602 VSS.n3515 VSS.n3514 0.4505
R2603 VSS.n3529 VSS.n3526 0.4505
R2604 VSS.n2647 VSS.n2646 0.4505
R2605 VSS.n3800 VSS.n3799 0.4505
R2606 VSS.n3802 VSS.n3801 0.4505
R2607 VSS.n3793 VSS.n3792 0.4505
R2608 VSS.n3809 VSS.n3808 0.4505
R2609 VSS.n3810 VSS.n3791 0.4505
R2610 VSS.n3812 VSS.n3811 0.4505
R2611 VSS.n3738 VSS.n3736 0.4505
R2612 VSS.n4159 VSS.n4158 0.4505
R2613 VSS.n4157 VSS.n3737 0.4505
R2614 VSS.n4156 VSS.n4155 0.4505
R2615 VSS.n3740 VSS.n3739 0.4505
R2616 VSS.n3874 VSS.n3873 0.4505
R2617 VSS.n3765 VSS.n3763 0.4505
R2618 VSS.n4141 VSS.n4140 0.4505
R2619 VSS.n4139 VSS.n3764 0.4505
R2620 VSS.n4138 VSS.n4137 0.4505
R2621 VSS.n3767 VSS.n3766 0.4505
R2622 VSS.n3917 VSS.n3916 0.4505
R2623 VSS.n3934 VSS.n3933 0.4505
R2624 VSS.n3935 VSS.n3913 0.4505
R2625 VSS.n3938 VSS.n3937 0.4505
R2626 VSS.n3936 VSS.n3915 0.4505
R2627 VSS.n3896 VSS.n3894 0.4505
R2628 VSS.n4112 VSS.n4111 0.4505
R2629 VSS.n4110 VSS.n3895 0.4505
R2630 VSS.n4109 VSS.n4108 0.4505
R2631 VSS.n3898 VSS.n3897 0.4505
R2632 VSS.n3961 VSS.n3959 0.4505
R2633 VSS.n4096 VSS.n4095 0.4505
R2634 VSS.n4094 VSS.n3960 0.4505
R2635 VSS.n4093 VSS.n4092 0.4505
R2636 VSS.n3963 VSS.n3962 0.4505
R2637 VSS.n4054 VSS.n4053 0.4505
R2638 VSS.n4052 VSS.n3967 0.4505
R2639 VSS.n4051 VSS.n4050 0.4505
R2640 VSS.n3969 VSS.n3968 0.4505
R2641 VSS.n4046 VSS.n4045 0.4505
R2642 VSS.n4044 VSS.n3971 0.4505
R2643 VSS.n4043 VSS.n4042 0.4505
R2644 VSS.n3973 VSS.n3972 0.4505
R2645 VSS.n4038 VSS.n4037 0.4505
R2646 VSS.n4036 VSS.n3975 0.4505
R2647 VSS.n4035 VSS.n4034 0.4505
R2648 VSS.n3977 VSS.n3976 0.4505
R2649 VSS.n4030 VSS.n4029 0.4505
R2650 VSS.n4028 VSS.n3979 0.4505
R2651 VSS.n4027 VSS.n4026 0.4505
R2652 VSS.n3981 VSS.n3980 0.4505
R2653 VSS.n4022 VSS.n4021 0.4505
R2654 VSS.n4020 VSS.n3983 0.4505
R2655 VSS.n4019 VSS.n4018 0.4505
R2656 VSS.n3985 VSS.n3984 0.4505
R2657 VSS.n4014 VSS.n4013 0.4505
R2658 VSS.n4012 VSS.n3987 0.4505
R2659 VSS.n4011 VSS.n4010 0.4505
R2660 VSS.n3989 VSS.n3988 0.4505
R2661 VSS.n4006 VSS.n4005 0.4505
R2662 VSS.n4004 VSS.n3991 0.4505
R2663 VSS.n4003 VSS.n4002 0.4505
R2664 VSS.n3993 VSS.n3992 0.4505
R2665 VSS.n3998 VSS.n3997 0.4505
R2666 VSS.n3996 VSS.n3995 0.4505
R2667 VSS.n4188 VSS.n4187 0.4505
R2668 VSS.n4186 VSS.n2640 0.4505
R2669 VSS.n4185 VSS.n4184 0.4505
R2670 VSS.n2642 VSS.n2641 0.4505
R2671 VSS.n4180 VSS.n4179 0.4505
R2672 VSS.n4178 VSS.n2645 0.4505
R2673 VSS.n4177 VSS.n4176 0.4505
R2674 VSS.n4380 VSS.n4379 0.4505
R2675 VSS.n4384 VSS.n4383 0.4505
R2676 VSS.n4385 VSS.n4378 0.4505
R2677 VSS.n4387 VSS.n4386 0.4505
R2678 VSS.n4376 VSS.n4375 0.4505
R2679 VSS.n4392 VSS.n4391 0.4505
R2680 VSS.n4393 VSS.n4374 0.4505
R2681 VSS.n4395 VSS.n4394 0.4505
R2682 VSS.n4372 VSS.n4371 0.4505
R2683 VSS.n4400 VSS.n4399 0.4505
R2684 VSS.n4401 VSS.n4370 0.4505
R2685 VSS.n4403 VSS.n4402 0.4505
R2686 VSS.n4368 VSS.n4367 0.4505
R2687 VSS.n4408 VSS.n4407 0.4505
R2688 VSS.n4409 VSS.n4366 0.4505
R2689 VSS.n4411 VSS.n4410 0.4505
R2690 VSS.n4364 VSS.n4363 0.4505
R2691 VSS.n4416 VSS.n4415 0.4505
R2692 VSS.n4417 VSS.n4362 0.4505
R2693 VSS.n4419 VSS.n4418 0.4505
R2694 VSS.n4360 VSS.n4359 0.4505
R2695 VSS.n4424 VSS.n4423 0.4505
R2696 VSS.n4425 VSS.n4358 0.4505
R2697 VSS.n4427 VSS.n4426 0.4505
R2698 VSS.n4356 VSS.n4355 0.4505
R2699 VSS.n4432 VSS.n4431 0.4505
R2700 VSS.n4433 VSS.n4351 0.4505
R2701 VSS.n4524 VSS.n2550 0.4505
R2702 VSS.n2553 VSS.n2549 0.4505
R2703 VSS.n4520 VSS.n4519 0.4505
R2704 VSS.n4518 VSS.n2552 0.4505
R2705 VSS.n4517 VSS.n4516 0.4505
R2706 VSS.n2555 VSS.n2554 0.4505
R2707 VSS.n4510 VSS.n4509 0.4505
R2708 VSS.n4508 VSS.n2570 0.4505
R2709 VSS.n4507 VSS.n4506 0.4505
R2710 VSS.n2572 VSS.n2571 0.4505
R2711 VSS.n4502 VSS.n4501 0.4505
R2712 VSS.n4500 VSS.n2574 0.4505
R2713 VSS.n4499 VSS.n4498 0.4505
R2714 VSS.n2576 VSS.n2575 0.4505
R2715 VSS.n4494 VSS.n4493 0.4505
R2716 VSS.n4492 VSS.n2578 0.4505
R2717 VSS.n4491 VSS.n4490 0.4505
R2718 VSS.n2580 VSS.n2579 0.4505
R2719 VSS.n4486 VSS.n4485 0.4505
R2720 VSS.n4484 VSS.n2582 0.4505
R2721 VSS.n4483 VSS.n4482 0.4505
R2722 VSS.n2584 VSS.n2583 0.4505
R2723 VSS.n4478 VSS.n4477 0.4505
R2724 VSS.n4476 VSS.n2586 0.4505
R2725 VSS.n4475 VSS.n4474 0.4505
R2726 VSS.n2588 VSS.n2587 0.4505
R2727 VSS.n4470 VSS.n4469 0.4505
R2728 VSS.n4468 VSS.n2590 0.4505
R2729 VSS.n4467 VSS.n4466 0.4505
R2730 VSS.n2592 VSS.n2591 0.4505
R2731 VSS.n4462 VSS.n4461 0.4505
R2732 VSS.n4460 VSS.n2594 0.4505
R2733 VSS.n4459 VSS.n4458 0.4505
R2734 VSS.n2596 VSS.n2595 0.4505
R2735 VSS.n4454 VSS.n4453 0.4505
R2736 VSS.n4452 VSS.n2598 0.4505
R2737 VSS.n4451 VSS.n4450 0.4505
R2738 VSS.n2600 VSS.n2599 0.4505
R2739 VSS.n4446 VSS.n4445 0.4505
R2740 VSS.n4444 VSS.n2602 0.4505
R2741 VSS.n4443 VSS.n4442 0.4505
R2742 VSS.n2604 VSS.n2603 0.4505
R2743 VSS.n4353 VSS.n4352 0.4505
R2744 VSS.n4354 VSS.n4350 0.4505
R2745 VSS.n4435 VSS.n4434 0.4505
R2746 VSS.n4351 VSS.n4349 0.4505
R2747 VSS.n4526 VSS.n4525 0.4505
R2748 VSS.n4431 VSS.n4430 0.4505
R2749 VSS.n4429 VSS.n4356 0.4505
R2750 VSS.n4428 VSS.n4427 0.4505
R2751 VSS.n4358 VSS.n4357 0.4505
R2752 VSS.n4423 VSS.n4422 0.4505
R2753 VSS.n4421 VSS.n4360 0.4505
R2754 VSS.n4420 VSS.n4419 0.4505
R2755 VSS.n4362 VSS.n4361 0.4505
R2756 VSS.n4415 VSS.n4414 0.4505
R2757 VSS.n4413 VSS.n4364 0.4505
R2758 VSS.n4412 VSS.n4411 0.4505
R2759 VSS.n4366 VSS.n4365 0.4505
R2760 VSS.n4407 VSS.n4406 0.4505
R2761 VSS.n4405 VSS.n4368 0.4505
R2762 VSS.n4404 VSS.n4403 0.4505
R2763 VSS.n4370 VSS.n4369 0.4505
R2764 VSS.n4399 VSS.n4398 0.4505
R2765 VSS.n4397 VSS.n4372 0.4505
R2766 VSS.n4396 VSS.n4395 0.4505
R2767 VSS.n4374 VSS.n4373 0.4505
R2768 VSS.n4391 VSS.n4390 0.4505
R2769 VSS.n4389 VSS.n4376 0.4505
R2770 VSS.n4388 VSS.n4387 0.4505
R2771 VSS.n4378 VSS.n4377 0.4505
R2772 VSS.n4383 VSS.n4382 0.4505
R2773 VSS.n4524 VSS.n4523 0.4505
R2774 VSS.n4522 VSS.n2549 0.4505
R2775 VSS.n4521 VSS.n4520 0.4505
R2776 VSS.n2552 VSS.n2551 0.4505
R2777 VSS.n4516 VSS.n4515 0.4505
R2778 VSS.n2562 VSS.n2555 0.4505
R2779 VSS.n4511 VSS.n4510 0.4505
R2780 VSS.n2570 VSS.n2569 0.4505
R2781 VSS.n4506 VSS.n4505 0.4505
R2782 VSS.n4504 VSS.n2572 0.4505
R2783 VSS.n4503 VSS.n4502 0.4505
R2784 VSS.n2574 VSS.n2573 0.4505
R2785 VSS.n4498 VSS.n4497 0.4505
R2786 VSS.n4496 VSS.n2576 0.4505
R2787 VSS.n4495 VSS.n4494 0.4505
R2788 VSS.n2578 VSS.n2577 0.4505
R2789 VSS.n4490 VSS.n4489 0.4505
R2790 VSS.n4488 VSS.n2580 0.4505
R2791 VSS.n4487 VSS.n4486 0.4505
R2792 VSS.n2582 VSS.n2581 0.4505
R2793 VSS.n4482 VSS.n4481 0.4505
R2794 VSS.n4480 VSS.n2584 0.4505
R2795 VSS.n4479 VSS.n4478 0.4505
R2796 VSS.n2586 VSS.n2585 0.4505
R2797 VSS.n4474 VSS.n4473 0.4505
R2798 VSS.n4472 VSS.n2588 0.4505
R2799 VSS.n4471 VSS.n4470 0.4505
R2800 VSS.n2590 VSS.n2589 0.4505
R2801 VSS.n4466 VSS.n4465 0.4505
R2802 VSS.n4464 VSS.n2592 0.4505
R2803 VSS.n4463 VSS.n4462 0.4505
R2804 VSS.n2594 VSS.n2593 0.4505
R2805 VSS.n4458 VSS.n4457 0.4505
R2806 VSS.n4456 VSS.n2596 0.4505
R2807 VSS.n4455 VSS.n4454 0.4505
R2808 VSS.n2598 VSS.n2597 0.4505
R2809 VSS.n4450 VSS.n4449 0.4505
R2810 VSS.n4448 VSS.n2600 0.4505
R2811 VSS.n4447 VSS.n4446 0.4505
R2812 VSS.n2602 VSS.n2601 0.4505
R2813 VSS.n4442 VSS.n4441 0.4505
R2814 VSS.n4440 VSS.n2604 0.4505
R2815 VSS.n4352 VSS.n2609 0.4505
R2816 VSS.n4350 VSS.n4348 0.4505
R2817 VSS.n4436 VSS.n4435 0.4505
R2818 VSS.n1837 VSS.n1829 0.4505
R2819 VSS.n1831 VSS.n1828 0.4505
R2820 VSS.n2060 VSS.n2059 0.4505
R2821 VSS.n2058 VSS.n1614 0.4505
R2822 VSS.n2057 VSS.n2056 0.4505
R2823 VSS.n1616 VSS.n1615 0.4505
R2824 VSS.n2052 VSS.n2051 0.4505
R2825 VSS.n2050 VSS.n1619 0.4505
R2826 VSS.n2049 VSS.n2048 0.4505
R2827 VSS.n1621 VSS.n1620 0.4505
R2828 VSS.n1637 VSS.n1635 0.4505
R2829 VSS.n2036 VSS.n2035 0.4505
R2830 VSS.n2034 VSS.n1636 0.4505
R2831 VSS.n2033 VSS.n2032 0.4505
R2832 VSS.n1639 VSS.n1638 0.4505
R2833 VSS.n2028 VSS.n2027 0.4505
R2834 VSS.n2026 VSS.n1645 0.4505
R2835 VSS.n2025 VSS.n2024 0.4505
R2836 VSS.n1647 VSS.n1646 0.4505
R2837 VSS.n1654 VSS.n1652 0.4505
R2838 VSS.n2016 VSS.n2015 0.4505
R2839 VSS.n2014 VSS.n1653 0.4505
R2840 VSS.n2013 VSS.n2012 0.4505
R2841 VSS.n1656 VSS.n1655 0.4505
R2842 VSS.n1668 VSS.n1666 0.4505
R2843 VSS.n2003 VSS.n2002 0.4505
R2844 VSS.n2001 VSS.n1667 0.4505
R2845 VSS.n2000 VSS.n1999 0.4505
R2846 VSS.n1670 VSS.n1669 0.4505
R2847 VSS.n1995 VSS.n1994 0.4505
R2848 VSS.n1993 VSS.n1672 0.4505
R2849 VSS.n1992 VSS.n1991 0.4505
R2850 VSS.n1674 VSS.n1673 0.4505
R2851 VSS.n1984 VSS.n1983 0.4505
R2852 VSS.n1982 VSS.n1679 0.4505
R2853 VSS.n1981 VSS.n1980 0.4505
R2854 VSS.n1681 VSS.n1680 0.4505
R2855 VSS.n1693 VSS.n1691 0.4505
R2856 VSS.n1971 VSS.n1970 0.4505
R2857 VSS.n1969 VSS.n1692 0.4505
R2858 VSS.n1968 VSS.n1967 0.4505
R2859 VSS.n1695 VSS.n1694 0.4505
R2860 VSS.n1963 VSS.n1962 0.4505
R2861 VSS.n1961 VSS.n1697 0.4505
R2862 VSS.n1960 VSS.n1959 0.4505
R2863 VSS.n1699 VSS.n1698 0.4505
R2864 VSS.n1711 VSS.n1709 0.4505
R2865 VSS.n1948 VSS.n1947 0.4505
R2866 VSS.n1946 VSS.n1710 0.4505
R2867 VSS.n1945 VSS.n1944 0.4505
R2868 VSS.n1713 VSS.n1712 0.4505
R2869 VSS.n1933 VSS.n1932 0.4505
R2870 VSS.n1931 VSS.n1717 0.4505
R2871 VSS.n1930 VSS.n1929 0.4505
R2872 VSS.n1719 VSS.n1718 0.4505
R2873 VSS.n1925 VSS.n1924 0.4505
R2874 VSS.n1923 VSS.n1721 0.4505
R2875 VSS.n1922 VSS.n1921 0.4505
R2876 VSS.n1723 VSS.n1722 0.4505
R2877 VSS.n1753 VSS.n1751 0.4505
R2878 VSS.n1910 VSS.n1909 0.4505
R2879 VSS.n1908 VSS.n1752 0.4505
R2880 VSS.n1907 VSS.n1906 0.4505
R2881 VSS.n1755 VSS.n1754 0.4505
R2882 VSS.n1895 VSS.n1894 0.4505
R2883 VSS.n1893 VSS.n1759 0.4505
R2884 VSS.n1892 VSS.n1891 0.4505
R2885 VSS.n1761 VSS.n1760 0.4505
R2886 VSS.n1887 VSS.n1886 0.4505
R2887 VSS.n1885 VSS.n1763 0.4505
R2888 VSS.n1884 VSS.n1883 0.4505
R2889 VSS.n1765 VSS.n1764 0.4505
R2890 VSS.n1781 VSS.n1779 0.4505
R2891 VSS.n1871 VSS.n1870 0.4505
R2892 VSS.n1869 VSS.n1780 0.4505
R2893 VSS.n1868 VSS.n1867 0.4505
R2894 VSS.n1783 VSS.n1782 0.4505
R2895 VSS.n1863 VSS.n1862 0.4505
R2896 VSS.n1861 VSS.n1789 0.4505
R2897 VSS.n1860 VSS.n1859 0.4505
R2898 VSS.n1791 VSS.n1790 0.4505
R2899 VSS.n1852 VSS.n1851 0.4505
R2900 VSS.n1850 VSS.n1822 0.4505
R2901 VSS.n1849 VSS.n1848 0.4505
R2902 VSS.n1824 VSS.n1823 0.4505
R2903 VSS.n1844 VSS.n1843 0.4505
R2904 VSS.n1842 VSS.n1826 0.4505
R2905 VSS.n1841 VSS.n1840 0.4505
R2906 VSS.n1839 VSS.n1827 0.4505
R2907 VSS.n1834 VSS.n1833 0.4505
R2908 VSS.n1835 VSS.n1828 0.4505
R2909 VSS.n1837 VSS.n1836 0.4505
R2910 VSS.n1613 VSS.n1603 0.4505
R2911 VSS.n2061 VSS.n2060 0.4505
R2912 VSS.n1617 VSS.n1614 0.4505
R2913 VSS.n2056 VSS.n2055 0.4505
R2914 VSS.n2054 VSS.n1616 0.4505
R2915 VSS.n2053 VSS.n2052 0.4505
R2916 VSS.n1622 VSS.n1619 0.4505
R2917 VSS.n2048 VSS.n2047 0.4505
R2918 VSS.n1624 VSS.n1621 0.4505
R2919 VSS.n1635 VSS.n1633 0.4505
R2920 VSS.n2037 VSS.n2036 0.4505
R2921 VSS.n1640 VSS.n1636 0.4505
R2922 VSS.n2032 VSS.n2031 0.4505
R2923 VSS.n2030 VSS.n1639 0.4505
R2924 VSS.n2029 VSS.n2028 0.4505
R2925 VSS.n1645 VSS.n1644 0.4505
R2926 VSS.n2024 VSS.n2023 0.4505
R2927 VSS.n2022 VSS.n1647 0.4505
R2928 VSS.n1652 VSS.n1648 0.4505
R2929 VSS.n2017 VSS.n2016 0.4505
R2930 VSS.n1657 VSS.n1653 0.4505
R2931 VSS.n2012 VSS.n2011 0.4505
R2932 VSS.n1659 VSS.n1656 0.4505
R2933 VSS.n1666 VSS.n1664 0.4505
R2934 VSS.n2004 VSS.n2003 0.4505
R2935 VSS.n1667 VSS.n1665 0.4505
R2936 VSS.n1999 VSS.n1998 0.4505
R2937 VSS.n1997 VSS.n1670 0.4505
R2938 VSS.n1996 VSS.n1995 0.4505
R2939 VSS.n1672 VSS.n1671 0.4505
R2940 VSS.n1991 VSS.n1990 0.4505
R2941 VSS.n1675 VSS.n1674 0.4505
R2942 VSS.n1985 VSS.n1984 0.4505
R2943 VSS.n1682 VSS.n1679 0.4505
R2944 VSS.n1980 VSS.n1979 0.4505
R2945 VSS.n1684 VSS.n1681 0.4505
R2946 VSS.n1691 VSS.n1689 0.4505
R2947 VSS.n1972 VSS.n1971 0.4505
R2948 VSS.n1692 VSS.n1690 0.4505
R2949 VSS.n1967 VSS.n1966 0.4505
R2950 VSS.n1965 VSS.n1695 0.4505
R2951 VSS.n1964 VSS.n1963 0.4505
R2952 VSS.n1697 VSS.n1696 0.4505
R2953 VSS.n1959 VSS.n1958 0.4505
R2954 VSS.n1701 VSS.n1699 0.4505
R2955 VSS.n1709 VSS.n1707 0.4505
R2956 VSS.n1949 VSS.n1948 0.4505
R2957 VSS.n1714 VSS.n1710 0.4505
R2958 VSS.n1944 VSS.n1943 0.4505
R2959 VSS.n1935 VSS.n1713 0.4505
R2960 VSS.n1934 VSS.n1933 0.4505
R2961 VSS.n1717 VSS.n1716 0.4505
R2962 VSS.n1929 VSS.n1928 0.4505
R2963 VSS.n1927 VSS.n1719 0.4505
R2964 VSS.n1926 VSS.n1925 0.4505
R2965 VSS.n1721 VSS.n1720 0.4505
R2966 VSS.n1921 VSS.n1920 0.4505
R2967 VSS.n1725 VSS.n1723 0.4505
R2968 VSS.n1751 VSS.n1749 0.4505
R2969 VSS.n1911 VSS.n1910 0.4505
R2970 VSS.n1756 VSS.n1752 0.4505
R2971 VSS.n1906 VSS.n1905 0.4505
R2972 VSS.n1897 VSS.n1755 0.4505
R2973 VSS.n1896 VSS.n1895 0.4505
R2974 VSS.n1759 VSS.n1758 0.4505
R2975 VSS.n1891 VSS.n1890 0.4505
R2976 VSS.n1889 VSS.n1761 0.4505
R2977 VSS.n1888 VSS.n1887 0.4505
R2978 VSS.n1766 VSS.n1763 0.4505
R2979 VSS.n1883 VSS.n1882 0.4505
R2980 VSS.n1768 VSS.n1765 0.4505
R2981 VSS.n1779 VSS.n1777 0.4505
R2982 VSS.n1872 VSS.n1871 0.4505
R2983 VSS.n1784 VSS.n1780 0.4505
R2984 VSS.n1867 VSS.n1866 0.4505
R2985 VSS.n1865 VSS.n1783 0.4505
R2986 VSS.n1864 VSS.n1863 0.4505
R2987 VSS.n1789 VSS.n1788 0.4505
R2988 VSS.n1859 VSS.n1858 0.4505
R2989 VSS.n1798 VSS.n1791 0.4505
R2990 VSS.n1853 VSS.n1852 0.4505
R2991 VSS.n1822 VSS.n1821 0.4505
R2992 VSS.n1848 VSS.n1847 0.4505
R2993 VSS.n1846 VSS.n1824 0.4505
R2994 VSS.n1845 VSS.n1844 0.4505
R2995 VSS.n1826 VSS.n1825 0.4505
R2996 VSS.n1840 VSS.n23 0.4505
R2997 VSS.n1839 VSS.n1838 0.4505
R2998 VSS.n1585 VSS.n1584 0.4505
R2999 VSS.n1583 VSS.n1301 0.4505
R3000 VSS.n1582 VSS.n1581 0.4505
R3001 VSS.n1304 VSS.n1303 0.4505
R3002 VSS.n1577 VSS.n1576 0.4505
R3003 VSS.n1575 VSS.n1306 0.4505
R3004 VSS.n1574 VSS.n1573 0.4505
R3005 VSS.n1308 VSS.n1307 0.4505
R3006 VSS.n1569 VSS.n1568 0.4505
R3007 VSS.n1567 VSS.n1310 0.4505
R3008 VSS.n1566 VSS.n1565 0.4505
R3009 VSS.n1312 VSS.n1311 0.4505
R3010 VSS.n1561 VSS.n1560 0.4505
R3011 VSS.n1559 VSS.n1314 0.4505
R3012 VSS.n1558 VSS.n1557 0.4505
R3013 VSS.n1316 VSS.n1315 0.4505
R3014 VSS.n1553 VSS.n1552 0.4505
R3015 VSS.n1551 VSS.n1318 0.4505
R3016 VSS.n1550 VSS.n1549 0.4505
R3017 VSS.n1320 VSS.n1319 0.4505
R3018 VSS.n1545 VSS.n1544 0.4505
R3019 VSS.n1543 VSS.n1322 0.4505
R3020 VSS.n1542 VSS.n1541 0.4505
R3021 VSS.n1324 VSS.n1323 0.4505
R3022 VSS.n1537 VSS.n1536 0.4505
R3023 VSS.n1535 VSS.n1326 0.4505
R3024 VSS.n1534 VSS.n1533 0.4505
R3025 VSS.n1328 VSS.n1327 0.4505
R3026 VSS.n1529 VSS.n1528 0.4505
R3027 VSS.n1527 VSS.n1330 0.4505
R3028 VSS.n1526 VSS.n1525 0.4505
R3029 VSS.n1332 VSS.n1331 0.4505
R3030 VSS.n1521 VSS.n1520 0.4505
R3031 VSS.n1519 VSS.n1334 0.4505
R3032 VSS.n1518 VSS.n1517 0.4505
R3033 VSS.n1336 VSS.n1335 0.4505
R3034 VSS.n1513 VSS.n1512 0.4505
R3035 VSS.n1511 VSS.n1338 0.4505
R3036 VSS.n1510 VSS.n1509 0.4505
R3037 VSS.n1340 VSS.n1339 0.4505
R3038 VSS.n1505 VSS.n1504 0.4505
R3039 VSS.n1503 VSS.n1342 0.4505
R3040 VSS.n1502 VSS.n1501 0.4505
R3041 VSS.n1344 VSS.n1343 0.4505
R3042 VSS.n1497 VSS.n1496 0.4505
R3043 VSS.n1495 VSS.n1346 0.4505
R3044 VSS.n1494 VSS.n1493 0.4505
R3045 VSS.n1348 VSS.n1347 0.4505
R3046 VSS.n1489 VSS.n1488 0.4505
R3047 VSS.n1487 VSS.n1350 0.4505
R3048 VSS.n1486 VSS.n1485 0.4505
R3049 VSS.n1352 VSS.n1351 0.4505
R3050 VSS.n1481 VSS.n1480 0.4505
R3051 VSS.n1479 VSS.n1354 0.4505
R3052 VSS.n1478 VSS.n1477 0.4505
R3053 VSS.n1356 VSS.n1355 0.4505
R3054 VSS.n1473 VSS.n1472 0.4505
R3055 VSS.n1471 VSS.n1358 0.4505
R3056 VSS.n1470 VSS.n1469 0.4505
R3057 VSS.n1360 VSS.n1359 0.4505
R3058 VSS.n1465 VSS.n1464 0.4505
R3059 VSS.n1463 VSS.n1362 0.4505
R3060 VSS.n1462 VSS.n1461 0.4505
R3061 VSS.n1364 VSS.n1363 0.4505
R3062 VSS.n1457 VSS.n1456 0.4505
R3063 VSS.n1455 VSS.n1366 0.4505
R3064 VSS.n1454 VSS.n1453 0.4505
R3065 VSS.n1368 VSS.n1367 0.4505
R3066 VSS.n1449 VSS.n1448 0.4505
R3067 VSS.n1447 VSS.n1370 0.4505
R3068 VSS.n1446 VSS.n1445 0.4505
R3069 VSS.n1372 VSS.n1371 0.4505
R3070 VSS.n1441 VSS.n1440 0.4505
R3071 VSS.n1439 VSS.n1374 0.4505
R3072 VSS.n1438 VSS.n1437 0.4505
R3073 VSS.n1376 VSS.n1375 0.4505
R3074 VSS.n1433 VSS.n1432 0.4505
R3075 VSS.n1431 VSS.n1378 0.4505
R3076 VSS.n1430 VSS.n1429 0.4505
R3077 VSS.n1380 VSS.n1379 0.4505
R3078 VSS.n1425 VSS.n1424 0.4505
R3079 VSS.n1423 VSS.n1382 0.4505
R3080 VSS.n1422 VSS.n1421 0.4505
R3081 VSS.n1384 VSS.n1383 0.4505
R3082 VSS.n1417 VSS.n1416 0.4505
R3083 VSS.n1415 VSS.n1386 0.4505
R3084 VSS.n1414 VSS.n1413 0.4505
R3085 VSS.n1388 VSS.n1387 0.4505
R3086 VSS.n1409 VSS.n1408 0.4505
R3087 VSS.n1407 VSS.n1390 0.4505
R3088 VSS.n1406 VSS.n1405 0.4505
R3089 VSS.n1392 VSS.n1391 0.4505
R3090 VSS.n1401 VSS.n1400 0.4505
R3091 VSS.n1399 VSS.n1394 0.4505
R3092 VSS.n1398 VSS.n1397 0.4505
R3093 VSS.n1300 VSS.n1298 0.4505
R3094 VSS.n1586 VSS.n1585 0.4505
R3095 VSS.n1301 VSS.n1299 0.4505
R3096 VSS.n1581 VSS.n1580 0.4505
R3097 VSS.n1579 VSS.n1304 0.4505
R3098 VSS.n1578 VSS.n1577 0.4505
R3099 VSS.n1306 VSS.n1305 0.4505
R3100 VSS.n1573 VSS.n1572 0.4505
R3101 VSS.n1571 VSS.n1308 0.4505
R3102 VSS.n1570 VSS.n1569 0.4505
R3103 VSS.n1310 VSS.n1309 0.4505
R3104 VSS.n1565 VSS.n1564 0.4505
R3105 VSS.n1563 VSS.n1312 0.4505
R3106 VSS.n1562 VSS.n1561 0.4505
R3107 VSS.n1314 VSS.n1313 0.4505
R3108 VSS.n1557 VSS.n1556 0.4505
R3109 VSS.n1555 VSS.n1316 0.4505
R3110 VSS.n1554 VSS.n1553 0.4505
R3111 VSS.n1318 VSS.n1317 0.4505
R3112 VSS.n1549 VSS.n1548 0.4505
R3113 VSS.n1547 VSS.n1320 0.4505
R3114 VSS.n1546 VSS.n1545 0.4505
R3115 VSS.n1322 VSS.n1321 0.4505
R3116 VSS.n1541 VSS.n1540 0.4505
R3117 VSS.n1539 VSS.n1324 0.4505
R3118 VSS.n1538 VSS.n1537 0.4505
R3119 VSS.n1326 VSS.n1325 0.4505
R3120 VSS.n1533 VSS.n1532 0.4505
R3121 VSS.n1531 VSS.n1328 0.4505
R3122 VSS.n1530 VSS.n1529 0.4505
R3123 VSS.n1330 VSS.n1329 0.4505
R3124 VSS.n1525 VSS.n1524 0.4505
R3125 VSS.n1523 VSS.n1332 0.4505
R3126 VSS.n1522 VSS.n1521 0.4505
R3127 VSS.n1334 VSS.n1333 0.4505
R3128 VSS.n1517 VSS.n1516 0.4505
R3129 VSS.n1515 VSS.n1336 0.4505
R3130 VSS.n1514 VSS.n1513 0.4505
R3131 VSS.n1338 VSS.n1337 0.4505
R3132 VSS.n1509 VSS.n1508 0.4505
R3133 VSS.n1507 VSS.n1340 0.4505
R3134 VSS.n1506 VSS.n1505 0.4505
R3135 VSS.n1342 VSS.n1341 0.4505
R3136 VSS.n1501 VSS.n1500 0.4505
R3137 VSS.n1499 VSS.n1344 0.4505
R3138 VSS.n1498 VSS.n1497 0.4505
R3139 VSS.n1346 VSS.n1345 0.4505
R3140 VSS.n1493 VSS.n1492 0.4505
R3141 VSS.n1491 VSS.n1348 0.4505
R3142 VSS.n1490 VSS.n1489 0.4505
R3143 VSS.n1350 VSS.n1349 0.4505
R3144 VSS.n1485 VSS.n1484 0.4505
R3145 VSS.n1483 VSS.n1352 0.4505
R3146 VSS.n1482 VSS.n1481 0.4505
R3147 VSS.n1354 VSS.n1353 0.4505
R3148 VSS.n1477 VSS.n1476 0.4505
R3149 VSS.n1475 VSS.n1356 0.4505
R3150 VSS.n1474 VSS.n1473 0.4505
R3151 VSS.n1358 VSS.n1357 0.4505
R3152 VSS.n1469 VSS.n1468 0.4505
R3153 VSS.n1467 VSS.n1360 0.4505
R3154 VSS.n1466 VSS.n1465 0.4505
R3155 VSS.n1362 VSS.n1361 0.4505
R3156 VSS.n1461 VSS.n1460 0.4505
R3157 VSS.n1459 VSS.n1364 0.4505
R3158 VSS.n1458 VSS.n1457 0.4505
R3159 VSS.n1366 VSS.n1365 0.4505
R3160 VSS.n1453 VSS.n1452 0.4505
R3161 VSS.n1451 VSS.n1368 0.4505
R3162 VSS.n1450 VSS.n1449 0.4505
R3163 VSS.n1370 VSS.n1369 0.4505
R3164 VSS.n1445 VSS.n1444 0.4505
R3165 VSS.n1443 VSS.n1372 0.4505
R3166 VSS.n1442 VSS.n1441 0.4505
R3167 VSS.n1374 VSS.n1373 0.4505
R3168 VSS.n1437 VSS.n1436 0.4505
R3169 VSS.n1435 VSS.n1376 0.4505
R3170 VSS.n1434 VSS.n1433 0.4505
R3171 VSS.n1378 VSS.n1377 0.4505
R3172 VSS.n1429 VSS.n1428 0.4505
R3173 VSS.n1427 VSS.n1380 0.4505
R3174 VSS.n1426 VSS.n1425 0.4505
R3175 VSS.n1382 VSS.n1381 0.4505
R3176 VSS.n1421 VSS.n1420 0.4505
R3177 VSS.n1419 VSS.n1384 0.4505
R3178 VSS.n1418 VSS.n1417 0.4505
R3179 VSS.n1386 VSS.n1385 0.4505
R3180 VSS.n1413 VSS.n1412 0.4505
R3181 VSS.n1411 VSS.n1388 0.4505
R3182 VSS.n1410 VSS.n1409 0.4505
R3183 VSS.n1390 VSS.n1389 0.4505
R3184 VSS.n1405 VSS.n1404 0.4505
R3185 VSS.n1403 VSS.n1392 0.4505
R3186 VSS.n1402 VSS.n1401 0.4505
R3187 VSS.n1394 VSS.n1393 0.4505
R3188 VSS.n1397 VSS.n1396 0.4505
R3189 VSS.n3999 VSS.n3998 0.4505
R3190 VSS.n4000 VSS.n3993 0.4505
R3191 VSS.n4002 VSS.n4001 0.4505
R3192 VSS.n3991 VSS.n3990 0.4505
R3193 VSS.n4007 VSS.n4006 0.4505
R3194 VSS.n4008 VSS.n3989 0.4505
R3195 VSS.n4010 VSS.n4009 0.4505
R3196 VSS.n3987 VSS.n3986 0.4505
R3197 VSS.n4015 VSS.n4014 0.4505
R3198 VSS.n4016 VSS.n3985 0.4505
R3199 VSS.n4018 VSS.n4017 0.4505
R3200 VSS.n3983 VSS.n3982 0.4505
R3201 VSS.n4023 VSS.n4022 0.4505
R3202 VSS.n4024 VSS.n3981 0.4505
R3203 VSS.n4026 VSS.n4025 0.4505
R3204 VSS.n3979 VSS.n3978 0.4505
R3205 VSS.n4031 VSS.n4030 0.4505
R3206 VSS.n4032 VSS.n3977 0.4505
R3207 VSS.n4034 VSS.n4033 0.4505
R3208 VSS.n3975 VSS.n3974 0.4505
R3209 VSS.n4039 VSS.n4038 0.4505
R3210 VSS.n4040 VSS.n3973 0.4505
R3211 VSS.n4042 VSS.n4041 0.4505
R3212 VSS.n3971 VSS.n3970 0.4505
R3213 VSS.n4047 VSS.n4046 0.4505
R3214 VSS.n4048 VSS.n3969 0.4505
R3215 VSS.n4050 VSS.n4049 0.4505
R3216 VSS.n3967 VSS.n3966 0.4505
R3217 VSS.n4055 VSS.n4054 0.4505
R3218 VSS.n4056 VSS.n3963 0.4505
R3219 VSS.n4092 VSS.n4091 0.4505
R3220 VSS.n4087 VSS.n3960 0.4505
R3221 VSS.n4097 VSS.n4096 0.4505
R3222 VSS.n3959 VSS.n3957 0.4505
R3223 VSS.n3901 VSS.n3898 0.4505
R3224 VSS.n4108 VSS.n4107 0.4505
R3225 VSS.n3899 VSS.n3895 0.4505
R3226 VSS.n4113 VSS.n4112 0.4505
R3227 VSS.n3894 VSS.n3891 0.4505
R3228 VSS.n3915 VSS.n3914 0.4505
R3229 VSS.n3939 VSS.n3938 0.4505
R3230 VSS.n3913 VSS.n3911 0.4505
R3231 VSS.n3933 VSS.n3932 0.4505
R3232 VSS.n3923 VSS.n3917 0.4505
R3233 VSS.n3770 VSS.n3767 0.4505
R3234 VSS.n4137 VSS.n4136 0.4505
R3235 VSS.n3764 VSS.n3762 0.4505
R3236 VSS.n4142 VSS.n4141 0.4505
R3237 VSS.n3763 VSS.n3761 0.4505
R3238 VSS.n3875 VSS.n3874 0.4505
R3239 VSS.n3743 VSS.n3740 0.4505
R3240 VSS.n4155 VSS.n4154 0.4505
R3241 VSS.n3741 VSS.n3737 0.4505
R3242 VSS.n4160 VSS.n4159 0.4505
R3243 VSS.n3736 VSS.n3734 0.4505
R3244 VSS.n3813 VSS.n3812 0.4505
R3245 VSS.n3791 VSS.n3790 0.4505
R3246 VSS.n2649 VSS.n2647 0.4505
R3247 VSS.n3799 VSS.n3798 0.4505
R3248 VSS.n3803 VSS.n3802 0.4505
R3249 VSS.n3794 VSS.n3793 0.4505
R3250 VSS.n3808 VSS.n3807 0.4505
R3251 VSS.n4190 VSS.n4189 0.4505
R3252 VSS.n4188 VSS.n2639 0.4505
R3253 VSS.n2643 VSS.n2640 0.4505
R3254 VSS.n4184 VSS.n4183 0.4505
R3255 VSS.n4182 VSS.n2642 0.4505
R3256 VSS.n4181 VSS.n4180 0.4505
R3257 VSS.n3826 VSS.n2645 0.4505
R3258 VSS.n4176 VSS.n4175 0.4505
R3259 VSS.n3708 VSS.n2677 0.4505
R3260 VSS.n5190 VSS.n5189 0.4505
R3261 VSS.n5192 VSS.n5191 0.4505
R3262 VSS.n5187 VSS.n5186 0.4505
R3263 VSS.n5197 VSS.n5196 0.4505
R3264 VSS.n5198 VSS.n5185 0.4505
R3265 VSS.n5200 VSS.n5199 0.4505
R3266 VSS.n2270 VSS.n2269 0.4505
R3267 VSS.n5205 VSS.n5204 0.4505
R3268 VSS.n5206 VSS.n2268 0.4505
R3269 VSS.n5208 VSS.n5207 0.4505
R3270 VSS.n2266 VSS.n2265 0.4505
R3271 VSS.n5213 VSS.n5212 0.4505
R3272 VSS.n5214 VSS.n2264 0.4505
R3273 VSS.n5216 VSS.n5215 0.4505
R3274 VSS.n2262 VSS.n2261 0.4505
R3275 VSS.n5221 VSS.n5220 0.4505
R3276 VSS.n5222 VSS.n2260 0.4505
R3277 VSS.n5224 VSS.n5223 0.4505
R3278 VSS.n2258 VSS.n2257 0.4505
R3279 VSS.n5229 VSS.n5228 0.4505
R3280 VSS.n5230 VSS.n2256 0.4505
R3281 VSS.n5232 VSS.n5231 0.4505
R3282 VSS.n2254 VSS.n2253 0.4505
R3283 VSS.n5237 VSS.n5236 0.4505
R3284 VSS.n5238 VSS.n2252 0.4505
R3285 VSS.n5240 VSS.n5239 0.4505
R3286 VSS.n2249 VSS.n2248 0.4505
R3287 VSS.n5245 VSS.n5244 0.4505
R3288 VSS.n5246 VSS.n2246 0.4505
R3289 VSS.n5248 VSS.n5247 0.4505
R3290 VSS.n2247 VSS.n2245 0.4505
R3291 VSS.n3660 VSS.n3659 0.4505
R3292 VSS.n3662 VSS.n3661 0.4505
R3293 VSS.n3657 VSS.n3656 0.4505
R3294 VSS.n3668 VSS.n3667 0.4505
R3295 VSS.n3669 VSS.n3628 0.4505
R3296 VSS.n3671 VSS.n3670 0.4505
R3297 VSS.n3655 VSS.n3627 0.4505
R3298 VSS.n3654 VSS.n3653 0.4505
R3299 VSS.n3630 VSS.n3629 0.4505
R3300 VSS.n3647 VSS.n3646 0.4505
R3301 VSS.n3645 VSS.n3632 0.4505
R3302 VSS.n3644 VSS.n3643 0.4505
R3303 VSS.n3634 VSS.n3633 0.4505
R3304 VSS.n3636 VSS.n3635 0.4505
R3305 VSS.n2691 VSS.n2690 0.4505
R3306 VSS.n3685 VSS.n3684 0.4505
R3307 VSS.n3686 VSS.n2689 0.4505
R3308 VSS.n3688 VSS.n3687 0.4505
R3309 VSS.n2687 VSS.n2686 0.4505
R3310 VSS.n3693 VSS.n3692 0.4505
R3311 VSS.n3694 VSS.n2685 0.4505
R3312 VSS.n3696 VSS.n3695 0.4505
R3313 VSS.n2683 VSS.n2682 0.4505
R3314 VSS.n3701 VSS.n3700 0.4505
R3315 VSS.n3702 VSS.n2680 0.4505
R3316 VSS.n3704 VSS.n3703 0.4505
R3317 VSS.n2681 VSS.n2678 0.4505
R3318 VSS.n3542 VSS.n3536 0.4505
R3319 VSS.n3559 VSS.n3558 0.4505
R3320 VSS.n3557 VSS.n3537 0.4505
R3321 VSS.n3556 VSS.n3555 0.4505
R3322 VSS.n3544 VSS.n3543 0.4505
R3323 VSS.n3550 VSS.n3549 0.4505
R3324 VSS.n3548 VSS.n3547 0.4505
R3325 VSS.n2722 VSS.n2721 0.4505
R3326 VSS.n3571 VSS.n3570 0.4505
R3327 VSS.n3572 VSS.n2720 0.4505
R3328 VSS.n3574 VSS.n3573 0.4505
R3329 VSS.n2718 VSS.n2717 0.4505
R3330 VSS.n3580 VSS.n3579 0.4505
R3331 VSS.n3581 VSS.n2716 0.4505
R3332 VSS.n3583 VSS.n3582 0.4505
R3333 VSS.n2714 VSS.n2713 0.4505
R3334 VSS.n3590 VSS.n3589 0.4505
R3335 VSS.n3591 VSS.n2711 0.4505
R3336 VSS.n3597 VSS.n3596 0.4505
R3337 VSS.n3595 VSS.n2712 0.4505
R3338 VSS.n3594 VSS.n3593 0.4505
R3339 VSS.n2676 VSS.n2674 0.4505
R3340 VSS.n3713 VSS.n3712 0.4505
R3341 VSS.n3711 VSS.n2675 0.4505
R3342 VSS.n3710 VSS.n3709 0.4505
R3343 VSS.n3653 VSS.n3652 0.4505
R3344 VSS.n2693 VSS.n2691 0.4505
R3345 VSS.n3637 VSS.n3636 0.4505
R3346 VSS.n3638 VSS.n3634 0.4505
R3347 VSS.n3643 VSS.n3642 0.4505
R3348 VSS.n3632 VSS.n3631 0.4505
R3349 VSS.n3648 VSS.n3647 0.4505
R3350 VSS.n3649 VSS.n3630 0.4505
R3351 VSS.n3627 VSS.n3625 0.4505
R3352 VSS.n3672 VSS.n3671 0.4505
R3353 VSS.n3628 VSS.n3626 0.4505
R3354 VSS.n3667 VSS.n3666 0.4505
R3355 VSS.n3665 VSS.n3657 0.4505
R3356 VSS.n3663 VSS.n3662 0.4505
R3357 VSS.n3659 VSS.n3658 0.4505
R3358 VSS.n2245 VSS.n2243 0.4505
R3359 VSS.n5249 VSS.n5248 0.4505
R3360 VSS.n2250 VSS.n2246 0.4505
R3361 VSS.n5244 VSS.n5243 0.4505
R3362 VSS.n5242 VSS.n2249 0.4505
R3363 VSS.n5241 VSS.n5240 0.4505
R3364 VSS.n2252 VSS.n2251 0.4505
R3365 VSS.n5236 VSS.n5235 0.4505
R3366 VSS.n5234 VSS.n2254 0.4505
R3367 VSS.n5233 VSS.n5232 0.4505
R3368 VSS.n2256 VSS.n2255 0.4505
R3369 VSS.n5228 VSS.n5227 0.4505
R3370 VSS.n5226 VSS.n2258 0.4505
R3371 VSS.n5225 VSS.n5224 0.4505
R3372 VSS.n2260 VSS.n2259 0.4505
R3373 VSS.n5220 VSS.n5219 0.4505
R3374 VSS.n5218 VSS.n2262 0.4505
R3375 VSS.n5217 VSS.n5216 0.4505
R3376 VSS.n2264 VSS.n2263 0.4505
R3377 VSS.n5212 VSS.n5211 0.4505
R3378 VSS.n5210 VSS.n2266 0.4505
R3379 VSS.n5209 VSS.n5208 0.4505
R3380 VSS.n2268 VSS.n2267 0.4505
R3381 VSS.n5204 VSS.n5203 0.4505
R3382 VSS.n5202 VSS.n2270 0.4505
R3383 VSS.n5201 VSS.n5200 0.4505
R3384 VSS.n5185 VSS.n5184 0.4505
R3385 VSS.n5196 VSS.n5195 0.4505
R3386 VSS.n5194 VSS.n5187 0.4505
R3387 VSS.n5193 VSS.n5192 0.4505
R3388 VSS.n3684 VSS.n3683 0.4505
R3389 VSS.n3708 VSS.n3707 0.4505
R3390 VSS.n3706 VSS.n2678 0.4505
R3391 VSS.n3705 VSS.n3704 0.4505
R3392 VSS.n2680 VSS.n2679 0.4505
R3393 VSS.n3700 VSS.n3699 0.4505
R3394 VSS.n3698 VSS.n2683 0.4505
R3395 VSS.n3697 VSS.n3696 0.4505
R3396 VSS.n2685 VSS.n2684 0.4505
R3397 VSS.n3692 VSS.n3691 0.4505
R3398 VSS.n3690 VSS.n2687 0.4505
R3399 VSS.n3689 VSS.n3688 0.4505
R3400 VSS.n2692 VSS.n2689 0.4505
R3401 VSS.n3540 VSS.n3539 0.4505
R3402 VSS.n3536 VSS.n3534 0.4505
R3403 VSS.n3560 VSS.n3559 0.4505
R3404 VSS.n3537 VSS.n3535 0.4505
R3405 VSS.n3555 VSS.n3554 0.4505
R3406 VSS.n3552 VSS.n3544 0.4505
R3407 VSS.n3551 VSS.n3550 0.4505
R3408 VSS.n3547 VSS.n3546 0.4505
R3409 VSS.n3545 VSS.n2722 0.4505
R3410 VSS.n3570 VSS.n3569 0.4505
R3411 VSS.n2724 VSS.n2720 0.4505
R3412 VSS.n3575 VSS.n3574 0.4505
R3413 VSS.n3576 VSS.n2718 0.4505
R3414 VSS.n3579 VSS.n3578 0.4505
R3415 VSS.n3577 VSS.n2716 0.4505
R3416 VSS.n3584 VSS.n3583 0.4505
R3417 VSS.n3585 VSS.n2714 0.4505
R3418 VSS.n3589 VSS.n3588 0.4505
R3419 VSS.n2711 VSS.n2709 0.4505
R3420 VSS.n3598 VSS.n3597 0.4505
R3421 VSS.n2712 VSS.n2710 0.4505
R3422 VSS.n3593 VSS.n3592 0.4505
R3423 VSS.n2674 VSS.n2670 0.4505
R3424 VSS.n3714 VSS.n3713 0.4505
R3425 VSS.n2675 VSS.n2656 0.4505
R3426 VSS.n3709 VSS.n2661 0.4505
R3427 VSS.n3365 VSS.n3364 0.4505
R3428 VSS.n3366 VSS.n3359 0.4505
R3429 VSS.n3368 VSS.n3367 0.4505
R3430 VSS.n3374 VSS.n3373 0.4505
R3431 VSS.n3375 VSS.n2422 0.4505
R3432 VSS.n2737 VSS.n2735 0.4505
R3433 VSS.n3511 VSS.n3510 0.4505
R3434 VSS.n3509 VSS.n3292 0.4505
R3435 VSS.n3508 VSS.n3507 0.4505
R3436 VSS.n3294 VSS.n3293 0.4505
R3437 VSS.n3503 VSS.n3502 0.4505
R3438 VSS.n3501 VSS.n3296 0.4505
R3439 VSS.n3500 VSS.n3499 0.4505
R3440 VSS.n3298 VSS.n3297 0.4505
R3441 VSS.n3495 VSS.n3494 0.4505
R3442 VSS.n3493 VSS.n3300 0.4505
R3443 VSS.n3492 VSS.n3491 0.4505
R3444 VSS.n3302 VSS.n3301 0.4505
R3445 VSS.n3487 VSS.n3486 0.4505
R3446 VSS.n3485 VSS.n3304 0.4505
R3447 VSS.n3484 VSS.n3483 0.4505
R3448 VSS.n3306 VSS.n3305 0.4505
R3449 VSS.n3479 VSS.n3478 0.4505
R3450 VSS.n3477 VSS.n3308 0.4505
R3451 VSS.n3476 VSS.n3475 0.4505
R3452 VSS.n3310 VSS.n3309 0.4505
R3453 VSS.n3471 VSS.n3470 0.4505
R3454 VSS.n3469 VSS.n3312 0.4505
R3455 VSS.n3468 VSS.n3467 0.4505
R3456 VSS.n3314 VSS.n3313 0.4505
R3457 VSS.n3463 VSS.n3462 0.4505
R3458 VSS.n3461 VSS.n3316 0.4505
R3459 VSS.n3460 VSS.n3459 0.4505
R3460 VSS.n3318 VSS.n3317 0.4505
R3461 VSS.n3455 VSS.n3454 0.4505
R3462 VSS.n3453 VSS.n3320 0.4505
R3463 VSS.n3452 VSS.n3451 0.4505
R3464 VSS.n3322 VSS.n3321 0.4505
R3465 VSS.n3447 VSS.n3446 0.4505
R3466 VSS.n3445 VSS.n3324 0.4505
R3467 VSS.n3444 VSS.n3443 0.4505
R3468 VSS.n3326 VSS.n3325 0.4505
R3469 VSS.n3439 VSS.n3438 0.4505
R3470 VSS.n3437 VSS.n3328 0.4505
R3471 VSS.n3436 VSS.n3435 0.4505
R3472 VSS.n3330 VSS.n3329 0.4505
R3473 VSS.n3431 VSS.n3430 0.4505
R3474 VSS.n3429 VSS.n3332 0.4505
R3475 VSS.n3428 VSS.n3427 0.4505
R3476 VSS.n3334 VSS.n3333 0.4505
R3477 VSS.n3423 VSS.n3422 0.4505
R3478 VSS.n3421 VSS.n3336 0.4505
R3479 VSS.n3420 VSS.n3419 0.4505
R3480 VSS.n3338 VSS.n3337 0.4505
R3481 VSS.n3415 VSS.n3414 0.4505
R3482 VSS.n3413 VSS.n3340 0.4505
R3483 VSS.n3412 VSS.n3411 0.4505
R3484 VSS.n3342 VSS.n3341 0.4505
R3485 VSS.n3407 VSS.n3406 0.4505
R3486 VSS.n3405 VSS.n3344 0.4505
R3487 VSS.n3404 VSS.n3403 0.4505
R3488 VSS.n3346 VSS.n3345 0.4505
R3489 VSS.n3399 VSS.n3398 0.4505
R3490 VSS.n3397 VSS.n3348 0.4505
R3491 VSS.n3396 VSS.n3395 0.4505
R3492 VSS.n3350 VSS.n3349 0.4505
R3493 VSS.n3391 VSS.n3390 0.4505
R3494 VSS.n3389 VSS.n3352 0.4505
R3495 VSS.n3388 VSS.n3387 0.4505
R3496 VSS.n3354 VSS.n3353 0.4505
R3497 VSS.n3383 VSS.n3382 0.4505
R3498 VSS.n3381 VSS.n3356 0.4505
R3499 VSS.n3380 VSS.n3379 0.4505
R3500 VSS.n3357 VSS.n2417 0.4505
R3501 VSS.n2767 VSS.n2763 0.4505
R3502 VSS.n2769 VSS.n2768 0.4505
R3503 VSS.n2761 VSS.n2760 0.4505
R3504 VSS.n2774 VSS.n2773 0.4505
R3505 VSS.n2775 VSS.n2759 0.4505
R3506 VSS.n2777 VSS.n2776 0.4505
R3507 VSS.n2757 VSS.n2756 0.4505
R3508 VSS.n2782 VSS.n2781 0.4505
R3509 VSS.n2783 VSS.n2755 0.4505
R3510 VSS.n2785 VSS.n2784 0.4505
R3511 VSS.n2753 VSS.n2752 0.4505
R3512 VSS.n2790 VSS.n2789 0.4505
R3513 VSS.n3262 VSS.n2751 0.4505
R3514 VSS.n3264 VSS.n3263 0.4505
R3515 VSS.n2749 VSS.n2748 0.4505
R3516 VSS.n3269 VSS.n3268 0.4505
R3517 VSS.n3270 VSS.n2747 0.4505
R3518 VSS.n3272 VSS.n3271 0.4505
R3519 VSS.n2745 VSS.n2744 0.4505
R3520 VSS.n3277 VSS.n3276 0.4505
R3521 VSS.n3278 VSS.n2743 0.4505
R3522 VSS.n3280 VSS.n3279 0.4505
R3523 VSS.n2741 VSS.n2740 0.4505
R3524 VSS.n3285 VSS.n3284 0.4505
R3525 VSS.n3286 VSS.n2739 0.4505
R3526 VSS.n3288 VSS.n3287 0.4505
R3527 VSS.n2736 VSS.n2734 0.4505
R3528 VSS.n3516 VSS.n3515 0.4505
R3529 VSS.n5716 VSS.n5 0.4505
R3530 VSS.n5718 VSS.n5717 0.4505
R3531 VSS.n6 VSS.n2 0.4505
R3532 VSS.n5723 VSS.n5722 0.4505
R3533 VSS.n4824 VSS.n4823 0.4505
R3534 VSS.n4822 VSS.n2432 0.4505
R3535 VSS.n4816 VSS.n2433 0.4505
R3536 VSS.n4818 VSS.n4817 0.4505
R3537 VSS.n4815 VSS.n2435 0.4505
R3538 VSS.n4814 VSS.n4813 0.4505
R3539 VSS.n2437 VSS.n2436 0.4505
R3540 VSS.n4809 VSS.n4808 0.4505
R3541 VSS.n4807 VSS.n2439 0.4505
R3542 VSS.n4806 VSS.n4805 0.4505
R3543 VSS.n2441 VSS.n2440 0.4505
R3544 VSS.n4801 VSS.n4800 0.4505
R3545 VSS.n4799 VSS.n2443 0.4505
R3546 VSS.n4798 VSS.n4797 0.4505
R3547 VSS.n2445 VSS.n2444 0.4505
R3548 VSS.n4793 VSS.n4792 0.4505
R3549 VSS.n4791 VSS.n2447 0.4505
R3550 VSS.n4790 VSS.n4789 0.4505
R3551 VSS.n2449 VSS.n2448 0.4505
R3552 VSS.n4785 VSS.n4784 0.4505
R3553 VSS.n4783 VSS.n2451 0.4505
R3554 VSS.n4782 VSS.n4781 0.4505
R3555 VSS.n2453 VSS.n2452 0.4505
R3556 VSS.n4777 VSS.n4776 0.4505
R3557 VSS.n4775 VSS.n2455 0.4505
R3558 VSS.n4774 VSS.n4773 0.4505
R3559 VSS.n2457 VSS.n2456 0.4505
R3560 VSS.n4769 VSS.n4768 0.4505
R3561 VSS.n4767 VSS.n2459 0.4505
R3562 VSS.n4766 VSS.n4765 0.4505
R3563 VSS.n2461 VSS.n2460 0.4505
R3564 VSS.n4761 VSS.n4760 0.4505
R3565 VSS.n4759 VSS.n2463 0.4505
R3566 VSS.n4758 VSS.n4757 0.4505
R3567 VSS.n2465 VSS.n2464 0.4505
R3568 VSS.n4753 VSS.n4752 0.4505
R3569 VSS.n4751 VSS.n2467 0.4505
R3570 VSS.n4749 VSS.n4748 0.4505
R3571 VSS.n2469 VSS.n2468 0.4505
R3572 VSS.n4744 VSS.n4743 0.4505
R3573 VSS.n4742 VSS.n2471 0.4505
R3574 VSS.n4741 VSS.n4740 0.4505
R3575 VSS.n2473 VSS.n2472 0.4505
R3576 VSS.n4736 VSS.n4735 0.4505
R3577 VSS.n4734 VSS.n2475 0.4505
R3578 VSS.n4733 VSS.n4732 0.4505
R3579 VSS.n2477 VSS.n2476 0.4505
R3580 VSS.n4728 VSS.n4727 0.4505
R3581 VSS.n4726 VSS.n2479 0.4505
R3582 VSS.n4725 VSS.n4724 0.4505
R3583 VSS.n2481 VSS.n2480 0.4505
R3584 VSS.n4720 VSS.n4719 0.4505
R3585 VSS.n4718 VSS.n2483 0.4505
R3586 VSS.n4717 VSS.n4716 0.4505
R3587 VSS.n2485 VSS.n2484 0.4505
R3588 VSS.n4712 VSS.n4711 0.4505
R3589 VSS.n4710 VSS.n2487 0.4505
R3590 VSS.n4709 VSS.n4708 0.4505
R3591 VSS.n2489 VSS.n2488 0.4505
R3592 VSS.n4704 VSS.n4703 0.4505
R3593 VSS.n4702 VSS.n2491 0.4505
R3594 VSS.n4701 VSS.n4700 0.4505
R3595 VSS.n2493 VSS.n2492 0.4505
R3596 VSS.n4696 VSS.n4695 0.4505
R3597 VSS.n4694 VSS.n2495 0.4505
R3598 VSS.n4693 VSS.n4692 0.4505
R3599 VSS.n2497 VSS.n2496 0.4505
R3600 VSS.n4688 VSS.n4687 0.4505
R3601 VSS.n2500 VSS.n2499 0.4505
R3602 VSS.n4683 VSS.n4682 0.4505
R3603 VSS.n2507 VSS.n2503 0.4505
R3604 VSS.n4678 VSS.n4677 0.4505
R3605 VSS.n4278 VSS.n2505 0.4505
R3606 VSS.n4282 VSS.n4281 0.4505
R3607 VSS.n4276 VSS.n4275 0.4505
R3608 VSS.n4287 VSS.n4286 0.4505
R3609 VSS.n4273 VSS.n4272 0.4505
R3610 VSS.n4292 VSS.n4291 0.4505
R3611 VSS.n4293 VSS.n4271 0.4505
R3612 VSS.n4295 VSS.n4294 0.4505
R3613 VSS.n4222 VSS.n4220 0.4505
R3614 VSS.n4300 VSS.n4299 0.4505
R3615 VSS.n4240 VSS.n4239 0.4505
R3616 VSS.n4241 VSS.n4236 0.4505
R3617 VSS.n4243 VSS.n4242 0.4505
R3618 VSS.n4234 VSS.n4233 0.4505
R3619 VSS.n4248 VSS.n4247 0.4505
R3620 VSS.n4249 VSS.n4232 0.4505
R3621 VSS.n4251 VSS.n4250 0.4505
R3622 VSS.n4230 VSS.n4229 0.4505
R3623 VSS.n4256 VSS.n4255 0.4505
R3624 VSS.n4257 VSS.n4228 0.4505
R3625 VSS.n4259 VSS.n4258 0.4505
R3626 VSS.n4226 VSS.n4225 0.4505
R3627 VSS.n4264 VSS.n4263 0.4505
R3628 VSS.n4265 VSS.n4224 0.4505
R3629 VSS.n4267 VSS.n4266 0.4505
R3630 VSS.n4299 VSS.n4298 0.4505
R3631 VSS.n4297 VSS.n4222 0.4505
R3632 VSS.n4296 VSS.n4295 0.4505
R3633 VSS.n4271 VSS.n4270 0.4505
R3634 VSS.n4291 VSS.n4290 0.4505
R3635 VSS.n4289 VSS.n4273 0.4505
R3636 VSS.n4288 VSS.n4287 0.4505
R3637 VSS.n4275 VSS.n4274 0.4505
R3638 VSS.n4281 VSS.n4280 0.4505
R3639 VSS.n2505 VSS.n2504 0.4505
R3640 VSS.n4679 VSS.n4678 0.4505
R3641 VSS.n4680 VSS.n2503 0.4505
R3642 VSS.n4682 VSS.n4681 0.4505
R3643 VSS.n2499 VSS.n2498 0.4505
R3644 VSS.n4689 VSS.n4688 0.4505
R3645 VSS.n4690 VSS.n2497 0.4505
R3646 VSS.n4692 VSS.n4691 0.4505
R3647 VSS.n2495 VSS.n2494 0.4505
R3648 VSS.n4697 VSS.n4696 0.4505
R3649 VSS.n4698 VSS.n2493 0.4505
R3650 VSS.n4700 VSS.n4699 0.4505
R3651 VSS.n2491 VSS.n2490 0.4505
R3652 VSS.n4705 VSS.n4704 0.4505
R3653 VSS.n4706 VSS.n2489 0.4505
R3654 VSS.n4708 VSS.n4707 0.4505
R3655 VSS.n2487 VSS.n2486 0.4505
R3656 VSS.n4713 VSS.n4712 0.4505
R3657 VSS.n4714 VSS.n2485 0.4505
R3658 VSS.n4716 VSS.n4715 0.4505
R3659 VSS.n2483 VSS.n2482 0.4505
R3660 VSS.n4721 VSS.n4720 0.4505
R3661 VSS.n4722 VSS.n2481 0.4505
R3662 VSS.n4724 VSS.n4723 0.4505
R3663 VSS.n2479 VSS.n2478 0.4505
R3664 VSS.n4729 VSS.n4728 0.4505
R3665 VSS.n4730 VSS.n2477 0.4505
R3666 VSS.n4732 VSS.n4731 0.4505
R3667 VSS.n2475 VSS.n2474 0.4505
R3668 VSS.n4737 VSS.n4736 0.4505
R3669 VSS.n4738 VSS.n2473 0.4505
R3670 VSS.n4740 VSS.n4739 0.4505
R3671 VSS.n2471 VSS.n2470 0.4505
R3672 VSS.n4745 VSS.n4744 0.4505
R3673 VSS.n4746 VSS.n2469 0.4505
R3674 VSS.n4748 VSS.n4747 0.4505
R3675 VSS.n2467 VSS.n2466 0.4505
R3676 VSS.n4754 VSS.n4753 0.4505
R3677 VSS.n4755 VSS.n2465 0.4505
R3678 VSS.n4757 VSS.n4756 0.4505
R3679 VSS.n2463 VSS.n2462 0.4505
R3680 VSS.n4762 VSS.n4761 0.4505
R3681 VSS.n4763 VSS.n2461 0.4505
R3682 VSS.n4765 VSS.n4764 0.4505
R3683 VSS.n2459 VSS.n2458 0.4505
R3684 VSS.n4770 VSS.n4769 0.4505
R3685 VSS.n4771 VSS.n2457 0.4505
R3686 VSS.n4773 VSS.n4772 0.4505
R3687 VSS.n2455 VSS.n2454 0.4505
R3688 VSS.n4778 VSS.n4777 0.4505
R3689 VSS.n4779 VSS.n2453 0.4505
R3690 VSS.n4781 VSS.n4780 0.4505
R3691 VSS.n2451 VSS.n2450 0.4505
R3692 VSS.n4786 VSS.n4785 0.4505
R3693 VSS.n4787 VSS.n2449 0.4505
R3694 VSS.n4789 VSS.n4788 0.4505
R3695 VSS.n2447 VSS.n2446 0.4505
R3696 VSS.n4794 VSS.n4793 0.4505
R3697 VSS.n4795 VSS.n2445 0.4505
R3698 VSS.n4797 VSS.n4796 0.4505
R3699 VSS.n2443 VSS.n2442 0.4505
R3700 VSS.n4802 VSS.n4801 0.4505
R3701 VSS.n4803 VSS.n2441 0.4505
R3702 VSS.n4805 VSS.n4804 0.4505
R3703 VSS.n2439 VSS.n2438 0.4505
R3704 VSS.n4810 VSS.n4809 0.4505
R3705 VSS.n4811 VSS.n2437 0.4505
R3706 VSS.n4813 VSS.n4812 0.4505
R3707 VSS.n2435 VSS.n2434 0.4505
R3708 VSS.n4819 VSS.n4818 0.4505
R3709 VSS.n4820 VSS.n2433 0.4505
R3710 VSS.n4822 VSS.n4821 0.4505
R3711 VSS.n4823 VSS.n3 0.4505
R3712 VSS.n5722 VSS.n5721 0.4505
R3713 VSS.n5720 VSS.n2 0.4505
R3714 VSS.n5719 VSS.n5718 0.4505
R3715 VSS.n4236 VSS.n4235 0.4505
R3716 VSS.n4244 VSS.n4243 0.4505
R3717 VSS.n4245 VSS.n4234 0.4505
R3718 VSS.n4247 VSS.n4246 0.4505
R3719 VSS.n4232 VSS.n4231 0.4505
R3720 VSS.n4252 VSS.n4251 0.4505
R3721 VSS.n4253 VSS.n4230 0.4505
R3722 VSS.n4255 VSS.n4254 0.4505
R3723 VSS.n4228 VSS.n4227 0.4505
R3724 VSS.n4260 VSS.n4259 0.4505
R3725 VSS.n4261 VSS.n4226 0.4505
R3726 VSS.n4263 VSS.n4262 0.4505
R3727 VSS.n4224 VSS.n4223 0.4505
R3728 VSS.n4268 VSS.n4267 0.4505
R3729 VSS.n4269 VSS.n4221 0.4505
R3730 VSS.n4221 VSS.n4219 0.4505
R3731 VSS.n5420 DVSS 0.449176
R3732 VSS.n5325 DVSS 0.449176
R3733 VSS.n5325 DVSS 0.449176
R3734 VSS.n5256 VSS.n5255 0.441235
R3735 VSS.n5695 VSS.n5694 0.439524
R3736 VSS.n1590 VSS.n1170 0.439458
R3737 VSS.n5329 VSS.n2127 0.420329
R3738 VSS.n4668 VSS.n2095 0.41962
R3739 VSS.n4209 VSS.n4208 0.4165
R3740 VSS.n4214 VSS.n4213 0.4165
R3741 VSS.n4207 VSS.n2625 0.412794
R3742 VSS.n4197 VSS.n4196 0.409053
R3743 VSS.n4202 VSS.n2632 0.409053
R3744 VSS.n4530 VSS.n4529 0.40882
R3745 VSS.n3678 DVSS 0.402853
R3746 VSS.n5261 DVSS 0.402853
R3747 VSS.n3519 DVSS 0.402853
R3748 DVSS VSS.n3564 0.402853
R3749 VSS.n4122 VSS.n4121 0.388068
R3750 VSS.n3882 VSS.n3870 0.387662
R3751 VSS.n5420 DVSS 0.384324
R3752 VSS.n4531 VSS.n4530 0.382451
R3753 VSS.n3259 VSS.n2733 0.375755
R3754 VSS.n3869 VSS.n3868 0.3755
R3755 VSS.n4120 VSS.n3783 0.3755
R3756 VSS.n4674 VSS.n4673 0.3755
R3757 VSS.n3680 VSS.n3679 0.368789
R3758 VSS.n3678 VSS.n2696 0.368789
R3759 VSS.n3677 VSS.n3623 0.368789
R3760 VSS.n3675 VSS.n3674 0.368789
R3761 VSS.n5261 VSS.n2241 0.368789
R3762 VSS.n5260 VSS.n5259 0.368789
R3763 VSS.n3586 VSS.n2708 0.368789
R3764 VSS.n3519 VSS.n3518 0.368789
R3765 VSS.n2727 VSS.n2726 0.368789
R3766 VSS.n3565 VSS.n2728 0.368789
R3767 VSS.n3564 VSS.n2729 0.368789
R3768 VSS.n3563 VSS.n3562 0.368789
R3769 VSS.n5284 VSS.n2218 0.367935
R3770 VSS.n5284 VSS.n5281 0.367935
R3771 VSS.n2233 VSS.n2205 0.367935
R3772 VSS.n2219 VSS.n2205 0.367935
R3773 VSS.n2234 VSS.n2206 0.367935
R3774 VSS.n2220 VSS.n2206 0.367935
R3775 VSS.n2235 VSS.n2207 0.367935
R3776 VSS.n2221 VSS.n2207 0.367935
R3777 VSS.n2236 VSS.n2208 0.367935
R3778 VSS.n2222 VSS.n2208 0.367935
R3779 VSS.n5270 VSS.n5269 0.367935
R3780 VSS.n2231 VSS.n2209 0.367935
R3781 VSS.n2222 VSS.n2210 0.367935
R3782 VSS.n2221 VSS.n2211 0.367935
R3783 VSS.n2220 VSS.n2212 0.367935
R3784 VSS.n2219 VSS.n2213 0.367935
R3785 VSS.n5281 VSS.n2214 0.367935
R3786 VSS.n5269 VSS.n2210 0.367935
R3787 VSS.n2236 VSS.n2211 0.367935
R3788 VSS.n2235 VSS.n2212 0.367935
R3789 VSS.n2234 VSS.n2213 0.367935
R3790 VSS.n2233 VSS.n2214 0.367935
R3791 VSS.n5287 VSS.n2218 0.367935
R3792 VSS.n5270 VSS.n2209 0.367935
R3793 VSS.n3524 VSS.n3523 0.36232
R3794 VSS.n3526 VSS.n3525 0.36232
R3795 VSS.n4331 DVSS 0.358788
R3796 VSS.n4528 VSS.n2547 0.346654
R3797 VSS.n4528 VSS.n4527 0.346654
R3798 VSS.n5322 VSS.n2134 0.342906
R3799 VSS.n5135 VSS.n2271 0.338834
R3800 VSS.n3531 VSS.n3530 0.335984
R3801 VSS.n1773 VSS.n1772 0.328381
R3802 VSS.n1786 VSS.n1774 0.328381
R3803 VSS.n1916 VSS.n1726 0.328381
R3804 VSS.n1903 VSS.n1902 0.328381
R3805 VSS.n1954 VSS.n1702 0.328381
R3806 VSS.n1941 VSS.n1940 0.328381
R3807 VSS.n1988 VSS.n1676 0.328381
R3808 VSS.n1975 VSS.n1974 0.328381
R3809 VSS.n2020 VSS.n1649 0.328381
R3810 VSS.n2007 VSS.n2006 0.328381
R3811 VSS.n1629 VSS.n1628 0.328381
R3812 VSS.n1642 VSS.n1630 0.328381
R3813 VSS.n5180 VSS.n5179 0.3255
R3814 VSS.n5179 VSS.n5178 0.3255
R3815 VSS.n5181 VSS.n2272 0.316244
R3816 VSS.n3841 VSS.n3840 0.311888
R3817 VSS.n4070 VSS.n4069 0.311888
R3818 VSS.n3529 VSS.n3528 0.309579
R3819 VSS.n2733 VSS.n2732 0.309579
R3820 VSS.n3258 VSS.n2792 0.309579
R3821 VSS.n3257 VSS.n2794 0.309579
R3822 VSS.n3530 VSS.n2733 0.307559
R3823 VSS.n5405 VSS.n5404 0.297643
R3824 VSS.n5348 VSS.n5347 0.297643
R3825 VSS.n5441 VSS.n5440 0.297643
R3826 VSS.n2530 VSS.n2100 0.297643
R3827 VSS.n1006 VSS.n1005 0.28175
R3828 VSS.n523 VSS.n375 0.28175
R3829 DVSS VSS.n2227 0.273784
R3830 VSS.n4305 VSS.n4304 0.273147
R3831 VSS.n4216 VSS.n2629 0.273147
R3832 VSS.n5336 VSS.n2127 0.271399
R3833 VSS.n5430 VSS.n2095 0.271321
R3834 VSS.n3606 VSS.n3605 0.268132
R3835 VSS.n5343 VSS.n2173 0.266421
R3836 VSS.n265 VSS.n222 0.265206
R3837 VSS.n381 VSS.n380 0.265206
R3838 VSS.n5413 VSS.n2107 0.265206
R3839 VSS.n5413 VSS.n5412 0.265206
R3840 VSS.n5389 VSS.n2127 0.264882
R3841 VSS.n4544 VSS.n2095 0.264797
R3842 VSS.n5344 VSS.n5343 0.2605
R3843 VSS.n5415 VSS.n5414 0.2605
R3844 VSS.n5447 VSS.n5446 0.2605
R3845 VSS.n2518 VSS 0.258658
R3846 VSS.n5296 VSS.n2199 0.254359
R3847 VSS.n5313 VSS.n5311 0.249324
R3848 VSS.n5309 VSS.n5308 0.249324
R3849 VSS.n4848 VSS.n4847 0.249324
R3850 VSS.n3530 VSS.n3529 0.238735
R3851 VSS.n4238 VSS.n4235 0.233167
R3852 VSS.n3868 VSS.n3867 0.231484
R3853 VSS.n4071 VSS.n3783 0.231484
R3854 VSS.n5719 VSS.n4 0.231338
R3855 VSS.n2770 VSS.n2762 0.231338
R3856 VSS.n3363 VSS.n3362 0.231338
R3857 VSS.n1832 VSS.n1831 0.231338
R3858 VSS.n3868 VSS.n3782 0.229569
R3859 VSS VSS.n5310 0.229471
R3860 VSS.n5310 VSS 0.229471
R3861 VSS.n4124 VSS.n3783 0.228851
R3862 VSS.n2518 VSS.n2517 0.224316
R3863 VSS.n1080 VSS.n1079 0.219756
R3864 VSS.n2168 VSS.n2167 0.219756
R3865 VSS.n1029 VSS.n37 0.217409
R3866 VSS.n1138 VSS.n1137 0.217409
R3867 VSS.n170 VSS.n95 0.214786
R3868 VSS.n581 VSS.n366 0.214786
R3869 VSS.n2170 VSS.n2166 0.214786
R3870 VSS.n2165 VSS.n2162 0.214786
R3871 VSS.n5355 VSS.n2161 0.214786
R3872 VSS.n5356 VSS.n2160 0.214786
R3873 VSS.n5357 VSS.n2159 0.214786
R3874 VSS.n2158 VSS.n2156 0.214786
R3875 VSS.n5361 VSS.n2155 0.214786
R3876 VSS.n5362 VSS.n2154 0.214786
R3877 VSS.n5363 VSS.n2153 0.214786
R3878 VSS.n2152 VSS.n2150 0.214786
R3879 VSS.n5367 VSS.n2149 0.214786
R3880 VSS.n5368 VSS.n2148 0.214786
R3881 VSS.n5369 VSS.n2147 0.214786
R3882 VSS.n2146 VSS.n2144 0.214786
R3883 VSS.n5373 VSS.n2143 0.214786
R3884 VSS.n5374 VSS.n2142 0.214786
R3885 VSS.n5375 VSS.n2141 0.214786
R3886 VSS.n2140 VSS.n2138 0.214786
R3887 VSS.n5379 VSS.n2137 0.214786
R3888 VSS.n5380 VSS.n2136 0.214786
R3889 VSS.n2135 VSS.n2133 0.214786
R3890 VSS.n5384 VSS.n2132 0.214786
R3891 VSS.n5385 VSS.n2131 0.214786
R3892 VSS.n5386 VSS.n2130 0.214786
R3893 VSS.n2129 VSS.n2126 0.214786
R3894 VSS.n5391 VSS.n2125 0.214786
R3895 VSS.n5392 VSS.n2124 0.214786
R3896 VSS.n5393 VSS.n2123 0.214786
R3897 VSS.n2122 VSS.n2120 0.214786
R3898 VSS.n5397 VSS.n2119 0.214786
R3899 VSS.n5398 VSS.n2118 0.214786
R3900 VSS.n4534 VSS.n4533 0.214786
R3901 VSS.n2543 VSS.n2542 0.214786
R3902 VSS.n4539 VSS.n4538 0.214786
R3903 VSS.n4540 VSS.n2541 0.214786
R3904 VSS.n4542 VSS.n4541 0.214786
R3905 VSS.n2539 VSS.n2538 0.214786
R3906 VSS.n4548 VSS.n4547 0.214786
R3907 VSS.n4549 VSS.n2537 0.214786
R3908 VSS.n4551 VSS.n4550 0.214786
R3909 VSS.n2535 VSS.n2534 0.214786
R3910 VSS.n4556 VSS.n4555 0.214786
R3911 VSS.n4557 VSS.n2533 0.214786
R3912 VSS.n4662 VSS.n4558 0.214786
R3913 VSS.n4661 VSS.n4559 0.214786
R3914 VSS.n4660 VSS.n4560 0.214786
R3915 VSS.n4563 VSS.n4561 0.214786
R3916 VSS.n4656 VSS.n4564 0.214786
R3917 VSS.n4655 VSS.n4565 0.214786
R3918 VSS.n4654 VSS.n4566 0.214786
R3919 VSS.n4569 VSS.n4567 0.214786
R3920 VSS.n4650 VSS.n4570 0.214786
R3921 VSS.n4649 VSS.n4571 0.214786
R3922 VSS.n4648 VSS.n4572 0.214786
R3923 VSS.n4576 VSS.n4573 0.214786
R3924 VSS.n4644 VSS.n4577 0.214786
R3925 VSS.n4643 VSS.n4578 0.214786
R3926 VSS.n4642 VSS.n4579 0.214786
R3927 VSS.n4582 VSS.n4580 0.214786
R3928 VSS.n4638 VSS.n4583 0.214786
R3929 VSS.n4637 VSS.n4584 0.214786
R3930 VSS.n4636 VSS.n4585 0.214786
R3931 VSS.n4588 VSS.n4586 0.214786
R3932 VSS.n4632 VSS.n4589 0.214786
R3933 VSS.n4631 VSS.n4590 0.214786
R3934 VSS.n4630 VSS.n4591 0.214786
R3935 VSS.n4594 VSS.n4592 0.214786
R3936 VSS.n4626 VSS.n4595 0.214786
R3937 VSS.n4625 VSS.n4596 0.214786
R3938 VSS.n4624 VSS.n4597 0.214786
R3939 VSS.n4600 VSS.n4598 0.214786
R3940 VSS.n4620 VSS.n4601 0.214786
R3941 VSS.n4619 VSS.n4602 0.214786
R3942 VSS.n4618 VSS.n4603 0.214786
R3943 VSS.n4606 VSS.n4604 0.214786
R3944 VSS.n4614 VSS.n4607 0.214786
R3945 VSS.n4613 VSS.n4608 0.214786
R3946 VSS.n4612 VSS.n4610 0.214786
R3947 VSS.n4609 VSS.n2116 0.214786
R3948 VSS.n5399 VSS.n2117 0.214786
R3949 VSS.n1031 VSS.n1028 0.214786
R3950 VSS.n1027 VSS.n1026 0.214786
R3951 VSS.n1035 VSS.n1025 0.214786
R3952 VSS.n1036 VSS.n1024 0.214786
R3953 VSS.n1023 VSS.n1022 0.214786
R3954 VSS.n1040 VSS.n1021 0.214786
R3955 VSS.n1041 VSS.n1020 0.214786
R3956 VSS.n1042 VSS.n1019 0.214786
R3957 VSS.n1018 VSS.n1016 0.214786
R3958 VSS.n1046 VSS.n1015 0.214786
R3959 VSS.n1047 VSS.n1014 0.214786
R3960 VSS.n1048 VSS.n1013 0.214786
R3961 VSS.n1011 VSS.n1010 0.214786
R3962 VSS.n1053 VSS.n1052 0.214786
R3963 VSS.n1009 VSS.n1008 0.214786
R3964 VSS.n102 VSS.n101 0.214786
R3965 VSS.n1001 VSS.n1000 0.214786
R3966 VSS.n999 VSS.n107 0.214786
R3967 VSS.n998 VSS.n997 0.214786
R3968 VSS.n109 VSS.n108 0.214786
R3969 VSS.n993 VSS.n992 0.214786
R3970 VSS.n991 VSS.n111 0.214786
R3971 VSS.n990 VSS.n989 0.214786
R3972 VSS.n113 VSS.n112 0.214786
R3973 VSS.n985 VSS.n984 0.214786
R3974 VSS.n983 VSS.n115 0.214786
R3975 VSS.n982 VSS.n981 0.214786
R3976 VSS.n117 VSS.n116 0.214786
R3977 VSS.n977 VSS.n976 0.214786
R3978 VSS.n975 VSS.n119 0.214786
R3979 VSS.n974 VSS.n973 0.214786
R3980 VSS.n121 VSS.n120 0.214786
R3981 VSS.n969 VSS.n968 0.214786
R3982 VSS.n967 VSS.n123 0.214786
R3983 VSS.n966 VSS.n965 0.214786
R3984 VSS.n125 VSS.n124 0.214786
R3985 VSS.n960 VSS.n959 0.214786
R3986 VSS.n958 VSS.n127 0.214786
R3987 VSS.n956 VSS.n955 0.214786
R3988 VSS.n130 VSS.n129 0.214786
R3989 VSS.n456 VSS.n455 0.214786
R3990 VSS.n459 VSS.n454 0.214786
R3991 VSS.n460 VSS.n453 0.214786
R3992 VSS.n461 VSS.n452 0.214786
R3993 VSS.n451 VSS.n449 0.214786
R3994 VSS.n465 VSS.n448 0.214786
R3995 VSS.n466 VSS.n447 0.214786
R3996 VSS.n467 VSS.n446 0.214786
R3997 VSS.n445 VSS.n443 0.214786
R3998 VSS.n471 VSS.n442 0.214786
R3999 VSS.n472 VSS.n441 0.214786
R4000 VSS.n473 VSS.n440 0.214786
R4001 VSS.n439 VSS.n437 0.214786
R4002 VSS.n477 VSS.n436 0.214786
R4003 VSS.n478 VSS.n435 0.214786
R4004 VSS.n479 VSS.n434 0.214786
R4005 VSS.n433 VSS.n431 0.214786
R4006 VSS.n483 VSS.n430 0.214786
R4007 VSS.n484 VSS.n429 0.214786
R4008 VSS.n485 VSS.n428 0.214786
R4009 VSS.n427 VSS.n424 0.214786
R4010 VSS.n489 VSS.n423 0.214786
R4011 VSS.n491 VSS.n422 0.214786
R4012 VSS.n492 VSS.n421 0.214786
R4013 VSS.n420 VSS.n418 0.214786
R4014 VSS.n496 VSS.n417 0.214786
R4015 VSS.n497 VSS.n416 0.214786
R4016 VSS.n415 VSS.n414 0.214786
R4017 VSS.n501 VSS.n413 0.214786
R4018 VSS.n502 VSS.n412 0.214786
R4019 VSS.n503 VSS.n411 0.214786
R4020 VSS.n410 VSS.n408 0.214786
R4021 VSS.n507 VSS.n407 0.214786
R4022 VSS.n508 VSS.n406 0.214786
R4023 VSS.n509 VSS.n405 0.214786
R4024 VSS.n404 VSS.n402 0.214786
R4025 VSS.n513 VSS.n401 0.214786
R4026 VSS.n514 VSS.n400 0.214786
R4027 VSS.n515 VSS.n399 0.214786
R4028 VSS.n398 VSS.n396 0.214786
R4029 VSS.n519 VSS.n395 0.214786
R4030 VSS.n520 VSS.n394 0.214786
R4031 VSS.n521 VSS.n393 0.214786
R4032 VSS.n392 VSS.n390 0.214786
R4033 VSS.n576 VSS.n388 0.214786
R4034 VSS.n575 VSS.n389 0.214786
R4035 VSS.n1136 VSS.n1135 0.214786
R4036 VSS.n80 VSS.n79 0.214786
R4037 VSS.n1131 VSS.n1130 0.214786
R4038 VSS.n1129 VSS.n82 0.214786
R4039 VSS.n1128 VSS.n1127 0.214786
R4040 VSS.n84 VSS.n83 0.214786
R4041 VSS.n1123 VSS.n1122 0.214786
R4042 VSS.n1121 VSS.n86 0.214786
R4043 VSS.n1120 VSS.n1119 0.214786
R4044 VSS.n88 VSS.n87 0.214786
R4045 VSS.n1115 VSS.n1114 0.214786
R4046 VSS.n1113 VSS.n90 0.214786
R4047 VSS.n1112 VSS.n1111 0.214786
R4048 VSS.n92 VSS.n91 0.214786
R4049 VSS.n1106 VSS.n97 0.214786
R4050 VSS.n168 VSS.n96 0.214786
R4051 VSS.n919 VSS.n169 0.214786
R4052 VSS.n920 VSS.n167 0.214786
R4053 VSS.n921 VSS.n166 0.214786
R4054 VSS.n165 VSS.n163 0.214786
R4055 VSS.n925 VSS.n162 0.214786
R4056 VSS.n926 VSS.n161 0.214786
R4057 VSS.n927 VSS.n160 0.214786
R4058 VSS.n159 VSS.n157 0.214786
R4059 VSS.n931 VSS.n156 0.214786
R4060 VSS.n932 VSS.n155 0.214786
R4061 VSS.n933 VSS.n154 0.214786
R4062 VSS.n153 VSS.n151 0.214786
R4063 VSS.n937 VSS.n150 0.214786
R4064 VSS.n938 VSS.n149 0.214786
R4065 VSS.n939 VSS.n148 0.214786
R4066 VSS.n147 VSS.n145 0.214786
R4067 VSS.n943 VSS.n144 0.214786
R4068 VSS.n944 VSS.n143 0.214786
R4069 VSS.n142 VSS.n140 0.214786
R4070 VSS.n948 VSS.n139 0.214786
R4071 VSS.n949 VSS.n138 0.214786
R4072 VSS.n950 VSS.n137 0.214786
R4073 VSS.n805 VSS.n804 0.214786
R4074 VSS.n807 VSS.n803 0.214786
R4075 VSS.n808 VSS.n802 0.214786
R4076 VSS.n809 VSS.n801 0.214786
R4077 VSS.n800 VSS.n798 0.214786
R4078 VSS.n813 VSS.n797 0.214786
R4079 VSS.n814 VSS.n796 0.214786
R4080 VSS.n815 VSS.n795 0.214786
R4081 VSS.n794 VSS.n792 0.214786
R4082 VSS.n819 VSS.n791 0.214786
R4083 VSS.n820 VSS.n790 0.214786
R4084 VSS.n821 VSS.n789 0.214786
R4085 VSS.n788 VSS.n308 0.214786
R4086 VSS.n787 VSS.n786 0.214786
R4087 VSS.n310 VSS.n309 0.214786
R4088 VSS.n782 VSS.n781 0.214786
R4089 VSS.n780 VSS.n312 0.214786
R4090 VSS.n779 VSS.n778 0.214786
R4091 VSS.n314 VSS.n313 0.214786
R4092 VSS.n774 VSS.n773 0.214786
R4093 VSS.n772 VSS.n316 0.214786
R4094 VSS.n771 VSS.n770 0.214786
R4095 VSS.n318 VSS.n317 0.214786
R4096 VSS.n766 VSS.n765 0.214786
R4097 VSS.n763 VSS.n762 0.214786
R4098 VSS.n324 VSS.n323 0.214786
R4099 VSS.n758 VSS.n757 0.214786
R4100 VSS.n756 VSS.n326 0.214786
R4101 VSS.n755 VSS.n754 0.214786
R4102 VSS.n328 VSS.n327 0.214786
R4103 VSS.n608 VSS.n606 0.214786
R4104 VSS.n609 VSS.n605 0.214786
R4105 VSS.n610 VSS.n604 0.214786
R4106 VSS.n603 VSS.n601 0.214786
R4107 VSS.n614 VSS.n600 0.214786
R4108 VSS.n615 VSS.n599 0.214786
R4109 VSS.n616 VSS.n598 0.214786
R4110 VSS.n597 VSS.n595 0.214786
R4111 VSS.n620 VSS.n594 0.214786
R4112 VSS.n621 VSS.n593 0.214786
R4113 VSS.n622 VSS.n592 0.214786
R4114 VSS.n591 VSS.n589 0.214786
R4115 VSS.n626 VSS.n588 0.214786
R4116 VSS.n627 VSS.n587 0.214786
R4117 VSS.n628 VSS.n586 0.214786
R4118 VSS.n585 VSS.n369 0.214786
R4119 VSS.n584 VSS.n583 0.214786
R4120 VSS.n371 VSS.n370 0.214786
R4121 VSS.n1082 VSS.n1077 0.214786
R4122 VSS.n1076 VSS.n1074 0.214786
R4123 VSS.n1086 VSS.n1073 0.214786
R4124 VSS.n1087 VSS.n1072 0.214786
R4125 VSS.n1071 VSS.n1070 0.214786
R4126 VSS.n1091 VSS.n1069 0.214786
R4127 VSS.n1092 VSS.n1068 0.214786
R4128 VSS.n1093 VSS.n1067 0.214786
R4129 VSS.n1066 VSS.n1064 0.214786
R4130 VSS.n1097 VSS.n1063 0.214786
R4131 VSS.n1098 VSS.n1062 0.214786
R4132 VSS.n1099 VSS.n1061 0.214786
R4133 VSS.n1060 VSS.n1058 0.214786
R4134 VSS.n1103 VSS.n1057 0.214786
R4135 VSS.n100 VSS.n99 0.214786
R4136 VSS.n898 VSS.n897 0.214786
R4137 VSS.n899 VSS.n896 0.214786
R4138 VSS.n895 VSS.n267 0.214786
R4139 VSS.n894 VSS.n893 0.214786
R4140 VSS.n269 VSS.n268 0.214786
R4141 VSS.n889 VSS.n888 0.214786
R4142 VSS.n887 VSS.n271 0.214786
R4143 VSS.n886 VSS.n885 0.214786
R4144 VSS.n273 VSS.n272 0.214786
R4145 VSS.n881 VSS.n880 0.214786
R4146 VSS.n879 VSS.n275 0.214786
R4147 VSS.n878 VSS.n877 0.214786
R4148 VSS.n277 VSS.n276 0.214786
R4149 VSS.n873 VSS.n872 0.214786
R4150 VSS.n871 VSS.n279 0.214786
R4151 VSS.n870 VSS.n869 0.214786
R4152 VSS.n281 VSS.n280 0.214786
R4153 VSS.n865 VSS.n864 0.214786
R4154 VSS.n863 VSS.n284 0.214786
R4155 VSS.n862 VSS.n861 0.214786
R4156 VSS.n286 VSS.n285 0.214786
R4157 VSS.n856 VSS.n855 0.214786
R4158 VSS.n854 VSS.n288 0.214786
R4159 VSS.n852 VSS.n851 0.214786
R4160 VSS.n290 VSS.n289 0.214786
R4161 VSS.n847 VSS.n846 0.214786
R4162 VSS.n845 VSS.n293 0.214786
R4163 VSS.n844 VSS.n843 0.214786
R4164 VSS.n295 VSS.n294 0.214786
R4165 VSS.n839 VSS.n838 0.214786
R4166 VSS.n837 VSS.n297 0.214786
R4167 VSS.n836 VSS.n835 0.214786
R4168 VSS.n299 VSS.n298 0.214786
R4169 VSS.n831 VSS.n830 0.214786
R4170 VSS.n829 VSS.n301 0.214786
R4171 VSS.n828 VSS.n827 0.214786
R4172 VSS.n303 VSS.n302 0.214786
R4173 VSS.n728 VSS.n727 0.214786
R4174 VSS.n729 VSS.n726 0.214786
R4175 VSS.n725 VSS.n723 0.214786
R4176 VSS.n733 VSS.n722 0.214786
R4177 VSS.n734 VSS.n721 0.214786
R4178 VSS.n735 VSS.n720 0.214786
R4179 VSS.n719 VSS.n717 0.214786
R4180 VSS.n739 VSS.n716 0.214786
R4181 VSS.n740 VSS.n715 0.214786
R4182 VSS.n741 VSS.n714 0.214786
R4183 VSS.n711 VSS.n710 0.214786
R4184 VSS.n746 VSS.n709 0.214786
R4185 VSS.n747 VSS.n708 0.214786
R4186 VSS.n748 VSS.n707 0.214786
R4187 VSS.n706 VSS.n333 0.214786
R4188 VSS.n705 VSS.n704 0.214786
R4189 VSS.n335 VSS.n334 0.214786
R4190 VSS.n700 VSS.n699 0.214786
R4191 VSS.n698 VSS.n337 0.214786
R4192 VSS.n697 VSS.n696 0.214786
R4193 VSS.n339 VSS.n338 0.214786
R4194 VSS.n692 VSS.n691 0.214786
R4195 VSS.n690 VSS.n341 0.214786
R4196 VSS.n689 VSS.n688 0.214786
R4197 VSS.n343 VSS.n342 0.214786
R4198 VSS.n684 VSS.n683 0.214786
R4199 VSS.n682 VSS.n345 0.214786
R4200 VSS.n681 VSS.n680 0.214786
R4201 VSS.n347 VSS.n346 0.214786
R4202 VSS.n676 VSS.n675 0.214786
R4203 VSS.n674 VSS.n349 0.214786
R4204 VSS.n673 VSS.n672 0.214786
R4205 VSS.n351 VSS.n350 0.214786
R4206 VSS.n384 VSS.n383 0.214786
R4207 VSS.n333 VSS.n331 0.214786
R4208 VSS.n1081 VSS.n1075 0.214786
R4209 VSS.n1083 VSS.n1082 0.214786
R4210 VSS.n1084 VSS.n1074 0.214786
R4211 VSS.n1086 VSS.n1085 0.214786
R4212 VSS.n1088 VSS.n1087 0.214786
R4213 VSS.n1089 VSS.n1070 0.214786
R4214 VSS.n1091 VSS.n1090 0.214786
R4215 VSS.n1092 VSS.n1065 0.214786
R4216 VSS.n1094 VSS.n1093 0.214786
R4217 VSS.n1095 VSS.n1064 0.214786
R4218 VSS.n1097 VSS.n1096 0.214786
R4219 VSS.n1098 VSS.n1059 0.214786
R4220 VSS.n1100 VSS.n1099 0.214786
R4221 VSS.n1101 VSS.n1058 0.214786
R4222 VSS.n1103 VSS.n1102 0.214786
R4223 VSS.n264 VSS.n99 0.214786
R4224 VSS.n898 VSS.n266 0.214786
R4225 VSS.n900 VSS.n899 0.214786
R4226 VSS.n267 VSS.n263 0.214786
R4227 VSS.n893 VSS.n892 0.214786
R4228 VSS.n891 VSS.n269 0.214786
R4229 VSS.n890 VSS.n889 0.214786
R4230 VSS.n271 VSS.n270 0.214786
R4231 VSS.n885 VSS.n884 0.214786
R4232 VSS.n883 VSS.n273 0.214786
R4233 VSS.n882 VSS.n881 0.214786
R4234 VSS.n275 VSS.n274 0.214786
R4235 VSS.n877 VSS.n876 0.214786
R4236 VSS.n875 VSS.n277 0.214786
R4237 VSS.n874 VSS.n873 0.214786
R4238 VSS.n279 VSS.n278 0.214786
R4239 VSS.n869 VSS.n868 0.214786
R4240 VSS.n867 VSS.n281 0.214786
R4241 VSS.n866 VSS.n865 0.214786
R4242 VSS.n859 VSS.n284 0.214786
R4243 VSS.n861 VSS.n860 0.214786
R4244 VSS.n858 VSS.n286 0.214786
R4245 VSS.n857 VSS.n856 0.214786
R4246 VSS.n288 VSS.n287 0.214786
R4247 VSS.n851 VSS.n850 0.214786
R4248 VSS.n849 VSS.n290 0.214786
R4249 VSS.n848 VSS.n847 0.214786
R4250 VSS.n293 VSS.n292 0.214786
R4251 VSS.n843 VSS.n842 0.214786
R4252 VSS.n841 VSS.n295 0.214786
R4253 VSS.n840 VSS.n839 0.214786
R4254 VSS.n297 VSS.n296 0.214786
R4255 VSS.n835 VSS.n834 0.214786
R4256 VSS.n833 VSS.n299 0.214786
R4257 VSS.n832 VSS.n831 0.214786
R4258 VSS.n301 VSS.n300 0.214786
R4259 VSS.n827 VSS.n826 0.214786
R4260 VSS.n304 VSS.n303 0.214786
R4261 VSS.n728 VSS.n724 0.214786
R4262 VSS.n730 VSS.n729 0.214786
R4263 VSS.n731 VSS.n723 0.214786
R4264 VSS.n733 VSS.n732 0.214786
R4265 VSS.n734 VSS.n718 0.214786
R4266 VSS.n736 VSS.n735 0.214786
R4267 VSS.n737 VSS.n717 0.214786
R4268 VSS.n739 VSS.n738 0.214786
R4269 VSS.n740 VSS.n712 0.214786
R4270 VSS.n742 VSS.n741 0.214786
R4271 VSS.n744 VSS.n711 0.214786
R4272 VSS.n746 VSS.n745 0.214786
R4273 VSS.n747 VSS.n332 0.214786
R4274 VSS.n749 VSS.n748 0.214786
R4275 VSS.n704 VSS.n703 0.214786
R4276 VSS.n702 VSS.n335 0.214786
R4277 VSS.n701 VSS.n700 0.214786
R4278 VSS.n337 VSS.n336 0.214786
R4279 VSS.n696 VSS.n695 0.214786
R4280 VSS.n694 VSS.n339 0.214786
R4281 VSS.n693 VSS.n692 0.214786
R4282 VSS.n341 VSS.n340 0.214786
R4283 VSS.n688 VSS.n687 0.214786
R4284 VSS.n686 VSS.n343 0.214786
R4285 VSS.n685 VSS.n684 0.214786
R4286 VSS.n345 VSS.n344 0.214786
R4287 VSS.n680 VSS.n679 0.214786
R4288 VSS.n678 VSS.n347 0.214786
R4289 VSS.n677 VSS.n676 0.214786
R4290 VSS.n349 VSS.n348 0.214786
R4291 VSS.n672 VSS.n671 0.214786
R4292 VSS.n352 VSS.n351 0.214786
R4293 VSS.n383 VSS.n382 0.214786
R4294 VSS.n78 VSS.n57 0.214786
R4295 VSS.n1135 VSS.n1134 0.214786
R4296 VSS.n1133 VSS.n80 0.214786
R4297 VSS.n1132 VSS.n1131 0.214786
R4298 VSS.n82 VSS.n81 0.214786
R4299 VSS.n1127 VSS.n1126 0.214786
R4300 VSS.n1125 VSS.n84 0.214786
R4301 VSS.n1124 VSS.n1123 0.214786
R4302 VSS.n86 VSS.n85 0.214786
R4303 VSS.n1119 VSS.n1118 0.214786
R4304 VSS.n1117 VSS.n88 0.214786
R4305 VSS.n1116 VSS.n1115 0.214786
R4306 VSS.n90 VSS.n89 0.214786
R4307 VSS.n1111 VSS.n1110 0.214786
R4308 VSS.n1109 VSS.n92 0.214786
R4309 VSS.n1107 VSS.n1106 0.214786
R4310 VSS.n917 VSS.n96 0.214786
R4311 VSS.n919 VSS.n918 0.214786
R4312 VSS.n920 VSS.n164 0.214786
R4313 VSS.n922 VSS.n921 0.214786
R4314 VSS.n923 VSS.n163 0.214786
R4315 VSS.n925 VSS.n924 0.214786
R4316 VSS.n926 VSS.n158 0.214786
R4317 VSS.n928 VSS.n927 0.214786
R4318 VSS.n929 VSS.n157 0.214786
R4319 VSS.n931 VSS.n930 0.214786
R4320 VSS.n932 VSS.n152 0.214786
R4321 VSS.n934 VSS.n933 0.214786
R4322 VSS.n935 VSS.n151 0.214786
R4323 VSS.n937 VSS.n936 0.214786
R4324 VSS.n938 VSS.n146 0.214786
R4325 VSS.n940 VSS.n939 0.214786
R4326 VSS.n941 VSS.n145 0.214786
R4327 VSS.n943 VSS.n942 0.214786
R4328 VSS.n945 VSS.n944 0.214786
R4329 VSS.n946 VSS.n140 0.214786
R4330 VSS.n948 VSS.n947 0.214786
R4331 VSS.n949 VSS.n135 0.214786
R4332 VSS.n951 VSS.n950 0.214786
R4333 VSS.n805 VSS.n134 0.214786
R4334 VSS.n807 VSS.n806 0.214786
R4335 VSS.n808 VSS.n799 0.214786
R4336 VSS.n810 VSS.n809 0.214786
R4337 VSS.n811 VSS.n798 0.214786
R4338 VSS.n813 VSS.n812 0.214786
R4339 VSS.n814 VSS.n793 0.214786
R4340 VSS.n816 VSS.n815 0.214786
R4341 VSS.n817 VSS.n792 0.214786
R4342 VSS.n819 VSS.n818 0.214786
R4343 VSS.n820 VSS.n307 0.214786
R4344 VSS.n822 VSS.n821 0.214786
R4345 VSS.n308 VSS.n306 0.214786
R4346 VSS.n786 VSS.n785 0.214786
R4347 VSS.n784 VSS.n310 0.214786
R4348 VSS.n783 VSS.n782 0.214786
R4349 VSS.n312 VSS.n311 0.214786
R4350 VSS.n778 VSS.n777 0.214786
R4351 VSS.n776 VSS.n314 0.214786
R4352 VSS.n775 VSS.n774 0.214786
R4353 VSS.n316 VSS.n315 0.214786
R4354 VSS.n770 VSS.n769 0.214786
R4355 VSS.n768 VSS.n318 0.214786
R4356 VSS.n767 VSS.n766 0.214786
R4357 VSS.n762 VSS.n761 0.214786
R4358 VSS.n760 VSS.n324 0.214786
R4359 VSS.n759 VSS.n758 0.214786
R4360 VSS.n326 VSS.n325 0.214786
R4361 VSS.n754 VSS.n753 0.214786
R4362 VSS.n329 VSS.n328 0.214786
R4363 VSS.n608 VSS.n607 0.214786
R4364 VSS.n609 VSS.n602 0.214786
R4365 VSS.n611 VSS.n610 0.214786
R4366 VSS.n612 VSS.n601 0.214786
R4367 VSS.n614 VSS.n613 0.214786
R4368 VSS.n615 VSS.n596 0.214786
R4369 VSS.n617 VSS.n616 0.214786
R4370 VSS.n618 VSS.n595 0.214786
R4371 VSS.n620 VSS.n619 0.214786
R4372 VSS.n621 VSS.n590 0.214786
R4373 VSS.n623 VSS.n622 0.214786
R4374 VSS.n624 VSS.n589 0.214786
R4375 VSS.n626 VSS.n625 0.214786
R4376 VSS.n627 VSS.n368 0.214786
R4377 VSS.n629 VSS.n628 0.214786
R4378 VSS.n369 VSS.n367 0.214786
R4379 VSS.n583 VSS.n582 0.214786
R4380 VSS.n580 VSS.n371 0.214786
R4381 VSS.n1030 VSS.n36 0.214786
R4382 VSS.n1032 VSS.n1031 0.214786
R4383 VSS.n1033 VSS.n1026 0.214786
R4384 VSS.n1035 VSS.n1034 0.214786
R4385 VSS.n1037 VSS.n1036 0.214786
R4386 VSS.n1038 VSS.n1022 0.214786
R4387 VSS.n1040 VSS.n1039 0.214786
R4388 VSS.n1041 VSS.n1017 0.214786
R4389 VSS.n1043 VSS.n1042 0.214786
R4390 VSS.n1044 VSS.n1016 0.214786
R4391 VSS.n1046 VSS.n1045 0.214786
R4392 VSS.n1047 VSS.n1012 0.214786
R4393 VSS.n1049 VSS.n1048 0.214786
R4394 VSS.n1050 VSS.n1011 0.214786
R4395 VSS.n1052 VSS.n1051 0.214786
R4396 VSS.n1008 VSS.n1007 0.214786
R4397 VSS.n103 VSS.n102 0.214786
R4398 VSS.n1002 VSS.n1001 0.214786
R4399 VSS.n107 VSS.n106 0.214786
R4400 VSS.n997 VSS.n996 0.214786
R4401 VSS.n995 VSS.n109 0.214786
R4402 VSS.n994 VSS.n993 0.214786
R4403 VSS.n111 VSS.n110 0.214786
R4404 VSS.n989 VSS.n988 0.214786
R4405 VSS.n987 VSS.n113 0.214786
R4406 VSS.n986 VSS.n985 0.214786
R4407 VSS.n115 VSS.n114 0.214786
R4408 VSS.n981 VSS.n980 0.214786
R4409 VSS.n979 VSS.n117 0.214786
R4410 VSS.n978 VSS.n977 0.214786
R4411 VSS.n119 VSS.n118 0.214786
R4412 VSS.n973 VSS.n972 0.214786
R4413 VSS.n971 VSS.n121 0.214786
R4414 VSS.n970 VSS.n969 0.214786
R4415 VSS.n963 VSS.n123 0.214786
R4416 VSS.n965 VSS.n964 0.214786
R4417 VSS.n962 VSS.n125 0.214786
R4418 VSS.n961 VSS.n960 0.214786
R4419 VSS.n127 VSS.n126 0.214786
R4420 VSS.n955 VSS.n954 0.214786
R4421 VSS.n132 VSS.n130 0.214786
R4422 VSS.n457 VSS.n456 0.214786
R4423 VSS.n459 VSS.n458 0.214786
R4424 VSS.n460 VSS.n450 0.214786
R4425 VSS.n462 VSS.n461 0.214786
R4426 VSS.n463 VSS.n449 0.214786
R4427 VSS.n465 VSS.n464 0.214786
R4428 VSS.n466 VSS.n444 0.214786
R4429 VSS.n468 VSS.n467 0.214786
R4430 VSS.n469 VSS.n443 0.214786
R4431 VSS.n471 VSS.n470 0.214786
R4432 VSS.n472 VSS.n438 0.214786
R4433 VSS.n474 VSS.n473 0.214786
R4434 VSS.n475 VSS.n437 0.214786
R4435 VSS.n477 VSS.n476 0.214786
R4436 VSS.n478 VSS.n432 0.214786
R4437 VSS.n480 VSS.n479 0.214786
R4438 VSS.n481 VSS.n431 0.214786
R4439 VSS.n483 VSS.n482 0.214786
R4440 VSS.n484 VSS.n426 0.214786
R4441 VSS.n486 VSS.n485 0.214786
R4442 VSS.n487 VSS.n424 0.214786
R4443 VSS.n489 VSS.n488 0.214786
R4444 VSS.n491 VSS.n419 0.214786
R4445 VSS.n493 VSS.n492 0.214786
R4446 VSS.n494 VSS.n418 0.214786
R4447 VSS.n496 VSS.n495 0.214786
R4448 VSS.n498 VSS.n497 0.214786
R4449 VSS.n499 VSS.n414 0.214786
R4450 VSS.n501 VSS.n500 0.214786
R4451 VSS.n502 VSS.n409 0.214786
R4452 VSS.n504 VSS.n503 0.214786
R4453 VSS.n505 VSS.n408 0.214786
R4454 VSS.n507 VSS.n506 0.214786
R4455 VSS.n508 VSS.n403 0.214786
R4456 VSS.n510 VSS.n509 0.214786
R4457 VSS.n511 VSS.n402 0.214786
R4458 VSS.n513 VSS.n512 0.214786
R4459 VSS.n514 VSS.n397 0.214786
R4460 VSS.n516 VSS.n515 0.214786
R4461 VSS.n517 VSS.n396 0.214786
R4462 VSS.n519 VSS.n518 0.214786
R4463 VSS.n520 VSS.n391 0.214786
R4464 VSS.n522 VSS.n521 0.214786
R4465 VSS.n573 VSS.n390 0.214786
R4466 VSS.n577 VSS.n576 0.214786
R4467 VSS.n575 VSS.n574 0.214786
R4468 VSS.n4543 VSS.n4542 0.214786
R4469 VSS.n2169 VSS.n2164 0.214786
R4470 VSS.n2171 VSS.n2170 0.214786
R4471 VSS.n2163 VSS.n2162 0.214786
R4472 VSS.n5355 VSS.n5354 0.214786
R4473 VSS.n5356 VSS.n2157 0.214786
R4474 VSS.n5358 VSS.n5357 0.214786
R4475 VSS.n5359 VSS.n2156 0.214786
R4476 VSS.n5361 VSS.n5360 0.214786
R4477 VSS.n5362 VSS.n2151 0.214786
R4478 VSS.n5364 VSS.n5363 0.214786
R4479 VSS.n5365 VSS.n2150 0.214786
R4480 VSS.n5367 VSS.n5366 0.214786
R4481 VSS.n5368 VSS.n2145 0.214786
R4482 VSS.n5370 VSS.n5369 0.214786
R4483 VSS.n5371 VSS.n2144 0.214786
R4484 VSS.n5373 VSS.n5372 0.214786
R4485 VSS.n5374 VSS.n2139 0.214786
R4486 VSS.n5376 VSS.n5375 0.214786
R4487 VSS.n5377 VSS.n2138 0.214786
R4488 VSS.n5379 VSS.n5378 0.214786
R4489 VSS.n5381 VSS.n5380 0.214786
R4490 VSS.n5382 VSS.n2133 0.214786
R4491 VSS.n5384 VSS.n5383 0.214786
R4492 VSS.n5385 VSS.n2128 0.214786
R4493 VSS.n5387 VSS.n5386 0.214786
R4494 VSS.n5388 VSS.n2126 0.214786
R4495 VSS.n5398 VSS.n2115 0.214786
R4496 VSS.n5397 VSS.n5396 0.214786
R4497 VSS.n5395 VSS.n2120 0.214786
R4498 VSS.n5394 VSS.n5393 0.214786
R4499 VSS.n5392 VSS.n2121 0.214786
R4500 VSS.n5391 VSS.n5390 0.214786
R4501 VSS.n2545 VSS.n2544 0.214786
R4502 VSS.n4535 VSS.n4534 0.214786
R4503 VSS.n4536 VSS.n2543 0.214786
R4504 VSS.n4538 VSS.n4537 0.214786
R4505 VSS.n2541 VSS.n2540 0.214786
R4506 VSS.n4545 VSS.n2539 0.214786
R4507 VSS.n4547 VSS.n4546 0.214786
R4508 VSS.n2537 VSS.n2536 0.214786
R4509 VSS.n4552 VSS.n4551 0.214786
R4510 VSS.n4553 VSS.n2535 0.214786
R4511 VSS.n4555 VSS.n4554 0.214786
R4512 VSS.n2533 VSS.n2531 0.214786
R4513 VSS.n4663 VSS.n4662 0.214786
R4514 VSS.n4661 VSS.n2532 0.214786
R4515 VSS.n4660 VSS.n4659 0.214786
R4516 VSS.n4658 VSS.n4561 0.214786
R4517 VSS.n4657 VSS.n4656 0.214786
R4518 VSS.n4655 VSS.n4562 0.214786
R4519 VSS.n4654 VSS.n4653 0.214786
R4520 VSS.n4652 VSS.n4567 0.214786
R4521 VSS.n4651 VSS.n4650 0.214786
R4522 VSS.n4649 VSS.n4568 0.214786
R4523 VSS.n4648 VSS.n4647 0.214786
R4524 VSS.n4646 VSS.n4573 0.214786
R4525 VSS.n4645 VSS.n4644 0.214786
R4526 VSS.n4643 VSS.n4575 0.214786
R4527 VSS.n4642 VSS.n4641 0.214786
R4528 VSS.n4640 VSS.n4580 0.214786
R4529 VSS.n4639 VSS.n4638 0.214786
R4530 VSS.n4637 VSS.n4581 0.214786
R4531 VSS.n4636 VSS.n4635 0.214786
R4532 VSS.n4634 VSS.n4586 0.214786
R4533 VSS.n4633 VSS.n4632 0.214786
R4534 VSS.n4631 VSS.n4587 0.214786
R4535 VSS.n4630 VSS.n4629 0.214786
R4536 VSS.n4628 VSS.n4592 0.214786
R4537 VSS.n4627 VSS.n4626 0.214786
R4538 VSS.n4625 VSS.n4593 0.214786
R4539 VSS.n4624 VSS.n4623 0.214786
R4540 VSS.n4622 VSS.n4598 0.214786
R4541 VSS.n4621 VSS.n4620 0.214786
R4542 VSS.n4619 VSS.n4599 0.214786
R4543 VSS.n4618 VSS.n4617 0.214786
R4544 VSS.n4616 VSS.n4604 0.214786
R4545 VSS.n4615 VSS.n4614 0.214786
R4546 VSS.n4613 VSS.n4605 0.214786
R4547 VSS.n4612 VSS.n4611 0.214786
R4548 VSS.n2116 VSS.n2114 0.214786
R4549 VSS.n5400 VSS.n5399 0.214786
R4550 VSS.n5436 VSS.n2084 0.212265
R4551 VSS.n5696 VSS.n5695 0.201836
R4552 VSS.n5175 DVSS 0.194818
R4553 VSS.n5445 VSS.n5444 0.192412
R4554 VSS VSS.n3615 0.189765
R4555 VSS.n3615 VSS 0.189765
R4556 VSS.n5330 VSS.n5329 0.186214
R4557 VSS.n5331 VSS.n5330 0.186214
R4558 VSS.n4669 VSS.n4668 0.186214
R4559 VSS.n4670 VSS.n4669 0.186214
R4560 VSS.n1590 VSS.n1589 0.185484
R4561 VSS VSS.n4303 0.17855
R4562 VSS.n2232 VSS.n2231 0.178408
R4563 VSS.n2231 VSS.n2230 0.178408
R4564 VSS.n5284 VSS.n5282 0.178408
R4565 VSS.n2231 VSS.n2229 0.178408
R4566 VSS.n5284 VSS.n5283 0.178408
R4567 VSS.n2231 VSS.n2228 0.178408
R4568 VSS.n5284 VSS.n2204 0.178408
R4569 VSS.n2515 VSS.n2514 0.175807
R4570 VSS.n5259 DVSS 0.175804
R4571 VSS.n3680 DVSS 0.175804
R4572 VSS.n3623 DVSS 0.175804
R4573 VSS.n3674 DVSS 0.175804
R4574 VSS.n3562 DVSS 0.175804
R4575 VSS.n3586 DVSS 0.175804
R4576 VSS.n2726 DVSS 0.175804
R4577 VSS.n2728 DVSS 0.175804
R4578 VSS.n2696 DVSS 0.175729
R4579 VSS.n2241 DVSS 0.175729
R4580 VSS.n3518 DVSS 0.175729
R4581 VSS.n2729 DVSS 0.175729
R4582 VSS.n902 VSS.n901 0.173577
R4583 VSS.n670 VSS.n669 0.173577
R4584 VSS.n4529 DVSS 0.172116
R4585 VSS.n5352 DVSS 0.172116
R4586 VSS.n5321 DVSS 0.172116
R4587 VSS.n5402 DVSS 0.172116
R4588 VSS.n4665 DVSS 0.172116
R4589 VSS VSS.n4202 0.169912
R4590 VSS.n4284 VSS.n4277 0.168658
R4591 VSS.n4277 VSS.n2508 0.168658
R4592 VSS.n4675 VSS.n2501 0.168658
R4593 VSS.n4685 VSS.n2501 0.168658
R4594 VSS.n4673 VSS.n4672 0.166289
R4595 VSS.n282 VSS.n141 0.163909
R4596 VSS.n824 VSS.n823 0.163909
R4597 VSS.n752 VSS.n751 0.163909
R4598 VSS.n535 VSS.n365 0.161214
R4599 VSS.n217 VSS.n216 0.161214
R4600 VSS.n1141 VSS.n1140 0.149124
R4601 VSS.n3259 VSS.n3258 0.145461
R4602 VSS.n5149 DVSS 0.144526
R4603 VSS.n4213 DVSS 0.144421
R4604 VSS.n4209 DVSS 0.144187
R4605 VSS.n4212 DVSS 0.1436
R4606 DVSS VSS.n4211 0.1436
R4607 VSS.n4211 DVSS 0.1436
R4608 DVSS VSS.n4210 0.1436
R4609 DVSS VSS.n3677 0.143441
R4610 VSS.n3675 DVSS 0.143441
R4611 DVSS VSS.n2727 0.143441
R4612 VSS.n3565 DVSS 0.143441
R4613 VSS.n1004 VSS.n1003 0.141125
R4614 VSS.n572 VSS.n571 0.141125
R4615 VSS.n3677 VSS.n3676 0.140794
R4616 VSS.n3676 VSS.n3675 0.140794
R4617 VSS.n3566 VSS.n2727 0.140794
R4618 VSS.n3566 VSS.n3565 0.140794
R4619 VSS.n3609 VSS 0.139932
R4620 DVSS VSS.n5174 0.139047
R4621 VSS.n4193 DVSS 0.138622
R4622 VSS.n1005 VSS.n104 0.137596
R4623 VSS.n569 VSS.n523 0.137559
R4624 VSS.n4196 VSS 0.1355
R4625 VSS.n3528 VSS 0.1355
R4626 VSS.n2732 VSS 0.1355
R4627 VSS.n2792 VSS 0.1355
R4628 VSS.n2794 VSS 0.1355
R4629 DVSS VSS.n2101 0.1355
R4630 VSS.n2632 VSS 0.1355
R4631 VSS.n2705 DVSS 0.132383
R4632 VSS.n906 VSS.n222 0.130943
R4633 VSS.n3994 DVSS 0.130618
R4634 VSS.n380 VSS.n221 0.130587
R4635 VSS.n4381 DVSS 0.130161
R4636 VSS.n5188 DVSS 0.130161
R4637 VSS.n1302 VSS.n1297 0.129009
R4638 VSS.n3883 VSS.n3882 0.128608
R4639 VSS.n4122 VSS.n3883 0.128203
R4640 VSS.n1395 DVSS 0.125798
R4641 VSS.n5174 VSS.n5173 0.122865
R4642 VSS.n1395 VSS.n33 0.12265
R4643 VSS.n5253 DVSS 0.115647
R4644 VSS.n3820 VSS.n3786 0.114824
R4645 VSS.n4068 VSS.n3885 0.114824
R4646 VSS VSS.n2413 0.113
R4647 VSS.n3616 VSS 0.113
R4648 VSS VSS.n3252 0.113
R4649 VSS.n5149 DVSS 0.111845
R4650 VSS.n4207 DVSS 0.111373
R4651 VSS.n2168 VSS.n2166 0.110634
R4652 VSS.n1080 VSS.n1077 0.110634
R4653 VSS.n1137 VSS.n1136 0.110634
R4654 VSS.n1029 VSS.n1028 0.110634
R4655 VSS.n3524 VSS 0.110353
R4656 VSS.n4129 VSS.n3758 0.109959
R4657 VSS.n4130 VSS.n4129 0.109959
R4658 VSS.n916 VSS.n915 0.107643
R4659 VSS.n631 VSS.n630 0.107643
R4660 DVSS VSS.n4207 0.107291
R4661 VSS.n4674 VSS.n2508 0.107079
R4662 VSS.n2529 VSS.n2528 0.105895
R4663 VSS.n1584 VSS.n1302 0.102277
R4664 VSS.n4211 DVSS 0.102157
R4665 VSS.n5690 VSS.n8 0.101471
R4666 VSS.n5454 VSS.n5453 0.101471
R4667 DVSS VSS.n4381 0.101206
R4668 VSS.n5188 DVSS 0.101206
R4669 VSS.n3994 DVSS 0.10093
R4670 VSS.n5181 VSS.n5180 0.100383
R4671 DVSS VSS.n2624 0.0991804
R4672 VSS.n1589 VSS.n1296 0.0985668
R4673 VSS.n1589 VSS.n1588 0.0984658
R4674 VSS.n2516 VSS 0.0939292
R4675 VSS.n2626 VSS 0.0939292
R4676 VSS.n2628 VSS 0.0939292
R4677 VSS.n2188 VSS 0.0939292
R4678 VSS.n2190 VSS 0.0939292
R4679 VSS.n4846 VSS 0.0939292
R4680 VSS.n5175 DVSS 0.0938582
R4681 VSS.n4673 VSS 0.0928684
R4682 VSS.n2938 VSS.n2937 0.0923483
R4683 VSS.n5444 VSS.n5443 0.0891765
R4684 VSS.n5297 VSS.n5296 0.0883604
R4685 VSS.n4207 DVSS 0.0837012
R4686 VSS.n4324 VSS.n2199 0.08175
R4687 VSS.n4331 VSS.n2201 0.08175
R4688 DVSS VSS.n5419 0.0812353
R4689 DVSS VSS.n5323 0.0812353
R4690 DVSS VSS.n5324 0.0812353
R4691 VSS.n3918 VSS.n3768 0.077375
R4692 VSS.n4145 VSS.n3760 0.077375
R4693 DVSS VSS.n5436 0.0772647
R4694 VSS.n5264 VSS.n2238 0.0769706
R4695 VSS.n5264 VSS.n5263 0.0769706
R4696 VSS.n3541 VSS.n3538 0.0766156
R4697 VSS.n4125 VSS.n4124 0.0763777
R4698 VSS.n5069 DVSS 0.0761
R4699 VSS.n5060 DVSS 0.0761
R4700 VSS.n4981 DVSS 0.0761
R4701 DVSS VSS.n4980 0.0761
R4702 VSS.n4918 DVSS 0.0761
R4703 VSS.n4909 DVSS 0.0761
R4704 VSS.n3186 DVSS 0.0761
R4705 VSS.n3242 DVSS 0.0761
R4706 VSS.n3121 DVSS 0.0761
R4707 DVSS VSS.n2845 0.0761
R4708 DVSS VSS.n2882 0.0761
R4709 VSS.n3003 DVSS 0.0761
R4710 DVSS VSS.n2915 0.0761
R4711 VSS.n2960 DVSS 0.0761
R4712 VSS.n4125 VSS.n3782 0.0756596
R4713 VSS.n4212 DVSS 0.0748392
R4714 VSS.n4210 DVSS 0.0746758
R4715 VSS.n2939 VSS.n2938 0.07437
R4716 VSS.n2065 VSS.n1598 0.0741096
R4717 VSS.n4527 VSS.n2548 0.0728571
R4718 VSS.n4191 VSS.n2638 0.0693638
R4719 VSS.n4201 VSS.n2633 0.0668158
R4720 VSS.n4303 VSS.n4217 0.0656316
R4721 VSS.n5176 DVSS 0.064306
R4722 VSS.n2059 VSS.n1598 0.0624601
R4723 VSS.n4675 VSS.n4674 0.0620789
R4724 VSS.n3542 VSS.n3541 0.0602043
R4725 VSS.n38 VSS.n35 0.0597445
R4726 VSS.n40 VSS.n39 0.0597445
R4727 VSS.n42 VSS.n41 0.0597445
R4728 VSS.n44 VSS.n43 0.0597445
R4729 VSS.n46 VSS.n45 0.0597445
R4730 VSS.n48 VSS.n47 0.0597445
R4731 VSS.n50 VSS.n49 0.0597445
R4732 VSS.n52 VSS.n51 0.0597445
R4733 VSS.n54 VSS.n53 0.0597445
R4734 VSS.n67 VSS.n56 0.0597445
R4735 VSS.n76 VSS.n66 0.0597445
R4736 VSS.n75 VSS.n65 0.0597445
R4737 VSS.n74 VSS.n64 0.0597445
R4738 VSS.n73 VSS.n63 0.0597445
R4739 VSS.n72 VSS.n62 0.0597445
R4740 VSS.n71 VSS.n61 0.0597445
R4741 VSS.n70 VSS.n60 0.0597445
R4742 VSS.n69 VSS.n59 0.0597445
R4743 VSS.n68 VSS.n58 0.0597445
R4744 VSS.n1143 VSS.n35 0.0597445
R4745 VSS.n39 VSS.n38 0.0597445
R4746 VSS.n41 VSS.n40 0.0597445
R4747 VSS.n43 VSS.n42 0.0597445
R4748 VSS.n45 VSS.n44 0.0597445
R4749 VSS.n47 VSS.n46 0.0597445
R4750 VSS.n49 VSS.n48 0.0597445
R4751 VSS.n51 VSS.n50 0.0597445
R4752 VSS.n53 VSS.n52 0.0597445
R4753 VSS.n55 VSS.n54 0.0597445
R4754 VSS.n76 VSS.n67 0.0597445
R4755 VSS.n75 VSS.n66 0.0597445
R4756 VSS.n74 VSS.n65 0.0597445
R4757 VSS.n73 VSS.n64 0.0597445
R4758 VSS.n72 VSS.n63 0.0597445
R4759 VSS.n71 VSS.n62 0.0597445
R4760 VSS.n70 VSS.n61 0.0597445
R4761 VSS.n69 VSS.n60 0.0597445
R4762 VSS.n68 VSS.n59 0.0597445
R4763 VSS.n2077 VSS.n2076 0.0588383
R4764 VSS.n4123 VSS.n3784 0.058625
R4765 VSS.n3881 VSS.n3880 0.058625
R4766 VSS.n4187 VSS.n2638 0.0585457
R4767 VSS.n2550 VSS.n2548 0.058308
R4768 DVSS VSS.n2624 0.0574691
R4769 VSS.n5173 DVSS 0.0569179
R4770 DVSS VSS.n2272 0.0569179
R4771 VSS.n5707 VSS.n16 0.0562784
R4772 VSS.n3883 VSS.n3778 0.0546667
R4773 VSS.n4127 VSS.n3778 0.0546667
R4774 VSS.n4129 VSS.n4128 0.0546667
R4775 VSS.n4128 VSS.n4127 0.0546667
R4776 VSS.n3920 VSS.n3919 0.0544368
R4777 VSS.n3921 VSS.n3920 0.0544368
R4778 VSS.n3878 VSS.n3877 0.0544368
R4779 VSS.n3878 VSS.n3871 0.0544368
R4780 VSS.n3523 VSS 0.0537197
R4781 VSS.n3525 VSS 0.0537197
R4782 VSS.n4171 VSS.n2652 0.0532027
R4783 VSS.n4061 VSS.n4058 0.0532027
R4784 VSS.n5707 VSS.n5706 0.0500653
R4785 VSS.n4328 VSS.n4327 0.0495566
R4786 VSS.n5295 VSS.n5294 0.0495566
R4787 VSS.n4332 VSS.n4331 0.0486793
R4788 VSS.n2513 VSS 0.0456808
R4789 VSS.n4857 VSS 0.0456808
R4790 VSS.n2700 VSS 0.0456808
R4791 VSS.n2699 VSS 0.0456808
R4792 VSS.n3253 VSS 0.0456808
R4793 VSS.n3943 VSS.n3942 0.0450872
R4794 VSS.n3752 VSS.n3750 0.0450872
R4795 VSS.n4101 VSS.n4100 0.0450872
R4796 VSS.n3831 VSS.n3830 0.0450872
R4797 VSS.n3866 VSS.n3839 0.0450872
R4798 VSS.n3721 VSS.n2653 0.0450718
R4799 VSS.n3723 VSS.n3721 0.0450718
R4800 VSS.n3728 VSS.n3727 0.0450718
R4801 VSS.n3729 VSS.n3728 0.0450718
R4802 VSS.n3947 VSS.n3906 0.0450718
R4803 VSS.n3906 VSS.n3904 0.0450718
R4804 VSS.n4080 VSS.n4064 0.0442838
R4805 VSS.n4073 VSS.n4072 0.0442838
R4806 VSS.n4082 VSS.n4081 0.0442838
R4807 VSS.n4081 VSS.n4065 0.0442838
R4808 VSS.n4075 VSS.n4074 0.0442838
R4809 VSS.n3832 VSS.n3824 0.0442838
R4810 VSS.n3833 VSS.n3832 0.0442838
R4811 VSS.n3838 VSS.n3837 0.0442838
R4812 VSS.n4171 VSS.n4170 0.0442838
R4813 VSS.n4168 VSS.n4167 0.0442838
R4814 VSS.n4167 VSS.n3724 0.0442838
R4815 VSS.n3747 VSS.n3746 0.0442838
R4816 VSS.n3748 VSS.n3747 0.0442838
R4817 VSS.n3753 VSS.n3748 0.0442838
R4818 VSS.n3754 VSS.n3753 0.0442838
R4819 VSS.n4150 VSS.n3754 0.0442838
R4820 VSS.n4150 VSS.n4149 0.0442838
R4821 VSS.n4149 VSS.n3755 0.0442838
R4822 VSS.n3926 VSS.n3774 0.0442838
R4823 VSS.n3928 VSS.n3926 0.0442838
R4824 VSS.n3928 VSS.n3927 0.0442838
R4825 VSS.n3927 VSS.n3909 0.0442838
R4826 VSS.n3944 VSS.n3909 0.0442838
R4827 VSS.n3945 VSS.n3944 0.0442838
R4828 VSS.n3945 VSS.n3907 0.0442838
R4829 VSS.n3953 VSS.n3952 0.0442838
R4830 VSS.n4103 VSS.n3953 0.0442838
R4831 VSS.n4103 VSS.n4102 0.0442838
R4832 VSS.n4102 VSS.n3954 0.0442838
R4833 VSS.n4060 VSS.n3954 0.0442838
R4834 VSS.n4061 VSS.n4060 0.0442838
R4835 VSS.n2568 VSS.n2199 0.0432989
R4836 VSS.n3946 VSS.n3908 0.0430229
R4837 VSS.n3749 VSS.n3725 0.0430229
R4838 VSS.n3834 VSS.n3823 0.0426101
R4839 VSS.n4104 VSS.n3903 0.0421972
R4840 VSS.n4163 VSS.n3732 0.0418677
R4841 VSS.n3948 VSS.n3890 0.0418677
R4842 VSS.n4079 VSS.n4078 0.0418514
R4843 VSS.n5708 VSS.n5707 0.0417698
R4844 VSS.n5709 VSS.n5708 0.0417698
R4845 VSS.n2078 VSS.n2077 0.0417698
R4846 VSS.n2079 VSS.n2078 0.0417698
R4847 VSS.n3929 VSS.n3925 0.0405459
R4848 VSS.n4151 VSS.n3745 0.0405459
R4849 VSS.n3244 VSS.n3243 0.0398939
R4850 VSS.n3245 VSS.n3244 0.0398939
R4851 VSS.n4173 VSS.n4172 0.0397202
R4852 VSS.n4075 VSS.n4067 0.0382027
R4853 VSS.n3837 VSS.n3822 0.0382027
R4854 VSS.n4126 VSS.n4125 0.0381812
R4855 VSS.n4127 VSS.n4126 0.0381812
R4856 VSS.n4064 VSS.n3965 0.0373919
R4857 VSS.n4532 VSS.n4531 0.0359178
R4858 VSS.n4330 VSS.n4329 0.0357988
R4859 VSS.n4872 VSS.n4871 0.0349371
R4860 VSS.n4871 VSS.n4870 0.0349371
R4861 VSS.n2517 VSS 0.0348421
R4862 VSS.n4099 VSS.n3955 0.0339404
R4863 VSS.n377 VSS.n372 0.0336863
R4864 VSS.n579 VSS.n373 0.0336863
R4865 VSS.n5429 VSS.n5428 0.0336579
R4866 VSS.n5335 VSS.n2181 0.0336579
R4867 VSS.n5338 VSS.n5337 0.0336579
R4868 VSS.n5432 VSS.n5431 0.0336579
R4869 VSS.n578 VSS.n374 0.0332409
R4870 VSS.n3941 VSS.n3910 0.0331147
R4871 VSS.n3751 VSS.n3744 0.0331147
R4872 VSS.n1877 VSS.n14 0.033
R4873 VSS.n14 VSS.n13 0.033
R4874 VSS.n1746 VSS.n1745 0.033
R4875 VSS.n1745 VSS.n1744 0.033
R4876 VSS.n1728 VSS.n1704 0.033
R4877 VSS.n1743 VSS.n1728 0.033
R4878 VSS.n1741 VSS.n1740 0.033
R4879 VSS.n1742 VSS.n1741 0.033
R4880 VSS.n1735 VSS.n1734 0.033
R4881 VSS.n1735 VSS.n1729 0.033
R4882 VSS.n2042 VSS.n1295 0.033
R4883 VSS.n1295 VSS.n1293 0.033
R4884 VSS.n5424 VSS.n2101 0.0322647
R4885 VSS.n5180 DVSS 0.0320421
R4886 VSS.n3869 VSS.n3819 0.031778
R4887 VSS.n4120 VSS.n4119 0.031778
R4888 VSS.n2949 VSS.n2948 0.0315
R4889 VSS.n2992 VSS.n2903 0.0315
R4890 VSS.n2996 VSS.n2903 0.0315
R4891 VSS.n3047 VSS.n3046 0.0315
R4892 VSS.n3100 VSS.n3099 0.0315
R4893 VSS.n3147 VSS.n2839 0.0315
R4894 VSS.n3188 VSS.n2804 0.0315
R4895 VSS.n4874 VSS.n2396 0.0315
R4896 VSS.n4944 VSS.n4943 0.0315
R4897 VSS.n4983 VSS.n2353 0.0315
R4898 VSS.n5026 VSS.n2322 0.0315
R4899 VSS.n5091 VSS.n2302 0.0315
R4900 VSS.n5092 VSS.n5091 0.0315
R4901 VSS.n5111 VSS.n5110 0.0315
R4902 VSS.n2933 VSS.n2932 0.0315
R4903 VSS.n2961 VSS.n2901 0.0315
R4904 VSS.n3000 VSS.n2901 0.0315
R4905 VSS.n3006 VSS.n3005 0.0315
R4906 VSS.n3067 VSS.n3066 0.0315
R4907 VSS.n3134 VSS.n3133 0.0315
R4908 VSS.n3240 VSS.n2800 0.0315
R4909 VSS.n3211 VSS.n3210 0.0315
R4910 VSS.n4903 VSS.n4902 0.0315
R4911 VSS.n4976 VSS.n4975 0.0315
R4912 VSS.n5011 VSS.n5010 0.0315
R4913 VSS.n5056 VSS.n2304 0.0315
R4914 VSS.n5053 VSS.n2304 0.0315
R4915 VSS.n5124 VSS.n2284 0.0315
R4916 VSS.n3836 VSS.n3821 0.0310505
R4917 VSS.n2947 VSS.n2925 0.031
R4918 VSS.n3050 VSS.n2881 0.031
R4919 VSS.n5027 VSS.n2332 0.031
R4920 VSS.n5171 VSS.n2276 0.031
R4921 VSS.n2936 VSS.n2927 0.031
R4922 VSS.n3054 VSS.n2879 0.031
R4923 VSS.n5013 VSS.n2331 0.031
R4924 VSS.n5125 VSS.n2278 0.031
R4925 VSS.n4074 VSS.n4068 0.0309054
R4926 VSS.n3838 VSS.n3820 0.0309054
R4927 VSS.n387 VSS.n374 0.0309017
R4928 VSS.n4063 VSS.n4062 0.0306376
R4929 VSS.n4076 VSS.n4066 0.0305
R4930 VSS.n3103 VSS.n2859 0.0305
R4931 VSS.n4963 VSS.n4962 0.0305
R4932 VSS.n3063 VSS.n3058 0.0305
R4933 VSS.n4974 VSS.n4973 0.0305
R4934 VSS.n385 VSS.n377 0.0304416
R4935 VSS.n386 VSS.n373 0.0304416
R4936 VSS.n4166 VSS.n4165 0.0302248
R4937 VSS.n3950 VSS.n3902 0.0302248
R4938 VSS.n1144 VSS.n1143 0.0301222
R4939 VSS.n1141 VSS.n55 0.0301222
R4940 VSS.n1140 VSS.n56 0.0301222
R4941 VSS.n1078 VSS.n58 0.0301222
R4942 VSS.n5176 VSS.n5175 0.0300522
R4943 VSS.n3148 VSS.n2829 0.03
R4944 VSS.n4942 VSS.n2376 0.03
R4945 VSS.n3130 VSS.n2838 0.03
R4946 VSS.n4905 VSS.n2378 0.03
R4947 VSS.n4533 VSS.n4532 0.0298971
R4948 VSS.n3237 VSS.n3236 0.0295
R4949 VSS.n4875 VSS.n2406 0.0295
R4950 VSS.n3239 VSS.n2801 0.0295
R4951 VSS.n3213 VSS.n2405 0.0295
R4952 VSS.n3189 VSS.n2818 0.029
R4953 VSS.n4890 VSS.n4889 0.029
R4954 VSS.n3174 VSS.n2817 0.029
R4955 VSS.n2399 VSS.n2398 0.029
R4956 VSS.n3836 VSS.n3835 0.0285734
R4957 VSS.n3143 VSS.n3142 0.0285
R4958 VSS.n4947 VSS.n2374 0.0285
R4959 VSS.n3137 VSS.n2844 0.0285
R4960 VSS.n4901 VSS.n2370 0.0285
R4961 VSS.n184 VSS.n105 0.0283304
R4962 VSS.n185 VSS.n184 0.0283304
R4963 VSS.n186 VSS.n185 0.0283304
R4964 VSS.n186 VSS.n181 0.0283304
R4965 VSS.n190 VSS.n181 0.0283304
R4966 VSS.n191 VSS.n190 0.0283304
R4967 VSS.n192 VSS.n191 0.0283304
R4968 VSS.n192 VSS.n179 0.0283304
R4969 VSS.n196 VSS.n179 0.0283304
R4970 VSS.n197 VSS.n196 0.0283304
R4971 VSS.n198 VSS.n197 0.0283304
R4972 VSS.n198 VSS.n177 0.0283304
R4973 VSS.n202 VSS.n177 0.0283304
R4974 VSS.n203 VSS.n202 0.0283304
R4975 VSS.n204 VSS.n203 0.0283304
R4976 VSS.n204 VSS.n175 0.0283304
R4977 VSS.n208 VSS.n175 0.0283304
R4978 VSS.n209 VSS.n208 0.0283304
R4979 VSS.n210 VSS.n209 0.0283304
R4980 VSS.n210 VSS.n173 0.0283304
R4981 VSS.n214 VSS.n173 0.0283304
R4982 VSS.n215 VSS.n214 0.0283304
R4983 VSS.n914 VSS.n171 0.0283304
R4984 VSS.n233 VSS.n171 0.0283304
R4985 VSS.n234 VSS.n233 0.0283304
R4986 VSS.n234 VSS.n232 0.0283304
R4987 VSS.n238 VSS.n232 0.0283304
R4988 VSS.n239 VSS.n238 0.0283304
R4989 VSS.n240 VSS.n239 0.0283304
R4990 VSS.n240 VSS.n230 0.0283304
R4991 VSS.n244 VSS.n230 0.0283304
R4992 VSS.n245 VSS.n244 0.0283304
R4993 VSS.n246 VSS.n245 0.0283304
R4994 VSS.n246 VSS.n228 0.0283304
R4995 VSS.n250 VSS.n228 0.0283304
R4996 VSS.n251 VSS.n250 0.0283304
R4997 VSS.n252 VSS.n251 0.0283304
R4998 VSS.n252 VSS.n226 0.0283304
R4999 VSS.n256 VSS.n226 0.0283304
R5000 VSS.n257 VSS.n256 0.0283304
R5001 VSS.n258 VSS.n257 0.0283304
R5002 VSS.n258 VSS.n224 0.0283304
R5003 VSS.n262 VSS.n224 0.0283304
R5004 VSS.n904 VSS.n903 0.0283304
R5005 VSS.n4105 VSS.n3902 0.0281606
R5006 VSS.n4077 VSS.n4076 0.0280676
R5007 VSS.n3096 VSS.n2860 0.028
R5008 VSS.n4984 VSS.n2343 0.028
R5009 VSS.n3069 VSS.n3068 0.028
R5010 VSS.n4978 VSS.n2352 0.028
R5011 VSS.n3097 VSS.n2861 0.0279877
R5012 VSS.n3165 VSS.n2828 0.0279877
R5013 VSS.n5025 VSS.n5024 0.0279877
R5014 VSS.n3072 VSS.n3070 0.0279877
R5015 VSS.n3131 VSS.n2824 0.0279877
R5016 VSS.n5014 VSS.n5012 0.0279877
R5017 VSS.n2930 VSS.n2924 0.0279877
R5018 VSS.n2950 VSS.n2924 0.0279877
R5019 VSS.n2952 VSS.n2950 0.0279877
R5020 VSS.n2952 VSS.n2951 0.0279877
R5021 VSS.n2975 VSS.n2974 0.0279877
R5022 VSS.n2975 VSS.n2904 0.0279877
R5023 VSS.n2993 VSS.n2904 0.0279877
R5024 VSS.n2994 VSS.n2993 0.0279877
R5025 VSS.n2995 VSS.n2994 0.0279877
R5026 VSS.n2995 VSS.n2895 0.0279877
R5027 VSS.n3021 VSS.n2895 0.0279877
R5028 VSS.n3022 VSS.n2884 0.0279877
R5029 VSS.n3044 VSS.n2884 0.0279877
R5030 VSS.n3045 VSS.n3044 0.0279877
R5031 VSS.n3049 VSS.n3048 0.0279877
R5032 VSS.n3049 VSS.n2873 0.0279877
R5033 VSS.n3082 VSS.n2873 0.0279877
R5034 VSS.n3083 VSS.n3082 0.0279877
R5035 VSS.n3083 VSS.n2861 0.0279877
R5036 VSS.n3098 VSS.n3097 0.0279877
R5037 VSS.n3102 VSS.n3101 0.0279877
R5038 VSS.n3102 VSS.n2849 0.0279877
R5039 VSS.n3120 VSS.n2849 0.0279877
R5040 VSS.n3122 VSS.n2840 0.0279877
R5041 VSS.n3144 VSS.n2840 0.0279877
R5042 VSS.n3145 VSS.n3144 0.0279877
R5043 VSS.n3146 VSS.n3145 0.0279877
R5044 VSS.n3146 VSS.n2828 0.0279877
R5045 VSS.n3166 VSS.n3165 0.0279877
R5046 VSS.n3184 VSS.n2819 0.0279877
R5047 VSS.n3185 VSS.n3184 0.0279877
R5048 VSS.n3187 VSS.n3185 0.0279877
R5049 VSS.n3235 VSS.n2806 0.0279877
R5050 VSS.n3235 VSS.n3234 0.0279877
R5051 VSS.n3234 VSS.n2807 0.0279877
R5052 VSS.n3222 VSS.n2807 0.0279877
R5053 VSS.n3223 VSS.n3222 0.0279877
R5054 VSS.n3223 VSS.n2407 0.0279877
R5055 VSS.n4891 VSS.n2395 0.0279877
R5056 VSS.n4892 VSS.n4891 0.0279877
R5057 VSS.n4892 VSS.n2386 0.0279877
R5058 VSS.n4917 VSS.n2386 0.0279877
R5059 VSS.n4920 VSS.n4919 0.0279877
R5060 VSS.n4919 VSS.n2375 0.0279877
R5061 VSS.n4945 VSS.n2375 0.0279877
R5062 VSS.n4946 VSS.n4945 0.0279877
R5063 VSS.n4946 VSS.n2365 0.0279877
R5064 VSS.n4960 VSS.n2365 0.0279877
R5065 VSS.n4965 VSS.n4961 0.0279877
R5066 VSS.n4965 VSS.n4964 0.0279877
R5067 VSS.n4964 VSS.n2354 0.0279877
R5068 VSS.n4982 VSS.n2354 0.0279877
R5069 VSS.n5000 VSS.n2342 0.0279877
R5070 VSS.n5001 VSS.n5000 0.0279877
R5071 VSS.n5001 VSS.n2333 0.0279877
R5072 VSS.n5023 VSS.n2333 0.0279877
R5073 VSS.n5024 VSS.n5023 0.0279877
R5074 VSS.n5043 VSS.n2321 0.0279877
R5075 VSS.n5044 VSS.n5043 0.0279877
R5076 VSS.n5044 VSS.n2312 0.0279877
R5077 VSS.n5068 VSS.n2312 0.0279877
R5078 VSS.n5071 VSS.n5070 0.0279877
R5079 VSS.n5070 VSS.n2301 0.0279877
R5080 VSS.n5093 VSS.n2301 0.0279877
R5081 VSS.n5094 VSS.n5093 0.0279877
R5082 VSS.n5094 VSS.n2291 0.0279877
R5083 VSS.n5108 VSS.n2291 0.0279877
R5084 VSS.n5113 VSS.n5109 0.0279877
R5085 VSS.n5113 VSS.n5112 0.0279877
R5086 VSS.n5112 VSS.n2275 0.0279877
R5087 VSS.n5172 VSS.n2275 0.0279877
R5088 VSS.n2935 VSS.n2934 0.0279877
R5089 VSS.n2934 VSS.n2920 0.0279877
R5090 VSS.n2958 VSS.n2920 0.0279877
R5091 VSS.n2959 VSS.n2958 0.0279877
R5092 VSS.n2967 VSS.n2966 0.0279877
R5093 VSS.n2966 VSS.n2964 0.0279877
R5094 VSS.n2964 VSS.n2962 0.0279877
R5095 VSS.n2962 VSS.n2900 0.0279877
R5096 VSS.n3001 VSS.n2900 0.0279877
R5097 VSS.n3002 VSS.n3001 0.0279877
R5098 VSS.n3014 VSS.n3002 0.0279877
R5099 VSS.n3013 VSS.n3011 0.0279877
R5100 VSS.n3011 VSS.n3009 0.0279877
R5101 VSS.n3009 VSS.n3004 0.0279877
R5102 VSS.n3055 VSS.n2878 0.0279877
R5103 VSS.n3056 VSS.n3055 0.0279877
R5104 VSS.n3075 VSS.n3056 0.0279877
R5105 VSS.n3075 VSS.n3074 0.0279877
R5106 VSS.n3074 VSS.n3072 0.0279877
R5107 VSS.n3070 VSS.n3057 0.0279877
R5108 VSS.n3065 VSS.n3064 0.0279877
R5109 VSS.n3064 VSS.n3062 0.0279877
R5110 VSS.n3062 VSS.n3060 0.0279877
R5111 VSS.n3129 VSS.n3128 0.0279877
R5112 VSS.n3136 VSS.n3129 0.0279877
R5113 VSS.n3136 VSS.n3135 0.0279877
R5114 VSS.n3135 VSS.n3132 0.0279877
R5115 VSS.n3132 VSS.n3131 0.0279877
R5116 VSS.n3172 VSS.n2824 0.0279877
R5117 VSS.n3176 VSS.n3173 0.0279877
R5118 VSS.n3176 VSS.n3175 0.0279877
R5119 VSS.n3175 VSS.n2798 0.0279877
R5120 VSS.n3241 VSS.n2799 0.0279877
R5121 VSS.n3204 VSS.n2799 0.0279877
R5122 VSS.n3207 VSS.n3204 0.0279877
R5123 VSS.n3208 VSS.n3207 0.0279877
R5124 VSS.n3215 VSS.n3208 0.0279877
R5125 VSS.n3215 VSS.n3214 0.0279877
R5126 VSS.n3214 VSS.n3212 0.0279877
R5127 VSS.n3209 VSS.n2391 0.0279877
R5128 VSS.n4898 VSS.n2391 0.0279877
R5129 VSS.n4899 VSS.n4898 0.0279877
R5130 VSS.n4910 VSS.n4899 0.0279877
R5131 VSS.n4908 VSS.n4906 0.0279877
R5132 VSS.n4906 VSS.n4904 0.0279877
R5133 VSS.n4904 VSS.n4900 0.0279877
R5134 VSS.n4900 VSS.n2369 0.0279877
R5135 VSS.n4953 VSS.n2369 0.0279877
R5136 VSS.n4954 VSS.n4953 0.0279877
R5137 VSS.n4971 VSS.n2357 0.0279877
R5138 VSS.n4972 VSS.n4971 0.0279877
R5139 VSS.n4972 VSS.n2355 0.0279877
R5140 VSS.n4977 VSS.n2355 0.0279877
R5141 VSS.n4979 VSS.n2338 0.0279877
R5142 VSS.n5007 VSS.n2338 0.0279877
R5143 VSS.n5008 VSS.n5007 0.0279877
R5144 VSS.n5015 VSS.n5008 0.0279877
R5145 VSS.n5015 VSS.n5014 0.0279877
R5146 VSS.n5009 VSS.n2317 0.0279877
R5147 VSS.n5050 VSS.n2317 0.0279877
R5148 VSS.n5051 VSS.n5050 0.0279877
R5149 VSS.n5061 VSS.n5051 0.0279877
R5150 VSS.n5059 VSS.n5057 0.0279877
R5151 VSS.n5057 VSS.n5055 0.0279877
R5152 VSS.n5055 VSS.n5054 0.0279877
R5153 VSS.n5054 VSS.n2295 0.0279877
R5154 VSS.n5101 VSS.n2295 0.0279877
R5155 VSS.n5102 VSS.n5101 0.0279877
R5156 VSS.n5120 VSS.n2285 0.0279877
R5157 VSS.n5121 VSS.n5120 0.0279877
R5158 VSS.n5123 VSS.n5121 0.0279877
R5159 VSS.n5123 VSS.n5122 0.0279877
R5160 VSS.n4920 VSS.n4918 0.0275443
R5161 VSS.n4909 VSS.n4908 0.0275443
R5162 VSS.n2953 VSS.n2923 0.0275
R5163 VSS.n3043 VSS.n2883 0.0275
R5164 VSS.n5042 VSS.n5041 0.0275
R5165 VSS.n5114 VSS.n2290 0.0275
R5166 VSS.n2957 VSS.n2921 0.0275
R5167 VSS.n3008 VSS.n3007 0.0275
R5168 VSS.n2325 VSS.n2324 0.0275
R5169 VSS.n5119 VSS.n5118 0.0275
R5170 VSS.n3921 VSS.n3784 0.0274684
R5171 VSS.n3919 VSS.n3918 0.0274684
R5172 VSS.n3880 VSS.n3871 0.0274684
R5173 VSS.n3877 VSS.n3760 0.0274684
R5174 VSS.n904 VSS.n222 0.0272082
R5175 VSS.n2991 VSS.n2905 0.027
R5176 VSS.n2997 VSS.n2896 0.027
R5177 VSS.n5073 VSS.n5072 0.027
R5178 VSS.n5095 VSS.n2300 0.027
R5179 VSS.n2963 VSS.n2907 0.027
R5180 VSS.n2999 VSS.n2898 0.027
R5181 VSS.n5058 VSS.n2310 0.027
R5182 VSS.n5052 VSS.n2296 0.027
R5183 VSS.n3858 VSS.n3855 0.026913
R5184 VSS.n3855 VSS.n3854 0.026913
R5185 VSS.n3854 VSS.n3852 0.026913
R5186 VSS.n3852 VSS.n3850 0.026913
R5187 VSS.n3850 VSS.n3848 0.026913
R5188 VSS.n3848 VSS.n3845 0.026913
R5189 VSS.n3845 VSS.n3844 0.026913
R5190 VSS.n3844 VSS.n3842 0.026913
R5191 VSS.n3842 VSS.n2568 0.026913
R5192 VSS.n4346 VSS.n4330 0.026913
R5193 VSS.n4346 VSS.n4345 0.026913
R5194 VSS.n4345 VSS.n4343 0.026913
R5195 VSS.n4343 VSS.n4340 0.026913
R5196 VSS.n4340 VSS.n4339 0.026913
R5197 VSS.n4339 VSS.n4337 0.026913
R5198 VSS.n4337 VSS.n4335 0.026913
R5199 VSS.n4335 VSS.n4332 0.026913
R5200 VSS.n2615 VSS.n2613 0.026913
R5201 VSS.n4342 VSS.n4341 0.026913
R5202 VSS.n4334 VSS.n4333 0.026913
R5203 VSS.n4525 VSS.n2548 0.0267204
R5204 VSS.n4189 VSS.n2638 0.0267108
R5205 VSS.n3930 VSS.n3910 0.0265092
R5206 VSS.n4152 VSS.n3744 0.0265092
R5207 VSS.n3051 VSS.n2874 0.0265
R5208 VSS.n5022 VSS.n5021 0.0265
R5209 VSS.n3053 VSS.n2876 0.0265
R5210 VSS.n5016 VSS.n2337 0.0265
R5211 VSS.n4872 VSS.n2407 0.0262143
R5212 VSS.n4853 VSS.n4852 0.02615
R5213 VSS.n3104 VSS.n2850 0.026
R5214 VSS.n4966 VSS.n2364 0.026
R5215 VSS.n3061 VSS.n2858 0.026
R5216 VSS.n4970 VSS.n2356 0.026
R5217 VSS.n3541 VSS.n3540 0.0258812
R5218 VSS.n3187 VSS.n3186 0.0257709
R5219 VSS.n570 VSS.n524 0.0257489
R5220 VSS.n566 VSS.n524 0.0257489
R5221 VSS.n566 VSS.n565 0.0257489
R5222 VSS.n565 VSS.n564 0.0257489
R5223 VSS.n564 VSS.n526 0.0257489
R5224 VSS.n560 VSS.n526 0.0257489
R5225 VSS.n560 VSS.n559 0.0257489
R5226 VSS.n559 VSS.n558 0.0257489
R5227 VSS.n558 VSS.n528 0.0257489
R5228 VSS.n554 VSS.n528 0.0257489
R5229 VSS.n554 VSS.n553 0.0257489
R5230 VSS.n553 VSS.n552 0.0257489
R5231 VSS.n552 VSS.n530 0.0257489
R5232 VSS.n548 VSS.n530 0.0257489
R5233 VSS.n548 VSS.n547 0.0257489
R5234 VSS.n547 VSS.n546 0.0257489
R5235 VSS.n546 VSS.n532 0.0257489
R5236 VSS.n542 VSS.n532 0.0257489
R5237 VSS.n542 VSS.n541 0.0257489
R5238 VSS.n541 VSS.n540 0.0257489
R5239 VSS.n540 VSS.n534 0.0257489
R5240 VSS.n536 VSS.n534 0.0257489
R5241 VSS.n632 VSS.n364 0.0257489
R5242 VSS.n637 VSS.n364 0.0257489
R5243 VSS.n638 VSS.n637 0.0257489
R5244 VSS.n639 VSS.n638 0.0257489
R5245 VSS.n639 VSS.n362 0.0257489
R5246 VSS.n643 VSS.n362 0.0257489
R5247 VSS.n644 VSS.n643 0.0257489
R5248 VSS.n645 VSS.n644 0.0257489
R5249 VSS.n645 VSS.n360 0.0257489
R5250 VSS.n649 VSS.n360 0.0257489
R5251 VSS.n650 VSS.n649 0.0257489
R5252 VSS.n651 VSS.n650 0.0257489
R5253 VSS.n651 VSS.n358 0.0257489
R5254 VSS.n655 VSS.n358 0.0257489
R5255 VSS.n656 VSS.n655 0.0257489
R5256 VSS.n657 VSS.n656 0.0257489
R5257 VSS.n657 VSS.n356 0.0257489
R5258 VSS.n661 VSS.n356 0.0257489
R5259 VSS.n662 VSS.n661 0.0257489
R5260 VSS.n663 VSS.n662 0.0257489
R5261 VSS.n663 VSS.n353 0.0257489
R5262 VSS.n668 VSS.n354 0.0257489
R5263 VSS.n4059 VSS.n3955 0.0256835
R5264 VSS.n3022 DVSS 0.0255493
R5265 DVSS VSS.n3013 0.0255493
R5266 VSS.n3164 VSS.n3163 0.0255
R5267 VSS.n4922 VSS.n4921 0.0255
R5268 VSS.n2832 VSS.n2831 0.0255
R5269 VSS.n4907 VSS.n2384 0.0255
R5270 VSS.n3233 VSS.n2805 0.025
R5271 VSS.n3224 VSS.n3221 0.025
R5272 VSS.n3203 VSS.n3202 0.025
R5273 VSS.n3216 VSS.n3200 0.025
R5274 VSS.n903 VSS.n902 0.0249638
R5275 VSS.n4981 VSS.n2342 0.0248842
R5276 VSS.n4980 VSS.n4979 0.0248842
R5277 VSS.n1613 VSS.n1598 0.0248508
R5278 VSS.n2938 VSS.n2929 0.0248045
R5279 VSS.n380 VSS.n354 0.0247308
R5280 VSS.n3183 VSS.n3182 0.0245
R5281 VSS.n4893 VSS.n2394 0.0245
R5282 VSS.n3177 VSS.n2823 0.0245
R5283 VSS.n4897 VSS.n2392 0.0245
R5284 VSS.n5324 VSS.n5319 0.0242837
R5285 VSS.n5323 VSS.n5320 0.0242837
R5286 VSS.n2706 DVSS 0.0241842
R5287 VSS.n3141 VSS.n2841 0.024
R5288 VSS.n4949 VSS.n4948 0.024
R5289 VSS.n3138 VSS.n2843 0.024
R5290 VSS.n4952 VSS.n4951 0.024
R5291 VSS.n3095 VSS.n2862 0.0235
R5292 VSS.n4999 VSS.n4998 0.0235
R5293 VSS.n3071 VSS.n2864 0.0235
R5294 VSS.n2346 VSS.n2345 0.0235
R5295 VSS.n3121 VSS.n3120 0.0231108
R5296 VSS.n3060 VSS.n2845 0.0231108
R5297 VSS.n2954 VSS.n2916 0.023
R5298 VSS.n3042 VSS.n2885 0.023
R5299 VSS.n5045 VSS.n2320 0.023
R5300 VSS.n5115 VSS.n2289 0.023
R5301 VSS.n2956 VSS.n2918 0.023
R5302 VSS.n3010 VSS.n2887 0.023
R5303 VSS.n5049 VSS.n2318 0.023
R5304 VSS.n5117 VSS.n2286 0.023
R5305 VSS.n3101 DVSS 0.0228892
R5306 VSS.n3065 DVSS 0.0228892
R5307 VSS.n3829 VSS.n2650 0.0227936
R5308 VSS.n4168 VSS.n3723 0.0227859
R5309 VSS.n3746 VSS.n3729 0.0227859
R5310 VSS.n3757 VSS.n3755 0.0227859
R5311 VSS.n4130 VSS.n3772 0.0227859
R5312 VSS.n3952 VSS.n3904 0.0227859
R5313 VSS.n3758 VSS.n3757 0.0227859
R5314 VSS.n3774 VSS.n3772 0.0227859
R5315 VSS.n3947 VSS.n3907 0.0227859
R5316 VSS.n3727 VSS.n3724 0.0227859
R5317 VSS.n4170 VSS.n2653 0.0227859
R5318 VSS.n4344 VSS.n2610 0.0227554
R5319 VSS.n4338 VSS.n2607 0.0227554
R5320 VSS.n669 VSS.n668 0.0226946
R5321 VSS.n2977 VSS.n2976 0.0225
R5322 VSS.n3020 VSS.n3019 0.0225
R5323 VSS.n5067 VSS.n2311 0.0225
R5324 VSS.n5097 VSS.n5096 0.0225
R5325 VSS.n2965 VSS.n2913 0.0225
R5326 VSS.n3016 VSS.n3015 0.0225
R5327 VSS.n5062 VSS.n2316 0.0225
R5328 VSS.n5100 VSS.n5099 0.0225
R5329 VSS.n4086 VSS.n4063 0.0223919
R5330 VSS.n4084 VSS.n4063 0.0223919
R5331 VSS.n3825 VSS.n2652 0.0223919
R5332 VSS.n4083 VSS.n4058 0.0223919
R5333 VSS.n4085 VSS.n4083 0.0223919
R5334 VSS.n3829 VSS.n3828 0.0223807
R5335 VSS.n3830 VSS.n3829 0.0223807
R5336 VSS.n5071 VSS.n5069 0.0222241
R5337 VSS.n5060 VSS.n5059 0.0222241
R5338 VSS.n3081 VSS.n3080 0.022
R5339 VSS.n5020 VSS.n2334 0.022
R5340 VSS.n3077 VSS.n3076 0.022
R5341 VSS.n5017 VSS.n2336 0.022
R5342 VSS.n5419 VSS.n5418 0.0216765
R5343 VSS.n4132 VSS.n3773 0.021555
R5344 VSS.n4166 VSS.n3722 0.021555
R5345 VSS.n906 VSS.n905 0.0215113
R5346 VSS.n3119 VSS.n3118 0.0215
R5347 VSS.n4967 VSS.n2361 0.0215
R5348 VSS.n3059 VSS.n2852 0.0215
R5349 VSS.n4969 VSS.n2358 0.0215
R5350 VSS.n4438 VSS.n4347 0.021288
R5351 VSS.n4336 VSS.n2606 0.021288
R5352 VSS.n5452 VSS.n1287 0.021205
R5353 VSS.n5459 VSS.n1287 0.021205
R5354 VSS.n5460 VSS.n5459 0.021205
R5355 VSS.n5461 VSS.n5460 0.021205
R5356 VSS.n5461 VSS.n1283 0.021205
R5357 VSS.n5467 VSS.n1283 0.021205
R5358 VSS.n5468 VSS.n5467 0.021205
R5359 VSS.n5469 VSS.n5468 0.021205
R5360 VSS.n5469 VSS.n1279 0.021205
R5361 VSS.n5475 VSS.n1279 0.021205
R5362 VSS.n5476 VSS.n5475 0.021205
R5363 VSS.n5477 VSS.n5476 0.021205
R5364 VSS.n5477 VSS.n1275 0.021205
R5365 VSS.n5483 VSS.n1275 0.021205
R5366 VSS.n5484 VSS.n5483 0.021205
R5367 VSS.n5485 VSS.n5484 0.021205
R5368 VSS.n5485 VSS.n1271 0.021205
R5369 VSS.n5491 VSS.n1271 0.021205
R5370 VSS.n5492 VSS.n5491 0.021205
R5371 VSS.n5493 VSS.n5492 0.021205
R5372 VSS.n5493 VSS.n1267 0.021205
R5373 VSS.n5499 VSS.n1267 0.021205
R5374 VSS.n5500 VSS.n5499 0.021205
R5375 VSS.n5501 VSS.n5500 0.021205
R5376 VSS.n5501 VSS.n1263 0.021205
R5377 VSS.n5507 VSS.n1263 0.021205
R5378 VSS.n5508 VSS.n5507 0.021205
R5379 VSS.n5509 VSS.n5508 0.021205
R5380 VSS.n5509 VSS.n1259 0.021205
R5381 VSS.n5515 VSS.n1259 0.021205
R5382 VSS.n5516 VSS.n5515 0.021205
R5383 VSS.n5517 VSS.n5516 0.021205
R5384 VSS.n5517 VSS.n1255 0.021205
R5385 VSS.n5523 VSS.n1255 0.021205
R5386 VSS.n5524 VSS.n5523 0.021205
R5387 VSS.n5525 VSS.n5524 0.021205
R5388 VSS.n5525 VSS.n1251 0.021205
R5389 VSS.n5531 VSS.n1251 0.021205
R5390 VSS.n5532 VSS.n5531 0.021205
R5391 VSS.n5533 VSS.n5532 0.021205
R5392 VSS.n5533 VSS.n1247 0.021205
R5393 VSS.n5539 VSS.n1247 0.021205
R5394 VSS.n5540 VSS.n5539 0.021205
R5395 VSS.n5541 VSS.n5540 0.021205
R5396 VSS.n5541 VSS.n1243 0.021205
R5397 VSS.n5547 VSS.n1243 0.021205
R5398 VSS.n5548 VSS.n5547 0.021205
R5399 VSS.n5549 VSS.n5548 0.021205
R5400 VSS.n5549 VSS.n1239 0.021205
R5401 VSS.n5555 VSS.n1239 0.021205
R5402 VSS.n5556 VSS.n5555 0.021205
R5403 VSS.n5557 VSS.n5556 0.021205
R5404 VSS.n5557 VSS.n1235 0.021205
R5405 VSS.n5563 VSS.n1235 0.021205
R5406 VSS.n5564 VSS.n5563 0.021205
R5407 VSS.n5566 VSS.n5564 0.021205
R5408 VSS.n5566 VSS.n5565 0.021205
R5409 VSS.n5574 VSS.n5573 0.021205
R5410 VSS.n5575 VSS.n5574 0.021205
R5411 VSS.n5575 VSS.n1227 0.021205
R5412 VSS.n5581 VSS.n1227 0.021205
R5413 VSS.n5582 VSS.n5581 0.021205
R5414 VSS.n5583 VSS.n5582 0.021205
R5415 VSS.n5583 VSS.n1223 0.021205
R5416 VSS.n5589 VSS.n1223 0.021205
R5417 VSS.n5590 VSS.n5589 0.021205
R5418 VSS.n5591 VSS.n5590 0.021205
R5419 VSS.n5591 VSS.n1219 0.021205
R5420 VSS.n5597 VSS.n1219 0.021205
R5421 VSS.n5598 VSS.n5597 0.021205
R5422 VSS.n5599 VSS.n5598 0.021205
R5423 VSS.n5599 VSS.n1215 0.021205
R5424 VSS.n5605 VSS.n1215 0.021205
R5425 VSS.n5606 VSS.n5605 0.021205
R5426 VSS.n5607 VSS.n5606 0.021205
R5427 VSS.n5607 VSS.n1211 0.021205
R5428 VSS.n5613 VSS.n1211 0.021205
R5429 VSS.n5614 VSS.n5613 0.021205
R5430 VSS.n5615 VSS.n5614 0.021205
R5431 VSS.n5615 VSS.n1207 0.021205
R5432 VSS.n5621 VSS.n1207 0.021205
R5433 VSS.n5622 VSS.n5621 0.021205
R5434 VSS.n5623 VSS.n5622 0.021205
R5435 VSS.n5623 VSS.n1203 0.021205
R5436 VSS.n5629 VSS.n1203 0.021205
R5437 VSS.n5630 VSS.n5629 0.021205
R5438 VSS.n5631 VSS.n5630 0.021205
R5439 VSS.n5631 VSS.n1199 0.021205
R5440 VSS.n5637 VSS.n1199 0.021205
R5441 VSS.n5638 VSS.n5637 0.021205
R5442 VSS.n5639 VSS.n5638 0.021205
R5443 VSS.n5639 VSS.n1195 0.021205
R5444 VSS.n5645 VSS.n1195 0.021205
R5445 VSS.n5646 VSS.n5645 0.021205
R5446 VSS.n5647 VSS.n5646 0.021205
R5447 VSS.n5647 VSS.n1191 0.021205
R5448 VSS.n5653 VSS.n1191 0.021205
R5449 VSS.n5654 VSS.n5653 0.021205
R5450 VSS.n5655 VSS.n5654 0.021205
R5451 VSS.n5655 VSS.n1187 0.021205
R5452 VSS.n5661 VSS.n1187 0.021205
R5453 VSS.n5662 VSS.n5661 0.021205
R5454 VSS.n5663 VSS.n5662 0.021205
R5455 VSS.n5663 VSS.n1183 0.021205
R5456 VSS.n5669 VSS.n1183 0.021205
R5457 VSS.n5670 VSS.n5669 0.021205
R5458 VSS.n5671 VSS.n5670 0.021205
R5459 VSS.n5671 VSS.n1179 0.021205
R5460 VSS.n5677 VSS.n1179 0.021205
R5461 VSS.n5678 VSS.n5677 0.021205
R5462 VSS.n5679 VSS.n5678 0.021205
R5463 VSS.n5679 VSS.n1175 0.021205
R5464 VSS.n5685 VSS.n1175 0.021205
R5465 VSS.n5686 VSS.n5685 0.021205
R5466 VSS.n5687 VSS.n5686 0.021205
R5467 VSS.n4083 VSS.n4082 0.0211757
R5468 VSS.n3825 VSS.n3824 0.0211757
R5469 VSS.n4148 VSS.n4147 0.0211422
R5470 VSS.n3167 VSS.n2827 0.021
R5471 VSS.n4916 VSS.n2385 0.021
R5472 VSS.n3171 VSS.n2825 0.021
R5473 VSS.n4911 VSS.n2390 0.021
R5474 VSS.n4133 VSS.n4132 0.02075
R5475 VSS.n4132 VSS.n4131 0.02075
R5476 VSS.n4147 VSS.n3756 0.02075
R5477 VSS.n4147 VSS.n4146 0.02075
R5478 VSS.n3243 VSS.n2798 0.0206724
R5479 VSS.n666 VSS.n221 0.0206158
R5480 VSS.n3232 VSS.n2808 0.0205
R5481 VSS.n3225 VSS.n3220 0.0205
R5482 VSS.n3206 VSS.n2810 0.0205
R5483 VSS.n3217 VSS.n3199 0.0205
R5484 VSS.n3045 VSS.n2882 0.0204507
R5485 VSS.n3004 VSS.n3003 0.0204507
R5486 DVSS VSS.n2819 0.0202291
R5487 VSS.n3173 DVSS 0.0202291
R5488 VSS.n911 VSS.n910 0.020197
R5489 VSS.n3181 VSS.n2820 0.02
R5490 VSS.n4894 VSS.n2387 0.02
R5491 VSS.n3178 VSS.n2822 0.02
R5492 VSS.n4896 VSS.n2389 0.02
R5493 VSS.n4062 VSS.n4059 0.0199037
R5494 VSS.n4172 VSS.n2651 0.0199037
R5495 VSS.n5700 VSS.n5699 0.0195912
R5496 VSS.n5699 VSS.n5698 0.0195912
R5497 VSS.n5698 VSS.n5697 0.0195912
R5498 VSS.n1149 VSS.n1148 0.0195912
R5499 VSS.n1148 VSS.n1147 0.0195912
R5500 VSS.n1147 VSS.n1146 0.0195912
R5501 VSS.n3124 VSS.n3123 0.0195
R5502 VSS.n4959 VSS.n2366 0.0195
R5503 VSS.n3127 VSS.n3126 0.0195
R5504 VSS.n4955 VSS.n2368 0.0195
R5505 VSS.n216 VSS.n215 0.0191284
R5506 VSS.n3930 VSS.n3929 0.019078
R5507 VSS.n4152 VSS.n4151 0.019078
R5508 VSS.n3085 VSS.n3084 0.019
R5509 VSS.n5002 VSS.n2341 0.019
R5510 VSS.n3073 VSS.n2871 0.019
R5511 VSS.n5006 VSS.n2339 0.019
R5512 DVSS VSS.n5108 0.018899
R5513 VSS.n5102 DVSS 0.018899
R5514 VSS.n2973 VSS.n2972 0.0185
R5515 VSS.n3024 VSS.n3023 0.0185
R5516 VSS.n5046 VSS.n2313 0.0185
R5517 VSS.n5107 VSS.n5106 0.0185
R5518 VSS.n2969 VSS.n2968 0.0185
R5519 VSS.n3012 VSS.n2893 0.0185
R5520 VSS.n5048 VSS.n2315 0.0185
R5521 VSS.n5104 VSS.n5103 0.0185
R5522 VSS.n1397 VSS.n1395 0.018166
R5523 VSS.n2973 VSS.n2914 0.018
R5524 VSS.n3023 VSS.n2894 0.018
R5525 VSS.n5066 VSS.n2313 0.018
R5526 VSS.n5107 VSS.n2292 0.018
R5527 VSS.n2968 VSS.n2919 0.018
R5528 VSS.n3012 VSS.n2899 0.018
R5529 VSS.n5063 VSS.n2315 0.018
R5530 VSS.n5103 VSS.n2294 0.018
R5531 VSS.n3722 VSS.n2651 0.0178394
R5532 VSS.n2951 VSS.n2915 0.0177906
R5533 VSS.n2960 VSS.n2959 0.0177906
R5534 VSS.n2074 VSS.n2066 0.0176
R5535 VSS.n1820 VSS.n1819 0.0176
R5536 DVSS VSS.n2395 0.017569
R5537 VSS.n3209 DVSS 0.017569
R5538 VSS.n3084 VSS.n2872 0.0175
R5539 VSS.n5003 VSS.n5002 0.0175
R5540 VSS.n3073 VSS.n2877 0.0175
R5541 VSS.n5006 VSS.n5005 0.0175
R5542 VSS.n4105 VSS.n4104 0.0174266
R5543 VSS.n536 VSS.n535 0.0174005
R5544 VSS.n1818 VSS.n1811 0.0172066
R5545 VSS.n2764 VSS.n9 0.0171667
R5546 VSS.n4869 VSS.n9 0.0171667
R5547 VSS.n1231 VSS.n10 0.0171667
R5548 VSS.n5570 VSS.n10 0.0171667
R5549 VSS.n3835 VSS.n3834 0.0170138
R5550 VSS.n3123 VSS.n2848 0.017
R5551 VSS.n4959 VSS.n4958 0.017
R5552 VSS.n3127 VSS.n2846 0.017
R5553 VSS.n4956 VSS.n4955 0.017
R5554 VSS.n2424 VSS.n2415 0.0169185
R5555 VSS.n2424 VSS.n2423 0.0169185
R5556 VSS.n3369 VSS.n2426 0.0169185
R5557 VSS.n2426 VSS.n2425 0.0169185
R5558 VSS.n3370 VSS.n2428 0.0169185
R5559 VSS.n2428 VSS.n2427 0.0169185
R5560 VSS.n3371 VSS.n2430 0.0169185
R5561 VSS.n2430 VSS.n2429 0.0169185
R5562 VSS.n4854 VSS.n2431 0.0169185
R5563 VSS.n4841 VSS.n4840 0.0169185
R5564 VSS.n4839 VSS.n4838 0.0169185
R5565 VSS.n4837 VSS.n4836 0.0169185
R5566 VSS.n4836 VSS.n4835 0.0169185
R5567 VSS.n4834 VSS.n4833 0.0169185
R5568 VSS.n4831 VSS.n4830 0.0169185
R5569 VSS.n4830 VSS.n4829 0.0169185
R5570 VSS.n4827 VSS.n4826 0.0169185
R5571 VSS.n1602 VSS.n1596 0.0169185
R5572 VSS.n1604 VSS.n1602 0.0169185
R5573 VSS.n1612 VSS.n1601 0.0169185
R5574 VSS.n1606 VSS.n1601 0.0169185
R5575 VSS.n1611 VSS.n1600 0.0169185
R5576 VSS.n1608 VSS.n1600 0.0169185
R5577 VSS.n1610 VSS.n1599 0.0169185
R5578 VSS.n2063 VSS.n1599 0.0169185
R5579 VSS.n2066 VSS.n1596 0.0169185
R5580 VSS.n1605 VSS.n1604 0.0169185
R5581 VSS.n1612 VSS.n1605 0.0169185
R5582 VSS.n1607 VSS.n1606 0.0169185
R5583 VSS.n1611 VSS.n1607 0.0169185
R5584 VSS.n1609 VSS.n1608 0.0169185
R5585 VSS.n1610 VSS.n1609 0.0169185
R5586 VSS.n2064 VSS.n2063 0.0169185
R5587 VSS.n1807 VSS.n1796 0.0169185
R5588 VSS.n1808 VSS.n1806 0.0169185
R5589 VSS.n1804 VSS.n1795 0.0169185
R5590 VSS.n1805 VSS.n1803 0.0169185
R5591 VSS.n1801 VSS.n1794 0.0169185
R5592 VSS.n1802 VSS.n1800 0.0169185
R5593 VSS.n1799 VSS.n1793 0.0169185
R5594 VSS.n1856 VSS.n1855 0.0169185
R5595 VSS.n1820 VSS.n1796 0.0169185
R5596 VSS.n1808 VSS.n1807 0.0169185
R5597 VSS.n1806 VSS.n1795 0.0169185
R5598 VSS.n1805 VSS.n1804 0.0169185
R5599 VSS.n1803 VSS.n1794 0.0169185
R5600 VSS.n1802 VSS.n1801 0.0169185
R5601 VSS.n1800 VSS.n1793 0.0169185
R5602 VSS.n1855 VSS.n1799 0.0169185
R5603 VSS.n3717 VSS.n3716 0.0169185
R5604 VSS.n2669 VSS.n2668 0.0169185
R5605 VSS.n2671 VSS.n2669 0.0169185
R5606 VSS.n2667 VSS.n2666 0.0169185
R5607 VSS.n2672 VSS.n2667 0.0169185
R5608 VSS.n2665 VSS.n2664 0.0169185
R5609 VSS.n2673 VSS.n2665 0.0169185
R5610 VSS.n2663 VSS.n2662 0.0169185
R5611 VSS.n2663 VSS.n2655 0.0169185
R5612 VSS.n3719 VSS.n2655 0.0169185
R5613 VSS.n2673 VSS.n2660 0.0169185
R5614 VSS.n2662 VSS.n2660 0.0169185
R5615 VSS.n2672 VSS.n2659 0.0169185
R5616 VSS.n2664 VSS.n2659 0.0169185
R5617 VSS.n2671 VSS.n2658 0.0169185
R5618 VSS.n2666 VSS.n2658 0.0169185
R5619 VSS.n3716 VSS.n2657 0.0169185
R5620 VSS.n2668 VSS.n2657 0.0169185
R5621 VSS.n4856 VSS.n2415 0.0169185
R5622 VSS.n2423 VSS.n2421 0.0169185
R5623 VSS.n3369 VSS.n2421 0.0169185
R5624 VSS.n2425 VSS.n2420 0.0169185
R5625 VSS.n3370 VSS.n2420 0.0169185
R5626 VSS.n2427 VSS.n2419 0.0169185
R5627 VSS.n3371 VSS.n2419 0.0169185
R5628 VSS.n2429 VSS.n2418 0.0169185
R5629 VSS.n2431 VSS.n2418 0.0169185
R5630 VSS.n4842 VSS.n4841 0.0169185
R5631 VSS.n4840 VSS.n4839 0.0169185
R5632 VSS.n4838 VSS.n4837 0.0169185
R5633 VSS.n4835 VSS.n4834 0.0169185
R5634 VSS.n4833 VSS.n4832 0.0169185
R5635 VSS.n4832 VSS.n4831 0.0169185
R5636 VSS.n4829 VSS.n4828 0.0169185
R5637 VSS.n4828 VSS.n4827 0.0169185
R5638 VSS.n4078 VSS.n4077 0.0167162
R5639 VSS.n908 VSS.n907 0.0166994
R5640 VSS.n909 VSS.n908 0.0166994
R5641 VSS.n3168 VSS.n2820 0.0165
R5642 VSS.n4915 VSS.n2387 0.0165
R5643 VSS.n3170 VSS.n2822 0.0165
R5644 VSS.n4912 VSS.n2389 0.0165
R5645 VSS.n5173 VSS.n5172 0.0164606
R5646 VSS.n5122 VSS.n2272 0.0164606
R5647 VSS.n5025 DVSS 0.0162389
R5648 VSS.n5012 DVSS 0.0162389
R5649 VSS.n3219 VSS.n2808 0.016
R5650 VSS.n3220 VSS.n3219 0.016
R5651 VSS.n3206 VSS.n3205 0.016
R5652 VSS.n3205 VSS.n3199 0.016
R5653 VSS.n3168 VSS.n3167 0.0155
R5654 VSS.n4916 VSS.n4915 0.0155
R5655 VSS.n3171 VSS.n3170 0.0155
R5656 VSS.n4912 VSS.n4911 0.0155
R5657 VSS.n5150 VSS.n5149 0.0154891
R5658 VSS.n2074 VSS.n1595 0.01535
R5659 VSS.n1819 VSS.n1797 0.01535
R5660 VSS.n3817 VSS.n3815 0.0152819
R5661 VSS.n3817 VSS.n3816 0.0152819
R5662 VSS.n3819 VSS.n3787 0.0152819
R5663 VSS.n3815 VSS.n3732 0.0152819
R5664 VSS.n3816 VSS.n3789 0.0152819
R5665 VSS.n3789 VSS.n3787 0.0152819
R5666 VSS.n4117 VSS.n4115 0.0152819
R5667 VSS.n4117 VSS.n4116 0.0152819
R5668 VSS.n4119 VSS.n3886 0.0152819
R5669 VSS.n4115 VSS.n3890 0.0152819
R5670 VSS.n4116 VSS.n3889 0.0152819
R5671 VSS.n3889 VSS.n3886 0.0152819
R5672 VSS.n635 VSS.n220 0.0152727
R5673 VSS.n3119 VSS.n2848 0.015
R5674 VSS.n4958 VSS.n2361 0.015
R5675 VSS.n3059 VSS.n2846 0.015
R5676 VSS.n4956 VSS.n2358 0.015
R5677 VSS.n4173 VSS.n2650 0.0149495
R5678 VSS.n4961 DVSS 0.0149089
R5679 DVSS VSS.n2357 0.0149089
R5680 VSS.n2072 VSS.n1592 0.0149069
R5681 VSS.n2071 VSS.n2070 0.0149069
R5682 VSS.n2071 VSS.n1593 0.0149069
R5683 VSS.n2068 VSS.n1593 0.0149069
R5684 VSS.n2067 VSS.n1592 0.0149069
R5685 VSS.n2070 VSS.n2067 0.0149069
R5686 VSS.n1816 VSS.n1815 0.0149069
R5687 VSS.n1814 VSS.n1813 0.0149069
R5688 VSS.n1812 VSS.n1810 0.0149069
R5689 VSS.n1813 VSS.n1812 0.0149069
R5690 VSS.n1815 VSS.n1814 0.0149069
R5691 VSS.n1817 VSS.n1816 0.0149069
R5692 VSS.n5706 VSS.n17 0.0145462
R5693 VSS.n1151 VSS.n17 0.0145462
R5694 VSS.n1153 VSS.n1151 0.0145462
R5695 VSS.n1155 VSS.n1153 0.0145462
R5696 VSS.n1156 VSS.n1155 0.0145462
R5697 VSS.n1159 VSS.n1156 0.0145462
R5698 VSS.n1161 VSS.n1159 0.0145462
R5699 VSS.n1163 VSS.n1161 0.0145462
R5700 VSS.n1164 VSS.n1163 0.0145462
R5701 VSS.n1167 VSS.n1164 0.0145462
R5702 VSS.n1168 VSS.n1167 0.0145462
R5703 VSS.n3839 VSS.n3821 0.0145367
R5704 VSS.n3081 VSS.n2872 0.0145
R5705 VSS.n5003 VSS.n2334 0.0145
R5706 VSS.n3076 VSS.n2877 0.0145
R5707 VSS.n5005 VSS.n2336 0.0145
R5708 VSS.n4347 VSS.n2608 0.0144402
R5709 VSS.n4336 VSS.n2611 0.0144402
R5710 VSS.n1302 VSS.n1300 0.0144028
R5711 VSS.n3995 VSS.n3994 0.0142903
R5712 VSS.n4073 VSS.n4066 0.0142838
R5713 VSS.n4381 VSS.n4380 0.0142814
R5714 VSS.n5189 VSS.n5188 0.0142814
R5715 VSS.n3861 VSS.n3859 0.0141679
R5716 VSS.n3862 VSS.n2616 0.0141679
R5717 VSS.n3862 VSS.n3859 0.0141679
R5718 VSS.n3864 VSS.n3861 0.0141679
R5719 VSS.n2976 VSS.n2914 0.014
R5720 VSS.n3020 VSS.n2894 0.014
R5721 VSS.n5067 VSS.n5066 0.014
R5722 VSS.n5096 VSS.n2292 0.014
R5723 VSS.n2965 VSS.n2919 0.014
R5724 VSS.n3015 VSS.n2899 0.014
R5725 VSS.n5063 VSS.n5062 0.014
R5726 VSS.n5100 VSS.n2294 0.014
R5727 VSS.n1150 VSS.n21 0.0136707
R5728 VSS.n1158 VSS.n1157 0.0136707
R5729 VSS.n1166 VSS.n1165 0.0136707
R5730 DVSS VSS.n4960 0.0135788
R5731 VSS.n4954 DVSS 0.0135788
R5732 VSS.n2068 VSS.n1595 0.01355
R5733 VSS.n1810 VSS.n1797 0.01355
R5734 VSS.n4532 VSS.n2545 0.0135392
R5735 VSS.n2972 VSS.n2916 0.0135
R5736 VSS.n3024 VSS.n2885 0.0135
R5737 VSS.n5046 VSS.n5045 0.0135
R5738 VSS.n5106 VSS.n2289 0.0135
R5739 VSS.n2969 VSS.n2918 0.0135
R5740 VSS.n3010 VSS.n2893 0.0135
R5741 VSS.n5049 VSS.n5048 0.0135
R5742 VSS.n5104 VSS.n2286 0.0135
R5743 VSS.n3841 VSS.n3820 0.0134255
R5744 VSS.n3867 VSS.n3820 0.0134255
R5745 VSS.n4071 VSS.n4068 0.0134255
R5746 VSS.n4070 VSS.n4068 0.0134255
R5747 VSS.n3857 VSS.n3856 0.0133402
R5748 VSS.n3847 VSS.n3846 0.0133402
R5749 VSS.n3085 VSS.n2862 0.013
R5750 VSS.n4999 VSS.n2341 0.013
R5751 VSS.n3071 VSS.n2871 0.013
R5752 VSS.n2345 VSS.n2339 0.013
R5753 VSS.n3853 VSS.n2564 0.0129835
R5754 VSS.n3849 VSS.n2558 0.0129835
R5755 VSS.n4344 VSS.n2608 0.0129728
R5756 VSS.n4338 VSS.n2611 0.0129728
R5757 VSS.n183 VSS.n104 0.0129415
R5758 VSS.n183 VSS.n182 0.0129415
R5759 VSS.n187 VSS.n182 0.0129415
R5760 VSS.n188 VSS.n187 0.0129415
R5761 VSS.n189 VSS.n188 0.0129415
R5762 VSS.n189 VSS.n180 0.0129415
R5763 VSS.n193 VSS.n180 0.0129415
R5764 VSS.n194 VSS.n193 0.0129415
R5765 VSS.n195 VSS.n194 0.0129415
R5766 VSS.n195 VSS.n178 0.0129415
R5767 VSS.n199 VSS.n178 0.0129415
R5768 VSS.n200 VSS.n199 0.0129415
R5769 VSS.n201 VSS.n200 0.0129415
R5770 VSS.n201 VSS.n176 0.0129415
R5771 VSS.n205 VSS.n176 0.0129415
R5772 VSS.n206 VSS.n205 0.0129415
R5773 VSS.n207 VSS.n206 0.0129415
R5774 VSS.n207 VSS.n174 0.0129415
R5775 VSS.n211 VSS.n174 0.0129415
R5776 VSS.n212 VSS.n211 0.0129415
R5777 VSS.n213 VSS.n212 0.0129415
R5778 VSS.n213 VSS.n172 0.0129415
R5779 VSS.n913 VSS.n912 0.0129415
R5780 VSS.n235 VSS.n218 0.0129415
R5781 VSS.n236 VSS.n235 0.0129415
R5782 VSS.n237 VSS.n236 0.0129415
R5783 VSS.n237 VSS.n231 0.0129415
R5784 VSS.n241 VSS.n231 0.0129415
R5785 VSS.n242 VSS.n241 0.0129415
R5786 VSS.n243 VSS.n242 0.0129415
R5787 VSS.n243 VSS.n229 0.0129415
R5788 VSS.n247 VSS.n229 0.0129415
R5789 VSS.n248 VSS.n247 0.0129415
R5790 VSS.n249 VSS.n248 0.0129415
R5791 VSS.n249 VSS.n227 0.0129415
R5792 VSS.n253 VSS.n227 0.0129415
R5793 VSS.n254 VSS.n253 0.0129415
R5794 VSS.n255 VSS.n254 0.0129415
R5795 VSS.n255 VSS.n225 0.0129415
R5796 VSS.n259 VSS.n225 0.0129415
R5797 VSS.n260 VSS.n259 0.0129415
R5798 VSS.n261 VSS.n260 0.0129415
R5799 VSS.n261 VSS.n223 0.0129415
R5800 VSS.n905 VSS.n223 0.0129415
R5801 VSS.n378 VSS.n373 0.0127609
R5802 VSS.n379 VSS.n377 0.0127609
R5803 VSS.n376 VSS.n374 0.0127528
R5804 VSS.n4169 VSS.n3722 0.01265
R5805 VSS.n3795 VSS.n3722 0.01265
R5806 VSS.n3124 VSS.n2841 0.0125
R5807 VSS.n4948 VSS.n2366 0.0125
R5808 VSS.n3126 VSS.n2843 0.0125
R5809 VSS.n4952 VSS.n2368 0.0125
R5810 VSS.n3942 VSS.n3941 0.0124725
R5811 VSS.n3752 VSS.n3751 0.0124725
R5812 VSS.n569 VSS.n568 0.0123471
R5813 VSS.n568 VSS.n567 0.0123471
R5814 VSS.n567 VSS.n525 0.0123471
R5815 VSS.n563 VSS.n525 0.0123471
R5816 VSS.n563 VSS.n562 0.0123471
R5817 VSS.n562 VSS.n561 0.0123471
R5818 VSS.n561 VSS.n527 0.0123471
R5819 VSS.n557 VSS.n527 0.0123471
R5820 VSS.n557 VSS.n556 0.0123471
R5821 VSS.n556 VSS.n555 0.0123471
R5822 VSS.n555 VSS.n529 0.0123471
R5823 VSS.n551 VSS.n529 0.0123471
R5824 VSS.n551 VSS.n550 0.0123471
R5825 VSS.n550 VSS.n549 0.0123471
R5826 VSS.n549 VSS.n531 0.0123471
R5827 VSS.n545 VSS.n531 0.0123471
R5828 VSS.n545 VSS.n544 0.0123471
R5829 VSS.n544 VSS.n543 0.0123471
R5830 VSS.n543 VSS.n533 0.0123471
R5831 VSS.n539 VSS.n533 0.0123471
R5832 VSS.n539 VSS.n538 0.0123471
R5833 VSS.n538 VSS.n537 0.0123471
R5834 VSS.n634 VSS.n633 0.0123471
R5835 VSS.n636 VSS.n363 0.0123471
R5836 VSS.n640 VSS.n363 0.0123471
R5837 VSS.n641 VSS.n640 0.0123471
R5838 VSS.n642 VSS.n641 0.0123471
R5839 VSS.n642 VSS.n361 0.0123471
R5840 VSS.n646 VSS.n361 0.0123471
R5841 VSS.n647 VSS.n646 0.0123471
R5842 VSS.n648 VSS.n647 0.0123471
R5843 VSS.n648 VSS.n359 0.0123471
R5844 VSS.n652 VSS.n359 0.0123471
R5845 VSS.n653 VSS.n652 0.0123471
R5846 VSS.n654 VSS.n653 0.0123471
R5847 VSS.n654 VSS.n357 0.0123471
R5848 VSS.n658 VSS.n357 0.0123471
R5849 VSS.n659 VSS.n658 0.0123471
R5850 VSS.n660 VSS.n659 0.0123471
R5851 VSS.n660 VSS.n355 0.0123471
R5852 VSS.n664 VSS.n355 0.0123471
R5853 VSS.n665 VSS.n664 0.0123471
R5854 VSS.n667 VSS.n665 0.0123471
R5855 VSS.n667 VSS.n666 0.0123471
R5856 VSS.n5705 VSS.n5704 0.0123293
R5857 VSS.n31 VSS.n27 0.0123293
R5858 VSS.n3860 VSS.n2561 0.0122701
R5859 VSS.n4513 VSS.n2567 0.0122701
R5860 DVSS VSS.n2321 0.0122488
R5861 VSS.n5009 DVSS 0.0122488
R5862 VSS.n3183 VSS.n3181 0.012
R5863 VSS.n4894 VSS.n4893 0.012
R5864 VSS.n3178 VSS.n3177 0.012
R5865 VSS.n4897 VSS.n4896 0.012
R5866 VSS.n4100 VSS.n4099 0.0116468
R5867 VSS.n5286 VSS.n2227 0.0116
R5868 VSS.n1154 VSS.n30 0.0115976
R5869 VSS.n1160 VSS.n26 0.0115976
R5870 VSS.n3233 VSS.n3232 0.0115
R5871 VSS.n3225 VSS.n3224 0.0115
R5872 VSS.n3203 VSS.n2810 0.0115
R5873 VSS.n3217 VSS.n3216 0.0115
R5874 VSS.n4165 VSS.n3726 0.0113969
R5875 VSS.n4165 VSS.n4164 0.0113969
R5876 VSS.n3951 VSS.n3950 0.0113969
R5877 VSS.n3950 VSS.n3949 0.0113969
R5878 VSS.n1771 VSS.n1769 0.0112561
R5879 VSS.n1785 VSS.n1775 0.0112561
R5880 VSS.n1918 VSS.n1917 0.0112561
R5881 VSS.n1901 VSS.n1898 0.0112561
R5882 VSS.n1956 VSS.n1955 0.0112561
R5883 VSS.n1939 VSS.n1936 0.0112561
R5884 VSS.n1987 VSS.n1677 0.0112561
R5885 VSS.n1976 VSS.n1686 0.0112561
R5886 VSS.n2019 VSS.n1650 0.0112561
R5887 VSS.n2008 VSS.n1661 0.0112561
R5888 VSS.n1627 VSS.n1625 0.0112561
R5889 VSS.n1641 VSS.n1631 0.0112561
R5890 VSS.n5311 VSS 0.0110882
R5891 VSS VSS.n5309 0.0110882
R5892 VSS.n4847 VSS 0.0110882
R5893 VSS.n5573 VSS.n1231 0.0110195
R5894 VSS.n3164 VSS.n2827 0.011
R5895 VSS.n4921 VSS.n2385 0.011
R5896 VSS.n2831 VSS.n2825 0.011
R5897 VSS.n4907 VSS.n2390 0.011
R5898 VSS.n4311 VSS.n4310 0.0109694
R5899 VSS.n4312 VSS.n4311 0.0109694
R5900 VSS.n4312 VSS.n2620 0.0109694
R5901 VSS.n4318 VSS.n2620 0.0109694
R5902 VSS.n4319 VSS.n4318 0.0109694
R5903 VSS.n4320 VSS.n4319 0.0109694
R5904 VSS.n4320 VSS.n2198 0.0109694
R5905 VSS.n5298 VSS.n2198 0.0109694
R5906 VSS.n5298 VSS.n5297 0.0109694
R5907 VSS.n4873 DVSS 0.0109187
R5908 VSS.n3212 DVSS 0.0109187
R5909 VSS.n5286 VSS.n5285 0.0109
R5910 VSS.n5285 VSS.n5280 0.0109
R5911 VSS.n5280 VSS.n5279 0.0109
R5912 VSS.n5279 VSS.n5278 0.0109
R5913 VSS.n5278 VSS.n5277 0.0109
R5914 VSS.n5277 VSS.n5276 0.0109
R5915 VSS.n5276 VSS.n5275 0.0109
R5916 VSS.n5275 VSS.n5274 0.0109
R5917 VSS.n5274 VSS.n5273 0.0109
R5918 VSS.n5273 VSS.n5272 0.0109
R5919 VSS.n5272 VSS.n5271 0.0109
R5920 VSS.n1152 VSS.n29 0.0108659
R5921 VSS.n1162 VSS.n24 0.0108659
R5922 VSS.n2974 VSS.n2915 0.010697
R5923 VSS.n2967 VSS.n2960 0.010697
R5924 VSS.n5565 VSS.n1231 0.0106855
R5925 VSS.n3118 VSS.n2850 0.0105
R5926 VSS.n4967 VSS.n4966 0.0105
R5927 VSS.n3061 VSS.n2852 0.0105
R5928 VSS.n4970 VSS.n4969 0.0105
R5929 VSS.n2944 VSS.n2929 0.0105
R5930 VSS.n2944 VSS.n2943 0.0105
R5931 VSS.n2943 VSS.n2942 0.0105
R5932 VSS.n2942 VSS.n2911 0.0105
R5933 VSS.n2980 VSS.n2911 0.0105
R5934 VSS.n2980 VSS.n2909 0.0105
R5935 VSS.n2988 VSS.n2909 0.0105
R5936 VSS.n2988 VSS.n2987 0.0105
R5937 VSS.n2987 VSS.n2986 0.0105
R5938 VSS.n2986 VSS.n2891 0.0105
R5939 VSS.n3027 VSS.n2891 0.0105
R5940 VSS.n3027 VSS.n2889 0.0105
R5941 VSS.n3039 VSS.n2889 0.0105
R5942 VSS.n3039 VSS.n3038 0.0105
R5943 VSS.n3038 VSS.n3035 0.0105
R5944 VSS.n3035 VSS.n3034 0.0105
R5945 VSS.n3034 VSS.n2869 0.0105
R5946 VSS.n3088 VSS.n2869 0.0105
R5947 VSS.n3088 VSS.n2867 0.0105
R5948 VSS.n3092 VSS.n2867 0.0105
R5949 VSS.n3092 VSS.n2856 0.0105
R5950 VSS.n3107 VSS.n2856 0.0105
R5951 VSS.n3107 VSS.n2854 0.0105
R5952 VSS.n3115 VSS.n2854 0.0105
R5953 VSS.n3115 VSS.n3114 0.0105
R5954 VSS.n3114 VSS.n3113 0.0105
R5955 VSS.n3113 VSS.n2836 0.0105
R5956 VSS.n3151 VSS.n2836 0.0105
R5957 VSS.n3151 VSS.n2834 0.0105
R5958 VSS.n3160 VSS.n2834 0.0105
R5959 VSS.n3160 VSS.n3159 0.0105
R5960 VSS.n3159 VSS.n3158 0.0105
R5961 VSS.n3158 VSS.n2814 0.0105
R5962 VSS.n3192 VSS.n2814 0.0105
R5963 VSS.n3193 VSS.n3192 0.0105
R5964 VSS.n3194 VSS.n3193 0.0105
R5965 VSS.n3194 VSS.n2812 0.0105
R5966 VSS.n3229 VSS.n2812 0.0105
R5967 VSS.n3229 VSS.n3228 0.0105
R5968 VSS.n3228 VSS.n2403 0.0105
R5969 VSS.n4878 VSS.n2403 0.0105
R5970 VSS.n4878 VSS.n2401 0.0105
R5971 VSS.n4886 VSS.n2401 0.0105
R5972 VSS.n4886 VSS.n4885 0.0105
R5973 VSS.n4885 VSS.n4884 0.0105
R5974 VSS.n4884 VSS.n2382 0.0105
R5975 VSS.n4925 VSS.n2382 0.0105
R5976 VSS.n4925 VSS.n2380 0.0105
R5977 VSS.n4939 VSS.n2380 0.0105
R5978 VSS.n4939 VSS.n4938 0.0105
R5979 VSS.n4938 VSS.n4937 0.0105
R5980 VSS.n4937 VSS.n4936 0.0105
R5981 VSS.n4936 VSS.n4935 0.0105
R5982 VSS.n4935 VSS.n4934 0.0105
R5983 VSS.n4934 VSS.n2350 0.0105
R5984 VSS.n4987 VSS.n2350 0.0105
R5985 VSS.n4987 VSS.n2348 0.0105
R5986 VSS.n4995 VSS.n2348 0.0105
R5987 VSS.n4995 VSS.n4994 0.0105
R5988 VSS.n4994 VSS.n4993 0.0105
R5989 VSS.n4993 VSS.n2329 0.0105
R5990 VSS.n5030 VSS.n2329 0.0105
R5991 VSS.n5030 VSS.n2327 0.0105
R5992 VSS.n5038 VSS.n2327 0.0105
R5993 VSS.n5038 VSS.n5037 0.0105
R5994 VSS.n5037 VSS.n5036 0.0105
R5995 VSS.n5036 VSS.n2308 0.0105
R5996 VSS.n5076 VSS.n2308 0.0105
R5997 VSS.n5076 VSS.n2306 0.0105
R5998 VSS.n5088 VSS.n2306 0.0105
R5999 VSS.n5088 VSS.n5087 0.0105
R6000 VSS.n5087 VSS.n5086 0.0105
R6001 VSS.n5086 VSS.n5085 0.0105
R6002 VSS.n5085 VSS.n5084 0.0105
R6003 VSS.n5084 VSS.n2282 0.0105
R6004 VSS.n5128 VSS.n2282 0.0105
R6005 VSS.n5128 VSS.n2280 0.0105
R6006 VSS.n5168 VSS.n2280 0.0105
R6007 VSS.n5168 VSS.n5167 0.0105
R6008 VSS.n5167 VSS.n5166 0.0105
R6009 VSS.n5166 VSS.n5134 0.0105
R6010 VSS.n5162 VSS.n5134 0.0105
R6011 VSS.n5162 VSS.n5161 0.0105
R6012 VSS.n5161 VSS.n5139 0.0105
R6013 VSS.n5157 VSS.n5139 0.0105
R6014 VSS.n5157 VSS.n5156 0.0105
R6015 VSS.n5156 VSS.n5155 0.0105
R6016 VSS.n5155 VSS.n5145 0.0105
R6017 VSS.n5151 VSS.n5145 0.0105
R6018 VSS.n5169 VSS.n2279 0.0105
R6019 VSS.n5165 VSS.n2279 0.0105
R6020 VSS.n5165 VSS.n5164 0.0105
R6021 VSS.n5164 VSS.n5163 0.0105
R6022 VSS.n5160 VSS.n5159 0.0105
R6023 VSS.n5159 VSS.n5158 0.0105
R6024 VSS.n5158 VSS.n5140 0.0105
R6025 VSS.n5154 VSS.n5140 0.0105
R6026 VSS.n5154 VSS.n5153 0.0105
R6027 VSS.n5153 VSS.n5152 0.0105
R6028 VSS.n5160 VSS.n5135 0.0104296
R6029 VSS.n1772 VSS.n1771 0.0101185
R6030 VSS.n1786 VSS.n1785 0.0101185
R6031 VSS.n1918 VSS.n1726 0.0101185
R6032 VSS.n1903 VSS.n1898 0.0101185
R6033 VSS.n1956 VSS.n1702 0.0101185
R6034 VSS.n1941 VSS.n1936 0.0101185
R6035 VSS.n1988 VSS.n1987 0.0101185
R6036 VSS.n1974 VSS.n1686 0.0101185
R6037 VSS.n2020 VSS.n2019 0.0101185
R6038 VSS.n2006 VSS.n1661 0.0101185
R6039 VSS.n1628 VSS.n1627 0.0101185
R6040 VSS.n1642 VSS.n1641 0.0101185
R6041 VSS.n5696 VSS.n1149 0.0100456
R6042 VSS.n5701 VSS.n5700 0.0100456
R6043 VSS.n5697 VSS.n5696 0.0100456
R6044 VSS.n1146 VSS.n1145 0.0100456
R6045 VSS.n3080 VSS.n2874 0.01
R6046 VSS.n5022 VSS.n5020 0.01
R6047 VSS.n3077 VSS.n2876 0.01
R6048 VSS.n5017 VSS.n5016 0.01
R6049 VSS.n3604 DVSS 0.00997368
R6050 VSS.n3863 VSS.n2560 0.00965456
R6051 VSS.n3843 VSS.n2566 0.00965456
R6052 VSS.n2769 VSS.n2763 0.00962857
R6053 VSS.n2769 VSS.n2761 0.00962857
R6054 VSS.n2773 VSS.n2761 0.00962857
R6055 VSS.n2773 VSS.n2759 0.00962857
R6056 VSS.n2777 VSS.n2759 0.00962857
R6057 VSS.n2777 VSS.n2757 0.00962857
R6058 VSS.n2781 VSS.n2757 0.00962857
R6059 VSS.n2781 VSS.n2755 0.00962857
R6060 VSS.n2785 VSS.n2755 0.00962857
R6061 VSS.n2785 VSS.n2753 0.00962857
R6062 VSS.n2789 VSS.n2753 0.00962857
R6063 VSS.n2789 VSS.n2751 0.00962857
R6064 VSS.n3264 VSS.n2751 0.00962857
R6065 VSS.n3264 VSS.n2749 0.00962857
R6066 VSS.n3268 VSS.n2749 0.00962857
R6067 VSS.n3268 VSS.n2747 0.00962857
R6068 VSS.n3272 VSS.n2747 0.00962857
R6069 VSS.n3272 VSS.n2745 0.00962857
R6070 VSS.n3276 VSS.n2745 0.00962857
R6071 VSS.n3276 VSS.n2743 0.00962857
R6072 VSS.n3280 VSS.n2743 0.00962857
R6073 VSS.n3280 VSS.n2741 0.00962857
R6074 VSS.n3284 VSS.n2741 0.00962857
R6075 VSS.n3284 VSS.n2739 0.00962857
R6076 VSS.n3288 VSS.n2739 0.00962857
R6077 VSS.n3288 VSS.n2736 0.00962857
R6078 VSS.n3515 VSS.n2736 0.00962857
R6079 VSS.n3515 VSS.n2737 0.00962857
R6080 VSS.n3511 VSS.n2737 0.00962857
R6081 VSS.n3511 VSS.n3292 0.00962857
R6082 VSS.n3507 VSS.n3292 0.00962857
R6083 VSS.n3507 VSS.n3294 0.00962857
R6084 VSS.n3503 VSS.n3294 0.00962857
R6085 VSS.n3503 VSS.n3296 0.00962857
R6086 VSS.n3499 VSS.n3296 0.00962857
R6087 VSS.n3499 VSS.n3298 0.00962857
R6088 VSS.n3495 VSS.n3298 0.00962857
R6089 VSS.n3495 VSS.n3300 0.00962857
R6090 VSS.n3491 VSS.n3300 0.00962857
R6091 VSS.n3491 VSS.n3302 0.00962857
R6092 VSS.n3487 VSS.n3302 0.00962857
R6093 VSS.n3487 VSS.n3304 0.00962857
R6094 VSS.n3483 VSS.n3304 0.00962857
R6095 VSS.n3483 VSS.n3306 0.00962857
R6096 VSS.n3479 VSS.n3306 0.00962857
R6097 VSS.n3479 VSS.n3308 0.00962857
R6098 VSS.n3475 VSS.n3308 0.00962857
R6099 VSS.n3475 VSS.n3310 0.00962857
R6100 VSS.n3471 VSS.n3310 0.00962857
R6101 VSS.n3471 VSS.n3312 0.00962857
R6102 VSS.n3467 VSS.n3312 0.00962857
R6103 VSS.n3467 VSS.n3314 0.00962857
R6104 VSS.n3463 VSS.n3314 0.00962857
R6105 VSS.n3463 VSS.n3316 0.00962857
R6106 VSS.n3459 VSS.n3316 0.00962857
R6107 VSS.n3459 VSS.n3318 0.00962857
R6108 VSS.n3455 VSS.n3318 0.00962857
R6109 VSS.n3455 VSS.n3320 0.00962857
R6110 VSS.n3451 VSS.n3320 0.00962857
R6111 VSS.n3451 VSS.n3322 0.00962857
R6112 VSS.n3447 VSS.n3322 0.00962857
R6113 VSS.n3447 VSS.n3324 0.00962857
R6114 VSS.n3443 VSS.n3324 0.00962857
R6115 VSS.n3443 VSS.n3326 0.00962857
R6116 VSS.n3439 VSS.n3326 0.00962857
R6117 VSS.n3439 VSS.n3328 0.00962857
R6118 VSS.n3435 VSS.n3328 0.00962857
R6119 VSS.n3435 VSS.n3330 0.00962857
R6120 VSS.n3431 VSS.n3330 0.00962857
R6121 VSS.n3431 VSS.n3332 0.00962857
R6122 VSS.n3427 VSS.n3332 0.00962857
R6123 VSS.n3427 VSS.n3334 0.00962857
R6124 VSS.n3423 VSS.n3334 0.00962857
R6125 VSS.n3423 VSS.n3336 0.00962857
R6126 VSS.n3419 VSS.n3336 0.00962857
R6127 VSS.n3419 VSS.n3338 0.00962857
R6128 VSS.n3415 VSS.n3338 0.00962857
R6129 VSS.n3415 VSS.n3340 0.00962857
R6130 VSS.n3411 VSS.n3340 0.00962857
R6131 VSS.n3411 VSS.n3342 0.00962857
R6132 VSS.n3407 VSS.n3342 0.00962857
R6133 VSS.n3407 VSS.n3344 0.00962857
R6134 VSS.n3403 VSS.n3344 0.00962857
R6135 VSS.n3403 VSS.n3346 0.00962857
R6136 VSS.n3399 VSS.n3346 0.00962857
R6137 VSS.n3399 VSS.n3348 0.00962857
R6138 VSS.n3395 VSS.n3348 0.00962857
R6139 VSS.n3395 VSS.n3350 0.00962857
R6140 VSS.n3391 VSS.n3350 0.00962857
R6141 VSS.n3391 VSS.n3352 0.00962857
R6142 VSS.n3387 VSS.n3352 0.00962857
R6143 VSS.n3387 VSS.n3354 0.00962857
R6144 VSS.n3383 VSS.n3354 0.00962857
R6145 VSS.n3383 VSS.n3356 0.00962857
R6146 VSS.n3379 VSS.n3356 0.00962857
R6147 VSS.n3379 VSS.n3357 0.00962857
R6148 VSS.n3375 VSS.n3357 0.00962857
R6149 VSS.n3374 VSS.n3368 0.00962857
R6150 VSS.n3368 VSS.n3359 0.00962857
R6151 VSS.n3364 VSS.n3359 0.00962857
R6152 VSS.n4189 VSS.n4188 0.00962857
R6153 VSS.n4188 VSS.n2640 0.00962857
R6154 VSS.n4184 VSS.n2640 0.00962857
R6155 VSS.n4184 VSS.n2642 0.00962857
R6156 VSS.n4180 VSS.n2642 0.00962857
R6157 VSS.n4180 VSS.n2645 0.00962857
R6158 VSS.n4176 VSS.n2645 0.00962857
R6159 VSS.n4176 VSS.n2647 0.00962857
R6160 VSS.n3799 VSS.n2647 0.00962857
R6161 VSS.n3802 VSS.n3799 0.00962857
R6162 VSS.n3802 VSS.n3793 0.00962857
R6163 VSS.n3808 VSS.n3793 0.00962857
R6164 VSS.n3808 VSS.n3791 0.00962857
R6165 VSS.n3812 VSS.n3791 0.00962857
R6166 VSS.n3812 VSS.n3736 0.00962857
R6167 VSS.n4159 VSS.n3736 0.00962857
R6168 VSS.n4159 VSS.n3737 0.00962857
R6169 VSS.n4155 VSS.n3737 0.00962857
R6170 VSS.n4155 VSS.n3740 0.00962857
R6171 VSS.n3874 VSS.n3740 0.00962857
R6172 VSS.n3874 VSS.n3763 0.00962857
R6173 VSS.n4141 VSS.n3763 0.00962857
R6174 VSS.n4141 VSS.n3764 0.00962857
R6175 VSS.n4137 VSS.n3764 0.00962857
R6176 VSS.n4137 VSS.n3767 0.00962857
R6177 VSS.n3917 VSS.n3767 0.00962857
R6178 VSS.n3933 VSS.n3917 0.00962857
R6179 VSS.n3933 VSS.n3913 0.00962857
R6180 VSS.n3938 VSS.n3913 0.00962857
R6181 VSS.n3938 VSS.n3915 0.00962857
R6182 VSS.n3915 VSS.n3894 0.00962857
R6183 VSS.n4112 VSS.n3894 0.00962857
R6184 VSS.n4112 VSS.n3895 0.00962857
R6185 VSS.n4108 VSS.n3895 0.00962857
R6186 VSS.n4108 VSS.n3898 0.00962857
R6187 VSS.n3959 VSS.n3898 0.00962857
R6188 VSS.n4096 VSS.n3959 0.00962857
R6189 VSS.n4096 VSS.n3960 0.00962857
R6190 VSS.n4092 VSS.n3960 0.00962857
R6191 VSS.n4092 VSS.n3963 0.00962857
R6192 VSS.n4054 VSS.n3963 0.00962857
R6193 VSS.n4054 VSS.n3967 0.00962857
R6194 VSS.n4050 VSS.n3967 0.00962857
R6195 VSS.n4050 VSS.n3969 0.00962857
R6196 VSS.n4046 VSS.n3969 0.00962857
R6197 VSS.n4046 VSS.n3971 0.00962857
R6198 VSS.n4042 VSS.n3971 0.00962857
R6199 VSS.n4042 VSS.n3973 0.00962857
R6200 VSS.n4038 VSS.n3973 0.00962857
R6201 VSS.n4038 VSS.n3975 0.00962857
R6202 VSS.n4034 VSS.n3975 0.00962857
R6203 VSS.n4034 VSS.n3977 0.00962857
R6204 VSS.n4030 VSS.n3977 0.00962857
R6205 VSS.n4030 VSS.n3979 0.00962857
R6206 VSS.n4026 VSS.n3979 0.00962857
R6207 VSS.n4026 VSS.n3981 0.00962857
R6208 VSS.n4022 VSS.n3981 0.00962857
R6209 VSS.n4022 VSS.n3983 0.00962857
R6210 VSS.n4018 VSS.n3983 0.00962857
R6211 VSS.n4018 VSS.n3985 0.00962857
R6212 VSS.n4014 VSS.n3985 0.00962857
R6213 VSS.n4014 VSS.n3987 0.00962857
R6214 VSS.n4010 VSS.n3987 0.00962857
R6215 VSS.n4010 VSS.n3989 0.00962857
R6216 VSS.n4006 VSS.n3989 0.00962857
R6217 VSS.n4006 VSS.n3991 0.00962857
R6218 VSS.n4002 VSS.n3991 0.00962857
R6219 VSS.n4002 VSS.n3993 0.00962857
R6220 VSS.n3998 VSS.n3993 0.00962857
R6221 VSS.n4525 VSS.n4524 0.00962857
R6222 VSS.n4524 VSS.n2549 0.00962857
R6223 VSS.n4520 VSS.n2549 0.00962857
R6224 VSS.n4520 VSS.n2552 0.00962857
R6225 VSS.n4516 VSS.n2552 0.00962857
R6226 VSS.n4516 VSS.n2555 0.00962857
R6227 VSS.n4510 VSS.n2555 0.00962857
R6228 VSS.n4510 VSS.n2570 0.00962857
R6229 VSS.n4506 VSS.n2570 0.00962857
R6230 VSS.n4506 VSS.n2572 0.00962857
R6231 VSS.n4502 VSS.n2572 0.00962857
R6232 VSS.n4502 VSS.n2574 0.00962857
R6233 VSS.n4498 VSS.n2574 0.00962857
R6234 VSS.n4498 VSS.n2576 0.00962857
R6235 VSS.n4494 VSS.n2576 0.00962857
R6236 VSS.n4494 VSS.n2578 0.00962857
R6237 VSS.n4490 VSS.n2578 0.00962857
R6238 VSS.n4490 VSS.n2580 0.00962857
R6239 VSS.n4486 VSS.n2580 0.00962857
R6240 VSS.n4486 VSS.n2582 0.00962857
R6241 VSS.n4482 VSS.n2582 0.00962857
R6242 VSS.n4482 VSS.n2584 0.00962857
R6243 VSS.n4478 VSS.n2584 0.00962857
R6244 VSS.n4478 VSS.n2586 0.00962857
R6245 VSS.n4474 VSS.n2586 0.00962857
R6246 VSS.n4474 VSS.n2588 0.00962857
R6247 VSS.n4470 VSS.n2588 0.00962857
R6248 VSS.n4470 VSS.n2590 0.00962857
R6249 VSS.n4466 VSS.n2590 0.00962857
R6250 VSS.n4466 VSS.n2592 0.00962857
R6251 VSS.n4462 VSS.n2592 0.00962857
R6252 VSS.n4462 VSS.n2594 0.00962857
R6253 VSS.n4458 VSS.n2594 0.00962857
R6254 VSS.n4458 VSS.n2596 0.00962857
R6255 VSS.n4454 VSS.n2596 0.00962857
R6256 VSS.n4454 VSS.n2598 0.00962857
R6257 VSS.n4450 VSS.n2598 0.00962857
R6258 VSS.n4450 VSS.n2600 0.00962857
R6259 VSS.n4446 VSS.n2600 0.00962857
R6260 VSS.n4446 VSS.n2602 0.00962857
R6261 VSS.n4442 VSS.n2602 0.00962857
R6262 VSS.n4442 VSS.n2604 0.00962857
R6263 VSS.n4352 VSS.n2604 0.00962857
R6264 VSS.n4352 VSS.n4350 0.00962857
R6265 VSS.n4435 VSS.n4350 0.00962857
R6266 VSS.n4435 VSS.n4351 0.00962857
R6267 VSS.n4431 VSS.n4351 0.00962857
R6268 VSS.n4431 VSS.n4356 0.00962857
R6269 VSS.n4427 VSS.n4356 0.00962857
R6270 VSS.n4427 VSS.n4358 0.00962857
R6271 VSS.n4423 VSS.n4358 0.00962857
R6272 VSS.n4423 VSS.n4360 0.00962857
R6273 VSS.n4419 VSS.n4360 0.00962857
R6274 VSS.n4419 VSS.n4362 0.00962857
R6275 VSS.n4415 VSS.n4362 0.00962857
R6276 VSS.n4415 VSS.n4364 0.00962857
R6277 VSS.n4411 VSS.n4364 0.00962857
R6278 VSS.n4411 VSS.n4366 0.00962857
R6279 VSS.n4407 VSS.n4366 0.00962857
R6280 VSS.n4407 VSS.n4368 0.00962857
R6281 VSS.n4403 VSS.n4368 0.00962857
R6282 VSS.n4403 VSS.n4370 0.00962857
R6283 VSS.n4399 VSS.n4370 0.00962857
R6284 VSS.n4399 VSS.n4372 0.00962857
R6285 VSS.n4395 VSS.n4372 0.00962857
R6286 VSS.n4395 VSS.n4374 0.00962857
R6287 VSS.n4391 VSS.n4374 0.00962857
R6288 VSS.n4391 VSS.n4376 0.00962857
R6289 VSS.n4387 VSS.n4376 0.00962857
R6290 VSS.n4387 VSS.n4378 0.00962857
R6291 VSS.n4383 VSS.n4378 0.00962857
R6292 VSS.n4523 VSS.n4522 0.00962857
R6293 VSS.n4522 VSS.n4521 0.00962857
R6294 VSS.n4521 VSS.n2551 0.00962857
R6295 VSS.n4511 VSS.n2569 0.00962857
R6296 VSS.n4505 VSS.n2569 0.00962857
R6297 VSS.n4505 VSS.n4504 0.00962857
R6298 VSS.n4504 VSS.n4503 0.00962857
R6299 VSS.n4503 VSS.n2573 0.00962857
R6300 VSS.n4497 VSS.n2573 0.00962857
R6301 VSS.n4497 VSS.n4496 0.00962857
R6302 VSS.n4496 VSS.n4495 0.00962857
R6303 VSS.n4495 VSS.n2577 0.00962857
R6304 VSS.n4489 VSS.n2577 0.00962857
R6305 VSS.n4489 VSS.n4488 0.00962857
R6306 VSS.n4488 VSS.n4487 0.00962857
R6307 VSS.n4487 VSS.n2581 0.00962857
R6308 VSS.n4481 VSS.n2581 0.00962857
R6309 VSS.n4481 VSS.n4480 0.00962857
R6310 VSS.n4480 VSS.n4479 0.00962857
R6311 VSS.n4479 VSS.n2585 0.00962857
R6312 VSS.n4473 VSS.n2585 0.00962857
R6313 VSS.n4473 VSS.n4472 0.00962857
R6314 VSS.n4472 VSS.n4471 0.00962857
R6315 VSS.n4471 VSS.n2589 0.00962857
R6316 VSS.n4465 VSS.n2589 0.00962857
R6317 VSS.n4465 VSS.n4464 0.00962857
R6318 VSS.n4464 VSS.n4463 0.00962857
R6319 VSS.n4463 VSS.n2593 0.00962857
R6320 VSS.n4457 VSS.n2593 0.00962857
R6321 VSS.n4457 VSS.n4456 0.00962857
R6322 VSS.n4456 VSS.n4455 0.00962857
R6323 VSS.n4455 VSS.n2597 0.00962857
R6324 VSS.n4449 VSS.n2597 0.00962857
R6325 VSS.n4449 VSS.n4448 0.00962857
R6326 VSS.n4448 VSS.n4447 0.00962857
R6327 VSS.n4447 VSS.n2601 0.00962857
R6328 VSS.n4441 VSS.n2601 0.00962857
R6329 VSS.n4441 VSS.n4440 0.00962857
R6330 VSS.n4436 VSS.n4349 0.00962857
R6331 VSS.n4430 VSS.n4349 0.00962857
R6332 VSS.n4430 VSS.n4429 0.00962857
R6333 VSS.n4429 VSS.n4428 0.00962857
R6334 VSS.n4428 VSS.n4357 0.00962857
R6335 VSS.n4422 VSS.n4357 0.00962857
R6336 VSS.n4422 VSS.n4421 0.00962857
R6337 VSS.n4421 VSS.n4420 0.00962857
R6338 VSS.n4420 VSS.n4361 0.00962857
R6339 VSS.n4414 VSS.n4361 0.00962857
R6340 VSS.n4414 VSS.n4413 0.00962857
R6341 VSS.n4413 VSS.n4412 0.00962857
R6342 VSS.n4412 VSS.n4365 0.00962857
R6343 VSS.n4406 VSS.n4365 0.00962857
R6344 VSS.n4406 VSS.n4405 0.00962857
R6345 VSS.n4405 VSS.n4404 0.00962857
R6346 VSS.n4404 VSS.n4369 0.00962857
R6347 VSS.n4398 VSS.n4369 0.00962857
R6348 VSS.n4398 VSS.n4397 0.00962857
R6349 VSS.n4397 VSS.n4396 0.00962857
R6350 VSS.n4396 VSS.n4373 0.00962857
R6351 VSS.n4390 VSS.n4373 0.00962857
R6352 VSS.n4390 VSS.n4389 0.00962857
R6353 VSS.n4389 VSS.n4388 0.00962857
R6354 VSS.n4388 VSS.n4377 0.00962857
R6355 VSS.n4382 VSS.n4377 0.00962857
R6356 VSS.n2060 VSS.n1613 0.00962857
R6357 VSS.n2060 VSS.n1614 0.00962857
R6358 VSS.n2056 VSS.n1614 0.00962857
R6359 VSS.n2056 VSS.n1616 0.00962857
R6360 VSS.n2052 VSS.n1616 0.00962857
R6361 VSS.n2052 VSS.n1619 0.00962857
R6362 VSS.n2048 VSS.n1619 0.00962857
R6363 VSS.n2048 VSS.n1621 0.00962857
R6364 VSS.n1635 VSS.n1621 0.00962857
R6365 VSS.n2036 VSS.n1635 0.00962857
R6366 VSS.n2036 VSS.n1636 0.00962857
R6367 VSS.n2032 VSS.n1636 0.00962857
R6368 VSS.n2032 VSS.n1639 0.00962857
R6369 VSS.n2028 VSS.n1639 0.00962857
R6370 VSS.n2028 VSS.n1645 0.00962857
R6371 VSS.n2024 VSS.n1645 0.00962857
R6372 VSS.n2024 VSS.n1647 0.00962857
R6373 VSS.n1652 VSS.n1647 0.00962857
R6374 VSS.n2016 VSS.n1652 0.00962857
R6375 VSS.n2016 VSS.n1653 0.00962857
R6376 VSS.n2012 VSS.n1653 0.00962857
R6377 VSS.n2012 VSS.n1656 0.00962857
R6378 VSS.n1666 VSS.n1656 0.00962857
R6379 VSS.n2003 VSS.n1666 0.00962857
R6380 VSS.n2003 VSS.n1667 0.00962857
R6381 VSS.n1999 VSS.n1667 0.00962857
R6382 VSS.n1999 VSS.n1670 0.00962857
R6383 VSS.n1995 VSS.n1670 0.00962857
R6384 VSS.n1995 VSS.n1672 0.00962857
R6385 VSS.n1991 VSS.n1672 0.00962857
R6386 VSS.n1991 VSS.n1674 0.00962857
R6387 VSS.n1984 VSS.n1674 0.00962857
R6388 VSS.n1984 VSS.n1679 0.00962857
R6389 VSS.n1980 VSS.n1679 0.00962857
R6390 VSS.n1980 VSS.n1681 0.00962857
R6391 VSS.n1691 VSS.n1681 0.00962857
R6392 VSS.n1971 VSS.n1691 0.00962857
R6393 VSS.n1971 VSS.n1692 0.00962857
R6394 VSS.n1967 VSS.n1692 0.00962857
R6395 VSS.n1967 VSS.n1695 0.00962857
R6396 VSS.n1963 VSS.n1695 0.00962857
R6397 VSS.n1963 VSS.n1697 0.00962857
R6398 VSS.n1959 VSS.n1697 0.00962857
R6399 VSS.n1959 VSS.n1699 0.00962857
R6400 VSS.n1709 VSS.n1699 0.00962857
R6401 VSS.n1948 VSS.n1709 0.00962857
R6402 VSS.n1948 VSS.n1710 0.00962857
R6403 VSS.n1944 VSS.n1710 0.00962857
R6404 VSS.n1944 VSS.n1713 0.00962857
R6405 VSS.n1933 VSS.n1713 0.00962857
R6406 VSS.n1933 VSS.n1717 0.00962857
R6407 VSS.n1929 VSS.n1717 0.00962857
R6408 VSS.n1929 VSS.n1719 0.00962857
R6409 VSS.n1925 VSS.n1719 0.00962857
R6410 VSS.n1925 VSS.n1721 0.00962857
R6411 VSS.n1921 VSS.n1721 0.00962857
R6412 VSS.n1921 VSS.n1723 0.00962857
R6413 VSS.n1751 VSS.n1723 0.00962857
R6414 VSS.n1910 VSS.n1751 0.00962857
R6415 VSS.n1910 VSS.n1752 0.00962857
R6416 VSS.n1906 VSS.n1752 0.00962857
R6417 VSS.n1906 VSS.n1755 0.00962857
R6418 VSS.n1895 VSS.n1755 0.00962857
R6419 VSS.n1895 VSS.n1759 0.00962857
R6420 VSS.n1891 VSS.n1759 0.00962857
R6421 VSS.n1891 VSS.n1761 0.00962857
R6422 VSS.n1887 VSS.n1761 0.00962857
R6423 VSS.n1887 VSS.n1763 0.00962857
R6424 VSS.n1883 VSS.n1763 0.00962857
R6425 VSS.n1883 VSS.n1765 0.00962857
R6426 VSS.n1779 VSS.n1765 0.00962857
R6427 VSS.n1871 VSS.n1779 0.00962857
R6428 VSS.n1871 VSS.n1780 0.00962857
R6429 VSS.n1867 VSS.n1780 0.00962857
R6430 VSS.n1867 VSS.n1783 0.00962857
R6431 VSS.n1863 VSS.n1783 0.00962857
R6432 VSS.n1863 VSS.n1789 0.00962857
R6433 VSS.n1859 VSS.n1789 0.00962857
R6434 VSS.n1859 VSS.n1791 0.00962857
R6435 VSS.n1852 VSS.n1791 0.00962857
R6436 VSS.n1852 VSS.n1822 0.00962857
R6437 VSS.n1848 VSS.n1822 0.00962857
R6438 VSS.n1848 VSS.n1824 0.00962857
R6439 VSS.n1844 VSS.n1824 0.00962857
R6440 VSS.n1844 VSS.n1826 0.00962857
R6441 VSS.n1840 VSS.n1826 0.00962857
R6442 VSS.n1839 VSS.n1837 0.00962857
R6443 VSS.n1837 VSS.n1828 0.00962857
R6444 VSS.n1833 VSS.n1828 0.00962857
R6445 VSS.n2055 VSS.n1617 0.00962857
R6446 VSS.n2055 VSS.n2054 0.00962857
R6447 VSS.n2054 VSS.n2053 0.00962857
R6448 VSS.n2031 VSS.n2030 0.00962857
R6449 VSS.n2030 VSS.n2029 0.00962857
R6450 VSS.n2029 VSS.n1644 0.00962857
R6451 VSS.n2023 VSS.n1644 0.00962857
R6452 VSS.n2023 VSS.n2022 0.00962857
R6453 VSS.n2004 VSS.n1665 0.00962857
R6454 VSS.n1998 VSS.n1665 0.00962857
R6455 VSS.n1998 VSS.n1997 0.00962857
R6456 VSS.n1997 VSS.n1996 0.00962857
R6457 VSS.n1996 VSS.n1671 0.00962857
R6458 VSS.n1990 VSS.n1671 0.00962857
R6459 VSS.n1972 VSS.n1690 0.00962857
R6460 VSS.n1966 VSS.n1690 0.00962857
R6461 VSS.n1966 VSS.n1965 0.00962857
R6462 VSS.n1965 VSS.n1964 0.00962857
R6463 VSS.n1964 VSS.n1696 0.00962857
R6464 VSS.n1935 VSS.n1934 0.00962857
R6465 VSS.n1934 VSS.n1716 0.00962857
R6466 VSS.n1928 VSS.n1716 0.00962857
R6467 VSS.n1928 VSS.n1927 0.00962857
R6468 VSS.n1927 VSS.n1926 0.00962857
R6469 VSS.n1926 VSS.n1720 0.00962857
R6470 VSS.n1897 VSS.n1896 0.00962857
R6471 VSS.n1896 VSS.n1758 0.00962857
R6472 VSS.n1890 VSS.n1758 0.00962857
R6473 VSS.n1890 VSS.n1889 0.00962857
R6474 VSS.n1889 VSS.n1888 0.00962857
R6475 VSS.n1866 VSS.n1865 0.00962857
R6476 VSS.n1865 VSS.n1864 0.00962857
R6477 VSS.n1864 VSS.n1788 0.00962857
R6478 VSS.n1853 VSS.n1821 0.00962857
R6479 VSS.n1847 VSS.n1821 0.00962857
R6480 VSS.n1847 VSS.n1846 0.00962857
R6481 VSS.n1846 VSS.n1845 0.00962857
R6482 VSS.n1845 VSS.n1825 0.00962857
R6483 VSS.n1825 VSS.n23 0.00962857
R6484 VSS.n1836 VSS.n1835 0.00962857
R6485 VSS.n1835 VSS.n1834 0.00962857
R6486 VSS.n1585 VSS.n1300 0.00962857
R6487 VSS.n1585 VSS.n1301 0.00962857
R6488 VSS.n1581 VSS.n1301 0.00962857
R6489 VSS.n1581 VSS.n1304 0.00962857
R6490 VSS.n1577 VSS.n1304 0.00962857
R6491 VSS.n1577 VSS.n1306 0.00962857
R6492 VSS.n1573 VSS.n1306 0.00962857
R6493 VSS.n1573 VSS.n1308 0.00962857
R6494 VSS.n1569 VSS.n1308 0.00962857
R6495 VSS.n1569 VSS.n1310 0.00962857
R6496 VSS.n1565 VSS.n1310 0.00962857
R6497 VSS.n1565 VSS.n1312 0.00962857
R6498 VSS.n1561 VSS.n1312 0.00962857
R6499 VSS.n1561 VSS.n1314 0.00962857
R6500 VSS.n1557 VSS.n1314 0.00962857
R6501 VSS.n1557 VSS.n1316 0.00962857
R6502 VSS.n1553 VSS.n1316 0.00962857
R6503 VSS.n1553 VSS.n1318 0.00962857
R6504 VSS.n1549 VSS.n1318 0.00962857
R6505 VSS.n1549 VSS.n1320 0.00962857
R6506 VSS.n1545 VSS.n1320 0.00962857
R6507 VSS.n1545 VSS.n1322 0.00962857
R6508 VSS.n1541 VSS.n1322 0.00962857
R6509 VSS.n1541 VSS.n1324 0.00962857
R6510 VSS.n1537 VSS.n1324 0.00962857
R6511 VSS.n1537 VSS.n1326 0.00962857
R6512 VSS.n1533 VSS.n1326 0.00962857
R6513 VSS.n1533 VSS.n1328 0.00962857
R6514 VSS.n1529 VSS.n1328 0.00962857
R6515 VSS.n1529 VSS.n1330 0.00962857
R6516 VSS.n1525 VSS.n1330 0.00962857
R6517 VSS.n1525 VSS.n1332 0.00962857
R6518 VSS.n1521 VSS.n1332 0.00962857
R6519 VSS.n1521 VSS.n1334 0.00962857
R6520 VSS.n1517 VSS.n1334 0.00962857
R6521 VSS.n1517 VSS.n1336 0.00962857
R6522 VSS.n1513 VSS.n1336 0.00962857
R6523 VSS.n1513 VSS.n1338 0.00962857
R6524 VSS.n1509 VSS.n1338 0.00962857
R6525 VSS.n1509 VSS.n1340 0.00962857
R6526 VSS.n1505 VSS.n1340 0.00962857
R6527 VSS.n1505 VSS.n1342 0.00962857
R6528 VSS.n1501 VSS.n1342 0.00962857
R6529 VSS.n1501 VSS.n1344 0.00962857
R6530 VSS.n1497 VSS.n1344 0.00962857
R6531 VSS.n1497 VSS.n1346 0.00962857
R6532 VSS.n1493 VSS.n1346 0.00962857
R6533 VSS.n1493 VSS.n1348 0.00962857
R6534 VSS.n1489 VSS.n1348 0.00962857
R6535 VSS.n1489 VSS.n1350 0.00962857
R6536 VSS.n1485 VSS.n1350 0.00962857
R6537 VSS.n1485 VSS.n1352 0.00962857
R6538 VSS.n1481 VSS.n1352 0.00962857
R6539 VSS.n1481 VSS.n1354 0.00962857
R6540 VSS.n1477 VSS.n1354 0.00962857
R6541 VSS.n1477 VSS.n1356 0.00962857
R6542 VSS.n1473 VSS.n1356 0.00962857
R6543 VSS.n1473 VSS.n1358 0.00962857
R6544 VSS.n1469 VSS.n1358 0.00962857
R6545 VSS.n1469 VSS.n1360 0.00962857
R6546 VSS.n1465 VSS.n1360 0.00962857
R6547 VSS.n1465 VSS.n1362 0.00962857
R6548 VSS.n1461 VSS.n1362 0.00962857
R6549 VSS.n1461 VSS.n1364 0.00962857
R6550 VSS.n1457 VSS.n1364 0.00962857
R6551 VSS.n1457 VSS.n1366 0.00962857
R6552 VSS.n1453 VSS.n1366 0.00962857
R6553 VSS.n1453 VSS.n1368 0.00962857
R6554 VSS.n1449 VSS.n1368 0.00962857
R6555 VSS.n1449 VSS.n1370 0.00962857
R6556 VSS.n1445 VSS.n1370 0.00962857
R6557 VSS.n1445 VSS.n1372 0.00962857
R6558 VSS.n1441 VSS.n1372 0.00962857
R6559 VSS.n1441 VSS.n1374 0.00962857
R6560 VSS.n1437 VSS.n1374 0.00962857
R6561 VSS.n1437 VSS.n1376 0.00962857
R6562 VSS.n1433 VSS.n1376 0.00962857
R6563 VSS.n1433 VSS.n1378 0.00962857
R6564 VSS.n1429 VSS.n1378 0.00962857
R6565 VSS.n1429 VSS.n1380 0.00962857
R6566 VSS.n1425 VSS.n1380 0.00962857
R6567 VSS.n1425 VSS.n1382 0.00962857
R6568 VSS.n1421 VSS.n1382 0.00962857
R6569 VSS.n1421 VSS.n1384 0.00962857
R6570 VSS.n1417 VSS.n1384 0.00962857
R6571 VSS.n1417 VSS.n1386 0.00962857
R6572 VSS.n1413 VSS.n1386 0.00962857
R6573 VSS.n1413 VSS.n1388 0.00962857
R6574 VSS.n1409 VSS.n1388 0.00962857
R6575 VSS.n1409 VSS.n1390 0.00962857
R6576 VSS.n1405 VSS.n1390 0.00962857
R6577 VSS.n1405 VSS.n1392 0.00962857
R6578 VSS.n1401 VSS.n1392 0.00962857
R6579 VSS.n1401 VSS.n1394 0.00962857
R6580 VSS.n1586 VSS.n1299 0.00962857
R6581 VSS.n1580 VSS.n1299 0.00962857
R6582 VSS.n1580 VSS.n1579 0.00962857
R6583 VSS.n1579 VSS.n1578 0.00962857
R6584 VSS.n1578 VSS.n1305 0.00962857
R6585 VSS.n1572 VSS.n1305 0.00962857
R6586 VSS.n1572 VSS.n1571 0.00962857
R6587 VSS.n1571 VSS.n1570 0.00962857
R6588 VSS.n1570 VSS.n1309 0.00962857
R6589 VSS.n1564 VSS.n1309 0.00962857
R6590 VSS.n1564 VSS.n1563 0.00962857
R6591 VSS.n1563 VSS.n1562 0.00962857
R6592 VSS.n1562 VSS.n1313 0.00962857
R6593 VSS.n1556 VSS.n1313 0.00962857
R6594 VSS.n1556 VSS.n1555 0.00962857
R6595 VSS.n1555 VSS.n1554 0.00962857
R6596 VSS.n1554 VSS.n1317 0.00962857
R6597 VSS.n1548 VSS.n1317 0.00962857
R6598 VSS.n1548 VSS.n1547 0.00962857
R6599 VSS.n1547 VSS.n1546 0.00962857
R6600 VSS.n1546 VSS.n1321 0.00962857
R6601 VSS.n1540 VSS.n1321 0.00962857
R6602 VSS.n1540 VSS.n1539 0.00962857
R6603 VSS.n1539 VSS.n1538 0.00962857
R6604 VSS.n1538 VSS.n1325 0.00962857
R6605 VSS.n1532 VSS.n1325 0.00962857
R6606 VSS.n1532 VSS.n1531 0.00962857
R6607 VSS.n1531 VSS.n1530 0.00962857
R6608 VSS.n1530 VSS.n1329 0.00962857
R6609 VSS.n1524 VSS.n1329 0.00962857
R6610 VSS.n1524 VSS.n1523 0.00962857
R6611 VSS.n1523 VSS.n1522 0.00962857
R6612 VSS.n1522 VSS.n1333 0.00962857
R6613 VSS.n1516 VSS.n1333 0.00962857
R6614 VSS.n1516 VSS.n1515 0.00962857
R6615 VSS.n1515 VSS.n1514 0.00962857
R6616 VSS.n1514 VSS.n1337 0.00962857
R6617 VSS.n1508 VSS.n1337 0.00962857
R6618 VSS.n1508 VSS.n1507 0.00962857
R6619 VSS.n1507 VSS.n1506 0.00962857
R6620 VSS.n1506 VSS.n1341 0.00962857
R6621 VSS.n1500 VSS.n1341 0.00962857
R6622 VSS.n1500 VSS.n1499 0.00962857
R6623 VSS.n1499 VSS.n1498 0.00962857
R6624 VSS.n1498 VSS.n1345 0.00962857
R6625 VSS.n1492 VSS.n1345 0.00962857
R6626 VSS.n1492 VSS.n1491 0.00962857
R6627 VSS.n1491 VSS.n1490 0.00962857
R6628 VSS.n1490 VSS.n1349 0.00962857
R6629 VSS.n1484 VSS.n1349 0.00962857
R6630 VSS.n1484 VSS.n1483 0.00962857
R6631 VSS.n1483 VSS.n1482 0.00962857
R6632 VSS.n1482 VSS.n1353 0.00962857
R6633 VSS.n1476 VSS.n1353 0.00962857
R6634 VSS.n1476 VSS.n1475 0.00962857
R6635 VSS.n1475 VSS.n1474 0.00962857
R6636 VSS.n1474 VSS.n1357 0.00962857
R6637 VSS.n1468 VSS.n1357 0.00962857
R6638 VSS.n1468 VSS.n1467 0.00962857
R6639 VSS.n1467 VSS.n1466 0.00962857
R6640 VSS.n1466 VSS.n1361 0.00962857
R6641 VSS.n1460 VSS.n1361 0.00962857
R6642 VSS.n1460 VSS.n1459 0.00962857
R6643 VSS.n1459 VSS.n1458 0.00962857
R6644 VSS.n1458 VSS.n1365 0.00962857
R6645 VSS.n1452 VSS.n1365 0.00962857
R6646 VSS.n1452 VSS.n1451 0.00962857
R6647 VSS.n1451 VSS.n1450 0.00962857
R6648 VSS.n1450 VSS.n1369 0.00962857
R6649 VSS.n1444 VSS.n1369 0.00962857
R6650 VSS.n1444 VSS.n1443 0.00962857
R6651 VSS.n1443 VSS.n1442 0.00962857
R6652 VSS.n1442 VSS.n1373 0.00962857
R6653 VSS.n1436 VSS.n1373 0.00962857
R6654 VSS.n1436 VSS.n1435 0.00962857
R6655 VSS.n1435 VSS.n1434 0.00962857
R6656 VSS.n1434 VSS.n1377 0.00962857
R6657 VSS.n1428 VSS.n1377 0.00962857
R6658 VSS.n1428 VSS.n1427 0.00962857
R6659 VSS.n1427 VSS.n1426 0.00962857
R6660 VSS.n1426 VSS.n1381 0.00962857
R6661 VSS.n1420 VSS.n1381 0.00962857
R6662 VSS.n1420 VSS.n1419 0.00962857
R6663 VSS.n1419 VSS.n1418 0.00962857
R6664 VSS.n1418 VSS.n1385 0.00962857
R6665 VSS.n1412 VSS.n1385 0.00962857
R6666 VSS.n1412 VSS.n1411 0.00962857
R6667 VSS.n1411 VSS.n1410 0.00962857
R6668 VSS.n1410 VSS.n1389 0.00962857
R6669 VSS.n1404 VSS.n1389 0.00962857
R6670 VSS.n1404 VSS.n1403 0.00962857
R6671 VSS.n1403 VSS.n1402 0.00962857
R6672 VSS.n1402 VSS.n1393 0.00962857
R6673 VSS.n4190 VSS.n2639 0.00962857
R6674 VSS.n4183 VSS.n2643 0.00962857
R6675 VSS.n4183 VSS.n4182 0.00962857
R6676 VSS.n4182 VSS.n4181 0.00962857
R6677 VSS.n4142 VSS.n3762 0.00962857
R6678 VSS.n4136 VSS.n3762 0.00962857
R6679 VSS.n4056 VSS.n4055 0.00962857
R6680 VSS.n4055 VSS.n3966 0.00962857
R6681 VSS.n4049 VSS.n3966 0.00962857
R6682 VSS.n4049 VSS.n4048 0.00962857
R6683 VSS.n4048 VSS.n4047 0.00962857
R6684 VSS.n4047 VSS.n3970 0.00962857
R6685 VSS.n4041 VSS.n3970 0.00962857
R6686 VSS.n4041 VSS.n4040 0.00962857
R6687 VSS.n4040 VSS.n4039 0.00962857
R6688 VSS.n4039 VSS.n3974 0.00962857
R6689 VSS.n4033 VSS.n3974 0.00962857
R6690 VSS.n4033 VSS.n4032 0.00962857
R6691 VSS.n4032 VSS.n4031 0.00962857
R6692 VSS.n4031 VSS.n3978 0.00962857
R6693 VSS.n4025 VSS.n3978 0.00962857
R6694 VSS.n4025 VSS.n4024 0.00962857
R6695 VSS.n4024 VSS.n4023 0.00962857
R6696 VSS.n4023 VSS.n3982 0.00962857
R6697 VSS.n4017 VSS.n3982 0.00962857
R6698 VSS.n4017 VSS.n4016 0.00962857
R6699 VSS.n4016 VSS.n4015 0.00962857
R6700 VSS.n4015 VSS.n3986 0.00962857
R6701 VSS.n4009 VSS.n3986 0.00962857
R6702 VSS.n4009 VSS.n4008 0.00962857
R6703 VSS.n4008 VSS.n4007 0.00962857
R6704 VSS.n4007 VSS.n3990 0.00962857
R6705 VSS.n4001 VSS.n3990 0.00962857
R6706 VSS.n4001 VSS.n4000 0.00962857
R6707 VSS.n4000 VSS.n3999 0.00962857
R6708 VSS.n3540 VSS.n3536 0.00962857
R6709 VSS.n3559 VSS.n3536 0.00962857
R6710 VSS.n3559 VSS.n3537 0.00962857
R6711 VSS.n3555 VSS.n3537 0.00962857
R6712 VSS.n3555 VSS.n3544 0.00962857
R6713 VSS.n3550 VSS.n3544 0.00962857
R6714 VSS.n3550 VSS.n3547 0.00962857
R6715 VSS.n3547 VSS.n2722 0.00962857
R6716 VSS.n3570 VSS.n2722 0.00962857
R6717 VSS.n3570 VSS.n2720 0.00962857
R6718 VSS.n3574 VSS.n2720 0.00962857
R6719 VSS.n3574 VSS.n2718 0.00962857
R6720 VSS.n3579 VSS.n2718 0.00962857
R6721 VSS.n3579 VSS.n2716 0.00962857
R6722 VSS.n3583 VSS.n2716 0.00962857
R6723 VSS.n3583 VSS.n2714 0.00962857
R6724 VSS.n3589 VSS.n2714 0.00962857
R6725 VSS.n3589 VSS.n2711 0.00962857
R6726 VSS.n3597 VSS.n2711 0.00962857
R6727 VSS.n3597 VSS.n2712 0.00962857
R6728 VSS.n3593 VSS.n2712 0.00962857
R6729 VSS.n3593 VSS.n2674 0.00962857
R6730 VSS.n3713 VSS.n2674 0.00962857
R6731 VSS.n3713 VSS.n2675 0.00962857
R6732 VSS.n3709 VSS.n2675 0.00962857
R6733 VSS.n3709 VSS.n3708 0.00962857
R6734 VSS.n3708 VSS.n2678 0.00962857
R6735 VSS.n3704 VSS.n2678 0.00962857
R6736 VSS.n3704 VSS.n2680 0.00962857
R6737 VSS.n3700 VSS.n2680 0.00962857
R6738 VSS.n3700 VSS.n2683 0.00962857
R6739 VSS.n3696 VSS.n2683 0.00962857
R6740 VSS.n3696 VSS.n2685 0.00962857
R6741 VSS.n3692 VSS.n2685 0.00962857
R6742 VSS.n3692 VSS.n2687 0.00962857
R6743 VSS.n3688 VSS.n2687 0.00962857
R6744 VSS.n3688 VSS.n2689 0.00962857
R6745 VSS.n3684 VSS.n2689 0.00962857
R6746 VSS.n3684 VSS.n2691 0.00962857
R6747 VSS.n3636 VSS.n2691 0.00962857
R6748 VSS.n3636 VSS.n3634 0.00962857
R6749 VSS.n3643 VSS.n3634 0.00962857
R6750 VSS.n3643 VSS.n3632 0.00962857
R6751 VSS.n3647 VSS.n3632 0.00962857
R6752 VSS.n3647 VSS.n3630 0.00962857
R6753 VSS.n3653 VSS.n3630 0.00962857
R6754 VSS.n3653 VSS.n3627 0.00962857
R6755 VSS.n3671 VSS.n3627 0.00962857
R6756 VSS.n3671 VSS.n3628 0.00962857
R6757 VSS.n3667 VSS.n3628 0.00962857
R6758 VSS.n3667 VSS.n3657 0.00962857
R6759 VSS.n3662 VSS.n3657 0.00962857
R6760 VSS.n3662 VSS.n3659 0.00962857
R6761 VSS.n3659 VSS.n2245 0.00962857
R6762 VSS.n5248 VSS.n2245 0.00962857
R6763 VSS.n5248 VSS.n2246 0.00962857
R6764 VSS.n5244 VSS.n2246 0.00962857
R6765 VSS.n5244 VSS.n2249 0.00962857
R6766 VSS.n5240 VSS.n2249 0.00962857
R6767 VSS.n5240 VSS.n2252 0.00962857
R6768 VSS.n5236 VSS.n2252 0.00962857
R6769 VSS.n5236 VSS.n2254 0.00962857
R6770 VSS.n5232 VSS.n2254 0.00962857
R6771 VSS.n5232 VSS.n2256 0.00962857
R6772 VSS.n5228 VSS.n2256 0.00962857
R6773 VSS.n5228 VSS.n2258 0.00962857
R6774 VSS.n5224 VSS.n2258 0.00962857
R6775 VSS.n5224 VSS.n2260 0.00962857
R6776 VSS.n5220 VSS.n2260 0.00962857
R6777 VSS.n5220 VSS.n2262 0.00962857
R6778 VSS.n5216 VSS.n2262 0.00962857
R6779 VSS.n5216 VSS.n2264 0.00962857
R6780 VSS.n5212 VSS.n2264 0.00962857
R6781 VSS.n5212 VSS.n2266 0.00962857
R6782 VSS.n5208 VSS.n2266 0.00962857
R6783 VSS.n5208 VSS.n2268 0.00962857
R6784 VSS.n5204 VSS.n2268 0.00962857
R6785 VSS.n5204 VSS.n2270 0.00962857
R6786 VSS.n5200 VSS.n2270 0.00962857
R6787 VSS.n5200 VSS.n5185 0.00962857
R6788 VSS.n5196 VSS.n5185 0.00962857
R6789 VSS.n5196 VSS.n5187 0.00962857
R6790 VSS.n5192 VSS.n5187 0.00962857
R6791 VSS.n3539 VSS.n3534 0.00962857
R6792 VSS.n3560 VSS.n3535 0.00962857
R6793 VSS.n3554 VSS.n3535 0.00962857
R6794 VSS.n3552 VSS.n3551 0.00962857
R6795 VSS.n3551 VSS.n3546 0.00962857
R6796 VSS.n3546 VSS.n3545 0.00962857
R6797 VSS.n3576 VSS.n3575 0.00962857
R6798 VSS.n3578 VSS.n3576 0.00962857
R6799 VSS.n3578 VSS.n3577 0.00962857
R6800 VSS.n3585 VSS.n3584 0.00962857
R6801 VSS.n3588 VSS.n3585 0.00962857
R6802 VSS.n3598 VSS.n2710 0.00962857
R6803 VSS.n3592 VSS.n2710 0.00962857
R6804 VSS.n3592 VSS.n2670 0.00962857
R6805 VSS.n3707 VSS.n2661 0.00962857
R6806 VSS.n3707 VSS.n3706 0.00962857
R6807 VSS.n3706 VSS.n3705 0.00962857
R6808 VSS.n3705 VSS.n2679 0.00962857
R6809 VSS.n3699 VSS.n2679 0.00962857
R6810 VSS.n3699 VSS.n3698 0.00962857
R6811 VSS.n3698 VSS.n3697 0.00962857
R6812 VSS.n3697 VSS.n2684 0.00962857
R6813 VSS.n3691 VSS.n2684 0.00962857
R6814 VSS.n3691 VSS.n3690 0.00962857
R6815 VSS.n3690 VSS.n3689 0.00962857
R6816 VSS.n3683 VSS.n2692 0.00962857
R6817 VSS.n3637 VSS.n2693 0.00962857
R6818 VSS.n3638 VSS.n3637 0.00962857
R6819 VSS.n3642 VSS.n3631 0.00962857
R6820 VSS.n3648 VSS.n3631 0.00962857
R6821 VSS.n3649 VSS.n3648 0.00962857
R6822 VSS.n3672 VSS.n3626 0.00962857
R6823 VSS.n3666 VSS.n3626 0.00962857
R6824 VSS.n3666 VSS.n3665 0.00962857
R6825 VSS.n3663 VSS.n3658 0.00962857
R6826 VSS.n3658 VSS.n2243 0.00962857
R6827 VSS.n5243 VSS.n2250 0.00962857
R6828 VSS.n5243 VSS.n5242 0.00962857
R6829 VSS.n5242 VSS.n5241 0.00962857
R6830 VSS.n5241 VSS.n2251 0.00962857
R6831 VSS.n5235 VSS.n2251 0.00962857
R6832 VSS.n5235 VSS.n5234 0.00962857
R6833 VSS.n5234 VSS.n5233 0.00962857
R6834 VSS.n5233 VSS.n2255 0.00962857
R6835 VSS.n5227 VSS.n2255 0.00962857
R6836 VSS.n5227 VSS.n5226 0.00962857
R6837 VSS.n5226 VSS.n5225 0.00962857
R6838 VSS.n5225 VSS.n2259 0.00962857
R6839 VSS.n5219 VSS.n2259 0.00962857
R6840 VSS.n5219 VSS.n5218 0.00962857
R6841 VSS.n5218 VSS.n5217 0.00962857
R6842 VSS.n5217 VSS.n2263 0.00962857
R6843 VSS.n5211 VSS.n2263 0.00962857
R6844 VSS.n5211 VSS.n5210 0.00962857
R6845 VSS.n5210 VSS.n5209 0.00962857
R6846 VSS.n5209 VSS.n2267 0.00962857
R6847 VSS.n5203 VSS.n5202 0.00962857
R6848 VSS.n5202 VSS.n5201 0.00962857
R6849 VSS.n5201 VSS.n5184 0.00962857
R6850 VSS.n5195 VSS.n5184 0.00962857
R6851 VSS.n5195 VSS.n5194 0.00962857
R6852 VSS.n5194 VSS.n5193 0.00962857
R6853 VSS.n2767 VSS.n2766 0.00962857
R6854 VSS.n2768 VSS.n2767 0.00962857
R6855 VSS.n2768 VSS.n2760 0.00962857
R6856 VSS.n2774 VSS.n2760 0.00962857
R6857 VSS.n2775 VSS.n2774 0.00962857
R6858 VSS.n2776 VSS.n2775 0.00962857
R6859 VSS.n2776 VSS.n2756 0.00962857
R6860 VSS.n2782 VSS.n2756 0.00962857
R6861 VSS.n2783 VSS.n2782 0.00962857
R6862 VSS.n2784 VSS.n2783 0.00962857
R6863 VSS.n2784 VSS.n2752 0.00962857
R6864 VSS.n2790 VSS.n2752 0.00962857
R6865 VSS.n3263 VSS.n3262 0.00962857
R6866 VSS.n3263 VSS.n2748 0.00962857
R6867 VSS.n3269 VSS.n2748 0.00962857
R6868 VSS.n3270 VSS.n3269 0.00962857
R6869 VSS.n3271 VSS.n3270 0.00962857
R6870 VSS.n3271 VSS.n2744 0.00962857
R6871 VSS.n3277 VSS.n2744 0.00962857
R6872 VSS.n3278 VSS.n3277 0.00962857
R6873 VSS.n3279 VSS.n3278 0.00962857
R6874 VSS.n3279 VSS.n2740 0.00962857
R6875 VSS.n3285 VSS.n2740 0.00962857
R6876 VSS.n3286 VSS.n3285 0.00962857
R6877 VSS.n3287 VSS.n3286 0.00962857
R6878 VSS.n3287 VSS.n2734 0.00962857
R6879 VSS.n3516 VSS.n2735 0.00962857
R6880 VSS.n3510 VSS.n2735 0.00962857
R6881 VSS.n3510 VSS.n3509 0.00962857
R6882 VSS.n3509 VSS.n3508 0.00962857
R6883 VSS.n3508 VSS.n3293 0.00962857
R6884 VSS.n3502 VSS.n3293 0.00962857
R6885 VSS.n3502 VSS.n3501 0.00962857
R6886 VSS.n3501 VSS.n3500 0.00962857
R6887 VSS.n3500 VSS.n3297 0.00962857
R6888 VSS.n3494 VSS.n3297 0.00962857
R6889 VSS.n3494 VSS.n3493 0.00962857
R6890 VSS.n3493 VSS.n3492 0.00962857
R6891 VSS.n3492 VSS.n3301 0.00962857
R6892 VSS.n3486 VSS.n3301 0.00962857
R6893 VSS.n3486 VSS.n3485 0.00962857
R6894 VSS.n3485 VSS.n3484 0.00962857
R6895 VSS.n3484 VSS.n3305 0.00962857
R6896 VSS.n3478 VSS.n3305 0.00962857
R6897 VSS.n3478 VSS.n3477 0.00962857
R6898 VSS.n3477 VSS.n3476 0.00962857
R6899 VSS.n3476 VSS.n3309 0.00962857
R6900 VSS.n3470 VSS.n3309 0.00962857
R6901 VSS.n3470 VSS.n3469 0.00962857
R6902 VSS.n3469 VSS.n3468 0.00962857
R6903 VSS.n3468 VSS.n3313 0.00962857
R6904 VSS.n3462 VSS.n3313 0.00962857
R6905 VSS.n3462 VSS.n3461 0.00962857
R6906 VSS.n3461 VSS.n3460 0.00962857
R6907 VSS.n3460 VSS.n3317 0.00962857
R6908 VSS.n3454 VSS.n3317 0.00962857
R6909 VSS.n3454 VSS.n3453 0.00962857
R6910 VSS.n3453 VSS.n3452 0.00962857
R6911 VSS.n3452 VSS.n3321 0.00962857
R6912 VSS.n3446 VSS.n3321 0.00962857
R6913 VSS.n3446 VSS.n3445 0.00962857
R6914 VSS.n3445 VSS.n3444 0.00962857
R6915 VSS.n3444 VSS.n3325 0.00962857
R6916 VSS.n3438 VSS.n3325 0.00962857
R6917 VSS.n3438 VSS.n3437 0.00962857
R6918 VSS.n3437 VSS.n3436 0.00962857
R6919 VSS.n3436 VSS.n3329 0.00962857
R6920 VSS.n3430 VSS.n3329 0.00962857
R6921 VSS.n3430 VSS.n3429 0.00962857
R6922 VSS.n3429 VSS.n3428 0.00962857
R6923 VSS.n3428 VSS.n3333 0.00962857
R6924 VSS.n3422 VSS.n3333 0.00962857
R6925 VSS.n3422 VSS.n3421 0.00962857
R6926 VSS.n3421 VSS.n3420 0.00962857
R6927 VSS.n3420 VSS.n3337 0.00962857
R6928 VSS.n3414 VSS.n3337 0.00962857
R6929 VSS.n3414 VSS.n3413 0.00962857
R6930 VSS.n3413 VSS.n3412 0.00962857
R6931 VSS.n3412 VSS.n3341 0.00962857
R6932 VSS.n3406 VSS.n3341 0.00962857
R6933 VSS.n3406 VSS.n3405 0.00962857
R6934 VSS.n3405 VSS.n3404 0.00962857
R6935 VSS.n3404 VSS.n3345 0.00962857
R6936 VSS.n3398 VSS.n3345 0.00962857
R6937 VSS.n3398 VSS.n3397 0.00962857
R6938 VSS.n3397 VSS.n3396 0.00962857
R6939 VSS.n3396 VSS.n3349 0.00962857
R6940 VSS.n3390 VSS.n3349 0.00962857
R6941 VSS.n3390 VSS.n3389 0.00962857
R6942 VSS.n3389 VSS.n3388 0.00962857
R6943 VSS.n3388 VSS.n3353 0.00962857
R6944 VSS.n3382 VSS.n3353 0.00962857
R6945 VSS.n3382 VSS.n3381 0.00962857
R6946 VSS.n3381 VSS.n3380 0.00962857
R6947 VSS.n3380 VSS.n2417 0.00962857
R6948 VSS.n3367 VSS.n3366 0.00962857
R6949 VSS.n3366 VSS.n3365 0.00962857
R6950 VSS.n3365 VSS.n3361 0.00962857
R6951 VSS.n4240 VSS.n4237 0.00962857
R6952 VSS.n4241 VSS.n4240 0.00962857
R6953 VSS.n4242 VSS.n4241 0.00962857
R6954 VSS.n4242 VSS.n4233 0.00962857
R6955 VSS.n4248 VSS.n4233 0.00962857
R6956 VSS.n4249 VSS.n4248 0.00962857
R6957 VSS.n4250 VSS.n4249 0.00962857
R6958 VSS.n4250 VSS.n4229 0.00962857
R6959 VSS.n4256 VSS.n4229 0.00962857
R6960 VSS.n4257 VSS.n4256 0.00962857
R6961 VSS.n4258 VSS.n4257 0.00962857
R6962 VSS.n4258 VSS.n4225 0.00962857
R6963 VSS.n4264 VSS.n4225 0.00962857
R6964 VSS.n4265 VSS.n4264 0.00962857
R6965 VSS.n4266 VSS.n4265 0.00962857
R6966 VSS.n4300 VSS.n4220 0.00962857
R6967 VSS.n4294 VSS.n4220 0.00962857
R6968 VSS.n4294 VSS.n4293 0.00962857
R6969 VSS.n4293 VSS.n4292 0.00962857
R6970 VSS.n4292 VSS.n4272 0.00962857
R6971 VSS.n4286 VSS.n4272 0.00962857
R6972 VSS.n4687 VSS.n2496 0.00962857
R6973 VSS.n4693 VSS.n2496 0.00962857
R6974 VSS.n4694 VSS.n4693 0.00962857
R6975 VSS.n4695 VSS.n4694 0.00962857
R6976 VSS.n4695 VSS.n2492 0.00962857
R6977 VSS.n4701 VSS.n2492 0.00962857
R6978 VSS.n4702 VSS.n4701 0.00962857
R6979 VSS.n4703 VSS.n4702 0.00962857
R6980 VSS.n4703 VSS.n2488 0.00962857
R6981 VSS.n4709 VSS.n2488 0.00962857
R6982 VSS.n4710 VSS.n4709 0.00962857
R6983 VSS.n4711 VSS.n4710 0.00962857
R6984 VSS.n4711 VSS.n2484 0.00962857
R6985 VSS.n4717 VSS.n2484 0.00962857
R6986 VSS.n4718 VSS.n4717 0.00962857
R6987 VSS.n4719 VSS.n4718 0.00962857
R6988 VSS.n4719 VSS.n2480 0.00962857
R6989 VSS.n4725 VSS.n2480 0.00962857
R6990 VSS.n4726 VSS.n4725 0.00962857
R6991 VSS.n4727 VSS.n4726 0.00962857
R6992 VSS.n4727 VSS.n2476 0.00962857
R6993 VSS.n4733 VSS.n2476 0.00962857
R6994 VSS.n4734 VSS.n4733 0.00962857
R6995 VSS.n4735 VSS.n4734 0.00962857
R6996 VSS.n4735 VSS.n2472 0.00962857
R6997 VSS.n4741 VSS.n2472 0.00962857
R6998 VSS.n4742 VSS.n4741 0.00962857
R6999 VSS.n4743 VSS.n4742 0.00962857
R7000 VSS.n4743 VSS.n2468 0.00962857
R7001 VSS.n4749 VSS.n2468 0.00962857
R7002 VSS.n4752 VSS.n4751 0.00962857
R7003 VSS.n4752 VSS.n2464 0.00962857
R7004 VSS.n4758 VSS.n2464 0.00962857
R7005 VSS.n4759 VSS.n4758 0.00962857
R7006 VSS.n4760 VSS.n4759 0.00962857
R7007 VSS.n4760 VSS.n2460 0.00962857
R7008 VSS.n4766 VSS.n2460 0.00962857
R7009 VSS.n4767 VSS.n4766 0.00962857
R7010 VSS.n4768 VSS.n4767 0.00962857
R7011 VSS.n4768 VSS.n2456 0.00962857
R7012 VSS.n4774 VSS.n2456 0.00962857
R7013 VSS.n4775 VSS.n4774 0.00962857
R7014 VSS.n4776 VSS.n4775 0.00962857
R7015 VSS.n4776 VSS.n2452 0.00962857
R7016 VSS.n4782 VSS.n2452 0.00962857
R7017 VSS.n4783 VSS.n4782 0.00962857
R7018 VSS.n4784 VSS.n4783 0.00962857
R7019 VSS.n4784 VSS.n2448 0.00962857
R7020 VSS.n4790 VSS.n2448 0.00962857
R7021 VSS.n4791 VSS.n4790 0.00962857
R7022 VSS.n4792 VSS.n4791 0.00962857
R7023 VSS.n4792 VSS.n2444 0.00962857
R7024 VSS.n4798 VSS.n2444 0.00962857
R7025 VSS.n4799 VSS.n4798 0.00962857
R7026 VSS.n4800 VSS.n4799 0.00962857
R7027 VSS.n4800 VSS.n2440 0.00962857
R7028 VSS.n4806 VSS.n2440 0.00962857
R7029 VSS.n4807 VSS.n4806 0.00962857
R7030 VSS.n4808 VSS.n4807 0.00962857
R7031 VSS.n4808 VSS.n2436 0.00962857
R7032 VSS.n4814 VSS.n2436 0.00962857
R7033 VSS.n4815 VSS.n4814 0.00962857
R7034 VSS.n4817 VSS.n4815 0.00962857
R7035 VSS.n4817 VSS.n4816 0.00962857
R7036 VSS.n4816 VSS.n2432 0.00962857
R7037 VSS.n5717 VSS.n6 0.00962857
R7038 VSS.n5717 VSS.n5716 0.00962857
R7039 VSS.n5716 VSS.n5715 0.00962857
R7040 VSS.n4239 VSS.n4236 0.00962857
R7041 VSS.n4243 VSS.n4236 0.00962857
R7042 VSS.n4243 VSS.n4234 0.00962857
R7043 VSS.n4247 VSS.n4234 0.00962857
R7044 VSS.n4247 VSS.n4232 0.00962857
R7045 VSS.n4251 VSS.n4232 0.00962857
R7046 VSS.n4251 VSS.n4230 0.00962857
R7047 VSS.n4255 VSS.n4230 0.00962857
R7048 VSS.n4255 VSS.n4228 0.00962857
R7049 VSS.n4259 VSS.n4228 0.00962857
R7050 VSS.n4259 VSS.n4226 0.00962857
R7051 VSS.n4263 VSS.n4226 0.00962857
R7052 VSS.n4263 VSS.n4224 0.00962857
R7053 VSS.n4267 VSS.n4224 0.00962857
R7054 VSS.n4267 VSS.n4221 0.00962857
R7055 VSS.n4299 VSS.n4221 0.00962857
R7056 VSS.n4299 VSS.n4222 0.00962857
R7057 VSS.n4295 VSS.n4222 0.00962857
R7058 VSS.n4295 VSS.n4271 0.00962857
R7059 VSS.n4291 VSS.n4271 0.00962857
R7060 VSS.n4291 VSS.n4273 0.00962857
R7061 VSS.n4287 VSS.n4273 0.00962857
R7062 VSS.n4287 VSS.n4275 0.00962857
R7063 VSS.n4281 VSS.n4275 0.00962857
R7064 VSS.n4281 VSS.n2505 0.00962857
R7065 VSS.n4678 VSS.n2505 0.00962857
R7066 VSS.n4678 VSS.n2503 0.00962857
R7067 VSS.n4682 VSS.n2503 0.00962857
R7068 VSS.n4682 VSS.n2499 0.00962857
R7069 VSS.n4688 VSS.n2499 0.00962857
R7070 VSS.n4688 VSS.n2497 0.00962857
R7071 VSS.n4692 VSS.n2497 0.00962857
R7072 VSS.n4692 VSS.n2495 0.00962857
R7073 VSS.n4696 VSS.n2495 0.00962857
R7074 VSS.n4696 VSS.n2493 0.00962857
R7075 VSS.n4700 VSS.n2493 0.00962857
R7076 VSS.n4700 VSS.n2491 0.00962857
R7077 VSS.n4704 VSS.n2491 0.00962857
R7078 VSS.n4704 VSS.n2489 0.00962857
R7079 VSS.n4708 VSS.n2489 0.00962857
R7080 VSS.n4708 VSS.n2487 0.00962857
R7081 VSS.n4712 VSS.n2487 0.00962857
R7082 VSS.n4712 VSS.n2485 0.00962857
R7083 VSS.n4716 VSS.n2485 0.00962857
R7084 VSS.n4716 VSS.n2483 0.00962857
R7085 VSS.n4720 VSS.n2483 0.00962857
R7086 VSS.n4720 VSS.n2481 0.00962857
R7087 VSS.n4724 VSS.n2481 0.00962857
R7088 VSS.n4724 VSS.n2479 0.00962857
R7089 VSS.n4728 VSS.n2479 0.00962857
R7090 VSS.n4728 VSS.n2477 0.00962857
R7091 VSS.n4732 VSS.n2477 0.00962857
R7092 VSS.n4732 VSS.n2475 0.00962857
R7093 VSS.n4736 VSS.n2475 0.00962857
R7094 VSS.n4736 VSS.n2473 0.00962857
R7095 VSS.n4740 VSS.n2473 0.00962857
R7096 VSS.n4740 VSS.n2471 0.00962857
R7097 VSS.n4744 VSS.n2471 0.00962857
R7098 VSS.n4744 VSS.n2469 0.00962857
R7099 VSS.n4748 VSS.n2469 0.00962857
R7100 VSS.n4748 VSS.n2467 0.00962857
R7101 VSS.n4753 VSS.n2467 0.00962857
R7102 VSS.n4753 VSS.n2465 0.00962857
R7103 VSS.n4757 VSS.n2465 0.00962857
R7104 VSS.n4757 VSS.n2463 0.00962857
R7105 VSS.n4761 VSS.n2463 0.00962857
R7106 VSS.n4761 VSS.n2461 0.00962857
R7107 VSS.n4765 VSS.n2461 0.00962857
R7108 VSS.n4765 VSS.n2459 0.00962857
R7109 VSS.n4769 VSS.n2459 0.00962857
R7110 VSS.n4769 VSS.n2457 0.00962857
R7111 VSS.n4773 VSS.n2457 0.00962857
R7112 VSS.n4773 VSS.n2455 0.00962857
R7113 VSS.n4777 VSS.n2455 0.00962857
R7114 VSS.n4777 VSS.n2453 0.00962857
R7115 VSS.n4781 VSS.n2453 0.00962857
R7116 VSS.n4781 VSS.n2451 0.00962857
R7117 VSS.n4785 VSS.n2451 0.00962857
R7118 VSS.n4785 VSS.n2449 0.00962857
R7119 VSS.n4789 VSS.n2449 0.00962857
R7120 VSS.n4789 VSS.n2447 0.00962857
R7121 VSS.n4793 VSS.n2447 0.00962857
R7122 VSS.n4793 VSS.n2445 0.00962857
R7123 VSS.n4797 VSS.n2445 0.00962857
R7124 VSS.n4797 VSS.n2443 0.00962857
R7125 VSS.n4801 VSS.n2443 0.00962857
R7126 VSS.n4801 VSS.n2441 0.00962857
R7127 VSS.n4805 VSS.n2441 0.00962857
R7128 VSS.n4805 VSS.n2439 0.00962857
R7129 VSS.n4809 VSS.n2439 0.00962857
R7130 VSS.n4809 VSS.n2437 0.00962857
R7131 VSS.n4813 VSS.n2437 0.00962857
R7132 VSS.n4813 VSS.n2435 0.00962857
R7133 VSS.n4818 VSS.n2435 0.00962857
R7134 VSS.n4818 VSS.n2433 0.00962857
R7135 VSS.n4822 VSS.n2433 0.00962857
R7136 VSS.n4823 VSS.n4822 0.00962857
R7137 VSS.n5722 VSS.n2 0.00962857
R7138 VSS.n5718 VSS.n2 0.00962857
R7139 VSS.n5718 VSS.n5 0.00962857
R7140 VSS.n5109 DVSS 0.00958867
R7141 DVSS VSS.n2285 0.00958867
R7142 VSS.n3950 VSS.n3946 0.00958257
R7143 VSS.n4165 VSS.n3725 0.00958257
R7144 VSS.n5203 VSS.n5183 0.00956429
R7145 VSS.n911 VSS.n218 0.0095301
R7146 VSS.n4174 VSS.n2649 0.0095
R7147 VSS.n3798 VSS.n3797 0.0095
R7148 VSS.n3804 VSS.n3803 0.0095
R7149 VSS.n3796 VSS.n3794 0.0095
R7150 VSS.n3807 VSS.n3806 0.0095
R7151 VSS.n4162 VSS.n4160 0.0095
R7152 VSS.n3741 VSS.n3735 0.0095
R7153 VSS.n4154 VSS.n3742 0.0095
R7154 VSS.n4153 VSS.n3743 0.0095
R7155 VSS.n4144 VSS.n4142 0.0095
R7156 VSS.n3932 VSS.n3924 0.0095
R7157 VSS.n3931 VSS.n3911 0.0095
R7158 VSS.n3940 VSS.n3939 0.0095
R7159 VSS.n3914 VSS.n3912 0.0095
R7160 VSS.n4107 VSS.n3900 0.0095
R7161 VSS.n4106 VSS.n3901 0.0095
R7162 VSS.n3957 VSS.n3956 0.0095
R7163 VSS.n4098 VSS.n4097 0.0095
R7164 VSS.n4087 VSS.n3958 0.0095
R7165 VSS.n2977 VSS.n2905 0.0095
R7166 VSS.n3019 VSS.n2896 0.0095
R7167 VSS.n5072 VSS.n2311 0.0095
R7168 VSS.n5097 VSS.n5095 0.0095
R7169 VSS.n2963 VSS.n2913 0.0095
R7170 VSS.n3016 VSS.n2898 0.0095
R7171 VSS.n5058 VSS.n2316 0.0095
R7172 VSS.n5099 VSS.n2296 0.0095
R7173 VSS.n5694 VSS.n5693 0.00934354
R7174 VSS.n5693 VSS.n5692 0.00934354
R7175 VSS.n2076 VSS.n2075 0.00933782
R7176 VSS.n2069 VSS.n1594 0.00933782
R7177 VSS.n2075 VSS.n1594 0.00933782
R7178 VSS.n2073 VSS.n2069 0.00933782
R7179 VSS.n1809 VSS.n16 0.00933782
R7180 VSS.n1811 VSS.n1809 0.00933782
R7181 VSS.n1880 VSS.n1879 0.00928049
R7182 VSS.n1875 VSS.n1874 0.00928049
R7183 VSS.n1914 VSS.n1727 0.00928049
R7184 VSS.n1900 VSS.n1747 0.00928049
R7185 VSS.n1952 VSS.n1703 0.00928049
R7186 VSS.n1938 VSS.n1705 0.00928049
R7187 VSS.n1738 VSS.n1736 0.00928049
R7188 VSS.n1977 VSS.n1685 0.00928049
R7189 VSS.n1732 VSS.n1730 0.00928049
R7190 VSS.n2009 VSS.n1660 0.00928049
R7191 VSS.n2045 VSS.n2044 0.00928049
R7192 VSS.n2040 VSS.n2039 0.00928049
R7193 VSS.n1396 VSS.n33 0.00924286
R7194 VSS.n5451 VSS.n5450 0.00910927
R7195 VSS.n5713 VSS.n5712 0.00910927
R7196 VSS.n636 VSS.n635 0.00909873
R7197 VSS.n2954 VSS.n2953 0.009
R7198 VSS.n3043 VSS.n3042 0.009
R7199 VSS.n5042 VSS.n2320 0.009
R7200 VSS.n5115 VSS.n5114 0.009
R7201 VSS.n2957 VSS.n2956 0.009
R7202 VSS.n3008 VSS.n2887 0.009
R7203 VSS.n2324 VSS.n2318 0.009
R7204 VSS.n5119 VSS.n5117 0.009
R7205 VSS.n3851 VSS.n2559 0.00894122
R7206 VSS.n3851 VSS.n2565 0.00894122
R7207 VSS.n3652 VSS.n3650 0.00892143
R7208 VSS.n3664 VSS.n3663 0.00892143
R7209 VSS.n4266 VSS.n4218 0.00892143
R7210 VSS.n4301 VSS.n4219 0.00892143
R7211 VSS.n217 VSS.n172 0.00882776
R7212 VSS.n4239 VSS.n4238 0.00880017
R7213 VSS.n4440 VSS.n4439 0.00879286
R7214 VSS.n2614 VSS.n2609 0.00879286
R7215 VSS.n4437 VSS.n4348 0.00879286
R7216 VSS.n3599 VSS.n2709 0.00879286
R7217 VSS.n4181 VSS.n2644 0.0086
R7218 VSS.n4515 VSS.n2556 0.00853571
R7219 VSS.n4514 VSS.n2562 0.00853571
R7220 VSS.n4512 VSS.n4511 0.00853571
R7221 VSS.n1920 VSS.n1724 0.00853571
R7222 VSS.n1919 VSS.n1725 0.00853571
R7223 VSS.n1749 VSS.n1748 0.00853571
R7224 VSS.n1912 VSS.n1911 0.00853571
R7225 VSS.n1756 VSS.n1750 0.00853571
R7226 VSS.n1905 VSS.n1757 0.00853571
R7227 VSS.n1904 VSS.n1897 0.00853571
R7228 VSS.n3689 VSS.n2688 0.00853571
R7229 VSS.n5151 DVSS 0.00852817
R7230 VSS.n5152 DVSS 0.00852817
R7231 VSS.n3096 VSS.n3095 0.0085
R7232 VSS.n4998 VSS.n2343 0.0085
R7233 VSS.n3069 VSS.n2864 0.0085
R7234 VSS.n4978 VSS.n2346 0.0085
R7235 VSS.n1830 VSS.n20 0.00847143
R7236 VSS.n3827 VSS.n2648 0.00847143
R7237 VSS.n4286 VSS.n4285 0.00847143
R7238 VSS.n4283 VSS.n4276 0.00847143
R7239 VSS.n4282 VSS.n4279 0.00847143
R7240 VSS.n4278 VSS.n2506 0.00847143
R7241 VSS.n4677 VSS.n4676 0.00847143
R7242 VSS.n2507 VSS.n2502 0.00847143
R7243 VSS.n4684 VSS.n4683 0.00847143
R7244 VSS.n4686 VSS.n2500 0.00847143
R7245 VSS.n537 VSS.n365 0.00842994
R7246 VSS.n4091 VSS.n3964 0.00834286
R7247 VSS.n4057 VSS.n4056 0.00834286
R7248 VSS.n3569 VSS.n2723 0.00827857
R7249 VSS.n3584 VSS.n2715 0.00827857
R7250 VSS.n3166 DVSS 0.00825862
R7251 DVSS VSS.n3172 0.00825862
R7252 VSS.n4213 VSS.n4212 0.00823128
R7253 VSS.n3863 VSS.n2563 0.00822787
R7254 VSS.n3843 VSS.n2557 0.00822787
R7255 VSS.n4210 VSS.n4209 0.00821429
R7256 VSS.n5249 VSS.n2244 0.00815
R7257 VSS.n3048 VSS.n2882 0.00803695
R7258 VSS.n3003 VSS.n2878 0.00803695
R7259 VSS.n2946 VSS.n2926 0.00803521
R7260 VSS.n2945 VSS.n2928 0.00803521
R7261 VSS.n2955 VSS.n2922 0.00803521
R7262 VSS.n2971 VSS.n2917 0.00803521
R7263 VSS.n2970 VSS.n2912 0.00803521
R7264 VSS.n2979 VSS.n2978 0.00803521
R7265 VSS.n2990 VSS.n2906 0.00803521
R7266 VSS.n2989 VSS.n2908 0.00803521
R7267 VSS.n2998 VSS.n2902 0.00803521
R7268 VSS.n3018 VSS.n2897 0.00803521
R7269 VSS.n3017 VSS.n2892 0.00803521
R7270 VSS.n3026 VSS.n3025 0.00803521
R7271 VSS.n3041 VSS.n2886 0.00803521
R7272 VSS.n3040 VSS.n2888 0.00803521
R7273 VSS.n3037 VSS.n3036 0.00803521
R7274 VSS.n3052 VSS.n2880 0.00803521
R7275 VSS.n3079 VSS.n2875 0.00803521
R7276 VSS.n3078 VSS.n2870 0.00803521
R7277 VSS.n3087 VSS.n3086 0.00803521
R7278 VSS.n3094 VSS.n2863 0.00803521
R7279 VSS.n3093 VSS.n2866 0.00803521
R7280 VSS.n2865 VSS.n2857 0.00803521
R7281 VSS.n3106 VSS.n3105 0.00803521
R7282 VSS.n3117 VSS.n2851 0.00803521
R7283 VSS.n3116 VSS.n2853 0.00803521
R7284 VSS.n3125 VSS.n2847 0.00803521
R7285 VSS.n3140 VSS.n2842 0.00803521
R7286 VSS.n3139 VSS.n2837 0.00803521
R7287 VSS.n3150 VSS.n3149 0.00803521
R7288 VSS.n3162 VSS.n2830 0.00803521
R7289 VSS.n3161 VSS.n2833 0.00803521
R7290 VSS.n3169 VSS.n2826 0.00803521
R7291 VSS.n3180 VSS.n2821 0.00803521
R7292 VSS.n3179 VSS.n2816 0.00803521
R7293 VSS.n3191 VSS.n3190 0.00803521
R7294 VSS.n3238 VSS.n2802 0.00803521
R7295 VSS.n3201 VSS.n2803 0.00803521
R7296 VSS.n3231 VSS.n2809 0.00803521
R7297 VSS.n3230 VSS.n2811 0.00803521
R7298 VSS.n3227 VSS.n3226 0.00803521
R7299 VSS.n3218 VSS.n2404 0.00803521
R7300 VSS.n4877 VSS.n4876 0.00803521
R7301 VSS.n4888 VSS.n2397 0.00803521
R7302 VSS.n4887 VSS.n2400 0.00803521
R7303 VSS.n4895 VSS.n2393 0.00803521
R7304 VSS.n4914 VSS.n2388 0.00803521
R7305 VSS.n4913 VSS.n2383 0.00803521
R7306 VSS.n4924 VSS.n4923 0.00803521
R7307 VSS.n4941 VSS.n2377 0.00803521
R7308 VSS.n4940 VSS.n2379 0.00803521
R7309 VSS.n4950 VSS.n2371 0.00803521
R7310 VSS.n2373 VSS.n2372 0.00803521
R7311 VSS.n4957 VSS.n2367 0.00803521
R7312 VSS.n4968 VSS.n2359 0.00803521
R7313 VSS.n2363 VSS.n2360 0.00803521
R7314 VSS.n2362 VSS.n2351 0.00803521
R7315 VSS.n4986 VSS.n4985 0.00803521
R7316 VSS.n4997 VSS.n2344 0.00803521
R7317 VSS.n4996 VSS.n2347 0.00803521
R7318 VSS.n5004 VSS.n2340 0.00803521
R7319 VSS.n5019 VSS.n2335 0.00803521
R7320 VSS.n5018 VSS.n2330 0.00803521
R7321 VSS.n5029 VSS.n5028 0.00803521
R7322 VSS.n5040 VSS.n2323 0.00803521
R7323 VSS.n5039 VSS.n2326 0.00803521
R7324 VSS.n5047 VSS.n2319 0.00803521
R7325 VSS.n5065 VSS.n2314 0.00803521
R7326 VSS.n5064 VSS.n2309 0.00803521
R7327 VSS.n5075 VSS.n5074 0.00803521
R7328 VSS.n5090 VSS.n2303 0.00803521
R7329 VSS.n5089 VSS.n2305 0.00803521
R7330 VSS.n5098 VSS.n2297 0.00803521
R7331 VSS.n2299 VSS.n2298 0.00803521
R7332 VSS.n5105 VSS.n2293 0.00803521
R7333 VSS.n5116 VSS.n2287 0.00803521
R7334 VSS.n2288 VSS.n2283 0.00803521
R7335 VSS.n5127 VSS.n5126 0.00803521
R7336 VSS.n5170 VSS.n2277 0.00803521
R7337 VSS.n3143 VSS.n3141 0.008
R7338 VSS.n4949 VSS.n4947 0.008
R7339 VSS.n3138 VSS.n3137 0.008
R7340 VSS.n4951 VSS.n2370 0.008
R7341 VSS.n4855 VSS.n2422 0.00789286
R7342 VSS.n3367 VSS.n2416 0.00789286
R7343 VSS.n4825 VSS.n4824 0.00789286
R7344 VSS.n6 VSS.n1 0.00789286
R7345 VSS.n3375 VSS 0.00782857
R7346 VSS.n3998 DVSS 0.00782857
R7347 VSS.n4383 DVSS 0.00782857
R7348 VSS.n4382 DVSS 0.00782857
R7349 VSS.n1840 DVSS 0.00782857
R7350 DVSS VSS.n1394 0.00782857
R7351 VSS.n1393 DVSS 0.00782857
R7352 VSS.n3999 DVSS 0.00782857
R7353 VSS.n5192 DVSS 0.00782857
R7354 VSS.n5193 DVSS 0.00782857
R7355 VSS.n4823 VSS 0.00782857
R7356 VSS.n3682 VSS.n2693 0.00776429
R7357 VSS.n1878 VSS.n1773 0.00761735
R7358 VSS.n1876 VSS.n1774 0.00761735
R7359 VSS.n1916 VSS.n1915 0.00761735
R7360 VSS.n1902 VSS.n1899 0.00761735
R7361 VSS.n1954 VSS.n1953 0.00761735
R7362 VSS.n1940 VSS.n1937 0.00761735
R7363 VSS.n1739 VSS.n1676 0.00761735
R7364 VSS.n1975 VSS.n1687 0.00761735
R7365 VSS.n1733 VSS.n1649 0.00761735
R7366 VSS.n2007 VSS.n1662 0.00761735
R7367 VSS.n2043 VSS.n1629 0.00761735
R7368 VSS.n2041 VSS.n1630 0.00761735
R7369 VSS.n2022 VSS.n2021 0.00757143
R7370 VSS.n2018 VSS.n1648 0.00757143
R7371 VSS.n2017 VSS.n1651 0.00757143
R7372 VSS.n1658 VSS.n1657 0.00757143
R7373 VSS.n2011 VSS.n2010 0.00757143
R7374 VSS.n1663 VSS.n1659 0.00757143
R7375 VSS.n2005 VSS.n1664 0.00757143
R7376 VSS.n3879 VSS.n3872 0.00757143
R7377 VSS.n3876 VSS.n3759 0.00757143
R7378 VSS.n1989 VSS.n1675 0.00750714
R7379 VSS.n1986 VSS.n1985 0.00750714
R7380 VSS.n1682 VSS.n1678 0.00750714
R7381 VSS.n1979 VSS.n1683 0.00750714
R7382 VSS.n1978 VSS.n1684 0.00750714
R7383 VSS.n1689 VSS.n1688 0.00750714
R7384 VSS.n1973 VSS.n1972 0.00750714
R7385 VSS.n1792 VSS.n1788 0.00750714
R7386 VSS.n1858 VSS.n1857 0.00750714
R7387 VSS.n1854 VSS.n1798 0.00750714
R7388 VSS.n3770 VSS.n3769 0.00750714
R7389 VSS.n3923 VSS.n3922 0.00750714
R7390 VSS.n3182 VSS.n2818 0.0075
R7391 VSS.n4890 VSS.n2394 0.0075
R7392 VSS.n3174 VSS.n2823 0.0075
R7393 VSS.n2398 VSS.n2392 0.0075
R7394 VSS.n1152 VSS.n25 0.00745122
R7395 VSS.n1162 VSS.n28 0.00745122
R7396 VSS.n4089 VSS.n4086 0.00739189
R7397 VSS.n4084 VSS.n3965 0.00739189
R7398 VSS.n1879 VSS.n1770 0.00730488
R7399 VSS.n1875 VSS.n1770 0.00730488
R7400 VSS.n1914 VSS.n1913 0.00730488
R7401 VSS.n1913 VSS.n1747 0.00730488
R7402 VSS.n1952 VSS.n1951 0.00730488
R7403 VSS.n1951 VSS.n1705 0.00730488
R7404 VSS.n1738 VSS.n1737 0.00730488
R7405 VSS.n1737 VSS.n1685 0.00730488
R7406 VSS.n1732 VSS.n1731 0.00730488
R7407 VSS.n1731 VSS.n1660 0.00730488
R7408 VSS.n2044 VSS.n1626 0.00730488
R7409 VSS.n2040 VSS.n1626 0.00730488
R7410 VSS.n2940 VSS.n2939 0.00716667
R7411 VSS.n2941 VSS.n2940 0.00716667
R7412 VSS.n2941 VSS.n2910 0.00716667
R7413 VSS.n2981 VSS.n2910 0.00716667
R7414 VSS.n2982 VSS.n2981 0.00716667
R7415 VSS.n2983 VSS.n2982 0.00716667
R7416 VSS.n2984 VSS.n2983 0.00716667
R7417 VSS.n2985 VSS.n2984 0.00716667
R7418 VSS.n2985 VSS.n2890 0.00716667
R7419 VSS.n3028 VSS.n2890 0.00716667
R7420 VSS.n3029 VSS.n3028 0.00716667
R7421 VSS.n3030 VSS.n3029 0.00716667
R7422 VSS.n3031 VSS.n3030 0.00716667
R7423 VSS.n3032 VSS.n3031 0.00716667
R7424 VSS.n3033 VSS.n3032 0.00716667
R7425 VSS.n3033 VSS.n2868 0.00716667
R7426 VSS.n3089 VSS.n2868 0.00716667
R7427 VSS.n3090 VSS.n3089 0.00716667
R7428 VSS.n3091 VSS.n3090 0.00716667
R7429 VSS.n3091 VSS.n2855 0.00716667
R7430 VSS.n3108 VSS.n2855 0.00716667
R7431 VSS.n3109 VSS.n3108 0.00716667
R7432 VSS.n3110 VSS.n3109 0.00716667
R7433 VSS.n3111 VSS.n3110 0.00716667
R7434 VSS.n3112 VSS.n3111 0.00716667
R7435 VSS.n3112 VSS.n2835 0.00716667
R7436 VSS.n3152 VSS.n2835 0.00716667
R7437 VSS.n3153 VSS.n3152 0.00716667
R7438 VSS.n3154 VSS.n3153 0.00716667
R7439 VSS.n3155 VSS.n3154 0.00716667
R7440 VSS.n3157 VSS.n3155 0.00716667
R7441 VSS.n3157 VSS.n3156 0.00716667
R7442 VSS.n3156 VSS.n2815 0.00716667
R7443 VSS.n2815 VSS.n2813 0.00716667
R7444 VSS.n3195 VSS.n2813 0.00716667
R7445 VSS.n3196 VSS.n3195 0.00716667
R7446 VSS.n3197 VSS.n3196 0.00716667
R7447 VSS.n3198 VSS.n3197 0.00716667
R7448 VSS.n3198 VSS.n2402 0.00716667
R7449 VSS.n4879 VSS.n2402 0.00716667
R7450 VSS.n4880 VSS.n4879 0.00716667
R7451 VSS.n4881 VSS.n4880 0.00716667
R7452 VSS.n4882 VSS.n4881 0.00716667
R7453 VSS.n4883 VSS.n4882 0.00716667
R7454 VSS.n4883 VSS.n2381 0.00716667
R7455 VSS.n4926 VSS.n2381 0.00716667
R7456 VSS.n4927 VSS.n4926 0.00716667
R7457 VSS.n4928 VSS.n4927 0.00716667
R7458 VSS.n4929 VSS.n4928 0.00716667
R7459 VSS.n4930 VSS.n4929 0.00716667
R7460 VSS.n4931 VSS.n4930 0.00716667
R7461 VSS.n4932 VSS.n4931 0.00716667
R7462 VSS.n4933 VSS.n4932 0.00716667
R7463 VSS.n4933 VSS.n2349 0.00716667
R7464 VSS.n4988 VSS.n2349 0.00716667
R7465 VSS.n4989 VSS.n4988 0.00716667
R7466 VSS.n4990 VSS.n4989 0.00716667
R7467 VSS.n4991 VSS.n4990 0.00716667
R7468 VSS.n4992 VSS.n4991 0.00716667
R7469 VSS.n4992 VSS.n2328 0.00716667
R7470 VSS.n5031 VSS.n2328 0.00716667
R7471 VSS.n5032 VSS.n5031 0.00716667
R7472 VSS.n5033 VSS.n5032 0.00716667
R7473 VSS.n5034 VSS.n5033 0.00716667
R7474 VSS.n5035 VSS.n5034 0.00716667
R7475 VSS.n5035 VSS.n2307 0.00716667
R7476 VSS.n5077 VSS.n2307 0.00716667
R7477 VSS.n5078 VSS.n5077 0.00716667
R7478 VSS.n5079 VSS.n5078 0.00716667
R7479 VSS.n5080 VSS.n5079 0.00716667
R7480 VSS.n5081 VSS.n5080 0.00716667
R7481 VSS.n5082 VSS.n5081 0.00716667
R7482 VSS.n5083 VSS.n5082 0.00716667
R7483 VSS.n5083 VSS.n2281 0.00716667
R7484 VSS.n5129 VSS.n2281 0.00716667
R7485 VSS.n5130 VSS.n5129 0.00716667
R7486 VSS.n5131 VSS.n5130 0.00716667
R7487 VSS.n5132 VSS.n5131 0.00716667
R7488 VSS.n5133 VSS.n5132 0.00716667
R7489 VSS.n5136 VSS.n5133 0.00716667
R7490 VSS.n5137 VSS.n5136 0.00716667
R7491 VSS.n5138 VSS.n5137 0.00716667
R7492 VSS.n5141 VSS.n5138 0.00716667
R7493 VSS.n5142 VSS.n5141 0.00716667
R7494 VSS.n5143 VSS.n5142 0.00716667
R7495 VSS.n5144 VSS.n5143 0.00716667
R7496 VSS.n5146 VSS.n5144 0.00716667
R7497 VSS.n5147 VSS.n5146 0.00716667
R7498 VSS.n5148 VSS.n5147 0.00716667
R7499 VSS.n5703 VSS.n23 0.00712143
R7500 VSS.n1838 VSS.n19 0.00712143
R7501 VSS.n1298 VSS.n1297 0.00712143
R7502 VSS.n1587 VSS.n1586 0.00712143
R7503 VSS.n3561 VSS.n3560 0.00712143
R7504 VSS.n3715 VSS.n2670 0.00705714
R7505 VSS.n3714 VSS.n2654 0.00705714
R7506 VSS.n3718 VSS.n2656 0.00705714
R7507 VSS.n1004 VSS.n105 0.00700873
R7508 VSS.n3236 VSS.n2805 0.007
R7509 VSS.n3221 VSS.n2406 0.007
R7510 VSS.n3202 VSS.n2801 0.007
R7511 VSS.n3213 VSS.n3200 0.007
R7512 VSS.n3554 VSS.n3553 0.00699286
R7513 VSS.n2724 VSS.n2719 0.00699286
R7514 VSS.n3517 VSS.n2734 0.00692857
R7515 VSS.n4134 VSS.n4133 0.006875
R7516 VSS.n4131 VSS.n3768 0.006875
R7517 VSS.n4143 VSS.n3756 0.006875
R7518 VSS.n4146 VSS.n4145 0.006875
R7519 VSS.n4852 VSS.n4842 0.0068
R7520 VSS.n1700 VSS.n1696 0.0068
R7521 VSS.n1958 VSS.n1957 0.0068
R7522 VSS.n1706 VSS.n1701 0.0068
R7523 VSS.n1950 VSS.n1707 0.0068
R7524 VSS.n1949 VSS.n1708 0.0068
R7525 VSS.n1715 VSS.n1714 0.0068
R7526 VSS.n1943 VSS.n1942 0.0068
R7527 VSS.n4750 VSS.n4749 0.0068
R7528 VSS.n1154 VSS.n25 0.00671951
R7529 VSS.n1160 VSS.n28 0.00671951
R7530 VSS.n4244 VSS.n4235 0.00658571
R7531 VSS.n4245 VSS.n4244 0.00658571
R7532 VSS.n4246 VSS.n4245 0.00658571
R7533 VSS.n4246 VSS.n4231 0.00658571
R7534 VSS.n4252 VSS.n4231 0.00658571
R7535 VSS.n4253 VSS.n4252 0.00658571
R7536 VSS.n4254 VSS.n4253 0.00658571
R7537 VSS.n4254 VSS.n4227 0.00658571
R7538 VSS.n4260 VSS.n4227 0.00658571
R7539 VSS.n4261 VSS.n4260 0.00658571
R7540 VSS.n4262 VSS.n4261 0.00658571
R7541 VSS.n4262 VSS.n4223 0.00658571
R7542 VSS.n4268 VSS.n4223 0.00658571
R7543 VSS.n4269 VSS.n4268 0.00658571
R7544 VSS.n4298 VSS.n4269 0.00658571
R7545 VSS.n4298 VSS.n4297 0.00658571
R7546 VSS.n4297 VSS.n4296 0.00658571
R7547 VSS.n4296 VSS.n4270 0.00658571
R7548 VSS.n4290 VSS.n4270 0.00658571
R7549 VSS.n4290 VSS.n4289 0.00658571
R7550 VSS.n4289 VSS.n4288 0.00658571
R7551 VSS.n4288 VSS.n4274 0.00658571
R7552 VSS.n4280 VSS.n4274 0.00658571
R7553 VSS.n4280 VSS.n2504 0.00658571
R7554 VSS.n4679 VSS.n2504 0.00658571
R7555 VSS.n4680 VSS.n4679 0.00658571
R7556 VSS.n4681 VSS.n4680 0.00658571
R7557 VSS.n4681 VSS.n2498 0.00658571
R7558 VSS.n4689 VSS.n2498 0.00658571
R7559 VSS.n4690 VSS.n4689 0.00658571
R7560 VSS.n4691 VSS.n4690 0.00658571
R7561 VSS.n4691 VSS.n2494 0.00658571
R7562 VSS.n4697 VSS.n2494 0.00658571
R7563 VSS.n4698 VSS.n4697 0.00658571
R7564 VSS.n4699 VSS.n4698 0.00658571
R7565 VSS.n4699 VSS.n2490 0.00658571
R7566 VSS.n4705 VSS.n2490 0.00658571
R7567 VSS.n4706 VSS.n4705 0.00658571
R7568 VSS.n4707 VSS.n4706 0.00658571
R7569 VSS.n4707 VSS.n2486 0.00658571
R7570 VSS.n4713 VSS.n2486 0.00658571
R7571 VSS.n4714 VSS.n4713 0.00658571
R7572 VSS.n4715 VSS.n4714 0.00658571
R7573 VSS.n4715 VSS.n2482 0.00658571
R7574 VSS.n4721 VSS.n2482 0.00658571
R7575 VSS.n4722 VSS.n4721 0.00658571
R7576 VSS.n4723 VSS.n4722 0.00658571
R7577 VSS.n4723 VSS.n2478 0.00658571
R7578 VSS.n4729 VSS.n2478 0.00658571
R7579 VSS.n4730 VSS.n4729 0.00658571
R7580 VSS.n4731 VSS.n4730 0.00658571
R7581 VSS.n4731 VSS.n2474 0.00658571
R7582 VSS.n4737 VSS.n2474 0.00658571
R7583 VSS.n4738 VSS.n4737 0.00658571
R7584 VSS.n4739 VSS.n4738 0.00658571
R7585 VSS.n4739 VSS.n2470 0.00658571
R7586 VSS.n4745 VSS.n2470 0.00658571
R7587 VSS.n4746 VSS.n4745 0.00658571
R7588 VSS.n4747 VSS.n4746 0.00658571
R7589 VSS.n4747 VSS.n2466 0.00658571
R7590 VSS.n4754 VSS.n2466 0.00658571
R7591 VSS.n4755 VSS.n4754 0.00658571
R7592 VSS.n4756 VSS.n4755 0.00658571
R7593 VSS.n4756 VSS.n2462 0.00658571
R7594 VSS.n4762 VSS.n2462 0.00658571
R7595 VSS.n4763 VSS.n4762 0.00658571
R7596 VSS.n4764 VSS.n4763 0.00658571
R7597 VSS.n4764 VSS.n2458 0.00658571
R7598 VSS.n4770 VSS.n2458 0.00658571
R7599 VSS.n4771 VSS.n4770 0.00658571
R7600 VSS.n4772 VSS.n4771 0.00658571
R7601 VSS.n4772 VSS.n2454 0.00658571
R7602 VSS.n4778 VSS.n2454 0.00658571
R7603 VSS.n4779 VSS.n4778 0.00658571
R7604 VSS.n4780 VSS.n4779 0.00658571
R7605 VSS.n4780 VSS.n2450 0.00658571
R7606 VSS.n4786 VSS.n2450 0.00658571
R7607 VSS.n4787 VSS.n4786 0.00658571
R7608 VSS.n4788 VSS.n4787 0.00658571
R7609 VSS.n4788 VSS.n2446 0.00658571
R7610 VSS.n4794 VSS.n2446 0.00658571
R7611 VSS.n4795 VSS.n4794 0.00658571
R7612 VSS.n4796 VSS.n4795 0.00658571
R7613 VSS.n4796 VSS.n2442 0.00658571
R7614 VSS.n4802 VSS.n2442 0.00658571
R7615 VSS.n4803 VSS.n4802 0.00658571
R7616 VSS.n4804 VSS.n4803 0.00658571
R7617 VSS.n4804 VSS.n2438 0.00658571
R7618 VSS.n4810 VSS.n2438 0.00658571
R7619 VSS.n4811 VSS.n4810 0.00658571
R7620 VSS.n4812 VSS.n4811 0.00658571
R7621 VSS.n4812 VSS.n2434 0.00658571
R7622 VSS.n4819 VSS.n2434 0.00658571
R7623 VSS.n4820 VSS.n4819 0.00658571
R7624 VSS.n4821 VSS.n4820 0.00658571
R7625 VSS.n4821 VSS.n3 0.00658571
R7626 VSS.n5721 VSS.n3 0.00658571
R7627 VSS.n5720 VSS.n5719 0.00658571
R7628 VSS.n2771 VSS.n2770 0.00658571
R7629 VSS.n2772 VSS.n2771 0.00658571
R7630 VSS.n2772 VSS.n2758 0.00658571
R7631 VSS.n2778 VSS.n2758 0.00658571
R7632 VSS.n2779 VSS.n2778 0.00658571
R7633 VSS.n2780 VSS.n2779 0.00658571
R7634 VSS.n2780 VSS.n2754 0.00658571
R7635 VSS.n2786 VSS.n2754 0.00658571
R7636 VSS.n2787 VSS.n2786 0.00658571
R7637 VSS.n2788 VSS.n2787 0.00658571
R7638 VSS.n2788 VSS.n2750 0.00658571
R7639 VSS.n3265 VSS.n2750 0.00658571
R7640 VSS.n3266 VSS.n3265 0.00658571
R7641 VSS.n3267 VSS.n3266 0.00658571
R7642 VSS.n3267 VSS.n2746 0.00658571
R7643 VSS.n3273 VSS.n2746 0.00658571
R7644 VSS.n3274 VSS.n3273 0.00658571
R7645 VSS.n3275 VSS.n3274 0.00658571
R7646 VSS.n3275 VSS.n2742 0.00658571
R7647 VSS.n3281 VSS.n2742 0.00658571
R7648 VSS.n3282 VSS.n3281 0.00658571
R7649 VSS.n3283 VSS.n3282 0.00658571
R7650 VSS.n3283 VSS.n2738 0.00658571
R7651 VSS.n3289 VSS.n2738 0.00658571
R7652 VSS.n3290 VSS.n3289 0.00658571
R7653 VSS.n3514 VSS.n3290 0.00658571
R7654 VSS.n3514 VSS.n3513 0.00658571
R7655 VSS.n3513 VSS.n3512 0.00658571
R7656 VSS.n3512 VSS.n3291 0.00658571
R7657 VSS.n3506 VSS.n3291 0.00658571
R7658 VSS.n3506 VSS.n3505 0.00658571
R7659 VSS.n3505 VSS.n3504 0.00658571
R7660 VSS.n3504 VSS.n3295 0.00658571
R7661 VSS.n3498 VSS.n3295 0.00658571
R7662 VSS.n3498 VSS.n3497 0.00658571
R7663 VSS.n3497 VSS.n3496 0.00658571
R7664 VSS.n3496 VSS.n3299 0.00658571
R7665 VSS.n3490 VSS.n3299 0.00658571
R7666 VSS.n3490 VSS.n3489 0.00658571
R7667 VSS.n3489 VSS.n3488 0.00658571
R7668 VSS.n3488 VSS.n3303 0.00658571
R7669 VSS.n3482 VSS.n3303 0.00658571
R7670 VSS.n3482 VSS.n3481 0.00658571
R7671 VSS.n3481 VSS.n3480 0.00658571
R7672 VSS.n3480 VSS.n3307 0.00658571
R7673 VSS.n3474 VSS.n3307 0.00658571
R7674 VSS.n3474 VSS.n3473 0.00658571
R7675 VSS.n3473 VSS.n3472 0.00658571
R7676 VSS.n3472 VSS.n3311 0.00658571
R7677 VSS.n3466 VSS.n3311 0.00658571
R7678 VSS.n3466 VSS.n3465 0.00658571
R7679 VSS.n3465 VSS.n3464 0.00658571
R7680 VSS.n3464 VSS.n3315 0.00658571
R7681 VSS.n3458 VSS.n3315 0.00658571
R7682 VSS.n3458 VSS.n3457 0.00658571
R7683 VSS.n3457 VSS.n3456 0.00658571
R7684 VSS.n3456 VSS.n3319 0.00658571
R7685 VSS.n3450 VSS.n3319 0.00658571
R7686 VSS.n3450 VSS.n3449 0.00658571
R7687 VSS.n3449 VSS.n3448 0.00658571
R7688 VSS.n3448 VSS.n3323 0.00658571
R7689 VSS.n3442 VSS.n3323 0.00658571
R7690 VSS.n3442 VSS.n3441 0.00658571
R7691 VSS.n3441 VSS.n3440 0.00658571
R7692 VSS.n3440 VSS.n3327 0.00658571
R7693 VSS.n3434 VSS.n3327 0.00658571
R7694 VSS.n3434 VSS.n3433 0.00658571
R7695 VSS.n3433 VSS.n3432 0.00658571
R7696 VSS.n3432 VSS.n3331 0.00658571
R7697 VSS.n3426 VSS.n3331 0.00658571
R7698 VSS.n3426 VSS.n3425 0.00658571
R7699 VSS.n3425 VSS.n3424 0.00658571
R7700 VSS.n3424 VSS.n3335 0.00658571
R7701 VSS.n3418 VSS.n3335 0.00658571
R7702 VSS.n3418 VSS.n3417 0.00658571
R7703 VSS.n3417 VSS.n3416 0.00658571
R7704 VSS.n3416 VSS.n3339 0.00658571
R7705 VSS.n3410 VSS.n3339 0.00658571
R7706 VSS.n3410 VSS.n3409 0.00658571
R7707 VSS.n3409 VSS.n3408 0.00658571
R7708 VSS.n3408 VSS.n3343 0.00658571
R7709 VSS.n3402 VSS.n3343 0.00658571
R7710 VSS.n3402 VSS.n3401 0.00658571
R7711 VSS.n3401 VSS.n3400 0.00658571
R7712 VSS.n3400 VSS.n3347 0.00658571
R7713 VSS.n3394 VSS.n3347 0.00658571
R7714 VSS.n3394 VSS.n3393 0.00658571
R7715 VSS.n3393 VSS.n3392 0.00658571
R7716 VSS.n3392 VSS.n3351 0.00658571
R7717 VSS.n3386 VSS.n3351 0.00658571
R7718 VSS.n3386 VSS.n3385 0.00658571
R7719 VSS.n3385 VSS.n3384 0.00658571
R7720 VSS.n3384 VSS.n3355 0.00658571
R7721 VSS.n3378 VSS.n3355 0.00658571
R7722 VSS.n3378 VSS.n3377 0.00658571
R7723 VSS.n3377 VSS.n3376 0.00658571
R7724 VSS.n3376 VSS.n3358 0.00658571
R7725 VSS.n3362 VSS.n3360 0.00658571
R7726 VSS.n4187 VSS.n4186 0.00658571
R7727 VSS.n4186 VSS.n4185 0.00658571
R7728 VSS.n4185 VSS.n2641 0.00658571
R7729 VSS.n4179 VSS.n2641 0.00658571
R7730 VSS.n4179 VSS.n4178 0.00658571
R7731 VSS.n4178 VSS.n4177 0.00658571
R7732 VSS.n4177 VSS.n2646 0.00658571
R7733 VSS.n3800 VSS.n2646 0.00658571
R7734 VSS.n3801 VSS.n3800 0.00658571
R7735 VSS.n3801 VSS.n3792 0.00658571
R7736 VSS.n3809 VSS.n3792 0.00658571
R7737 VSS.n3810 VSS.n3809 0.00658571
R7738 VSS.n3811 VSS.n3810 0.00658571
R7739 VSS.n3811 VSS.n3738 0.00658571
R7740 VSS.n4158 VSS.n3738 0.00658571
R7741 VSS.n4158 VSS.n4157 0.00658571
R7742 VSS.n4157 VSS.n4156 0.00658571
R7743 VSS.n4156 VSS.n3739 0.00658571
R7744 VSS.n3873 VSS.n3739 0.00658571
R7745 VSS.n3873 VSS.n3765 0.00658571
R7746 VSS.n4140 VSS.n3765 0.00658571
R7747 VSS.n4140 VSS.n4139 0.00658571
R7748 VSS.n4139 VSS.n4138 0.00658571
R7749 VSS.n4138 VSS.n3766 0.00658571
R7750 VSS.n3916 VSS.n3766 0.00658571
R7751 VSS.n3934 VSS.n3916 0.00658571
R7752 VSS.n3935 VSS.n3934 0.00658571
R7753 VSS.n3937 VSS.n3935 0.00658571
R7754 VSS.n3937 VSS.n3936 0.00658571
R7755 VSS.n3936 VSS.n3896 0.00658571
R7756 VSS.n4111 VSS.n3896 0.00658571
R7757 VSS.n4111 VSS.n4110 0.00658571
R7758 VSS.n4110 VSS.n4109 0.00658571
R7759 VSS.n4109 VSS.n3897 0.00658571
R7760 VSS.n3961 VSS.n3897 0.00658571
R7761 VSS.n4095 VSS.n3961 0.00658571
R7762 VSS.n4095 VSS.n4094 0.00658571
R7763 VSS.n4094 VSS.n4093 0.00658571
R7764 VSS.n4093 VSS.n3962 0.00658571
R7765 VSS.n4053 VSS.n3962 0.00658571
R7766 VSS.n4053 VSS.n4052 0.00658571
R7767 VSS.n4052 VSS.n4051 0.00658571
R7768 VSS.n4051 VSS.n3968 0.00658571
R7769 VSS.n4045 VSS.n3968 0.00658571
R7770 VSS.n4045 VSS.n4044 0.00658571
R7771 VSS.n4044 VSS.n4043 0.00658571
R7772 VSS.n4043 VSS.n3972 0.00658571
R7773 VSS.n4037 VSS.n3972 0.00658571
R7774 VSS.n4037 VSS.n4036 0.00658571
R7775 VSS.n4036 VSS.n4035 0.00658571
R7776 VSS.n4035 VSS.n3976 0.00658571
R7777 VSS.n4029 VSS.n3976 0.00658571
R7778 VSS.n4029 VSS.n4028 0.00658571
R7779 VSS.n4028 VSS.n4027 0.00658571
R7780 VSS.n4027 VSS.n3980 0.00658571
R7781 VSS.n4021 VSS.n3980 0.00658571
R7782 VSS.n4021 VSS.n4020 0.00658571
R7783 VSS.n4020 VSS.n4019 0.00658571
R7784 VSS.n4019 VSS.n3984 0.00658571
R7785 VSS.n4013 VSS.n3984 0.00658571
R7786 VSS.n4013 VSS.n4012 0.00658571
R7787 VSS.n4012 VSS.n4011 0.00658571
R7788 VSS.n4011 VSS.n3988 0.00658571
R7789 VSS.n4005 VSS.n3988 0.00658571
R7790 VSS.n4005 VSS.n4004 0.00658571
R7791 VSS.n4004 VSS.n4003 0.00658571
R7792 VSS.n4003 VSS.n3992 0.00658571
R7793 VSS.n3997 VSS.n3992 0.00658571
R7794 VSS.n3997 VSS.n3996 0.00658571
R7795 VSS.n2553 VSS.n2550 0.00658571
R7796 VSS.n4519 VSS.n2553 0.00658571
R7797 VSS.n4519 VSS.n4518 0.00658571
R7798 VSS.n4518 VSS.n4517 0.00658571
R7799 VSS.n4517 VSS.n2554 0.00658571
R7800 VSS.n4509 VSS.n2554 0.00658571
R7801 VSS.n4509 VSS.n4508 0.00658571
R7802 VSS.n4508 VSS.n4507 0.00658571
R7803 VSS.n4507 VSS.n2571 0.00658571
R7804 VSS.n4501 VSS.n2571 0.00658571
R7805 VSS.n4501 VSS.n4500 0.00658571
R7806 VSS.n4500 VSS.n4499 0.00658571
R7807 VSS.n4499 VSS.n2575 0.00658571
R7808 VSS.n4493 VSS.n2575 0.00658571
R7809 VSS.n4493 VSS.n4492 0.00658571
R7810 VSS.n4492 VSS.n4491 0.00658571
R7811 VSS.n4491 VSS.n2579 0.00658571
R7812 VSS.n4485 VSS.n2579 0.00658571
R7813 VSS.n4485 VSS.n4484 0.00658571
R7814 VSS.n4484 VSS.n4483 0.00658571
R7815 VSS.n4483 VSS.n2583 0.00658571
R7816 VSS.n4477 VSS.n2583 0.00658571
R7817 VSS.n4477 VSS.n4476 0.00658571
R7818 VSS.n4476 VSS.n4475 0.00658571
R7819 VSS.n4475 VSS.n2587 0.00658571
R7820 VSS.n4469 VSS.n2587 0.00658571
R7821 VSS.n4469 VSS.n4468 0.00658571
R7822 VSS.n4468 VSS.n4467 0.00658571
R7823 VSS.n4467 VSS.n2591 0.00658571
R7824 VSS.n4461 VSS.n2591 0.00658571
R7825 VSS.n4461 VSS.n4460 0.00658571
R7826 VSS.n4460 VSS.n4459 0.00658571
R7827 VSS.n4459 VSS.n2595 0.00658571
R7828 VSS.n4453 VSS.n2595 0.00658571
R7829 VSS.n4453 VSS.n4452 0.00658571
R7830 VSS.n4452 VSS.n4451 0.00658571
R7831 VSS.n4451 VSS.n2599 0.00658571
R7832 VSS.n4445 VSS.n2599 0.00658571
R7833 VSS.n4445 VSS.n4444 0.00658571
R7834 VSS.n4444 VSS.n4443 0.00658571
R7835 VSS.n4443 VSS.n2603 0.00658571
R7836 VSS.n4353 VSS.n2603 0.00658571
R7837 VSS.n4354 VSS.n4353 0.00658571
R7838 VSS.n4434 VSS.n4354 0.00658571
R7839 VSS.n4434 VSS.n4433 0.00658571
R7840 VSS.n4433 VSS.n4432 0.00658571
R7841 VSS.n4432 VSS.n4355 0.00658571
R7842 VSS.n4426 VSS.n4355 0.00658571
R7843 VSS.n4426 VSS.n4425 0.00658571
R7844 VSS.n4425 VSS.n4424 0.00658571
R7845 VSS.n4424 VSS.n4359 0.00658571
R7846 VSS.n4418 VSS.n4359 0.00658571
R7847 VSS.n4418 VSS.n4417 0.00658571
R7848 VSS.n4417 VSS.n4416 0.00658571
R7849 VSS.n4416 VSS.n4363 0.00658571
R7850 VSS.n4410 VSS.n4363 0.00658571
R7851 VSS.n4410 VSS.n4409 0.00658571
R7852 VSS.n4409 VSS.n4408 0.00658571
R7853 VSS.n4408 VSS.n4367 0.00658571
R7854 VSS.n4402 VSS.n4367 0.00658571
R7855 VSS.n4402 VSS.n4401 0.00658571
R7856 VSS.n4401 VSS.n4400 0.00658571
R7857 VSS.n4400 VSS.n4371 0.00658571
R7858 VSS.n4394 VSS.n4371 0.00658571
R7859 VSS.n4394 VSS.n4393 0.00658571
R7860 VSS.n4393 VSS.n4392 0.00658571
R7861 VSS.n4392 VSS.n4375 0.00658571
R7862 VSS.n4386 VSS.n4375 0.00658571
R7863 VSS.n4386 VSS.n4385 0.00658571
R7864 VSS.n4385 VSS.n4384 0.00658571
R7865 VSS.n4384 VSS.n4379 0.00658571
R7866 VSS.n2059 VSS.n2058 0.00658571
R7867 VSS.n2058 VSS.n2057 0.00658571
R7868 VSS.n2057 VSS.n1615 0.00658571
R7869 VSS.n2051 VSS.n1615 0.00658571
R7870 VSS.n2051 VSS.n2050 0.00658571
R7871 VSS.n2050 VSS.n2049 0.00658571
R7872 VSS.n2049 VSS.n1620 0.00658571
R7873 VSS.n1637 VSS.n1620 0.00658571
R7874 VSS.n2035 VSS.n1637 0.00658571
R7875 VSS.n2035 VSS.n2034 0.00658571
R7876 VSS.n2034 VSS.n2033 0.00658571
R7877 VSS.n2033 VSS.n1638 0.00658571
R7878 VSS.n2027 VSS.n1638 0.00658571
R7879 VSS.n2027 VSS.n2026 0.00658571
R7880 VSS.n2026 VSS.n2025 0.00658571
R7881 VSS.n2025 VSS.n1646 0.00658571
R7882 VSS.n1654 VSS.n1646 0.00658571
R7883 VSS.n2015 VSS.n1654 0.00658571
R7884 VSS.n2015 VSS.n2014 0.00658571
R7885 VSS.n2014 VSS.n2013 0.00658571
R7886 VSS.n2013 VSS.n1655 0.00658571
R7887 VSS.n1668 VSS.n1655 0.00658571
R7888 VSS.n2002 VSS.n1668 0.00658571
R7889 VSS.n2002 VSS.n2001 0.00658571
R7890 VSS.n2001 VSS.n2000 0.00658571
R7891 VSS.n2000 VSS.n1669 0.00658571
R7892 VSS.n1994 VSS.n1669 0.00658571
R7893 VSS.n1994 VSS.n1993 0.00658571
R7894 VSS.n1993 VSS.n1992 0.00658571
R7895 VSS.n1992 VSS.n1673 0.00658571
R7896 VSS.n1983 VSS.n1673 0.00658571
R7897 VSS.n1983 VSS.n1982 0.00658571
R7898 VSS.n1982 VSS.n1981 0.00658571
R7899 VSS.n1981 VSS.n1680 0.00658571
R7900 VSS.n1693 VSS.n1680 0.00658571
R7901 VSS.n1970 VSS.n1693 0.00658571
R7902 VSS.n1970 VSS.n1969 0.00658571
R7903 VSS.n1969 VSS.n1968 0.00658571
R7904 VSS.n1968 VSS.n1694 0.00658571
R7905 VSS.n1962 VSS.n1694 0.00658571
R7906 VSS.n1962 VSS.n1961 0.00658571
R7907 VSS.n1961 VSS.n1960 0.00658571
R7908 VSS.n1960 VSS.n1698 0.00658571
R7909 VSS.n1711 VSS.n1698 0.00658571
R7910 VSS.n1947 VSS.n1711 0.00658571
R7911 VSS.n1947 VSS.n1946 0.00658571
R7912 VSS.n1946 VSS.n1945 0.00658571
R7913 VSS.n1945 VSS.n1712 0.00658571
R7914 VSS.n1932 VSS.n1712 0.00658571
R7915 VSS.n1932 VSS.n1931 0.00658571
R7916 VSS.n1931 VSS.n1930 0.00658571
R7917 VSS.n1930 VSS.n1718 0.00658571
R7918 VSS.n1924 VSS.n1718 0.00658571
R7919 VSS.n1924 VSS.n1923 0.00658571
R7920 VSS.n1923 VSS.n1922 0.00658571
R7921 VSS.n1922 VSS.n1722 0.00658571
R7922 VSS.n1753 VSS.n1722 0.00658571
R7923 VSS.n1909 VSS.n1753 0.00658571
R7924 VSS.n1909 VSS.n1908 0.00658571
R7925 VSS.n1908 VSS.n1907 0.00658571
R7926 VSS.n1907 VSS.n1754 0.00658571
R7927 VSS.n1894 VSS.n1754 0.00658571
R7928 VSS.n1894 VSS.n1893 0.00658571
R7929 VSS.n1893 VSS.n1892 0.00658571
R7930 VSS.n1892 VSS.n1760 0.00658571
R7931 VSS.n1886 VSS.n1760 0.00658571
R7932 VSS.n1886 VSS.n1885 0.00658571
R7933 VSS.n1885 VSS.n1884 0.00658571
R7934 VSS.n1884 VSS.n1764 0.00658571
R7935 VSS.n1781 VSS.n1764 0.00658571
R7936 VSS.n1870 VSS.n1781 0.00658571
R7937 VSS.n1870 VSS.n1869 0.00658571
R7938 VSS.n1869 VSS.n1868 0.00658571
R7939 VSS.n1868 VSS.n1782 0.00658571
R7940 VSS.n1862 VSS.n1782 0.00658571
R7941 VSS.n1862 VSS.n1861 0.00658571
R7942 VSS.n1861 VSS.n1860 0.00658571
R7943 VSS.n1860 VSS.n1790 0.00658571
R7944 VSS.n1851 VSS.n1790 0.00658571
R7945 VSS.n1851 VSS.n1850 0.00658571
R7946 VSS.n1850 VSS.n1849 0.00658571
R7947 VSS.n1849 VSS.n1823 0.00658571
R7948 VSS.n1843 VSS.n1823 0.00658571
R7949 VSS.n1843 VSS.n1842 0.00658571
R7950 VSS.n1842 VSS.n1841 0.00658571
R7951 VSS.n1841 VSS.n1827 0.00658571
R7952 VSS.n1831 VSS.n1829 0.00658571
R7953 VSS.n1584 VSS.n1583 0.00658571
R7954 VSS.n1583 VSS.n1582 0.00658571
R7955 VSS.n1582 VSS.n1303 0.00658571
R7956 VSS.n1576 VSS.n1303 0.00658571
R7957 VSS.n1576 VSS.n1575 0.00658571
R7958 VSS.n1575 VSS.n1574 0.00658571
R7959 VSS.n1574 VSS.n1307 0.00658571
R7960 VSS.n1568 VSS.n1307 0.00658571
R7961 VSS.n1568 VSS.n1567 0.00658571
R7962 VSS.n1567 VSS.n1566 0.00658571
R7963 VSS.n1566 VSS.n1311 0.00658571
R7964 VSS.n1560 VSS.n1311 0.00658571
R7965 VSS.n1560 VSS.n1559 0.00658571
R7966 VSS.n1559 VSS.n1558 0.00658571
R7967 VSS.n1558 VSS.n1315 0.00658571
R7968 VSS.n1552 VSS.n1315 0.00658571
R7969 VSS.n1552 VSS.n1551 0.00658571
R7970 VSS.n1551 VSS.n1550 0.00658571
R7971 VSS.n1550 VSS.n1319 0.00658571
R7972 VSS.n1544 VSS.n1319 0.00658571
R7973 VSS.n1544 VSS.n1543 0.00658571
R7974 VSS.n1543 VSS.n1542 0.00658571
R7975 VSS.n1542 VSS.n1323 0.00658571
R7976 VSS.n1536 VSS.n1323 0.00658571
R7977 VSS.n1536 VSS.n1535 0.00658571
R7978 VSS.n1535 VSS.n1534 0.00658571
R7979 VSS.n1534 VSS.n1327 0.00658571
R7980 VSS.n1528 VSS.n1327 0.00658571
R7981 VSS.n1528 VSS.n1527 0.00658571
R7982 VSS.n1527 VSS.n1526 0.00658571
R7983 VSS.n1526 VSS.n1331 0.00658571
R7984 VSS.n1520 VSS.n1331 0.00658571
R7985 VSS.n1520 VSS.n1519 0.00658571
R7986 VSS.n1519 VSS.n1518 0.00658571
R7987 VSS.n1518 VSS.n1335 0.00658571
R7988 VSS.n1512 VSS.n1335 0.00658571
R7989 VSS.n1512 VSS.n1511 0.00658571
R7990 VSS.n1511 VSS.n1510 0.00658571
R7991 VSS.n1510 VSS.n1339 0.00658571
R7992 VSS.n1504 VSS.n1339 0.00658571
R7993 VSS.n1504 VSS.n1503 0.00658571
R7994 VSS.n1503 VSS.n1502 0.00658571
R7995 VSS.n1502 VSS.n1343 0.00658571
R7996 VSS.n1496 VSS.n1343 0.00658571
R7997 VSS.n1496 VSS.n1495 0.00658571
R7998 VSS.n1495 VSS.n1494 0.00658571
R7999 VSS.n1494 VSS.n1347 0.00658571
R8000 VSS.n1488 VSS.n1347 0.00658571
R8001 VSS.n1488 VSS.n1487 0.00658571
R8002 VSS.n1487 VSS.n1486 0.00658571
R8003 VSS.n1486 VSS.n1351 0.00658571
R8004 VSS.n1480 VSS.n1351 0.00658571
R8005 VSS.n1480 VSS.n1479 0.00658571
R8006 VSS.n1479 VSS.n1478 0.00658571
R8007 VSS.n1478 VSS.n1355 0.00658571
R8008 VSS.n1472 VSS.n1355 0.00658571
R8009 VSS.n1472 VSS.n1471 0.00658571
R8010 VSS.n1471 VSS.n1470 0.00658571
R8011 VSS.n1470 VSS.n1359 0.00658571
R8012 VSS.n1464 VSS.n1359 0.00658571
R8013 VSS.n1464 VSS.n1463 0.00658571
R8014 VSS.n1463 VSS.n1462 0.00658571
R8015 VSS.n1462 VSS.n1363 0.00658571
R8016 VSS.n1456 VSS.n1363 0.00658571
R8017 VSS.n1456 VSS.n1455 0.00658571
R8018 VSS.n1455 VSS.n1454 0.00658571
R8019 VSS.n1454 VSS.n1367 0.00658571
R8020 VSS.n1448 VSS.n1367 0.00658571
R8021 VSS.n1448 VSS.n1447 0.00658571
R8022 VSS.n1447 VSS.n1446 0.00658571
R8023 VSS.n1446 VSS.n1371 0.00658571
R8024 VSS.n1440 VSS.n1371 0.00658571
R8025 VSS.n1440 VSS.n1439 0.00658571
R8026 VSS.n1439 VSS.n1438 0.00658571
R8027 VSS.n1438 VSS.n1375 0.00658571
R8028 VSS.n1432 VSS.n1375 0.00658571
R8029 VSS.n1432 VSS.n1431 0.00658571
R8030 VSS.n1431 VSS.n1430 0.00658571
R8031 VSS.n1430 VSS.n1379 0.00658571
R8032 VSS.n1424 VSS.n1379 0.00658571
R8033 VSS.n1424 VSS.n1423 0.00658571
R8034 VSS.n1423 VSS.n1422 0.00658571
R8035 VSS.n1422 VSS.n1383 0.00658571
R8036 VSS.n1416 VSS.n1383 0.00658571
R8037 VSS.n1416 VSS.n1415 0.00658571
R8038 VSS.n1415 VSS.n1414 0.00658571
R8039 VSS.n1414 VSS.n1387 0.00658571
R8040 VSS.n1408 VSS.n1387 0.00658571
R8041 VSS.n1408 VSS.n1407 0.00658571
R8042 VSS.n1407 VSS.n1406 0.00658571
R8043 VSS.n1406 VSS.n1391 0.00658571
R8044 VSS.n1400 VSS.n1391 0.00658571
R8045 VSS.n1400 VSS.n1399 0.00658571
R8046 VSS.n1399 VSS.n1398 0.00658571
R8047 VSS.n3558 VSS.n3542 0.00658571
R8048 VSS.n3558 VSS.n3557 0.00658571
R8049 VSS.n3557 VSS.n3556 0.00658571
R8050 VSS.n3556 VSS.n3543 0.00658571
R8051 VSS.n3549 VSS.n3543 0.00658571
R8052 VSS.n3549 VSS.n3548 0.00658571
R8053 VSS.n3548 VSS.n2721 0.00658571
R8054 VSS.n3571 VSS.n2721 0.00658571
R8055 VSS.n3572 VSS.n3571 0.00658571
R8056 VSS.n3573 VSS.n3572 0.00658571
R8057 VSS.n3573 VSS.n2717 0.00658571
R8058 VSS.n3580 VSS.n2717 0.00658571
R8059 VSS.n3581 VSS.n3580 0.00658571
R8060 VSS.n3582 VSS.n3581 0.00658571
R8061 VSS.n3582 VSS.n2713 0.00658571
R8062 VSS.n3590 VSS.n2713 0.00658571
R8063 VSS.n3591 VSS.n3590 0.00658571
R8064 VSS.n3596 VSS.n3591 0.00658571
R8065 VSS.n3596 VSS.n3595 0.00658571
R8066 VSS.n3595 VSS.n3594 0.00658571
R8067 VSS.n3594 VSS.n2676 0.00658571
R8068 VSS.n3712 VSS.n2676 0.00658571
R8069 VSS.n3712 VSS.n3711 0.00658571
R8070 VSS.n3711 VSS.n3710 0.00658571
R8071 VSS.n3710 VSS.n2677 0.00658571
R8072 VSS.n2681 VSS.n2677 0.00658571
R8073 VSS.n3703 VSS.n2681 0.00658571
R8074 VSS.n3703 VSS.n3702 0.00658571
R8075 VSS.n3702 VSS.n3701 0.00658571
R8076 VSS.n3701 VSS.n2682 0.00658571
R8077 VSS.n3695 VSS.n2682 0.00658571
R8078 VSS.n3695 VSS.n3694 0.00658571
R8079 VSS.n3694 VSS.n3693 0.00658571
R8080 VSS.n3693 VSS.n2686 0.00658571
R8081 VSS.n3687 VSS.n2686 0.00658571
R8082 VSS.n3687 VSS.n3686 0.00658571
R8083 VSS.n3686 VSS.n3685 0.00658571
R8084 VSS.n3685 VSS.n2690 0.00658571
R8085 VSS.n3635 VSS.n2690 0.00658571
R8086 VSS.n3635 VSS.n3633 0.00658571
R8087 VSS.n3644 VSS.n3633 0.00658571
R8088 VSS.n3645 VSS.n3644 0.00658571
R8089 VSS.n3646 VSS.n3645 0.00658571
R8090 VSS.n3646 VSS.n3629 0.00658571
R8091 VSS.n3654 VSS.n3629 0.00658571
R8092 VSS.n3655 VSS.n3654 0.00658571
R8093 VSS.n3670 VSS.n3655 0.00658571
R8094 VSS.n3670 VSS.n3669 0.00658571
R8095 VSS.n3669 VSS.n3668 0.00658571
R8096 VSS.n3668 VSS.n3656 0.00658571
R8097 VSS.n3661 VSS.n3656 0.00658571
R8098 VSS.n3661 VSS.n3660 0.00658571
R8099 VSS.n3660 VSS.n2247 0.00658571
R8100 VSS.n5247 VSS.n2247 0.00658571
R8101 VSS.n5247 VSS.n5246 0.00658571
R8102 VSS.n5246 VSS.n5245 0.00658571
R8103 VSS.n5245 VSS.n2248 0.00658571
R8104 VSS.n5239 VSS.n2248 0.00658571
R8105 VSS.n5239 VSS.n5238 0.00658571
R8106 VSS.n5238 VSS.n5237 0.00658571
R8107 VSS.n5237 VSS.n2253 0.00658571
R8108 VSS.n5231 VSS.n2253 0.00658571
R8109 VSS.n5231 VSS.n5230 0.00658571
R8110 VSS.n5230 VSS.n5229 0.00658571
R8111 VSS.n5229 VSS.n2257 0.00658571
R8112 VSS.n5223 VSS.n2257 0.00658571
R8113 VSS.n5223 VSS.n5222 0.00658571
R8114 VSS.n5222 VSS.n5221 0.00658571
R8115 VSS.n5221 VSS.n2261 0.00658571
R8116 VSS.n5215 VSS.n2261 0.00658571
R8117 VSS.n5215 VSS.n5214 0.00658571
R8118 VSS.n5214 VSS.n5213 0.00658571
R8119 VSS.n5213 VSS.n2265 0.00658571
R8120 VSS.n5207 VSS.n2265 0.00658571
R8121 VSS.n5207 VSS.n5206 0.00658571
R8122 VSS.n5206 VSS.n5205 0.00658571
R8123 VSS.n5205 VSS.n2269 0.00658571
R8124 VSS.n5199 VSS.n2269 0.00658571
R8125 VSS.n5199 VSS.n5198 0.00658571
R8126 VSS.n5198 VSS.n5197 0.00658571
R8127 VSS.n5197 VSS.n5186 0.00658571
R8128 VSS.n5191 VSS.n5186 0.00658571
R8129 VSS.n5191 VSS.n5190 0.00658571
R8130 VSS.n4067 VSS.n4065 0.00658108
R8131 VSS.n3833 VSS.n3822 0.00658108
R8132 VSS.n1622 VSS.n1618 0.00654286
R8133 VSS.n2047 VSS.n1623 0.00654286
R8134 VSS.n2046 VSS.n1624 0.00654286
R8135 VSS.n1633 VSS.n1632 0.00654286
R8136 VSS.n2038 VSS.n2037 0.00654286
R8137 VSS.n1640 VSS.n1634 0.00654286
R8138 VSS.n2031 VSS.n1643 0.00654286
R8139 VSS.n425 VSS.n319 0.0065
R8140 VSS.n953 VSS.n952 0.0065
R8141 VSS.n379 VSS.n378 0.0065
R8142 VSS.n713 VSS.n320 0.0065
R8143 VSS.n1105 VSS.n98 0.0065
R8144 VSS.n490 VSS.n320 0.0065
R8145 VSS.n378 VSS.n376 0.0065
R8146 VSS.n136 VSS.n131 0.0065
R8147 VSS.n291 VSS.n136 0.0065
R8148 VSS.n1105 VSS.n1104 0.0065
R8149 VSS.n579 VSS.n372 0.0065
R8150 VSS.n743 VSS.n319 0.0065
R8151 VSS.n952 VSS.n133 0.0065
R8152 VSS.n1108 VSS.n93 0.0065
R8153 VSS.n1108 VSS.n94 0.0065
R8154 VSS.n579 VSS.n578 0.0065
R8155 VSS.n3163 VSS.n2829 0.0065
R8156 VSS.n4922 VSS.n2376 0.0065
R8157 VSS.n3130 VSS.n2832 0.0065
R8158 VSS.n4905 VSS.n2384 0.0065
R8159 VSS VSS.n5720 0.00641429
R8160 VSS.n3360 VSS 0.00641429
R8161 VSS.n1829 DVSS 0.00641429
R8162 VSS.n571 VSS.n570 0.00640498
R8163 VSS.n4191 VSS.n4190 0.00635
R8164 VSS.n3641 VSS.n3638 0.00635
R8165 VSS.n3651 VSS.n3625 0.00635
R8166 VSS.n3673 VSS.n3625 0.00635
R8167 VSS.n5069 VSS.n5068 0.00626355
R8168 VSS.n5061 VSS.n5060 0.00626355
R8169 VSS.n4438 VSS.n2613 0.006125
R8170 VSS.n4334 VSS.n2606 0.006125
R8171 VSS.n4526 VSS.n2547 0.00609286
R8172 VSS VSS.n3372 0.00609286
R8173 VSS VSS.n0 0.00609286
R8174 VSS.n2065 VSS.n1603 0.00602857
R8175 VSS.n2062 VSS.n2061 0.00602857
R8176 VSS.n1617 VSS.n1597 0.00602857
R8177 VSS.n3104 VSS.n3103 0.006
R8178 VSS.n4963 VSS.n2364 0.006
R8179 VSS.n3063 VSS.n2858 0.006
R8180 VSS.n4973 VSS.n2356 0.006
R8181 VSS.n5705 VSS.n18 0.0059878
R8182 VSS.n5702 VSS.n31 0.0059878
R8183 VSS.n1888 VSS.n1762 0.00596429
R8184 VSS.n1767 VSS.n1766 0.00596429
R8185 VSS.n1882 VSS.n1881 0.00596429
R8186 VSS.n1776 VSS.n1768 0.00596429
R8187 VSS.n1873 VSS.n1777 0.00596429
R8188 VSS.n1872 VSS.n1778 0.00596429
R8189 VSS.n1787 VSS.n1784 0.00596429
R8190 VSS.n3588 VSS.n3587 0.00583571
R8191 VSS.n3568 VSS.n2724 0.00570714
R8192 VSS.n3860 VSS.n2563 0.00561229
R8193 VSS.n2567 VSS.n2557 0.00561229
R8194 VSS.n3098 DVSS 0.00559852
R8195 DVSS VSS.n3057 0.00559852
R8196 VSS.n3243 VSS.n3242 0.00559852
R8197 VSS.n5693 VSS.n1171 0.00559091
R8198 VSS.n3818 VSS.n3731 0.00551429
R8199 VSS.n3814 VSS.n3733 0.00551429
R8200 VSS.n3788 VSS.n3730 0.00551429
R8201 VSS.n3051 VSS.n3050 0.0055
R8202 VSS.n5021 VSS.n2332 0.0055
R8203 VSS.n3054 VSS.n3053 0.0055
R8204 VSS.n5013 VSS.n2337 0.0055
R8205 VSS.n3364 VSS.n3363 0.00548841
R8206 VSS.n2763 VSS.n2762 0.00548841
R8207 VSS.n1833 VSS.n1832 0.00548841
R8208 VSS.n5 VSS.n4 0.00548841
R8209 VSS.n4118 VSS.n3891 0.00538571
R8210 VSS.n4114 VSS.n4113 0.00538571
R8211 VSS.n3899 VSS.n3887 0.00538571
R8212 VSS.n3122 VSS.n3121 0.00537685
R8213 VSS.n3128 VSS.n2845 0.00537685
R8214 VSS.n1880 VSS.n1769 0.00532927
R8215 VSS.n1874 VSS.n1775 0.00532927
R8216 VSS.n1917 VSS.n1727 0.00532927
R8217 VSS.n1901 VSS.n1900 0.00532927
R8218 VSS.n1955 VSS.n1703 0.00532927
R8219 VSS.n1939 VSS.n1938 0.00532927
R8220 VSS.n1736 VSS.n1677 0.00532927
R8221 VSS.n1977 VSS.n1976 0.00532927
R8222 VSS.n1730 VSS.n1650 0.00532927
R8223 VSS.n2009 VSS.n2008 0.00532927
R8224 VSS.n2045 VSS.n1625 0.00532927
R8225 VSS.n2039 VSS.n1631 0.00532927
R8226 VSS.n2639 VSS.n2546 0.00519286
R8227 VSS.n5250 VSS.n2243 0.00519286
R8228 VSS.n3262 VSS.n3261 0.00519286
R8229 VSS.n3859 VSS.n3858 0.00514674
R8230 VSS.n1169 VSS.n15 0.00505741
R8231 VSS.n15 VSS.n12 0.00505741
R8232 VSS.n1591 VSS.n1294 0.00505741
R8233 VSS.n1294 VSS.n1292 0.00505741
R8234 VSS.n3925 VSS.n3773 0.00504128
R8235 VSS.n4148 VSS.n3745 0.00504128
R8236 VSS.n2992 VSS.n2991 0.005
R8237 VSS.n2997 VSS.n2996 0.005
R8238 VSS.n5073 VSS.n2302 0.005
R8239 VSS.n5092 VSS.n2300 0.005
R8240 VSS.n2961 VSS.n2907 0.005
R8241 VSS.n3000 VSS.n2999 0.005
R8242 VSS.n5056 VSS.n2310 0.005
R8243 VSS.n5053 VSS.n5052 0.005
R8244 VSS.n915 VSS.n914 0.00498878
R8245 VSS.n1171 VSS.n1170 0.0049789
R8246 VSS.n1172 VSS.n1171 0.0049789
R8247 VSS.n2643 VSS.n2546 0.00493571
R8248 VSS.n5250 VSS.n5249 0.00493571
R8249 VSS.n3261 VSS.n2790 0.00493571
R8250 VSS.n3853 VSS.n2559 0.00489894
R8251 VSS.n3849 VSS.n2565 0.00489894
R8252 VSS.n4534 VSS.n2545 0.00476
R8253 VSS.n4534 VSS.n2543 0.00476
R8254 VSS.n4538 VSS.n2543 0.00476
R8255 VSS.n4538 VSS.n2541 0.00476
R8256 VSS.n4542 VSS.n2541 0.00476
R8257 VSS.n4542 VSS.n2539 0.00476
R8258 VSS.n4547 VSS.n2539 0.00476
R8259 VSS.n4547 VSS.n2537 0.00476
R8260 VSS.n4551 VSS.n2537 0.00476
R8261 VSS.n4551 VSS.n2535 0.00476
R8262 VSS.n4555 VSS.n2535 0.00476
R8263 VSS.n4555 VSS.n2533 0.00476
R8264 VSS.n4662 VSS.n2533 0.00476
R8265 VSS.n4662 VSS.n4661 0.00476
R8266 VSS.n4661 VSS.n4660 0.00476
R8267 VSS.n4660 VSS.n4561 0.00476
R8268 VSS.n4656 VSS.n4561 0.00476
R8269 VSS.n4656 VSS.n4655 0.00476
R8270 VSS.n4655 VSS.n4654 0.00476
R8271 VSS.n4654 VSS.n4567 0.00476
R8272 VSS.n4650 VSS.n4567 0.00476
R8273 VSS.n4650 VSS.n4649 0.00476
R8274 VSS.n4649 VSS.n4648 0.00476
R8275 VSS.n4648 VSS.n4573 0.00476
R8276 VSS.n4644 VSS.n4573 0.00476
R8277 VSS.n4644 VSS.n4643 0.00476
R8278 VSS.n4643 VSS.n4642 0.00476
R8279 VSS.n4642 VSS.n4580 0.00476
R8280 VSS.n4638 VSS.n4580 0.00476
R8281 VSS.n4638 VSS.n4637 0.00476
R8282 VSS.n4637 VSS.n4636 0.00476
R8283 VSS.n4636 VSS.n4586 0.00476
R8284 VSS.n4632 VSS.n4586 0.00476
R8285 VSS.n4632 VSS.n4631 0.00476
R8286 VSS.n4631 VSS.n4630 0.00476
R8287 VSS.n4630 VSS.n4592 0.00476
R8288 VSS.n4626 VSS.n4592 0.00476
R8289 VSS.n4626 VSS.n4625 0.00476
R8290 VSS.n4625 VSS.n4624 0.00476
R8291 VSS.n4624 VSS.n4598 0.00476
R8292 VSS.n4620 VSS.n4598 0.00476
R8293 VSS.n4620 VSS.n4619 0.00476
R8294 VSS.n4619 VSS.n4618 0.00476
R8295 VSS.n4618 VSS.n4604 0.00476
R8296 VSS.n4614 VSS.n4604 0.00476
R8297 VSS.n4614 VSS.n4613 0.00476
R8298 VSS.n4613 VSS.n4612 0.00476
R8299 VSS.n4612 VSS.n2116 0.00476
R8300 VSS.n5399 VSS.n2116 0.00476
R8301 VSS.n5399 VSS.n5398 0.00476
R8302 VSS.n5398 VSS.n5397 0.00476
R8303 VSS.n5397 VSS.n2120 0.00476
R8304 VSS.n5393 VSS.n2120 0.00476
R8305 VSS.n5393 VSS.n5392 0.00476
R8306 VSS.n5392 VSS.n5391 0.00476
R8307 VSS.n5391 VSS.n2126 0.00476
R8308 VSS.n5386 VSS.n2126 0.00476
R8309 VSS.n5386 VSS.n5385 0.00476
R8310 VSS.n5385 VSS.n5384 0.00476
R8311 VSS.n5384 VSS.n2133 0.00476
R8312 VSS.n5380 VSS.n2133 0.00476
R8313 VSS.n5380 VSS.n5379 0.00476
R8314 VSS.n5379 VSS.n2138 0.00476
R8315 VSS.n5375 VSS.n2138 0.00476
R8316 VSS.n5375 VSS.n5374 0.00476
R8317 VSS.n5374 VSS.n5373 0.00476
R8318 VSS.n5373 VSS.n2144 0.00476
R8319 VSS.n5369 VSS.n2144 0.00476
R8320 VSS.n5369 VSS.n5368 0.00476
R8321 VSS.n5368 VSS.n5367 0.00476
R8322 VSS.n5367 VSS.n2150 0.00476
R8323 VSS.n5363 VSS.n2150 0.00476
R8324 VSS.n5363 VSS.n5362 0.00476
R8325 VSS.n5362 VSS.n5361 0.00476
R8326 VSS.n5361 VSS.n2156 0.00476
R8327 VSS.n5357 VSS.n2156 0.00476
R8328 VSS.n5357 VSS.n5356 0.00476
R8329 VSS.n5355 VSS.n2162 0.00476
R8330 VSS.n2170 VSS.n2162 0.00476
R8331 VSS.n2170 VSS.n2169 0.00476
R8332 VSS.n576 VSS.n575 0.00476
R8333 VSS.n575 VSS.n390 0.00476
R8334 VSS.n521 VSS.n390 0.00476
R8335 VSS.n521 VSS.n520 0.00476
R8336 VSS.n520 VSS.n519 0.00476
R8337 VSS.n519 VSS.n396 0.00476
R8338 VSS.n515 VSS.n396 0.00476
R8339 VSS.n515 VSS.n514 0.00476
R8340 VSS.n514 VSS.n513 0.00476
R8341 VSS.n513 VSS.n402 0.00476
R8342 VSS.n509 VSS.n402 0.00476
R8343 VSS.n509 VSS.n508 0.00476
R8344 VSS.n508 VSS.n507 0.00476
R8345 VSS.n507 VSS.n408 0.00476
R8346 VSS.n503 VSS.n408 0.00476
R8347 VSS.n503 VSS.n502 0.00476
R8348 VSS.n502 VSS.n501 0.00476
R8349 VSS.n501 VSS.n414 0.00476
R8350 VSS.n497 VSS.n414 0.00476
R8351 VSS.n497 VSS.n496 0.00476
R8352 VSS.n496 VSS.n418 0.00476
R8353 VSS.n492 VSS.n418 0.00476
R8354 VSS.n492 VSS.n491 0.00476
R8355 VSS.n489 VSS.n424 0.00476
R8356 VSS.n485 VSS.n424 0.00476
R8357 VSS.n485 VSS.n484 0.00476
R8358 VSS.n484 VSS.n483 0.00476
R8359 VSS.n483 VSS.n431 0.00476
R8360 VSS.n479 VSS.n431 0.00476
R8361 VSS.n479 VSS.n478 0.00476
R8362 VSS.n478 VSS.n477 0.00476
R8363 VSS.n477 VSS.n437 0.00476
R8364 VSS.n473 VSS.n437 0.00476
R8365 VSS.n473 VSS.n472 0.00476
R8366 VSS.n472 VSS.n471 0.00476
R8367 VSS.n471 VSS.n443 0.00476
R8368 VSS.n467 VSS.n443 0.00476
R8369 VSS.n467 VSS.n466 0.00476
R8370 VSS.n466 VSS.n465 0.00476
R8371 VSS.n465 VSS.n449 0.00476
R8372 VSS.n461 VSS.n449 0.00476
R8373 VSS.n461 VSS.n460 0.00476
R8374 VSS.n460 VSS.n459 0.00476
R8375 VSS.n459 VSS.n456 0.00476
R8376 VSS.n456 VSS.n130 0.00476
R8377 VSS.n955 VSS.n130 0.00476
R8378 VSS.n960 VSS.n127 0.00476
R8379 VSS.n960 VSS.n125 0.00476
R8380 VSS.n965 VSS.n125 0.00476
R8381 VSS.n965 VSS.n123 0.00476
R8382 VSS.n969 VSS.n123 0.00476
R8383 VSS.n969 VSS.n121 0.00476
R8384 VSS.n973 VSS.n121 0.00476
R8385 VSS.n973 VSS.n119 0.00476
R8386 VSS.n977 VSS.n119 0.00476
R8387 VSS.n977 VSS.n117 0.00476
R8388 VSS.n981 VSS.n117 0.00476
R8389 VSS.n981 VSS.n115 0.00476
R8390 VSS.n985 VSS.n115 0.00476
R8391 VSS.n985 VSS.n113 0.00476
R8392 VSS.n989 VSS.n113 0.00476
R8393 VSS.n989 VSS.n111 0.00476
R8394 VSS.n993 VSS.n111 0.00476
R8395 VSS.n993 VSS.n109 0.00476
R8396 VSS.n997 VSS.n109 0.00476
R8397 VSS.n997 VSS.n107 0.00476
R8398 VSS.n1001 VSS.n107 0.00476
R8399 VSS.n1001 VSS.n102 0.00476
R8400 VSS.n1008 VSS.n102 0.00476
R8401 VSS.n1052 VSS.n1011 0.00476
R8402 VSS.n1048 VSS.n1011 0.00476
R8403 VSS.n1048 VSS.n1047 0.00476
R8404 VSS.n1047 VSS.n1046 0.00476
R8405 VSS.n1046 VSS.n1016 0.00476
R8406 VSS.n1042 VSS.n1016 0.00476
R8407 VSS.n1042 VSS.n1041 0.00476
R8408 VSS.n1041 VSS.n1040 0.00476
R8409 VSS.n1040 VSS.n1022 0.00476
R8410 VSS.n1036 VSS.n1022 0.00476
R8411 VSS.n1035 VSS.n1026 0.00476
R8412 VSS.n1031 VSS.n1026 0.00476
R8413 VSS.n1031 VSS.n1030 0.00476
R8414 VSS.n583 VSS.n371 0.00476
R8415 VSS.n583 VSS.n369 0.00476
R8416 VSS.n628 VSS.n369 0.00476
R8417 VSS.n628 VSS.n627 0.00476
R8418 VSS.n627 VSS.n626 0.00476
R8419 VSS.n626 VSS.n589 0.00476
R8420 VSS.n622 VSS.n589 0.00476
R8421 VSS.n622 VSS.n621 0.00476
R8422 VSS.n621 VSS.n620 0.00476
R8423 VSS.n620 VSS.n595 0.00476
R8424 VSS.n616 VSS.n595 0.00476
R8425 VSS.n616 VSS.n615 0.00476
R8426 VSS.n615 VSS.n614 0.00476
R8427 VSS.n614 VSS.n601 0.00476
R8428 VSS.n610 VSS.n601 0.00476
R8429 VSS.n610 VSS.n609 0.00476
R8430 VSS.n609 VSS.n608 0.00476
R8431 VSS.n608 VSS.n328 0.00476
R8432 VSS.n754 VSS.n328 0.00476
R8433 VSS.n754 VSS.n326 0.00476
R8434 VSS.n758 VSS.n326 0.00476
R8435 VSS.n758 VSS.n324 0.00476
R8436 VSS.n762 VSS.n324 0.00476
R8437 VSS.n766 VSS.n318 0.00476
R8438 VSS.n770 VSS.n318 0.00476
R8439 VSS.n770 VSS.n316 0.00476
R8440 VSS.n774 VSS.n316 0.00476
R8441 VSS.n774 VSS.n314 0.00476
R8442 VSS.n778 VSS.n314 0.00476
R8443 VSS.n778 VSS.n312 0.00476
R8444 VSS.n782 VSS.n312 0.00476
R8445 VSS.n782 VSS.n310 0.00476
R8446 VSS.n786 VSS.n310 0.00476
R8447 VSS.n786 VSS.n308 0.00476
R8448 VSS.n821 VSS.n308 0.00476
R8449 VSS.n821 VSS.n820 0.00476
R8450 VSS.n820 VSS.n819 0.00476
R8451 VSS.n819 VSS.n792 0.00476
R8452 VSS.n815 VSS.n792 0.00476
R8453 VSS.n815 VSS.n814 0.00476
R8454 VSS.n814 VSS.n813 0.00476
R8455 VSS.n813 VSS.n798 0.00476
R8456 VSS.n809 VSS.n798 0.00476
R8457 VSS.n809 VSS.n808 0.00476
R8458 VSS.n808 VSS.n807 0.00476
R8459 VSS.n807 VSS.n805 0.00476
R8460 VSS.n950 VSS.n949 0.00476
R8461 VSS.n949 VSS.n948 0.00476
R8462 VSS.n948 VSS.n140 0.00476
R8463 VSS.n944 VSS.n140 0.00476
R8464 VSS.n944 VSS.n943 0.00476
R8465 VSS.n943 VSS.n145 0.00476
R8466 VSS.n939 VSS.n145 0.00476
R8467 VSS.n939 VSS.n938 0.00476
R8468 VSS.n938 VSS.n937 0.00476
R8469 VSS.n937 VSS.n151 0.00476
R8470 VSS.n933 VSS.n151 0.00476
R8471 VSS.n933 VSS.n932 0.00476
R8472 VSS.n932 VSS.n931 0.00476
R8473 VSS.n931 VSS.n157 0.00476
R8474 VSS.n927 VSS.n157 0.00476
R8475 VSS.n927 VSS.n926 0.00476
R8476 VSS.n926 VSS.n925 0.00476
R8477 VSS.n925 VSS.n163 0.00476
R8478 VSS.n921 VSS.n163 0.00476
R8479 VSS.n921 VSS.n920 0.00476
R8480 VSS.n920 VSS.n919 0.00476
R8481 VSS.n919 VSS.n96 0.00476
R8482 VSS.n1106 VSS.n96 0.00476
R8483 VSS.n1111 VSS.n92 0.00476
R8484 VSS.n1111 VSS.n90 0.00476
R8485 VSS.n1115 VSS.n90 0.00476
R8486 VSS.n1115 VSS.n88 0.00476
R8487 VSS.n1119 VSS.n88 0.00476
R8488 VSS.n1119 VSS.n86 0.00476
R8489 VSS.n1123 VSS.n86 0.00476
R8490 VSS.n1123 VSS.n84 0.00476
R8491 VSS.n1127 VSS.n84 0.00476
R8492 VSS.n1127 VSS.n82 0.00476
R8493 VSS.n1131 VSS.n82 0.00476
R8494 VSS.n1135 VSS.n80 0.00476
R8495 VSS.n1135 VSS.n78 0.00476
R8496 VSS.n383 VSS.n351 0.00476
R8497 VSS.n672 VSS.n351 0.00476
R8498 VSS.n672 VSS.n349 0.00476
R8499 VSS.n676 VSS.n349 0.00476
R8500 VSS.n676 VSS.n347 0.00476
R8501 VSS.n680 VSS.n347 0.00476
R8502 VSS.n680 VSS.n345 0.00476
R8503 VSS.n684 VSS.n345 0.00476
R8504 VSS.n684 VSS.n343 0.00476
R8505 VSS.n688 VSS.n343 0.00476
R8506 VSS.n688 VSS.n341 0.00476
R8507 VSS.n692 VSS.n341 0.00476
R8508 VSS.n692 VSS.n339 0.00476
R8509 VSS.n696 VSS.n339 0.00476
R8510 VSS.n696 VSS.n337 0.00476
R8511 VSS.n700 VSS.n337 0.00476
R8512 VSS.n700 VSS.n335 0.00476
R8513 VSS.n704 VSS.n335 0.00476
R8514 VSS.n704 VSS.n333 0.00476
R8515 VSS.n748 VSS.n333 0.00476
R8516 VSS.n748 VSS.n747 0.00476
R8517 VSS.n747 VSS.n746 0.00476
R8518 VSS.n746 VSS.n711 0.00476
R8519 VSS.n741 VSS.n740 0.00476
R8520 VSS.n740 VSS.n739 0.00476
R8521 VSS.n739 VSS.n717 0.00476
R8522 VSS.n735 VSS.n717 0.00476
R8523 VSS.n735 VSS.n734 0.00476
R8524 VSS.n734 VSS.n733 0.00476
R8525 VSS.n733 VSS.n723 0.00476
R8526 VSS.n729 VSS.n723 0.00476
R8527 VSS.n729 VSS.n728 0.00476
R8528 VSS.n728 VSS.n303 0.00476
R8529 VSS.n827 VSS.n303 0.00476
R8530 VSS.n827 VSS.n301 0.00476
R8531 VSS.n831 VSS.n301 0.00476
R8532 VSS.n831 VSS.n299 0.00476
R8533 VSS.n835 VSS.n299 0.00476
R8534 VSS.n835 VSS.n297 0.00476
R8535 VSS.n839 VSS.n297 0.00476
R8536 VSS.n839 VSS.n295 0.00476
R8537 VSS.n843 VSS.n295 0.00476
R8538 VSS.n843 VSS.n293 0.00476
R8539 VSS.n847 VSS.n293 0.00476
R8540 VSS.n847 VSS.n290 0.00476
R8541 VSS.n851 VSS.n290 0.00476
R8542 VSS.n856 VSS.n288 0.00476
R8543 VSS.n856 VSS.n286 0.00476
R8544 VSS.n861 VSS.n286 0.00476
R8545 VSS.n861 VSS.n284 0.00476
R8546 VSS.n865 VSS.n284 0.00476
R8547 VSS.n865 VSS.n281 0.00476
R8548 VSS.n869 VSS.n281 0.00476
R8549 VSS.n869 VSS.n279 0.00476
R8550 VSS.n873 VSS.n279 0.00476
R8551 VSS.n873 VSS.n277 0.00476
R8552 VSS.n877 VSS.n277 0.00476
R8553 VSS.n877 VSS.n275 0.00476
R8554 VSS.n881 VSS.n275 0.00476
R8555 VSS.n881 VSS.n273 0.00476
R8556 VSS.n885 VSS.n273 0.00476
R8557 VSS.n885 VSS.n271 0.00476
R8558 VSS.n889 VSS.n271 0.00476
R8559 VSS.n889 VSS.n269 0.00476
R8560 VSS.n893 VSS.n269 0.00476
R8561 VSS.n893 VSS.n267 0.00476
R8562 VSS.n899 VSS.n267 0.00476
R8563 VSS.n899 VSS.n898 0.00476
R8564 VSS.n898 VSS.n99 0.00476
R8565 VSS.n1103 VSS.n1058 0.00476
R8566 VSS.n1099 VSS.n1058 0.00476
R8567 VSS.n1099 VSS.n1098 0.00476
R8568 VSS.n1098 VSS.n1097 0.00476
R8569 VSS.n1097 VSS.n1064 0.00476
R8570 VSS.n1093 VSS.n1064 0.00476
R8571 VSS.n1093 VSS.n1092 0.00476
R8572 VSS.n1092 VSS.n1091 0.00476
R8573 VSS.n1091 VSS.n1070 0.00476
R8574 VSS.n1087 VSS.n1070 0.00476
R8575 VSS.n1086 VSS.n1074 0.00476
R8576 VSS.n1082 VSS.n1074 0.00476
R8577 VSS.n1082 VSS.n1081 0.00476
R8578 VSS.n671 VSS.n352 0.00476
R8579 VSS.n677 VSS.n348 0.00476
R8580 VSS.n678 VSS.n677 0.00476
R8581 VSS.n679 VSS.n678 0.00476
R8582 VSS.n679 VSS.n344 0.00476
R8583 VSS.n685 VSS.n344 0.00476
R8584 VSS.n686 VSS.n685 0.00476
R8585 VSS.n687 VSS.n686 0.00476
R8586 VSS.n687 VSS.n340 0.00476
R8587 VSS.n693 VSS.n340 0.00476
R8588 VSS.n694 VSS.n693 0.00476
R8589 VSS.n695 VSS.n694 0.00476
R8590 VSS.n695 VSS.n336 0.00476
R8591 VSS.n701 VSS.n336 0.00476
R8592 VSS.n702 VSS.n701 0.00476
R8593 VSS.n703 VSS.n702 0.00476
R8594 VSS.n703 VSS.n331 0.00476
R8595 VSS.n749 VSS.n332 0.00476
R8596 VSS.n745 VSS.n332 0.00476
R8597 VSS.n745 VSS.n744 0.00476
R8598 VSS.n742 VSS.n712 0.00476
R8599 VSS.n738 VSS.n712 0.00476
R8600 VSS.n738 VSS.n737 0.00476
R8601 VSS.n737 VSS.n736 0.00476
R8602 VSS.n736 VSS.n718 0.00476
R8603 VSS.n732 VSS.n718 0.00476
R8604 VSS.n732 VSS.n731 0.00476
R8605 VSS.n731 VSS.n730 0.00476
R8606 VSS.n730 VSS.n724 0.00476
R8607 VSS.n724 VSS.n304 0.00476
R8608 VSS.n826 VSS.n304 0.00476
R8609 VSS.n832 VSS.n300 0.00476
R8610 VSS.n833 VSS.n832 0.00476
R8611 VSS.n834 VSS.n833 0.00476
R8612 VSS.n834 VSS.n296 0.00476
R8613 VSS.n840 VSS.n296 0.00476
R8614 VSS.n841 VSS.n840 0.00476
R8615 VSS.n842 VSS.n841 0.00476
R8616 VSS.n842 VSS.n292 0.00476
R8617 VSS.n848 VSS.n292 0.00476
R8618 VSS.n849 VSS.n848 0.00476
R8619 VSS.n850 VSS.n849 0.00476
R8620 VSS.n857 VSS.n287 0.00476
R8621 VSS.n858 VSS.n857 0.00476
R8622 VSS.n860 VSS.n858 0.00476
R8623 VSS.n860 VSS.n859 0.00476
R8624 VSS.n867 VSS.n866 0.00476
R8625 VSS.n868 VSS.n867 0.00476
R8626 VSS.n868 VSS.n278 0.00476
R8627 VSS.n874 VSS.n278 0.00476
R8628 VSS.n875 VSS.n874 0.00476
R8629 VSS.n876 VSS.n875 0.00476
R8630 VSS.n876 VSS.n274 0.00476
R8631 VSS.n882 VSS.n274 0.00476
R8632 VSS.n883 VSS.n882 0.00476
R8633 VSS.n884 VSS.n883 0.00476
R8634 VSS.n884 VSS.n270 0.00476
R8635 VSS.n890 VSS.n270 0.00476
R8636 VSS.n891 VSS.n890 0.00476
R8637 VSS.n892 VSS.n891 0.00476
R8638 VSS.n892 VSS.n263 0.00476
R8639 VSS.n900 VSS.n266 0.00476
R8640 VSS.n1102 VSS.n1101 0.00476
R8641 VSS.n1101 VSS.n1100 0.00476
R8642 VSS.n1100 VSS.n1059 0.00476
R8643 VSS.n1096 VSS.n1059 0.00476
R8644 VSS.n1096 VSS.n1095 0.00476
R8645 VSS.n1095 VSS.n1094 0.00476
R8646 VSS.n1094 VSS.n1065 0.00476
R8647 VSS.n1090 VSS.n1065 0.00476
R8648 VSS.n1090 VSS.n1089 0.00476
R8649 VSS.n1089 VSS.n1088 0.00476
R8650 VSS.n1085 VSS.n1084 0.00476
R8651 VSS.n1084 VSS.n1083 0.00476
R8652 VSS.n1083 VSS.n1075 0.00476
R8653 VSS.n582 VSS.n367 0.00476
R8654 VSS.n629 VSS.n368 0.00476
R8655 VSS.n625 VSS.n368 0.00476
R8656 VSS.n625 VSS.n624 0.00476
R8657 VSS.n624 VSS.n623 0.00476
R8658 VSS.n623 VSS.n590 0.00476
R8659 VSS.n619 VSS.n590 0.00476
R8660 VSS.n619 VSS.n618 0.00476
R8661 VSS.n618 VSS.n617 0.00476
R8662 VSS.n617 VSS.n596 0.00476
R8663 VSS.n613 VSS.n596 0.00476
R8664 VSS.n613 VSS.n612 0.00476
R8665 VSS.n612 VSS.n611 0.00476
R8666 VSS.n611 VSS.n602 0.00476
R8667 VSS.n607 VSS.n602 0.00476
R8668 VSS.n607 VSS.n329 0.00476
R8669 VSS.n753 VSS.n329 0.00476
R8670 VSS.n759 VSS.n325 0.00476
R8671 VSS.n760 VSS.n759 0.00476
R8672 VSS.n761 VSS.n760 0.00476
R8673 VSS.n768 VSS.n767 0.00476
R8674 VSS.n769 VSS.n768 0.00476
R8675 VSS.n769 VSS.n315 0.00476
R8676 VSS.n775 VSS.n315 0.00476
R8677 VSS.n776 VSS.n775 0.00476
R8678 VSS.n777 VSS.n776 0.00476
R8679 VSS.n777 VSS.n311 0.00476
R8680 VSS.n783 VSS.n311 0.00476
R8681 VSS.n784 VSS.n783 0.00476
R8682 VSS.n785 VSS.n784 0.00476
R8683 VSS.n785 VSS.n306 0.00476
R8684 VSS.n822 VSS.n307 0.00476
R8685 VSS.n818 VSS.n307 0.00476
R8686 VSS.n818 VSS.n817 0.00476
R8687 VSS.n817 VSS.n816 0.00476
R8688 VSS.n816 VSS.n793 0.00476
R8689 VSS.n812 VSS.n793 0.00476
R8690 VSS.n812 VSS.n811 0.00476
R8691 VSS.n811 VSS.n810 0.00476
R8692 VSS.n810 VSS.n799 0.00476
R8693 VSS.n806 VSS.n799 0.00476
R8694 VSS.n806 VSS.n134 0.00476
R8695 VSS.n951 VSS.n135 0.00476
R8696 VSS.n947 VSS.n135 0.00476
R8697 VSS.n947 VSS.n946 0.00476
R8698 VSS.n946 VSS.n945 0.00476
R8699 VSS.n942 VSS.n941 0.00476
R8700 VSS.n941 VSS.n940 0.00476
R8701 VSS.n940 VSS.n146 0.00476
R8702 VSS.n936 VSS.n146 0.00476
R8703 VSS.n936 VSS.n935 0.00476
R8704 VSS.n935 VSS.n934 0.00476
R8705 VSS.n934 VSS.n152 0.00476
R8706 VSS.n930 VSS.n152 0.00476
R8707 VSS.n930 VSS.n929 0.00476
R8708 VSS.n929 VSS.n928 0.00476
R8709 VSS.n928 VSS.n158 0.00476
R8710 VSS.n924 VSS.n158 0.00476
R8711 VSS.n924 VSS.n923 0.00476
R8712 VSS.n923 VSS.n922 0.00476
R8713 VSS.n922 VSS.n164 0.00476
R8714 VSS.n918 VSS.n917 0.00476
R8715 VSS.n1110 VSS.n1109 0.00476
R8716 VSS.n1110 VSS.n89 0.00476
R8717 VSS.n1116 VSS.n89 0.00476
R8718 VSS.n1117 VSS.n1116 0.00476
R8719 VSS.n1118 VSS.n1117 0.00476
R8720 VSS.n1118 VSS.n85 0.00476
R8721 VSS.n1124 VSS.n85 0.00476
R8722 VSS.n1125 VSS.n1124 0.00476
R8723 VSS.n1126 VSS.n1125 0.00476
R8724 VSS.n1126 VSS.n81 0.00476
R8725 VSS.n1132 VSS.n81 0.00476
R8726 VSS.n1134 VSS.n1133 0.00476
R8727 VSS.n1134 VSS.n57 0.00476
R8728 VSS.n574 VSS.n573 0.00476
R8729 VSS.n522 VSS.n391 0.00476
R8730 VSS.n518 VSS.n391 0.00476
R8731 VSS.n518 VSS.n517 0.00476
R8732 VSS.n517 VSS.n516 0.00476
R8733 VSS.n516 VSS.n397 0.00476
R8734 VSS.n512 VSS.n397 0.00476
R8735 VSS.n512 VSS.n511 0.00476
R8736 VSS.n511 VSS.n510 0.00476
R8737 VSS.n510 VSS.n403 0.00476
R8738 VSS.n506 VSS.n403 0.00476
R8739 VSS.n506 VSS.n505 0.00476
R8740 VSS.n505 VSS.n504 0.00476
R8741 VSS.n504 VSS.n409 0.00476
R8742 VSS.n500 VSS.n409 0.00476
R8743 VSS.n500 VSS.n499 0.00476
R8744 VSS.n499 VSS.n498 0.00476
R8745 VSS.n495 VSS.n494 0.00476
R8746 VSS.n494 VSS.n493 0.00476
R8747 VSS.n493 VSS.n419 0.00476
R8748 VSS.n488 VSS.n487 0.00476
R8749 VSS.n487 VSS.n486 0.00476
R8750 VSS.n486 VSS.n426 0.00476
R8751 VSS.n482 VSS.n426 0.00476
R8752 VSS.n482 VSS.n481 0.00476
R8753 VSS.n481 VSS.n480 0.00476
R8754 VSS.n480 VSS.n432 0.00476
R8755 VSS.n476 VSS.n432 0.00476
R8756 VSS.n476 VSS.n475 0.00476
R8757 VSS.n475 VSS.n474 0.00476
R8758 VSS.n474 VSS.n438 0.00476
R8759 VSS.n470 VSS.n469 0.00476
R8760 VSS.n469 VSS.n468 0.00476
R8761 VSS.n468 VSS.n444 0.00476
R8762 VSS.n464 VSS.n444 0.00476
R8763 VSS.n464 VSS.n463 0.00476
R8764 VSS.n463 VSS.n462 0.00476
R8765 VSS.n462 VSS.n450 0.00476
R8766 VSS.n458 VSS.n450 0.00476
R8767 VSS.n458 VSS.n457 0.00476
R8768 VSS.n457 VSS.n132 0.00476
R8769 VSS.n954 VSS.n132 0.00476
R8770 VSS.n961 VSS.n126 0.00476
R8771 VSS.n962 VSS.n961 0.00476
R8772 VSS.n964 VSS.n962 0.00476
R8773 VSS.n964 VSS.n963 0.00476
R8774 VSS.n971 VSS.n970 0.00476
R8775 VSS.n972 VSS.n971 0.00476
R8776 VSS.n972 VSS.n118 0.00476
R8777 VSS.n978 VSS.n118 0.00476
R8778 VSS.n979 VSS.n978 0.00476
R8779 VSS.n980 VSS.n979 0.00476
R8780 VSS.n980 VSS.n114 0.00476
R8781 VSS.n986 VSS.n114 0.00476
R8782 VSS.n987 VSS.n986 0.00476
R8783 VSS.n988 VSS.n987 0.00476
R8784 VSS.n988 VSS.n110 0.00476
R8785 VSS.n994 VSS.n110 0.00476
R8786 VSS.n995 VSS.n994 0.00476
R8787 VSS.n996 VSS.n995 0.00476
R8788 VSS.n996 VSS.n106 0.00476
R8789 VSS.n1002 VSS.n103 0.00476
R8790 VSS.n1051 VSS.n1050 0.00476
R8791 VSS.n1050 VSS.n1049 0.00476
R8792 VSS.n1049 VSS.n1012 0.00476
R8793 VSS.n1045 VSS.n1012 0.00476
R8794 VSS.n1045 VSS.n1044 0.00476
R8795 VSS.n1044 VSS.n1043 0.00476
R8796 VSS.n1043 VSS.n1017 0.00476
R8797 VSS.n1039 VSS.n1017 0.00476
R8798 VSS.n1039 VSS.n1038 0.00476
R8799 VSS.n1038 VSS.n1037 0.00476
R8800 VSS.n1034 VSS.n1033 0.00476
R8801 VSS.n1033 VSS.n1032 0.00476
R8802 VSS.n1032 VSS.n36 0.00476
R8803 VSS.n4535 VSS.n2544 0.00476
R8804 VSS.n4536 VSS.n4535 0.00476
R8805 VSS.n4537 VSS.n4536 0.00476
R8806 VSS.n4537 VSS.n2540 0.00476
R8807 VSS.n4543 VSS.n2540 0.00476
R8808 VSS.n4546 VSS.n4545 0.00476
R8809 VSS.n4546 VSS.n2536 0.00476
R8810 VSS.n4552 VSS.n2536 0.00476
R8811 VSS.n4553 VSS.n4552 0.00476
R8812 VSS.n4554 VSS.n4553 0.00476
R8813 VSS.n4554 VSS.n2531 0.00476
R8814 VSS.n4663 VSS.n2532 0.00476
R8815 VSS.n4659 VSS.n2532 0.00476
R8816 VSS.n4659 VSS.n4658 0.00476
R8817 VSS.n4658 VSS.n4657 0.00476
R8818 VSS.n4657 VSS.n4562 0.00476
R8819 VSS.n4653 VSS.n4562 0.00476
R8820 VSS.n4653 VSS.n4652 0.00476
R8821 VSS.n4652 VSS.n4651 0.00476
R8822 VSS.n4651 VSS.n4568 0.00476
R8823 VSS.n4647 VSS.n4646 0.00476
R8824 VSS.n4646 VSS.n4645 0.00476
R8825 VSS.n4645 VSS.n4575 0.00476
R8826 VSS.n4641 VSS.n4575 0.00476
R8827 VSS.n4641 VSS.n4640 0.00476
R8828 VSS.n4640 VSS.n4639 0.00476
R8829 VSS.n4639 VSS.n4581 0.00476
R8830 VSS.n4635 VSS.n4581 0.00476
R8831 VSS.n4635 VSS.n4634 0.00476
R8832 VSS.n4634 VSS.n4633 0.00476
R8833 VSS.n4633 VSS.n4587 0.00476
R8834 VSS.n4629 VSS.n4587 0.00476
R8835 VSS.n4629 VSS.n4628 0.00476
R8836 VSS.n4628 VSS.n4627 0.00476
R8837 VSS.n4627 VSS.n4593 0.00476
R8838 VSS.n4623 VSS.n4593 0.00476
R8839 VSS.n4623 VSS.n4622 0.00476
R8840 VSS.n4622 VSS.n4621 0.00476
R8841 VSS.n4621 VSS.n4599 0.00476
R8842 VSS.n4617 VSS.n4599 0.00476
R8843 VSS.n4617 VSS.n4616 0.00476
R8844 VSS.n4616 VSS.n4615 0.00476
R8845 VSS.n4615 VSS.n4605 0.00476
R8846 VSS.n4611 VSS.n4605 0.00476
R8847 VSS.n4611 VSS.n2114 0.00476
R8848 VSS.n5400 VSS.n2115 0.00476
R8849 VSS.n5396 VSS.n2115 0.00476
R8850 VSS.n5396 VSS.n5395 0.00476
R8851 VSS.n5395 VSS.n5394 0.00476
R8852 VSS.n5394 VSS.n2121 0.00476
R8853 VSS.n5390 VSS.n2121 0.00476
R8854 VSS.n5388 VSS.n5387 0.00476
R8855 VSS.n5387 VSS.n2128 0.00476
R8856 VSS.n5383 VSS.n2128 0.00476
R8857 VSS.n5383 VSS.n5382 0.00476
R8858 VSS.n5382 VSS.n5381 0.00476
R8859 VSS.n5378 VSS.n5377 0.00476
R8860 VSS.n5377 VSS.n5376 0.00476
R8861 VSS.n5376 VSS.n2139 0.00476
R8862 VSS.n5372 VSS.n2139 0.00476
R8863 VSS.n5372 VSS.n5371 0.00476
R8864 VSS.n5371 VSS.n5370 0.00476
R8865 VSS.n5370 VSS.n2145 0.00476
R8866 VSS.n5366 VSS.n2145 0.00476
R8867 VSS.n5366 VSS.n5365 0.00476
R8868 VSS.n5365 VSS.n5364 0.00476
R8869 VSS.n5364 VSS.n2151 0.00476
R8870 VSS.n5360 VSS.n2151 0.00476
R8871 VSS.n5360 VSS.n5359 0.00476
R8872 VSS.n5359 VSS.n5358 0.00476
R8873 VSS.n5358 VSS.n2157 0.00476
R8874 VSS.n2171 VSS.n2164 0.00476
R8875 VSS.n4342 VSS.n2610 0.00465761
R8876 VSS.n4341 VSS.n2607 0.00465761
R8877 VSS.n4118 VSS.n3888 0.00461429
R8878 VSS.n4114 VSS.n3892 0.00461429
R8879 VSS.n3893 VSS.n3887 0.00461429
R8880 VSS.n913 VSS.n217 0.00461371
R8881 VSS.n1087 DVSS 0.00458
R8882 VSS.n1088 DVSS 0.00458
R8883 VSS.n632 VSS.n631 0.0045724
R8884 VSS.n764 VSS.n321 0.0045
R8885 VSS.n957 VSS.n128 0.0045
R8886 VSS.n386 VSS.n385 0.0045
R8887 VSS.n764 VSS.n322 0.0045
R8888 VSS.n853 VSS.n128 0.0045
R8889 VSS.n1055 VSS.n1054 0.0045
R8890 VSS.n1056 VSS.n1055 0.0045
R8891 VSS.n387 VSS.n386 0.0045
R8892 VSS.n2949 VSS.n2923 0.0045
R8893 VSS.n3046 VSS.n2883 0.0045
R8894 VSS.n5041 VSS.n2322 0.0045
R8895 VSS.n5111 VSS.n2290 0.0045
R8896 VSS.n2932 VSS.n2921 0.0045
R8897 VSS.n3007 VSS.n3006 0.0045
R8898 VSS.n5010 VSS.n2325 0.0045
R8899 VSS.n5118 VSS.n2284 0.0045
R8900 VSS.n3818 VSS.n3790 0.00448571
R8901 VSS.n3814 VSS.n3813 0.00448571
R8902 VSS.n3788 VSS.n3734 0.00448571
R8903 VSS.n3569 VSS.n3568 0.00442143
R8904 VSS.n633 VSS.n365 0.0044172
R8905 VSS.n382 VSS.n381 0.00434
R8906 VSS.n581 VSS.n580 0.00434
R8907 VSS.n577 VSS.n375 0.00434
R8908 VSS.n4169 VSS.n3720 0.004325
R8909 VSS.n3805 VSS.n3795 0.004325
R8910 VSS.n3587 VSS.n2709 0.00429286
R8911 VSS.n1878 VSS.n1877 0.00428827
R8912 VSS.n1915 VSS.n1746 0.00428827
R8913 VSS.n1953 VSS.n1704 0.00428827
R8914 VSS.n1740 VSS.n1739 0.00428827
R8915 VSS.n1734 VSS.n1733 0.00428827
R8916 VSS.n2043 VSS.n2042 0.00428827
R8917 VSS.n750 VSS.n749 0.00425
R8918 VSS.n752 VSS.n325 0.00425
R8919 VSS.n495 VSS.n330 0.00425
R8920 VSS.n1139 VSS.n1138 0.00422
R8921 VSS.n1142 VSS.n37 0.00422
R8922 VSS.n5401 VSS.n2114 0.00419
R8923 VSS.n2172 VSS.n2163 0.00419
R8924 VSS.n3857 VSS.n2560 0.0041856
R8925 VSS.n3846 VSS.n2566 0.0041856
R8926 VSS.n1766 VSS.n1762 0.00416429
R8927 VSS.n1882 VSS.n1767 0.00416429
R8928 VSS.n1881 VSS.n1768 0.00416429
R8929 VSS.n1777 VSS.n1776 0.00416429
R8930 VSS.n1873 VSS.n1872 0.00416429
R8931 VSS.n1784 VSS.n1778 0.00416429
R8932 VSS.n1866 VSS.n1787 0.00416429
R8933 VSS.n2062 VSS.n1603 0.0041
R8934 VSS.n2061 VSS.n1597 0.0041
R8935 VSS.n4544 VSS.n4543 0.00407
R8936 VSS.n4664 VSS.n4663 0.00407
R8937 VSS.n1052 VSS.n98 0.00404
R8938 VSS.n1105 VSS.n92 0.00404
R8939 VSS.n1104 VSS.n1103 0.00404
R8940 VSS.n1102 VSS.n94 0.00404
R8941 VSS.n1109 VSS.n1108 0.00404
R8942 VSS.n1051 VSS.n93 0.00404
R8943 VSS.n4523 VSS.n2547 0.00403571
R8944 VSS.n3099 VSS.n2860 0.004
R8945 VSS.n4984 VSS.n4983 0.004
R8946 VSS.n3068 VSS.n3067 0.004
R8947 VSS.n4976 VSS.n2352 0.004
R8948 VSS.n866 VSS.n283 0.00395
R8949 VSS.n942 VSS.n141 0.00395
R8950 VSS.n970 VSS.n122 0.00395
R8951 VSS.n5389 VSS.n5388 0.00395
R8952 VSS.n5353 VSS.n2163 0.00395
R8953 VSS.n4161 VSS.n3726 0.00393049
R8954 VSS.n4164 VSS.n4163 0.00393049
R8955 VSS.n3951 VSS.n3905 0.00393049
R8956 VSS.n3949 VSS.n3948 0.00393049
R8957 VSS.n5356 DVSS 0.00392
R8958 VSS.n1036 DVSS 0.00392
R8959 VSS.n1037 DVSS 0.00392
R8960 DVSS VSS.n2157 0.00392
R8961 VSS.n912 VSS.n911 0.00391137
R8962 VSS.n902 VSS.n262 0.00386658
R8963 VSS.n1877 VSS.n1876 0.00382908
R8964 VSS.n1899 VSS.n1746 0.00382908
R8965 VSS.n1937 VSS.n1704 0.00382908
R8966 VSS.n1740 VSS.n1687 0.00382908
R8967 VSS.n1734 VSS.n1662 0.00382908
R8968 VSS.n2042 VSS.n2041 0.00382908
R8969 VSS.n131 VSS.n127 0.0038
R8970 VSS.n950 VSS.n136 0.0038
R8971 VSS.n291 VSS.n288 0.0038
R8972 VSS.n287 VSS.n133 0.0038
R8973 VSS.n952 VSS.n951 0.0038
R8974 VSS.n953 VSS.n126 0.0038
R8975 VSS.n4647 VSS.n4574 0.0038
R8976 VSS.n3642 VSS.n3641 0.00377857
R8977 VSS.n3652 VSS.n3651 0.00377857
R8978 VSS.n3673 VSS.n3672 0.00377857
R8979 VSS.n635 VSS.n634 0.00374841
R8980 VSS.n4310 VSS.n2624 0.00362245
R8981 VSS.n4982 VSS.n4981 0.00360345
R8982 VSS.n4980 VSS.n4977 0.00360345
R8983 VSS.n901 VSS.n263 0.00359
R8984 VSS.n916 VSS.n164 0.00359
R8985 VSS.n1003 VSS.n106 0.00359
R8986 VSS.n2053 VSS.n1618 0.00358571
R8987 VSS.n1623 VSS.n1622 0.00358571
R8988 VSS.n2047 VSS.n2046 0.00358571
R8989 VSS.n1632 VSS.n1624 0.00358571
R8990 VSS.n2038 VSS.n1633 0.00358571
R8991 VSS.n2037 VSS.n1634 0.00358571
R8992 VSS.n1643 VSS.n1640 0.00358571
R8993 VSS.n490 VSS.n489 0.00356
R8994 VSS.n766 VSS.n320 0.00356
R8995 VSS.n741 VSS.n713 0.00356
R8996 VSS.n743 VSS.n742 0.00356
R8997 VSS.n767 VSS.n319 0.00356
R8998 VSS.n488 VSS.n425 0.00356
R8999 VSS.n669 VSS.n353 0.0035543
R9000 DVSS VSS.n80 0.00353
R9001 VSS.n1133 DVSS 0.00353
R9002 VSS.n3142 VSS.n2839 0.0035
R9003 VSS.n4944 VSS.n2374 0.0035
R9004 VSS.n3134 VSS.n2844 0.0035
R9005 VSS.n4902 VSS.n4901 0.0035
R9006 VSS.n1005 VSS.n1004 0.00341771
R9007 VSS.n4101 VSS.n3903 0.00338991
R9008 VSS.n1079 VSS.n1075 0.00338166
R9009 VSS.n2167 VSS.n2164 0.00338166
R9010 VSS.n4533 VSS.n2542 0.00334
R9011 VSS.n4539 VSS.n2542 0.00334
R9012 VSS.n4540 VSS.n4539 0.00334
R9013 VSS.n4541 VSS.n4540 0.00334
R9014 VSS.n4541 VSS.n2538 0.00334
R9015 VSS.n4548 VSS.n2538 0.00334
R9016 VSS.n4549 VSS.n4548 0.00334
R9017 VSS.n4550 VSS.n4549 0.00334
R9018 VSS.n4550 VSS.n2534 0.00334
R9019 VSS.n4556 VSS.n2534 0.00334
R9020 VSS.n4557 VSS.n4556 0.00334
R9021 VSS.n4558 VSS.n4557 0.00334
R9022 VSS.n4559 VSS.n4558 0.00334
R9023 VSS.n4560 VSS.n4559 0.00334
R9024 VSS.n4563 VSS.n4560 0.00334
R9025 VSS.n4564 VSS.n4563 0.00334
R9026 VSS.n4565 VSS.n4564 0.00334
R9027 VSS.n4566 VSS.n4565 0.00334
R9028 VSS.n4569 VSS.n4566 0.00334
R9029 VSS.n4570 VSS.n4569 0.00334
R9030 VSS.n4571 VSS.n4570 0.00334
R9031 VSS.n4572 VSS.n4571 0.00334
R9032 VSS.n4576 VSS.n4572 0.00334
R9033 VSS.n4577 VSS.n4576 0.00334
R9034 VSS.n4578 VSS.n4577 0.00334
R9035 VSS.n4579 VSS.n4578 0.00334
R9036 VSS.n4582 VSS.n4579 0.00334
R9037 VSS.n4583 VSS.n4582 0.00334
R9038 VSS.n4584 VSS.n4583 0.00334
R9039 VSS.n4585 VSS.n4584 0.00334
R9040 VSS.n4588 VSS.n4585 0.00334
R9041 VSS.n4589 VSS.n4588 0.00334
R9042 VSS.n4590 VSS.n4589 0.00334
R9043 VSS.n4591 VSS.n4590 0.00334
R9044 VSS.n4594 VSS.n4591 0.00334
R9045 VSS.n4595 VSS.n4594 0.00334
R9046 VSS.n4596 VSS.n4595 0.00334
R9047 VSS.n4597 VSS.n4596 0.00334
R9048 VSS.n4600 VSS.n4597 0.00334
R9049 VSS.n4601 VSS.n4600 0.00334
R9050 VSS.n4602 VSS.n4601 0.00334
R9051 VSS.n4603 VSS.n4602 0.00334
R9052 VSS.n4606 VSS.n4603 0.00334
R9053 VSS.n4607 VSS.n4606 0.00334
R9054 VSS.n4608 VSS.n4607 0.00334
R9055 VSS.n4610 VSS.n4608 0.00334
R9056 VSS.n4610 VSS.n4609 0.00334
R9057 VSS.n4609 VSS.n2117 0.00334
R9058 VSS.n2118 VSS.n2117 0.00334
R9059 VSS.n2119 VSS.n2118 0.00334
R9060 VSS.n2122 VSS.n2119 0.00334
R9061 VSS.n2123 VSS.n2122 0.00334
R9062 VSS.n2124 VSS.n2123 0.00334
R9063 VSS.n2125 VSS.n2124 0.00334
R9064 VSS.n2129 VSS.n2125 0.00334
R9065 VSS.n2130 VSS.n2129 0.00334
R9066 VSS.n2131 VSS.n2130 0.00334
R9067 VSS.n2132 VSS.n2131 0.00334
R9068 VSS.n2135 VSS.n2132 0.00334
R9069 VSS.n2136 VSS.n2135 0.00334
R9070 VSS.n2137 VSS.n2136 0.00334
R9071 VSS.n2140 VSS.n2137 0.00334
R9072 VSS.n2141 VSS.n2140 0.00334
R9073 VSS.n2142 VSS.n2141 0.00334
R9074 VSS.n2143 VSS.n2142 0.00334
R9075 VSS.n2146 VSS.n2143 0.00334
R9076 VSS.n2147 VSS.n2146 0.00334
R9077 VSS.n2148 VSS.n2147 0.00334
R9078 VSS.n2149 VSS.n2148 0.00334
R9079 VSS.n2152 VSS.n2149 0.00334
R9080 VSS.n2153 VSS.n2152 0.00334
R9081 VSS.n2154 VSS.n2153 0.00334
R9082 VSS.n2155 VSS.n2154 0.00334
R9083 VSS.n2158 VSS.n2155 0.00334
R9084 VSS.n2159 VSS.n2158 0.00334
R9085 VSS.n2160 VSS.n2159 0.00334
R9086 VSS.n2166 VSS.n2165 0.00334
R9087 VSS.n384 VSS.n350 0.00334
R9088 VSS.n673 VSS.n350 0.00334
R9089 VSS.n674 VSS.n673 0.00334
R9090 VSS.n675 VSS.n674 0.00334
R9091 VSS.n675 VSS.n346 0.00334
R9092 VSS.n681 VSS.n346 0.00334
R9093 VSS.n682 VSS.n681 0.00334
R9094 VSS.n683 VSS.n682 0.00334
R9095 VSS.n683 VSS.n342 0.00334
R9096 VSS.n689 VSS.n342 0.00334
R9097 VSS.n690 VSS.n689 0.00334
R9098 VSS.n691 VSS.n690 0.00334
R9099 VSS.n691 VSS.n338 0.00334
R9100 VSS.n697 VSS.n338 0.00334
R9101 VSS.n698 VSS.n697 0.00334
R9102 VSS.n699 VSS.n698 0.00334
R9103 VSS.n699 VSS.n334 0.00334
R9104 VSS.n705 VSS.n334 0.00334
R9105 VSS.n706 VSS.n705 0.00334
R9106 VSS.n707 VSS.n706 0.00334
R9107 VSS.n708 VSS.n707 0.00334
R9108 VSS.n709 VSS.n708 0.00334
R9109 VSS.n710 VSS.n709 0.00334
R9110 VSS.n715 VSS.n714 0.00334
R9111 VSS.n716 VSS.n715 0.00334
R9112 VSS.n719 VSS.n716 0.00334
R9113 VSS.n720 VSS.n719 0.00334
R9114 VSS.n721 VSS.n720 0.00334
R9115 VSS.n722 VSS.n721 0.00334
R9116 VSS.n725 VSS.n722 0.00334
R9117 VSS.n726 VSS.n725 0.00334
R9118 VSS.n727 VSS.n726 0.00334
R9119 VSS.n727 VSS.n302 0.00334
R9120 VSS.n828 VSS.n302 0.00334
R9121 VSS.n829 VSS.n828 0.00334
R9122 VSS.n830 VSS.n829 0.00334
R9123 VSS.n830 VSS.n298 0.00334
R9124 VSS.n836 VSS.n298 0.00334
R9125 VSS.n837 VSS.n836 0.00334
R9126 VSS.n838 VSS.n837 0.00334
R9127 VSS.n838 VSS.n294 0.00334
R9128 VSS.n844 VSS.n294 0.00334
R9129 VSS.n845 VSS.n844 0.00334
R9130 VSS.n846 VSS.n845 0.00334
R9131 VSS.n846 VSS.n289 0.00334
R9132 VSS.n852 VSS.n289 0.00334
R9133 VSS.n855 VSS.n854 0.00334
R9134 VSS.n855 VSS.n285 0.00334
R9135 VSS.n862 VSS.n285 0.00334
R9136 VSS.n863 VSS.n862 0.00334
R9137 VSS.n864 VSS.n863 0.00334
R9138 VSS.n864 VSS.n280 0.00334
R9139 VSS.n870 VSS.n280 0.00334
R9140 VSS.n871 VSS.n870 0.00334
R9141 VSS.n872 VSS.n871 0.00334
R9142 VSS.n872 VSS.n276 0.00334
R9143 VSS.n878 VSS.n276 0.00334
R9144 VSS.n879 VSS.n878 0.00334
R9145 VSS.n880 VSS.n879 0.00334
R9146 VSS.n880 VSS.n272 0.00334
R9147 VSS.n886 VSS.n272 0.00334
R9148 VSS.n887 VSS.n886 0.00334
R9149 VSS.n888 VSS.n887 0.00334
R9150 VSS.n888 VSS.n268 0.00334
R9151 VSS.n894 VSS.n268 0.00334
R9152 VSS.n895 VSS.n894 0.00334
R9153 VSS.n896 VSS.n895 0.00334
R9154 VSS.n897 VSS.n896 0.00334
R9155 VSS.n897 VSS.n100 0.00334
R9156 VSS.n1060 VSS.n1057 0.00334
R9157 VSS.n1061 VSS.n1060 0.00334
R9158 VSS.n1062 VSS.n1061 0.00334
R9159 VSS.n1063 VSS.n1062 0.00334
R9160 VSS.n1066 VSS.n1063 0.00334
R9161 VSS.n1067 VSS.n1066 0.00334
R9162 VSS.n1068 VSS.n1067 0.00334
R9163 VSS.n1069 VSS.n1068 0.00334
R9164 VSS.n1071 VSS.n1069 0.00334
R9165 VSS.n1072 VSS.n1071 0.00334
R9166 VSS.n1073 VSS.n1072 0.00334
R9167 VSS.n1077 VSS.n1076 0.00334
R9168 VSS.n584 VSS.n370 0.00334
R9169 VSS.n585 VSS.n584 0.00334
R9170 VSS.n586 VSS.n585 0.00334
R9171 VSS.n587 VSS.n586 0.00334
R9172 VSS.n588 VSS.n587 0.00334
R9173 VSS.n591 VSS.n588 0.00334
R9174 VSS.n592 VSS.n591 0.00334
R9175 VSS.n593 VSS.n592 0.00334
R9176 VSS.n594 VSS.n593 0.00334
R9177 VSS.n597 VSS.n594 0.00334
R9178 VSS.n598 VSS.n597 0.00334
R9179 VSS.n599 VSS.n598 0.00334
R9180 VSS.n600 VSS.n599 0.00334
R9181 VSS.n603 VSS.n600 0.00334
R9182 VSS.n604 VSS.n603 0.00334
R9183 VSS.n605 VSS.n604 0.00334
R9184 VSS.n606 VSS.n605 0.00334
R9185 VSS.n606 VSS.n327 0.00334
R9186 VSS.n755 VSS.n327 0.00334
R9187 VSS.n756 VSS.n755 0.00334
R9188 VSS.n757 VSS.n756 0.00334
R9189 VSS.n757 VSS.n323 0.00334
R9190 VSS.n763 VSS.n323 0.00334
R9191 VSS.n765 VSS.n317 0.00334
R9192 VSS.n771 VSS.n317 0.00334
R9193 VSS.n772 VSS.n771 0.00334
R9194 VSS.n773 VSS.n772 0.00334
R9195 VSS.n773 VSS.n313 0.00334
R9196 VSS.n779 VSS.n313 0.00334
R9197 VSS.n780 VSS.n779 0.00334
R9198 VSS.n781 VSS.n780 0.00334
R9199 VSS.n781 VSS.n309 0.00334
R9200 VSS.n787 VSS.n309 0.00334
R9201 VSS.n788 VSS.n787 0.00334
R9202 VSS.n789 VSS.n788 0.00334
R9203 VSS.n790 VSS.n789 0.00334
R9204 VSS.n791 VSS.n790 0.00334
R9205 VSS.n794 VSS.n791 0.00334
R9206 VSS.n795 VSS.n794 0.00334
R9207 VSS.n796 VSS.n795 0.00334
R9208 VSS.n797 VSS.n796 0.00334
R9209 VSS.n800 VSS.n797 0.00334
R9210 VSS.n801 VSS.n800 0.00334
R9211 VSS.n802 VSS.n801 0.00334
R9212 VSS.n803 VSS.n802 0.00334
R9213 VSS.n804 VSS.n803 0.00334
R9214 VSS.n138 VSS.n137 0.00334
R9215 VSS.n139 VSS.n138 0.00334
R9216 VSS.n142 VSS.n139 0.00334
R9217 VSS.n143 VSS.n142 0.00334
R9218 VSS.n144 VSS.n143 0.00334
R9219 VSS.n147 VSS.n144 0.00334
R9220 VSS.n148 VSS.n147 0.00334
R9221 VSS.n149 VSS.n148 0.00334
R9222 VSS.n150 VSS.n149 0.00334
R9223 VSS.n153 VSS.n150 0.00334
R9224 VSS.n154 VSS.n153 0.00334
R9225 VSS.n155 VSS.n154 0.00334
R9226 VSS.n156 VSS.n155 0.00334
R9227 VSS.n159 VSS.n156 0.00334
R9228 VSS.n160 VSS.n159 0.00334
R9229 VSS.n161 VSS.n160 0.00334
R9230 VSS.n162 VSS.n161 0.00334
R9231 VSS.n165 VSS.n162 0.00334
R9232 VSS.n166 VSS.n165 0.00334
R9233 VSS.n167 VSS.n166 0.00334
R9234 VSS.n169 VSS.n167 0.00334
R9235 VSS.n169 VSS.n168 0.00334
R9236 VSS.n168 VSS.n97 0.00334
R9237 VSS.n1112 VSS.n91 0.00334
R9238 VSS.n1113 VSS.n1112 0.00334
R9239 VSS.n1114 VSS.n1113 0.00334
R9240 VSS.n1114 VSS.n87 0.00334
R9241 VSS.n1120 VSS.n87 0.00334
R9242 VSS.n1121 VSS.n1120 0.00334
R9243 VSS.n1122 VSS.n1121 0.00334
R9244 VSS.n1122 VSS.n83 0.00334
R9245 VSS.n1128 VSS.n83 0.00334
R9246 VSS.n1129 VSS.n1128 0.00334
R9247 VSS.n1130 VSS.n1129 0.00334
R9248 VSS.n1136 VSS.n79 0.00334
R9249 VSS.n389 VSS.n388 0.00334
R9250 VSS.n392 VSS.n389 0.00334
R9251 VSS.n393 VSS.n392 0.00334
R9252 VSS.n394 VSS.n393 0.00334
R9253 VSS.n395 VSS.n394 0.00334
R9254 VSS.n398 VSS.n395 0.00334
R9255 VSS.n399 VSS.n398 0.00334
R9256 VSS.n400 VSS.n399 0.00334
R9257 VSS.n401 VSS.n400 0.00334
R9258 VSS.n404 VSS.n401 0.00334
R9259 VSS.n405 VSS.n404 0.00334
R9260 VSS.n406 VSS.n405 0.00334
R9261 VSS.n407 VSS.n406 0.00334
R9262 VSS.n410 VSS.n407 0.00334
R9263 VSS.n411 VSS.n410 0.00334
R9264 VSS.n412 VSS.n411 0.00334
R9265 VSS.n413 VSS.n412 0.00334
R9266 VSS.n415 VSS.n413 0.00334
R9267 VSS.n416 VSS.n415 0.00334
R9268 VSS.n417 VSS.n416 0.00334
R9269 VSS.n420 VSS.n417 0.00334
R9270 VSS.n421 VSS.n420 0.00334
R9271 VSS.n422 VSS.n421 0.00334
R9272 VSS.n427 VSS.n423 0.00334
R9273 VSS.n428 VSS.n427 0.00334
R9274 VSS.n429 VSS.n428 0.00334
R9275 VSS.n430 VSS.n429 0.00334
R9276 VSS.n433 VSS.n430 0.00334
R9277 VSS.n434 VSS.n433 0.00334
R9278 VSS.n435 VSS.n434 0.00334
R9279 VSS.n436 VSS.n435 0.00334
R9280 VSS.n439 VSS.n436 0.00334
R9281 VSS.n440 VSS.n439 0.00334
R9282 VSS.n441 VSS.n440 0.00334
R9283 VSS.n442 VSS.n441 0.00334
R9284 VSS.n445 VSS.n442 0.00334
R9285 VSS.n446 VSS.n445 0.00334
R9286 VSS.n447 VSS.n446 0.00334
R9287 VSS.n448 VSS.n447 0.00334
R9288 VSS.n451 VSS.n448 0.00334
R9289 VSS.n452 VSS.n451 0.00334
R9290 VSS.n453 VSS.n452 0.00334
R9291 VSS.n454 VSS.n453 0.00334
R9292 VSS.n455 VSS.n454 0.00334
R9293 VSS.n455 VSS.n129 0.00334
R9294 VSS.n956 VSS.n129 0.00334
R9295 VSS.n959 VSS.n958 0.00334
R9296 VSS.n959 VSS.n124 0.00334
R9297 VSS.n966 VSS.n124 0.00334
R9298 VSS.n967 VSS.n966 0.00334
R9299 VSS.n968 VSS.n967 0.00334
R9300 VSS.n968 VSS.n120 0.00334
R9301 VSS.n974 VSS.n120 0.00334
R9302 VSS.n975 VSS.n974 0.00334
R9303 VSS.n976 VSS.n975 0.00334
R9304 VSS.n976 VSS.n116 0.00334
R9305 VSS.n982 VSS.n116 0.00334
R9306 VSS.n983 VSS.n982 0.00334
R9307 VSS.n984 VSS.n983 0.00334
R9308 VSS.n984 VSS.n112 0.00334
R9309 VSS.n990 VSS.n112 0.00334
R9310 VSS.n991 VSS.n990 0.00334
R9311 VSS.n992 VSS.n991 0.00334
R9312 VSS.n992 VSS.n108 0.00334
R9313 VSS.n998 VSS.n108 0.00334
R9314 VSS.n999 VSS.n998 0.00334
R9315 VSS.n1000 VSS.n999 0.00334
R9316 VSS.n1000 VSS.n101 0.00334
R9317 VSS.n1009 VSS.n101 0.00334
R9318 VSS.n1053 VSS.n1010 0.00334
R9319 VSS.n1013 VSS.n1010 0.00334
R9320 VSS.n1014 VSS.n1013 0.00334
R9321 VSS.n1015 VSS.n1014 0.00334
R9322 VSS.n1018 VSS.n1015 0.00334
R9323 VSS.n1019 VSS.n1018 0.00334
R9324 VSS.n1020 VSS.n1019 0.00334
R9325 VSS.n1021 VSS.n1020 0.00334
R9326 VSS.n1023 VSS.n1021 0.00334
R9327 VSS.n1024 VSS.n1023 0.00334
R9328 VSS.n1025 VSS.n1024 0.00334
R9329 VSS.n1028 VSS.n1027 0.00334
R9330 VSS.n1958 VSS.n1700 0.00332857
R9331 VSS.n1957 VSS.n1701 0.00332857
R9332 VSS.n1707 VSS.n1706 0.00332857
R9333 VSS.n1950 VSS.n1949 0.00332857
R9334 VSS.n1714 VSS.n1708 0.00332857
R9335 VSS.n1943 VSS.n1715 0.00332857
R9336 VSS.n1942 VSS.n1935 0.00332857
R9337 VSS.n4751 VSS.n4750 0.00332857
R9338 VSS.n576 VSS.n376 0.00332
R9339 VSS.n378 VSS.n371 0.00332
R9340 VSS.n383 VSS.n379 0.00332
R9341 VSS.n382 VSS.n372 0.00332
R9342 VSS.n580 VSS.n579 0.00332
R9343 VSS.n578 VSS.n577 0.00332
R9344 VSS.n1150 VSS.n29 0.00330488
R9345 VSS.n1165 VSS.n24 0.00330488
R9346 VSS.n826 VSS.n825 0.00329
R9347 VSS.n823 VSS.n306 0.00329
R9348 VSS.n438 VSS.n305 0.00329
R9349 VSS.n2165 DVSS 0.00326
R9350 VSS.n1027 DVSS 0.00326
R9351 VSS.n4527 VSS.n4526 0.0032
R9352 VSS.n3517 VSS.n3516 0.0032
R9353 VSS.n915 VSS.n170 0.00319327
R9354 VSS.n2615 VSS.n2605 0.00319022
R9355 VSS.n4333 VSS.n2612 0.00319022
R9356 VSS.n4304 VSS 0.00314706
R9357 VSS VSS.n2629 0.00314706
R9358 VSS.n571 VSS.n523 0.00314706
R9359 VSS.n3553 VSS.n3552 0.00313571
R9360 VSS.n3575 VSS.n2719 0.00313571
R9361 VSS.n671 VSS.n670 0.00311
R9362 VSS.n630 VSS.n367 0.00311
R9363 VSS.n573 VSS.n572 0.00311
R9364 VSS.n2169 VSS.n2168 0.00309529
R9365 VSS.n1030 VSS.n1029 0.00309529
R9366 VSS.n1137 VSS.n78 0.00309529
R9367 VSS.n1081 VSS.n1080 0.00309529
R9368 VSS.n3715 VSS.n3714 0.00307143
R9369 VSS.n2656 VSS.n2654 0.00307143
R9370 VSS.n3718 VSS.n2661 0.00307143
R9371 VSS.n1836 VSS.n19 0.00300714
R9372 VSS.n1587 VSS.n1298 0.00300714
R9373 VSS.n3561 VSS.n3534 0.00300714
R9374 VSS.n3189 VSS.n3188 0.003
R9375 VSS.n4889 VSS.n2396 0.003
R9376 VSS.n2817 VSS.n2800 0.003
R9377 VSS.n3210 VSS.n2399 0.003
R9378 VSS.n3831 VSS.n3823 0.00297706
R9379 VSS.n2937 VSS.n2926 0.00296479
R9380 VSS.n2946 VSS.n2945 0.00296479
R9381 VSS.n2928 VSS.n2922 0.00296479
R9382 VSS.n2955 VSS.n2917 0.00296479
R9383 VSS.n2971 VSS.n2970 0.00296479
R9384 VSS.n2979 VSS.n2912 0.00296479
R9385 VSS.n2978 VSS.n2906 0.00296479
R9386 VSS.n2990 VSS.n2989 0.00296479
R9387 VSS.n2908 VSS.n2902 0.00296479
R9388 VSS.n2998 VSS.n2897 0.00296479
R9389 VSS.n3018 VSS.n3017 0.00296479
R9390 VSS.n3026 VSS.n2892 0.00296479
R9391 VSS.n3025 VSS.n2886 0.00296479
R9392 VSS.n3041 VSS.n3040 0.00296479
R9393 VSS.n3037 VSS.n2888 0.00296479
R9394 VSS.n3036 VSS.n2880 0.00296479
R9395 VSS.n3052 VSS.n2875 0.00296479
R9396 VSS.n3079 VSS.n3078 0.00296479
R9397 VSS.n3087 VSS.n2870 0.00296479
R9398 VSS.n3086 VSS.n2863 0.00296479
R9399 VSS.n3094 VSS.n3093 0.00296479
R9400 VSS.n2866 VSS.n2865 0.00296479
R9401 VSS.n3106 VSS.n2857 0.00296479
R9402 VSS.n3105 VSS.n2851 0.00296479
R9403 VSS.n3117 VSS.n3116 0.00296479
R9404 VSS.n2853 VSS.n2847 0.00296479
R9405 VSS.n3125 VSS.n2842 0.00296479
R9406 VSS.n3140 VSS.n3139 0.00296479
R9407 VSS.n3150 VSS.n2837 0.00296479
R9408 VSS.n3149 VSS.n2830 0.00296479
R9409 VSS.n3162 VSS.n3161 0.00296479
R9410 VSS.n2833 VSS.n2826 0.00296479
R9411 VSS.n3169 VSS.n2821 0.00296479
R9412 VSS.n3180 VSS.n3179 0.00296479
R9413 VSS.n3191 VSS.n2816 0.00296479
R9414 VSS.n3190 VSS.n2802 0.00296479
R9415 VSS.n3238 VSS.n2803 0.00296479
R9416 VSS.n3201 VSS.n2809 0.00296479
R9417 VSS.n3231 VSS.n3230 0.00296479
R9418 VSS.n3227 VSS.n2811 0.00296479
R9419 VSS.n3226 VSS.n3218 0.00296479
R9420 VSS.n4877 VSS.n2404 0.00296479
R9421 VSS.n4876 VSS.n2397 0.00296479
R9422 VSS.n4888 VSS.n4887 0.00296479
R9423 VSS.n2400 VSS.n2393 0.00296479
R9424 VSS.n4895 VSS.n2388 0.00296479
R9425 VSS.n4914 VSS.n4913 0.00296479
R9426 VSS.n4924 VSS.n2383 0.00296479
R9427 VSS.n4923 VSS.n2377 0.00296479
R9428 VSS.n4941 VSS.n4940 0.00296479
R9429 VSS.n2379 VSS.n2371 0.00296479
R9430 VSS.n4950 VSS.n2373 0.00296479
R9431 VSS.n2372 VSS.n2367 0.00296479
R9432 VSS.n4957 VSS.n2359 0.00296479
R9433 VSS.n4968 VSS.n2360 0.00296479
R9434 VSS.n2363 VSS.n2362 0.00296479
R9435 VSS.n4986 VSS.n2351 0.00296479
R9436 VSS.n4985 VSS.n2344 0.00296479
R9437 VSS.n4997 VSS.n4996 0.00296479
R9438 VSS.n2347 VSS.n2340 0.00296479
R9439 VSS.n5004 VSS.n2335 0.00296479
R9440 VSS.n5019 VSS.n5018 0.00296479
R9441 VSS.n5029 VSS.n2330 0.00296479
R9442 VSS.n5028 VSS.n2323 0.00296479
R9443 VSS.n5040 VSS.n5039 0.00296479
R9444 VSS.n2326 VSS.n2319 0.00296479
R9445 VSS.n5047 VSS.n2314 0.00296479
R9446 VSS.n5065 VSS.n5064 0.00296479
R9447 VSS.n5075 VSS.n2309 0.00296479
R9448 VSS.n5074 VSS.n2303 0.00296479
R9449 VSS.n5090 VSS.n5089 0.00296479
R9450 VSS.n2305 VSS.n2297 0.00296479
R9451 VSS.n5098 VSS.n2299 0.00296479
R9452 VSS.n2298 VSS.n2293 0.00296479
R9453 VSS.n5105 VSS.n2287 0.00296479
R9454 VSS.n5116 VSS.n2288 0.00296479
R9455 VSS.n5127 VSS.n2283 0.00296479
R9456 VSS.n5126 VSS.n2277 0.00296479
R9457 VSS.n5170 VSS.n5169 0.00296479
R9458 VSS.n631 VSS.n366 0.00294344
R9459 DVSS VSS.n3021 0.00293842
R9460 VSS.n3014 DVSS 0.00293842
R9461 VSS.n4080 VSS.n4079 0.00293243
R9462 VSS.n265 VSS.n264 0.0029
R9463 VSS.n1107 VSS.n95 0.0029
R9464 VSS.n1007 VSS.n1006 0.0029
R9465 VSS.n5445 DVSS 0.00286842
R9466 DVSS VSS.n5351 0.00286842
R9467 VSS.n5412 DVSS 0.00286842
R9468 VSS.n2107 DVSS 0.00286842
R9469 VSS VSS.n2515 0.00286842
R9470 VSS.n1057 VSS.n1056 0.00286
R9471 VSS.n1055 VSS.n91 0.00286
R9472 VSS.n1054 VSS.n1053 0.00286
R9473 VSS.n1076 DVSS 0.00282
R9474 VSS.n2087 DVSS 0.00279616
R9475 VSS.n2174 DVSS 0.00279616
R9476 VSS.n5410 DVSS 0.00279616
R9477 VSS.n2526 DVSS 0.00279616
R9478 DVSS VSS.n2160 0.00278
R9479 VSS.n3186 VSS.n2806 0.00271675
R9480 VSS.n3242 VSS.n3241 0.00271675
R9481 VSS.n854 VSS.n853 0.0027
R9482 VSS.n137 VSS.n128 0.0027
R9483 VSS.n958 VSS.n957 0.0027
R9484 VSS.n5381 VSS.n2134 0.00269
R9485 VSS.n1990 VSS.n1989 0.00262143
R9486 VSS.n1986 VSS.n1675 0.00262143
R9487 VSS.n1985 VSS.n1678 0.00262143
R9488 VSS.n1683 VSS.n1682 0.00262143
R9489 VSS.n1979 VSS.n1978 0.00262143
R9490 VSS.n1688 VSS.n1684 0.00262143
R9491 VSS.n1973 VSS.n1689 0.00262143
R9492 VSS.n1858 VSS.n1792 0.00262143
R9493 VSS.n1857 VSS.n1798 0.00262143
R9494 VSS.n1854 VSS.n1853 0.00262143
R9495 VSS.n1157 VSS.n30 0.00257317
R9496 VSS.n1158 VSS.n26 0.00257317
R9497 VSS.n4531 VSS.n2544 0.00257
R9498 VSS.n5378 VSS.n2134 0.00257
R9499 VSS.n3943 VSS.n3908 0.00256422
R9500 VSS.n3750 VSS.n3749 0.00256422
R9501 VSS.n2021 VSS.n1648 0.00255714
R9502 VSS.n2018 VSS.n2017 0.00255714
R9503 VSS.n1657 VSS.n1651 0.00255714
R9504 VSS.n2011 VSS.n1658 0.00255714
R9505 VSS.n2010 VSS.n1659 0.00255714
R9506 VSS.n1664 VSS.n1663 0.00255714
R9507 VSS.n2005 VSS.n2004 0.00255714
R9508 VSS.n714 VSS.n322 0.00254
R9509 VSS.n765 VSS.n764 0.00254
R9510 VSS.n423 VSS.n321 0.00254
R9511 VSS.n216 VSS.n170 0.00251995
R9512 VSS.n3237 VSS.n2804 0.0025
R9513 VSS.n4875 VSS.n4874 0.0025
R9514 VSS.n3240 VSS.n3239 0.0025
R9515 VSS.n3211 VSS.n2405 0.0025
R9516 VSS.n4135 VSS.n3769 0.00249286
R9517 VSS.n3922 VSS.n3771 0.00249286
R9518 DVSS VSS.n5150 0.00247183
R9519 VSS.n3879 VSS.n3875 0.00242857
R9520 VSS.n3876 VSS.n3761 0.00242857
R9521 VSS.n385 VSS.n384 0.00238
R9522 VSS.n386 VSS.n370 0.00238
R9523 VSS.n388 VSS.n387 0.00238
R9524 VSS.n3683 VSS.n3682 0.00236429
R9525 VSS.n266 VSS.n265 0.00236
R9526 VSS.n917 VSS.n95 0.00236
R9527 VSS.n1006 VSS.n103 0.00236
R9528 VSS.n535 VSS.n366 0.00233258
R9529 VSS VSS.n3374 0.0023
R9530 VSS.n3995 DVSS 0.0023
R9531 VSS.n4380 DVSS 0.0023
R9532 DVSS VSS.n1839 0.0023
R9533 VSS.n1838 DVSS 0.0023
R9534 VSS.n1397 DVSS 0.0023
R9535 VSS.n5189 DVSS 0.0023
R9536 VSS.n3373 VSS 0.0023
R9537 VSS VSS.n5723 0.0023
R9538 VSS.n5722 VSS 0.0023
R9539 VSS.n4873 VSS.n4872 0.0022734
R9540 VSS.n4855 VSS.n2417 0.00223571
R9541 VSS.n3372 VSS.n2422 0.00223571
R9542 VSS.n3373 VSS.n2416 0.00223571
R9543 VSS.n4825 VSS.n2432 0.00223571
R9544 VSS.n4824 VSS.n0 0.00223571
R9545 VSS.n5723 VSS.n1 0.00223571
R9546 VSS.n670 VSS.n348 0.00215
R9547 VSS.n630 VSS.n629 0.00215
R9548 VSS.n572 VSS.n522 0.00215
R9549 VSS.n3148 VSS.n3147 0.002
R9550 VSS.n4943 VSS.n4942 0.002
R9551 VSS.n3133 VSS.n2838 0.002
R9552 VSS.n4903 VSS.n2378 0.002
R9553 VSS.n2250 VSS.n2244 0.00197857
R9554 VSS.n825 VSS.n300 0.00197
R9555 VSS.n823 VSS.n822 0.00197
R9556 VSS.n470 VSS.n305 0.00197
R9557 VSS.n1130 DVSS 0.00196
R9558 DVSS VSS.n32 0.00191429
R9559 DVSS VSS.n79 0.00188
R9560 VSS.n3545 VSS.n2723 0.00185
R9561 VSS.n3577 VSS.n2715 0.00185
R9562 VSS.n5704 VSS.n21 0.00184146
R9563 VSS.n1166 VSS.n27 0.00184146
R9564 VSS.n5252 DVSS 0.00179393
R9565 VSS.n1131 DVSS 0.00173
R9566 DVSS VSS.n1132 0.00173
R9567 VSS.n491 VSS.n490 0.0017
R9568 VSS.n762 VSS.n320 0.0017
R9569 VSS.n713 VSS.n711 0.0017
R9570 VSS.n744 VSS.n743 0.0017
R9571 VSS.n761 VSS.n319 0.0017
R9572 VSS.n425 VSS.n419 0.0017
R9573 VSS.n901 VSS.n900 0.00167
R9574 VSS.n918 VSS.n916 0.00167
R9575 VSS.n1003 VSS.n1002 0.00167
R9576 VSS.n1834 VSS.n20 0.00165714
R9577 VSS.n1830 VSS.n22 0.00165714
R9578 VSS.n4088 VSS.n3964 0.00165714
R9579 VSS.n4090 VSS.n4057 0.00165714
R9580 VSS.n4285 VSS.n4276 0.00165714
R9581 VSS.n4283 VSS.n4282 0.00165714
R9582 VSS.n4279 VSS.n4278 0.00165714
R9583 VSS.n4677 VSS.n2506 0.00165714
R9584 VSS.n4676 VSS.n2507 0.00165714
R9585 VSS.n4683 VSS.n2502 0.00165714
R9586 VSS.n4684 VSS.n2500 0.00165714
R9587 VSS.n4687 VSS.n4686 0.00165714
R9588 VSS.n2556 VSS.n2551 0.00159286
R9589 VSS.n4515 VSS.n4514 0.00159286
R9590 VSS.n4512 VSS.n2562 0.00159286
R9591 VSS.n1724 VSS.n1720 0.00159286
R9592 VSS.n1920 VSS.n1919 0.00159286
R9593 VSS.n1748 VSS.n1725 0.00159286
R9594 VSS.n1912 VSS.n1749 0.00159286
R9595 VSS.n1911 VSS.n1750 0.00159286
R9596 VSS.n1757 VSS.n1756 0.00159286
R9597 VSS.n1905 VSS.n1904 0.00159286
R9598 VSS.n2692 VSS.n2688 0.00159286
R9599 VSS.n3865 VSS.n2561 0.00157001
R9600 VSS.n3826 VSS.n2644 0.00152857
R9601 VSS.n4175 VSS.n2648 0.00152857
R9602 VSS.n3100 VSS.n2859 0.0015
R9603 VSS.n4962 VSS.n2353 0.0015
R9604 VSS.n3066 VSS.n3058 0.0015
R9605 VSS.n4975 VSS.n4974 0.0015
R9606 VSS.n955 VSS.n131 0.00146
R9607 VSS.n805 VSS.n136 0.00146
R9608 VSS.n851 VSS.n291 0.00146
R9609 VSS.n850 VSS.n133 0.00146
R9610 VSS.n952 VSS.n134 0.00146
R9611 VSS.n954 VSS.n953 0.00146
R9612 VSS.n4574 VSS.n4568 0.00146
R9613 DVSS VSS.n5355 0.00134
R9614 DVSS VSS.n1035 0.00134
R9615 VSS.n1034 DVSS 0.00134
R9616 VSS.n5354 DVSS 0.00134
R9617 VSS.n4439 VSS.n2609 0.00133571
R9618 VSS.n4348 VSS.n2614 0.00133571
R9619 VSS.n4437 VSS.n4436 0.00133571
R9620 VSS.n3599 VSS.n3598 0.00133571
R9621 VSS.n859 VSS.n283 0.00131
R9622 VSS.n945 VSS.n141 0.00131
R9623 VSS.n963 VSS.n122 0.00131
R9624 VSS.n5390 VSS.n5389 0.00131
R9625 VSS.n5354 VSS.n5353 0.00131
R9626 VSS.n710 VSS.n322 0.0013
R9627 VSS.n764 VSS.n763 0.0013
R9628 VSS.n422 VSS.n321 0.0013
R9629 VSS.n1008 VSS.n98 0.00122
R9630 VSS.n1106 VSS.n1105 0.00122
R9631 VSS.n1104 VSS.n99 0.00122
R9632 VSS.n264 VSS.n94 0.00122
R9633 VSS.n1108 VSS.n1107 0.00122
R9634 VSS.n1007 VSS.n93 0.00122
R9635 VSS.n5703 DVSS 0.00120714
R9636 VSS.n3650 VSS.n3649 0.00120714
R9637 VSS.n3665 VSS.n3664 0.00120714
R9638 VSS.n4219 VSS.n4218 0.00120714
R9639 VSS.n4301 VSS.n4300 0.00120714
R9640 VSS.n4545 VSS.n4544 0.00119
R9641 VSS.n4664 VSS.n2531 0.00119
R9642 VSS.n853 VSS.n852 0.00114
R9643 VSS.n804 VSS.n128 0.00114
R9644 VSS.n957 VSS.n956 0.00114
R9645 VSS.n5401 VSS.n5400 0.00107
R9646 VSS.n2172 VSS.n2171 0.00107
R9647 VSS.n2161 DVSS 0.00106
R9648 VSS.n1139 VSS.n57 0.00104
R9649 VSS.n1138 VSS.n77 0.00104
R9650 VSS.n1142 VSS.n36 0.00104
R9651 VSS.n37 VSS.n34 0.00104
R9652 DVSS VSS.n1073 0.00102
R9653 VSS.n750 VSS.n331 0.00101
R9654 VSS.n753 VSS.n752 0.00101
R9655 VSS.n498 VSS.n330 0.00101
R9656 VSS.n2948 VSS.n2947 0.001
R9657 VSS.n3047 VSS.n2881 0.001
R9658 VSS.n5027 VSS.n5026 0.001
R9659 VSS.n5110 VSS.n2276 0.001
R9660 VSS.n2933 VSS.n2927 0.001
R9661 VSS.n3005 VSS.n2879 0.001
R9662 VSS.n5011 VSS.n2331 0.001
R9663 VSS.n5125 VSS.n5124 0.001
R9664 VSS.n1056 VSS.n100 0.00098
R9665 VSS.n1055 VSS.n97 0.00098
R9666 VSS.n1054 VSS.n1009 0.00098
R9667 VSS.n3539 VSS.n3538 0.00095
R9668 VSS.n4918 VSS.n4917 0.00094335
R9669 VSS.n4910 VSS.n4909 0.00094335
R9670 VSS.n381 VSS.n352 0.00092
R9671 VSS.n582 VSS.n581 0.00092
R9672 VSS.n574 VSS.n375 0.00092
R9673 VSS.n1396 VSS.n32 0.000885714
R9674 VSS.n3856 VSS.n2564 0.000856671
R9675 VSS.n3847 VSS.n2558 0.000856671
R9676 DVSS VSS.n2930 0.000721675
R9677 VSS.n2935 DVSS 0.000721675
R9678 DVSS VSS.n5148 0.000687793
R9679 DVSS VSS.n1086 0.00068
R9680 VSS.n1085 DVSS 0.00068
R9681 VSS.n5721 VSS 0.000671429
R9682 VSS VSS.n3358 0.000671429
R9683 VSS.n3996 DVSS 0.000671429
R9684 DVSS VSS.n4379 0.000671429
R9685 DVSS VSS.n1827 0.000671429
R9686 VSS.n1398 DVSS 0.000671429
R9687 VSS.n5190 DVSS 0.000671429
R9688 VSS.n3827 VSS.n3826 0.000628571
R9689 VSS.n4175 VSS.n4174 0.000628571
R9690 VSS.n3797 VSS.n2649 0.000628571
R9691 VSS.n3804 VSS.n3798 0.000628571
R9692 VSS.n3803 VSS.n3796 0.000628571
R9693 VSS.n3806 VSS.n3794 0.000628571
R9694 VSS.n3807 VSS.n3731 0.000628571
R9695 VSS.n3790 VSS.n3733 0.000628571
R9696 VSS.n3813 VSS.n3730 0.000628571
R9697 VSS.n4162 VSS.n3734 0.000628571
R9698 VSS.n4160 VSS.n3735 0.000628571
R9699 VSS.n3742 VSS.n3741 0.000628571
R9700 VSS.n4154 VSS.n4153 0.000628571
R9701 VSS.n3872 VSS.n3743 0.000628571
R9702 VSS.n3875 VSS.n3759 0.000628571
R9703 VSS.n4144 VSS.n3761 0.000628571
R9704 VSS.n4136 VSS.n4135 0.000628571
R9705 VSS.n3771 VSS.n3770 0.000628571
R9706 VSS.n3924 VSS.n3923 0.000628571
R9707 VSS.n3932 VSS.n3931 0.000628571
R9708 VSS.n3940 VSS.n3911 0.000628571
R9709 VSS.n3939 VSS.n3912 0.000628571
R9710 VSS.n3914 VSS.n3888 0.000628571
R9711 VSS.n3892 VSS.n3891 0.000628571
R9712 VSS.n4113 VSS.n3893 0.000628571
R9713 VSS.n3900 VSS.n3899 0.000628571
R9714 VSS.n4107 VSS.n4106 0.000628571
R9715 VSS.n3956 VSS.n3901 0.000628571
R9716 VSS.n4098 VSS.n3957 0.000628571
R9717 VSS.n4097 VSS.n3958 0.000628571
R9718 VSS.n4088 VSS.n4087 0.000628571
R9719 VSS.n4091 VSS.n4090 0.000628571
R9720 DVSS VSS.n2161 0.00058
R9721 DVSS VSS.n1025 0.00058
R9722 VSS.n5163 VSS.n5135 0.000570422
R9723 VSS.n5694 VSS.n1170 0.000566519
R9724 VSS.n5183 VSS.n2267 0.000564286
R9725 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t4 37.5434
R9726 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t5 37.5434
R9727 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t2 25.3941
R9728 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t3 25.3941
R9729 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.n0 8.44221
R9730 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.n1 4.93097
R9731 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t1 2.6373
R9732 CS.n0 CS.t1 35.9269
R9733 CS.n0 CS.t2 30.9212
R9734 CS.n2 CS 18.5934
R9735 CS CS.n0 4.0005
R9736 CS.n2 CS.n1 2.4573
R9737 CS.n1 CS.t0 1.30145
R9738 CS CS.n2 0.840105
R9739 CS.n1 CS 0.01495
R9740 VDD.n442 VDD.n295 512.403
R9741 VDD VDD.t8 378.373
R9742 VDD.n594 VDD.t56 352.072
R9743 VDD.t43 VDD.t28 321.485
R9744 VDD.t8 VDD.t33 321.485
R9745 VDD.t32 VDD.t56 321.485
R9746 VDD.n650 VDD.t15 314.901
R9747 VDD.n597 VDD.t61 280.788
R9748 VDD.t10 VDD.n583 280.702
R9749 VDD.t4 VDD.n578 278.981
R9750 VDD.n578 VDD.t2 278.981
R9751 VDD.t45 VDD.n374 264.098
R9752 VDD.t0 VDD.n364 264.098
R9753 VDD.t13 VDD.n357 263.524
R9754 VDD.n357 VDD.t63 263.524
R9755 VDD.n662 VDD.t41 248.441
R9756 VDD.n218 VDD.n207 227.274
R9757 VDD.n224 VDD.n201 227.274
R9758 VDD.n872 VDD.t6 224.88
R9759 VDD.n233 VDD.t50 223.204
R9760 VDD.n233 VDD.t58 223.204
R9761 VDD.n876 VDD.t24 202.791
R9762 VDD.n195 VDD.t22 202.791
R9763 VDD.t52 VDD.n926 202.791
R9764 VDD.t20 VDD.n122 201.413
R9765 VDD.t15 VDD.t34 188.564
R9766 VDD.t34 VDD.t30 188.564
R9767 VDD.t30 VDD.t17 188.564
R9768 VDD.t17 VDD.t26 188.564
R9769 VDD.t37 VDD.t43 188.564
R9770 VDD.t39 VDD.t37 188.564
R9771 VDD.t41 VDD.t39 188.564
R9772 VDD.n129 VDD.t47 187.478
R9773 VDD.n122 VDD.t54 183.157
R9774 VDD.n580 VDD.t32 173.88
R9775 VDD.t33 VDD.n580 147.605
R9776 VDD.n661 VDD.t26 139.105
R9777 VDD.n218 VDD.t60 113.636
R9778 VDD.t60 VDD.n201 113.636
R9779 VDD.n77 VDD.n54 105.84
R9780 VDD.t19 VDD.n54 105.84
R9781 VDD.t19 VDD.n45 105.84
R9782 VDD.n96 VDD.n45 105.84
R9783 VDD.n584 VDD.t10 94.2818
R9784 VDD.n584 VDD.t4 94.2818
R9785 VDD.n596 VDD.t2 94.2818
R9786 VDD.t61 VDD.n596 94.2818
R9787 VDD.t24 VDD.n875 82.4504
R9788 VDD.n232 VDD.t22 82.4504
R9789 VDD.n927 VDD.t52 82.4504
R9790 VDD.n386 VDD.n312 75.7185
R9791 VDD.n386 VDD.t36 75.7185
R9792 VDD.n400 VDD.t36 75.7185
R9793 VDD.n400 VDD.n295 75.7185
R9794 VDD.n442 VDD.n300 75.7185
R9795 VDD.t12 VDD.n300 75.7185
R9796 VDD.t12 VDD.n427 75.7185
R9797 VDD.n427 VDD.n289 75.7185
R9798 VDD.n128 VDD.t54 73.6165
R9799 VDD.n123 VDD.n121 70.1484
R9800 VDD.t47 VDD.n128 70.083
R9801 VDD.n875 VDD.t6 61.249
R9802 VDD.t50 VDD.n232 61.249
R9803 VDD.n927 VDD.t58 61.249
R9804 VDD.n376 VDD.n374 53.6905
R9805 VDD.n364 VDD.n361 53.6905
R9806 VDD.t28 VDD.n661 49.4595
R9807 VDD.n197 VDD.t65 46.7726
R9808 VDD.n375 VDD.n373 45.0389
R9809 VDD.n349 VDD.n343 45.0389
R9810 VDD.n359 VDD.n358 45.0389
R9811 VDD.n366 VDD.n365 45.0389
R9812 VDD.n197 VDD.t49 41.2455
R9813 VDD.n356 VDD.n355 29.7505
R9814 VDD.n355 VDD.n348 23.9405
R9815 VDD.n355 VDD.n354 23.9405
R9816 VDD.n219 VDD.n206 10.5005
R9817 VDD.n219 VDD.n203 10.5005
R9818 VDD.n223 VDD.n203 10.5005
R9819 VDD.n213 VDD.n212 10.5005
R9820 VDD.n217 VDD.n208 10.5005
R9821 VDD.n217 VDD.n200 10.5005
R9822 VDD.n225 VDD.n200 10.5005
R9823 VDD.n330 VDD.n329 10.1505
R9824 VDD.n333 VDD.n330 10.1505
R9825 VDD.n320 VDD.n314 10.1505
R9826 VDD.n317 VDD.n314 10.1505
R9827 VDD.n452 VDD.n451 10.1505
R9828 VDD.n441 VDD.n435 10.1505
R9829 VDD.n435 VDD.n433 10.1505
R9830 VDD.n433 VDD.n288 10.1505
R9831 VDD.n454 VDD.n288 10.1505
R9832 VDD.n432 VDD.n429 10.1505
R9833 VDD.n430 VDD.n290 10.1505
R9834 VDD.n438 VDD.n437 10.1505
R9835 VDD.n385 VDD.n325 10.1505
R9836 VDD.n385 VDD.n304 10.1505
R9837 VDD.n401 VDD.n304 10.1505
R9838 VDD.n402 VDD.n401 10.1505
R9839 VDD.n328 VDD.n313 10.1505
R9840 VDD.n328 VDD.n305 10.1505
R9841 VDD.n338 VDD.n337 10.1505
R9842 VDD.n444 VDD.n294 10.1505
R9843 VDD.n414 VDD.n299 10.1505
R9844 VDD.n414 VDD.n407 10.1505
R9845 VDD.n408 VDD.n407 10.1505
R9846 VDD.n417 VDD.n408 10.1505
R9847 VDD.n422 VDD.n421 10.1505
R9848 VDD.n421 VDD.n420 10.1505
R9849 VDD.n406 VDD.n405 10.1505
R9850 VDD.n426 VDD.n425 10.1505
R9851 VDD.n324 VDD.n322 10.1505
R9852 VDD.n399 VDD.n307 10.1505
R9853 VDD.n396 VDD.n308 10.1505
R9854 VDD.n387 VDD.n311 10.1505
R9855 VDD.n388 VDD.n387 10.1505
R9856 VDD.n388 VDD.n306 10.1505
R9857 VDD.n391 VDD.n306 10.1505
R9858 VDD.n65 VDD.n63 10.1505
R9859 VDD.n72 VDD.n71 10.1505
R9860 VDD.n71 VDD.n61 10.1505
R9861 VDD.n75 VDD.n53 10.1505
R9862 VDD.n91 VDD.n53 10.1505
R9863 VDD.n91 VDD.n50 10.1505
R9864 VDD.n94 VDD.n50 10.1505
R9865 VDD.n69 VDD.n64 10.1505
R9866 VDD.n64 VDD.n55 10.1505
R9867 VDD.n55 VDD.n43 10.1505
R9868 VDD.n98 VDD.n43 10.1505
R9869 VDD.n85 VDD.n44 10.1505
R9870 VDD.n49 VDD.n48 10.1505
R9871 VDD.n82 VDD.n48 10.1505
R9872 VDD.n79 VDD.n56 10.1505
R9873 VDD.n90 VDD.n56 10.1505
R9874 VDD.n90 VDD.n57 10.1505
R9875 VDD.n84 VDD.n57 10.1505
R9876 VDD.n223 VDD.n202 7.3505
R9877 VDD.n449 VDD.n290 7.0005
R9878 VDD.n441 VDD.n440 7.0005
R9879 VDD.n340 VDD.n325 7.0005
R9880 VDD.n411 VDD.n299 7.0005
R9881 VDD.n393 VDD.n391 7.0005
R9882 VDD.n79 VDD.n60 7.0005
R9883 VDD.n86 VDD.n84 7.0005
R9884 VDD.n228 VDD.n227 6.78118
R9885 VDD.n425 VDD.n424 6.3005
R9886 VDD.n427 VDD.n426 6.3005
R9887 VDD.t12 VDD.n406 6.3005
R9888 VDD.n405 VDD.n300 6.3005
R9889 VDD.n445 VDD.n444 6.3005
R9890 VDD.n294 VDD 6.3005
R9891 VDD.n412 VDD.n411 6.3005
R9892 VDD.n420 VDD.n419 6.3005
R9893 VDD.n421 VDD 6.3005
R9894 VDD.n421 VDD.n289 6.3005
R9895 VDD.n423 VDD.n422 6.3005
R9896 VDD.n418 VDD.n417 6.3005
R9897 VDD.n416 VDD.n408 6.3005
R9898 VDD.n427 VDD.n408 6.3005
R9899 VDD VDD.n407 6.3005
R9900 VDD.t12 VDD.n407 6.3005
R9901 VDD.n415 VDD.n414 6.3005
R9902 VDD.n414 VDD.n300 6.3005
R9903 VDD.n413 VDD.n299 6.3005
R9904 VDD.n442 VDD.n299 6.3005
R9905 VDD.n341 VDD.n340 6.3005
R9906 VDD.n338 VDD 6.3005
R9907 VDD.n337 VDD.n336 6.3005
R9908 VDD.n440 VDD.n439 6.3005
R9909 VDD VDD.n438 6.3005
R9910 VDD.n437 VDD.n436 6.3005
R9911 VDD.n449 VDD.n448 6.3005
R9912 VDD.n451 VDD 6.3005
R9913 VDD.n452 VDD.n286 6.3005
R9914 VDD.n447 VDD.n290 6.3005
R9915 VDD.n290 VDD.n289 6.3005
R9916 VDD.n430 VDD.n427 6.3005
R9917 VDD.t12 VDD.n432 6.3005
R9918 VDD.n429 VDD.n300 6.3005
R9919 VDD.n391 VDD.n390 6.3005
R9920 VDD.n391 VDD.n295 6.3005
R9921 VDD.n389 VDD.n306 6.3005
R9922 VDD.n400 VDD.n306 6.3005
R9923 VDD VDD.n388 6.3005
R9924 VDD.n388 VDD.t36 6.3005
R9925 VDD.n387 VDD.n310 6.3005
R9926 VDD.n387 VDD.n386 6.3005
R9927 VDD.n315 VDD.n311 6.3005
R9928 VDD.n394 VDD.n393 6.3005
R9929 VDD VDD.n308 6.3005
R9930 VDD.n396 VDD.n395 6.3005
R9931 VDD.n320 VDD.n319 6.3005
R9932 VDD VDD.n314 6.3005
R9933 VDD.n314 VDD.n312 6.3005
R9934 VDD.n318 VDD.n317 6.3005
R9935 VDD.n400 VDD.n399 6.3005
R9936 VDD.n307 VDD.t36 6.3005
R9937 VDD.n386 VDD.n324 6.3005
R9938 VDD.n322 VDD 6.3005
R9939 VDD.n400 VDD.n305 6.3005
R9940 VDD VDD.n328 6.3005
R9941 VDD.n328 VDD.t36 6.3005
R9942 VDD.n386 VDD.n313 6.3005
R9943 VDD.n334 VDD.n333 6.3005
R9944 VDD.n330 VDD 6.3005
R9945 VDD.n330 VDD.n295 6.3005
R9946 VDD.n329 VDD.n301 6.3005
R9947 VDD.n403 VDD.n402 6.3005
R9948 VDD.n401 VDD.n302 6.3005
R9949 VDD.n401 VDD.n400 6.3005
R9950 VDD VDD.n304 6.3005
R9951 VDD.t36 VDD.n304 6.3005
R9952 VDD.n385 VDD.n384 6.3005
R9953 VDD.n386 VDD.n385 6.3005
R9954 VDD.n383 VDD.n325 6.3005
R9955 VDD.n325 VDD.n312 6.3005
R9956 VDD.n288 VDD.n287 6.3005
R9957 VDD.n427 VDD.n288 6.3005
R9958 VDD VDD.n433 6.3005
R9959 VDD.n433 VDD.t12 6.3005
R9960 VDD.n435 VDD.n434 6.3005
R9961 VDD.n435 VDD.n300 6.3005
R9962 VDD.n441 VDD.n404 6.3005
R9963 VDD.n442 VDD.n441 6.3005
R9964 VDD.n455 VDD.n454 6.3005
R9965 VDD.n94 VDD.n93 6.3005
R9966 VDD.n92 VDD.n50 6.3005
R9967 VDD.n50 VDD.n45 6.3005
R9968 VDD VDD.n91 6.3005
R9969 VDD.n91 VDD.t19 6.3005
R9970 VDD.n53 VDD.n52 6.3005
R9971 VDD.n54 VDD.n53 6.3005
R9972 VDD.n75 VDD.n74 6.3005
R9973 VDD.n73 VDD.n72 6.3005
R9974 VDD VDD.n71 6.3005
R9975 VDD.n77 VDD.n71 6.3005
R9976 VDD.n61 VDD.n59 6.3005
R9977 VDD.n60 VDD.n58 6.3005
R9978 VDD VDD.n65 6.3005
R9979 VDD.n66 VDD.n63 6.3005
R9980 VDD.n43 VDD.n42 6.3005
R9981 VDD.n45 VDD.n43 6.3005
R9982 VDD VDD.n55 6.3005
R9983 VDD.t19 VDD.n55 6.3005
R9984 VDD.n67 VDD.n64 6.3005
R9985 VDD.n64 VDD.n54 6.3005
R9986 VDD.n69 VDD.n68 6.3005
R9987 VDD.n83 VDD.n82 6.3005
R9988 VDD VDD.n48 6.3005
R9989 VDD.n96 VDD.n48 6.3005
R9990 VDD.n51 VDD.n49 6.3005
R9991 VDD.n88 VDD.n84 6.3005
R9992 VDD.n89 VDD.n57 6.3005
R9993 VDD.n57 VDD.n45 6.3005
R9994 VDD.n90 VDD 6.3005
R9995 VDD.t19 VDD.n90 6.3005
R9996 VDD.n81 VDD.n56 6.3005
R9997 VDD.n56 VDD.n54 6.3005
R9998 VDD.n80 VDD.n79 6.3005
R9999 VDD VDD.n85 6.3005
R10000 VDD.n87 VDD.n86 6.3005
R10001 VDD.n44 VDD.n41 6.3005
R10002 VDD.n99 VDD.n98 6.3005
R10003 VDD.n214 VDD.n213 6.3005
R10004 VDD.n212 VDD.n211 6.3005
R10005 VDD.n204 VDD.n202 6.3005
R10006 VDD.n223 VDD.n222 6.3005
R10007 VDD.n224 VDD.n223 6.3005
R10008 VDD.n221 VDD.n203 6.3005
R10009 VDD.n203 VDD.n201 6.3005
R10010 VDD.n220 VDD.n219 6.3005
R10011 VDD.n219 VDD.n218 6.3005
R10012 VDD.n206 VDD.n205 6.3005
R10013 VDD.n200 VDD.n198 6.3005
R10014 VDD.n201 VDD.n200 6.3005
R10015 VDD.n217 VDD.n216 6.3005
R10016 VDD.n218 VDD.n217 6.3005
R10017 VDD.n215 VDD.n208 6.3005
R10018 VDD.n225 VDD.n224 6.3005
R10019 VDD.n367 VDD.n366 5.80576
R10020 VDD.n226 VDD.n199 5.18619
R10021 VDD.n332 VDD.n331 5.06227
R10022 VDD.n443 VDD.n292 5.06227
R10023 VDD.n428 VDD.n297 5.06227
R10024 VDD.n398 VDD.n397 5.06227
R10025 VDD.n327 VDD.n326 5.06227
R10026 VDD.n587 VDD.n577 4.62839
R10027 VDD.n593 VDD.n592 4.62839
R10028 VDD.n372 VDD.n371 4.58103
R10029 VDD.n589 VDD.n577 4.5005
R10030 VDD.n592 VDD.n591 4.5005
R10031 VDD.n468 VDD.n274 4.5005
R10032 VDD.n817 VDD.n468 4.5005
R10033 VDD.n817 VDD.n471 4.5005
R10034 VDD.n817 VDD.n279 4.5005
R10035 VDD.n817 VDD.n473 4.5005
R10036 VDD.n817 VDD.n278 4.5005
R10037 VDD.n817 VDD.n475 4.5005
R10038 VDD.n817 VDD.n277 4.5005
R10039 VDD.n817 VDD.n816 4.5005
R10040 VDD.n817 VDD.n276 4.5005
R10041 VDD.n818 VDD.n274 4.5005
R10042 VDD.n818 VDD.n817 4.5005
R10043 VDD.n459 VDD.n458 4.5005
R10044 VDD.n459 VDD.n456 4.5005
R10045 VDD.n462 VDD.n456 4.5005
R10046 VDD.n463 VDD.n281 4.5005
R10047 VDD.n464 VDD.n463 4.5005
R10048 VDD.n465 VDD.n464 4.5005
R10049 VDD.n870 VDD.n820 4.5005
R10050 VDD.n870 VDD.n869 4.5005
R10051 VDD.n869 VDD.n828 4.5005
R10052 VDD.n869 VDD.n825 4.5005
R10053 VDD.n869 VDD.n830 4.5005
R10054 VDD.n869 VDD.n824 4.5005
R10055 VDD.n869 VDD.n832 4.5005
R10056 VDD.n869 VDD.n823 4.5005
R10057 VDD.n869 VDD.n834 4.5005
R10058 VDD.n869 VDD.n822 4.5005
R10059 VDD.n868 VDD.n820 4.5005
R10060 VDD.n869 VDD.n868 4.5005
R10061 VDD.n598 VDD.n597 4.14897
R10062 VDD.n119 VDD.n100 4.13212
R10063 VDD.n228 VDD.n197 4.0005
R10064 VDD.n202 VDD.n199 2.86464
R10065 VDD.n450 VDD.n449 2.81177
R10066 VDD.n429 VDD.n428 2.81177
R10067 VDD.n431 VDD.n430 2.81177
R10068 VDD.n440 VDD.n296 2.81177
R10069 VDD.n327 VDD.n313 2.81177
R10070 VDD.n340 VDD.n339 2.81177
R10071 VDD.n298 VDD.n294 2.81177
R10072 VDD.n405 VDD.n292 2.81177
R10073 VDD.n426 VDD.n293 2.81177
R10074 VDD.n406 VDD.n293 2.81177
R10075 VDD.n411 VDD.n298 2.81177
R10076 VDD.n339 VDD.n338 2.81177
R10077 VDD.n438 VDD.n296 2.81177
R10078 VDD.n451 VDD.n450 2.81177
R10079 VDD.n432 VDD.n431 2.81177
R10080 VDD.n323 VDD.n307 2.81177
R10081 VDD.n392 VDD.n308 2.81177
R10082 VDD.n393 VDD.n392 2.81177
R10083 VDD.n399 VDD.n398 2.81177
R10084 VDD.n324 VDD.n323 2.81177
R10085 VDD.n331 VDD.n305 2.81177
R10086 VDD.n62 VDD.n60 2.81177
R10087 VDD.n65 VDD.n62 2.81177
R10088 VDD.n86 VDD.n47 2.81177
R10089 VDD.n85 VDD.n47 2.81177
R10090 VDD.n658 VDD.t44 2.46086
R10091 VDD.n556 VDD.t42 2.46086
R10092 VDD.n124 VDD.t21 2.36071
R10093 VDD.n226 VDD.n225 2.32205
R10094 VDD.n213 VDD.n209 2.32205
R10095 VDD.n212 VDD.n210 2.32205
R10096 VDD.n210 VDD.n206 2.32205
R10097 VDD.n209 VDD.n208 2.32205
R10098 VDD.n461 VDD.n460 2.25705
R10099 VDD.n402 VDD.n303 2.251
R10100 VDD.n321 VDD.n320 2.251
R10101 VDD.n316 VDD.n311 2.251
R10102 VDD.n453 VDD.n452 2.251
R10103 VDD.n437 VDD.n297 2.251
R10104 VDD.n337 VDD.n326 2.251
R10105 VDD.n425 VDD.n409 2.251
R10106 VDD.n420 VDD.n410 2.251
R10107 VDD.n444 VDD.n443 2.251
R10108 VDD.n422 VDD.n409 2.251
R10109 VDD.n417 VDD.n410 2.251
R10110 VDD.n397 VDD.n396 2.251
R10111 VDD.n317 VDD.n316 2.251
R10112 VDD.n322 VDD.n321 2.251
R10113 VDD.n333 VDD.n332 2.251
R10114 VDD.n329 VDD.n303 2.251
R10115 VDD.n454 VDD.n453 2.251
R10116 VDD.n70 VDD.n63 2.251
R10117 VDD.n76 VDD.n75 2.251
R10118 VDD.n78 VDD.n61 2.251
R10119 VDD.n76 VDD.n72 2.251
R10120 VDD.n70 VDD.n69 2.251
R10121 VDD.n97 VDD.n44 2.251
R10122 VDD.n95 VDD.n94 2.251
R10123 VDD.n82 VDD.n46 2.251
R10124 VDD.n95 VDD.n49 2.251
R10125 VDD.n84 VDD.n46 2.251
R10126 VDD.n79 VDD.n78 2.251
R10127 VDD.n98 VDD.n97 2.251
R10128 VDD.n462 VDD.n461 2.24475
R10129 VDD.n467 VDD.n280 2.24475
R10130 VDD.n457 VDD.n285 2.24475
R10131 VDD.n466 VDD.n281 2.24405
R10132 VDD.n283 VDD.n282 2.24405
R10133 VDD.n813 VDD.n479 2.24304
R10134 VDD.n470 VDD.n274 2.24304
R10135 VDD.n813 VDD.n478 2.24304
R10136 VDD.n472 VDD.n274 2.24304
R10137 VDD.n813 VDD.n477 2.24304
R10138 VDD.n474 VDD.n274 2.24304
R10139 VDD.n814 VDD.n813 2.24304
R10140 VDD.n815 VDD.n274 2.24304
R10141 VDD.n813 VDD.n273 2.24304
R10142 VDD.n827 VDD.n820 2.24304
R10143 VDD.n866 VDD.n819 2.24304
R10144 VDD.n829 VDD.n820 2.24304
R10145 VDD.n866 VDD.n863 2.24304
R10146 VDD.n831 VDD.n820 2.24304
R10147 VDD.n866 VDD.n864 2.24304
R10148 VDD.n833 VDD.n820 2.24304
R10149 VDD.n866 VDD.n865 2.24304
R10150 VDD.n867 VDD.n866 2.24304
R10151 VDD.n362 VDD.t1 2.12386
R10152 VDD.n581 VDD.t9 2.12292
R10153 VDD.n871 VDD.n818 2.10965
R10154 VDD.n590 VDD.t57 2.08373
R10155 VDD.n409 VDD.n289 2.026
R10156 VDD.n443 VDD.n442 2.026
R10157 VDD.n410 VDD.n289 2.026
R10158 VDD.n326 VDD.n312 2.026
R10159 VDD.n442 VDD.n297 2.026
R10160 VDD.n453 VDD.n289 2.026
R10161 VDD.n316 VDD.n312 2.026
R10162 VDD.n321 VDD.n312 2.026
R10163 VDD.n397 VDD.n295 2.026
R10164 VDD.n332 VDD.n295 2.026
R10165 VDD.n303 VDD.n295 2.026
R10166 VDD.n96 VDD.n95 2.026
R10167 VDD.n77 VDD.n76 2.026
R10168 VDD.n78 VDD.n77 2.026
R10169 VDD.n77 VDD.n70 2.026
R10170 VDD.n96 VDD.n46 2.026
R10171 VDD.n97 VDD.n96 2.026
R10172 VDD.n209 VDD.n207 1.99047
R10173 VDD.n210 VDD.n207 1.99047
R10174 VDD.n227 VDD.n226 1.99047
R10175 VDD.n575 VDD.t62 1.96281
R10176 VDD.n873 VDD.t7 1.96281
R10177 VDD.n272 VDD.t25 1.96281
R10178 VDD.n126 VDD.t55 1.96281
R10179 VDD.n40 VDD.t48 1.96281
R10180 VDD.n1 VDD.t53 1.96281
R10181 VDD.n929 VDD.t59 1.96281
R10182 VDD.n196 VDD.t23 1.96281
R10183 VDD.n576 VDD.t3 1.92255
R10184 VDD.n586 VDD.t5 1.92255
R10185 VDD.n582 VDD.t11 1.92255
R10186 VDD.n195 VDD.n194 1.8507
R10187 VDD.n926 VDD.n925 1.8507
R10188 VDD.n877 VDD.n876 1.8228
R10189 VDD.n375 VDD.t45 1.81731
R10190 VDD.n358 VDD.t13 1.81731
R10191 VDD.n349 VDD.t63 1.81731
R10192 VDD.n365 VDD.t0 1.81731
R10193 VDD.n663 VDD.n662 1.80879
R10194 VDD.n650 VDD.n649 1.8024
R10195 VDD.n128 VDD.n127 1.8005
R10196 VDD.n651 VDD.t16 1.78389
R10197 VDD.n659 VDD.t29 1.78389
R10198 VDD VDD.n293 1.74562
R10199 VDD VDD.n292 1.74562
R10200 VDD.n442 VDD.n298 1.74562
R10201 VDD.n339 VDD.n312 1.74562
R10202 VDD.n442 VDD.n296 1.74562
R10203 VDD.n450 VDD.n289 1.74562
R10204 VDD.n431 VDD 1.74562
R10205 VDD.n428 VDD 1.74562
R10206 VDD.n392 VDD.n295 1.74562
R10207 VDD.n398 VDD 1.74562
R10208 VDD.n323 VDD 1.74562
R10209 VDD.n331 VDD 1.74562
R10210 VDD VDD.n327 1.74562
R10211 VDD.n77 VDD.n62 1.74562
R10212 VDD.n96 VDD.n47 1.74562
R10213 VDD.n657 VDD.n656 1.73286
R10214 VDD.n588 VDD.n578 1.72301
R10215 VDD.n224 VDD.n199 1.71918
R10216 VDD.n872 VDD.n871 1.70597
R10217 VDD.n344 VDD.t64 1.58219
R10218 VDD.n346 VDD.t14 1.58219
R10219 VDD.n380 VDD.t46 1.58219
R10220 VDD.n585 VDD.n584 1.5755
R10221 VDD.n596 VDD.n595 1.5755
R10222 VDD.n875 VDD.n874 1.5755
R10223 VDD.n928 VDD.n927 1.5755
R10224 VDD.n232 VDD.n231 1.5755
R10225 VDD.n599 VDD.n598 1.50189
R10226 VDD.n615 VDD.n598 1.50166
R10227 VDD.n235 VDD.n234 1.50061
R10228 VDD.n130 VDD.n129 1.46392
R10229 VDD.n229 VDD.t51 1.36414
R10230 VDD.n382 VDD.n381 1.32326
R10231 VDD VDD.n123 1.27477
R10232 VDD.n653 VDD.n652 1.26489
R10233 VDD.n655 VDD.n654 1.26489
R10234 VDD.n377 VDD.n376 1.2605
R10235 VDD.n354 VDD.n353 1.2605
R10236 VDD.n348 VDD.n347 1.2605
R10237 VDD.n361 VDD.n360 1.2605
R10238 VDD.n123 VDD.t20 1.24589
R10239 VDD.n364 VDD.n363 1.15029
R10240 VDD.n926 VDD.n1 1.10418
R10241 VDD.n196 VDD.n195 1.10418
R10242 VDD.n876 VDD.n272 1.1
R10243 VDD.n370 VDD.n344 1.07633
R10244 VDD.n368 VDD.n346 1.07633
R10245 VDD.n381 VDD.n380 1.07633
R10246 VDD.n129 VDD.n40 1.06559
R10247 VDD.n373 VDD.n372 1.06155
R10248 VDD.n371 VDD.n343 1.06155
R10249 VDD.n369 VDD.n345 1.06155
R10250 VDD.n367 VDD.n359 1.06155
R10251 VDD.n366 VDD.n360 0.973921
R10252 VDD.n377 VDD.n373 0.964726
R10253 VDD.n353 VDD.n343 0.964726
R10254 VDD.n359 VDD.n347 0.964726
R10255 VDD.n120 VDD.n119 0.921424
R10256 VDD.n229 VDD 0.869566
R10257 VDD.n234 VDD.n0 0.861978
R10258 VDD.n125 VDD.n120 0.857799
R10259 VDD.n234 VDD.n233 0.788
R10260 VDD.n662 VDD.n556 0.756026
R10261 VDD.n656 VDD.t38 0.7285
R10262 VDD.n656 VDD.t40 0.7285
R10263 VDD.n468 VDD.n467 0.671
R10264 VDD.n651 VDD.n650 0.651808
R10265 VDD.n580 VDD.n579 0.6005
R10266 VDD.n230 VDD.n229 0.600169
R10267 VDD.n356 VDD.n345 0.573227
R10268 VDD.n357 VDD.n356 0.573227
R10269 VDD.n374 VDD.n342 0.573227
R10270 VDD.n351 VDD.n345 0.557079
R10271 VDD.n378 VDD.n342 0.557079
R10272 VDD.n368 VDD.n367 0.555895
R10273 VDD.n371 VDD.n370 0.555895
R10274 VDD.n381 VDD.n372 0.555895
R10275 VDD.n653 VDD.n651 0.545794
R10276 VDD.n655 VDD.n653 0.545794
R10277 VDD.n658 VDD.n657 0.545794
R10278 VDD.n657 VDD.n556 0.545794
R10279 VDD.n352 VDD.n344 0.542091
R10280 VDD.n350 VDD.n346 0.542091
R10281 VDD.n380 VDD.n379 0.542091
R10282 VDD.n119 VDD.n118 0.541547
R10283 VDD.n652 VDD.t35 0.5205
R10284 VDD.n652 VDD.t31 0.5205
R10285 VDD.n654 VDD.t18 0.5205
R10286 VDD.n654 VDD.t27 0.5205
R10287 VDD.n813 VDD.n812 0.456899
R10288 VDD.n860 VDD.n820 0.456899
R10289 VDD.n859 VDD.n835 0.4505
R10290 VDD.n858 VDD.n857 0.4505
R10291 VDD.n856 VDD.n836 0.4505
R10292 VDD.n853 VDD.n852 0.4505
R10293 VDD.n851 VDD.n838 0.4505
R10294 VDD.n850 VDD.n849 0.4505
R10295 VDD.n840 VDD.n839 0.4505
R10296 VDD.n845 VDD.n844 0.4505
R10297 VDD.n843 VDD.n842 0.4505
R10298 VDD.n270 VDD.n269 0.4505
R10299 VDD.n880 VDD.n879 0.4505
R10300 VDD.n881 VDD.n268 0.4505
R10301 VDD.n883 VDD.n882 0.4505
R10302 VDD.n266 VDD.n265 0.4505
R10303 VDD.n888 VDD.n887 0.4505
R10304 VDD.n889 VDD.n264 0.4505
R10305 VDD.n891 VDD.n890 0.4505
R10306 VDD.n262 VDD.n261 0.4505
R10307 VDD.n896 VDD.n895 0.4505
R10308 VDD.n897 VDD.n260 0.4505
R10309 VDD.n899 VDD.n898 0.4505
R10310 VDD.n258 VDD.n257 0.4505
R10311 VDD.n904 VDD.n903 0.4505
R10312 VDD.n905 VDD.n256 0.4505
R10313 VDD.n907 VDD.n906 0.4505
R10314 VDD.n254 VDD.n253 0.4505
R10315 VDD.n912 VDD.n911 0.4505
R10316 VDD.n913 VDD.n252 0.4505
R10317 VDD.n915 VDD.n914 0.4505
R10318 VDD.n250 VDD.n249 0.4505
R10319 VDD.n920 VDD.n919 0.4505
R10320 VDD.n921 VDD.n5 0.4505
R10321 VDD.n923 VDD.n922 0.4505
R10322 VDD.n248 VDD.n4 0.4505
R10323 VDD.n247 VDD.n246 0.4505
R10324 VDD.n7 VDD.n6 0.4505
R10325 VDD.n242 VDD.n241 0.4505
R10326 VDD.n240 VDD.n9 0.4505
R10327 VDD.n239 VDD.n238 0.4505
R10328 VDD.n11 VDD.n10 0.4505
R10329 VDD.n181 VDD.n180 0.4505
R10330 VDD.n182 VDD.n179 0.4505
R10331 VDD.n184 VDD.n183 0.4505
R10332 VDD.n177 VDD.n176 0.4505
R10333 VDD.n189 VDD.n188 0.4505
R10334 VDD.n190 VDD.n16 0.4505
R10335 VDD.n115 VDD.n114 0.4505
R10336 VDD.n113 VDD.n103 0.4505
R10337 VDD.n112 VDD.n111 0.4505
R10338 VDD.n107 VDD.n104 0.4505
R10339 VDD.n106 VDD.n105 0.4505
R10340 VDD.n38 VDD.n37 0.4505
R10341 VDD.n134 VDD.n133 0.4505
R10342 VDD.n135 VDD.n36 0.4505
R10343 VDD.n137 VDD.n136 0.4505
R10344 VDD.n34 VDD.n33 0.4505
R10345 VDD.n142 VDD.n141 0.4505
R10346 VDD.n143 VDD.n32 0.4505
R10347 VDD.n145 VDD.n144 0.4505
R10348 VDD.n30 VDD.n29 0.4505
R10349 VDD.n150 VDD.n149 0.4505
R10350 VDD.n151 VDD.n28 0.4505
R10351 VDD.n153 VDD.n152 0.4505
R10352 VDD.n26 VDD.n25 0.4505
R10353 VDD.n158 VDD.n157 0.4505
R10354 VDD.n159 VDD.n24 0.4505
R10355 VDD.n161 VDD.n160 0.4505
R10356 VDD.n22 VDD.n21 0.4505
R10357 VDD.n166 VDD.n165 0.4505
R10358 VDD.n167 VDD.n20 0.4505
R10359 VDD.n169 VDD.n168 0.4505
R10360 VDD.n18 VDD.n17 0.4505
R10361 VDD.n174 VDD.n173 0.4505
R10362 VDD.n175 VDD.n15 0.4505
R10363 VDD.n192 VDD.n191 0.4505
R10364 VDD.n811 VDD.n810 0.4505
R10365 VDD.n809 VDD.n481 0.4505
R10366 VDD.n808 VDD.n482 0.4505
R10367 VDD.n805 VDD.n804 0.4505
R10368 VDD.n803 VDD.n484 0.4505
R10369 VDD.n802 VDD.n801 0.4505
R10370 VDD.n486 VDD.n485 0.4505
R10371 VDD.n797 VDD.n796 0.4505
R10372 VDD.n795 VDD.n488 0.4505
R10373 VDD.n794 VDD.n793 0.4505
R10374 VDD.n490 VDD.n489 0.4505
R10375 VDD.n789 VDD.n788 0.4505
R10376 VDD.n787 VDD.n492 0.4505
R10377 VDD.n786 VDD.n785 0.4505
R10378 VDD.n494 VDD.n493 0.4505
R10379 VDD.n781 VDD.n780 0.4505
R10380 VDD.n779 VDD.n496 0.4505
R10381 VDD.n778 VDD.n777 0.4505
R10382 VDD.n498 VDD.n497 0.4505
R10383 VDD.n773 VDD.n772 0.4505
R10384 VDD.n771 VDD.n500 0.4505
R10385 VDD.n770 VDD.n769 0.4505
R10386 VDD.n502 VDD.n501 0.4505
R10387 VDD.n765 VDD.n764 0.4505
R10388 VDD.n763 VDD.n504 0.4505
R10389 VDD.n762 VDD.n761 0.4505
R10390 VDD.n506 VDD.n505 0.4505
R10391 VDD.n757 VDD.n756 0.4505
R10392 VDD.n755 VDD.n508 0.4505
R10393 VDD.n754 VDD.n753 0.4505
R10394 VDD.n510 VDD.n509 0.4505
R10395 VDD.n749 VDD.n748 0.4505
R10396 VDD.n747 VDD.n512 0.4505
R10397 VDD.n746 VDD.n745 0.4505
R10398 VDD.n514 VDD.n513 0.4505
R10399 VDD.n741 VDD.n740 0.4505
R10400 VDD.n739 VDD.n516 0.4505
R10401 VDD.n738 VDD.n737 0.4505
R10402 VDD.n518 VDD.n517 0.4505
R10403 VDD.n733 VDD.n732 0.4505
R10404 VDD.n731 VDD.n520 0.4505
R10405 VDD.n730 VDD.n729 0.4505
R10406 VDD.n522 VDD.n521 0.4505
R10407 VDD.n725 VDD.n724 0.4505
R10408 VDD.n723 VDD.n524 0.4505
R10409 VDD.n722 VDD.n721 0.4505
R10410 VDD.n526 VDD.n525 0.4505
R10411 VDD.n717 VDD.n716 0.4505
R10412 VDD.n715 VDD.n528 0.4505
R10413 VDD.n714 VDD.n713 0.4505
R10414 VDD.n530 VDD.n529 0.4505
R10415 VDD.n709 VDD.n708 0.4505
R10416 VDD.n707 VDD.n532 0.4505
R10417 VDD.n706 VDD.n705 0.4505
R10418 VDD.n534 VDD.n533 0.4505
R10419 VDD.n701 VDD.n700 0.4505
R10420 VDD.n699 VDD.n536 0.4505
R10421 VDD.n698 VDD.n697 0.4505
R10422 VDD.n538 VDD.n537 0.4505
R10423 VDD.n693 VDD.n692 0.4505
R10424 VDD.n691 VDD.n540 0.4505
R10425 VDD.n690 VDD.n689 0.4505
R10426 VDD.n542 VDD.n541 0.4505
R10427 VDD.n685 VDD.n684 0.4505
R10428 VDD.n683 VDD.n544 0.4505
R10429 VDD.n682 VDD.n681 0.4505
R10430 VDD.n546 VDD.n545 0.4505
R10431 VDD.n677 VDD.n676 0.4505
R10432 VDD.n675 VDD.n548 0.4505
R10433 VDD.n674 VDD.n673 0.4505
R10434 VDD.n550 VDD.n549 0.4505
R10435 VDD.n669 VDD.n668 0.4505
R10436 VDD.n667 VDD.n552 0.4505
R10437 VDD.n646 VDD.n645 0.4505
R10438 VDD.n644 VDD.n559 0.4505
R10439 VDD.n643 VDD.n642 0.4505
R10440 VDD.n561 VDD.n560 0.4505
R10441 VDD.n638 VDD.n637 0.4505
R10442 VDD.n636 VDD.n564 0.4505
R10443 VDD.n635 VDD.n634 0.4505
R10444 VDD.n566 VDD.n565 0.4505
R10445 VDD.n630 VDD.n629 0.4505
R10446 VDD.n628 VDD.n568 0.4505
R10447 VDD.n627 VDD.n626 0.4505
R10448 VDD.n570 VDD.n569 0.4505
R10449 VDD.n622 VDD.n621 0.4505
R10450 VDD.n620 VDD.n572 0.4505
R10451 VDD.n619 VDD.n618 0.4505
R10452 VDD.n574 VDD.n573 0.4505
R10453 VDD.n613 VDD.n612 0.4505
R10454 VDD.n611 VDD.n600 0.4505
R10455 VDD.n610 VDD.n609 0.4505
R10456 VDD.n602 VDD.n601 0.4505
R10457 VDD.n605 VDD.n604 0.4505
R10458 VDD.n554 VDD.n553 0.4505
R10459 VDD.n666 VDD.n665 0.4505
R10460 VDD.n809 VDD.n275 0.4505
R10461 VDD.n480 VDD.n476 0.4505
R10462 VDD.n552 VDD.n551 0.4505
R10463 VDD.n670 VDD.n669 0.4505
R10464 VDD.n671 VDD.n550 0.4505
R10465 VDD.n673 VDD.n672 0.4505
R10466 VDD.n548 VDD.n547 0.4505
R10467 VDD.n678 VDD.n677 0.4505
R10468 VDD.n679 VDD.n546 0.4505
R10469 VDD.n681 VDD.n680 0.4505
R10470 VDD.n544 VDD.n543 0.4505
R10471 VDD.n686 VDD.n685 0.4505
R10472 VDD.n687 VDD.n542 0.4505
R10473 VDD.n689 VDD.n688 0.4505
R10474 VDD.n540 VDD.n539 0.4505
R10475 VDD.n694 VDD.n693 0.4505
R10476 VDD.n695 VDD.n538 0.4505
R10477 VDD.n697 VDD.n696 0.4505
R10478 VDD.n536 VDD.n535 0.4505
R10479 VDD.n702 VDD.n701 0.4505
R10480 VDD.n703 VDD.n534 0.4505
R10481 VDD.n705 VDD.n704 0.4505
R10482 VDD.n532 VDD.n531 0.4505
R10483 VDD.n710 VDD.n709 0.4505
R10484 VDD.n711 VDD.n530 0.4505
R10485 VDD.n713 VDD.n712 0.4505
R10486 VDD.n528 VDD.n527 0.4505
R10487 VDD.n718 VDD.n717 0.4505
R10488 VDD.n719 VDD.n526 0.4505
R10489 VDD.n721 VDD.n720 0.4505
R10490 VDD.n524 VDD.n523 0.4505
R10491 VDD.n726 VDD.n725 0.4505
R10492 VDD.n727 VDD.n522 0.4505
R10493 VDD.n729 VDD.n728 0.4505
R10494 VDD.n520 VDD.n519 0.4505
R10495 VDD.n734 VDD.n733 0.4505
R10496 VDD.n735 VDD.n518 0.4505
R10497 VDD.n737 VDD.n736 0.4505
R10498 VDD.n516 VDD.n515 0.4505
R10499 VDD.n742 VDD.n741 0.4505
R10500 VDD.n743 VDD.n514 0.4505
R10501 VDD.n745 VDD.n744 0.4505
R10502 VDD.n512 VDD.n511 0.4505
R10503 VDD.n750 VDD.n749 0.4505
R10504 VDD.n751 VDD.n510 0.4505
R10505 VDD.n753 VDD.n752 0.4505
R10506 VDD.n508 VDD.n507 0.4505
R10507 VDD.n758 VDD.n757 0.4505
R10508 VDD.n759 VDD.n506 0.4505
R10509 VDD.n761 VDD.n760 0.4505
R10510 VDD.n504 VDD.n503 0.4505
R10511 VDD.n766 VDD.n765 0.4505
R10512 VDD.n767 VDD.n502 0.4505
R10513 VDD.n769 VDD.n768 0.4505
R10514 VDD.n500 VDD.n499 0.4505
R10515 VDD.n774 VDD.n773 0.4505
R10516 VDD.n775 VDD.n498 0.4505
R10517 VDD.n777 VDD.n776 0.4505
R10518 VDD.n496 VDD.n495 0.4505
R10519 VDD.n782 VDD.n781 0.4505
R10520 VDD.n783 VDD.n494 0.4505
R10521 VDD.n785 VDD.n784 0.4505
R10522 VDD.n492 VDD.n491 0.4505
R10523 VDD.n790 VDD.n789 0.4505
R10524 VDD.n791 VDD.n490 0.4505
R10525 VDD.n793 VDD.n792 0.4505
R10526 VDD.n488 VDD.n487 0.4505
R10527 VDD.n798 VDD.n797 0.4505
R10528 VDD.n799 VDD.n486 0.4505
R10529 VDD.n801 VDD.n800 0.4505
R10530 VDD.n484 VDD.n483 0.4505
R10531 VDD.n806 VDD.n805 0.4505
R10532 VDD.n808 VDD.n807 0.4505
R10533 VDD.n810 VDD.n469 0.4505
R10534 VDD.n648 VDD.n647 0.4505
R10535 VDD.n646 VDD.n558 0.4505
R10536 VDD.n562 VDD.n559 0.4505
R10537 VDD.n642 VDD.n641 0.4505
R10538 VDD.n640 VDD.n561 0.4505
R10539 VDD.n639 VDD.n638 0.4505
R10540 VDD.n564 VDD.n563 0.4505
R10541 VDD.n634 VDD.n633 0.4505
R10542 VDD.n632 VDD.n566 0.4505
R10543 VDD.n631 VDD.n630 0.4505
R10544 VDD.n568 VDD.n567 0.4505
R10545 VDD.n626 VDD.n625 0.4505
R10546 VDD.n624 VDD.n570 0.4505
R10547 VDD.n623 VDD.n622 0.4505
R10548 VDD.n572 VDD.n571 0.4505
R10549 VDD.n618 VDD.n617 0.4505
R10550 VDD.n616 VDD.n574 0.4505
R10551 VDD.n614 VDD.n613 0.4505
R10552 VDD.n603 VDD.n600 0.4505
R10553 VDD.n609 VDD.n608 0.4505
R10554 VDD.n607 VDD.n602 0.4505
R10555 VDD.n606 VDD.n605 0.4505
R10556 VDD.n555 VDD.n554 0.4505
R10557 VDD.n665 VDD.n664 0.4505
R10558 VDD.n862 VDD.n861 0.4505
R10559 VDD.n835 VDD.n826 0.4505
R10560 VDD.n857 VDD.n821 0.4505
R10561 VDD.n856 VDD.n855 0.4505
R10562 VDD.n854 VDD.n853 0.4505
R10563 VDD.n838 VDD.n837 0.4505
R10564 VDD.n849 VDD.n848 0.4505
R10565 VDD.n847 VDD.n840 0.4505
R10566 VDD.n846 VDD.n845 0.4505
R10567 VDD.n842 VDD.n841 0.4505
R10568 VDD.n271 VDD.n270 0.4505
R10569 VDD.n879 VDD.n878 0.4505
R10570 VDD.n268 VDD.n267 0.4505
R10571 VDD.n884 VDD.n883 0.4505
R10572 VDD.n885 VDD.n266 0.4505
R10573 VDD.n887 VDD.n886 0.4505
R10574 VDD.n264 VDD.n263 0.4505
R10575 VDD.n892 VDD.n891 0.4505
R10576 VDD.n893 VDD.n262 0.4505
R10577 VDD.n895 VDD.n894 0.4505
R10578 VDD.n260 VDD.n259 0.4505
R10579 VDD.n900 VDD.n899 0.4505
R10580 VDD.n901 VDD.n258 0.4505
R10581 VDD.n903 VDD.n902 0.4505
R10582 VDD.n256 VDD.n255 0.4505
R10583 VDD.n908 VDD.n907 0.4505
R10584 VDD.n909 VDD.n254 0.4505
R10585 VDD.n911 VDD.n910 0.4505
R10586 VDD.n252 VDD.n251 0.4505
R10587 VDD.n916 VDD.n915 0.4505
R10588 VDD.n917 VDD.n250 0.4505
R10589 VDD.n919 VDD.n918 0.4505
R10590 VDD.n5 VDD.n3 0.4505
R10591 VDD.n924 VDD.n923 0.4505
R10592 VDD.n4 VDD.n2 0.4505
R10593 VDD.n246 VDD.n245 0.4505
R10594 VDD.n244 VDD.n7 0.4505
R10595 VDD.n243 VDD.n242 0.4505
R10596 VDD.n9 VDD.n8 0.4505
R10597 VDD.n238 VDD.n237 0.4505
R10598 VDD.n16 VDD.n14 0.4505
R10599 VDD.n188 VDD.n187 0.4505
R10600 VDD.n186 VDD.n177 0.4505
R10601 VDD.n185 VDD.n184 0.4505
R10602 VDD.n179 VDD.n178 0.4505
R10603 VDD.n180 VDD.n12 0.4505
R10604 VDD.n236 VDD.n11 0.4505
R10605 VDD.n117 VDD.n116 0.4505
R10606 VDD.n115 VDD.n102 0.4505
R10607 VDD.n108 VDD.n103 0.4505
R10608 VDD.n111 VDD.n110 0.4505
R10609 VDD.n109 VDD.n107 0.4505
R10610 VDD.n106 VDD.n39 0.4505
R10611 VDD.n131 VDD.n38 0.4505
R10612 VDD.n133 VDD.n132 0.4505
R10613 VDD.n36 VDD.n35 0.4505
R10614 VDD.n138 VDD.n137 0.4505
R10615 VDD.n139 VDD.n34 0.4505
R10616 VDD.n141 VDD.n140 0.4505
R10617 VDD.n32 VDD.n31 0.4505
R10618 VDD.n146 VDD.n145 0.4505
R10619 VDD.n147 VDD.n30 0.4505
R10620 VDD.n149 VDD.n148 0.4505
R10621 VDD.n28 VDD.n27 0.4505
R10622 VDD.n154 VDD.n153 0.4505
R10623 VDD.n155 VDD.n26 0.4505
R10624 VDD.n157 VDD.n156 0.4505
R10625 VDD.n24 VDD.n23 0.4505
R10626 VDD.n162 VDD.n161 0.4505
R10627 VDD.n163 VDD.n22 0.4505
R10628 VDD.n165 VDD.n164 0.4505
R10629 VDD.n20 VDD.n19 0.4505
R10630 VDD.n170 VDD.n169 0.4505
R10631 VDD.n171 VDD.n18 0.4505
R10632 VDD.n173 VDD.n172 0.4505
R10633 VDD.n15 VDD.n13 0.4505
R10634 VDD.n193 VDD.n192 0.4505
R10635 VDD.n661 VDD.n660 0.406952
R10636 VDD.n383 VDD.n382 0.397872
R10637 VDD.n121 VDD.n120 0.39425
R10638 VDD.n122 VDD.n121 0.39425
R10639 VDD.n583 VDD.n581 0.341837
R10640 VDD.n874 VDD.n272 0.296971
R10641 VDD.n928 VDD.n1 0.296971
R10642 VDD.n231 VDD.n196 0.296971
R10643 VDD.n127 VDD.n126 0.277118
R10644 VDD.n595 VDD.n575 0.273147
R10645 VDD.n447 VDD.n446 0.273
R10646 VDD.n127 VDD.n40 0.269176
R10647 VDD.n369 VDD.n368 0.264579
R10648 VDD.n370 VDD.n369 0.255105
R10649 VDD.n873 VDD 0.250647
R10650 VDD.n230 VDD 0.250647
R10651 VDD VDD.n929 0.250647
R10652 VDD.n874 VDD.n873 0.249324
R10653 VDD.n929 VDD.n928 0.249324
R10654 VDD.n231 VDD.n230 0.249324
R10655 VDD.n125 VDD.n124 0.241382
R10656 VDD.n363 VDD.n362 0.240059
R10657 VDD.n860 VDD.n859 0.231338
R10658 VDD.n812 VDD.n811 0.231338
R10659 VDD VDD.n655 0.226824
R10660 VDD.n424 VDD.n284 0.22175
R10661 VDD.n376 VDD.n375 0.212524
R10662 VDD.n354 VDD.n349 0.212524
R10663 VDD.n358 VDD.n348 0.212524
R10664 VDD.n365 VDD.n361 0.212524
R10665 VDD.n595 VDD.n594 0.208294
R10666 VDD.n660 VDD.n659 0.196382
R10667 VDD.n351 VDD.n350 0.195059
R10668 VDD.n379 VDD.n378 0.195059
R10669 VDD.n404 VDD.n403 0.187099
R10670 VDD.n352 VDD.n351 0.184471
R10671 VDD.n597 VDD.n575 0.181824
R10672 VDD.n446 VDD.n291 0.176791
R10673 VDD.n220 VDD.n205 0.1505
R10674 VDD.n222 VDD.n221 0.1505
R10675 VDD.n216 VDD.n215 0.1505
R10676 VDD.n463 VDD.n462 0.149225
R10677 VDD.n341 VDD 0.1455
R10678 VDD.n336 VDD 0.1455
R10679 VDD.n439 VDD 0.1455
R10680 VDD VDD.n436 0.1455
R10681 VDD.n445 VDD 0.1455
R10682 VDD.n412 VDD 0.1455
R10683 VDD.n415 VDD.n413 0.1455
R10684 VDD VDD.n415 0.1455
R10685 VDD.n416 VDD 0.1455
R10686 VDD.n418 VDD.n416 0.1455
R10687 VDD VDD.n286 0.1455
R10688 VDD.n448 VDD 0.1455
R10689 VDD.n448 VDD.n447 0.1455
R10690 VDD.n424 VDD.n423 0.1455
R10691 VDD.n423 VDD 0.1455
R10692 VDD.n419 VDD 0.1455
R10693 VDD.n315 VDD.n310 0.1455
R10694 VDD VDD.n310 0.1455
R10695 VDD.n389 VDD 0.1455
R10696 VDD.n390 VDD.n389 0.1455
R10697 VDD.n395 VDD 0.1455
R10698 VDD VDD.n394 0.1455
R10699 VDD.n319 VDD 0.1455
R10700 VDD VDD.n318 0.1455
R10701 VDD VDD.n301 0.1455
R10702 VDD.n334 VDD 0.1455
R10703 VDD VDD.n58 0.1455
R10704 VDD.n66 VDD 0.1455
R10705 VDD.n73 VDD 0.1455
R10706 VDD VDD.n59 0.1455
R10707 VDD VDD.n51 0.1455
R10708 VDD.n83 VDD 0.1455
R10709 VDD.n74 VDD.n52 0.1455
R10710 VDD VDD.n52 0.1455
R10711 VDD.n92 VDD 0.1455
R10712 VDD.n93 VDD.n92 0.1455
R10713 VDD.n68 VDD.n67 0.1455
R10714 VDD.n67 VDD 0.1455
R10715 VDD VDD.n42 0.1455
R10716 VDD.n81 VDD.n80 0.1455
R10717 VDD VDD.n81 0.1455
R10718 VDD VDD.n89 0.1455
R10719 VDD.n89 VDD.n88 0.1455
R10720 VDD.n87 VDD 0.1455
R10721 VDD VDD.n41 0.143658
R10722 VDD.n126 VDD 0.138147
R10723 VDD.n581 VDD 0.1355
R10724 VDD.n592 VDD.n577 0.128395
R10725 VDD.n659 VDD.n658 0.127559
R10726 VDD.n871 VDD.n870 0.1238
R10727 VDD.n660 VDD 0.123588
R10728 VDD.n227 VDD.n198 0.1235
R10729 VDD.n379 VDD.n377 0.113
R10730 VDD.n353 VDD.n352 0.113
R10731 VDD.n350 VDD.n347 0.113
R10732 VDD.n362 VDD.n360 0.113
R10733 VDD.n649 VDD.n557 0.107523
R10734 VDD.n436 VDD 0.107483
R10735 VDD VDD.n445 0.107483
R10736 VDD.n222 VDD.n204 0.1055
R10737 VDD.n215 VDD.n214 0.1055
R10738 VDD.n211 VDD.n205 0.1055
R10739 VDD.n383 VDD.n341 0.1005
R10740 VDD.n336 VDD.n335 0.1005
R10741 VDD.n439 VDD.n404 0.1005
R10742 VDD.n413 VDD.n412 0.1005
R10743 VDD.n455 VDD.n286 0.1005
R10744 VDD.n419 VDD.n418 0.1005
R10745 VDD.n395 VDD.n309 0.1005
R10746 VDD.n394 VDD.n390 0.1005
R10747 VDD.n319 VDD.n309 0.1005
R10748 VDD.n318 VDD.n315 0.1005
R10749 VDD.n403 VDD.n301 0.1005
R10750 VDD.n335 VDD.n334 0.1005
R10751 VDD.n80 VDD.n58 0.1005
R10752 VDD.n68 VDD.n66 0.1005
R10753 VDD.n74 VDD.n73 0.1005
R10754 VDD.n80 VDD.n59 0.1005
R10755 VDD.n93 VDD.n51 0.1005
R10756 VDD.n88 VDD.n83 0.1005
R10757 VDD.n99 VDD.n42 0.1005
R10758 VDD.n88 VDD.n87 0.1005
R10759 VDD.n456 VDD.n455 0.091309
R10760 VDD.n645 VDD.n557 0.0896854
R10761 VDD.n464 VDD.n284 0.0840281
R10762 VDD.n204 VDD 0.0755
R10763 VDD VDD.n220 0.0755
R10764 VDD.n221 VDD 0.0755
R10765 VDD.n214 VDD 0.0755
R10766 VDD.n211 VDD 0.0755
R10767 VDD.n216 VDD 0.0755
R10768 VDD VDD.n198 0.0755
R10769 VDD.n100 VDD.n41 0.0739211
R10770 VDD.n118 VDD.n101 0.0699284
R10771 VDD.n100 VDD.n99 0.0644474
R10772 VDD.n124 VDD 0.0627059
R10773 VDD VDD.n125 0.0627059
R10774 VDD.n114 VDD.n101 0.0585915
R10775 VDD.n446 VDD.n284 0.05175
R10776 VDD.n227 VDD 0.0455
R10777 VDD.n446 VDD 0.0427845
R10778 VDD.n446 VDD 0.0427845
R10779 VDD VDD.n872 0.0402059
R10780 VDD VDD.n0 0.0402059
R10781 VDD VDD.n0 0.0402059
R10782 VDD.n586 VDD.n585 0.037532
R10783 VDD VDD.n291 0.0371045
R10784 VDD VDD.n291 0.0371045
R10785 VDD VDD.n582 0.0322201
R10786 VDD.n587 VDD.n586 0.0284258
R10787 VDD.n462 VDD.n285 0.0284
R10788 VDD.n116 VDD.n101 0.026687
R10789 VDD.n282 VDD.n281 0.0255787
R10790 VDD.n582 VDD.n579 0.0253904
R10791 VDD.n384 VDD.n383 0.0239607
R10792 VDD.n384 VDD 0.0239607
R10793 VDD VDD.n302 0.0239607
R10794 VDD.n403 VDD.n302 0.0239607
R10795 VDD.n434 VDD.n404 0.0239607
R10796 VDD.n434 VDD 0.0239607
R10797 VDD VDD.n287 0.0239607
R10798 VDD.n455 VDD.n287 0.0239607
R10799 VDD.n363 VDD 0.0216765
R10800 VDD.n479 VDD.n471 0.0169185
R10801 VDD.n470 VDD.n279 0.0169185
R10802 VDD.n478 VDD.n473 0.0169185
R10803 VDD.n472 VDD.n278 0.0169185
R10804 VDD.n477 VDD.n475 0.0169185
R10805 VDD.n474 VDD.n277 0.0169185
R10806 VDD.n816 VDD.n814 0.0169185
R10807 VDD.n815 VDD.n276 0.0169185
R10808 VDD.n818 VDD.n273 0.0169185
R10809 VDD.n828 VDD.n819 0.0169185
R10810 VDD.n828 VDD.n827 0.0169185
R10811 VDD.n863 VDD.n830 0.0169185
R10812 VDD.n830 VDD.n829 0.0169185
R10813 VDD.n864 VDD.n832 0.0169185
R10814 VDD.n832 VDD.n831 0.0169185
R10815 VDD.n865 VDD.n834 0.0169185
R10816 VDD.n834 VDD.n833 0.0169185
R10817 VDD.n868 VDD.n867 0.0169185
R10818 VDD.n479 VDD.n468 0.0169185
R10819 VDD.n471 VDD.n470 0.0169185
R10820 VDD.n478 VDD.n279 0.0169185
R10821 VDD.n473 VDD.n472 0.0169185
R10822 VDD.n477 VDD.n278 0.0169185
R10823 VDD.n475 VDD.n474 0.0169185
R10824 VDD.n814 VDD.n277 0.0169185
R10825 VDD.n816 VDD.n815 0.0169185
R10826 VDD.n276 VDD.n273 0.0169185
R10827 VDD.n870 VDD.n819 0.0169185
R10828 VDD.n827 VDD.n825 0.0169185
R10829 VDD.n863 VDD.n825 0.0169185
R10830 VDD.n829 VDD.n824 0.0169185
R10831 VDD.n864 VDD.n824 0.0169185
R10832 VDD.n831 VDD.n823 0.0169185
R10833 VDD.n865 VDD.n823 0.0169185
R10834 VDD.n833 VDD.n822 0.0169185
R10835 VDD.n867 VDD.n822 0.0169185
R10836 VDD.n591 VDD.n589 0.0168912
R10837 VDD.n647 VDD.n557 0.0166877
R10838 VDD.n460 VDD.n459 0.0149069
R10839 VDD.n465 VDD.n283 0.0149069
R10840 VDD.n466 VDD.n465 0.0149069
R10841 VDD.n460 VDD.n285 0.0149069
R10842 VDD.n463 VDD.n283 0.0149069
R10843 VDD.n467 VDD.n466 0.0149069
R10844 VDD.n282 VDD.n280 0.0135045
R10845 VDD.n461 VDD.n458 0.0135045
R10846 VDD.n464 VDD.n280 0.0135045
R10847 VDD.n458 VDD.n457 0.0135045
R10848 VDD.n457 VDD.n456 0.0135045
R10849 VDD.n585 VDD.n579 0.0126417
R10850 VDD.n116 VDD.n115 0.00962857
R10851 VDD.n115 VDD.n103 0.00962857
R10852 VDD.n111 VDD.n103 0.00962857
R10853 VDD.n111 VDD.n107 0.00962857
R10854 VDD.n107 VDD.n106 0.00962857
R10855 VDD.n106 VDD.n38 0.00962857
R10856 VDD.n133 VDD.n38 0.00962857
R10857 VDD.n133 VDD.n36 0.00962857
R10858 VDD.n137 VDD.n36 0.00962857
R10859 VDD.n137 VDD.n34 0.00962857
R10860 VDD.n141 VDD.n34 0.00962857
R10861 VDD.n141 VDD.n32 0.00962857
R10862 VDD.n145 VDD.n32 0.00962857
R10863 VDD.n145 VDD.n30 0.00962857
R10864 VDD.n149 VDD.n30 0.00962857
R10865 VDD.n149 VDD.n28 0.00962857
R10866 VDD.n153 VDD.n28 0.00962857
R10867 VDD.n153 VDD.n26 0.00962857
R10868 VDD.n157 VDD.n26 0.00962857
R10869 VDD.n157 VDD.n24 0.00962857
R10870 VDD.n161 VDD.n24 0.00962857
R10871 VDD.n161 VDD.n22 0.00962857
R10872 VDD.n165 VDD.n22 0.00962857
R10873 VDD.n165 VDD.n20 0.00962857
R10874 VDD.n169 VDD.n20 0.00962857
R10875 VDD.n169 VDD.n18 0.00962857
R10876 VDD.n173 VDD.n18 0.00962857
R10877 VDD.n173 VDD.n15 0.00962857
R10878 VDD.n192 VDD.n15 0.00962857
R10879 VDD.n192 VDD.n16 0.00962857
R10880 VDD.n188 VDD.n16 0.00962857
R10881 VDD.n188 VDD.n177 0.00962857
R10882 VDD.n184 VDD.n177 0.00962857
R10883 VDD.n184 VDD.n179 0.00962857
R10884 VDD.n180 VDD.n179 0.00962857
R10885 VDD.n180 VDD.n11 0.00962857
R10886 VDD.n238 VDD.n11 0.00962857
R10887 VDD.n238 VDD.n9 0.00962857
R10888 VDD.n242 VDD.n9 0.00962857
R10889 VDD.n242 VDD.n7 0.00962857
R10890 VDD.n246 VDD.n7 0.00962857
R10891 VDD.n246 VDD.n4 0.00962857
R10892 VDD.n923 VDD.n4 0.00962857
R10893 VDD.n923 VDD.n5 0.00962857
R10894 VDD.n919 VDD.n5 0.00962857
R10895 VDD.n919 VDD.n250 0.00962857
R10896 VDD.n915 VDD.n250 0.00962857
R10897 VDD.n915 VDD.n252 0.00962857
R10898 VDD.n911 VDD.n252 0.00962857
R10899 VDD.n911 VDD.n254 0.00962857
R10900 VDD.n907 VDD.n254 0.00962857
R10901 VDD.n907 VDD.n256 0.00962857
R10902 VDD.n903 VDD.n256 0.00962857
R10903 VDD.n903 VDD.n258 0.00962857
R10904 VDD.n899 VDD.n258 0.00962857
R10905 VDD.n899 VDD.n260 0.00962857
R10906 VDD.n895 VDD.n260 0.00962857
R10907 VDD.n895 VDD.n262 0.00962857
R10908 VDD.n891 VDD.n262 0.00962857
R10909 VDD.n891 VDD.n264 0.00962857
R10910 VDD.n887 VDD.n264 0.00962857
R10911 VDD.n887 VDD.n266 0.00962857
R10912 VDD.n883 VDD.n266 0.00962857
R10913 VDD.n883 VDD.n268 0.00962857
R10914 VDD.n879 VDD.n268 0.00962857
R10915 VDD.n879 VDD.n270 0.00962857
R10916 VDD.n842 VDD.n270 0.00962857
R10917 VDD.n845 VDD.n842 0.00962857
R10918 VDD.n845 VDD.n840 0.00962857
R10919 VDD.n849 VDD.n840 0.00962857
R10920 VDD.n849 VDD.n838 0.00962857
R10921 VDD.n853 VDD.n838 0.00962857
R10922 VDD.n857 VDD.n856 0.00962857
R10923 VDD.n857 VDD.n835 0.00962857
R10924 VDD.n861 VDD.n835 0.00962857
R10925 VDD.n647 VDD.n646 0.00962857
R10926 VDD.n646 VDD.n559 0.00962857
R10927 VDD.n642 VDD.n559 0.00962857
R10928 VDD.n642 VDD.n561 0.00962857
R10929 VDD.n638 VDD.n561 0.00962857
R10930 VDD.n638 VDD.n564 0.00962857
R10931 VDD.n634 VDD.n564 0.00962857
R10932 VDD.n634 VDD.n566 0.00962857
R10933 VDD.n630 VDD.n566 0.00962857
R10934 VDD.n630 VDD.n568 0.00962857
R10935 VDD.n626 VDD.n568 0.00962857
R10936 VDD.n626 VDD.n570 0.00962857
R10937 VDD.n622 VDD.n570 0.00962857
R10938 VDD.n622 VDD.n572 0.00962857
R10939 VDD.n618 VDD.n572 0.00962857
R10940 VDD.n618 VDD.n574 0.00962857
R10941 VDD.n613 VDD.n574 0.00962857
R10942 VDD.n613 VDD.n600 0.00962857
R10943 VDD.n609 VDD.n600 0.00962857
R10944 VDD.n609 VDD.n602 0.00962857
R10945 VDD.n605 VDD.n602 0.00962857
R10946 VDD.n605 VDD.n554 0.00962857
R10947 VDD.n665 VDD.n554 0.00962857
R10948 VDD.n665 VDD.n552 0.00962857
R10949 VDD.n669 VDD.n552 0.00962857
R10950 VDD.n669 VDD.n550 0.00962857
R10951 VDD.n673 VDD.n550 0.00962857
R10952 VDD.n673 VDD.n548 0.00962857
R10953 VDD.n677 VDD.n548 0.00962857
R10954 VDD.n677 VDD.n546 0.00962857
R10955 VDD.n681 VDD.n546 0.00962857
R10956 VDD.n681 VDD.n544 0.00962857
R10957 VDD.n685 VDD.n544 0.00962857
R10958 VDD.n685 VDD.n542 0.00962857
R10959 VDD.n689 VDD.n542 0.00962857
R10960 VDD.n689 VDD.n540 0.00962857
R10961 VDD.n693 VDD.n540 0.00962857
R10962 VDD.n693 VDD.n538 0.00962857
R10963 VDD.n697 VDD.n538 0.00962857
R10964 VDD.n697 VDD.n536 0.00962857
R10965 VDD.n701 VDD.n536 0.00962857
R10966 VDD.n701 VDD.n534 0.00962857
R10967 VDD.n705 VDD.n534 0.00962857
R10968 VDD.n705 VDD.n532 0.00962857
R10969 VDD.n709 VDD.n532 0.00962857
R10970 VDD.n709 VDD.n530 0.00962857
R10971 VDD.n713 VDD.n530 0.00962857
R10972 VDD.n713 VDD.n528 0.00962857
R10973 VDD.n717 VDD.n528 0.00962857
R10974 VDD.n717 VDD.n526 0.00962857
R10975 VDD.n721 VDD.n526 0.00962857
R10976 VDD.n721 VDD.n524 0.00962857
R10977 VDD.n725 VDD.n524 0.00962857
R10978 VDD.n725 VDD.n522 0.00962857
R10979 VDD.n729 VDD.n522 0.00962857
R10980 VDD.n729 VDD.n520 0.00962857
R10981 VDD.n733 VDD.n520 0.00962857
R10982 VDD.n733 VDD.n518 0.00962857
R10983 VDD.n737 VDD.n518 0.00962857
R10984 VDD.n737 VDD.n516 0.00962857
R10985 VDD.n741 VDD.n516 0.00962857
R10986 VDD.n741 VDD.n514 0.00962857
R10987 VDD.n745 VDD.n514 0.00962857
R10988 VDD.n745 VDD.n512 0.00962857
R10989 VDD.n749 VDD.n512 0.00962857
R10990 VDD.n749 VDD.n510 0.00962857
R10991 VDD.n753 VDD.n510 0.00962857
R10992 VDD.n753 VDD.n508 0.00962857
R10993 VDD.n757 VDD.n508 0.00962857
R10994 VDD.n757 VDD.n506 0.00962857
R10995 VDD.n761 VDD.n506 0.00962857
R10996 VDD.n761 VDD.n504 0.00962857
R10997 VDD.n765 VDD.n504 0.00962857
R10998 VDD.n765 VDD.n502 0.00962857
R10999 VDD.n769 VDD.n502 0.00962857
R11000 VDD.n769 VDD.n500 0.00962857
R11001 VDD.n773 VDD.n500 0.00962857
R11002 VDD.n773 VDD.n498 0.00962857
R11003 VDD.n777 VDD.n498 0.00962857
R11004 VDD.n777 VDD.n496 0.00962857
R11005 VDD.n781 VDD.n496 0.00962857
R11006 VDD.n781 VDD.n494 0.00962857
R11007 VDD.n785 VDD.n494 0.00962857
R11008 VDD.n785 VDD.n492 0.00962857
R11009 VDD.n789 VDD.n492 0.00962857
R11010 VDD.n789 VDD.n490 0.00962857
R11011 VDD.n793 VDD.n490 0.00962857
R11012 VDD.n793 VDD.n488 0.00962857
R11013 VDD.n797 VDD.n488 0.00962857
R11014 VDD.n797 VDD.n486 0.00962857
R11015 VDD.n801 VDD.n486 0.00962857
R11016 VDD.n801 VDD.n484 0.00962857
R11017 VDD.n805 VDD.n484 0.00962857
R11018 VDD.n809 VDD.n808 0.00962857
R11019 VDD.n810 VDD.n809 0.00962857
R11020 VDD.n810 VDD.n480 0.00962857
R11021 VDD.n648 VDD.n558 0.00962857
R11022 VDD.n562 VDD.n558 0.00962857
R11023 VDD.n641 VDD.n562 0.00962857
R11024 VDD.n641 VDD.n640 0.00962857
R11025 VDD.n640 VDD.n639 0.00962857
R11026 VDD.n639 VDD.n563 0.00962857
R11027 VDD.n633 VDD.n563 0.00962857
R11028 VDD.n633 VDD.n632 0.00962857
R11029 VDD.n632 VDD.n631 0.00962857
R11030 VDD.n631 VDD.n567 0.00962857
R11031 VDD.n625 VDD.n567 0.00962857
R11032 VDD.n625 VDD.n624 0.00962857
R11033 VDD.n624 VDD.n623 0.00962857
R11034 VDD.n623 VDD.n571 0.00962857
R11035 VDD.n617 VDD.n571 0.00962857
R11036 VDD.n617 VDD.n616 0.00962857
R11037 VDD.n608 VDD.n603 0.00962857
R11038 VDD.n608 VDD.n607 0.00962857
R11039 VDD.n607 VDD.n606 0.00962857
R11040 VDD.n606 VDD.n555 0.00962857
R11041 VDD.n664 VDD.n551 0.00962857
R11042 VDD.n670 VDD.n551 0.00962857
R11043 VDD.n671 VDD.n670 0.00962857
R11044 VDD.n672 VDD.n671 0.00962857
R11045 VDD.n672 VDD.n547 0.00962857
R11046 VDD.n678 VDD.n547 0.00962857
R11047 VDD.n679 VDD.n678 0.00962857
R11048 VDD.n680 VDD.n679 0.00962857
R11049 VDD.n680 VDD.n543 0.00962857
R11050 VDD.n686 VDD.n543 0.00962857
R11051 VDD.n687 VDD.n686 0.00962857
R11052 VDD.n688 VDD.n687 0.00962857
R11053 VDD.n688 VDD.n539 0.00962857
R11054 VDD.n694 VDD.n539 0.00962857
R11055 VDD.n695 VDD.n694 0.00962857
R11056 VDD.n696 VDD.n695 0.00962857
R11057 VDD.n696 VDD.n535 0.00962857
R11058 VDD.n702 VDD.n535 0.00962857
R11059 VDD.n703 VDD.n702 0.00962857
R11060 VDD.n704 VDD.n703 0.00962857
R11061 VDD.n704 VDD.n531 0.00962857
R11062 VDD.n710 VDD.n531 0.00962857
R11063 VDD.n711 VDD.n710 0.00962857
R11064 VDD.n712 VDD.n711 0.00962857
R11065 VDD.n712 VDD.n527 0.00962857
R11066 VDD.n718 VDD.n527 0.00962857
R11067 VDD.n719 VDD.n718 0.00962857
R11068 VDD.n720 VDD.n719 0.00962857
R11069 VDD.n720 VDD.n523 0.00962857
R11070 VDD.n726 VDD.n523 0.00962857
R11071 VDD.n727 VDD.n726 0.00962857
R11072 VDD.n728 VDD.n727 0.00962857
R11073 VDD.n728 VDD.n519 0.00962857
R11074 VDD.n734 VDD.n519 0.00962857
R11075 VDD.n735 VDD.n734 0.00962857
R11076 VDD.n736 VDD.n735 0.00962857
R11077 VDD.n736 VDD.n515 0.00962857
R11078 VDD.n742 VDD.n515 0.00962857
R11079 VDD.n743 VDD.n742 0.00962857
R11080 VDD.n744 VDD.n743 0.00962857
R11081 VDD.n744 VDD.n511 0.00962857
R11082 VDD.n750 VDD.n511 0.00962857
R11083 VDD.n751 VDD.n750 0.00962857
R11084 VDD.n752 VDD.n751 0.00962857
R11085 VDD.n752 VDD.n507 0.00962857
R11086 VDD.n758 VDD.n507 0.00962857
R11087 VDD.n759 VDD.n758 0.00962857
R11088 VDD.n760 VDD.n759 0.00962857
R11089 VDD.n760 VDD.n503 0.00962857
R11090 VDD.n766 VDD.n503 0.00962857
R11091 VDD.n767 VDD.n766 0.00962857
R11092 VDD.n768 VDD.n767 0.00962857
R11093 VDD.n768 VDD.n499 0.00962857
R11094 VDD.n774 VDD.n499 0.00962857
R11095 VDD.n775 VDD.n774 0.00962857
R11096 VDD.n776 VDD.n775 0.00962857
R11097 VDD.n776 VDD.n495 0.00962857
R11098 VDD.n782 VDD.n495 0.00962857
R11099 VDD.n783 VDD.n782 0.00962857
R11100 VDD.n784 VDD.n783 0.00962857
R11101 VDD.n784 VDD.n491 0.00962857
R11102 VDD.n790 VDD.n491 0.00962857
R11103 VDD.n791 VDD.n790 0.00962857
R11104 VDD.n792 VDD.n791 0.00962857
R11105 VDD.n792 VDD.n487 0.00962857
R11106 VDD.n798 VDD.n487 0.00962857
R11107 VDD.n799 VDD.n798 0.00962857
R11108 VDD.n800 VDD.n799 0.00962857
R11109 VDD.n800 VDD.n483 0.00962857
R11110 VDD.n806 VDD.n483 0.00962857
R11111 VDD.n807 VDD.n275 0.00962857
R11112 VDD.n117 VDD.n102 0.00962857
R11113 VDD.n108 VDD.n102 0.00962857
R11114 VDD.n110 VDD.n108 0.00962857
R11115 VDD.n110 VDD.n109 0.00962857
R11116 VDD.n109 VDD.n39 0.00962857
R11117 VDD.n132 VDD.n131 0.00962857
R11118 VDD.n132 VDD.n35 0.00962857
R11119 VDD.n138 VDD.n35 0.00962857
R11120 VDD.n139 VDD.n138 0.00962857
R11121 VDD.n140 VDD.n139 0.00962857
R11122 VDD.n140 VDD.n31 0.00962857
R11123 VDD.n146 VDD.n31 0.00962857
R11124 VDD.n147 VDD.n146 0.00962857
R11125 VDD.n148 VDD.n147 0.00962857
R11126 VDD.n148 VDD.n27 0.00962857
R11127 VDD.n154 VDD.n27 0.00962857
R11128 VDD.n155 VDD.n154 0.00962857
R11129 VDD.n156 VDD.n155 0.00962857
R11130 VDD.n156 VDD.n23 0.00962857
R11131 VDD.n162 VDD.n23 0.00962857
R11132 VDD.n163 VDD.n162 0.00962857
R11133 VDD.n164 VDD.n163 0.00962857
R11134 VDD.n164 VDD.n19 0.00962857
R11135 VDD.n170 VDD.n19 0.00962857
R11136 VDD.n171 VDD.n170 0.00962857
R11137 VDD.n172 VDD.n171 0.00962857
R11138 VDD.n172 VDD.n13 0.00962857
R11139 VDD.n193 VDD.n14 0.00962857
R11140 VDD.n187 VDD.n14 0.00962857
R11141 VDD.n187 VDD.n186 0.00962857
R11142 VDD.n186 VDD.n185 0.00962857
R11143 VDD.n185 VDD.n178 0.00962857
R11144 VDD.n178 VDD.n12 0.00962857
R11145 VDD.n237 VDD.n236 0.00962857
R11146 VDD.n237 VDD.n8 0.00962857
R11147 VDD.n243 VDD.n8 0.00962857
R11148 VDD.n244 VDD.n243 0.00962857
R11149 VDD.n245 VDD.n244 0.00962857
R11150 VDD.n245 VDD.n2 0.00962857
R11151 VDD.n924 VDD.n3 0.00962857
R11152 VDD.n918 VDD.n3 0.00962857
R11153 VDD.n918 VDD.n917 0.00962857
R11154 VDD.n917 VDD.n916 0.00962857
R11155 VDD.n916 VDD.n251 0.00962857
R11156 VDD.n910 VDD.n251 0.00962857
R11157 VDD.n910 VDD.n909 0.00962857
R11158 VDD.n909 VDD.n908 0.00962857
R11159 VDD.n908 VDD.n255 0.00962857
R11160 VDD.n902 VDD.n255 0.00962857
R11161 VDD.n902 VDD.n901 0.00962857
R11162 VDD.n901 VDD.n900 0.00962857
R11163 VDD.n900 VDD.n259 0.00962857
R11164 VDD.n894 VDD.n259 0.00962857
R11165 VDD.n894 VDD.n893 0.00962857
R11166 VDD.n893 VDD.n892 0.00962857
R11167 VDD.n892 VDD.n263 0.00962857
R11168 VDD.n886 VDD.n263 0.00962857
R11169 VDD.n886 VDD.n885 0.00962857
R11170 VDD.n885 VDD.n884 0.00962857
R11171 VDD.n884 VDD.n267 0.00962857
R11172 VDD.n878 VDD.n267 0.00962857
R11173 VDD.n841 VDD.n271 0.00962857
R11174 VDD.n846 VDD.n841 0.00962857
R11175 VDD.n847 VDD.n846 0.00962857
R11176 VDD.n848 VDD.n847 0.00962857
R11177 VDD.n848 VDD.n837 0.00962857
R11178 VDD.n854 VDD.n837 0.00962857
R11179 VDD.n855 VDD.n821 0.00962857
R11180 VDD.n616 VDD.n615 0.00956429
R11181 VDD.n594 VDD.n593 0.00915093
R11182 VDD.n588 VDD.n587 0.00884739
R11183 VDD.n194 VDD.n13 0.0086
R11184 VDD.n649 VDD.n648 0.00853571
R11185 VDD.n817 VDD.n275 0.00827857
R11186 VDD.n469 VDD.n274 0.00827857
R11187 VDD.n813 VDD.n476 0.00827857
R11188 VDD.n869 VDD.n821 0.00827857
R11189 VDD.n866 VDD.n826 0.00827857
R11190 VDD.n862 VDD.n820 0.00827857
R11191 VDD.n878 VDD.n877 0.00795714
R11192 VDD.n853 VDD 0.00782857
R11193 VDD.n805 VDD 0.00782857
R11194 VDD VDD.n806 0.00782857
R11195 VDD VDD.n854 0.00782857
R11196 VDD.n614 VDD.n599 0.00763571
R11197 VDD.n663 VDD.n555 0.00692857
R11198 VDD.n235 VDD.n12 0.0068
R11199 VDD.n114 VDD.n113 0.00658571
R11200 VDD.n113 VDD.n112 0.00658571
R11201 VDD.n112 VDD.n104 0.00658571
R11202 VDD.n105 VDD.n104 0.00658571
R11203 VDD.n105 VDD.n37 0.00658571
R11204 VDD.n134 VDD.n37 0.00658571
R11205 VDD.n135 VDD.n134 0.00658571
R11206 VDD.n136 VDD.n135 0.00658571
R11207 VDD.n136 VDD.n33 0.00658571
R11208 VDD.n142 VDD.n33 0.00658571
R11209 VDD.n143 VDD.n142 0.00658571
R11210 VDD.n144 VDD.n143 0.00658571
R11211 VDD.n144 VDD.n29 0.00658571
R11212 VDD.n150 VDD.n29 0.00658571
R11213 VDD.n151 VDD.n150 0.00658571
R11214 VDD.n152 VDD.n151 0.00658571
R11215 VDD.n152 VDD.n25 0.00658571
R11216 VDD.n158 VDD.n25 0.00658571
R11217 VDD.n159 VDD.n158 0.00658571
R11218 VDD.n160 VDD.n159 0.00658571
R11219 VDD.n160 VDD.n21 0.00658571
R11220 VDD.n166 VDD.n21 0.00658571
R11221 VDD.n167 VDD.n166 0.00658571
R11222 VDD.n168 VDD.n167 0.00658571
R11223 VDD.n168 VDD.n17 0.00658571
R11224 VDD.n174 VDD.n17 0.00658571
R11225 VDD.n175 VDD.n174 0.00658571
R11226 VDD.n191 VDD.n175 0.00658571
R11227 VDD.n191 VDD.n190 0.00658571
R11228 VDD.n190 VDD.n189 0.00658571
R11229 VDD.n189 VDD.n176 0.00658571
R11230 VDD.n183 VDD.n176 0.00658571
R11231 VDD.n183 VDD.n182 0.00658571
R11232 VDD.n182 VDD.n181 0.00658571
R11233 VDD.n181 VDD.n10 0.00658571
R11234 VDD.n239 VDD.n10 0.00658571
R11235 VDD.n240 VDD.n239 0.00658571
R11236 VDD.n241 VDD.n240 0.00658571
R11237 VDD.n241 VDD.n6 0.00658571
R11238 VDD.n247 VDD.n6 0.00658571
R11239 VDD.n248 VDD.n247 0.00658571
R11240 VDD.n922 VDD.n248 0.00658571
R11241 VDD.n922 VDD.n921 0.00658571
R11242 VDD.n921 VDD.n920 0.00658571
R11243 VDD.n920 VDD.n249 0.00658571
R11244 VDD.n914 VDD.n249 0.00658571
R11245 VDD.n914 VDD.n913 0.00658571
R11246 VDD.n913 VDD.n912 0.00658571
R11247 VDD.n912 VDD.n253 0.00658571
R11248 VDD.n906 VDD.n253 0.00658571
R11249 VDD.n906 VDD.n905 0.00658571
R11250 VDD.n905 VDD.n904 0.00658571
R11251 VDD.n904 VDD.n257 0.00658571
R11252 VDD.n898 VDD.n257 0.00658571
R11253 VDD.n898 VDD.n897 0.00658571
R11254 VDD.n897 VDD.n896 0.00658571
R11255 VDD.n896 VDD.n261 0.00658571
R11256 VDD.n890 VDD.n261 0.00658571
R11257 VDD.n890 VDD.n889 0.00658571
R11258 VDD.n889 VDD.n888 0.00658571
R11259 VDD.n888 VDD.n265 0.00658571
R11260 VDD.n882 VDD.n265 0.00658571
R11261 VDD.n882 VDD.n881 0.00658571
R11262 VDD.n881 VDD.n880 0.00658571
R11263 VDD.n880 VDD.n269 0.00658571
R11264 VDD.n843 VDD.n269 0.00658571
R11265 VDD.n844 VDD.n843 0.00658571
R11266 VDD.n844 VDD.n839 0.00658571
R11267 VDD.n850 VDD.n839 0.00658571
R11268 VDD.n851 VDD.n850 0.00658571
R11269 VDD.n852 VDD.n851 0.00658571
R11270 VDD.n852 VDD.n836 0.00658571
R11271 VDD.n859 VDD.n858 0.00658571
R11272 VDD.n645 VDD.n644 0.00658571
R11273 VDD.n644 VDD.n643 0.00658571
R11274 VDD.n643 VDD.n560 0.00658571
R11275 VDD.n637 VDD.n560 0.00658571
R11276 VDD.n637 VDD.n636 0.00658571
R11277 VDD.n636 VDD.n635 0.00658571
R11278 VDD.n635 VDD.n565 0.00658571
R11279 VDD.n629 VDD.n565 0.00658571
R11280 VDD.n629 VDD.n628 0.00658571
R11281 VDD.n628 VDD.n627 0.00658571
R11282 VDD.n627 VDD.n569 0.00658571
R11283 VDD.n621 VDD.n569 0.00658571
R11284 VDD.n621 VDD.n620 0.00658571
R11285 VDD.n620 VDD.n619 0.00658571
R11286 VDD.n619 VDD.n573 0.00658571
R11287 VDD.n612 VDD.n573 0.00658571
R11288 VDD.n612 VDD.n611 0.00658571
R11289 VDD.n611 VDD.n610 0.00658571
R11290 VDD.n610 VDD.n601 0.00658571
R11291 VDD.n604 VDD.n601 0.00658571
R11292 VDD.n604 VDD.n553 0.00658571
R11293 VDD.n666 VDD.n553 0.00658571
R11294 VDD.n667 VDD.n666 0.00658571
R11295 VDD.n668 VDD.n667 0.00658571
R11296 VDD.n668 VDD.n549 0.00658571
R11297 VDD.n674 VDD.n549 0.00658571
R11298 VDD.n675 VDD.n674 0.00658571
R11299 VDD.n676 VDD.n675 0.00658571
R11300 VDD.n676 VDD.n545 0.00658571
R11301 VDD.n682 VDD.n545 0.00658571
R11302 VDD.n683 VDD.n682 0.00658571
R11303 VDD.n684 VDD.n683 0.00658571
R11304 VDD.n684 VDD.n541 0.00658571
R11305 VDD.n690 VDD.n541 0.00658571
R11306 VDD.n691 VDD.n690 0.00658571
R11307 VDD.n692 VDD.n691 0.00658571
R11308 VDD.n692 VDD.n537 0.00658571
R11309 VDD.n698 VDD.n537 0.00658571
R11310 VDD.n699 VDD.n698 0.00658571
R11311 VDD.n700 VDD.n699 0.00658571
R11312 VDD.n700 VDD.n533 0.00658571
R11313 VDD.n706 VDD.n533 0.00658571
R11314 VDD.n707 VDD.n706 0.00658571
R11315 VDD.n708 VDD.n707 0.00658571
R11316 VDD.n708 VDD.n529 0.00658571
R11317 VDD.n714 VDD.n529 0.00658571
R11318 VDD.n715 VDD.n714 0.00658571
R11319 VDD.n716 VDD.n715 0.00658571
R11320 VDD.n716 VDD.n525 0.00658571
R11321 VDD.n722 VDD.n525 0.00658571
R11322 VDD.n723 VDD.n722 0.00658571
R11323 VDD.n724 VDD.n723 0.00658571
R11324 VDD.n724 VDD.n521 0.00658571
R11325 VDD.n730 VDD.n521 0.00658571
R11326 VDD.n731 VDD.n730 0.00658571
R11327 VDD.n732 VDD.n731 0.00658571
R11328 VDD.n732 VDD.n517 0.00658571
R11329 VDD.n738 VDD.n517 0.00658571
R11330 VDD.n739 VDD.n738 0.00658571
R11331 VDD.n740 VDD.n739 0.00658571
R11332 VDD.n740 VDD.n513 0.00658571
R11333 VDD.n746 VDD.n513 0.00658571
R11334 VDD.n747 VDD.n746 0.00658571
R11335 VDD.n748 VDD.n747 0.00658571
R11336 VDD.n748 VDD.n509 0.00658571
R11337 VDD.n754 VDD.n509 0.00658571
R11338 VDD.n755 VDD.n754 0.00658571
R11339 VDD.n756 VDD.n755 0.00658571
R11340 VDD.n756 VDD.n505 0.00658571
R11341 VDD.n762 VDD.n505 0.00658571
R11342 VDD.n763 VDD.n762 0.00658571
R11343 VDD.n764 VDD.n763 0.00658571
R11344 VDD.n764 VDD.n501 0.00658571
R11345 VDD.n770 VDD.n501 0.00658571
R11346 VDD.n771 VDD.n770 0.00658571
R11347 VDD.n772 VDD.n771 0.00658571
R11348 VDD.n772 VDD.n497 0.00658571
R11349 VDD.n778 VDD.n497 0.00658571
R11350 VDD.n779 VDD.n778 0.00658571
R11351 VDD.n780 VDD.n779 0.00658571
R11352 VDD.n780 VDD.n493 0.00658571
R11353 VDD.n786 VDD.n493 0.00658571
R11354 VDD.n787 VDD.n786 0.00658571
R11355 VDD.n788 VDD.n787 0.00658571
R11356 VDD.n788 VDD.n489 0.00658571
R11357 VDD.n794 VDD.n489 0.00658571
R11358 VDD.n795 VDD.n794 0.00658571
R11359 VDD.n796 VDD.n795 0.00658571
R11360 VDD.n796 VDD.n485 0.00658571
R11361 VDD.n802 VDD.n485 0.00658571
R11362 VDD.n803 VDD.n802 0.00658571
R11363 VDD.n804 VDD.n803 0.00658571
R11364 VDD.n811 VDD.n481 0.00658571
R11365 VDD.n335 VDD 0.00654478
R11366 VDD.n309 VDD 0.00654478
R11367 VDD.n351 VDD 0.00642105
R11368 VDD.n378 VDD 0.00642105
R11369 VDD.n657 VDD 0.00642105
R11370 VDD.n591 VDD.n590 0.00641906
R11371 VDD.n590 VDD.n576 0.00641906
R11372 VDD.n858 VDD 0.00641429
R11373 VDD VDD.n481 0.00641429
R11374 VDD.n118 VDD.n117 0.00583571
R11375 VDD.n130 VDD.n39 0.00564286
R11376 VDD.n861 VDD.n860 0.00548841
R11377 VDD.n812 VDD.n480 0.00548841
R11378 VDD.n804 VDD 0.00538571
R11379 VDD.n925 VDD.n924 0.00512857
R11380 VDD.n583 VDD 0.00505312
R11381 VDD VDD.n588 0.00505312
R11382 VDD.n593 VDD.n576 0.00505312
R11383 VDD.n925 VDD.n2 0.005
R11384 VDD.n131 VDD.n130 0.00448571
R11385 VDD.n589 VDD 0.00399073
R11386 VDD.n236 VDD.n235 0.00332857
R11387 VDD.n664 VDD.n663 0.0032
R11388 VDD.n382 VDD.n342 0.00286842
R11389 VDD.n603 VDD.n599 0.00249286
R11390 VDD.n856 VDD 0.0023
R11391 VDD.n808 VDD 0.0023
R11392 VDD.n807 VDD 0.0023
R11393 VDD.n855 VDD 0.0023
R11394 VDD.n877 VDD.n271 0.00217143
R11395 VDD VDD.n228 0.002
R11396 VDD.n817 VDD.n469 0.00185
R11397 VDD.n476 VDD.n274 0.00185
R11398 VDD.n869 VDD.n826 0.00185
R11399 VDD.n866 VDD.n862 0.00185
R11400 VDD VDD.n482 0.0017
R11401 VDD.n194 VDD.n193 0.00152857
R11402 VDD.n836 VDD 0.000671429
R11403 VDD.n482 VDD 0.000671429
R11404 VDD.n615 VDD.n614 0.000564286
R11405 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t9 82.0028
R11406 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t5 82.0028
R11407 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t8 82.0028
R11408 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t3 82.0028
R11409 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t7 42.2319
R11410 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t4 42.2319
R11411 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t6 42.2319
R11412 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t2 42.2319
R11413 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 10.5577
R11414 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 10.4346
R11415 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 6.98616
R11416 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.n0 4.85103
R11417 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.n2 4.69358
R11418 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 4.47707
R11419 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.n1 2.2505
R11420 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t1 2.04837
R11421 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t0 1.49421
R11422 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t6 80.4772
R11423 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t7 80.4772
R11424 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t3 62.5719
R11425 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t8 62.5719
R11426 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t4 45.4098
R11427 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t5 34.4148
R11428 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n1 8.06816
R11429 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n0 8.06816
R11430 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n2 6.31953
R11431 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n4 6.08116
R11432 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n3 4.80357
R11433 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t1 4.54043
R11434 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t2 1.1409
R11435 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 0.702585
R11436 DVSS.n1730 DVSS.n1516 196056
R11437 DVSS.n3592 DVSS.n3591 37210.9
R11438 DVSS.n4944 DVSS.n1169 32551.1
R11439 DVSS.n4488 DVSS.n4487 32385.4
R11440 DVSS.n3590 DVSS.n3589 30893.3
R11441 DVSS.n5353 DVSS.n5352 27088.7
R11442 DVSS.n5112 DVSS.n960 25861.7
R11443 DVSS.n3943 DVSS.n1516 21519.5
R11444 DVSS.n5352 DVSS.n962 20471.6
R11445 DVSS.n3983 DVSS.n1439 19823.1
R11446 DVSS.n5113 DVSS.n5112 19552.7
R11447 DVSS.n1492 DVSS.n1491 17654
R11448 DVSS.n4925 DVSS.n961 16516.8
R11449 DVSS.n4489 DVSS.n1273 16516.8
R11450 DVSS.n1491 DVSS.n1158 16432
R11451 DVSS.n3590 DVSS.n1438 16400
R11452 DVSS.n1863 DVSS.n1862 16252.3
R11453 DVSS.n5353 DVSS.n961 16242.7
R11454 DVSS.n1273 DVSS.n960 16242.7
R11455 DVSS.n4953 DVSS.n1166 16230.9
R11456 DVSS.n4968 DVSS.n1158 16230.9
R11457 DVSS.n1491 DVSS.n1490 16230.9
R11458 DVSS.n1492 DVSS.n1481 16230.9
R11459 DVSS.n4467 DVSS.n1286 16230.9
R11460 DVSS.n3589 DVSS.n2235 15030.2
R11461 DVSS.n2253 DVSS.n2235 14984.7
R11462 DVSS.n3985 DVSS.n3983 14824
R11463 DVSS.n1863 DVSS.n1438 14824
R11464 DVSS.n5354 DVSS.n5353 14769.2
R11465 DVSS.n5355 DVSS.n960 14767.1
R11466 DVSS.n3592 DVSS.n3590 13915.8
R11467 DVSS.n2660 DVSS.n2263 12369.1
R11468 DVSS.n3558 DVSS.n2238 12369.1
R11469 DVSS.n3567 DVSS.n3559 12369.1
R11470 DVSS.n3760 DVSS.n1694 12369.1
R11471 DVSS.n3985 DVSS.n3984 11473.2
R11472 DVSS.n3984 DVSS.n1166 10835.5
R11473 DVSS.n3591 DVSS.n1167 10290.4
R11474 DVSS.n3591 DVSS.n1166 8547.5
R11475 DVSS.n3589 DVSS.n3588 7940.47
R11476 DVSS.n4487 DVSS.n1274 7811.82
R11477 DVSS.n3943 DVSS.n3942 7328.63
R11478 DVSS.n3648 DVSS.n3647 6939.76
R11479 DVSS.n1862 DVSS.n1861 6651.3
R11480 DVSS.n3976 DVSS.n1493 6538.35
R11481 DVSS.n3559 DVSS.n3558 6519.88
R11482 DVSS.n2658 DVSS.n1694 6104.43
R11483 DVSS.n3645 DVSS.n3592 5387.7
R11484 DVSS.n4967 DVSS.n1159 4902.86
R11485 DVSS.n4954 DVSS.n1165 4902.86
R11486 DVSS.n1482 DVSS.n1304 4902.86
R11487 DVSS.n1493 DVSS.n1286 4526.71
R11488 DVSS.n2254 DVSS.n2253 4493.06
R11489 DVSS.n1862 DVSS.n1516 3491.91
R11490 DVSS.n3986 DVSS.n3985 3437.85
R11491 DVSS.n3986 DVSS.n1438 3435.27
R11492 DVSS.n1922 DVSS.t19 3354.59
R11493 DVSS.n2161 DVSS.t19 3354.59
R11494 DVSS.n1493 DVSS.n1492 3311.99
R11495 DVSS.n3944 DVSS.n3943 3307.91
R11496 DVSS.n3559 DVSS.n2254 3136.7
R11497 DVSS.n1861 DVSS.n1439 3086.59
R11498 DVSS.n3750 DVSS.n1694 2581.97
R11499 DVSS.n3942 DVSS.n1517 2507.4
R11500 DVSS.n2657 DVSS.n1024 2402.48
R11501 DVSS.n5231 DVSS.n1024 2401.2
R11502 DVSS.n2657 DVSS.n1023 2400.01
R11503 DVSS.n5231 DVSS.n1023 2398.73
R11504 DVSS.n3558 DVSS.n3557 2395.26
R11505 DVSS.n4924 DVSS.n4923 2286.22
R11506 DVSS.n4677 DVSS.n4676 2282.35
R11507 DVSS.n4677 DVSS.n1216 2282.35
R11508 DVSS.n4676 DVSS.n4675 2278.48
R11509 DVSS.n4923 DVSS.n1216 2277.19
R11510 DVSS.n1511 DVSS.n1286 2219.8
R11511 DVSS.n4926 DVSS.n4924 2185.59
R11512 DVSS.n4675 DVSS.n4490 2179.14
R11513 DVSS.n3984 DVSS.n1158 2099.5
R11514 DVSS.n1862 DVSS.n1494 1819.86
R11515 DVSS.n2235 DVSS.n2234 1783.15
R11516 DVSS.n4946 DVSS.n4945 1674.85
R11517 DVSS.n3557 DVSS.n2660 1508.72
R11518 DVSS.n4384 DVSS.t32 1472.87
R11519 DVSS.n4388 DVSS.t37 1472.87
R11520 DVSS.n1454 DVSS.t40 1472.87
R11521 DVSS.n1456 DVSS.t44 1472.87
R11522 DVSS.n4963 DVSS.n1163 1449.32
R11523 DVSS.n4977 DVSS.n1156 1375
R11524 DVSS.n2234 DVSS.n2233 1219.32
R11525 DVSS.n1489 DVSS.n1157 1124.46
R11526 DVSS.n4977 DVSS.n1157 1124.46
R11527 DVSS.n4977 DVSS.n4976 1124.46
R11528 DVSS.n4976 DVSS.n4969 1124.46
R11529 DVSS.n3749 DVSS.n1700 1105.19
R11530 DVSS.t181 DVSS.n1302 1075.57
R11531 DVSS.n4966 DVSS.t96 1075.57
R11532 DVSS.t194 DVSS.n4955 1075.57
R11533 DVSS.n3751 DVSS.n3750 1047.22
R11534 DVSS.n4946 DVSS.n1167 1041.24
R11535 DVSS.n3648 DVSS.n1700 1024.12
R11536 DVSS.n4490 DVSS.n4489 967.646
R11537 DVSS.n4926 DVSS.n4925 967.646
R11538 DVSS.n3945 DVSS.n3944 835.686
R11539 DVSS.n3750 DVSS.n3749 826.212
R11540 DVSS.t136 DVSS.n4963 824.14
R11541 DVSS.n4963 DVSS.t81 824.14
R11542 DVSS.n4952 DVSS.n1167 796.203
R11543 DVSS.n2230 DVSS.t107 782.032
R11544 DVSS.n2235 DVSS.n1517 724.26
R11545 DVSS.n1490 DVSS.n1489 693.769
R11546 DVSS.n4969 DVSS.n4968 693.769
R11547 DVSS.n4953 DVSS.n4952 693.769
R11548 DVSS.t50 DVSS.t185 640.298
R11549 DVSS.t87 DVSS.t141 640.298
R11550 DVSS.t117 DVSS.t92 640.298
R11551 DVSS.t53 DVSS.t20 640.298
R11552 DVSS.n2233 DVSS.n1730 614.245
R11553 DVSS.n4489 DVSS.n4488 608.972
R11554 DVSS.n4925 DVSS.n1169 608.972
R11555 DVSS.n3622 DVSS.t9 587.904
R11556 DVSS.n2661 DVSS.n1701 586.833
R11557 DVSS.n2253 DVSS.n2252 562.811
R11558 DVSS.n1482 DVSS.n1302 547.1
R11559 DVSS.n4967 DVSS.n4966 547.1
R11560 DVSS.n4955 DVSS.n4954 547.1
R11561 DVSS.n3556 DVSS.n2661 517.379
R11562 DVSS.n4384 DVSS.n1312 488.243
R11563 DVSS.n4389 DVSS.n4388 488.243
R11564 DVSS.n1454 DVSS.n1287 488.243
R11565 DVSS.n1456 DVSS.n1295 488.243
R11566 DVSS.n3950 DVSS.n1504 486.896
R11567 DVSS.n3556 DVSS.n1702 478.878
R11568 DVSS.n3956 DVSS.n1504 472.783
R11569 DVSS.t188 DVSS.t98 463.173
R11570 DVSS.n3748 DVSS.n1701 447.923
R11571 DVSS.n4964 DVSS.t136 409.743
R11572 DVSS.n4956 DVSS.t81 409.743
R11573 DVSS.t70 DVSS.n4445 400.822
R11574 DVSS.n3752 DVSS.t11 367.289
R11575 DVSS.n3569 DVSS.n2249 344.332
R11576 DVSS.n3569 DVSS.n3568 344.332
R11577 DVSS.n3579 DVSS.n2244 344.332
R11578 DVSS.n3759 DVSS.n1695 344.332
R11579 DVSS.t150 DVSS.n1159 320.659
R11580 DVSS.t124 DVSS.n1586 306.072
R11581 DVSS.n1586 DVSS.t179 306.072
R11582 DVSS.t32 DVSS.n4383 303.188
R11583 DVSS.n4383 DVSS.t37 303.188
R11584 DVSS.n3568 DVSS.n3567 300.031
R11585 DVSS.n3567 DVSS.n3566 300.031
R11586 DVSS.n275 DVSS.t50 298.296
R11587 DVSS.n3621 DVSS.n3604 290.733
R11588 DVSS.n2246 DVSS.t105 287.95
R11589 DVSS.n3951 DVSS.n3950 285.283
R11590 DVSS.n5726 DVSS.t53 282.926
R11591 DVSS.n2241 DVSS.n2237 278.889
R11592 DVSS.n3957 DVSS.n1502 273.185
R11593 DVSS.t192 DVSS.t120 271.668
R11594 DVSS.t139 DVSS.t148 271.668
R11595 DVSS.t111 DVSS.t204 271.668
R11596 DVSS.t113 DVSS.t109 271.668
R11597 DVSS.t109 DVSS.t83 271.668
R11598 DVSS.t171 DVSS.n4430 271.668
R11599 DVSS.t152 DVSS.t171 271.668
R11600 DVSS.t32 DVSS.t99 271.668
R11601 DVSS.t190 DVSS.t169 271.668
R11602 DVSS.t169 DVSS.n4404 271.668
R11603 DVSS.t200 DVSS.t80 271.668
R11604 DVSS.n1511 DVSS.n1274 271
R11605 DVSS.n2263 DVSS.t62 270.834
R11606 DVSS.t204 DVSS.n1304 269.442
R11607 DVSS.n2660 DVSS.n2659 266.361
R11608 DVSS.n2255 DVSS.t15 256.738
R11609 DVSS.n3944 DVSS.n1515 255.427
R11610 DVSS.t120 DVSS.t200 252.742
R11611 DVSS.n4446 DVSS.t70 250.514
R11612 DVSS.n3566 DVSS.n3565 248.684
R11613 DVSS.t132 DVSS.t134 245.663
R11614 DVSS.t122 DVSS.t124 245.663
R11615 DVSS.t146 DVSS.t154 245.663
R11616 DVSS.t13 DVSS.t6 245.663
R11617 DVSS.t16 DVSS.t0 245.663
R11618 DVSS.t29 DVSS.t27 245.663
R11619 DVSS.n4486 DVSS.t161 241.587
R11620 DVSS.n3789 DVSS.t5 238.615
R11621 DVSS.t157 DVSS.n1695 235.595
R11622 DVSS.n1922 DVSS.n1921 233.749
R11623 DVSS.n2161 DVSS.n2160 233.749
R11624 DVSS.n4945 DVSS.n4944 232.701
R11625 DVSS.n3580 DVSS.n2243 227.541
R11626 DVSS.t37 DVSS.n1163 226.019
R11627 DVSS.n3978 DVSS.n1439 224.798
R11628 DVSS.n3623 DVSS.n3622 219.064
R11629 DVSS.n2262 DVSS.t18 216.465
R11630 DVSS.n2260 DVSS.t8 210.424
R11631 DVSS.n1481 DVSS.n1480 199.98
R11632 DVSS.t3 DVSS.n3760 192.303
R11633 DVSS.n4430 DVSS.t156 191.505
R11634 DVSS.n1447 DVSS.t95 188.571
R11635 DVSS.n2661 DVSS.n2254 187.429
R11636 DVSS.t196 DVSS.n2260 180.22
R11637 DVSS.t126 DVSS.t115 170.153
R11638 DVSS.t128 DVSS.t25 170.153
R11639 DVSS.n2229 DVSS.n1730 169.606
R11640 DVSS.n3603 DVSS.t17 169.145
R11641 DVSS.n4945 DVSS.t148 168.124
R11642 DVSS.n3903 DVSS.t179 166.125
R11643 DVSS.n4431 DVSS.t152 165.897
R11644 DVSS.n4405 DVSS.t190 165.897
R11645 DVSS.n3751 DVSS.t9 164.453
R11646 DVSS.n4479 DVSS.t167 163.742
R11647 DVSS.t44 DVSS.t100 163.742
R11648 DVSS.t72 DVSS.t76 163.742
R11649 DVSS.t185 DVSS.t87 161.953
R11650 DVSS.t20 DVSS.t117 161.953
R11651 DVSS.n4457 DVSS.t173 161.728
R11652 DVSS.n4964 DVSS.t96 158.31
R11653 DVSS.n4956 DVSS.t194 158.31
R11654 DVSS.t197 DVSS.t63 154.043
R11655 DVSS.t144 DVSS.t173 153.675
R11656 DVSS.n4471 DVSS.t161 152.333
R11657 DVSS.n4488 DVSS.n1023 152.252
R11658 DVSS.n1169 DVSS.n1024 152.252
R11659 DVSS.t103 DVSS.n3587 151.023
R11660 DVSS.t156 DVSS.n1156 150.309
R11661 DVSS.n2659 DVSS.n2658 149.083
R11662 DVSS.n1490 DVSS.n1482 146.669
R11663 DVSS.n4968 DVSS.n4967 146.669
R11664 DVSS.n4954 DVSS.n4953 146.669
R11665 DVSS.n4478 DVSS.t202 145.624
R11666 DVSS.t99 DVSS.n1159 142.516
R11667 DVSS.t25 DVSS.n3761 137.935
R11668 DVSS.n3951 DVSS.n1274 137.097
R11669 DVSS.n1170 DVSS.t192 135.834
R11670 DVSS.n1170 DVSS.t139 135.834
R11671 DVSS.n4433 DVSS.t111 135.834
R11672 DVSS.n4433 DVSS.t113 135.834
R11673 DVSS.n2255 DVSS.t8 133.906
R11674 DVSS.n1478 DVSS.n1477 132.07
R11675 DVSS.n4445 DVSS.n1304 131.381
R11676 DVSS.n4465 DVSS.n1275 129.345
R11677 DVSS.n4406 DVSS.n1171 129.345
R11678 DVSS.n4459 DVSS.n1296 129.345
R11679 DVSS.n4434 DVSS.n4432 129.345
R11680 DVSS.n4485 DVSS.n1275 128.957
R11681 DVSS.n4943 DVSS.n1171 128.957
R11682 DVSS.t165 DVSS.t85 125.49
R11683 DVSS.n1587 DVSS.t122 123.838
R11684 DVSS.t78 DVSS.n3902 123.838
R11685 DVSS.n3762 DVSS.t23 123.838
R11686 DVSS.t40 DVSS.n1453 122.806
R11687 DVSS.t134 DVSS.n1587 121.826
R11688 DVSS.n3902 DVSS.t154 121.826
R11689 DVSS.n3790 DVSS.t183 121.826
R11690 DVSS.n3762 DVSS.t126 121.826
R11691 DVSS.t83 DVSS.n1156 121.361
R11692 DVSS.n2263 DVSS.t196 119.811
R11693 DVSS.n4404 DVSS.n1165 118.02
R11694 DVSS.n3960 DVSS.n1502 114.919
R11695 DVSS.n3966 DVSS.n1498 114.919
R11696 DVSS.n3967 DVSS.n3966 114.919
R11697 DVSS.n3969 DVSS.n3967 114.919
R11698 DVSS.n3969 DVSS.n3968 114.919
R11699 DVSS.n3978 DVSS.n3977 114.919
R11700 DVSS.n1477 DVSS.n1445 112.962
R11701 DVSS.n3976 DVSS.n3975 112.903
R11702 DVSS.n3968 DVSS.n1494 111.895
R11703 DVSS.n1708 DVSS.n1702 110.056
R11704 DVSS.n3752 DVSS.t157 108.737
R11705 DVSS.n3761 DVSS.t3 107.73
R11706 DVSS.t85 DVSS.n4454 106.701
R11707 DVSS.n4431 DVSS.t150 105.773
R11708 DVSS.n4405 DVSS.t188 105.773
R11709 DVSS.n3624 DVSS.n3623 102.416
R11710 DVSS.n4386 DVSS.n4381 102.356
R11711 DVSS.n1476 DVSS.n1458 102.356
R11712 DVSS.t163 DVSS.t56 101.332
R11713 DVSS.t177 DVSS.t199 101.332
R11714 DVSS.n4458 DVSS.t66 99.9902
R11715 DVSS.n4928 DVSS.n959 99.728
R11716 DVSS.n5356 DVSS.n958 99.7229
R11717 DVSS.n3960 DVSS.n3959 98.7908
R11718 DVSS.t18 DVSS.t197 91.6207
R11719 DVSS.t63 DVSS.t183 91.6207
R11720 DVSS.t31 DVSS.t13 91.6207
R11721 DVSS.n2246 DVSS.n2243 90.6139
R11722 DVSS.n1447 DVSS.t64 90.5952
R11723 DVSS.t40 DVSS.n1445 89.3577
R11724 DVSS.t92 DVSS.n5725 87.8106
R11725 DVSS.t15 DVSS.n2244 87.5934
R11726 DVSS.t11 DVSS.n3751 86.3383
R11727 DVSS.n5726 DVSS.n59 86.0408
R11728 DVSS.n4455 DVSS.t138 85.2266
R11729 DVSS.n3587 DVSS.n2238 82.5594
R11730 DVSS.n4472 DVSS.t130 81.8712
R11731 DVSS.t159 DVSS.n4472 81.8712
R11732 DVSS.n275 DVSS.n59 80.8661
R11733 DVSS.n4473 DVSS.t1 80.5291
R11734 DVSS.n3903 DVSS.t78 79.5389
R11735 DVSS.t115 DVSS.t128 75.5117
R11736 DVSS.n5725 DVSS.t141 74.1437
R11737 DVSS.t80 DVSS.n1165 73.4846
R11738 DVSS.n2163 DVSS.n1803 73.4718
R11739 DVSS.n2163 DVSS.n2162 73.4718
R11740 DVSS.n1924 DVSS.n1806 73.2997
R11741 DVSS.n1924 DVSS.n1923 73.2997
R11742 DVSS.n4444 DVSS.n1305 72.4894
R11743 DVSS.n1478 DVSS.t44 70.25
R11744 DVSS.n4491 DVSS.n958 69.3341
R11745 DVSS.n4928 DVSS.n4927 69.3341
R11746 DVSS.t60 DVSS.t5 67.4571
R11747 DVSS.t17 DVSS.t23 67.4571
R11748 DVSS.n1303 DVSS.t90 65.0944
R11749 DVSS.n3945 DVSS.n1274 64.5166
R11750 DVSS.n4466 DVSS.t64 63.7523
R11751 DVSS.n4458 DVSS.t68 63.7523
R11752 DVSS.t56 DVSS.t159 62.4102
R11753 DVSS.t1 DVSS.t163 62.4102
R11754 DVSS.t101 DVSS.t177 62.4102
R11755 DVSS.t199 DVSS.t175 62.4102
R11756 DVSS.n4386 DVSS.n4385 61.1338
R11757 DVSS.n4387 DVSS.n4386 61.1338
R11758 DVSS.n1458 DVSS.n1455 61.1338
R11759 DVSS.n1458 DVSS.n1457 61.1338
R11760 DVSS.n1452 DVSS.n1446 59.6561
R11761 DVSS.n2230 DVSS.n1731 59.6561
R11762 DVSS.n3753 DVSS.n1696 59.6561
R11763 DVSS.n3570 DVSS.n2248 59.6561
R11764 DVSS.n3565 DVSS.t132 59.4026
R11765 DVSS.n5724 DVSS.n59 58.4662
R11766 DVSS.n4454 DVSS.t76 57.0416
R11767 DVSS.n1305 DVSS.n1296 56.4672
R11768 DVSS.n4434 DVSS.n1305 56.4672
R11769 DVSS.n3758 DVSS.n1696 56.0005
R11770 DVSS.n2259 DVSS.n2256 56.0005
R11771 DVSS.n3570 DVSS.n2247 56.0005
R11772 DVSS.t202 DVSS.n4467 54.3573
R11773 DVSS.t6 DVSS.t16 53.3617
R11774 DVSS.n3760 DVSS.t29 53.3617
R11775 DVSS.n4479 DVSS.t175 53.0152
R11776 DVSS.n4447 DVSS.n1303 53.0152
R11777 DVSS.n3588 DVSS.t103 46.314
R11778 DVSS.t98 DVSS.n1163 45.6497
R11779 DVSS.n4467 DVSS.n4466 45.6334
R11780 DVSS.n1480 DVSS.t100 44.9623
R11781 DVSS.n1453 DVSS.t95 40.9359
R11782 DVSS.n4465 DVSS.n1287 40.8338
R11783 DVSS.n4406 DVSS.n4389 40.8338
R11784 DVSS.n4432 DVSS.n1312 40.8338
R11785 DVSS.n4459 DVSS.n1295 40.8338
R11786 DVSS.n1867 DVSS.n1814 40.2769
R11787 DVSS.n1867 DVSS.n1804 40.2769
R11788 DVSS.n3623 DVSS.n1721 39.6013
R11789 DVSS.n3748 DVSS.n1702 38.5005
R11790 DVSS.t138 DVSS.t165 38.2516
R11791 DVSS.n2252 DVSS.n2249 37.2527
R11792 DVSS.n1481 DVSS.t68 34.2252
R11793 DVSS.n3574 DVSS.n2245 33.0561
R11794 DVSS.n3790 DVSS.t31 32.2186
R11795 DVSS.n4455 DVSS.n1300 30.1987
R11796 DVSS.n5119 DVSS.n1079 29.2479
R11797 DVSS.n5120 DVSS.n5119 29.2479
R11798 DVSS.n5121 DVSS.n5120 29.2479
R11799 DVSS.n5121 DVSS.n1075 29.2479
R11800 DVSS.n5127 DVSS.n1075 29.2479
R11801 DVSS.n5128 DVSS.n5127 29.2479
R11802 DVSS.n5129 DVSS.n5128 29.2479
R11803 DVSS.n5129 DVSS.n1071 29.2479
R11804 DVSS.n5135 DVSS.n1071 29.2479
R11805 DVSS.n5136 DVSS.n5135 29.2479
R11806 DVSS.n5137 DVSS.n5136 29.2479
R11807 DVSS.n5137 DVSS.n1067 29.2479
R11808 DVSS.n5143 DVSS.n1067 29.2479
R11809 DVSS.n5144 DVSS.n5143 29.2479
R11810 DVSS.n5145 DVSS.n5144 29.2479
R11811 DVSS.n5145 DVSS.n1063 29.2479
R11812 DVSS.n5151 DVSS.n1063 29.2479
R11813 DVSS.n5152 DVSS.n5151 29.2479
R11814 DVSS.n5153 DVSS.n5152 29.2479
R11815 DVSS.n5153 DVSS.n1059 29.2479
R11816 DVSS.n5159 DVSS.n1059 29.2479
R11817 DVSS.n5160 DVSS.n5159 29.2479
R11818 DVSS.n5161 DVSS.n5160 29.2479
R11819 DVSS.n5161 DVSS.n1055 29.2479
R11820 DVSS.n5167 DVSS.n1055 29.2479
R11821 DVSS.n5168 DVSS.n5167 29.2479
R11822 DVSS.n5169 DVSS.n5168 29.2479
R11823 DVSS.n5169 DVSS.n1051 29.2479
R11824 DVSS.n5175 DVSS.n1051 29.2479
R11825 DVSS.n5176 DVSS.n5175 29.2479
R11826 DVSS.n5177 DVSS.n5176 29.2479
R11827 DVSS.n5177 DVSS.n1047 29.2479
R11828 DVSS.n5183 DVSS.n1047 29.2479
R11829 DVSS.n5184 DVSS.n5183 29.2479
R11830 DVSS.n5185 DVSS.n5184 29.2479
R11831 DVSS.n5185 DVSS.n1043 29.2479
R11832 DVSS.n5191 DVSS.n1043 29.2479
R11833 DVSS.n5192 DVSS.n5191 29.2479
R11834 DVSS.n5193 DVSS.n5192 29.2479
R11835 DVSS.n5193 DVSS.n1039 29.2479
R11836 DVSS.n5199 DVSS.n1039 29.2479
R11837 DVSS.n5200 DVSS.n5199 29.2479
R11838 DVSS.n5201 DVSS.n5200 29.2479
R11839 DVSS.n5201 DVSS.n1035 29.2479
R11840 DVSS.n5207 DVSS.n1035 29.2479
R11841 DVSS.n5208 DVSS.n5207 29.2479
R11842 DVSS.n5209 DVSS.n5208 29.2479
R11843 DVSS.n5209 DVSS.n1031 29.2479
R11844 DVSS.n5215 DVSS.n1031 29.2479
R11845 DVSS.n5216 DVSS.n5215 29.2479
R11846 DVSS.n5217 DVSS.n5216 29.2479
R11847 DVSS.n5217 DVSS.n1027 29.2479
R11848 DVSS.n5224 DVSS.n1027 29.2479
R11849 DVSS.n5225 DVSS.n5224 29.2479
R11850 DVSS.n5226 DVSS.n5225 29.2479
R11851 DVSS.n5226 DVSS.n1022 29.2479
R11852 DVSS.n5234 DVSS.n5233 29.2479
R11853 DVSS.n5234 DVSS.n1018 29.2479
R11854 DVSS.n5240 DVSS.n1018 29.2479
R11855 DVSS.n5241 DVSS.n5240 29.2479
R11856 DVSS.n5242 DVSS.n5241 29.2479
R11857 DVSS.n5242 DVSS.n1014 29.2479
R11858 DVSS.n5248 DVSS.n1014 29.2479
R11859 DVSS.n5249 DVSS.n5248 29.2479
R11860 DVSS.n5250 DVSS.n5249 29.2479
R11861 DVSS.n5250 DVSS.n1010 29.2479
R11862 DVSS.n5256 DVSS.n1010 29.2479
R11863 DVSS.n5257 DVSS.n5256 29.2479
R11864 DVSS.n5258 DVSS.n5257 29.2479
R11865 DVSS.n5258 DVSS.n1006 29.2479
R11866 DVSS.n5264 DVSS.n1006 29.2479
R11867 DVSS.n5265 DVSS.n5264 29.2479
R11868 DVSS.n5266 DVSS.n5265 29.2479
R11869 DVSS.n5266 DVSS.n1002 29.2479
R11870 DVSS.n5272 DVSS.n1002 29.2479
R11871 DVSS.n5273 DVSS.n5272 29.2479
R11872 DVSS.n5274 DVSS.n5273 29.2479
R11873 DVSS.n5274 DVSS.n998 29.2479
R11874 DVSS.n5280 DVSS.n998 29.2479
R11875 DVSS.n5281 DVSS.n5280 29.2479
R11876 DVSS.n5282 DVSS.n5281 29.2479
R11877 DVSS.n5282 DVSS.n994 29.2479
R11878 DVSS.n5288 DVSS.n994 29.2479
R11879 DVSS.n5289 DVSS.n5288 29.2479
R11880 DVSS.n5290 DVSS.n5289 29.2479
R11881 DVSS.n5290 DVSS.n990 29.2479
R11882 DVSS.n5296 DVSS.n990 29.2479
R11883 DVSS.n5297 DVSS.n5296 29.2479
R11884 DVSS.n5298 DVSS.n5297 29.2479
R11885 DVSS.n5298 DVSS.n986 29.2479
R11886 DVSS.n5304 DVSS.n986 29.2479
R11887 DVSS.n5305 DVSS.n5304 29.2479
R11888 DVSS.n5306 DVSS.n5305 29.2479
R11889 DVSS.n5306 DVSS.n982 29.2479
R11890 DVSS.n5312 DVSS.n982 29.2479
R11891 DVSS.n5313 DVSS.n5312 29.2479
R11892 DVSS.n5314 DVSS.n5313 29.2479
R11893 DVSS.n5314 DVSS.n978 29.2479
R11894 DVSS.n5320 DVSS.n978 29.2479
R11895 DVSS.n5321 DVSS.n5320 29.2479
R11896 DVSS.n5322 DVSS.n5321 29.2479
R11897 DVSS.n5322 DVSS.n974 29.2479
R11898 DVSS.n5328 DVSS.n974 29.2479
R11899 DVSS.n5329 DVSS.n5328 29.2479
R11900 DVSS.n5330 DVSS.n5329 29.2479
R11901 DVSS.n5330 DVSS.n970 29.2479
R11902 DVSS.n5336 DVSS.n970 29.2479
R11903 DVSS.n5337 DVSS.n5336 29.2479
R11904 DVSS.n5338 DVSS.n5337 29.2479
R11905 DVSS.n5338 DVSS.n966 29.2479
R11906 DVSS.n5345 DVSS.n966 29.2479
R11907 DVSS.n5346 DVSS.n5345 29.2479
R11908 DVSS.n5347 DVSS.n5346 29.2479
R11909 DVSS.n2241 DVSS.t146 29.1981
R11910 DVSS.t62 DVSS.n2262 29.1981
R11911 DVSS.n4447 DVSS.t74 28.8566
R11912 DVSS.n3578 DVSS.n2245 26.6005
R11913 DVSS.n2256 DVSS.n2245 26.6005
R11914 DVSS.n3580 DVSS.n3579 26.1777
R11915 DVSS.n5113 DVSS.n1079 21.9361
R11916 DVSS.n4487 DVSS.n4486 21.4748
R11917 DVSS.n4473 DVSS.t101 20.8037
R11918 DVSS.n3588 DVSS.n2237 20.1368
R11919 DVSS.n5349 DVSS.n962 19.8187
R11920 DVSS.t167 DVSS.n4478 18.1194
R11921 DVSS.t90 DVSS.t72 16.7773
R11922 DVSS.n3959 DVSS.n1498 16.1295
R11923 DVSS.n1279 DVSS.t207 15.9461
R11924 DVSS.n4435 DVSS.t209 15.9461
R11925 DVSS.n1461 DVSS.t208 15.9461
R11926 DVSS.n4397 DVSS.t206 15.9461
R11927 DVSS.n5351 DVSS.n963 14.9684
R11928 DVSS.n5233 DVSS.n5232 14.8601
R11929 DVSS.n5111 DVSS.n5110 14.6638
R11930 DVSS.n5232 DVSS.n1022 14.3883
R11931 DVSS.n3957 DVSS.n3956 14.1134
R11932 DVSS.n4189 DVSS.n4184 12.4433
R11933 DVSS.t105 DVSS.n2238 12.0823
R11934 DVSS.n5347 DVSS.n962 12.0297
R11935 DVSS.n3583 DVSS.n3582 11.7115
R11936 DVSS.t130 DVSS.n4471 11.4087
R11937 DVSS.n1487 VSS 10.8266
R11938 DVSS.n4973 VSS 10.8266
R11939 DVSS.n4950 VSS 10.8266
R11940 DVSS.n2655 DVSS.n2264 10.6065
R11941 DVSS.n5109 DVSS.n1081 10.6065
R11942 DVSS.n1479 DVSS.n1478 10.3873
R11943 DVSS.n1446 DVSS.n1445 10.1573
R11944 DVSS.n1300 DVSS.t144 10.0666
R11945 DVSS.n5114 DVSS.n5113 9.91235
R11946 DVSS.n3603 DVSS.t60 9.06184
R11947 DVSS.n3614 DVSS.t28 8.35531
R11948 DVSS.n3615 DVSS.t28 8.13558
R11949 DVSS.n2656 DVSS.n2655 8.06976
R11950 DVSS.n2656 DVSS.n1081 8.03441
R11951 DVSS.t74 DVSS.n4446 7.95592
R11952 DVSS.n1806 DVSS.n1804 7.77509
R11953 DVSS.n1923 DVSS.n1814 7.77509
R11954 DVSS.n4922 DVSS.n1194 7.61966
R11955 DVSS.n4678 DVSS.n1272 7.60677
R11956 DVSS.n4678 DVSS.n1217 7.60677
R11957 DVSS.n1814 DVSS.n1803 7.60296
R11958 DVSS.n2162 DVSS.n1804 7.60296
R11959 DVSS.n4674 DVSS.n1272 7.59387
R11960 DVSS.n4922 DVSS.n1217 7.58957
R11961 DVSS.n4927 DVSS.n1194 7.28428
R11962 DVSS.n4674 DVSS.n4491 7.26279
R11963 DVSS.t0 DVSS.n3789 7.04821
R11964 DVSS.n3573 DVSS.n3572 6.95655
R11965 DVSS.n1733 DVSS.n1732 6.3005
R11966 DVSS.n4426 DVSS.n4425 6.3005
R11967 DVSS.n1471 DVSS.n1470 6.3005
R11968 DVSS.n4187 DVSS.n4186 6.3005
R11969 DVSS.n3608 DVSS.n3607 6.3005
R11970 DVSS.n4392 DVSS.n4391 6.3005
R11971 DVSS.n4338 DVSS.n4337 6.3005
R11972 DVSS.n2264 DVSS.n963 6.19648
R11973 DVSS.n5110 DVSS.n5109 6.19648
R11974 DVSS.n3756 DVSS.n1698 5.57932
R11975 DVSS.n4933 DVSS.n4932 5.42247
R11976 VSS DVSS.n1486 5.2005
R11977 VSS DVSS.n1485 5.2005
R11978 VSS DVSS.n4972 5.2005
R11979 VSS DVSS.n4971 5.2005
R11980 VSS DVSS.n4949 5.2005
R11981 VSS DVSS.n4948 5.2005
R11982 DVSS.n3647 DVSS.n1715 5.2005
R11983 DVSS.n3647 DVSS.n3646 5.2005
R11984 DVSS.n1721 DVSS.n1715 5.2005
R11985 DVSS.n3594 DVSS.n1721 5.2005
R11986 DVSS.n1729 DVSS.n1721 5.2005
R11987 DVSS.n3595 DVSS.n1721 5.2005
R11988 DVSS.n1728 DVSS.n1721 5.2005
R11989 DVSS.n3596 DVSS.n1721 5.2005
R11990 DVSS.n1727 DVSS.n1721 5.2005
R11991 DVSS.n3597 DVSS.n1721 5.2005
R11992 DVSS.n1726 DVSS.n1721 5.2005
R11993 DVSS.n3644 DVSS.n1721 5.2005
R11994 DVSS.n3628 DVSS.n1721 5.2005
R11995 DVSS.n3646 DVSS.n1721 5.2005
R11996 DVSS.n1719 DVSS.n1715 5.2005
R11997 DVSS.n3594 DVSS.n1719 5.2005
R11998 DVSS.n1729 DVSS.n1719 5.2005
R11999 DVSS.n3595 DVSS.n1719 5.2005
R12000 DVSS.n1728 DVSS.n1719 5.2005
R12001 DVSS.n3596 DVSS.n1719 5.2005
R12002 DVSS.n1727 DVSS.n1719 5.2005
R12003 DVSS.n3597 DVSS.n1719 5.2005
R12004 DVSS.n1726 DVSS.n1719 5.2005
R12005 DVSS.n3644 DVSS.n1719 5.2005
R12006 DVSS.n3646 DVSS.n1719 5.2005
R12007 DVSS.n1722 DVSS.n1715 5.2005
R12008 DVSS.n3594 DVSS.n1722 5.2005
R12009 DVSS.n1729 DVSS.n1722 5.2005
R12010 DVSS.n3595 DVSS.n1722 5.2005
R12011 DVSS.n1728 DVSS.n1722 5.2005
R12012 DVSS.n3596 DVSS.n1722 5.2005
R12013 DVSS.n1727 DVSS.n1722 5.2005
R12014 DVSS.n3597 DVSS.n1722 5.2005
R12015 DVSS.n1726 DVSS.n1722 5.2005
R12016 DVSS.n3644 DVSS.n1722 5.2005
R12017 DVSS.n3646 DVSS.n1722 5.2005
R12018 DVSS.n1718 DVSS.n1715 5.2005
R12019 DVSS.n3594 DVSS.n1718 5.2005
R12020 DVSS.n1729 DVSS.n1718 5.2005
R12021 DVSS.n3595 DVSS.n1718 5.2005
R12022 DVSS.n1728 DVSS.n1718 5.2005
R12023 DVSS.n3596 DVSS.n1718 5.2005
R12024 DVSS.n1727 DVSS.n1718 5.2005
R12025 DVSS.n3597 DVSS.n1718 5.2005
R12026 DVSS.n1726 DVSS.n1718 5.2005
R12027 DVSS.n3644 DVSS.n1718 5.2005
R12028 DVSS.n3646 DVSS.n1718 5.2005
R12029 DVSS.n1723 DVSS.n1715 5.2005
R12030 DVSS.n3594 DVSS.n1723 5.2005
R12031 DVSS.n1729 DVSS.n1723 5.2005
R12032 DVSS.n3595 DVSS.n1723 5.2005
R12033 DVSS.n1728 DVSS.n1723 5.2005
R12034 DVSS.n3596 DVSS.n1723 5.2005
R12035 DVSS.n1727 DVSS.n1723 5.2005
R12036 DVSS.n3597 DVSS.n1723 5.2005
R12037 DVSS.n1726 DVSS.n1723 5.2005
R12038 DVSS.n3644 DVSS.n1723 5.2005
R12039 DVSS.n3646 DVSS.n1723 5.2005
R12040 DVSS.n1717 DVSS.n1715 5.2005
R12041 DVSS.n3594 DVSS.n1717 5.2005
R12042 DVSS.n1729 DVSS.n1717 5.2005
R12043 DVSS.n3595 DVSS.n1717 5.2005
R12044 DVSS.n1728 DVSS.n1717 5.2005
R12045 DVSS.n3596 DVSS.n1717 5.2005
R12046 DVSS.n1727 DVSS.n1717 5.2005
R12047 DVSS.n3597 DVSS.n1717 5.2005
R12048 DVSS.n1726 DVSS.n1717 5.2005
R12049 DVSS.n3644 DVSS.n1717 5.2005
R12050 DVSS.n3646 DVSS.n1717 5.2005
R12051 DVSS.n3645 DVSS.n3594 5.2005
R12052 DVSS.n3645 DVSS.n1729 5.2005
R12053 DVSS.n3645 DVSS.n3595 5.2005
R12054 DVSS.n3645 DVSS.n1728 5.2005
R12055 DVSS.n3645 DVSS.n3596 5.2005
R12056 DVSS.n3645 DVSS.n1727 5.2005
R12057 DVSS.n3645 DVSS.n3597 5.2005
R12058 DVSS.n3645 DVSS.n1726 5.2005
R12059 DVSS.n3645 DVSS.n3644 5.2005
R12060 DVSS.n3646 DVSS.n3645 5.2005
R12061 DVSS.n4184 DVSS.n1368 5.08553
R12062 DVSS.n3624 DVSS.n1716 4.84618
R12063 DVSS.n3632 DVSS.n1719 4.84618
R12064 DVSS.n3626 DVSS.n1722 4.84618
R12065 DVSS.n3631 DVSS.n1718 4.84618
R12066 DVSS.n3627 DVSS.n1723 4.84618
R12067 DVSS.n3630 DVSS.n1717 4.84618
R12068 DVSS.n3645 DVSS.n1725 4.84618
R12069 DVSS.n3647 DVSS.n1716 4.84618
R12070 DVSS.n3632 DVSS.n1721 4.84618
R12071 DVSS.n3626 DVSS.n1719 4.84618
R12072 DVSS.n3631 DVSS.n1722 4.84618
R12073 DVSS.n3627 DVSS.n1718 4.84618
R12074 DVSS.n3630 DVSS.n1723 4.84618
R12075 DVSS.n1725 DVSS.n1717 4.84618
R12076 DVSS.n3947 DVSS.n1101 4.82802
R12077 DVSS.n5057 DVSS.n1110 4.66866
R12078 DVSS.n5045 DVSS.n1121 4.66866
R12079 DVSS.n4821 DVSS.n4820 4.5005
R12080 DVSS.n4820 DVSS.n4812 4.5005
R12081 DVSS.n4820 DVSS.n4810 4.5005
R12082 DVSS.n4819 DVSS.n4814 4.5005
R12083 DVSS.n4820 DVSS.n4819 4.5005
R12084 DVSS.n4872 DVSS.n4807 4.5005
R12085 DVSS.n4830 DVSS.n4807 4.5005
R12086 DVSS.n4875 DVSS.n4807 4.5005
R12087 DVSS.n4872 DVSS.n4822 4.5005
R12088 DVSS.n4875 DVSS.n4822 4.5005
R12089 DVSS.n4875 DVSS.n4806 4.5005
R12090 DVSS.n4875 DVSS.n4823 4.5005
R12091 DVSS.n4875 DVSS.n4805 4.5005
R12092 DVSS.n4875 DVSS.n4824 4.5005
R12093 DVSS.n4875 DVSS.n4804 4.5005
R12094 DVSS.n4875 DVSS.n4825 4.5005
R12095 DVSS.n4875 DVSS.n4803 4.5005
R12096 DVSS.n4874 DVSS.n4830 4.5005
R12097 DVSS.n4875 DVSS.n4874 4.5005
R12098 DVSS.n4539 DVSS.n4509 4.5005
R12099 DVSS.n4544 DVSS.n4539 4.5005
R12100 DVSS.n4539 DVSS.n4511 4.5005
R12101 DVSS.n4527 DVSS.n4509 4.5005
R12102 DVSS.n4527 DVSS.n4511 4.5005
R12103 DVSS.n4523 DVSS.n4511 4.5005
R12104 DVSS.n4521 DVSS.n4511 4.5005
R12105 DVSS.n4519 DVSS.n4511 4.5005
R12106 DVSS.n4517 DVSS.n4511 4.5005
R12107 DVSS.n4515 DVSS.n4511 4.5005
R12108 DVSS.n4513 DVSS.n4511 4.5005
R12109 DVSS.n4541 DVSS.n4511 4.5005
R12110 DVSS.n4544 DVSS.n4543 4.5005
R12111 DVSS.n4543 DVSS.n4511 4.5005
R12112 DVSS.n4538 DVSS.n4537 4.5005
R12113 DVSS.n4537 DVSS.n4525 4.5005
R12114 DVSS.n4535 DVSS.n4525 4.5005
R12115 DVSS.n4535 DVSS.n4534 4.5005
R12116 DVSS.n4535 DVSS.n4532 4.5005
R12117 DVSS.n4537 DVSS.n4536 4.5005
R12118 DVSS.n4536 DVSS.n4535 4.5005
R12119 DVSS.n1855 DVSS.n1854 4.5005
R12120 DVSS.n1865 DVSS.n1858 4.5005
R12121 DVSS.n1866 DVSS.n1854 4.5005
R12122 DVSS.n1866 DVSS.n1853 4.5005
R12123 DVSS.n1866 DVSS.n1865 4.5005
R12124 DVSS.n4093 DVSS.n1430 4.5005
R12125 DVSS.n1436 DVSS.n1430 4.5005
R12126 DVSS.n4095 DVSS.n1430 4.5005
R12127 DVSS.n4093 DVSS.n1432 4.5005
R12128 DVSS.n1436 DVSS.n1432 4.5005
R12129 DVSS.n4095 DVSS.n1432 4.5005
R12130 DVSS.n4095 DVSS.n1429 4.5005
R12131 DVSS.n1436 DVSS.n1429 4.5005
R12132 DVSS.n4093 DVSS.n1429 4.5005
R12133 DVSS.n4095 DVSS.n1433 4.5005
R12134 DVSS.n1436 DVSS.n1433 4.5005
R12135 DVSS.n4093 DVSS.n1433 4.5005
R12136 DVSS.n4093 DVSS.n1428 4.5005
R12137 DVSS.n1436 DVSS.n1428 4.5005
R12138 DVSS.n4095 DVSS.n1428 4.5005
R12139 DVSS.n4095 DVSS.n1434 4.5005
R12140 DVSS.n1436 DVSS.n1434 4.5005
R12141 DVSS.n4093 DVSS.n1434 4.5005
R12142 DVSS.n4093 DVSS.n1427 4.5005
R12143 DVSS.n1436 DVSS.n1427 4.5005
R12144 DVSS.n4095 DVSS.n1427 4.5005
R12145 DVSS.n4095 DVSS.n4094 4.5005
R12146 DVSS.n4094 DVSS.n1436 4.5005
R12147 DVSS.n4094 DVSS.n4093 4.5005
R12148 DVSS.n1383 DVSS.n1378 4.5005
R12149 DVSS.n4170 DVSS.n1383 4.5005
R12150 DVSS.n4168 DVSS.n1383 4.5005
R12151 DVSS.n1385 DVSS.n1378 4.5005
R12152 DVSS.n4170 DVSS.n1385 4.5005
R12153 DVSS.n4168 DVSS.n1385 4.5005
R12154 DVSS.n4168 DVSS.n1382 4.5005
R12155 DVSS.n4170 DVSS.n1382 4.5005
R12156 DVSS.n1382 DVSS.n1378 4.5005
R12157 DVSS.n1386 DVSS.n1378 4.5005
R12158 DVSS.n4170 DVSS.n1386 4.5005
R12159 DVSS.n4168 DVSS.n1386 4.5005
R12160 DVSS.n1381 DVSS.n1378 4.5005
R12161 DVSS.n4170 DVSS.n1381 4.5005
R12162 DVSS.n4168 DVSS.n1381 4.5005
R12163 DVSS.n4168 DVSS.n1387 4.5005
R12164 DVSS.n4170 DVSS.n1387 4.5005
R12165 DVSS.n1387 DVSS.n1378 4.5005
R12166 DVSS.n4168 DVSS.n1380 4.5005
R12167 DVSS.n4170 DVSS.n1380 4.5005
R12168 DVSS.n1380 DVSS.n1378 4.5005
R12169 DVSS.n1388 DVSS.n1378 4.5005
R12170 DVSS.n4170 DVSS.n1388 4.5005
R12171 DVSS.n4168 DVSS.n1388 4.5005
R12172 DVSS.n4168 DVSS.n1379 4.5005
R12173 DVSS.n4170 DVSS.n1379 4.5005
R12174 DVSS.n1379 DVSS.n1378 4.5005
R12175 DVSS.n4169 DVSS.n4168 4.5005
R12176 DVSS.n4170 DVSS.n4169 4.5005
R12177 DVSS.n4169 DVSS.n1378 4.5005
R12178 DVSS.n2170 DVSS.n1796 4.5005
R12179 DVSS.n1799 DVSS.n1796 4.5005
R12180 DVSS.n2169 DVSS.n1799 4.5005
R12181 DVSS.n2170 DVSS.n2169 4.5005
R12182 DVSS.n2146 DVSS.n1797 4.5005
R12183 DVSS.n2150 DVSS.n1797 4.5005
R12184 DVSS.n1817 DVSS.n1744 4.5005
R12185 DVSS.n1831 DVSS.n1740 4.5005
R12186 DVSS.n1831 DVSS.n1744 4.5005
R12187 DVSS.n1819 DVSS.n1740 4.5005
R12188 DVSS.n1819 DVSS.n1744 4.5005
R12189 DVSS.n1817 DVSS.n1740 4.5005
R12190 DVSS.n1919 DVSS.n1740 4.5005
R12191 DVSS.n1919 DVSS.n1744 4.5005
R12192 DVSS.n2180 DVSS.n1787 4.5005
R12193 DVSS.n2180 DVSS.n2179 4.5005
R12194 DVSS.n2179 DVSS.n2178 4.5005
R12195 DVSS.n2178 DVSS.n1787 4.5005
R12196 DVSS.n1877 DVSS.n1788 4.5005
R12197 DVSS.n1878 DVSS.n1877 4.5005
R12198 DVSS.n1981 DVSS.n1959 4.5005
R12199 DVSS.n1960 DVSS.n1959 4.5005
R12200 DVSS.n1961 DVSS.n1959 4.5005
R12201 DVSS.n1983 DVSS.n1959 4.5005
R12202 DVSS.n1983 DVSS.n1982 4.5005
R12203 DVSS.n1982 DVSS.n1961 4.5005
R12204 DVSS.n1982 DVSS.n1960 4.5005
R12205 DVSS.n1982 DVSS.n1981 4.5005
R12206 DVSS.n1977 DVSS.n1965 4.5005
R12207 DVSS.n1980 DVSS.n1965 4.5005
R12208 DVSS.n1980 DVSS.n1979 4.5005
R12209 DVSS.n1980 DVSS.n1964 4.5005
R12210 DVSS.n1977 DVSS.n1812 4.5005
R12211 DVSS.n1980 DVSS.n1812 4.5005
R12212 DVSS.n2101 DVSS.n1809 4.5005
R12213 DVSS.n2101 DVSS.n1810 4.5005
R12214 DVSS.n2158 DVSS.n1809 4.5005
R12215 DVSS.n2158 DVSS.n1810 4.5005
R12216 DVSS.n2107 DVSS.n1810 4.5005
R12217 DVSS.n2107 DVSS.n1809 4.5005
R12218 DVSS.n2116 DVSS.n2086 4.5005
R12219 DVSS.n2088 DVSS.n2086 4.5005
R12220 DVSS.n2115 DVSS.n2088 4.5005
R12221 DVSS.n2116 DVSS.n2115 4.5005
R12222 DVSS.n2105 DVSS.n1810 4.5005
R12223 DVSS.n2105 DVSS.n1809 4.5005
R12224 DVSS.n2159 DVSS.n2158 4.5005
R12225 DVSS.n1920 DVSS.n1919 4.5005
R12226 DVSS.n1919 DVSS.n1918 4.5005
R12227 DVSS.n2158 DVSS.n2157 4.5005
R12228 DVSS.n2112 DVSS.n2089 4.5005
R12229 DVSS.n2113 DVSS.n2112 4.5005
R12230 DVSS.n1943 DVSS.n1941 4.5005
R12231 DVSS.n1949 DVSS.n1943 4.5005
R12232 DVSS.n2114 DVSS.n2089 4.5005
R12233 DVSS.n2114 DVSS.n2113 4.5005
R12234 DVSS.n2166 DVSS.n1802 4.5005
R12235 DVSS.n2166 DVSS.n2165 4.5005
R12236 DVSS.n2181 DVSS.n1786 4.5005
R12237 DVSS.n2181 DVSS.n1783 4.5005
R12238 DVSS.n1754 DVSS.n1751 4.5005
R12239 DVSS.n1774 DVSS.n1754 4.5005
R12240 DVSS.n2198 DVSS.n1759 4.5005
R12241 DVSS.n2198 DVSS.n1761 4.5005
R12242 DVSS.n2198 DVSS.n1758 4.5005
R12243 DVSS.n2198 DVSS.n2197 4.5005
R12244 DVSS.n2197 DVSS.n2196 4.5005
R12245 DVSS.n2196 DVSS.n1758 4.5005
R12246 DVSS.n2196 DVSS.n1761 4.5005
R12247 DVSS.n2196 DVSS.n1759 4.5005
R12248 DVSS.n1882 DVSS.n1760 4.5005
R12249 DVSS.n1913 DVSS.n1760 4.5005
R12250 DVSS.n1913 DVSS.n1912 4.5005
R12251 DVSS.n1913 DVSS.n1883 4.5005
R12252 DVSS.n1914 DVSS.n1882 4.5005
R12253 DVSS.n1914 DVSS.n1913 4.5005
R12254 DVSS.n2207 DVSS.n1749 4.5005
R12255 DVSS.n2203 DVSS.n1749 4.5005
R12256 DVSS.n1899 DVSS.n1889 4.5005
R12257 DVSS.n1891 DVSS.n1889 4.5005
R12258 DVSS.n1901 DVSS.n1889 4.5005
R12259 DVSS.n1901 DVSS.n1900 4.5005
R12260 DVSS.n1900 DVSS.n1891 4.5005
R12261 DVSS.n1900 DVSS.n1899 4.5005
R12262 DVSS.n1890 DVSS.n1620 4.5005
R12263 DVSS.n1890 DVSS.n1625 4.5005
R12264 DVSS.n1631 DVSS.n1620 4.5005
R12265 DVSS.n3840 DVSS.n1629 4.5005
R12266 DVSS.n3840 DVSS.n3831 4.5005
R12267 DVSS.n3840 DVSS.n1628 4.5005
R12268 DVSS.n3840 DVSS.n3834 4.5005
R12269 DVSS.n3840 DVSS.n1627 4.5005
R12270 DVSS.n3840 DVSS.n3837 4.5005
R12271 DVSS.n3840 DVSS.n1626 4.5005
R12272 DVSS.n3839 DVSS.n1625 4.5005
R12273 DVSS.n3840 DVSS.n3839 4.5005
R12274 DVSS.n1487 VSS 4.5005
R12275 DVSS.n4973 VSS 4.5005
R12276 DVSS.n5045 DVSS.n5044 4.5005
R12277 DVSS.n5047 DVSS.n5046 4.5005
R12278 DVSS.n1120 DVSS.n1118 4.5005
R12279 DVSS.n1113 DVSS.n1112 4.5005
R12280 DVSS.n5056 DVSS.n5055 4.5005
R12281 DVSS.n5058 DVSS.n5057 4.5005
R12282 DVSS.n2420 DVSS.n2278 4.5005
R12283 DVSS.n2420 DVSS.n2275 4.5005
R12284 DVSS.n2408 DVSS.n2278 4.5005
R12285 DVSS.n2419 DVSS.n2281 4.5005
R12286 DVSS.n2419 DVSS.n2406 4.5005
R12287 DVSS.n2419 DVSS.n2280 4.5005
R12288 DVSS.n2419 DVSS.n2408 4.5005
R12289 DVSS.n2420 DVSS.n2419 4.5005
R12290 DVSS.n2410 DVSS.n2275 4.5005
R12291 DVSS.n2412 DVSS.n2275 4.5005
R12292 DVSS.n2414 DVSS.n2275 4.5005
R12293 DVSS.n2416 DVSS.n2275 4.5005
R12294 DVSS.n2419 DVSS.n2418 4.5005
R12295 DVSS.n2418 DVSS.n2275 4.5005
R12296 DVSS.n4950 VSS 4.5005
R12297 DVSS.n2648 DVSS.n1699 4.5005
R12298 DVSS.n2646 DVSS.n1699 4.5005
R12299 DVSS.n2646 DVSS.n2637 4.5005
R12300 DVSS.n2646 DVSS.n2425 4.5005
R12301 DVSS.n2646 DVSS.n2638 4.5005
R12302 DVSS.n2646 DVSS.n2424 4.5005
R12303 DVSS.n2646 DVSS.n2639 4.5005
R12304 DVSS.n2646 DVSS.n2423 4.5005
R12305 DVSS.n2646 DVSS.n2645 4.5005
R12306 DVSS.n2646 DVSS.n2422 4.5005
R12307 DVSS.n2648 DVSS.n2647 4.5005
R12308 DVSS.n2647 DVSS.n2646 4.5005
R12309 DVSS.n4934 DVSS.n1185 4.5005
R12310 DVSS.n1185 DVSS.n1177 4.5005
R12311 DVSS.n1185 DVSS.n1178 4.5005
R12312 DVSS.n1185 DVSS.n1180 4.5005
R12313 DVSS.n1182 DVSS.n1178 4.5005
R12314 DVSS.n1182 DVSS.n1180 4.5005
R12315 DVSS.n4934 DVSS.n1186 4.5005
R12316 DVSS.n1186 DVSS.n1177 4.5005
R12317 DVSS.n1186 DVSS.n1178 4.5005
R12318 DVSS.n1186 DVSS.n1180 4.5005
R12319 DVSS.n4934 DVSS.n1184 4.5005
R12320 DVSS.n1184 DVSS.n1177 4.5005
R12321 DVSS.n1184 DVSS.n1178 4.5005
R12322 DVSS.n1184 DVSS.n1180 4.5005
R12323 DVSS.n1189 DVSS.n1178 4.5005
R12324 DVSS.n1189 DVSS.n1180 4.5005
R12325 DVSS.n1183 DVSS.n1178 4.5005
R12326 DVSS.n1183 DVSS.n1180 4.5005
R12327 DVSS.n4934 DVSS.n1187 4.5005
R12328 DVSS.n1187 DVSS.n1177 4.5005
R12329 DVSS.n1187 DVSS.n1178 4.5005
R12330 DVSS.n1187 DVSS.n1180 4.5005
R12331 DVSS.n1188 DVSS.n1178 4.5005
R12332 DVSS.n1188 DVSS.n1180 4.5005
R12333 DVSS.n4935 DVSS.n1178 4.5005
R12334 DVSS.n4935 DVSS.n1180 4.5005
R12335 DVSS.n4935 DVSS.n1177 4.5005
R12336 DVSS.n4935 DVSS.n4934 4.5005
R12337 DVSS.n1188 DVSS.n1177 4.5005
R12338 DVSS.n4934 DVSS.n1188 4.5005
R12339 DVSS.n1183 DVSS.n1177 4.5005
R12340 DVSS.n4934 DVSS.n1183 4.5005
R12341 DVSS.n1189 DVSS.n1177 4.5005
R12342 DVSS.n4934 DVSS.n1189 4.5005
R12343 DVSS.n1182 DVSS.n1177 4.5005
R12344 DVSS.n4934 DVSS.n1182 4.5005
R12345 DVSS.n4933 DVSS.n1180 4.5005
R12346 DVSS.n4933 DVSS.n1178 4.5005
R12347 DVSS.n4933 DVSS.n1177 4.5005
R12348 DVSS.n4934 DVSS.n4933 4.5005
R12349 DVSS.n5554 DVSS.n5553 4.5005
R12350 DVSS.n4932 DVSS.n855 4.5005
R12351 DVSS.n5557 DVSS.n6 4.5005
R12352 DVSS.n5812 DVSS.n5811 4.5005
R12353 DVSS.n5555 DVSS.n829 4.5005
R12354 DVSS.n5560 DVSS.n5559 4.5005
R12355 DVSS.n3755 DVSS.n1699 4.24863
R12356 DVSS.n3605 DVSS.t10 4.10856
R12357 DVSS.n3606 DVSS.t12 4.10856
R12358 DVSS.n5114 DVSS.n1080 4.05657
R12359 DVSS.n5118 DVSS.n1080 4.05657
R12360 DVSS.n5118 DVSS.n1078 4.05657
R12361 DVSS.n5122 DVSS.n1078 4.05657
R12362 DVSS.n5122 DVSS.n1076 4.05657
R12363 DVSS.n5126 DVSS.n1076 4.05657
R12364 DVSS.n5126 DVSS.n1074 4.05657
R12365 DVSS.n5130 DVSS.n1074 4.05657
R12366 DVSS.n5130 DVSS.n1072 4.05657
R12367 DVSS.n5134 DVSS.n1072 4.05657
R12368 DVSS.n5134 DVSS.n1070 4.05657
R12369 DVSS.n5138 DVSS.n1070 4.05657
R12370 DVSS.n5138 DVSS.n1068 4.05657
R12371 DVSS.n5142 DVSS.n1068 4.05657
R12372 DVSS.n5142 DVSS.n1066 4.05657
R12373 DVSS.n5146 DVSS.n1066 4.05657
R12374 DVSS.n5146 DVSS.n1064 4.05657
R12375 DVSS.n5150 DVSS.n1064 4.05657
R12376 DVSS.n5150 DVSS.n1062 4.05657
R12377 DVSS.n5154 DVSS.n1062 4.05657
R12378 DVSS.n5154 DVSS.n1060 4.05657
R12379 DVSS.n5158 DVSS.n1060 4.05657
R12380 DVSS.n5158 DVSS.n1058 4.05657
R12381 DVSS.n5162 DVSS.n1058 4.05657
R12382 DVSS.n5162 DVSS.n1056 4.05657
R12383 DVSS.n5166 DVSS.n1056 4.05657
R12384 DVSS.n5166 DVSS.n1054 4.05657
R12385 DVSS.n5170 DVSS.n1054 4.05657
R12386 DVSS.n5170 DVSS.n1052 4.05657
R12387 DVSS.n5174 DVSS.n1052 4.05657
R12388 DVSS.n5174 DVSS.n1050 4.05657
R12389 DVSS.n5178 DVSS.n1050 4.05657
R12390 DVSS.n5178 DVSS.n1048 4.05657
R12391 DVSS.n5182 DVSS.n1048 4.05657
R12392 DVSS.n5182 DVSS.n1046 4.05657
R12393 DVSS.n5186 DVSS.n1046 4.05657
R12394 DVSS.n5186 DVSS.n1044 4.05657
R12395 DVSS.n5190 DVSS.n1044 4.05657
R12396 DVSS.n5190 DVSS.n1042 4.05657
R12397 DVSS.n5194 DVSS.n1042 4.05657
R12398 DVSS.n5194 DVSS.n1040 4.05657
R12399 DVSS.n5198 DVSS.n1040 4.05657
R12400 DVSS.n5198 DVSS.n1038 4.05657
R12401 DVSS.n5202 DVSS.n1038 4.05657
R12402 DVSS.n5202 DVSS.n1036 4.05657
R12403 DVSS.n5206 DVSS.n1036 4.05657
R12404 DVSS.n5206 DVSS.n1034 4.05657
R12405 DVSS.n5210 DVSS.n1034 4.05657
R12406 DVSS.n5210 DVSS.n1032 4.05657
R12407 DVSS.n5214 DVSS.n1032 4.05657
R12408 DVSS.n5214 DVSS.n1030 4.05657
R12409 DVSS.n5218 DVSS.n1030 4.05657
R12410 DVSS.n5218 DVSS.n1028 4.05657
R12411 DVSS.n5223 DVSS.n1028 4.05657
R12412 DVSS.n5223 DVSS.n1026 4.05657
R12413 DVSS.n5227 DVSS.n1026 4.05657
R12414 DVSS.n5228 DVSS.n5227 4.05657
R12415 DVSS.n5228 DVSS.n1021 4.05657
R12416 DVSS.n5235 DVSS.n1021 4.05657
R12417 DVSS.n5235 DVSS.n1019 4.05657
R12418 DVSS.n5239 DVSS.n1019 4.05657
R12419 DVSS.n5239 DVSS.n1017 4.05657
R12420 DVSS.n5243 DVSS.n1017 4.05657
R12421 DVSS.n5243 DVSS.n1015 4.05657
R12422 DVSS.n5247 DVSS.n1015 4.05657
R12423 DVSS.n5247 DVSS.n1013 4.05657
R12424 DVSS.n5251 DVSS.n1013 4.05657
R12425 DVSS.n5251 DVSS.n1011 4.05657
R12426 DVSS.n5255 DVSS.n1011 4.05657
R12427 DVSS.n5255 DVSS.n1009 4.05657
R12428 DVSS.n5259 DVSS.n1009 4.05657
R12429 DVSS.n5259 DVSS.n1007 4.05657
R12430 DVSS.n5263 DVSS.n1007 4.05657
R12431 DVSS.n5263 DVSS.n1005 4.05657
R12432 DVSS.n5267 DVSS.n1005 4.05657
R12433 DVSS.n5267 DVSS.n1003 4.05657
R12434 DVSS.n5271 DVSS.n1003 4.05657
R12435 DVSS.n5271 DVSS.n1001 4.05657
R12436 DVSS.n5275 DVSS.n1001 4.05657
R12437 DVSS.n5275 DVSS.n999 4.05657
R12438 DVSS.n5279 DVSS.n999 4.05657
R12439 DVSS.n5279 DVSS.n997 4.05657
R12440 DVSS.n5283 DVSS.n997 4.05657
R12441 DVSS.n5283 DVSS.n995 4.05657
R12442 DVSS.n5287 DVSS.n995 4.05657
R12443 DVSS.n5287 DVSS.n993 4.05657
R12444 DVSS.n5291 DVSS.n993 4.05657
R12445 DVSS.n5291 DVSS.n991 4.05657
R12446 DVSS.n5295 DVSS.n991 4.05657
R12447 DVSS.n5295 DVSS.n989 4.05657
R12448 DVSS.n5299 DVSS.n989 4.05657
R12449 DVSS.n5299 DVSS.n987 4.05657
R12450 DVSS.n5303 DVSS.n987 4.05657
R12451 DVSS.n5303 DVSS.n985 4.05657
R12452 DVSS.n5307 DVSS.n985 4.05657
R12453 DVSS.n5307 DVSS.n983 4.05657
R12454 DVSS.n5311 DVSS.n983 4.05657
R12455 DVSS.n5311 DVSS.n981 4.05657
R12456 DVSS.n5315 DVSS.n981 4.05657
R12457 DVSS.n5315 DVSS.n979 4.05657
R12458 DVSS.n5319 DVSS.n979 4.05657
R12459 DVSS.n5319 DVSS.n977 4.05657
R12460 DVSS.n5323 DVSS.n977 4.05657
R12461 DVSS.n5323 DVSS.n975 4.05657
R12462 DVSS.n5327 DVSS.n975 4.05657
R12463 DVSS.n5327 DVSS.n973 4.05657
R12464 DVSS.n5331 DVSS.n973 4.05657
R12465 DVSS.n5331 DVSS.n971 4.05657
R12466 DVSS.n5335 DVSS.n971 4.05657
R12467 DVSS.n5335 DVSS.n969 4.05657
R12468 DVSS.n5339 DVSS.n969 4.05657
R12469 DVSS.n5339 DVSS.n967 4.05657
R12470 DVSS.n5344 DVSS.n967 4.05657
R12471 DVSS.n5344 DVSS.n965 4.05657
R12472 DVSS.n5348 DVSS.n965 4.05657
R12473 DVSS.n5349 DVSS.n5348 4.05657
R12474 DVSS.n3939 DVSS.n3938 3.8345
R12475 DVSS.n3755 DVSS.n3754 3.7805
R12476 DVSS.n3756 DVSS.n3755 3.77031
R12477 DVSS.n4962 DVSS.n1164 3.68022
R12478 DVSS.n3581 DVSS.n1648 3.3741
R12479 DVSS.n3607 DVSS 3.20629
R12480 DVSS.n1732 DVSS 3.18489
R12481 DVSS.n4468 DVSS.t176 3.17811
R12482 DVSS.n4474 DVSS.t57 3.17811
R12483 DVSS.n1657 DVSS.t198 3.17811
R12484 DVSS.n1671 DVSS.t7 3.17811
R12485 DVSS.n1689 DVSS.t129 3.17811
R12486 DVSS.n3763 DVSS.t61 3.17811
R12487 DVSS.n1589 DVSS.t133 3.17811
R12488 DVSS.n3856 DVSS.t147 3.17811
R12489 DVSS.n1578 DVSS.t180 3.17811
R12490 DVSS.n1581 DVSS.t125 3.17811
R12491 DVSS.n4446 DVSS.t181 3.126
R12492 DVSS.n3975 DVSS.n1494 3.02469
R12493 DVSS.n2647 DVSS.n2420 2.95295
R12494 DVSS.n4453 DVSS.n1301 2.90887
R12495 DVSS.n1488 DVSS.n1487 2.81187
R12496 DVSS.n4974 DVSS.n4973 2.81187
R12497 DVSS.n4951 DVSS.n4950 2.81187
R12498 DVSS.n3745 DVSS.n3744 2.75988
R12499 DVSS.n5350 DVSS.n5349 2.6005
R12500 DVSS.n5348 DVSS.n964 2.6005
R12501 DVSS.n5348 DVSS.n5347 2.6005
R12502 DVSS.n5342 DVSS.n965 2.6005
R12503 DVSS.n5346 DVSS.n965 2.6005
R12504 DVSS.n5344 DVSS.n5343 2.6005
R12505 DVSS.n5345 DVSS.n5344 2.6005
R12506 DVSS.n5341 DVSS.n967 2.6005
R12507 DVSS.n967 DVSS.n966 2.6005
R12508 DVSS.n5340 DVSS.n5339 2.6005
R12509 DVSS.n5339 DVSS.n5338 2.6005
R12510 DVSS.n969 DVSS.n968 2.6005
R12511 DVSS.n5337 DVSS.n969 2.6005
R12512 DVSS.n5335 DVSS.n5334 2.6005
R12513 DVSS.n5336 DVSS.n5335 2.6005
R12514 DVSS.n5333 DVSS.n971 2.6005
R12515 DVSS.n971 DVSS.n970 2.6005
R12516 DVSS.n5332 DVSS.n5331 2.6005
R12517 DVSS.n5331 DVSS.n5330 2.6005
R12518 DVSS.n973 DVSS.n972 2.6005
R12519 DVSS.n5329 DVSS.n973 2.6005
R12520 DVSS.n5327 DVSS.n5326 2.6005
R12521 DVSS.n5328 DVSS.n5327 2.6005
R12522 DVSS.n5325 DVSS.n975 2.6005
R12523 DVSS.n975 DVSS.n974 2.6005
R12524 DVSS.n5324 DVSS.n5323 2.6005
R12525 DVSS.n5323 DVSS.n5322 2.6005
R12526 DVSS.n977 DVSS.n976 2.6005
R12527 DVSS.n5321 DVSS.n977 2.6005
R12528 DVSS.n5319 DVSS.n5318 2.6005
R12529 DVSS.n5320 DVSS.n5319 2.6005
R12530 DVSS.n5317 DVSS.n979 2.6005
R12531 DVSS.n979 DVSS.n978 2.6005
R12532 DVSS.n5316 DVSS.n5315 2.6005
R12533 DVSS.n5315 DVSS.n5314 2.6005
R12534 DVSS.n981 DVSS.n980 2.6005
R12535 DVSS.n5313 DVSS.n981 2.6005
R12536 DVSS.n5311 DVSS.n5310 2.6005
R12537 DVSS.n5312 DVSS.n5311 2.6005
R12538 DVSS.n5309 DVSS.n983 2.6005
R12539 DVSS.n983 DVSS.n982 2.6005
R12540 DVSS.n5308 DVSS.n5307 2.6005
R12541 DVSS.n5307 DVSS.n5306 2.6005
R12542 DVSS.n985 DVSS.n984 2.6005
R12543 DVSS.n5305 DVSS.n985 2.6005
R12544 DVSS.n5303 DVSS.n5302 2.6005
R12545 DVSS.n5304 DVSS.n5303 2.6005
R12546 DVSS.n5301 DVSS.n987 2.6005
R12547 DVSS.n987 DVSS.n986 2.6005
R12548 DVSS.n5300 DVSS.n5299 2.6005
R12549 DVSS.n5299 DVSS.n5298 2.6005
R12550 DVSS.n989 DVSS.n988 2.6005
R12551 DVSS.n5297 DVSS.n989 2.6005
R12552 DVSS.n5295 DVSS.n5294 2.6005
R12553 DVSS.n5296 DVSS.n5295 2.6005
R12554 DVSS.n5293 DVSS.n991 2.6005
R12555 DVSS.n991 DVSS.n990 2.6005
R12556 DVSS.n5292 DVSS.n5291 2.6005
R12557 DVSS.n5291 DVSS.n5290 2.6005
R12558 DVSS.n993 DVSS.n992 2.6005
R12559 DVSS.n5289 DVSS.n993 2.6005
R12560 DVSS.n5287 DVSS.n5286 2.6005
R12561 DVSS.n5288 DVSS.n5287 2.6005
R12562 DVSS.n5285 DVSS.n995 2.6005
R12563 DVSS.n995 DVSS.n994 2.6005
R12564 DVSS.n5284 DVSS.n5283 2.6005
R12565 DVSS.n5283 DVSS.n5282 2.6005
R12566 DVSS.n997 DVSS.n996 2.6005
R12567 DVSS.n5281 DVSS.n997 2.6005
R12568 DVSS.n5279 DVSS.n5278 2.6005
R12569 DVSS.n5280 DVSS.n5279 2.6005
R12570 DVSS.n5277 DVSS.n999 2.6005
R12571 DVSS.n999 DVSS.n998 2.6005
R12572 DVSS.n5276 DVSS.n5275 2.6005
R12573 DVSS.n5275 DVSS.n5274 2.6005
R12574 DVSS.n1001 DVSS.n1000 2.6005
R12575 DVSS.n5273 DVSS.n1001 2.6005
R12576 DVSS.n5271 DVSS.n5270 2.6005
R12577 DVSS.n5272 DVSS.n5271 2.6005
R12578 DVSS.n5269 DVSS.n1003 2.6005
R12579 DVSS.n1003 DVSS.n1002 2.6005
R12580 DVSS.n5268 DVSS.n5267 2.6005
R12581 DVSS.n5267 DVSS.n5266 2.6005
R12582 DVSS.n1005 DVSS.n1004 2.6005
R12583 DVSS.n5265 DVSS.n1005 2.6005
R12584 DVSS.n5263 DVSS.n5262 2.6005
R12585 DVSS.n5264 DVSS.n5263 2.6005
R12586 DVSS.n5261 DVSS.n1007 2.6005
R12587 DVSS.n1007 DVSS.n1006 2.6005
R12588 DVSS.n5260 DVSS.n5259 2.6005
R12589 DVSS.n5259 DVSS.n5258 2.6005
R12590 DVSS.n1009 DVSS.n1008 2.6005
R12591 DVSS.n5257 DVSS.n1009 2.6005
R12592 DVSS.n5255 DVSS.n5254 2.6005
R12593 DVSS.n5256 DVSS.n5255 2.6005
R12594 DVSS.n5253 DVSS.n1011 2.6005
R12595 DVSS.n1011 DVSS.n1010 2.6005
R12596 DVSS.n5252 DVSS.n5251 2.6005
R12597 DVSS.n5251 DVSS.n5250 2.6005
R12598 DVSS.n1013 DVSS.n1012 2.6005
R12599 DVSS.n5249 DVSS.n1013 2.6005
R12600 DVSS.n5247 DVSS.n5246 2.6005
R12601 DVSS.n5248 DVSS.n5247 2.6005
R12602 DVSS.n5245 DVSS.n1015 2.6005
R12603 DVSS.n1015 DVSS.n1014 2.6005
R12604 DVSS.n5244 DVSS.n5243 2.6005
R12605 DVSS.n5243 DVSS.n5242 2.6005
R12606 DVSS.n1017 DVSS.n1016 2.6005
R12607 DVSS.n5241 DVSS.n1017 2.6005
R12608 DVSS.n5239 DVSS.n5238 2.6005
R12609 DVSS.n5240 DVSS.n5239 2.6005
R12610 DVSS.n5237 DVSS.n1019 2.6005
R12611 DVSS.n1019 DVSS.n1018 2.6005
R12612 DVSS.n5236 DVSS.n5235 2.6005
R12613 DVSS.n5235 DVSS.n5234 2.6005
R12614 DVSS.n1021 DVSS.n1020 2.6005
R12615 DVSS.n5233 DVSS.n1021 2.6005
R12616 DVSS.n5229 DVSS.n5228 2.6005
R12617 DVSS.n5228 DVSS.n1022 2.6005
R12618 DVSS.n5227 DVSS.n1025 2.6005
R12619 DVSS.n5227 DVSS.n5226 2.6005
R12620 DVSS.n5221 DVSS.n1026 2.6005
R12621 DVSS.n5225 DVSS.n1026 2.6005
R12622 DVSS.n5223 DVSS.n5222 2.6005
R12623 DVSS.n5224 DVSS.n5223 2.6005
R12624 DVSS.n5220 DVSS.n1028 2.6005
R12625 DVSS.n1028 DVSS.n1027 2.6005
R12626 DVSS.n5219 DVSS.n5218 2.6005
R12627 DVSS.n5218 DVSS.n5217 2.6005
R12628 DVSS.n1030 DVSS.n1029 2.6005
R12629 DVSS.n5216 DVSS.n1030 2.6005
R12630 DVSS.n5214 DVSS.n5213 2.6005
R12631 DVSS.n5215 DVSS.n5214 2.6005
R12632 DVSS.n5212 DVSS.n1032 2.6005
R12633 DVSS.n1032 DVSS.n1031 2.6005
R12634 DVSS.n5211 DVSS.n5210 2.6005
R12635 DVSS.n5210 DVSS.n5209 2.6005
R12636 DVSS.n1034 DVSS.n1033 2.6005
R12637 DVSS.n5208 DVSS.n1034 2.6005
R12638 DVSS.n5206 DVSS.n5205 2.6005
R12639 DVSS.n5207 DVSS.n5206 2.6005
R12640 DVSS.n5204 DVSS.n1036 2.6005
R12641 DVSS.n1036 DVSS.n1035 2.6005
R12642 DVSS.n5203 DVSS.n5202 2.6005
R12643 DVSS.n5202 DVSS.n5201 2.6005
R12644 DVSS.n1038 DVSS.n1037 2.6005
R12645 DVSS.n5200 DVSS.n1038 2.6005
R12646 DVSS.n5198 DVSS.n5197 2.6005
R12647 DVSS.n5199 DVSS.n5198 2.6005
R12648 DVSS.n5196 DVSS.n1040 2.6005
R12649 DVSS.n1040 DVSS.n1039 2.6005
R12650 DVSS.n5195 DVSS.n5194 2.6005
R12651 DVSS.n5194 DVSS.n5193 2.6005
R12652 DVSS.n1042 DVSS.n1041 2.6005
R12653 DVSS.n5192 DVSS.n1042 2.6005
R12654 DVSS.n5190 DVSS.n5189 2.6005
R12655 DVSS.n5191 DVSS.n5190 2.6005
R12656 DVSS.n5188 DVSS.n1044 2.6005
R12657 DVSS.n1044 DVSS.n1043 2.6005
R12658 DVSS.n5187 DVSS.n5186 2.6005
R12659 DVSS.n5186 DVSS.n5185 2.6005
R12660 DVSS.n1046 DVSS.n1045 2.6005
R12661 DVSS.n5184 DVSS.n1046 2.6005
R12662 DVSS.n5182 DVSS.n5181 2.6005
R12663 DVSS.n5183 DVSS.n5182 2.6005
R12664 DVSS.n5180 DVSS.n1048 2.6005
R12665 DVSS.n1048 DVSS.n1047 2.6005
R12666 DVSS.n5179 DVSS.n5178 2.6005
R12667 DVSS.n5178 DVSS.n5177 2.6005
R12668 DVSS.n1050 DVSS.n1049 2.6005
R12669 DVSS.n5176 DVSS.n1050 2.6005
R12670 DVSS.n5174 DVSS.n5173 2.6005
R12671 DVSS.n5175 DVSS.n5174 2.6005
R12672 DVSS.n5172 DVSS.n1052 2.6005
R12673 DVSS.n1052 DVSS.n1051 2.6005
R12674 DVSS.n5171 DVSS.n5170 2.6005
R12675 DVSS.n5170 DVSS.n5169 2.6005
R12676 DVSS.n1054 DVSS.n1053 2.6005
R12677 DVSS.n5168 DVSS.n1054 2.6005
R12678 DVSS.n5166 DVSS.n5165 2.6005
R12679 DVSS.n5167 DVSS.n5166 2.6005
R12680 DVSS.n5164 DVSS.n1056 2.6005
R12681 DVSS.n1056 DVSS.n1055 2.6005
R12682 DVSS.n5163 DVSS.n5162 2.6005
R12683 DVSS.n5162 DVSS.n5161 2.6005
R12684 DVSS.n1058 DVSS.n1057 2.6005
R12685 DVSS.n5160 DVSS.n1058 2.6005
R12686 DVSS.n5158 DVSS.n5157 2.6005
R12687 DVSS.n5159 DVSS.n5158 2.6005
R12688 DVSS.n5156 DVSS.n1060 2.6005
R12689 DVSS.n1060 DVSS.n1059 2.6005
R12690 DVSS.n5155 DVSS.n5154 2.6005
R12691 DVSS.n5154 DVSS.n5153 2.6005
R12692 DVSS.n1062 DVSS.n1061 2.6005
R12693 DVSS.n5152 DVSS.n1062 2.6005
R12694 DVSS.n5150 DVSS.n5149 2.6005
R12695 DVSS.n5151 DVSS.n5150 2.6005
R12696 DVSS.n5148 DVSS.n1064 2.6005
R12697 DVSS.n1064 DVSS.n1063 2.6005
R12698 DVSS.n5147 DVSS.n5146 2.6005
R12699 DVSS.n5146 DVSS.n5145 2.6005
R12700 DVSS.n1066 DVSS.n1065 2.6005
R12701 DVSS.n5144 DVSS.n1066 2.6005
R12702 DVSS.n5142 DVSS.n5141 2.6005
R12703 DVSS.n5143 DVSS.n5142 2.6005
R12704 DVSS.n5140 DVSS.n1068 2.6005
R12705 DVSS.n1068 DVSS.n1067 2.6005
R12706 DVSS.n5139 DVSS.n5138 2.6005
R12707 DVSS.n5138 DVSS.n5137 2.6005
R12708 DVSS.n1070 DVSS.n1069 2.6005
R12709 DVSS.n5136 DVSS.n1070 2.6005
R12710 DVSS.n5134 DVSS.n5133 2.6005
R12711 DVSS.n5135 DVSS.n5134 2.6005
R12712 DVSS.n5132 DVSS.n1072 2.6005
R12713 DVSS.n1072 DVSS.n1071 2.6005
R12714 DVSS.n5131 DVSS.n5130 2.6005
R12715 DVSS.n5130 DVSS.n5129 2.6005
R12716 DVSS.n1074 DVSS.n1073 2.6005
R12717 DVSS.n5128 DVSS.n1074 2.6005
R12718 DVSS.n5126 DVSS.n5125 2.6005
R12719 DVSS.n5127 DVSS.n5126 2.6005
R12720 DVSS.n5124 DVSS.n1076 2.6005
R12721 DVSS.n1076 DVSS.n1075 2.6005
R12722 DVSS.n5123 DVSS.n5122 2.6005
R12723 DVSS.n5122 DVSS.n5121 2.6005
R12724 DVSS.n1078 DVSS.n1077 2.6005
R12725 DVSS.n5120 DVSS.n1078 2.6005
R12726 DVSS.n5118 DVSS.n5117 2.6005
R12727 DVSS.n5119 DVSS.n5118 2.6005
R12728 DVSS.n5116 DVSS.n1080 2.6005
R12729 DVSS.n1080 DVSS.n1079 2.6005
R12730 DVSS.n5115 DVSS.n5114 2.6005
R12731 DVSS.n3614 DVSS.n3613 2.49974
R12732 DVSS.n3613 DVSS.n3610 2.49796
R12733 DVSS.n4936 DVSS.n4935 2.43717
R12734 DVSS.n3647 DVSS.n1714 2.41753
R12735 DVSS.n3647 DVSS.n1713 2.41753
R12736 DVSS.n3647 DVSS.n1712 2.41753
R12737 DVSS.n3647 DVSS.n1711 2.41753
R12738 DVSS.n3647 DVSS.n1710 2.41753
R12739 DVSS.n3624 DVSS.n3601 2.41753
R12740 DVSS.n3624 DVSS.n3600 2.41753
R12741 DVSS.n3624 DVSS.n3599 2.41753
R12742 DVSS.n3624 DVSS.n3598 2.41753
R12743 DVSS.n3625 DVSS.n3624 2.41753
R12744 DVSS.n3624 DVSS.n1720 2.41753
R12745 DVSS.n3645 DVSS.n3593 2.41753
R12746 DVSS.n4409 DVSS.n4377 2.41274
R12747 DVSS.n4409 DVSS.n4408 2.41274
R12748 DVSS.n4463 DVSS.n4462 2.41274
R12749 DVSS.n4462 DVSS.n4461 2.41274
R12750 DVSS.n3938 DVSS.n1519 2.311
R12751 DVSS.n3611 DVSS 2.30994
R12752 DVSS.n3609 DVSS 2.30994
R12753 DVSS.t107 DVSS.n2229 2.29246
R12754 DVSS.n1824 DVSS.n1821 2.2728
R12755 DVSS.n4966 DVSS.n4965 2.25682
R12756 DVSS.n4457 DVSS.n4456 2.25682
R12757 DVSS.n4448 DVSS.n1302 2.25682
R12758 DVSS.n4957 DVSS.n4955 2.25682
R12759 DVSS.n1466 DVSS.n1301 2.25392
R12760 DVSS.n3613 DVSS.n3612 2.25346
R12761 DVSS.n1962 DVSS.n1942 2.2505
R12762 DVSS.n2137 DVSS.n2136 2.2505
R12763 DVSS.n1937 DVSS.n1931 2.2505
R12764 DVSS.n1936 DVSS.n1926 2.2505
R12765 DVSS.n1777 DVSS.n1763 2.2505
R12766 DVSS.n1870 DVSS.n1773 2.2505
R12767 DVSS.n2188 DVSS.n2187 2.2505
R12768 DVSS.n1779 DVSS.n1770 2.2505
R12769 DVSS.n2090 DVSS.n2085 2.2505
R12770 DVSS.n2093 DVSS.n1953 2.2505
R12771 DVSS.n2125 DVSS.n2124 2.2505
R12772 DVSS.n1984 DVSS.n1945 2.2505
R12773 DVSS.n2110 DVSS.n2099 2.2505
R12774 DVSS.n2102 DVSS.n1808 2.2505
R12775 DVSS.n2104 DVSS.n2103 2.2505
R12776 DVSS.n2106 DVSS.n2100 2.2505
R12777 DVSS.n2109 DVSS.n2108 2.2505
R12778 DVSS.n1835 DVSS.n1834 2.2505
R12779 DVSS.n1833 DVSS.n1832 2.2505
R12780 DVSS.n1830 DVSS.n1829 2.2505
R12781 DVSS.n1828 DVSS.n1827 2.2505
R12782 DVSS.n1826 DVSS.n1820 2.2505
R12783 DVSS.n2097 DVSS.n2096 2.2505
R12784 DVSS.n2095 DVSS.n2094 2.2505
R12785 DVSS.n2092 DVSS.n2091 2.2505
R12786 DVSS.n1951 DVSS.n1950 2.2505
R12787 DVSS.n2127 DVSS.n2126 2.2505
R12788 DVSS.n2129 DVSS.n2128 2.2505
R12789 DVSS.n2132 DVSS.n2131 2.2505
R12790 DVSS.n2133 DVSS.n1934 2.2505
R12791 DVSS.n2135 DVSS.n2134 2.2505
R12792 DVSS.n1940 DVSS.n1933 2.2505
R12793 DVSS.n1939 DVSS.n1938 2.2505
R12794 DVSS.n1935 DVSS.n1801 2.2505
R12795 DVSS.n2184 DVSS.n2183 2.2505
R12796 DVSS.n2186 DVSS.n2185 2.2505
R12797 DVSS.n1782 DVSS.n1772 2.2505
R12798 DVSS.n1781 DVSS.n1780 2.2505
R12799 DVSS.n1778 DVSS.n1776 2.2505
R12800 DVSS.n1775 DVSS.n1753 2.2505
R12801 DVSS.n2202 DVSS.n2201 2.2505
R12802 DVSS.n1748 DVSS.n1746 2.2505
R12803 DVSS.n2209 DVSS.n2208 2.2505
R12804 DVSS.n1892 DVSS.n1747 2.2505
R12805 DVSS.n2211 DVSS.n2210 2.2505
R12806 DVSS.n1824 DVSS.n1823 2.2505
R12807 DVSS.n3938 DVSS.n3937 2.2505
R12808 DVSS.n294 DVSS.n265 2.2505
R12809 DVSS.n293 DVSS.n292 2.2505
R12810 DVSS.n291 DVSS.n266 2.2505
R12811 DVSS.n290 DVSS.n289 2.2505
R12812 DVSS.n288 DVSS.n267 2.2505
R12813 DVSS.n287 DVSS.n286 2.2505
R12814 DVSS.n285 DVSS.n268 2.2505
R12815 DVSS.n284 DVSS.n283 2.2505
R12816 DVSS.n282 DVSS.n269 2.2505
R12817 DVSS.n281 DVSS.n280 2.2505
R12818 DVSS.n279 DVSS.n270 2.2505
R12819 DVSS.n278 DVSS.n277 2.2505
R12820 DVSS.n274 DVSS.n271 2.2505
R12821 DVSS.n273 DVSS.n272 2.2505
R12822 DVSS.n429 DVSS.n428 2.2505
R12823 DVSS.n430 DVSS.n240 2.2505
R12824 DVSS.n432 DVSS.n431 2.2505
R12825 DVSS.n433 DVSS.n239 2.2505
R12826 DVSS.n435 DVSS.n434 2.2505
R12827 DVSS.n436 DVSS.n238 2.2505
R12828 DVSS.n438 DVSS.n437 2.2505
R12829 DVSS.n439 DVSS.n237 2.2505
R12830 DVSS.n441 DVSS.n440 2.2505
R12831 DVSS.n442 DVSS.n236 2.2505
R12832 DVSS.n444 DVSS.n443 2.2505
R12833 DVSS.n445 DVSS.n235 2.2505
R12834 DVSS.n447 DVSS.n446 2.2505
R12835 DVSS.n448 DVSS.n234 2.2505
R12836 DVSS.n450 DVSS.n449 2.2505
R12837 DVSS.n451 DVSS.n233 2.2505
R12838 DVSS.n453 DVSS.n452 2.2505
R12839 DVSS.n454 DVSS.n232 2.2505
R12840 DVSS.n456 DVSS.n455 2.2505
R12841 DVSS.n457 DVSS.n231 2.2505
R12842 DVSS.n459 DVSS.n458 2.2505
R12843 DVSS.n460 DVSS.n230 2.2505
R12844 DVSS.n462 DVSS.n461 2.2505
R12845 DVSS.n307 DVSS.n261 2.2505
R12846 DVSS.n309 DVSS.n308 2.2505
R12847 DVSS.n306 DVSS.n259 2.2505
R12848 DVSS.n305 DVSS.n304 2.2505
R12849 DVSS.n303 DVSS.n262 2.2505
R12850 DVSS.n302 DVSS.n301 2.2505
R12851 DVSS.n300 DVSS.n263 2.2505
R12852 DVSS.n299 DVSS.n298 2.2505
R12853 DVSS.n297 DVSS.n264 2.2505
R12854 DVSS.n296 DVSS.n295 2.2505
R12855 DVSS.n800 DVSS.n754 2.2505
R12856 DVSS.n799 DVSS.n798 2.2505
R12857 DVSS.n797 DVSS.n755 2.2505
R12858 DVSS.n796 DVSS.n795 2.2505
R12859 DVSS.n794 DVSS.n756 2.2505
R12860 DVSS.n793 DVSS.n792 2.2505
R12861 DVSS.n791 DVSS.n757 2.2505
R12862 DVSS.n790 DVSS.n789 2.2505
R12863 DVSS.n787 DVSS.n786 2.2505
R12864 DVSS.n785 DVSS.n759 2.2505
R12865 DVSS.n784 DVSS.n783 2.2505
R12866 DVSS.n782 DVSS.n760 2.2505
R12867 DVSS.n781 DVSS.n780 2.2505
R12868 DVSS.n779 DVSS.n761 2.2505
R12869 DVSS.n778 DVSS.n777 2.2505
R12870 DVSS.n776 DVSS.n762 2.2505
R12871 DVSS.n775 DVSS.n774 2.2505
R12872 DVSS.n773 DVSS.n763 2.2505
R12873 DVSS.n772 DVSS.n771 2.2505
R12874 DVSS.n770 DVSS.n764 2.2505
R12875 DVSS.n769 DVSS.n768 2.2505
R12876 DVSS.n767 DVSS.n766 2.2505
R12877 DVSS.n5730 DVSS.n5729 2.2505
R12878 DVSS.n5728 DVSS.n56 2.2505
R12879 DVSS.n72 DVSS.n58 2.2505
R12880 DVSS.n74 DVSS.n73 2.2505
R12881 DVSS.n75 DVSS.n71 2.2505
R12882 DVSS.n77 DVSS.n76 2.2505
R12883 DVSS.n78 DVSS.n70 2.2505
R12884 DVSS.n80 DVSS.n79 2.2505
R12885 DVSS.n81 DVSS.n69 2.2505
R12886 DVSS.n83 DVSS.n82 2.2505
R12887 DVSS.n84 DVSS.n68 2.2505
R12888 DVSS.n86 DVSS.n85 2.2505
R12889 DVSS.n87 DVSS.n67 2.2505
R12890 DVSS.n89 DVSS.n88 2.2505
R12891 DVSS.n90 DVSS.n66 2.2505
R12892 DVSS.n92 DVSS.n91 2.2505
R12893 DVSS.n93 DVSS.n65 2.2505
R12894 DVSS.n95 DVSS.n94 2.2505
R12895 DVSS.n96 DVSS.n64 2.2505
R12896 DVSS.n98 DVSS.n97 2.2505
R12897 DVSS.n99 DVSS.n63 2.2505
R12898 DVSS.n101 DVSS.n100 2.2505
R12899 DVSS.n5719 DVSS.n62 2.2505
R12900 DVSS.n5721 DVSS.n5720 2.2505
R12901 DVSS.n788 DVSS.n758 2.2505
R12902 DVSS.n4821 DVSS.n4809 2.24683
R12903 DVSS.n4815 DVSS.n4811 2.24683
R12904 DVSS.n4538 DVSS.n4526 2.24683
R12905 DVSS.n5553 DVSS.n852 2.24648
R12906 DVSS.n5553 DVSS.n851 2.24648
R12907 DVSS.n5553 DVSS.n850 2.24648
R12908 DVSS.n5553 DVSS.n849 2.24648
R12909 DVSS.n855 DVSS.n848 2.24648
R12910 DVSS.n855 DVSS.n853 2.24648
R12911 DVSS.n1191 DVSS.n855 2.24648
R12912 DVSS.n855 DVSS.n854 2.24648
R12913 DVSS.n1856 DVSS.n1855 2.24442
R12914 DVSS.n1858 DVSS.n1857 2.24442
R12915 DVSS.n4817 DVSS.n4816 2.24405
R12916 DVSS.n4814 DVSS.n4813 2.24405
R12917 DVSS.n4818 DVSS.n4817 2.24405
R12918 DVSS.n4533 DVSS.n4529 2.24405
R12919 DVSS.n4537 DVSS.n4530 2.24405
R12920 DVSS.n4531 DVSS.n4529 2.24405
R12921 DVSS.n1978 DVSS.n1977 2.24386
R12922 DVSS.n1976 DVSS.n1975 2.24386
R12923 DVSS.n1975 DVSS.n1974 2.24386
R12924 DVSS.n1911 DVSS.n1882 2.24386
R12925 DVSS.n1910 DVSS.n1909 2.24386
R12926 DVSS.n1909 DVSS.n1881 2.24386
R12927 DVSS.n4872 DVSS.n4834 2.24304
R12928 DVSS.n4830 DVSS.n4829 2.24304
R12929 DVSS.n4872 DVSS.n4833 2.24304
R12930 DVSS.n4830 DVSS.n4828 2.24304
R12931 DVSS.n4872 DVSS.n4832 2.24304
R12932 DVSS.n4830 DVSS.n4827 2.24304
R12933 DVSS.n4873 DVSS.n4872 2.24304
R12934 DVSS.n4830 DVSS.n4826 2.24304
R12935 DVSS.n4544 DVSS.n4524 2.24304
R12936 DVSS.n4522 DVSS.n4509 2.24304
R12937 DVSS.n4544 DVSS.n4520 2.24304
R12938 DVSS.n4518 DVSS.n4509 2.24304
R12939 DVSS.n4544 DVSS.n4516 2.24304
R12940 DVSS.n4514 DVSS.n4509 2.24304
R12941 DVSS.n4544 DVSS.n4512 2.24304
R12942 DVSS.n4542 DVSS.n4509 2.24304
R12943 DVSS.n3840 DVSS.n1632 2.24304
R12944 DVSS.n1630 DVSS.n1625 2.24304
R12945 DVSS.n3830 DVSS.n1620 2.24304
R12946 DVSS.n3829 DVSS.n1625 2.24304
R12947 DVSS.n3833 DVSS.n1620 2.24304
R12948 DVSS.n3832 DVSS.n1625 2.24304
R12949 DVSS.n3836 DVSS.n1620 2.24304
R12950 DVSS.n3835 DVSS.n1625 2.24304
R12951 DVSS.n3838 DVSS.n1620 2.24304
R12952 DVSS.n2407 DVSS.n2275 2.24304
R12953 DVSS.n2404 DVSS.n2278 2.24304
R12954 DVSS.n2405 DVSS.n2275 2.24304
R12955 DVSS.n2419 DVSS.n2411 2.24304
R12956 DVSS.n2409 DVSS.n2278 2.24304
R12957 DVSS.n2419 DVSS.n2415 2.24304
R12958 DVSS.n2413 DVSS.n2278 2.24304
R12959 DVSS.n2417 DVSS.n2278 2.24304
R12960 DVSS.n2648 DVSS.n2270 2.24304
R12961 DVSS.n2643 DVSS.n2640 2.24304
R12962 DVSS.n2648 DVSS.n2271 2.24304
R12963 DVSS.n2643 DVSS.n2641 2.24304
R12964 DVSS.n2648 DVSS.n2272 2.24304
R12965 DVSS.n2643 DVSS.n2642 2.24304
R12966 DVSS.n2648 DVSS.n2273 2.24304
R12967 DVSS.n2644 DVSS.n2643 2.24304
R12968 DVSS.n2643 DVSS.n2274 2.24304
R12969 DVSS.n1948 DVSS.n1944 2.24011
R12970 DVSS.n1946 DVSS.n1944 2.24011
R12971 DVSS.n2199 DVSS.n1757 2.24011
R12972 DVSS.n2199 DVSS.n1755 2.24011
R12973 DVSS.n2204 DVSS.n1750 2.24011
R12974 DVSS.n2206 DVSS.n1750 2.24011
R12975 DVSS.n1785 DVSS.n1784 2.24011
R12976 DVSS.n2168 DVSS.n1800 2.24011
R12977 DVSS.n1947 DVSS.n1943 2.24011
R12978 DVSS.n1756 DVSS.n1754 2.24011
R12979 DVSS.n2205 DVSS.n1749 2.24011
R12980 DVSS.n2147 DVSS.n2145 2.23777
R12981 DVSS.n2148 DVSS.n1797 2.23777
R12982 DVSS.n2149 DVSS.n2145 2.23777
R12983 DVSS.n1875 DVSS.n1874 2.23777
R12984 DVSS.n1877 DVSS.n1876 2.23777
R12985 DVSS.n1874 DVSS.n1869 2.23777
R12986 DVSS.n5812 DVSS.n25 2.23644
R12987 DVSS.n24 DVSS.n6 2.23644
R12988 DVSS.n5812 DVSS.n23 2.23644
R12989 DVSS.n22 DVSS.n6 2.23644
R12990 DVSS.n5812 DVSS.n21 2.23644
R12991 DVSS.n20 DVSS.n6 2.23644
R12992 DVSS.n5812 DVSS.n19 2.23644
R12993 DVSS.n18 DVSS.n6 2.23644
R12994 DVSS.n5812 DVSS.n17 2.23644
R12995 DVSS.n16 DVSS.n6 2.23644
R12996 DVSS.n5812 DVSS.n15 2.23644
R12997 DVSS.n14 DVSS.n6 2.23644
R12998 DVSS.n5812 DVSS.n13 2.23644
R12999 DVSS.n12 DVSS.n6 2.23644
R13000 DVSS.n5812 DVSS.n11 2.23644
R13001 DVSS.n10 DVSS.n6 2.23644
R13002 DVSS.n5812 DVSS.n9 2.23644
R13003 DVSS.n8 DVSS.n6 2.23644
R13004 DVSS.n5812 DVSS.n7 2.23644
R13005 DVSS.n5810 DVSS.n6 2.23644
R13006 DVSS.n5560 DVSS.n5556 2.23644
R13007 DVSS.n847 DVSS.n829 2.23644
R13008 DVSS.n5560 DVSS.n846 2.23644
R13009 DVSS.n845 DVSS.n829 2.23644
R13010 DVSS.n5560 DVSS.n844 2.23644
R13011 DVSS.n843 DVSS.n829 2.23644
R13012 DVSS.n5560 DVSS.n842 2.23644
R13013 DVSS.n841 DVSS.n829 2.23644
R13014 DVSS.n5560 DVSS.n840 2.23644
R13015 DVSS.n839 DVSS.n829 2.23644
R13016 DVSS.n5560 DVSS.n838 2.23644
R13017 DVSS.n837 DVSS.n829 2.23644
R13018 DVSS.n5560 DVSS.n836 2.23644
R13019 DVSS.n835 DVSS.n829 2.23644
R13020 DVSS.n5560 DVSS.n834 2.23644
R13021 DVSS.n833 DVSS.n829 2.23644
R13022 DVSS.n5560 DVSS.n832 2.23644
R13023 DVSS.n831 DVSS.n829 2.23644
R13024 DVSS.n5560 DVSS.n830 2.23644
R13025 DVSS.n5558 DVSS.n829 2.23644
R13026 DVSS.n3612 DVSS.n3611 2.18437
R13027 DVSS.n3610 DVSS.n3609 2.18437
R13028 DVSS.n3959 DVSS.n3958 2.16228
R13029 DVSS.n5355 DVSS.n5354 2.15282
R13030 DVSS.n3905 DVSS.n3904 2.12226
R13031 DVSS.n3793 DVSS.n1654 2.10421
R13032 DVSS.n2242 DVSS.n2241 2.10097
R13033 DVSS.n4470 DVSS.n4469 2.08611
R13034 DVSS.n1692 DVSS.n1691 2.08611
R13035 DVSS.n1656 DVSS.n1655 2.08611
R13036 DVSS.n1576 DVSS.n1575 2.08611
R13037 DVSS.n1584 DVSS.n1583 2.08611
R13038 DVSS.n1480 DVSS.n1479 2.07167
R13039 DVSS.n3583 DVSS.n3581 2.04166
R13040 DVSS.n3977 DVSS.n3976 2.01663
R13041 DVSS.t66 DVSS.n4457 2.01372
R13042 DVSS.n3769 DVSS.n1688 1.96906
R13043 DVSS.n1451 DVSS.n1447 1.94426
R13044 DVSS.n3577 DVSS.n2246 1.94426
R13045 DVSS.n2233 DVSS.n2232 1.91475
R13046 DVSS.n2234 DVSS.n1518 1.91081
R13047 DVSS.n2252 DVSS.n2251 1.89625
R13048 DVSS.n3653 DVSS.n3652 1.87995
R13049 DVSS.n4385 DVSS.n4382 1.81109
R13050 DVSS.n1455 DVSS.n1290 1.81109
R13051 DVSS.n4387 DVSS.n4378 1.81109
R13052 DVSS.n1457 DVSS.n1292 1.81109
R13053 DVSS.n4478 DVSS.n4477 1.80682
R13054 VSS DVSS.n3945 1.7864
R13055 DVSS.n3942 VSS 1.7864
R13056 DVSS.n1279 DVSS.n1275 1.73383
R13057 DVSS.n4472 DVSS.n1275 1.73383
R13058 DVSS.n4397 DVSS.n1171 1.73383
R13059 DVSS.n1171 DVSS.n1170 1.73383
R13060 DVSS.n1461 DVSS.n1296 1.73383
R13061 DVSS.n1303 DVSS.n1296 1.73383
R13062 DVSS.n4435 DVSS.n4434 1.73383
R13063 DVSS.n4434 DVSS.n4433 1.73383
R13064 DVSS.n5351 DVSS.n5350 1.69455
R13065 DVSS.n5723 DVSS.n5722 1.66284
R13066 DVSS.n4485 DVSS.n4484 1.66212
R13067 DVSS.n5723 DVSS.n60 1.64846
R13068 DVSS.n1489 DVSS.n1488 1.61108
R13069 DVSS.n4974 DVSS.n4969 1.61108
R13070 DVSS.n4952 DVSS.n4951 1.61108
R13071 DVSS.n1510 DVSS.t42 1.5965
R13072 DVSS.n1514 DVSS.t41 1.5965
R13073 DVSS.n3953 DVSS.t47 1.5965
R13074 DVSS.n1507 DVSS.t43 1.5965
R13075 DVSS.n1508 DVSS.t43 1.5965
R13076 DVSS.n1508 DVSS.t41 1.5965
R13077 DVSS.n1505 DVSS.t47 1.5965
R13078 DVSS.n1505 DVSS.t42 1.5965
R13079 DVSS.n3895 DVSS.n3894 1.59033
R13080 DVSS.n3886 DVSS.n1585 1.59033
R13081 DVSS.n3877 DVSS.n1582 1.59033
R13082 DVSS.n1605 DVSS.n1579 1.59033
R13083 DVSS.n1610 DVSS.n1577 1.59033
R13084 DVSS.n3858 DVSS.n3857 1.59033
R13085 DVSS.n1674 DVSS.n1673 1.59033
R13086 DVSS.n3764 DVSS.n1662 1.59033
R13087 DVSS.n1693 DVSS.n1682 1.59033
R13088 DVSS.n2258 DVSS.n1698 1.56129
R13089 DVSS.n3948 DVSS.n1504 1.52301
R13090 DVSS.n3584 DVSS.n3580 1.51243
R13091 DVSS.n4900 DVSS.n4899 1.50734
R13092 DVSS.n4885 DVSS.n4884 1.50734
R13093 DVSS.n4754 DVSS.n4753 1.50734
R13094 DVSS.n4770 DVSS.n4769 1.50734
R13095 DVSS.n1252 DVSS.n1251 1.50734
R13096 DVSS.n4736 DVSS.n4735 1.50734
R13097 DVSS.n4620 DVSS.n4619 1.50734
R13098 DVSS.n4696 DVSS.n4695 1.50734
R13099 DVSS.n4652 DVSS.n4651 1.50734
R13100 DVSS.n4637 DVSS.n4636 1.50734
R13101 DVSS.n4561 DVSS.n4560 1.50734
R13102 DVSS.n4577 DVSS.n4576 1.50734
R13103 DVSS.n2803 DVSS.n2789 1.5055
R13104 DVSS.n3419 DVSS.n3418 1.5055
R13105 DVSS.n2803 DVSS.n2802 1.5055
R13106 DVSS.n3418 DVSS.n3375 1.5055
R13107 DVSS.n4376 DVSS.n1316 1.50326
R13108 DVSS.n1475 DVSS.n1474 1.50326
R13109 DVSS.n4169 DVSS.n1390 1.50157
R13110 DVSS.n4575 DVSS.n4497 1.5005
R13111 DVSS.n4670 DVSS.n4669 1.5005
R13112 DVSS.n4567 DVSS.n4494 1.5005
R13113 DVSS.n4566 DVSS.n4565 1.5005
R13114 DVSS.n4505 DVSS.n4503 1.5005
R13115 DVSS.n4602 DVSS.n4595 1.5005
R13116 DVSS.n4641 DVSS.n4640 1.5005
R13117 DVSS.n4597 DVSS.n4592 1.5005
R13118 DVSS.n4596 DVSS.n4585 1.5005
R13119 DVSS.n4650 DVSS.n4649 1.5005
R13120 DVSS.n1265 DVSS.n1261 1.5005
R13121 DVSS.n4692 DVSS.n4691 1.5005
R13122 DVSS.n4683 DVSS.n4682 1.5005
R13123 DVSS.n1270 DVSS.n1269 1.5005
R13124 DVSS.n4618 DVSS.n4617 1.5005
R13125 DVSS.n1244 DVSS.n1240 1.5005
R13126 DVSS.n4732 DVSS.n4731 1.5005
R13127 DVSS.n4722 DVSS.n4721 1.5005
R13128 DVSS.n1250 DVSS.n1249 1.5005
R13129 DVSS.n4715 DVSS.n4714 1.5005
R13130 DVSS.n4768 DVSS.n1223 1.5005
R13131 DVSS.n4918 DVSS.n4917 1.5005
R13132 DVSS.n4760 DVSS.n1220 1.5005
R13133 DVSS.n4759 DVSS.n4758 1.5005
R13134 DVSS.n1231 DVSS.n1229 1.5005
R13135 DVSS.n4795 DVSS.n4788 1.5005
R13136 DVSS.n4889 DVSS.n4888 1.5005
R13137 DVSS.n4790 DVSS.n4785 1.5005
R13138 DVSS.n4789 DVSS.n4778 1.5005
R13139 DVSS.n4898 DVSS.n4897 1.5005
R13140 DVSS.n1836 DVSS.n1389 1.5005
R13141 DVSS.n1838 DVSS.n1837 1.5005
R13142 DVSS.n1840 DVSS.n1839 1.5005
R13143 DVSS.n1842 DVSS.n1841 1.5005
R13144 DVSS.n1844 DVSS.n1843 1.5005
R13145 DVSS.n1846 DVSS.n1845 1.5005
R13146 DVSS.n1848 DVSS.n1847 1.5005
R13147 DVSS.n1850 DVSS.n1849 1.5005
R13148 DVSS.n1852 DVSS.n1851 1.5005
R13149 DVSS.n3989 DVSS.n3988 1.5005
R13150 DVSS.n3991 DVSS.n3990 1.5005
R13151 DVSS.n3993 DVSS.n3992 1.5005
R13152 DVSS.n3995 DVSS.n3994 1.5005
R13153 DVSS.n3997 DVSS.n3996 1.5005
R13154 DVSS.n3999 DVSS.n3998 1.5005
R13155 DVSS.n4001 DVSS.n4000 1.5005
R13156 DVSS.n4003 DVSS.n4002 1.5005
R13157 DVSS.n1437 DVSS.n1435 1.5005
R13158 DVSS.n3423 DVSS.n3422 1.5005
R13159 DVSS.n3421 DVSS.n3239 1.5005
R13160 DVSS.n3420 DVSS.n3419 1.5005
R13161 DVSS.n3241 DVSS.n3238 1.5005
R13162 DVSS.n3240 DVSS.n3225 1.5005
R13163 DVSS.n3433 DVSS.n3432 1.5005
R13164 DVSS.n3436 DVSS.n3435 1.5005
R13165 DVSS.n3224 DVSS.n3221 1.5005
R13166 DVSS.n3223 DVSS.n3208 1.5005
R13167 DVSS.n3444 DVSS.n3207 1.5005
R13168 DVSS.n3446 DVSS.n3445 1.5005
R13169 DVSS.n3448 DVSS.n3447 1.5005
R13170 DVSS.n3205 DVSS.n3203 1.5005
R13171 DVSS.n3190 DVSS.n3189 1.5005
R13172 DVSS.n3458 DVSS.n3457 1.5005
R13173 DVSS.n3460 DVSS.n3459 1.5005
R13174 DVSS.n3188 DVSS.n3182 1.5005
R13175 DVSS.n3187 DVSS.n3186 1.5005
R13176 DVSS.n3170 DVSS.n3169 1.5005
R13177 DVSS.n3470 DVSS.n3469 1.5005
R13178 DVSS.n3472 DVSS.n3471 1.5005
R13179 DVSS.n3168 DVSS.n3166 1.5005
R13180 DVSS.n3153 DVSS.n3151 1.5005
R13181 DVSS.n3482 DVSS.n3481 1.5005
R13182 DVSS.n3484 DVSS.n3149 1.5005
R13183 DVSS.n3486 DVSS.n3485 1.5005
R13184 DVSS.n3150 DVSS.n3148 1.5005
R13185 DVSS.n3135 DVSS.n3134 1.5005
R13186 DVSS.n3496 DVSS.n3495 1.5005
R13187 DVSS.n3498 DVSS.n3497 1.5005
R13188 DVSS.n3132 DVSS.n3129 1.5005
R13189 DVSS.n3131 DVSS.n3116 1.5005
R13190 DVSS.n3507 DVSS.n3115 1.5005
R13191 DVSS.n3509 DVSS.n3508 1.5005
R13192 DVSS.n3511 DVSS.n3510 1.5005
R13193 DVSS.n3114 DVSS.n3112 1.5005
R13194 DVSS.n3099 DVSS.n3098 1.5005
R13195 DVSS.n3521 DVSS.n3520 1.5005
R13196 DVSS.n3523 DVSS.n3522 1.5005
R13197 DVSS.n3097 DVSS.n3091 1.5005
R13198 DVSS.n3096 DVSS.n3095 1.5005
R13199 DVSS.n3093 DVSS.n3079 1.5005
R13200 DVSS.n3533 DVSS.n3532 1.5005
R13201 DVSS.n3536 DVSS.n3535 1.5005
R13202 DVSS.n3077 DVSS.n3075 1.5005
R13203 DVSS.n2672 DVSS.n2671 1.5005
R13204 DVSS.n3546 DVSS.n3545 1.5005
R13205 DVSS.n3548 DVSS.n3547 1.5005
R13206 DVSS.n2670 DVSS.n2668 1.5005
R13207 DVSS.n3060 DVSS.n3059 1.5005
R13208 DVSS.n3057 DVSS.n2682 1.5005
R13209 DVSS.n3056 DVSS.n3055 1.5005
R13210 DVSS.n2684 DVSS.n2683 1.5005
R13211 DVSS.n3039 DVSS.n3038 1.5005
R13212 DVSS.n3037 DVSS.n3036 1.5005
R13213 DVSS.n3017 DVSS.n2693 1.5005
R13214 DVSS.n3019 DVSS.n3018 1.5005
R13215 DVSS.n3016 DVSS.n2703 1.5005
R13216 DVSS.n3015 DVSS.n3014 1.5005
R13217 DVSS.n2705 DVSS.n2704 1.5005
R13218 DVSS.n2993 DVSS.n2992 1.5005
R13219 DVSS.n2990 DVSS.n2989 1.5005
R13220 DVSS.n2714 DVSS.n2713 1.5005
R13221 DVSS.n2973 DVSS.n2972 1.5005
R13222 DVSS.n2971 DVSS.n2970 1.5005
R13223 DVSS.n2969 DVSS.n2968 1.5005
R13224 DVSS.n2967 DVSS.n2966 1.5005
R13225 DVSS.n2952 DVSS.n2726 1.5005
R13226 DVSS.n2954 DVSS.n2953 1.5005
R13227 DVSS.n2951 DVSS.n2950 1.5005
R13228 DVSS.n2738 DVSS.n2737 1.5005
R13229 DVSS.n2918 DVSS.n2917 1.5005
R13230 DVSS.n2916 DVSS.n2915 1.5005
R13231 DVSS.n2914 DVSS.n2913 1.5005
R13232 DVSS.n2912 DVSS.n2911 1.5005
R13233 DVSS.n2749 DVSS.n2748 1.5005
R13234 DVSS.n2891 DVSS.n2890 1.5005
R13235 DVSS.n2889 DVSS.n2888 1.5005
R13236 DVSS.n2760 DVSS.n2759 1.5005
R13237 DVSS.n2863 DVSS.n2862 1.5005
R13238 DVSS.n2860 DVSS.n2767 1.5005
R13239 DVSS.n2859 DVSS.n2858 1.5005
R13240 DVSS.n2769 DVSS.n2768 1.5005
R13241 DVSS.n2842 DVSS.n2841 1.5005
R13242 DVSS.n2840 DVSS.n2839 1.5005
R13243 DVSS.n2817 DVSS.n2780 1.5005
R13244 DVSS.n2819 DVSS.n2818 1.5005
R13245 DVSS.n2816 DVSS.n2815 1.5005
R13246 DVSS.n2814 DVSS.n2788 1.5005
R13247 DVSS.n2794 DVSS.n2789 1.5005
R13248 DVSS.n3372 DVSS.n3371 1.5005
R13249 DVSS.n3375 DVSS.n1704 1.5005
R13250 DVSS.n2802 DVSS.n2801 1.5005
R13251 DVSS.n2800 DVSS.n2799 1.5005
R13252 DVSS.n2798 DVSS.n2784 1.5005
R13253 DVSS.n2824 DVSS.n2823 1.5005
R13254 DVSS.n2825 DVSS.n2782 1.5005
R13255 DVSS.n2834 DVSS.n2833 1.5005
R13256 DVSS.n2832 DVSS.n2831 1.5005
R13257 DVSS.n2830 DVSS.n2829 1.5005
R13258 DVSS.n2828 DVSS.n2827 1.5005
R13259 DVSS.n2765 DVSS.n2764 1.5005
R13260 DVSS.n2868 DVSS.n2867 1.5005
R13261 DVSS.n2870 DVSS.n2762 1.5005
R13262 DVSS.n2883 DVSS.n2882 1.5005
R13263 DVSS.n2881 DVSS.n2880 1.5005
R13264 DVSS.n2879 DVSS.n2878 1.5005
R13265 DVSS.n2877 DVSS.n2876 1.5005
R13266 DVSS.n2874 DVSS.n2872 1.5005
R13267 DVSS.n2873 DVSS.n2742 1.5005
R13268 DVSS.n2923 DVSS.n2922 1.5005
R13269 DVSS.n2924 DVSS.n2740 1.5005
R13270 DVSS.n2945 DVSS.n2944 1.5005
R13271 DVSS.n2943 DVSS.n2942 1.5005
R13272 DVSS.n2941 DVSS.n2940 1.5005
R13273 DVSS.n2938 DVSS.n2937 1.5005
R13274 DVSS.n2935 DVSS.n2925 1.5005
R13275 DVSS.n2934 DVSS.n2933 1.5005
R13276 DVSS.n2932 DVSS.n2931 1.5005
R13277 DVSS.n2930 DVSS.n2929 1.5005
R13278 DVSS.n2928 DVSS.n2927 1.5005
R13279 DVSS.n2998 DVSS.n2997 1.5005
R13280 DVSS.n2999 DVSS.n2707 1.5005
R13281 DVSS.n3008 DVSS.n3007 1.5005
R13282 DVSS.n3006 DVSS.n3005 1.5005
R13283 DVSS.n3004 DVSS.n3003 1.5005
R13284 DVSS.n3002 DVSS.n3001 1.5005
R13285 DVSS.n2695 DVSS.n2688 1.5005
R13286 DVSS.n3044 DVSS.n3043 1.5005
R13287 DVSS.n3045 DVSS.n2686 1.5005
R13288 DVSS.n3049 DVSS.n3048 1.5005
R13289 DVSS.n3047 DVSS.n3046 1.5005
R13290 DVSS.n2664 DVSS.n2662 1.5005
R13291 DVSS.n3553 DVSS.n3552 1.5005
R13292 DVSS.n2665 DVSS.n2663 1.5005
R13293 DVSS.n3257 DVSS.n3256 1.5005
R13294 DVSS.n3259 DVSS.n3258 1.5005
R13295 DVSS.n3262 DVSS.n3261 1.5005
R13296 DVSS.n3264 DVSS.n3263 1.5005
R13297 DVSS.n3268 DVSS.n3267 1.5005
R13298 DVSS.n3270 DVSS.n3269 1.5005
R13299 DVSS.n3271 DVSS.n3252 1.5005
R13300 DVSS.n3274 DVSS.n3273 1.5005
R13301 DVSS.n3276 DVSS.n3275 1.5005
R13302 DVSS.n3280 DVSS.n3279 1.5005
R13303 DVSS.n3282 DVSS.n3281 1.5005
R13304 DVSS.n3285 DVSS.n3284 1.5005
R13305 DVSS.n3287 DVSS.n3286 1.5005
R13306 DVSS.n3290 DVSS.n3249 1.5005
R13307 DVSS.n3292 DVSS.n3291 1.5005
R13308 DVSS.n3294 DVSS.n3293 1.5005
R13309 DVSS.n3297 DVSS.n3296 1.5005
R13310 DVSS.n3300 DVSS.n3299 1.5005
R13311 DVSS.n3304 DVSS.n3303 1.5005
R13312 DVSS.n3306 DVSS.n3305 1.5005
R13313 DVSS.n3309 DVSS.n3308 1.5005
R13314 DVSS.n3310 DVSS.n3248 1.5005
R13315 DVSS.n3312 DVSS.n3311 1.5005
R13316 DVSS.n3316 DVSS.n3315 1.5005
R13317 DVSS.n3318 DVSS.n3317 1.5005
R13318 DVSS.n3321 DVSS.n3320 1.5005
R13319 DVSS.n3323 DVSS.n3322 1.5005
R13320 DVSS.n3327 DVSS.n3326 1.5005
R13321 DVSS.n3329 DVSS.n3328 1.5005
R13322 DVSS.n3332 DVSS.n3331 1.5005
R13323 DVSS.n3334 DVSS.n3333 1.5005
R13324 DVSS.n3336 DVSS.n3335 1.5005
R13325 DVSS.n3340 DVSS.n3339 1.5005
R13326 DVSS.n3342 DVSS.n3341 1.5005
R13327 DVSS.n3345 DVSS.n3344 1.5005
R13328 DVSS.n3348 DVSS.n3347 1.5005
R13329 DVSS.n3352 DVSS.n3351 1.5005
R13330 DVSS.n3353 DVSS.n3210 1.5005
R13331 DVSS.n3355 DVSS.n3354 1.5005
R13332 DVSS.n3358 DVSS.n3357 1.5005
R13333 DVSS.n3360 DVSS.n3359 1.5005
R13334 DVSS.n3364 DVSS.n3363 1.5005
R13335 DVSS.n3366 DVSS.n3365 1.5005
R13336 DVSS.n3369 DVSS.n3368 1.5005
R13337 DVSS.n3370 DVSS.n3244 1.5005
R13338 DVSS.n3374 DVSS.n3373 1.5005
R13339 DVSS.n3425 DVSS.n3235 1.5005
R13340 DVSS.n3367 DVSS.n3228 1.5005
R13341 DVSS.n3430 DVSS.n3227 1.5005
R13342 DVSS.n3362 DVSS.n3361 1.5005
R13343 DVSS.n3438 DVSS.n3218 1.5005
R13344 DVSS.n3356 DVSS.n3211 1.5005
R13345 DVSS.n3443 DVSS.n3210 1.5005
R13346 DVSS.n3350 DVSS.n3349 1.5005
R13347 DVSS.n3450 DVSS.n3200 1.5005
R13348 DVSS.n3343 DVSS.n3193 1.5005
R13349 DVSS.n3455 DVSS.n3192 1.5005
R13350 DVSS.n3338 DVSS.n3337 1.5005
R13351 DVSS.n3462 DVSS.n3180 1.5005
R13352 DVSS.n3246 DVSS.n3173 1.5005
R13353 DVSS.n3467 DVSS.n3172 1.5005
R13354 DVSS.n3325 DVSS.n3324 1.5005
R13355 DVSS.n3474 DVSS.n3163 1.5005
R13356 DVSS.n3319 DVSS.n3156 1.5005
R13357 DVSS.n3479 DVSS.n3155 1.5005
R13358 DVSS.n3314 DVSS.n3313 1.5005
R13359 DVSS.n3488 DVSS.n3145 1.5005
R13360 DVSS.n3307 DVSS.n3138 1.5005
R13361 DVSS.n3493 DVSS.n3137 1.5005
R13362 DVSS.n3302 DVSS.n3301 1.5005
R13363 DVSS.n3500 DVSS.n3126 1.5005
R13364 DVSS.n3295 DVSS.n3119 1.5005
R13365 DVSS.n3505 DVSS.n3118 1.5005
R13366 DVSS.n3289 DVSS.n3288 1.5005
R13367 DVSS.n3513 DVSS.n3109 1.5005
R13368 DVSS.n3283 DVSS.n3102 1.5005
R13369 DVSS.n3518 DVSS.n3101 1.5005
R13370 DVSS.n3278 DVSS.n3277 1.5005
R13371 DVSS.n3525 DVSS.n3089 1.5005
R13372 DVSS.n3272 DVSS.n3082 1.5005
R13373 DVSS.n3530 DVSS.n3081 1.5005
R13374 DVSS.n3266 DVSS.n3265 1.5005
R13375 DVSS.n3538 DVSS.n3072 1.5005
R13376 DVSS.n3260 DVSS.n2675 1.5005
R13377 DVSS.n3543 DVSS.n2674 1.5005
R13378 DVSS.n3255 DVSS.n3254 1.5005
R13379 DVSS.n3551 DVSS.n3550 1.5005
R13380 DVSS.n3062 DVSS.n2681 1.5005
R13381 DVSS.n2687 DVSS.n2680 1.5005
R13382 DVSS.n3052 DVSS.n3050 1.5005
R13383 DVSS.n3042 DVSS.n3041 1.5005
R13384 DVSS.n2697 DVSS.n2689 1.5005
R13385 DVSS.n3034 DVSS.n2696 1.5005
R13386 DVSS.n3021 DVSS.n2702 1.5005
R13387 DVSS.n2708 DVSS.n2701 1.5005
R13388 DVSS.n3011 DVSS.n3009 1.5005
R13389 DVSS.n2996 DVSS.n2995 1.5005
R13390 DVSS.n2717 DVSS.n2710 1.5005
R13391 DVSS.n2987 DVSS.n2716 1.5005
R13392 DVSS.n2975 DVSS.n2722 1.5005
R13393 DVSS.n2926 DVSS.n2721 1.5005
R13394 DVSS.n2936 DVSS.n2730 1.5005
R13395 DVSS.n2964 DVSS.n2728 1.5005
R13396 DVSS.n2956 DVSS.n2735 1.5005
R13397 DVSS.n2741 DVSS.n2734 1.5005
R13398 DVSS.n2948 DVSS.n2946 1.5005
R13399 DVSS.n2921 DVSS.n2920 1.5005
R13400 DVSS.n2904 DVSS.n2743 1.5005
R13401 DVSS.n2875 DVSS.n2752 1.5005
R13402 DVSS.n2909 DVSS.n2751 1.5005
R13403 DVSS.n2893 DVSS.n2757 1.5005
R13404 DVSS.n2763 DVSS.n2756 1.5005
R13405 DVSS.n2886 DVSS.n2884 1.5005
R13406 DVSS.n2866 DVSS.n2865 1.5005
R13407 DVSS.n2772 DVSS.n2765 1.5005
R13408 DVSS.n2856 DVSS.n2771 1.5005
R13409 DVSS.n2844 DVSS.n2777 1.5005
R13410 DVSS.n2783 DVSS.n2776 1.5005
R13411 DVSS.n2837 DVSS.n2835 1.5005
R13412 DVSS.n2822 DVSS.n2821 1.5005
R13413 DVSS.n2792 DVSS.n2785 1.5005
R13414 DVSS.n2812 DVSS.n2791 1.5005
R13415 DVSS.n3373 DVSS.n3242 1.5005
R13416 DVSS.n3425 DVSS.n3424 1.5005
R13417 DVSS.n3237 DVSS.n3228 1.5005
R13418 DVSS.n3431 DVSS.n3430 1.5005
R13419 DVSS.n3361 DVSS.n3222 1.5005
R13420 DVSS.n3438 DVSS.n3437 1.5005
R13421 DVSS.n3220 DVSS.n3211 1.5005
R13422 DVSS.n3444 DVSS.n3443 1.5005
R13423 DVSS.n3349 DVSS.n3204 1.5005
R13424 DVSS.n3450 DVSS.n3449 1.5005
R13425 DVSS.n3202 DVSS.n3193 1.5005
R13426 DVSS.n3456 DVSS.n3455 1.5005
R13427 DVSS.n3337 DVSS.n3183 1.5005
R13428 DVSS.n3462 DVSS.n3461 1.5005
R13429 DVSS.n3185 DVSS.n3173 1.5005
R13430 DVSS.n3468 DVSS.n3467 1.5005
R13431 DVSS.n3324 DVSS.n3167 1.5005
R13432 DVSS.n3474 DVSS.n3473 1.5005
R13433 DVSS.n3165 DVSS.n3156 1.5005
R13434 DVSS.n3480 DVSS.n3479 1.5005
R13435 DVSS.n3313 DVSS.n3152 1.5005
R13436 DVSS.n3488 DVSS.n3487 1.5005
R13437 DVSS.n3147 DVSS.n3138 1.5005
R13438 DVSS.n3494 DVSS.n3493 1.5005
R13439 DVSS.n3301 DVSS.n3130 1.5005
R13440 DVSS.n3500 DVSS.n3499 1.5005
R13441 DVSS.n3128 DVSS.n3119 1.5005
R13442 DVSS.n3506 DVSS.n3505 1.5005
R13443 DVSS.n3288 DVSS.n3113 1.5005
R13444 DVSS.n3513 DVSS.n3512 1.5005
R13445 DVSS.n3111 DVSS.n3102 1.5005
R13446 DVSS.n3519 DVSS.n3518 1.5005
R13447 DVSS.n3277 DVSS.n3092 1.5005
R13448 DVSS.n3525 DVSS.n3524 1.5005
R13449 DVSS.n3094 DVSS.n3082 1.5005
R13450 DVSS.n3531 DVSS.n3530 1.5005
R13451 DVSS.n3265 DVSS.n3076 1.5005
R13452 DVSS.n3538 DVSS.n3537 1.5005
R13453 DVSS.n3074 DVSS.n2675 1.5005
R13454 DVSS.n3544 DVSS.n3543 1.5005
R13455 DVSS.n3254 DVSS.n2669 1.5005
R13456 DVSS.n3550 DVSS.n3549 1.5005
R13457 DVSS.n3062 DVSS.n3061 1.5005
R13458 DVSS.n3054 DVSS.n2680 1.5005
R13459 DVSS.n3053 DVSS.n3052 1.5005
R13460 DVSS.n3041 DVSS.n3040 1.5005
R13461 DVSS.n2697 DVSS.n2691 1.5005
R13462 DVSS.n3035 DVSS.n3034 1.5005
R13463 DVSS.n3021 DVSS.n3020 1.5005
R13464 DVSS.n3013 DVSS.n2701 1.5005
R13465 DVSS.n3012 DVSS.n3011 1.5005
R13466 DVSS.n2995 DVSS.n2994 1.5005
R13467 DVSS.n2717 DVSS.n2712 1.5005
R13468 DVSS.n2988 DVSS.n2987 1.5005
R13469 DVSS.n2975 DVSS.n2974 1.5005
R13470 DVSS.n2723 DVSS.n2721 1.5005
R13471 DVSS.n2730 DVSS.n2724 1.5005
R13472 DVSS.n2965 DVSS.n2964 1.5005
R13473 DVSS.n2956 DVSS.n2955 1.5005
R13474 DVSS.n2736 DVSS.n2734 1.5005
R13475 DVSS.n2949 DVSS.n2948 1.5005
R13476 DVSS.n2920 DVSS.n2919 1.5005
R13477 DVSS.n2904 DVSS.n2745 1.5005
R13478 DVSS.n2752 DVSS.n2747 1.5005
R13479 DVSS.n2910 DVSS.n2909 1.5005
R13480 DVSS.n2893 DVSS.n2892 1.5005
R13481 DVSS.n2758 DVSS.n2756 1.5005
R13482 DVSS.n2887 DVSS.n2886 1.5005
R13483 DVSS.n2865 DVSS.n2864 1.5005
R13484 DVSS.n2772 DVSS.n2767 1.5005
R13485 DVSS.n2857 DVSS.n2856 1.5005
R13486 DVSS.n2844 DVSS.n2843 1.5005
R13487 DVSS.n2778 DVSS.n2776 1.5005
R13488 DVSS.n2838 DVSS.n2837 1.5005
R13489 DVSS.n2821 DVSS.n2820 1.5005
R13490 DVSS.n2792 DVSS.n2787 1.5005
R13491 DVSS.n2813 DVSS.n2812 1.5005
R13492 DVSS.n3746 DVSS.n3745 1.5005
R13493 DVSS.n1214 DVSS.n1179 1.5005
R13494 DVSS.n1213 DVSS.n1212 1.5005
R13495 DVSS.n1211 DVSS.n1210 1.5005
R13496 DVSS.n1209 DVSS.n1208 1.5005
R13497 DVSS.n1207 DVSS.n1206 1.5005
R13498 DVSS.n1205 DVSS.n1204 1.5005
R13499 DVSS.n1203 DVSS.n1202 1.5005
R13500 DVSS.n1201 DVSS.n1200 1.5005
R13501 DVSS.n1199 DVSS.n1198 1.5005
R13502 DVSS.n1197 DVSS.n1196 1.5005
R13503 DVSS.n1195 DVSS.n1190 1.5005
R13504 DVSS.n4931 DVSS.n4930 1.5005
R13505 DVSS.n1860 DVSS.n1859 1.49818
R13506 DVSS.n3585 DVSS.n2243 1.49138
R13507 DVSS.n2152 DVSS.n2151 1.44688
R13508 DVSS.n1879 DVSS.n1813 1.44688
R13509 DVSS DVSS.n1276 1.41642
R13510 DVSS.n1283 DVSS 1.41642
R13511 DVSS.n4426 DVSS 1.41642
R13512 DVSS.n1309 DVSS 1.41642
R13513 DVSS DVSS.n4440 1.41642
R13514 DVSS DVSS.n1306 1.41642
R13515 DVSS.n1459 DVSS 1.41642
R13516 DVSS.n1471 DVSS 1.41642
R13517 DVSS.n4186 DVSS 1.41642
R13518 DVSS.n4392 DVSS 1.41642
R13519 DVSS.n4395 DVSS 1.41642
R13520 DVSS.n4337 DVSS 1.41642
R13521 DVSS.n4444 DVSS.n4443 1.39741
R13522 DVSS.n5115 DVSS.n5111 1.38664
R13523 DVSS.n1921 DVSS.n1814 1.35477
R13524 DVSS.n2160 DVSS.n1804 1.35477
R13525 DVSS.n3575 DVSS.n3573 1.328
R13526 DVSS.n1594 DVSS.n1588 1.31286
R13527 DVSS.n2236 DVSS.n1615 1.31286
R13528 DVSS.n2261 DVSS.n1647 1.31286
R13529 DVSS.n3676 DVSS.n1690 1.31286
R13530 DVSS.n4947 DVSS.n4946 1.3005
R13531 DVSS.n3950 DVSS.n3949 1.3005
R13532 DVSS.n3958 DVSS.n3957 1.3005
R13533 DVSS.n1484 DVSS.n1157 1.3005
R13534 DVSS.n4976 DVSS.n4975 1.3005
R13535 DVSS.n4388 DVSS.n4387 1.3005
R13536 DVSS.n4385 DVSS.n4384 1.3005
R13537 DVSS.n1457 DVSS.n1456 1.3005
R13538 DVSS.n1455 DVSS.n1454 1.3005
R13539 DVSS.n4464 DVSS.n1289 1.29067
R13540 DVSS.n4460 DVSS.n1294 1.29067
R13541 DVSS.n4407 DVSS.n4380 1.29067
R13542 DVSS.n1315 DVSS.n1314 1.29067
R13543 DVSS.n2248 VSS 1.28985
R13544 DVSS.n4942 DVSS.n1172 1.26649
R13545 DVSS.n3875 DVSS.n1580 1.25594
R13546 DVSS.n3788 DVSS.n3787 1.25594
R13547 DVSS.n1515 DVSS.n1514 1.20054
R13548 DVSS.n1515 DVSS.n1507 1.19935
R13549 DVSS.n4979 DVSS.n4978 1.19925
R13550 DVSS.n4427 DVSS.n4426 1.16866
R13551 DVSS.n1472 DVSS.n1471 1.16866
R13552 DVSS.n4186 DVSS.n4185 1.16866
R13553 DVSS.n4393 DVSS.n4392 1.16866
R13554 DVSS.n4337 DVSS.n4336 1.16866
R13555 DVSS.n3616 DVSS.n1688 1.16402
R13556 DVSS.n4471 DVSS.n1278 1.15745
R13557 DVSS.n3587 DVSS.n3586 1.15606
R13558 DVSS.n4456 DVSS.n4455 1.15606
R13559 DVSS.n4448 DVSS.n4447 1.15606
R13560 DVSS.n4965 DVSS.n4964 1.15606
R13561 DVSS.n4957 DVSS.n4956 1.15606
R13562 DVSS.n2231 DVSS.n2228 1.13009
R13563 DVSS.n3617 DVSS.n3608 1.12941
R13564 DVSS.n3602 DVSS.n1654 1.10843
R13565 DVSS.n2262 DVSS.n2261 1.10563
R13566 DVSS.n3761 DVSS.n1690 1.10563
R13567 DVSS.n3566 DVSS.n1588 1.10563
R13568 DVSS.n2237 DVSS.n2236 1.10563
R13569 DVSS.n1732 DVSS.t108 1.0925
R13570 DVSS.n4469 DVSS.t2 1.0925
R13571 DVSS.n4469 DVSS.t178 1.0925
R13572 DVSS.n1691 DVSS.t24 1.0925
R13573 DVSS.n1691 DVSS.t127 1.0925
R13574 DVSS.n1655 DVSS.t184 1.0925
R13575 DVSS.n1655 DVSS.t14 1.0925
R13576 DVSS.n1575 DVSS.t79 1.0925
R13577 DVSS.n1575 DVSS.t155 1.0925
R13578 DVSS.n1583 DVSS.t135 1.0925
R13579 DVSS.n1583 DVSS.t123 1.0925
R13580 DVSS.n3607 DVSS.t158 1.0925
R13581 DVSS.n4394 DVSS.n1316 1.08844
R13582 DVSS.n4428 DVSS.n1316 1.08844
R13583 DVSS.n1474 DVSS.n1473 1.08844
R13584 DVSS.n1474 DVSS.n1285 1.08844
R13585 DVSS.n4429 DVSS.n4428 1.0805
R13586 DVSS.n1473 DVSS.n1468 1.0805
R13587 DVSS.n4480 DVSS.n1285 1.0805
R13588 DVSS.n4403 DVSS.n4394 1.0805
R13589 DVSS.n3602 DVSS.n1688 1.07932
R13590 DVSS.n4528 DVSS.n956 1.07349
R13591 DVSS.n1900 DVSS.n1890 1.05604
R13592 DVSS.n1281 DVSS.n1280 1.0505
R13593 DVSS.n4437 DVSS.n4436 1.0505
R13594 DVSS.n1463 DVSS.n1462 1.0505
R13595 DVSS.n4399 DVSS.n4398 1.0505
R13596 DVSS.n1449 DVSS.n1446 1.05029
R13597 DVSS.n3571 DVSS.n3570 1.0405
R13598 DVSS.n3570 DVSS.n3569 1.0405
R13599 DVSS.n3579 DVSS.n3578 1.0405
R13600 DVSS.n2257 DVSS.n2256 1.0405
R13601 DVSS.n2256 DVSS.n2255 1.0405
R13602 DVSS.n1697 DVSS.n1696 1.0405
R13603 DVSS.n1696 DVSS.n1695 1.0405
R13604 DVSS.n2229 DVSS.n1731 1.0405
R13605 DVSS.n1453 DVSS.n1452 1.0405
R13606 DVSS.n4407 DVSS.n4406 1.0405
R13607 DVSS.n4406 DVSS.n4405 1.0405
R13608 DVSS.n4460 DVSS.n4459 1.0405
R13609 DVSS.n4459 DVSS.n4458 1.0405
R13610 DVSS.n4432 DVSS.n1315 1.0405
R13611 DVSS.n4432 DVSS.n4431 1.0405
R13612 DVSS.n4465 DVSS.n4464 1.0405
R13613 DVSS.n4466 DVSS.n4465 1.0405
R13614 DVSS.n1161 DVSS.n1160 1.02439
R13615 DVSS.n1298 DVSS.n1297 1.02439
R13616 DVSS.n4450 DVSS.n4449 1.02439
R13617 DVSS.n4959 DVSS.n4958 1.02439
R13618 DVSS.t27 DVSS.n3759 1.00732
R13619 DVSS.n3789 DVSS.n3788 1.00517
R13620 DVSS.n1586 DVSS.n1580 1.00517
R13621 DVSS.n3904 VSS 1.00241
R13622 DVSS.n2232 DVSS.n1731 0.998488
R13623 DVSS.n3578 DVSS.n3577 0.996088
R13624 DVSS.n1452 DVSS.n1451 0.996088
R13625 DVSS.n3582 DVSS.t59 0.958395
R13626 DVSS.n3582 DVSS.t58 0.958395
R13627 DVSS.n3245 DVSS.t49 0.9581
R13628 DVSS.n3330 DVSS.t36 0.9581
R13629 DVSS.n3298 DVSS.t46 0.9581
R13630 DVSS.n3253 DVSS.t34 0.9581
R13631 DVSS.n3000 DVSS.t45 0.9581
R13632 DVSS.n2939 DVSS.t38 0.9581
R13633 DVSS.n2869 DVSS.t48 0.9581
R13634 DVSS.n2797 DVSS.t35 0.9581
R13635 DVSS.n1705 DVSS.t39 0.9581
R13636 DVSS.n1707 DVSS.t33 0.9581
R13637 DVSS.n1707 DVSS.t39 0.9581
R13638 DVSS.n3651 DVSS.t33 0.9581
R13639 DVSS.n3434 DVSS.t49 0.9581
R13640 DVSS.n3184 DVSS.t36 0.9581
R13641 DVSS.n3133 DVSS.t46 0.9581
R13642 DVSS.n3534 DVSS.t34 0.9581
R13643 DVSS.n2692 DVSS.t45 0.9581
R13644 DVSS.n2725 DVSS.t38 0.9581
R13645 DVSS.n2861 DVSS.t48 0.9581
R13646 DVSS.n2795 DVSS.t35 0.9581
R13647 DVSS.n2276 DVSS.n1167 0.945955
R13648 DVSS.n3904 DVSS.n3903 0.945955
R13649 DVSS.n4454 DVSS.n4453 0.945955
R13650 DVSS.n4978 DVSS.n4977 0.945955
R13651 DVSS.n4963 DVSS.n4962 0.945955
R13652 DVSS.n1277 DVSS.n1276 0.941532
R13653 DVSS.n4441 DVSS.n4440 0.941532
R13654 DVSS.n1307 DVSS.n1306 0.941532
R13655 DVSS.n1282 DVSS.n1281 0.941367
R13656 DVSS.n1284 DVSS.n1283 0.941367
R13657 DVSS.n1310 DVSS.n1309 0.941367
R13658 DVSS.n4438 DVSS.n4437 0.941367
R13659 DVSS.n1464 DVSS.n1463 0.941367
R13660 DVSS.n1460 DVSS.n1459 0.941367
R13661 DVSS.n4396 DVSS.n4395 0.941367
R13662 DVSS.n4400 DVSS.n4399 0.941367
R13663 DVSS.n2655 DVSS.n2654 0.922809
R13664 DVSS.n2396 DVSS.n2264 0.922714
R13665 DVSS.n1534 DVSS.n1081 0.922457
R13666 DVSS.n5109 DVSS.n5108 0.922457
R13667 DVSS.n3941 DVSS.n3940 0.910322
R13668 DVSS.n955 DVSS.n952 0.902366
R13669 DVSS.n5361 DVSS.n952 0.902313
R13670 DVSS.n5361 DVSS.n5360 0.902282
R13671 DVSS.n5360 DVSS.n955 0.901878
R13672 DVSS.n3745 DVSS.n3653 0.882658
R13673 DVSS.n5358 DVSS.n956 0.879171
R13674 DVSS.n4929 DVSS.n1193 0.879171
R13675 DVSS.n3793 DVSS.n3792 0.875366
R13676 DVSS.n3769 DVSS.n3768 0.875366
R13677 DVSS.n1658 DVSS.n1648 0.87493
R13678 DVSS.n4424 DVSS.n4423 0.8749
R13679 DVSS.n1469 DVSS.n1354 0.8749
R13680 DVSS.n4340 DVSS.n4339 0.8749
R13681 DVSS.n3939 DVSS.n1518 0.873402
R13682 DVSS.n1280 DVSS.n1279 0.872079
R13683 DVSS.n4436 DVSS.n4435 0.872079
R13684 DVSS.n1462 DVSS.n1461 0.872079
R13685 DVSS.n4398 DVSS.n4397 0.872079
R13686 DVSS.n4930 DVSS.n4929 0.870066
R13687 DVSS.n3897 DVSS.n1587 0.867167
R13688 DVSS.n3902 DVSS.n3901 0.867167
R13689 DVSS.n3791 DVSS.n3790 0.867167
R13690 DVSS.n3766 DVSS.n3762 0.867167
R13691 DVSS.n2258 DVSS.n2257 0.843937
R13692 DVSS.n3572 DVSS.n3571 0.843937
R13693 DVSS.n3757 DVSS.n1697 0.843937
R13694 DVSS.n3581 DVSS.n1654 0.827218
R13695 DVSS.n5555 DVSS.n5554 0.820816
R13696 DVSS.n3573 DVSS.n1698 0.815237
R13697 DVSS.n3616 DVSS.n3615 0.80914
R13698 DVSS.n4476 DVSS.n4473 0.8005
R13699 DVSS.n3961 DVSS.n1501 0.796907
R13700 DVSS.n3961 DVSS.n1499 0.796907
R13701 DVSS.n3965 DVSS.n1499 0.796907
R13702 DVSS.n3965 DVSS.n1497 0.796907
R13703 DVSS.n3970 DVSS.n1497 0.796907
R13704 DVSS.n3970 DVSS.n1495 0.796907
R13705 DVSS.n3974 DVSS.n1495 0.796907
R13706 DVSS.n3974 DVSS.n1442 0.796907
R13707 DVSS.n3979 DVSS.n1442 0.796907
R13708 DVSS.n2276 VSS 0.78605
R13709 DVSS.n1919 DVSS.n1866 0.778288
R13710 DVSS.n4238 DVSS.n1301 0.774059
R13711 DVSS.n4942 DVSS.n4941 0.752663
R13712 DVSS.n2240 DVSS.n2239 0.751952
R13713 DVSS.n3754 VSS 0.751638
R13714 DVSS.n1880 DVSS.n1879 0.7505
R13715 DVSS.n2151 DVSS.n1811 0.7505
R13716 DVSS DVSS.n2231 0.746344
R13717 DVSS.n5616 DVSS.n5615 0.745113
R13718 DVSS.n688 DVSS.n169 0.745113
R13719 DVSS.n620 DVSS.n194 0.745113
R13720 DVSS.n1923 DVSS.n1815 0.743357
R13721 DVSS.n1923 DVSS.n1922 0.743357
R13722 DVSS.n2162 DVSS.n1805 0.743357
R13723 DVSS.n2162 DVSS.n2161 0.743357
R13724 DVSS.n2153 DVSS.n1806 0.743357
R13725 DVSS.n2161 DVSS.n1806 0.743357
R13726 DVSS.n1818 DVSS.n1803 0.743357
R13727 DVSS.n1922 DVSS.n1803 0.743357
R13728 DVSS.n5616 DVSS.n123 0.736857
R13729 DVSS.n688 DVSS.n687 0.736857
R13730 DVSS.n621 DVSS.n620 0.736857
R13731 DVSS.n2155 DVSS.n2154 0.735937
R13732 DVSS.n1916 DVSS.n1915 0.735937
R13733 DVSS.n4483 DVSS.n1278 0.7304
R13734 DVSS.n3794 DVSS.n3793 0.71546
R13735 DVSS.n3770 DVSS.n3769 0.71546
R13736 DVSS.n3802 DVSS.n1648 0.71533
R13737 DVSS.n1468 DVSS.n1467 0.707265
R13738 DVSS.n3619 DVSS.n3605 0.696386
R13739 DVSS.n3618 DVSS.n3606 0.696386
R13740 DVSS.n4382 DVSS.n1312 0.693432
R13741 DVSS.n4389 DVSS.n4378 0.693432
R13742 DVSS.n1295 DVSS.n1292 0.693432
R13743 DVSS.n1290 DVSS.n1287 0.693432
R13744 DVSS.n4461 DVSS.n1292 0.682241
R13745 DVSS.n4408 DVSS.n4378 0.682241
R13746 DVSS.n4382 DVSS.n4377 0.682241
R13747 DVSS.n4463 DVSS.n1290 0.682241
R13748 DVSS.n1864 DVSS.n1860 0.666308
R13749 DVSS.n3982 DVSS.n3981 0.66242
R13750 DVSS.n4429 DVSS.n1311 0.662265
R13751 DVSS.n4481 DVSS.n4480 0.662265
R13752 DVSS.n4403 DVSS.n4402 0.662265
R13753 DVSS.n1865 DVSS.n1864 0.64762
R13754 DVSS.n3619 DVSS.n3618 0.646382
R13755 DVSS.n4777 DVSS.n4776 0.643357
R13756 DVSS.n4792 DVSS.n4791 0.643357
R13757 DVSS.n4794 DVSS.n4787 0.643357
R13758 DVSS.n4887 DVSS.n4886 0.643357
R13759 DVSS.n4756 DVSS.n4755 0.643357
R13760 DVSS.n4757 DVSS.n1218 0.643357
R13761 DVSS.n4920 DVSS.n4919 0.643357
R13762 DVSS.n1221 DVSS.n1219 0.643357
R13763 DVSS.n4717 DVSS.n4716 0.643357
R13764 DVSS.n4720 DVSS.n4719 0.643357
R13765 DVSS.n1242 DVSS.n1241 0.643357
R13766 DVSS.n4734 DVSS.n4733 0.643357
R13767 DVSS.n4615 DVSS.n1271 0.643357
R13768 DVSS.n4681 DVSS.n4680 0.643357
R13769 DVSS.n1263 DVSS.n1262 0.643357
R13770 DVSS.n4694 DVSS.n4693 0.643357
R13771 DVSS.n4584 DVSS.n4583 0.643357
R13772 DVSS.n4599 DVSS.n4598 0.643357
R13773 DVSS.n4601 DVSS.n4594 0.643357
R13774 DVSS.n4639 DVSS.n4638 0.643357
R13775 DVSS.n4563 DVSS.n4562 0.643357
R13776 DVSS.n4564 DVSS.n4492 0.643357
R13777 DVSS.n4672 DVSS.n4671 0.643357
R13778 DVSS.n4495 DVSS.n4493 0.643357
R13779 DVSS.n3949 DVSS.n3948 0.634889
R13780 DVSS.n1503 VSS 0.622069
R13781 DVSS.n3946 VSS 0.622069
R13782 DVSS.n1483 VSS 0.622069
R13783 DVSS.n4970 VSS 0.622069
R13784 DVSS.n1168 VSS 0.622069
R13785 DVSS.n3618 DVSS.n3617 0.618588
R13786 DVSS.n3649 DVSS.n3648 0.612265
R13787 DVSS.n3982 DVSS 0.600908
R13788 DVSS.n4482 DVSS.n1282 0.597759
R13789 DVSS.n4481 DVSS.n1284 0.597759
R13790 DVSS.n1311 DVSS.n1310 0.597759
R13791 DVSS.n4439 DVSS.n4438 0.597759
R13792 DVSS.n1465 DVSS.n1464 0.597759
R13793 DVSS.n4402 DVSS.n4396 0.597759
R13794 DVSS.n4401 DVSS.n4400 0.597759
R13795 DVSS DVSS.n1277 0.595564
R13796 DVSS DVSS.n4441 0.595564
R13797 DVSS DVSS.n1307 0.595564
R13798 DVSS.n3634 DVSS.n3633 0.588678
R13799 DVSS.n2259 DVSS.n2258 0.585632
R13800 DVSS.n3572 DVSS.n2247 0.585632
R13801 DVSS.n3758 DVSS.n3757 0.585632
R13802 DVSS.n2261 DVSS.n1659 0.584525
R13803 DVSS.n3767 DVSS.n1690 0.584525
R13804 DVSS.n3896 DVSS.n1588 0.584525
R13805 DVSS.n2236 DVSS.n1574 0.584525
R13806 DVSS.n1448 VSS 0.581806
R13807 DVSS.n3634 DVSS.n1715 0.578278
R13808 DVSS.n3635 DVSS.n3594 0.578278
R13809 DVSS.n3636 DVSS.n1729 0.578278
R13810 DVSS.n3637 DVSS.n3595 0.578278
R13811 DVSS.n3638 DVSS.n1728 0.578278
R13812 DVSS.n3639 DVSS.n3596 0.578278
R13813 DVSS.n3640 DVSS.n1727 0.578278
R13814 DVSS.n3641 DVSS.n3597 0.578278
R13815 DVSS.n3642 DVSS.n1726 0.578278
R13816 DVSS.n3644 DVSS.n3643 0.578278
R13817 DVSS.n3629 DVSS.n3628 0.578278
R13818 DVSS.n3646 DVSS.n1724 0.578278
R13819 DVSS.n3748 DVSS 0.578278
R13820 DVSS.n3749 DVSS.n3748 0.578278
R13821 DVSS.n2796 DVSS.n2661 0.578278
R13822 DVSS.n3980 DVSS.n3979 0.578278
R13823 DVSS.n3979 DVSS.n3978 0.578278
R13824 DVSS.n1442 DVSS.n1441 0.578278
R13825 DVSS.n3977 DVSS.n1442 0.578278
R13826 DVSS.n3974 DVSS.n3973 0.578278
R13827 DVSS.n3975 DVSS.n3974 0.578278
R13828 DVSS.n3972 DVSS.n1495 0.578278
R13829 DVSS.n3968 DVSS.n1495 0.578278
R13830 DVSS.n3971 DVSS.n3970 0.578278
R13831 DVSS.n3970 DVSS.n3969 0.578278
R13832 DVSS.n1497 DVSS.n1496 0.578278
R13833 DVSS.n3967 DVSS.n1497 0.578278
R13834 DVSS.n3965 DVSS.n3964 0.578278
R13835 DVSS.n3966 DVSS.n3965 0.578278
R13836 DVSS.n3963 DVSS.n1499 0.578278
R13837 DVSS.n1499 DVSS.n1498 0.578278
R13838 DVSS.n3962 DVSS.n3961 0.578278
R13839 DVSS.n3961 DVSS.n3960 0.578278
R13840 DVSS.n1501 DVSS.n1500 0.578278
R13841 DVSS.n1502 DVSS.n1501 0.578278
R13842 DVSS.n3757 DVSS.n3756 0.563
R13843 DVSS.n4453 DVSS.n4452 0.557079
R13844 DVSS.n3586 DVSS.n3585 0.557079
R13845 DVSS.n3576 DVSS.n3575 0.557079
R13846 DVSS.n4978 DVSS.n1155 0.557079
R13847 DVSS.n4962 DVSS.n4961 0.557079
R13848 DVSS.n1488 DVSS.n1484 0.553108
R13849 DVSS.n4975 DVSS.n4974 0.553108
R13850 DVSS.n4951 DVSS.n4947 0.553108
R13851 DVSS.n1467 DVSS.n1460 0.548022
R13852 DVSS.n1160 DVSS.t97 0.5465
R13853 DVSS.n1160 DVSS.t137 0.5465
R13854 DVSS.n1297 DVSS.t145 0.5465
R13855 DVSS.n1297 DVSS.t166 0.5465
R13856 DVSS.n4449 DVSS.t91 0.5465
R13857 DVSS.n4449 DVSS.t182 0.5465
R13858 DVSS.n4958 DVSS.t82 0.5465
R13859 DVSS.n4958 DVSS.t195 0.5465
R13860 DVSS.n3562 DVSS.n3561 0.545794
R13861 DVSS.n4477 DVSS.n4476 0.545794
R13862 DVSS.n4482 DVSS.n4481 0.545794
R13863 DVSS.n4439 DVSS.n1311 0.545794
R13864 DVSS.n4442 DVSS.n4439 0.545794
R13865 DVSS.n1465 DVSS.n1308 0.545794
R13866 DVSS.n3791 DVSS.n1659 0.545794
R13867 DVSS.n3767 DVSS.n3766 0.545794
R13868 DVSS.n3901 DVSS.n1574 0.545794
R13869 DVSS.n3897 DVSS.n3896 0.545794
R13870 DVSS.n4402 DVSS.n4401 0.545794
R13871 DVSS.n4401 DVSS.n1172 0.545794
R13872 DVSS.n4428 DVSS.n4427 0.5442
R13873 DVSS.n1473 DVSS.n1472 0.5442
R13874 DVSS.n4185 DVSS.n1285 0.5442
R13875 DVSS.n4394 DVSS.n4393 0.5442
R13876 DVSS.n1518 VSS 0.544091
R13877 DVSS.n3941 VSS 0.544091
R13878 DVSS.n2251 DVSS.n2250 0.543147
R13879 DVSS.n4336 DVSS 0.541831
R13880 DVSS.n2242 DVSS.n2240 0.536572
R13881 DVSS.n4390 DVSS.n1164 0.532494
R13882 DVSS.n1915 DVSS.n1815 0.5255
R13883 DVSS.n2154 DVSS.n2153 0.5255
R13884 DVSS.n3568 DVSS.n2247 0.5205
R13885 DVSS.n2260 DVSS.n2259 0.5205
R13886 DVSS.n3759 DVSS.n3758 0.5205
R13887 DVSS.n1162 DVSS.n1161 0.518873
R13888 DVSS.n1299 DVSS.n1298 0.518873
R13889 DVSS.n4451 DVSS.n4450 0.518873
R13890 DVSS.n4960 DVSS.n4959 0.518873
R13891 DVSS.n3611 DVSS.t4 0.512375
R13892 DVSS.n3611 DVSS.t30 0.512375
R13893 DVSS.n3609 DVSS.t116 0.512375
R13894 DVSS.n3609 DVSS.t26 0.512375
R13895 DVSS.n1450 VSS 0.50383
R13896 DVSS.n1289 DVSS.n1288 0.500875
R13897 DVSS.n1294 DVSS.n1293 0.500875
R13898 DVSS.n4380 DVSS.n4379 0.500875
R13899 DVSS.n1314 DVSS.n1313 0.500875
R13900 DVSS.n2810 DVSS.n2805 0.5005
R13901 DVSS.n2809 DVSS.n2806 0.5005
R13902 DVSS.n2808 DVSS.n2807 0.5005
R13903 DVSS.n2775 DVSS.n2774 0.5005
R13904 DVSS.n2847 DVSS.n2846 0.5005
R13905 DVSS.n2848 DVSS.n2773 0.5005
R13906 DVSS.n2854 DVSS.n2849 0.5005
R13907 DVSS.n2853 DVSS.n2850 0.5005
R13908 DVSS.n2852 DVSS.n2851 0.5005
R13909 DVSS.n2755 DVSS.n2754 0.5005
R13910 DVSS.n2896 DVSS.n2895 0.5005
R13911 DVSS.n2897 DVSS.n2753 0.5005
R13912 DVSS.n2907 DVSS.n2898 0.5005
R13913 DVSS.n2906 DVSS.n2899 0.5005
R13914 DVSS.n2903 DVSS.n2900 0.5005
R13915 DVSS.n2902 DVSS.n2901 0.5005
R13916 DVSS.n2733 DVSS.n2732 0.5005
R13917 DVSS.n2959 DVSS.n2958 0.5005
R13918 DVSS.n2960 DVSS.n2731 0.5005
R13919 DVSS.n2962 DVSS.n2961 0.5005
R13920 DVSS.n2720 DVSS.n2719 0.5005
R13921 DVSS.n2978 DVSS.n2977 0.5005
R13922 DVSS.n2979 DVSS.n2718 0.5005
R13923 DVSS.n2985 DVSS.n2980 0.5005
R13924 DVSS.n2984 DVSS.n2981 0.5005
R13925 DVSS.n2983 DVSS.n2982 0.5005
R13926 DVSS.n2700 DVSS.n2699 0.5005
R13927 DVSS.n3024 DVSS.n3023 0.5005
R13928 DVSS.n3025 DVSS.n2698 0.5005
R13929 DVSS.n3032 DVSS.n3026 0.5005
R13930 DVSS.n3031 DVSS.n3027 0.5005
R13931 DVSS.n3030 DVSS.n3029 0.5005
R13932 DVSS.n3028 DVSS.n2678 0.5005
R13933 DVSS.n3064 DVSS.n2679 0.5005
R13934 DVSS.n3065 DVSS.n2677 0.5005
R13935 DVSS.n3067 DVSS.n3066 0.5005
R13936 DVSS.n3068 DVSS.n2676 0.5005
R13937 DVSS.n3541 DVSS.n3069 0.5005
R13938 DVSS.n3540 DVSS.n3070 0.5005
R13939 DVSS.n3084 DVSS.n3071 0.5005
R13940 DVSS.n3085 DVSS.n3083 0.5005
R13941 DVSS.n3528 DVSS.n3086 0.5005
R13942 DVSS.n3527 DVSS.n3087 0.5005
R13943 DVSS.n3104 DVSS.n3088 0.5005
R13944 DVSS.n3105 DVSS.n3103 0.5005
R13945 DVSS.n3516 DVSS.n3106 0.5005
R13946 DVSS.n3515 DVSS.n3107 0.5005
R13947 DVSS.n3121 DVSS.n3108 0.5005
R13948 DVSS.n3122 DVSS.n3120 0.5005
R13949 DVSS.n3503 DVSS.n3123 0.5005
R13950 DVSS.n3502 DVSS.n3124 0.5005
R13951 DVSS.n3140 DVSS.n3125 0.5005
R13952 DVSS.n3141 DVSS.n3139 0.5005
R13953 DVSS.n3491 DVSS.n3142 0.5005
R13954 DVSS.n3490 DVSS.n3143 0.5005
R13955 DVSS.n3158 DVSS.n3144 0.5005
R13956 DVSS.n3159 DVSS.n3157 0.5005
R13957 DVSS.n3477 DVSS.n3160 0.5005
R13958 DVSS.n3476 DVSS.n3161 0.5005
R13959 DVSS.n3175 DVSS.n3162 0.5005
R13960 DVSS.n3176 DVSS.n3174 0.5005
R13961 DVSS.n3465 DVSS.n3177 0.5005
R13962 DVSS.n3464 DVSS.n3178 0.5005
R13963 DVSS.n3195 DVSS.n3179 0.5005
R13964 DVSS.n3196 DVSS.n3194 0.5005
R13965 DVSS.n3453 DVSS.n3197 0.5005
R13966 DVSS.n3452 DVSS.n3198 0.5005
R13967 DVSS.n3213 DVSS.n3199 0.5005
R13968 DVSS.n3214 DVSS.n3212 0.5005
R13969 DVSS.n3441 DVSS.n3215 0.5005
R13970 DVSS.n3440 DVSS.n3216 0.5005
R13971 DVSS.n3230 DVSS.n3217 0.5005
R13972 DVSS.n3231 DVSS.n3229 0.5005
R13973 DVSS.n3428 DVSS.n3232 0.5005
R13974 DVSS.n3427 DVSS.n3233 0.5005
R13975 DVSS.n3378 DVSS.n3234 0.5005
R13976 DVSS.n3379 DVSS.n3377 0.5005
R13977 DVSS.n3416 DVSS.n3380 0.5005
R13978 DVSS.n3415 DVSS.n3381 0.5005
R13979 DVSS.n3414 DVSS.n3382 0.5005
R13980 DVSS.n3384 DVSS.n3383 0.5005
R13981 DVSS.n3410 DVSS.n3385 0.5005
R13982 DVSS.n3409 DVSS.n3386 0.5005
R13983 DVSS.n3389 DVSS.n3387 0.5005
R13984 DVSS.n3405 DVSS.n3390 0.5005
R13985 DVSS.n3404 DVSS.n3391 0.5005
R13986 DVSS.n3403 DVSS.n3392 0.5005
R13987 DVSS.n3394 DVSS.n3393 0.5005
R13988 DVSS.n3399 DVSS.n3395 0.5005
R13989 DVSS.n3398 DVSS.n3396 0.5005
R13990 DVSS.n3411 DVSS.n3410 0.5005
R13991 DVSS.n3412 DVSS.n3383 0.5005
R13992 DVSS.n3414 DVSS.n3413 0.5005
R13993 DVSS.n3415 DVSS.n3376 0.5005
R13994 DVSS.n3417 DVSS.n3416 0.5005
R13995 DVSS.n3377 DVSS.n3243 0.5005
R13996 DVSS.n3236 DVSS.n3234 0.5005
R13997 DVSS.n3427 DVSS.n3426 0.5005
R13998 DVSS.n3429 DVSS.n3428 0.5005
R13999 DVSS.n3229 DVSS.n3226 0.5005
R14000 DVSS.n3219 DVSS.n3217 0.5005
R14001 DVSS.n3440 DVSS.n3439 0.5005
R14002 DVSS.n3442 DVSS.n3441 0.5005
R14003 DVSS.n3212 DVSS.n3209 0.5005
R14004 DVSS.n3201 DVSS.n3199 0.5005
R14005 DVSS.n3452 DVSS.n3451 0.5005
R14006 DVSS.n3454 DVSS.n3453 0.5005
R14007 DVSS.n3194 DVSS.n3191 0.5005
R14008 DVSS.n3181 DVSS.n3179 0.5005
R14009 DVSS.n3464 DVSS.n3463 0.5005
R14010 DVSS.n3466 DVSS.n3465 0.5005
R14011 DVSS.n3174 DVSS.n3171 0.5005
R14012 DVSS.n3164 DVSS.n3162 0.5005
R14013 DVSS.n3476 DVSS.n3475 0.5005
R14014 DVSS.n3478 DVSS.n3477 0.5005
R14015 DVSS.n3157 DVSS.n3154 0.5005
R14016 DVSS.n3146 DVSS.n3144 0.5005
R14017 DVSS.n3490 DVSS.n3489 0.5005
R14018 DVSS.n3492 DVSS.n3491 0.5005
R14019 DVSS.n3139 DVSS.n3136 0.5005
R14020 DVSS.n3127 DVSS.n3125 0.5005
R14021 DVSS.n3502 DVSS.n3501 0.5005
R14022 DVSS.n3504 DVSS.n3503 0.5005
R14023 DVSS.n3120 DVSS.n3117 0.5005
R14024 DVSS.n3110 DVSS.n3108 0.5005
R14025 DVSS.n3515 DVSS.n3514 0.5005
R14026 DVSS.n3517 DVSS.n3516 0.5005
R14027 DVSS.n3103 DVSS.n3100 0.5005
R14028 DVSS.n3090 DVSS.n3088 0.5005
R14029 DVSS.n3527 DVSS.n3526 0.5005
R14030 DVSS.n3529 DVSS.n3528 0.5005
R14031 DVSS.n3083 DVSS.n3080 0.5005
R14032 DVSS.n3073 DVSS.n3071 0.5005
R14033 DVSS.n3540 DVSS.n3539 0.5005
R14034 DVSS.n3542 DVSS.n3541 0.5005
R14035 DVSS.n2676 DVSS.n2673 0.5005
R14036 DVSS.n3066 DVSS.n2667 0.5005
R14037 DVSS.n3065 DVSS.n2666 0.5005
R14038 DVSS.n3064 DVSS.n3063 0.5005
R14039 DVSS.n3051 DVSS.n2678 0.5005
R14040 DVSS.n3030 DVSS.n2685 0.5005
R14041 DVSS.n3031 DVSS.n2690 0.5005
R14042 DVSS.n3033 DVSS.n3032 0.5005
R14043 DVSS.n2698 DVSS.n2694 0.5005
R14044 DVSS.n3023 DVSS.n3022 0.5005
R14045 DVSS.n3010 DVSS.n2700 0.5005
R14046 DVSS.n2983 DVSS.n2706 0.5005
R14047 DVSS.n2984 DVSS.n2711 0.5005
R14048 DVSS.n2986 DVSS.n2985 0.5005
R14049 DVSS.n2718 DVSS.n2715 0.5005
R14050 DVSS.n2977 DVSS.n2976 0.5005
R14051 DVSS.n2729 DVSS.n2720 0.5005
R14052 DVSS.n2963 DVSS.n2962 0.5005
R14053 DVSS.n2731 DVSS.n2727 0.5005
R14054 DVSS.n2958 DVSS.n2957 0.5005
R14055 DVSS.n2947 DVSS.n2733 0.5005
R14056 DVSS.n2902 DVSS.n2739 0.5005
R14057 DVSS.n2903 DVSS.n2744 0.5005
R14058 DVSS.n2906 DVSS.n2905 0.5005
R14059 DVSS.n2908 DVSS.n2907 0.5005
R14060 DVSS.n2753 DVSS.n2750 0.5005
R14061 DVSS.n2895 DVSS.n2894 0.5005
R14062 DVSS.n2885 DVSS.n2755 0.5005
R14063 DVSS.n2852 DVSS.n2761 0.5005
R14064 DVSS.n2853 DVSS.n2766 0.5005
R14065 DVSS.n2855 DVSS.n2854 0.5005
R14066 DVSS.n2773 DVSS.n2770 0.5005
R14067 DVSS.n2846 DVSS.n2845 0.5005
R14068 DVSS.n2836 DVSS.n2775 0.5005
R14069 DVSS.n2808 DVSS.n2781 0.5005
R14070 DVSS.n2809 DVSS.n2786 0.5005
R14071 DVSS.n2811 DVSS.n2810 0.5005
R14072 DVSS.n2793 DVSS.n2790 0.5005
R14073 DVSS.n3409 DVSS.n3408 0.5005
R14074 DVSS.n3407 DVSS.n3387 0.5005
R14075 DVSS.n3406 DVSS.n3405 0.5005
R14076 DVSS.n3404 DVSS.n3388 0.5005
R14077 DVSS.n3403 DVSS.n3402 0.5005
R14078 DVSS.n3401 DVSS.n3393 0.5005
R14079 DVSS.n3400 DVSS.n3399 0.5005
R14080 DVSS.n4477 DVSS.n4468 0.497977
R14081 DVSS.n4476 DVSS.n4470 0.497977
R14082 DVSS.n4475 DVSS.n4474 0.497977
R14083 DVSS.n3788 DVSS.n1660 0.497868
R14084 DVSS.n3899 DVSS.n1580 0.497868
R14085 DVSS.n3940 DVSS.n1517 0.495738
R14086 DVSS.n5811 DVSS.n5809 0.490418
R14087 DVSS.n3621 DVSS.n3620 0.477527
R14088 DVSS.n3622 DVSS.n3621 0.473227
R14089 DVSS.n2249 DVSS.n2248 0.473227
R14090 DVSS.n3575 DVSS.n3574 0.473227
R14091 DVSS.n3574 DVSS.n2244 0.473227
R14092 DVSS.n3754 DVSS.n3753 0.473227
R14093 DVSS.n3753 DVSS.n3752 0.473227
R14094 DVSS.n2231 DVSS.n2230 0.473227
R14095 DVSS.n4476 DVSS 0.469029
R14096 DVSS.n1466 DVSS.n1465 0.465755
R14097 DVSS.n4850 DVSS.n4848 0.455549
R14098 DVSS.n1535 DVSS.n1534 0.455549
R14099 DVSS.n2654 DVSS.n2653 0.455549
R14100 DVSS.n5108 DVSS.n1082 0.455549
R14101 DVSS.n2399 DVSS.n2396 0.455549
R14102 DVSS.n1101 DVSS.n1100 0.452884
R14103 DVSS.n2277 DVSS.n2276 0.452868
R14104 DVSS.n5075 DVSS.n1101 0.452744
R14105 DVSS.n950 DVSS.n949 0.4505
R14106 DVSS.n5365 DVSS.n5364 0.4505
R14107 DVSS.n5366 DVSS.n948 0.4505
R14108 DVSS.n5368 DVSS.n5367 0.4505
R14109 DVSS.n946 DVSS.n945 0.4505
R14110 DVSS.n5373 DVSS.n5372 0.4505
R14111 DVSS.n5374 DVSS.n944 0.4505
R14112 DVSS.n5376 DVSS.n5375 0.4505
R14113 DVSS.n942 DVSS.n941 0.4505
R14114 DVSS.n5381 DVSS.n5380 0.4505
R14115 DVSS.n5382 DVSS.n940 0.4505
R14116 DVSS.n5384 DVSS.n5383 0.4505
R14117 DVSS.n938 DVSS.n937 0.4505
R14118 DVSS.n5389 DVSS.n5388 0.4505
R14119 DVSS.n5390 DVSS.n936 0.4505
R14120 DVSS.n5392 DVSS.n5391 0.4505
R14121 DVSS.n934 DVSS.n933 0.4505
R14122 DVSS.n5397 DVSS.n5396 0.4505
R14123 DVSS.n5398 DVSS.n932 0.4505
R14124 DVSS.n5400 DVSS.n5399 0.4505
R14125 DVSS.n930 DVSS.n929 0.4505
R14126 DVSS.n5405 DVSS.n5404 0.4505
R14127 DVSS.n5406 DVSS.n928 0.4505
R14128 DVSS.n5408 DVSS.n5407 0.4505
R14129 DVSS.n926 DVSS.n925 0.4505
R14130 DVSS.n5413 DVSS.n5412 0.4505
R14131 DVSS.n5414 DVSS.n924 0.4505
R14132 DVSS.n5416 DVSS.n5415 0.4505
R14133 DVSS.n922 DVSS.n921 0.4505
R14134 DVSS.n5421 DVSS.n5420 0.4505
R14135 DVSS.n5422 DVSS.n920 0.4505
R14136 DVSS.n5424 DVSS.n5423 0.4505
R14137 DVSS.n918 DVSS.n917 0.4505
R14138 DVSS.n5429 DVSS.n5428 0.4505
R14139 DVSS.n5430 DVSS.n916 0.4505
R14140 DVSS.n5432 DVSS.n5431 0.4505
R14141 DVSS.n914 DVSS.n913 0.4505
R14142 DVSS.n5437 DVSS.n5436 0.4505
R14143 DVSS.n5438 DVSS.n912 0.4505
R14144 DVSS.n5440 DVSS.n5439 0.4505
R14145 DVSS.n910 DVSS.n909 0.4505
R14146 DVSS.n5445 DVSS.n5444 0.4505
R14147 DVSS.n5446 DVSS.n908 0.4505
R14148 DVSS.n5448 DVSS.n5447 0.4505
R14149 DVSS.n906 DVSS.n905 0.4505
R14150 DVSS.n5453 DVSS.n5452 0.4505
R14151 DVSS.n5454 DVSS.n904 0.4505
R14152 DVSS.n5456 DVSS.n5455 0.4505
R14153 DVSS.n902 DVSS.n901 0.4505
R14154 DVSS.n5461 DVSS.n5460 0.4505
R14155 DVSS.n5462 DVSS.n900 0.4505
R14156 DVSS.n5464 DVSS.n5463 0.4505
R14157 DVSS.n898 DVSS.n897 0.4505
R14158 DVSS.n5469 DVSS.n5468 0.4505
R14159 DVSS.n5470 DVSS.n896 0.4505
R14160 DVSS.n5472 DVSS.n5471 0.4505
R14161 DVSS.n894 DVSS.n893 0.4505
R14162 DVSS.n5477 DVSS.n5476 0.4505
R14163 DVSS.n5478 DVSS.n892 0.4505
R14164 DVSS.n5480 DVSS.n5479 0.4505
R14165 DVSS.n890 DVSS.n889 0.4505
R14166 DVSS.n5485 DVSS.n5484 0.4505
R14167 DVSS.n5486 DVSS.n888 0.4505
R14168 DVSS.n5488 DVSS.n5487 0.4505
R14169 DVSS.n886 DVSS.n885 0.4505
R14170 DVSS.n5493 DVSS.n5492 0.4505
R14171 DVSS.n5494 DVSS.n884 0.4505
R14172 DVSS.n5496 DVSS.n5495 0.4505
R14173 DVSS.n882 DVSS.n881 0.4505
R14174 DVSS.n5501 DVSS.n5500 0.4505
R14175 DVSS.n5502 DVSS.n880 0.4505
R14176 DVSS.n5504 DVSS.n5503 0.4505
R14177 DVSS.n878 DVSS.n877 0.4505
R14178 DVSS.n5509 DVSS.n5508 0.4505
R14179 DVSS.n5510 DVSS.n876 0.4505
R14180 DVSS.n5512 DVSS.n5511 0.4505
R14181 DVSS.n874 DVSS.n873 0.4505
R14182 DVSS.n5517 DVSS.n5516 0.4505
R14183 DVSS.n5518 DVSS.n872 0.4505
R14184 DVSS.n5520 DVSS.n5519 0.4505
R14185 DVSS.n870 DVSS.n869 0.4505
R14186 DVSS.n5525 DVSS.n5524 0.4505
R14187 DVSS.n5526 DVSS.n868 0.4505
R14188 DVSS.n5528 DVSS.n5527 0.4505
R14189 DVSS.n866 DVSS.n865 0.4505
R14190 DVSS.n5533 DVSS.n5532 0.4505
R14191 DVSS.n5534 DVSS.n864 0.4505
R14192 DVSS.n5536 DVSS.n5535 0.4505
R14193 DVSS.n862 DVSS.n861 0.4505
R14194 DVSS.n5541 DVSS.n5540 0.4505
R14195 DVSS.n5542 DVSS.n860 0.4505
R14196 DVSS.n5544 DVSS.n5543 0.4505
R14197 DVSS.n858 DVSS.n857 0.4505
R14198 DVSS.n5549 DVSS.n5548 0.4505
R14199 DVSS.n5551 DVSS.n5550 0.4505
R14200 DVSS.n953 DVSS.n951 0.4505
R14201 DVSS.n5362 DVSS.n950 0.4505
R14202 DVSS.n5364 DVSS.n5363 0.4505
R14203 DVSS.n948 DVSS.n947 0.4505
R14204 DVSS.n5369 DVSS.n5368 0.4505
R14205 DVSS.n5370 DVSS.n946 0.4505
R14206 DVSS.n5372 DVSS.n5371 0.4505
R14207 DVSS.n944 DVSS.n943 0.4505
R14208 DVSS.n5377 DVSS.n5376 0.4505
R14209 DVSS.n5378 DVSS.n942 0.4505
R14210 DVSS.n5380 DVSS.n5379 0.4505
R14211 DVSS.n940 DVSS.n939 0.4505
R14212 DVSS.n5385 DVSS.n5384 0.4505
R14213 DVSS.n5386 DVSS.n938 0.4505
R14214 DVSS.n5388 DVSS.n5387 0.4505
R14215 DVSS.n936 DVSS.n935 0.4505
R14216 DVSS.n5393 DVSS.n5392 0.4505
R14217 DVSS.n5394 DVSS.n934 0.4505
R14218 DVSS.n5396 DVSS.n5395 0.4505
R14219 DVSS.n932 DVSS.n931 0.4505
R14220 DVSS.n5401 DVSS.n5400 0.4505
R14221 DVSS.n5402 DVSS.n930 0.4505
R14222 DVSS.n5404 DVSS.n5403 0.4505
R14223 DVSS.n928 DVSS.n927 0.4505
R14224 DVSS.n5409 DVSS.n5408 0.4505
R14225 DVSS.n5410 DVSS.n926 0.4505
R14226 DVSS.n5412 DVSS.n5411 0.4505
R14227 DVSS.n924 DVSS.n923 0.4505
R14228 DVSS.n5417 DVSS.n5416 0.4505
R14229 DVSS.n5418 DVSS.n922 0.4505
R14230 DVSS.n5420 DVSS.n5419 0.4505
R14231 DVSS.n920 DVSS.n919 0.4505
R14232 DVSS.n5425 DVSS.n5424 0.4505
R14233 DVSS.n5426 DVSS.n918 0.4505
R14234 DVSS.n5428 DVSS.n5427 0.4505
R14235 DVSS.n916 DVSS.n915 0.4505
R14236 DVSS.n5433 DVSS.n5432 0.4505
R14237 DVSS.n5434 DVSS.n914 0.4505
R14238 DVSS.n5436 DVSS.n5435 0.4505
R14239 DVSS.n912 DVSS.n911 0.4505
R14240 DVSS.n5441 DVSS.n5440 0.4505
R14241 DVSS.n5442 DVSS.n910 0.4505
R14242 DVSS.n5444 DVSS.n5443 0.4505
R14243 DVSS.n908 DVSS.n907 0.4505
R14244 DVSS.n5449 DVSS.n5448 0.4505
R14245 DVSS.n5450 DVSS.n906 0.4505
R14246 DVSS.n5452 DVSS.n5451 0.4505
R14247 DVSS.n904 DVSS.n903 0.4505
R14248 DVSS.n5457 DVSS.n5456 0.4505
R14249 DVSS.n5458 DVSS.n902 0.4505
R14250 DVSS.n5460 DVSS.n5459 0.4505
R14251 DVSS.n900 DVSS.n899 0.4505
R14252 DVSS.n5465 DVSS.n5464 0.4505
R14253 DVSS.n5466 DVSS.n898 0.4505
R14254 DVSS.n5468 DVSS.n5467 0.4505
R14255 DVSS.n896 DVSS.n895 0.4505
R14256 DVSS.n5473 DVSS.n5472 0.4505
R14257 DVSS.n5474 DVSS.n894 0.4505
R14258 DVSS.n5476 DVSS.n5475 0.4505
R14259 DVSS.n892 DVSS.n891 0.4505
R14260 DVSS.n5481 DVSS.n5480 0.4505
R14261 DVSS.n5482 DVSS.n890 0.4505
R14262 DVSS.n5484 DVSS.n5483 0.4505
R14263 DVSS.n888 DVSS.n887 0.4505
R14264 DVSS.n5489 DVSS.n5488 0.4505
R14265 DVSS.n5490 DVSS.n886 0.4505
R14266 DVSS.n5492 DVSS.n5491 0.4505
R14267 DVSS.n884 DVSS.n883 0.4505
R14268 DVSS.n5497 DVSS.n5496 0.4505
R14269 DVSS.n5498 DVSS.n882 0.4505
R14270 DVSS.n5500 DVSS.n5499 0.4505
R14271 DVSS.n880 DVSS.n879 0.4505
R14272 DVSS.n5505 DVSS.n5504 0.4505
R14273 DVSS.n5506 DVSS.n878 0.4505
R14274 DVSS.n5508 DVSS.n5507 0.4505
R14275 DVSS.n876 DVSS.n875 0.4505
R14276 DVSS.n5513 DVSS.n5512 0.4505
R14277 DVSS.n5514 DVSS.n874 0.4505
R14278 DVSS.n5516 DVSS.n5515 0.4505
R14279 DVSS.n872 DVSS.n871 0.4505
R14280 DVSS.n5521 DVSS.n5520 0.4505
R14281 DVSS.n5522 DVSS.n870 0.4505
R14282 DVSS.n5524 DVSS.n5523 0.4505
R14283 DVSS.n868 DVSS.n867 0.4505
R14284 DVSS.n5529 DVSS.n5528 0.4505
R14285 DVSS.n5530 DVSS.n866 0.4505
R14286 DVSS.n5532 DVSS.n5531 0.4505
R14287 DVSS.n864 DVSS.n863 0.4505
R14288 DVSS.n5537 DVSS.n5536 0.4505
R14289 DVSS.n5538 DVSS.n862 0.4505
R14290 DVSS.n5540 DVSS.n5539 0.4505
R14291 DVSS.n860 DVSS.n859 0.4505
R14292 DVSS.n5545 DVSS.n5544 0.4505
R14293 DVSS.n5546 DVSS.n858 0.4505
R14294 DVSS.n5548 DVSS.n5547 0.4505
R14295 DVSS.n5552 DVSS.n5551 0.4505
R14296 DVSS.n4855 DVSS.n4847 0.4505
R14297 DVSS.n4849 DVSS.n4846 0.4505
R14298 DVSS.n4548 DVSS.n4510 0.4505
R14299 DVSS.n4550 DVSS.n4549 0.4505
R14300 DVSS.n4508 DVSS.n4507 0.4505
R14301 DVSS.n4555 DVSS.n4554 0.4505
R14302 DVSS.n4556 DVSS.n4506 0.4505
R14303 DVSS.n4558 DVSS.n4557 0.4505
R14304 DVSS.n4501 DVSS.n4500 0.4505
R14305 DVSS.n4570 DVSS.n4569 0.4505
R14306 DVSS.n4571 DVSS.n4498 0.4505
R14307 DVSS.n4667 DVSS.n4666 0.4505
R14308 DVSS.n4665 DVSS.n4499 0.4505
R14309 DVSS.n4664 DVSS.n4663 0.4505
R14310 DVSS.n4573 DVSS.n4572 0.4505
R14311 DVSS.n4659 DVSS.n4658 0.4505
R14312 DVSS.n4657 DVSS.n4579 0.4505
R14313 DVSS.n4656 DVSS.n4655 0.4505
R14314 DVSS.n4581 DVSS.n4580 0.4505
R14315 DVSS.n4588 DVSS.n4586 0.4505
R14316 DVSS.n4647 DVSS.n4646 0.4505
R14317 DVSS.n4645 DVSS.n4587 0.4505
R14318 DVSS.n4644 DVSS.n4643 0.4505
R14319 DVSS.n4590 DVSS.n4589 0.4505
R14320 DVSS.n4607 DVSS.n4605 0.4505
R14321 DVSS.n4634 DVSS.n4633 0.4505
R14322 DVSS.n4632 DVSS.n4606 0.4505
R14323 DVSS.n4631 DVSS.n4630 0.4505
R14324 DVSS.n4609 DVSS.n4608 0.4505
R14325 DVSS.n4626 DVSS.n4625 0.4505
R14326 DVSS.n4624 DVSS.n4611 0.4505
R14327 DVSS.n4623 DVSS.n4622 0.4505
R14328 DVSS.n4613 DVSS.n4612 0.4505
R14329 DVSS.n1268 DVSS.n1267 0.4505
R14330 DVSS.n4686 DVSS.n4685 0.4505
R14331 DVSS.n4687 DVSS.n1266 0.4505
R14332 DVSS.n4689 DVSS.n4688 0.4505
R14333 DVSS.n1259 DVSS.n1258 0.4505
R14334 DVSS.n4699 DVSS.n4698 0.4505
R14335 DVSS.n4700 DVSS.n1257 0.4505
R14336 DVSS.n4702 DVSS.n4701 0.4505
R14337 DVSS.n1255 DVSS.n1254 0.4505
R14338 DVSS.n4708 DVSS.n4707 0.4505
R14339 DVSS.n4709 DVSS.n1253 0.4505
R14340 DVSS.n4711 DVSS.n4710 0.4505
R14341 DVSS.n1248 DVSS.n1247 0.4505
R14342 DVSS.n4725 DVSS.n4724 0.4505
R14343 DVSS.n4726 DVSS.n1245 0.4505
R14344 DVSS.n4729 DVSS.n4728 0.4505
R14345 DVSS.n4727 DVSS.n1246 0.4505
R14346 DVSS.n1238 DVSS.n1237 0.4505
R14347 DVSS.n4740 DVSS.n4739 0.4505
R14348 DVSS.n4741 DVSS.n1236 0.4505
R14349 DVSS.n4743 DVSS.n4742 0.4505
R14350 DVSS.n1234 DVSS.n1233 0.4505
R14351 DVSS.n4748 DVSS.n4747 0.4505
R14352 DVSS.n4749 DVSS.n1232 0.4505
R14353 DVSS.n4751 DVSS.n4750 0.4505
R14354 DVSS.n1227 DVSS.n1226 0.4505
R14355 DVSS.n4763 DVSS.n4762 0.4505
R14356 DVSS.n4764 DVSS.n1224 0.4505
R14357 DVSS.n4915 DVSS.n4914 0.4505
R14358 DVSS.n4913 DVSS.n1225 0.4505
R14359 DVSS.n4912 DVSS.n4911 0.4505
R14360 DVSS.n4766 DVSS.n4765 0.4505
R14361 DVSS.n4907 DVSS.n4906 0.4505
R14362 DVSS.n4905 DVSS.n4772 0.4505
R14363 DVSS.n4904 DVSS.n4903 0.4505
R14364 DVSS.n4774 DVSS.n4773 0.4505
R14365 DVSS.n4781 DVSS.n4779 0.4505
R14366 DVSS.n4895 DVSS.n4894 0.4505
R14367 DVSS.n4893 DVSS.n4780 0.4505
R14368 DVSS.n4892 DVSS.n4891 0.4505
R14369 DVSS.n4783 DVSS.n4782 0.4505
R14370 DVSS.n4800 DVSS.n4798 0.4505
R14371 DVSS.n4882 DVSS.n4881 0.4505
R14372 DVSS.n4880 DVSS.n4799 0.4505
R14373 DVSS.n4879 DVSS.n4878 0.4505
R14374 DVSS.n4802 DVSS.n4801 0.4505
R14375 DVSS.n4839 DVSS.n4838 0.4505
R14376 DVSS.n4840 DVSS.n4836 0.4505
R14377 DVSS.n4870 DVSS.n4869 0.4505
R14378 DVSS.n4868 DVSS.n4837 0.4505
R14379 DVSS.n4867 DVSS.n4866 0.4505
R14380 DVSS.n4842 DVSS.n4841 0.4505
R14381 DVSS.n4862 DVSS.n4861 0.4505
R14382 DVSS.n4860 DVSS.n4844 0.4505
R14383 DVSS.n4859 DVSS.n4858 0.4505
R14384 DVSS.n4857 DVSS.n4845 0.4505
R14385 DVSS.n4852 DVSS.n4851 0.4505
R14386 DVSS.n4853 DVSS.n4846 0.4505
R14387 DVSS.n4855 DVSS.n4854 0.4505
R14388 DVSS.n4546 DVSS.n4545 0.4505
R14389 DVSS.n4540 DVSS.n4510 0.4505
R14390 DVSS.n4551 DVSS.n4550 0.4505
R14391 DVSS.n4552 DVSS.n4508 0.4505
R14392 DVSS.n4554 DVSS.n4553 0.4505
R14393 DVSS.n4506 DVSS.n4504 0.4505
R14394 DVSS.n4559 DVSS.n4558 0.4505
R14395 DVSS.n4502 DVSS.n4501 0.4505
R14396 DVSS.n4569 DVSS.n4568 0.4505
R14397 DVSS.n4498 DVSS.n4496 0.4505
R14398 DVSS.n4668 DVSS.n4667 0.4505
R14399 DVSS.n4574 DVSS.n4499 0.4505
R14400 DVSS.n4663 DVSS.n4662 0.4505
R14401 DVSS.n4661 DVSS.n4573 0.4505
R14402 DVSS.n4660 DVSS.n4659 0.4505
R14403 DVSS.n4579 DVSS.n4578 0.4505
R14404 DVSS.n4655 DVSS.n4654 0.4505
R14405 DVSS.n4653 DVSS.n4581 0.4505
R14406 DVSS.n4586 DVSS.n4582 0.4505
R14407 DVSS.n4648 DVSS.n4647 0.4505
R14408 DVSS.n4591 DVSS.n4587 0.4505
R14409 DVSS.n4643 DVSS.n4642 0.4505
R14410 DVSS.n4593 DVSS.n4590 0.4505
R14411 DVSS.n4605 DVSS.n4603 0.4505
R14412 DVSS.n4635 DVSS.n4634 0.4505
R14413 DVSS.n4606 DVSS.n4604 0.4505
R14414 DVSS.n4630 DVSS.n4629 0.4505
R14415 DVSS.n4628 DVSS.n4609 0.4505
R14416 DVSS.n4627 DVSS.n4626 0.4505
R14417 DVSS.n4611 DVSS.n4610 0.4505
R14418 DVSS.n4622 DVSS.n4621 0.4505
R14419 DVSS.n4614 DVSS.n4613 0.4505
R14420 DVSS.n4616 DVSS.n1268 0.4505
R14421 DVSS.n4685 DVSS.n4684 0.4505
R14422 DVSS.n1266 DVSS.n1264 0.4505
R14423 DVSS.n4690 DVSS.n4689 0.4505
R14424 DVSS.n1260 DVSS.n1259 0.4505
R14425 DVSS.n4698 DVSS.n4697 0.4505
R14426 DVSS.n1257 DVSS.n1256 0.4505
R14427 DVSS.n4703 DVSS.n4702 0.4505
R14428 DVSS.n4704 DVSS.n1255 0.4505
R14429 DVSS.n4707 DVSS.n4706 0.4505
R14430 DVSS.n4705 DVSS.n1253 0.4505
R14431 DVSS.n4712 DVSS.n4711 0.4505
R14432 DVSS.n4713 DVSS.n1248 0.4505
R14433 DVSS.n4724 DVSS.n4723 0.4505
R14434 DVSS.n1245 DVSS.n1243 0.4505
R14435 DVSS.n4730 DVSS.n4729 0.4505
R14436 DVSS.n1246 DVSS.n1239 0.4505
R14437 DVSS.n4737 DVSS.n1238 0.4505
R14438 DVSS.n4739 DVSS.n4738 0.4505
R14439 DVSS.n1236 DVSS.n1235 0.4505
R14440 DVSS.n4744 DVSS.n4743 0.4505
R14441 DVSS.n4745 DVSS.n1234 0.4505
R14442 DVSS.n4747 DVSS.n4746 0.4505
R14443 DVSS.n1232 DVSS.n1230 0.4505
R14444 DVSS.n4752 DVSS.n4751 0.4505
R14445 DVSS.n1228 DVSS.n1227 0.4505
R14446 DVSS.n4762 DVSS.n4761 0.4505
R14447 DVSS.n1224 DVSS.n1222 0.4505
R14448 DVSS.n4916 DVSS.n4915 0.4505
R14449 DVSS.n4767 DVSS.n1225 0.4505
R14450 DVSS.n4911 DVSS.n4910 0.4505
R14451 DVSS.n4909 DVSS.n4766 0.4505
R14452 DVSS.n4908 DVSS.n4907 0.4505
R14453 DVSS.n4772 DVSS.n4771 0.4505
R14454 DVSS.n4903 DVSS.n4902 0.4505
R14455 DVSS.n4901 DVSS.n4774 0.4505
R14456 DVSS.n4779 DVSS.n4775 0.4505
R14457 DVSS.n4896 DVSS.n4895 0.4505
R14458 DVSS.n4784 DVSS.n4780 0.4505
R14459 DVSS.n4891 DVSS.n4890 0.4505
R14460 DVSS.n4786 DVSS.n4783 0.4505
R14461 DVSS.n4798 DVSS.n4796 0.4505
R14462 DVSS.n4883 DVSS.n4882 0.4505
R14463 DVSS.n4799 DVSS.n4797 0.4505
R14464 DVSS.n4878 DVSS.n4877 0.4505
R14465 DVSS.n4876 DVSS.n4802 0.4505
R14466 DVSS.n4838 DVSS.n4808 0.4505
R14467 DVSS.n4836 DVSS.n4831 0.4505
R14468 DVSS.n4871 DVSS.n4870 0.4505
R14469 DVSS.n4837 DVSS.n4835 0.4505
R14470 DVSS.n4866 DVSS.n4865 0.4505
R14471 DVSS.n4864 DVSS.n4842 0.4505
R14472 DVSS.n4863 DVSS.n4862 0.4505
R14473 DVSS.n4844 DVSS.n4843 0.4505
R14474 DVSS.n4858 DVSS.n1181 0.4505
R14475 DVSS.n4857 DVSS.n4856 0.4505
R14476 DVSS.n2652 DVSS.n2651 0.4505
R14477 DVSS.n2268 DVSS.n2267 0.4505
R14478 DVSS.n2633 DVSS.n2632 0.4505
R14479 DVSS.n2635 DVSS.n2634 0.4505
R14480 DVSS.n2631 DVSS.n2426 0.4505
R14481 DVSS.n2630 DVSS.n2629 0.4505
R14482 DVSS.n2428 DVSS.n2427 0.4505
R14483 DVSS.n2625 DVSS.n2624 0.4505
R14484 DVSS.n2623 DVSS.n2430 0.4505
R14485 DVSS.n2622 DVSS.n2621 0.4505
R14486 DVSS.n2432 DVSS.n2431 0.4505
R14487 DVSS.n2617 DVSS.n2616 0.4505
R14488 DVSS.n2615 DVSS.n2434 0.4505
R14489 DVSS.n2614 DVSS.n2613 0.4505
R14490 DVSS.n2436 DVSS.n2435 0.4505
R14491 DVSS.n2609 DVSS.n2608 0.4505
R14492 DVSS.n2607 DVSS.n2438 0.4505
R14493 DVSS.n2606 DVSS.n2605 0.4505
R14494 DVSS.n2440 DVSS.n2439 0.4505
R14495 DVSS.n2601 DVSS.n2600 0.4505
R14496 DVSS.n2599 DVSS.n2442 0.4505
R14497 DVSS.n2598 DVSS.n2597 0.4505
R14498 DVSS.n2444 DVSS.n2443 0.4505
R14499 DVSS.n2593 DVSS.n2592 0.4505
R14500 DVSS.n2591 DVSS.n2446 0.4505
R14501 DVSS.n2590 DVSS.n2589 0.4505
R14502 DVSS.n2448 DVSS.n2447 0.4505
R14503 DVSS.n2585 DVSS.n2584 0.4505
R14504 DVSS.n2583 DVSS.n2450 0.4505
R14505 DVSS.n2582 DVSS.n2581 0.4505
R14506 DVSS.n2452 DVSS.n2451 0.4505
R14507 DVSS.n2577 DVSS.n2576 0.4505
R14508 DVSS.n2575 DVSS.n2454 0.4505
R14509 DVSS.n2574 DVSS.n2573 0.4505
R14510 DVSS.n2456 DVSS.n2455 0.4505
R14511 DVSS.n2569 DVSS.n2568 0.4505
R14512 DVSS.n2567 DVSS.n2458 0.4505
R14513 DVSS.n2566 DVSS.n2565 0.4505
R14514 DVSS.n2460 DVSS.n2459 0.4505
R14515 DVSS.n2561 DVSS.n2560 0.4505
R14516 DVSS.n2559 DVSS.n2462 0.4505
R14517 DVSS.n2558 DVSS.n2557 0.4505
R14518 DVSS.n2464 DVSS.n2463 0.4505
R14519 DVSS.n2553 DVSS.n2552 0.4505
R14520 DVSS.n2551 DVSS.n2466 0.4505
R14521 DVSS.n2550 DVSS.n2549 0.4505
R14522 DVSS.n2468 DVSS.n2467 0.4505
R14523 DVSS.n2545 DVSS.n2544 0.4505
R14524 DVSS.n2543 DVSS.n2470 0.4505
R14525 DVSS.n2542 DVSS.n2541 0.4505
R14526 DVSS.n2472 DVSS.n2471 0.4505
R14527 DVSS.n2537 DVSS.n2536 0.4505
R14528 DVSS.n2535 DVSS.n2474 0.4505
R14529 DVSS.n2534 DVSS.n2533 0.4505
R14530 DVSS.n2476 DVSS.n2475 0.4505
R14531 DVSS.n2529 DVSS.n2528 0.4505
R14532 DVSS.n2527 DVSS.n2478 0.4505
R14533 DVSS.n2526 DVSS.n2525 0.4505
R14534 DVSS.n2480 DVSS.n2479 0.4505
R14535 DVSS.n2521 DVSS.n2520 0.4505
R14536 DVSS.n2519 DVSS.n2482 0.4505
R14537 DVSS.n2518 DVSS.n2517 0.4505
R14538 DVSS.n2484 DVSS.n2483 0.4505
R14539 DVSS.n2513 DVSS.n2512 0.4505
R14540 DVSS.n2511 DVSS.n2486 0.4505
R14541 DVSS.n2510 DVSS.n2509 0.4505
R14542 DVSS.n2488 DVSS.n2487 0.4505
R14543 DVSS.n2505 DVSS.n2504 0.4505
R14544 DVSS.n2503 DVSS.n2490 0.4505
R14545 DVSS.n2502 DVSS.n2501 0.4505
R14546 DVSS.n2492 DVSS.n2491 0.4505
R14547 DVSS.n2497 DVSS.n2496 0.4505
R14548 DVSS.n2495 DVSS.n2494 0.4505
R14549 DVSS.n1533 DVSS.n1532 0.4505
R14550 DVSS.n1541 DVSS.n1540 0.4505
R14551 DVSS.n1542 DVSS.n1531 0.4505
R14552 DVSS.n1544 DVSS.n1543 0.4505
R14553 DVSS.n1529 DVSS.n1528 0.4505
R14554 DVSS.n1549 DVSS.n1548 0.4505
R14555 DVSS.n1550 DVSS.n1527 0.4505
R14556 DVSS.n1552 DVSS.n1551 0.4505
R14557 DVSS.n1525 DVSS.n1524 0.4505
R14558 DVSS.n1557 DVSS.n1556 0.4505
R14559 DVSS.n1558 DVSS.n1522 0.4505
R14560 DVSS.n3935 DVSS.n3934 0.4505
R14561 DVSS.n3933 DVSS.n1523 0.4505
R14562 DVSS.n3932 DVSS.n3931 0.4505
R14563 DVSS.n1560 DVSS.n1559 0.4505
R14564 DVSS.n3927 DVSS.n3926 0.4505
R14565 DVSS.n3925 DVSS.n1562 0.4505
R14566 DVSS.n3924 DVSS.n3923 0.4505
R14567 DVSS.n1564 DVSS.n1563 0.4505
R14568 DVSS.n3919 DVSS.n3918 0.4505
R14569 DVSS.n3917 DVSS.n1566 0.4505
R14570 DVSS.n3916 DVSS.n3915 0.4505
R14571 DVSS.n1568 DVSS.n1567 0.4505
R14572 DVSS.n3911 DVSS.n3910 0.4505
R14573 DVSS.n3909 DVSS.n1570 0.4505
R14574 DVSS.n3908 DVSS.n3907 0.4505
R14575 DVSS.n1572 DVSS.n1571 0.4505
R14576 DVSS.n3563 DVSS.n3562 0.4505
R14577 DVSS.n3826 DVSS.n1634 0.4505
R14578 DVSS.n3727 DVSS.n3726 0.4505
R14579 DVSS.n3731 DVSS.n3730 0.4505
R14580 DVSS.n3732 DVSS.n3725 0.4505
R14581 DVSS.n3734 DVSS.n3733 0.4505
R14582 DVSS.n3723 DVSS.n3722 0.4505
R14583 DVSS.n3739 DVSS.n3738 0.4505
R14584 DVSS.n3740 DVSS.n3657 0.4505
R14585 DVSS.n3742 DVSS.n3741 0.4505
R14586 DVSS.n3721 DVSS.n3656 0.4505
R14587 DVSS.n3720 DVSS.n3719 0.4505
R14588 DVSS.n3659 DVSS.n3658 0.4505
R14589 DVSS.n3715 DVSS.n3714 0.4505
R14590 DVSS.n3713 DVSS.n3661 0.4505
R14591 DVSS.n3712 DVSS.n3711 0.4505
R14592 DVSS.n3663 DVSS.n3662 0.4505
R14593 DVSS.n3707 DVSS.n3706 0.4505
R14594 DVSS.n3705 DVSS.n3665 0.4505
R14595 DVSS.n3704 DVSS.n3703 0.4505
R14596 DVSS.n3667 DVSS.n3666 0.4505
R14597 DVSS.n3699 DVSS.n3698 0.4505
R14598 DVSS.n3697 DVSS.n3669 0.4505
R14599 DVSS.n3696 DVSS.n3695 0.4505
R14600 DVSS.n3671 DVSS.n3670 0.4505
R14601 DVSS.n3691 DVSS.n3690 0.4505
R14602 DVSS.n3689 DVSS.n3673 0.4505
R14603 DVSS.n3688 DVSS.n3687 0.4505
R14604 DVSS.n3675 DVSS.n3674 0.4505
R14605 DVSS.n3683 DVSS.n3682 0.4505
R14606 DVSS.n3681 DVSS.n3678 0.4505
R14607 DVSS.n3680 DVSS.n3679 0.4505
R14608 DVSS.n1685 DVSS.n1684 0.4505
R14609 DVSS.n3774 DVSS.n3773 0.4505
R14610 DVSS.n3775 DVSS.n1683 0.4505
R14611 DVSS.n3777 DVSS.n3776 0.4505
R14612 DVSS.n1680 DVSS.n1679 0.4505
R14613 DVSS.n3782 DVSS.n3781 0.4505
R14614 DVSS.n3783 DVSS.n1664 0.4505
R14615 DVSS.n3785 DVSS.n3784 0.4505
R14616 DVSS.n1678 DVSS.n1663 0.4505
R14617 DVSS.n1677 DVSS.n1676 0.4505
R14618 DVSS.n1666 DVSS.n1665 0.4505
R14619 DVSS.n1668 DVSS.n1667 0.4505
R14620 DVSS.n1652 DVSS.n1651 0.4505
R14621 DVSS.n3797 DVSS.n3796 0.4505
R14622 DVSS.n3798 DVSS.n1650 0.4505
R14623 DVSS.n3800 DVSS.n3799 0.4505
R14624 DVSS.n1646 DVSS.n1645 0.4505
R14625 DVSS.n3806 DVSS.n3805 0.4505
R14626 DVSS.n3807 DVSS.n1644 0.4505
R14627 DVSS.n3809 DVSS.n3808 0.4505
R14628 DVSS.n1642 DVSS.n1641 0.4505
R14629 DVSS.n3814 DVSS.n3813 0.4505
R14630 DVSS.n3815 DVSS.n1640 0.4505
R14631 DVSS.n3817 DVSS.n3816 0.4505
R14632 DVSS.n1637 DVSS.n1636 0.4505
R14633 DVSS.n3822 DVSS.n3821 0.4505
R14634 DVSS.n3823 DVSS.n1635 0.4505
R14635 DVSS.n3825 DVSS.n3824 0.4505
R14636 DVSS.n1598 DVSS.n1592 0.4505
R14637 DVSS.n3892 DVSS.n3891 0.4505
R14638 DVSS.n3890 DVSS.n1593 0.4505
R14639 DVSS.n3889 DVSS.n3888 0.4505
R14640 DVSS.n1600 DVSS.n1599 0.4505
R14641 DVSS.n3883 DVSS.n3882 0.4505
R14642 DVSS.n3881 DVSS.n1602 0.4505
R14643 DVSS.n3880 DVSS.n3879 0.4505
R14644 DVSS.n1604 DVSS.n1603 0.4505
R14645 DVSS.n3873 DVSS.n3872 0.4505
R14646 DVSS.n3871 DVSS.n1606 0.4505
R14647 DVSS.n3870 DVSS.n3869 0.4505
R14648 DVSS.n1608 DVSS.n1607 0.4505
R14649 DVSS.n3865 DVSS.n3864 0.4505
R14650 DVSS.n3863 DVSS.n1611 0.4505
R14651 DVSS.n3862 DVSS.n3861 0.4505
R14652 DVSS.n1613 DVSS.n1612 0.4505
R14653 DVSS.n3854 DVSS.n3853 0.4505
R14654 DVSS.n3852 DVSS.n1616 0.4505
R14655 DVSS.n3851 DVSS.n3850 0.4505
R14656 DVSS.n1618 DVSS.n1617 0.4505
R14657 DVSS.n3846 DVSS.n3845 0.4505
R14658 DVSS.n3844 DVSS.n1621 0.4505
R14659 DVSS.n3843 DVSS.n3842 0.4505
R14660 DVSS.n1623 DVSS.n1622 0.4505
R14661 DVSS.n1743 DVSS.n1742 0.4505
R14662 DVSS.n1895 DVSS.n1894 0.4505
R14663 DVSS.n1897 DVSS.n1896 0.4505
R14664 DVSS.n1887 DVSS.n1886 0.4505
R14665 DVSS.n1904 DVSS.n1903 0.4505
R14666 DVSS.n1905 DVSS.n1885 0.4505
R14667 DVSS.n1907 DVSS.n1906 0.4505
R14668 DVSS.n1766 DVSS.n1764 0.4505
R14669 DVSS.n2194 DVSS.n2193 0.4505
R14670 DVSS.n2192 DVSS.n1765 0.4505
R14671 DVSS.n2191 DVSS.n2190 0.4505
R14672 DVSS.n1768 DVSS.n1767 0.4505
R14673 DVSS.n1872 DVSS.n1871 0.4505
R14674 DVSS.n1793 DVSS.n1791 0.4505
R14675 DVSS.n2176 DVSS.n2175 0.4505
R14676 DVSS.n2174 DVSS.n1792 0.4505
R14677 DVSS.n2173 DVSS.n2172 0.4505
R14678 DVSS.n1795 DVSS.n1794 0.4505
R14679 DVSS.n2143 DVSS.n2142 0.4505
R14680 DVSS.n2141 DVSS.n1927 0.4505
R14681 DVSS.n2140 DVSS.n2139 0.4505
R14682 DVSS.n1929 DVSS.n1928 0.4505
R14683 DVSS.n1969 DVSS.n1968 0.4505
R14684 DVSS.n1970 DVSS.n1967 0.4505
R14685 DVSS.n1972 DVSS.n1971 0.4505
R14686 DVSS.n1957 DVSS.n1956 0.4505
R14687 DVSS.n1987 DVSS.n1986 0.4505
R14688 DVSS.n1988 DVSS.n1954 0.4505
R14689 DVSS.n2122 DVSS.n2121 0.4505
R14690 DVSS.n2120 DVSS.n1955 0.4505
R14691 DVSS.n2119 DVSS.n2118 0.4505
R14692 DVSS.n2083 DVSS.n1989 0.4505
R14693 DVSS.n2082 DVSS.n1991 0.4505
R14694 DVSS.n1994 DVSS.n1990 0.4505
R14695 DVSS.n2078 DVSS.n2077 0.4505
R14696 DVSS.n2076 DVSS.n1993 0.4505
R14697 DVSS.n2075 DVSS.n2074 0.4505
R14698 DVSS.n1996 DVSS.n1995 0.4505
R14699 DVSS.n2070 DVSS.n2069 0.4505
R14700 DVSS.n2068 DVSS.n1998 0.4505
R14701 DVSS.n2067 DVSS.n2066 0.4505
R14702 DVSS.n2000 DVSS.n1999 0.4505
R14703 DVSS.n2062 DVSS.n2061 0.4505
R14704 DVSS.n2060 DVSS.n2002 0.4505
R14705 DVSS.n2059 DVSS.n2058 0.4505
R14706 DVSS.n2004 DVSS.n2003 0.4505
R14707 DVSS.n2054 DVSS.n2053 0.4505
R14708 DVSS.n2052 DVSS.n2006 0.4505
R14709 DVSS.n2051 DVSS.n2050 0.4505
R14710 DVSS.n2008 DVSS.n2007 0.4505
R14711 DVSS.n2046 DVSS.n2045 0.4505
R14712 DVSS.n2044 DVSS.n2010 0.4505
R14713 DVSS.n2043 DVSS.n2042 0.4505
R14714 DVSS.n2012 DVSS.n2011 0.4505
R14715 DVSS.n2038 DVSS.n2037 0.4505
R14716 DVSS.n2036 DVSS.n2014 0.4505
R14717 DVSS.n2035 DVSS.n2034 0.4505
R14718 DVSS.n2016 DVSS.n2015 0.4505
R14719 DVSS.n2030 DVSS.n2029 0.4505
R14720 DVSS.n2028 DVSS.n2018 0.4505
R14721 DVSS.n2027 DVSS.n2026 0.4505
R14722 DVSS.n2020 DVSS.n2019 0.4505
R14723 DVSS.n2022 DVSS.n2021 0.4505
R14724 DVSS.n2225 DVSS.n2224 0.4505
R14725 DVSS.n2223 DVSS.n1736 0.4505
R14726 DVSS.n2222 DVSS.n2221 0.4505
R14727 DVSS.n1738 DVSS.n1737 0.4505
R14728 DVSS.n2217 DVSS.n2216 0.4505
R14729 DVSS.n2215 DVSS.n1741 0.4505
R14730 DVSS.n2214 DVSS.n2213 0.4505
R14731 DVSS.n4036 DVSS.n4035 0.4505
R14732 DVSS.n4040 DVSS.n4039 0.4505
R14733 DVSS.n4041 DVSS.n4034 0.4505
R14734 DVSS.n4043 DVSS.n4042 0.4505
R14735 DVSS.n4032 DVSS.n4031 0.4505
R14736 DVSS.n4048 DVSS.n4047 0.4505
R14737 DVSS.n4049 DVSS.n4030 0.4505
R14738 DVSS.n4051 DVSS.n4050 0.4505
R14739 DVSS.n4028 DVSS.n4027 0.4505
R14740 DVSS.n4056 DVSS.n4055 0.4505
R14741 DVSS.n4057 DVSS.n4026 0.4505
R14742 DVSS.n4059 DVSS.n4058 0.4505
R14743 DVSS.n4024 DVSS.n4023 0.4505
R14744 DVSS.n4064 DVSS.n4063 0.4505
R14745 DVSS.n4065 DVSS.n4022 0.4505
R14746 DVSS.n4067 DVSS.n4066 0.4505
R14747 DVSS.n4020 DVSS.n4019 0.4505
R14748 DVSS.n4072 DVSS.n4071 0.4505
R14749 DVSS.n4073 DVSS.n4018 0.4505
R14750 DVSS.n4075 DVSS.n4074 0.4505
R14751 DVSS.n4016 DVSS.n4015 0.4505
R14752 DVSS.n4080 DVSS.n4079 0.4505
R14753 DVSS.n4081 DVSS.n4014 0.4505
R14754 DVSS.n4083 DVSS.n4082 0.4505
R14755 DVSS.n4012 DVSS.n4011 0.4505
R14756 DVSS.n4088 DVSS.n4087 0.4505
R14757 DVSS.n4089 DVSS.n4007 0.4505
R14758 DVSS.n4180 DVSS.n1372 0.4505
R14759 DVSS.n1375 DVSS.n1371 0.4505
R14760 DVSS.n4176 DVSS.n4175 0.4505
R14761 DVSS.n4174 DVSS.n1374 0.4505
R14762 DVSS.n4173 DVSS.n4172 0.4505
R14763 DVSS.n1377 DVSS.n1376 0.4505
R14764 DVSS.n4166 DVSS.n4165 0.4505
R14765 DVSS.n4164 DVSS.n1392 0.4505
R14766 DVSS.n4163 DVSS.n4162 0.4505
R14767 DVSS.n1394 DVSS.n1393 0.4505
R14768 DVSS.n4158 DVSS.n4157 0.4505
R14769 DVSS.n4156 DVSS.n1396 0.4505
R14770 DVSS.n4155 DVSS.n4154 0.4505
R14771 DVSS.n1398 DVSS.n1397 0.4505
R14772 DVSS.n4150 DVSS.n4149 0.4505
R14773 DVSS.n4148 DVSS.n1400 0.4505
R14774 DVSS.n4147 DVSS.n4146 0.4505
R14775 DVSS.n1402 DVSS.n1401 0.4505
R14776 DVSS.n4142 DVSS.n4141 0.4505
R14777 DVSS.n4140 DVSS.n1404 0.4505
R14778 DVSS.n4139 DVSS.n4138 0.4505
R14779 DVSS.n1406 DVSS.n1405 0.4505
R14780 DVSS.n4134 DVSS.n4133 0.4505
R14781 DVSS.n4132 DVSS.n1408 0.4505
R14782 DVSS.n4131 DVSS.n4130 0.4505
R14783 DVSS.n1410 DVSS.n1409 0.4505
R14784 DVSS.n4126 DVSS.n4125 0.4505
R14785 DVSS.n4124 DVSS.n1412 0.4505
R14786 DVSS.n4123 DVSS.n4122 0.4505
R14787 DVSS.n1414 DVSS.n1413 0.4505
R14788 DVSS.n4118 DVSS.n4117 0.4505
R14789 DVSS.n4116 DVSS.n1416 0.4505
R14790 DVSS.n4115 DVSS.n4114 0.4505
R14791 DVSS.n1418 DVSS.n1417 0.4505
R14792 DVSS.n4110 DVSS.n4109 0.4505
R14793 DVSS.n4108 DVSS.n1420 0.4505
R14794 DVSS.n4107 DVSS.n4106 0.4505
R14795 DVSS.n1422 DVSS.n1421 0.4505
R14796 DVSS.n4102 DVSS.n4101 0.4505
R14797 DVSS.n4100 DVSS.n1424 0.4505
R14798 DVSS.n4099 DVSS.n4098 0.4505
R14799 DVSS.n1426 DVSS.n1425 0.4505
R14800 DVSS.n4009 DVSS.n4008 0.4505
R14801 DVSS.n4010 DVSS.n4006 0.4505
R14802 DVSS.n4091 DVSS.n4090 0.4505
R14803 DVSS.n4007 DVSS.n4005 0.4505
R14804 DVSS.n4182 DVSS.n4181 0.4505
R14805 DVSS.n4087 DVSS.n4086 0.4505
R14806 DVSS.n4085 DVSS.n4012 0.4505
R14807 DVSS.n4084 DVSS.n4083 0.4505
R14808 DVSS.n4014 DVSS.n4013 0.4505
R14809 DVSS.n4079 DVSS.n4078 0.4505
R14810 DVSS.n4077 DVSS.n4016 0.4505
R14811 DVSS.n4076 DVSS.n4075 0.4505
R14812 DVSS.n4018 DVSS.n4017 0.4505
R14813 DVSS.n4071 DVSS.n4070 0.4505
R14814 DVSS.n4069 DVSS.n4020 0.4505
R14815 DVSS.n4068 DVSS.n4067 0.4505
R14816 DVSS.n4022 DVSS.n4021 0.4505
R14817 DVSS.n4063 DVSS.n4062 0.4505
R14818 DVSS.n4061 DVSS.n4024 0.4505
R14819 DVSS.n4060 DVSS.n4059 0.4505
R14820 DVSS.n4026 DVSS.n4025 0.4505
R14821 DVSS.n4055 DVSS.n4054 0.4505
R14822 DVSS.n4053 DVSS.n4028 0.4505
R14823 DVSS.n4052 DVSS.n4051 0.4505
R14824 DVSS.n4030 DVSS.n4029 0.4505
R14825 DVSS.n4047 DVSS.n4046 0.4505
R14826 DVSS.n4045 DVSS.n4032 0.4505
R14827 DVSS.n4044 DVSS.n4043 0.4505
R14828 DVSS.n4034 DVSS.n4033 0.4505
R14829 DVSS.n4039 DVSS.n4038 0.4505
R14830 DVSS.n4180 DVSS.n4179 0.4505
R14831 DVSS.n4178 DVSS.n1371 0.4505
R14832 DVSS.n4177 DVSS.n4176 0.4505
R14833 DVSS.n1374 DVSS.n1373 0.4505
R14834 DVSS.n4172 DVSS.n4171 0.4505
R14835 DVSS.n1384 DVSS.n1377 0.4505
R14836 DVSS.n4167 DVSS.n4166 0.4505
R14837 DVSS.n1392 DVSS.n1391 0.4505
R14838 DVSS.n4162 DVSS.n4161 0.4505
R14839 DVSS.n4160 DVSS.n1394 0.4505
R14840 DVSS.n4159 DVSS.n4158 0.4505
R14841 DVSS.n1396 DVSS.n1395 0.4505
R14842 DVSS.n4154 DVSS.n4153 0.4505
R14843 DVSS.n4152 DVSS.n1398 0.4505
R14844 DVSS.n4151 DVSS.n4150 0.4505
R14845 DVSS.n1400 DVSS.n1399 0.4505
R14846 DVSS.n4146 DVSS.n4145 0.4505
R14847 DVSS.n4144 DVSS.n1402 0.4505
R14848 DVSS.n4143 DVSS.n4142 0.4505
R14849 DVSS.n1404 DVSS.n1403 0.4505
R14850 DVSS.n4138 DVSS.n4137 0.4505
R14851 DVSS.n4136 DVSS.n1406 0.4505
R14852 DVSS.n4135 DVSS.n4134 0.4505
R14853 DVSS.n1408 DVSS.n1407 0.4505
R14854 DVSS.n4130 DVSS.n4129 0.4505
R14855 DVSS.n4128 DVSS.n1410 0.4505
R14856 DVSS.n4127 DVSS.n4126 0.4505
R14857 DVSS.n1412 DVSS.n1411 0.4505
R14858 DVSS.n4122 DVSS.n4121 0.4505
R14859 DVSS.n4120 DVSS.n1414 0.4505
R14860 DVSS.n4119 DVSS.n4118 0.4505
R14861 DVSS.n1416 DVSS.n1415 0.4505
R14862 DVSS.n4114 DVSS.n4113 0.4505
R14863 DVSS.n4112 DVSS.n1418 0.4505
R14864 DVSS.n4111 DVSS.n4110 0.4505
R14865 DVSS.n1420 DVSS.n1419 0.4505
R14866 DVSS.n4106 DVSS.n4105 0.4505
R14867 DVSS.n4104 DVSS.n1422 0.4505
R14868 DVSS.n4103 DVSS.n4102 0.4505
R14869 DVSS.n1424 DVSS.n1423 0.4505
R14870 DVSS.n4098 DVSS.n4097 0.4505
R14871 DVSS.n4096 DVSS.n1426 0.4505
R14872 DVSS.n4008 DVSS.n1431 0.4505
R14873 DVSS.n4006 DVSS.n4004 0.4505
R14874 DVSS.n4092 DVSS.n4091 0.4505
R14875 DVSS.n2024 DVSS.n2020 0.4505
R14876 DVSS.n2026 DVSS.n2025 0.4505
R14877 DVSS.n2018 DVSS.n2017 0.4505
R14878 DVSS.n2031 DVSS.n2030 0.4505
R14879 DVSS.n2032 DVSS.n2016 0.4505
R14880 DVSS.n2034 DVSS.n2033 0.4505
R14881 DVSS.n2014 DVSS.n2013 0.4505
R14882 DVSS.n2039 DVSS.n2038 0.4505
R14883 DVSS.n2040 DVSS.n2012 0.4505
R14884 DVSS.n2042 DVSS.n2041 0.4505
R14885 DVSS.n2010 DVSS.n2009 0.4505
R14886 DVSS.n2047 DVSS.n2046 0.4505
R14887 DVSS.n2048 DVSS.n2008 0.4505
R14888 DVSS.n2050 DVSS.n2049 0.4505
R14889 DVSS.n2006 DVSS.n2005 0.4505
R14890 DVSS.n2055 DVSS.n2054 0.4505
R14891 DVSS.n2056 DVSS.n2004 0.4505
R14892 DVSS.n2058 DVSS.n2057 0.4505
R14893 DVSS.n2002 DVSS.n2001 0.4505
R14894 DVSS.n2063 DVSS.n2062 0.4505
R14895 DVSS.n2064 DVSS.n2000 0.4505
R14896 DVSS.n2066 DVSS.n2065 0.4505
R14897 DVSS.n1998 DVSS.n1997 0.4505
R14898 DVSS.n2071 DVSS.n2070 0.4505
R14899 DVSS.n2072 DVSS.n1996 0.4505
R14900 DVSS.n2074 DVSS.n2073 0.4505
R14901 DVSS.n1993 DVSS.n1992 0.4505
R14902 DVSS.n2079 DVSS.n2078 0.4505
R14903 DVSS.n2080 DVSS.n1990 0.4505
R14904 DVSS.n2082 DVSS.n2081 0.4505
R14905 DVSS.n2087 DVSS.n2083 0.4505
R14906 DVSS.n2118 DVSS.n2117 0.4505
R14907 DVSS.n2084 DVSS.n1955 0.4505
R14908 DVSS.n2123 DVSS.n2122 0.4505
R14909 DVSS.n1954 DVSS.n1952 0.4505
R14910 DVSS.n1986 DVSS.n1985 0.4505
R14911 DVSS.n1958 DVSS.n1957 0.4505
R14912 DVSS.n1973 DVSS.n1972 0.4505
R14913 DVSS.n1967 DVSS.n1966 0.4505
R14914 DVSS.n1968 DVSS.n1963 0.4505
R14915 DVSS.n1932 DVSS.n1929 0.4505
R14916 DVSS.n2139 DVSS.n2138 0.4505
R14917 DVSS.n1930 DVSS.n1927 0.4505
R14918 DVSS.n2144 DVSS.n2143 0.4505
R14919 DVSS.n1798 DVSS.n1795 0.4505
R14920 DVSS.n2172 DVSS.n2171 0.4505
R14921 DVSS.n1792 DVSS.n1790 0.4505
R14922 DVSS.n2177 DVSS.n2176 0.4505
R14923 DVSS.n1791 DVSS.n1789 0.4505
R14924 DVSS.n1873 DVSS.n1872 0.4505
R14925 DVSS.n1771 DVSS.n1768 0.4505
R14926 DVSS.n2190 DVSS.n2189 0.4505
R14927 DVSS.n1769 DVSS.n1765 0.4505
R14928 DVSS.n2195 DVSS.n2194 0.4505
R14929 DVSS.n1764 DVSS.n1762 0.4505
R14930 DVSS.n1908 DVSS.n1907 0.4505
R14931 DVSS.n1885 DVSS.n1884 0.4505
R14932 DVSS.n1745 DVSS.n1743 0.4505
R14933 DVSS.n1894 DVSS.n1893 0.4505
R14934 DVSS.n1898 DVSS.n1897 0.4505
R14935 DVSS.n1888 DVSS.n1887 0.4505
R14936 DVSS.n1903 DVSS.n1902 0.4505
R14937 DVSS.n2227 DVSS.n2226 0.4505
R14938 DVSS.n2225 DVSS.n1735 0.4505
R14939 DVSS.n1739 DVSS.n1736 0.4505
R14940 DVSS.n2221 DVSS.n2220 0.4505
R14941 DVSS.n2219 DVSS.n1738 0.4505
R14942 DVSS.n2218 DVSS.n2217 0.4505
R14943 DVSS.n1822 DVSS.n1741 0.4505
R14944 DVSS.n2213 DVSS.n2212 0.4505
R14945 DVSS.n1663 DVSS.n1661 0.4505
R14946 DVSS.n3801 DVSS.n3800 0.4505
R14947 DVSS.n1650 DVSS.n1649 0.4505
R14948 DVSS.n3796 DVSS.n3795 0.4505
R14949 DVSS.n1653 DVSS.n1652 0.4505
R14950 DVSS.n1669 DVSS.n1668 0.4505
R14951 DVSS.n1670 DVSS.n1666 0.4505
R14952 DVSS.n1676 DVSS.n1675 0.4505
R14953 DVSS.n3786 DVSS.n3785 0.4505
R14954 DVSS.n1681 DVSS.n1664 0.4505
R14955 DVSS.n3781 DVSS.n3780 0.4505
R14956 DVSS.n3779 DVSS.n1680 0.4505
R14957 DVSS.n3778 DVSS.n3777 0.4505
R14958 DVSS.n1686 DVSS.n1683 0.4505
R14959 DVSS.n3773 DVSS.n3772 0.4505
R14960 DVSS.n3771 DVSS.n1685 0.4505
R14961 DVSS.n3679 DVSS.n1687 0.4505
R14962 DVSS.n3678 DVSS.n3677 0.4505
R14963 DVSS.n3684 DVSS.n3683 0.4505
R14964 DVSS.n3685 DVSS.n3675 0.4505
R14965 DVSS.n3687 DVSS.n3686 0.4505
R14966 DVSS.n3673 DVSS.n3672 0.4505
R14967 DVSS.n3692 DVSS.n3691 0.4505
R14968 DVSS.n3693 DVSS.n3671 0.4505
R14969 DVSS.n3695 DVSS.n3694 0.4505
R14970 DVSS.n3669 DVSS.n3668 0.4505
R14971 DVSS.n3700 DVSS.n3699 0.4505
R14972 DVSS.n3701 DVSS.n3667 0.4505
R14973 DVSS.n3703 DVSS.n3702 0.4505
R14974 DVSS.n3665 DVSS.n3664 0.4505
R14975 DVSS.n3708 DVSS.n3707 0.4505
R14976 DVSS.n3709 DVSS.n3663 0.4505
R14977 DVSS.n3711 DVSS.n3710 0.4505
R14978 DVSS.n3661 DVSS.n3660 0.4505
R14979 DVSS.n3716 DVSS.n3715 0.4505
R14980 DVSS.n3717 DVSS.n3659 0.4505
R14981 DVSS.n3719 DVSS.n3718 0.4505
R14982 DVSS.n3656 DVSS.n3654 0.4505
R14983 DVSS.n3743 DVSS.n3742 0.4505
R14984 DVSS.n3657 DVSS.n3655 0.4505
R14985 DVSS.n3738 DVSS.n3737 0.4505
R14986 DVSS.n3736 DVSS.n3723 0.4505
R14987 DVSS.n3735 DVSS.n3734 0.4505
R14988 DVSS.n3725 DVSS.n3724 0.4505
R14989 DVSS.n3730 DVSS.n3729 0.4505
R14990 DVSS.n3803 DVSS.n1646 0.4505
R14991 DVSS.n3827 DVSS.n3826 0.4505
R14992 DVSS.n3825 DVSS.n1633 0.4505
R14993 DVSS.n1638 DVSS.n1635 0.4505
R14994 DVSS.n3821 DVSS.n3820 0.4505
R14995 DVSS.n3819 DVSS.n1637 0.4505
R14996 DVSS.n3818 DVSS.n3817 0.4505
R14997 DVSS.n1640 DVSS.n1639 0.4505
R14998 DVSS.n3813 DVSS.n3812 0.4505
R14999 DVSS.n3811 DVSS.n1642 0.4505
R15000 DVSS.n3810 DVSS.n3809 0.4505
R15001 DVSS.n1644 DVSS.n1643 0.4505
R15002 DVSS.n3805 DVSS.n3804 0.4505
R15003 DVSS.n1596 DVSS.n1595 0.4505
R15004 DVSS.n1592 DVSS.n1590 0.4505
R15005 DVSS.n3893 DVSS.n3892 0.4505
R15006 DVSS.n1593 DVSS.n1591 0.4505
R15007 DVSS.n3888 DVSS.n3887 0.4505
R15008 DVSS.n3885 DVSS.n1600 0.4505
R15009 DVSS.n3884 DVSS.n3883 0.4505
R15010 DVSS.n1602 DVSS.n1601 0.4505
R15011 DVSS.n3879 DVSS.n3878 0.4505
R15012 DVSS.n3876 DVSS.n1604 0.4505
R15013 DVSS.n3874 DVSS.n3873 0.4505
R15014 DVSS.n1609 DVSS.n1606 0.4505
R15015 DVSS.n3869 DVSS.n3868 0.4505
R15016 DVSS.n3867 DVSS.n1608 0.4505
R15017 DVSS.n3866 DVSS.n3865 0.4505
R15018 DVSS.n1614 DVSS.n1611 0.4505
R15019 DVSS.n3861 DVSS.n3860 0.4505
R15020 DVSS.n3859 DVSS.n1613 0.4505
R15021 DVSS.n3855 DVSS.n3854 0.4505
R15022 DVSS.n1619 DVSS.n1616 0.4505
R15023 DVSS.n3850 DVSS.n3849 0.4505
R15024 DVSS.n3848 DVSS.n1618 0.4505
R15025 DVSS.n3847 DVSS.n3846 0.4505
R15026 DVSS.n1624 DVSS.n1621 0.4505
R15027 DVSS.n3842 DVSS.n3841 0.4505
R15028 DVSS.n3828 DVSS.n1623 0.4505
R15029 DVSS.n1099 DVSS.n1098 0.4505
R15030 DVSS.n5072 DVSS.n5071 0.4505
R15031 DVSS.n5070 DVSS.n1103 0.4505
R15032 DVSS.n5069 DVSS.n5068 0.4505
R15033 DVSS.n1105 DVSS.n1104 0.4505
R15034 DVSS.n5064 DVSS.n5063 0.4505
R15035 DVSS.n5062 DVSS.n1107 0.4505
R15036 DVSS.n5061 DVSS.n5060 0.4505
R15037 DVSS.n1109 DVSS.n1108 0.4505
R15038 DVSS.n5053 DVSS.n5052 0.4505
R15039 DVSS.n5051 DVSS.n1114 0.4505
R15040 DVSS.n5050 DVSS.n5049 0.4505
R15041 DVSS.n1116 DVSS.n1115 0.4505
R15042 DVSS.n5042 DVSS.n5041 0.4505
R15043 DVSS.n5040 DVSS.n1122 0.4505
R15044 DVSS.n5039 DVSS.n5038 0.4505
R15045 DVSS.n1124 DVSS.n1123 0.4505
R15046 DVSS.n5034 DVSS.n5033 0.4505
R15047 DVSS.n5032 DVSS.n1127 0.4505
R15048 DVSS.n5031 DVSS.n5030 0.4505
R15049 DVSS.n1129 DVSS.n1128 0.4505
R15050 DVSS.n5026 DVSS.n5025 0.4505
R15051 DVSS.n5024 DVSS.n1131 0.4505
R15052 DVSS.n5023 DVSS.n5022 0.4505
R15053 DVSS.n1133 DVSS.n1132 0.4505
R15054 DVSS.n5018 DVSS.n5017 0.4505
R15055 DVSS.n5016 DVSS.n1135 0.4505
R15056 DVSS.n5015 DVSS.n5014 0.4505
R15057 DVSS.n1137 DVSS.n1136 0.4505
R15058 DVSS.n5010 DVSS.n5009 0.4505
R15059 DVSS.n5008 DVSS.n1139 0.4505
R15060 DVSS.n5007 DVSS.n5006 0.4505
R15061 DVSS.n1141 DVSS.n1140 0.4505
R15062 DVSS.n5002 DVSS.n5001 0.4505
R15063 DVSS.n5000 DVSS.n1143 0.4505
R15064 DVSS.n4999 DVSS.n4998 0.4505
R15065 DVSS.n1145 DVSS.n1144 0.4505
R15066 DVSS.n4994 DVSS.n4993 0.4505
R15067 DVSS.n4992 DVSS.n1147 0.4505
R15068 DVSS.n4991 DVSS.n4990 0.4505
R15069 DVSS.n1149 DVSS.n1148 0.4505
R15070 DVSS.n4986 DVSS.n4985 0.4505
R15071 DVSS.n4984 DVSS.n1151 0.4505
R15072 DVSS.n4983 DVSS.n4982 0.4505
R15073 DVSS.n1153 DVSS.n1152 0.4505
R15074 DVSS.n2320 DVSS.n2319 0.4505
R15075 DVSS.n2322 DVSS.n2321 0.4505
R15076 DVSS.n2318 DVSS.n2317 0.4505
R15077 DVSS.n2327 DVSS.n2326 0.4505
R15078 DVSS.n2328 DVSS.n2316 0.4505
R15079 DVSS.n2330 DVSS.n2329 0.4505
R15080 DVSS.n2314 DVSS.n2313 0.4505
R15081 DVSS.n2335 DVSS.n2334 0.4505
R15082 DVSS.n2336 DVSS.n2312 0.4505
R15083 DVSS.n2338 DVSS.n2337 0.4505
R15084 DVSS.n2310 DVSS.n2309 0.4505
R15085 DVSS.n2343 DVSS.n2342 0.4505
R15086 DVSS.n2344 DVSS.n2308 0.4505
R15087 DVSS.n2346 DVSS.n2345 0.4505
R15088 DVSS.n2306 DVSS.n2305 0.4505
R15089 DVSS.n2351 DVSS.n2350 0.4505
R15090 DVSS.n2352 DVSS.n2304 0.4505
R15091 DVSS.n2354 DVSS.n2353 0.4505
R15092 DVSS.n2302 DVSS.n2301 0.4505
R15093 DVSS.n2359 DVSS.n2358 0.4505
R15094 DVSS.n2360 DVSS.n2300 0.4505
R15095 DVSS.n2362 DVSS.n2361 0.4505
R15096 DVSS.n2298 DVSS.n2297 0.4505
R15097 DVSS.n2367 DVSS.n2366 0.4505
R15098 DVSS.n2368 DVSS.n2296 0.4505
R15099 DVSS.n2370 DVSS.n2369 0.4505
R15100 DVSS.n2294 DVSS.n2293 0.4505
R15101 DVSS.n2375 DVSS.n2374 0.4505
R15102 DVSS.n2376 DVSS.n2292 0.4505
R15103 DVSS.n2378 DVSS.n2377 0.4505
R15104 DVSS.n2290 DVSS.n2289 0.4505
R15105 DVSS.n2383 DVSS.n2382 0.4505
R15106 DVSS.n2384 DVSS.n2288 0.4505
R15107 DVSS.n2387 DVSS.n2386 0.4505
R15108 DVSS.n2385 DVSS.n2286 0.4505
R15109 DVSS.n2391 DVSS.n2285 0.4505
R15110 DVSS.n2394 DVSS.n2393 0.4505
R15111 DVSS.n2395 DVSS.n2283 0.4505
R15112 DVSS.n2402 DVSS.n2401 0.4505
R15113 DVSS.n2400 DVSS.n2284 0.4505
R15114 DVSS.n5105 DVSS.n5104 0.4505
R15115 DVSS.n5103 DVSS.n1084 0.4505
R15116 DVSS.n5102 DVSS.n5101 0.4505
R15117 DVSS.n1086 DVSS.n1085 0.4505
R15118 DVSS.n5097 DVSS.n5096 0.4505
R15119 DVSS.n5095 DVSS.n1089 0.4505
R15120 DVSS.n5094 DVSS.n5093 0.4505
R15121 DVSS.n1091 DVSS.n1090 0.4505
R15122 DVSS.n5089 DVSS.n5088 0.4505
R15123 DVSS.n5087 DVSS.n1093 0.4505
R15124 DVSS.n5086 DVSS.n5085 0.4505
R15125 DVSS.n1095 DVSS.n1094 0.4505
R15126 DVSS.n5081 DVSS.n5080 0.4505
R15127 DVSS.n5079 DVSS.n1097 0.4505
R15128 DVSS.n5078 DVSS.n5077 0.4505
R15129 DVSS.n2398 DVSS.n2397 0.4505
R15130 DVSS.n2284 DVSS.n2282 0.4505
R15131 DVSS.n2403 DVSS.n2402 0.4505
R15132 DVSS.n2283 DVSS.n2279 0.4505
R15133 DVSS.n2393 DVSS.n2392 0.4505
R15134 DVSS.n2391 DVSS.n2390 0.4505
R15135 DVSS.n2389 DVSS.n2286 0.4505
R15136 DVSS.n2388 DVSS.n2387 0.4505
R15137 DVSS.n2288 DVSS.n2287 0.4505
R15138 DVSS.n2382 DVSS.n2381 0.4505
R15139 DVSS.n2380 DVSS.n2290 0.4505
R15140 DVSS.n2379 DVSS.n2378 0.4505
R15141 DVSS.n2292 DVSS.n2291 0.4505
R15142 DVSS.n2374 DVSS.n2373 0.4505
R15143 DVSS.n2372 DVSS.n2294 0.4505
R15144 DVSS.n2371 DVSS.n2370 0.4505
R15145 DVSS.n2296 DVSS.n2295 0.4505
R15146 DVSS.n2366 DVSS.n2365 0.4505
R15147 DVSS.n2364 DVSS.n2298 0.4505
R15148 DVSS.n2363 DVSS.n2362 0.4505
R15149 DVSS.n2300 DVSS.n2299 0.4505
R15150 DVSS.n2358 DVSS.n2357 0.4505
R15151 DVSS.n2356 DVSS.n2302 0.4505
R15152 DVSS.n2355 DVSS.n2354 0.4505
R15153 DVSS.n2304 DVSS.n2303 0.4505
R15154 DVSS.n2350 DVSS.n2349 0.4505
R15155 DVSS.n2348 DVSS.n2306 0.4505
R15156 DVSS.n2347 DVSS.n2346 0.4505
R15157 DVSS.n2308 DVSS.n2307 0.4505
R15158 DVSS.n2342 DVSS.n2341 0.4505
R15159 DVSS.n2340 DVSS.n2310 0.4505
R15160 DVSS.n2339 DVSS.n2338 0.4505
R15161 DVSS.n2312 DVSS.n2311 0.4505
R15162 DVSS.n2334 DVSS.n2333 0.4505
R15163 DVSS.n2332 DVSS.n2314 0.4505
R15164 DVSS.n2331 DVSS.n2330 0.4505
R15165 DVSS.n2316 DVSS.n2315 0.4505
R15166 DVSS.n2326 DVSS.n2325 0.4505
R15167 DVSS.n2324 DVSS.n2318 0.4505
R15168 DVSS.n2323 DVSS.n2322 0.4505
R15169 DVSS.n2319 DVSS.n1154 0.4505
R15170 DVSS.n4980 DVSS.n1153 0.4505
R15171 DVSS.n4982 DVSS.n4981 0.4505
R15172 DVSS.n1151 DVSS.n1150 0.4505
R15173 DVSS.n4987 DVSS.n4986 0.4505
R15174 DVSS.n4988 DVSS.n1149 0.4505
R15175 DVSS.n4990 DVSS.n4989 0.4505
R15176 DVSS.n1147 DVSS.n1146 0.4505
R15177 DVSS.n4995 DVSS.n4994 0.4505
R15178 DVSS.n4996 DVSS.n1145 0.4505
R15179 DVSS.n4998 DVSS.n4997 0.4505
R15180 DVSS.n1143 DVSS.n1142 0.4505
R15181 DVSS.n5003 DVSS.n5002 0.4505
R15182 DVSS.n5004 DVSS.n1141 0.4505
R15183 DVSS.n5006 DVSS.n5005 0.4505
R15184 DVSS.n1139 DVSS.n1138 0.4505
R15185 DVSS.n5011 DVSS.n5010 0.4505
R15186 DVSS.n5012 DVSS.n1137 0.4505
R15187 DVSS.n5014 DVSS.n5013 0.4505
R15188 DVSS.n1135 DVSS.n1134 0.4505
R15189 DVSS.n5019 DVSS.n5018 0.4505
R15190 DVSS.n5020 DVSS.n1133 0.4505
R15191 DVSS.n5022 DVSS.n5021 0.4505
R15192 DVSS.n1131 DVSS.n1130 0.4505
R15193 DVSS.n5027 DVSS.n5026 0.4505
R15194 DVSS.n5028 DVSS.n1129 0.4505
R15195 DVSS.n5030 DVSS.n5029 0.4505
R15196 DVSS.n1127 DVSS.n1126 0.4505
R15197 DVSS.n5035 DVSS.n5034 0.4505
R15198 DVSS.n5036 DVSS.n1124 0.4505
R15199 DVSS.n5038 DVSS.n5037 0.4505
R15200 DVSS.n1125 DVSS.n1122 0.4505
R15201 DVSS.n5043 DVSS.n5042 0.4505
R15202 DVSS.n1119 DVSS.n1116 0.4505
R15203 DVSS.n5049 DVSS.n5048 0.4505
R15204 DVSS.n1117 DVSS.n1114 0.4505
R15205 DVSS.n5054 DVSS.n5053 0.4505
R15206 DVSS.n1111 DVSS.n1109 0.4505
R15207 DVSS.n5060 DVSS.n5059 0.4505
R15208 DVSS.n1107 DVSS.n1106 0.4505
R15209 DVSS.n5065 DVSS.n5064 0.4505
R15210 DVSS.n5066 DVSS.n1105 0.4505
R15211 DVSS.n5068 DVSS.n5067 0.4505
R15212 DVSS.n1103 DVSS.n1102 0.4505
R15213 DVSS.n5073 DVSS.n5072 0.4505
R15214 DVSS.n5074 DVSS.n1099 0.4505
R15215 DVSS.n5107 DVSS.n5106 0.4505
R15216 DVSS.n5105 DVSS.n1083 0.4505
R15217 DVSS.n1087 DVSS.n1084 0.4505
R15218 DVSS.n5101 DVSS.n5100 0.4505
R15219 DVSS.n5099 DVSS.n1086 0.4505
R15220 DVSS.n5098 DVSS.n5097 0.4505
R15221 DVSS.n1089 DVSS.n1088 0.4505
R15222 DVSS.n5093 DVSS.n5092 0.4505
R15223 DVSS.n5091 DVSS.n1091 0.4505
R15224 DVSS.n5090 DVSS.n5089 0.4505
R15225 DVSS.n1093 DVSS.n1092 0.4505
R15226 DVSS.n5085 DVSS.n5084 0.4505
R15227 DVSS.n5083 DVSS.n1095 0.4505
R15228 DVSS.n5082 DVSS.n5081 0.4505
R15229 DVSS.n1097 DVSS.n1096 0.4505
R15230 DVSS.n5077 DVSS.n5076 0.4505
R15231 DVSS.n2266 DVSS.n2265 0.4505
R15232 DVSS.n2651 DVSS.n2650 0.4505
R15233 DVSS.n2649 DVSS.n2268 0.4505
R15234 DVSS.n2632 DVSS.n2269 0.4505
R15235 DVSS.n2636 DVSS.n2635 0.4505
R15236 DVSS.n2494 DVSS.n2493 0.4505
R15237 DVSS.n2498 DVSS.n2497 0.4505
R15238 DVSS.n2499 DVSS.n2492 0.4505
R15239 DVSS.n2501 DVSS.n2500 0.4505
R15240 DVSS.n2490 DVSS.n2489 0.4505
R15241 DVSS.n2506 DVSS.n2505 0.4505
R15242 DVSS.n2507 DVSS.n2488 0.4505
R15243 DVSS.n2509 DVSS.n2508 0.4505
R15244 DVSS.n2486 DVSS.n2485 0.4505
R15245 DVSS.n2514 DVSS.n2513 0.4505
R15246 DVSS.n2515 DVSS.n2484 0.4505
R15247 DVSS.n2517 DVSS.n2516 0.4505
R15248 DVSS.n2482 DVSS.n2481 0.4505
R15249 DVSS.n2522 DVSS.n2521 0.4505
R15250 DVSS.n2523 DVSS.n2480 0.4505
R15251 DVSS.n2525 DVSS.n2524 0.4505
R15252 DVSS.n2478 DVSS.n2477 0.4505
R15253 DVSS.n2530 DVSS.n2529 0.4505
R15254 DVSS.n2531 DVSS.n2476 0.4505
R15255 DVSS.n2533 DVSS.n2532 0.4505
R15256 DVSS.n2474 DVSS.n2473 0.4505
R15257 DVSS.n2538 DVSS.n2537 0.4505
R15258 DVSS.n2539 DVSS.n2472 0.4505
R15259 DVSS.n2541 DVSS.n2540 0.4505
R15260 DVSS.n2470 DVSS.n2469 0.4505
R15261 DVSS.n2546 DVSS.n2545 0.4505
R15262 DVSS.n2547 DVSS.n2468 0.4505
R15263 DVSS.n2549 DVSS.n2548 0.4505
R15264 DVSS.n2466 DVSS.n2465 0.4505
R15265 DVSS.n2554 DVSS.n2553 0.4505
R15266 DVSS.n2555 DVSS.n2464 0.4505
R15267 DVSS.n2557 DVSS.n2556 0.4505
R15268 DVSS.n2462 DVSS.n2461 0.4505
R15269 DVSS.n2562 DVSS.n2561 0.4505
R15270 DVSS.n2563 DVSS.n2460 0.4505
R15271 DVSS.n2565 DVSS.n2564 0.4505
R15272 DVSS.n2458 DVSS.n2457 0.4505
R15273 DVSS.n2570 DVSS.n2569 0.4505
R15274 DVSS.n2571 DVSS.n2456 0.4505
R15275 DVSS.n2573 DVSS.n2572 0.4505
R15276 DVSS.n2454 DVSS.n2453 0.4505
R15277 DVSS.n2578 DVSS.n2577 0.4505
R15278 DVSS.n2579 DVSS.n2452 0.4505
R15279 DVSS.n2581 DVSS.n2580 0.4505
R15280 DVSS.n2450 DVSS.n2449 0.4505
R15281 DVSS.n2586 DVSS.n2585 0.4505
R15282 DVSS.n2587 DVSS.n2448 0.4505
R15283 DVSS.n2589 DVSS.n2588 0.4505
R15284 DVSS.n2446 DVSS.n2445 0.4505
R15285 DVSS.n2594 DVSS.n2593 0.4505
R15286 DVSS.n2595 DVSS.n2444 0.4505
R15287 DVSS.n2597 DVSS.n2596 0.4505
R15288 DVSS.n2442 DVSS.n2441 0.4505
R15289 DVSS.n2602 DVSS.n2601 0.4505
R15290 DVSS.n2603 DVSS.n2440 0.4505
R15291 DVSS.n2605 DVSS.n2604 0.4505
R15292 DVSS.n2438 DVSS.n2437 0.4505
R15293 DVSS.n2610 DVSS.n2609 0.4505
R15294 DVSS.n2611 DVSS.n2436 0.4505
R15295 DVSS.n2613 DVSS.n2612 0.4505
R15296 DVSS.n2434 DVSS.n2433 0.4505
R15297 DVSS.n2618 DVSS.n2617 0.4505
R15298 DVSS.n2619 DVSS.n2432 0.4505
R15299 DVSS.n2621 DVSS.n2620 0.4505
R15300 DVSS.n2430 DVSS.n2429 0.4505
R15301 DVSS.n2626 DVSS.n2625 0.4505
R15302 DVSS.n2627 DVSS.n2428 0.4505
R15303 DVSS.n2629 DVSS.n2628 0.4505
R15304 DVSS.n2426 DVSS.n2421 0.4505
R15305 DVSS.n1537 DVSS.n1536 0.4505
R15306 DVSS.n1538 DVSS.n1533 0.4505
R15307 DVSS.n1540 DVSS.n1539 0.4505
R15308 DVSS.n1531 DVSS.n1530 0.4505
R15309 DVSS.n1545 DVSS.n1544 0.4505
R15310 DVSS.n1546 DVSS.n1529 0.4505
R15311 DVSS.n1548 DVSS.n1547 0.4505
R15312 DVSS.n1527 DVSS.n1526 0.4505
R15313 DVSS.n1553 DVSS.n1552 0.4505
R15314 DVSS.n1554 DVSS.n1525 0.4505
R15315 DVSS.n1556 DVSS.n1555 0.4505
R15316 DVSS.n1522 DVSS.n1520 0.4505
R15317 DVSS.n3936 DVSS.n3935 0.4505
R15318 DVSS.n1523 DVSS.n1521 0.4505
R15319 DVSS.n3931 DVSS.n3930 0.4505
R15320 DVSS.n3929 DVSS.n1560 0.4505
R15321 DVSS.n3928 DVSS.n3927 0.4505
R15322 DVSS.n1562 DVSS.n1561 0.4505
R15323 DVSS.n3923 DVSS.n3922 0.4505
R15324 DVSS.n3921 DVSS.n1564 0.4505
R15325 DVSS.n3920 DVSS.n3919 0.4505
R15326 DVSS.n1566 DVSS.n1565 0.4505
R15327 DVSS.n3915 DVSS.n3914 0.4505
R15328 DVSS.n3913 DVSS.n1568 0.4505
R15329 DVSS.n3912 DVSS.n3911 0.4505
R15330 DVSS.n1570 DVSS.n1569 0.4505
R15331 DVSS.n3907 DVSS.n3906 0.4505
R15332 DVSS.n1573 DVSS.n1572 0.4505
R15333 DVSS.n4452 DVSS 0.449176
R15334 DVSS.n4961 DVSS 0.449176
R15335 DVSS.n4961 DVSS 0.449176
R15336 DVSS.n3563 VSS 0.444617
R15337 DVSS.n2251 VSS 0.444617
R15338 DVSS.n3560 VSS 0.444542
R15339 DVSS.n2250 VSS 0.444542
R15340 DVSS.n3617 DVSS.n3616 0.441235
R15341 DVSS.n1193 DVSS.n957 0.439524
R15342 DVSS.n5358 DVSS.n5357 0.439458
R15343 DVSS.n2796 DVSS.n2795 0.429011
R15344 DVSS.n2797 DVSS.n2796 0.429011
R15345 DVSS.n4410 DVSS.n4376 0.41962
R15346 DVSS.n1475 DVSS.n1291 0.41962
R15347 DVSS.n1512 DVSS.n1511 0.4165
R15348 DVSS.n3952 DVSS.n3951 0.4165
R15349 DVSS.n3561 VSS 0.415539
R15350 DVSS.n3562 VSS 0.415539
R15351 DVSS.n3956 DVSS.n3955 0.412794
R15352 DVSS.n2239 DVSS.t104 0.41
R15353 DVSS.n2239 DVSS.t106 0.41
R15354 DVSS.n4189 DVSS.n4188 0.407769
R15355 DVSS.n3766 DVSS 0.402853
R15356 DVSS.n3791 DVSS 0.402853
R15357 DVSS.n3901 DVSS 0.402853
R15358 DVSS DVSS.n3897 0.402853
R15359 DVSS.n2154 DVSS.n2152 0.388068
R15360 DVSS.n1915 DVSS.n1813 0.387662
R15361 DVSS.n4452 DVSS 0.384324
R15362 DVSS.n4190 DVSS.n4189 0.38247
R15363 DVSS.n3560 DVSS.n1519 0.375755
R15364 DVSS.n2156 DVSS.n2155 0.3755
R15365 DVSS.n1917 DVSS.n1916 0.3755
R15366 DVSS.n1444 DVSS.n1443 0.3755
R15367 DVSS.n1659 DVSS.n1658 0.368789
R15368 DVSS.n3768 DVSS.n3767 0.368789
R15369 DVSS.n3766 DVSS.n1693 0.368789
R15370 DVSS.n3765 DVSS.n3764 0.368789
R15371 DVSS.n1673 DVSS.n1672 0.368789
R15372 DVSS.n3792 DVSS.n3791 0.368789
R15373 DVSS.n3857 DVSS.n1574 0.368789
R15374 DVSS.n3901 DVSS.n1577 0.368789
R15375 DVSS.n3900 DVSS.n1579 0.368789
R15376 DVSS.n3898 DVSS.n1582 0.368789
R15377 DVSS.n3897 DVSS.n1585 0.368789
R15378 DVSS.n3896 DVSS.n3895 0.368789
R15379 DVSS.n3628 DVSS.n1720 0.367935
R15380 DVSS.n3628 DVSS.n1710 0.367935
R15381 DVSS.n3625 DVSS.n1726 0.367935
R15382 DVSS.n1726 DVSS.n1711 0.367935
R15383 DVSS.n3598 DVSS.n1727 0.367935
R15384 DVSS.n1727 DVSS.n1712 0.367935
R15385 DVSS.n3599 DVSS.n1728 0.367935
R15386 DVSS.n1728 DVSS.n1713 0.367935
R15387 DVSS.n3600 DVSS.n1729 0.367935
R15388 DVSS.n1729 DVSS.n1714 0.367935
R15389 DVSS.n3601 DVSS.n1715 0.367935
R15390 DVSS.n3633 DVSS.n3593 0.367935
R15391 DVSS.n3594 DVSS.n1714 0.367935
R15392 DVSS.n3595 DVSS.n1713 0.367935
R15393 DVSS.n3596 DVSS.n1712 0.367935
R15394 DVSS.n3597 DVSS.n1711 0.367935
R15395 DVSS.n3644 DVSS.n1710 0.367935
R15396 DVSS.n3601 DVSS.n3594 0.367935
R15397 DVSS.n3600 DVSS.n3595 0.367935
R15398 DVSS.n3599 DVSS.n3596 0.367935
R15399 DVSS.n3598 DVSS.n3597 0.367935
R15400 DVSS.n3644 DVSS.n3625 0.367935
R15401 DVSS.n3646 DVSS.n1720 0.367935
R15402 DVSS.n3593 DVSS.n1715 0.367935
R15403 DVSS.n1280 DVSS 0.366421
R15404 DVSS.n4436 DVSS 0.366421
R15405 DVSS.n1462 DVSS 0.366421
R15406 DVSS.n4398 DVSS 0.366421
R15407 DVSS.n3987 DVSS 0.358788
R15408 DVSS.n4184 DVSS.n1369 0.346654
R15409 DVSS.n4184 DVSS.n4183 0.346654
R15410 DVSS.n1282 DVSS 0.346309
R15411 DVSS.n1284 DVSS 0.346309
R15412 DVSS.n1310 DVSS 0.346309
R15413 DVSS.n4438 DVSS 0.346309
R15414 DVSS.n1464 DVSS 0.346309
R15415 DVSS.n1460 DVSS 0.346309
R15416 DVSS.n4396 DVSS 0.346309
R15417 DVSS.n4400 DVSS 0.346309
R15418 DVSS.n1277 DVSS 0.346114
R15419 DVSS.n4441 DVSS 0.346114
R15420 DVSS.n1307 DVSS 0.346114
R15421 DVSS.n4307 DVSS.n1164 0.342906
R15422 DVSS.n3653 DVSS.n1706 0.338834
R15423 DVSS.n3565 DVSS.n3564 0.335984
R15424 DVSS.n4899 DVSS.n4776 0.328381
R15425 DVSS.n4886 DVSS.n4885 0.328381
R15426 DVSS.n4755 DVSS.n4754 0.328381
R15427 DVSS.n4769 DVSS.n1219 0.328381
R15428 DVSS.n4717 DVSS.n1251 0.328381
R15429 DVSS.n4735 DVSS.n4734 0.328381
R15430 DVSS.n4619 DVSS.n1271 0.328381
R15431 DVSS.n4695 DVSS.n4694 0.328381
R15432 DVSS.n4651 DVSS.n4583 0.328381
R15433 DVSS.n4638 DVSS.n4637 0.328381
R15434 DVSS.n4562 DVSS.n4561 0.328381
R15435 DVSS.n4576 DVSS.n4493 0.328381
R15436 DVSS.n1709 DVSS.n1708 0.3255
R15437 DVSS.n1708 DVSS.n1700 0.3255
R15438 DVSS.n3747 DVSS.n3746 0.316244
R15439 DVSS.n1921 DVSS.n1920 0.311888
R15440 DVSS.n2160 DVSS.n2159 0.311888
R15441 DVSS DVSS.n1733 0.309579
R15442 DVSS.n3564 DVSS.n3560 0.307559
R15443 DVSS.n4480 DVSS.n4479 0.297643
R15444 DVSS.n1468 DVSS.n1300 0.297643
R15445 DVSS.n4430 DVSS.n4429 0.297643
R15446 DVSS.n4404 DVSS.n4403 0.297643
R15447 DVSS.n804 DVSS.n803 0.28175
R15448 DVSS.n365 DVSS.n229 0.28175
R15449 DVSS.n3620 DVSS 0.273784
R15450 DVSS.n1288 DVSS.t168 0.2735
R15451 DVSS.n1288 DVSS.t203 0.2735
R15452 DVSS.n1293 DVSS.t67 0.2735
R15453 DVSS.n1293 DVSS.t174 0.2735
R15454 DVSS.n4186 DVSS.t65 0.2735
R15455 DVSS.n1276 DVSS.t162 0.2735
R15456 DVSS.n1281 DVSS.t131 0.2735
R15457 DVSS.n1281 DVSS.t160 0.2735
R15458 DVSS.n1283 DVSS.t164 0.2735
R15459 DVSS.n1283 DVSS.t102 0.2735
R15460 DVSS.n4379 DVSS.t191 0.2735
R15461 DVSS.n4379 DVSS.t170 0.2735
R15462 DVSS.n1313 DVSS.t172 0.2735
R15463 DVSS.n1313 DVSS.t153 0.2735
R15464 DVSS.n4426 DVSS.t151 0.2735
R15465 DVSS.n1309 DVSS.t110 0.2735
R15466 DVSS.n1309 DVSS.t84 0.2735
R15467 DVSS.n4437 DVSS.t112 0.2735
R15468 DVSS.n4437 DVSS.t114 0.2735
R15469 DVSS.n4440 DVSS.t205 0.2735
R15470 DVSS.n1306 DVSS.t71 0.2735
R15471 DVSS.n1463 DVSS.t73 0.2735
R15472 DVSS.n1463 DVSS.t75 0.2735
R15473 DVSS.n1459 DVSS.t86 0.2735
R15474 DVSS.n1459 DVSS.t77 0.2735
R15475 DVSS.n1471 DVSS.t69 0.2735
R15476 DVSS.n4392 DVSS.t189 0.2735
R15477 DVSS.n4395 DVSS.t201 0.2735
R15478 DVSS.n4395 DVSS.t121 0.2735
R15479 DVSS.n4399 DVSS.t193 0.2735
R15480 DVSS.n4399 DVSS.t140 0.2735
R15481 DVSS.n4337 DVSS.t149 0.2735
R15482 DVSS.n3958 DVSS.n1503 0.273147
R15483 DVSS.n3949 DVSS.n3946 0.273147
R15484 DVSS.n4462 DVSS.n1291 0.271321
R15485 DVSS.n4410 DVSS.n4409 0.271321
R15486 DVSS.n3585 DVSS.n3584 0.268132
R15487 DVSS.n4943 DVSS.n4942 0.266421
R15488 DVSS.n4443 DVSS.n1308 0.265206
R15489 DVSS.n4443 DVSS.n4442 0.265206
R15490 DVSS.n105 DVSS.n61 0.265206
R15491 DVSS.n260 DVSS.n252 0.265206
R15492 DVSS.n4203 DVSS.n1291 0.264797
R15493 DVSS.n4411 DVSS.n4410 0.264797
R15494 DVSS.n4486 DVSS.n4485 0.2605
R15495 DVSS.n4445 DVSS.n4444 0.2605
R15496 DVSS.n4944 DVSS.n4943 0.2605
R15497 VSS DVSS.n1449 0.258658
R15498 DVSS.n3981 DVSS.n1440 0.254359
R15499 DVSS.n1484 DVSS.n1483 0.249324
R15500 DVSS.n4975 DVSS.n4970 0.249324
R15501 DVSS.n4947 DVSS.n1168 0.249324
R15502 DVSS.n4427 DVSS.n4424 0.243385
R15503 DVSS.n1472 DVSS.n1469 0.243385
R15504 DVSS.n4188 DVSS.n4185 0.243385
R15505 DVSS.n4393 DVSS.n4390 0.243385
R15506 DVSS.n4339 DVSS.n4336 0.243385
R15507 DVSS.n3584 DVSS.n3583 0.242079
R15508 DVSS.n3564 DVSS.n3563 0.238735
R15509 DVSS.n5809 DVSS.n5808 0.232304
R15510 DVSS.n1918 DVSS.n1917 0.231484
R15511 DVSS.n2157 DVSS.n2156 0.231484
R15512 DVSS.n4850 DVSS.n4849 0.231338
R15513 DVSS.n1535 DVSS.n1532 0.231338
R15514 DVSS.n2653 DVSS.n2652 0.231338
R15515 DVSS.n5104 DVSS.n1082 0.231338
R15516 DVSS.n2400 DVSS.n2399 0.231338
R15517 DVSS.n5562 DVSS.n5561 0.229958
R15518 DVSS.n5814 DVSS.n5813 0.229958
R15519 DVSS.n1917 DVSS.n1880 0.229569
R15520 VSS DVSS.n1155 0.229471
R15521 VSS DVSS.n1155 0.229471
R15522 DVSS.n2156 DVSS.n1811 0.228851
R15523 DVSS.n1449 DVSS.n1448 0.224316
R15524 DVSS.n3608 DVSS 0.223543
R15525 DVSS.n4937 DVSS.n4936 0.219756
R15526 DVSS.n55 DVSS.n48 0.214786
R15527 DVSS.n426 DVSS.n425 0.214786
R15528 DVSS.n4939 DVSS.n1176 0.214786
R15529 DVSS.n4334 DVSS.n1175 0.214786
R15530 DVSS.n4342 DVSS.n4335 0.214786
R15531 DVSS.n4343 DVSS.n4333 0.214786
R15532 DVSS.n4344 DVSS.n4332 0.214786
R15533 DVSS.n4331 DVSS.n4329 0.214786
R15534 DVSS.n4348 DVSS.n4328 0.214786
R15535 DVSS.n4349 DVSS.n4327 0.214786
R15536 DVSS.n4350 DVSS.n4326 0.214786
R15537 DVSS.n4325 DVSS.n4323 0.214786
R15538 DVSS.n4354 DVSS.n4322 0.214786
R15539 DVSS.n4355 DVSS.n4321 0.214786
R15540 DVSS.n4356 DVSS.n4320 0.214786
R15541 DVSS.n4319 DVSS.n4317 0.214786
R15542 DVSS.n4360 DVSS.n4316 0.214786
R15543 DVSS.n4361 DVSS.n4315 0.214786
R15544 DVSS.n4362 DVSS.n4314 0.214786
R15545 DVSS.n4313 DVSS.n4311 0.214786
R15546 DVSS.n4366 DVSS.n4310 0.214786
R15547 DVSS.n4367 DVSS.n4309 0.214786
R15548 DVSS.n4308 DVSS.n4306 0.214786
R15549 DVSS.n4371 DVSS.n4305 0.214786
R15550 DVSS.n4372 DVSS.n4304 0.214786
R15551 DVSS.n4373 DVSS.n4303 0.214786
R15552 DVSS.n4302 DVSS.n4300 0.214786
R15553 DVSS.n4413 DVSS.n4299 0.214786
R15554 DVSS.n4414 DVSS.n4298 0.214786
R15555 DVSS.n4415 DVSS.n4297 0.214786
R15556 DVSS.n4296 DVSS.n4294 0.214786
R15557 DVSS.n4419 DVSS.n4293 0.214786
R15558 DVSS.n4420 DVSS.n4292 0.214786
R15559 DVSS.n4193 DVSS.n4192 0.214786
R15560 DVSS.n1365 DVSS.n1364 0.214786
R15561 DVSS.n4198 DVSS.n4197 0.214786
R15562 DVSS.n4199 DVSS.n1363 0.214786
R15563 DVSS.n4201 DVSS.n4200 0.214786
R15564 DVSS.n1361 DVSS.n1360 0.214786
R15565 DVSS.n4207 DVSS.n4206 0.214786
R15566 DVSS.n4208 DVSS.n1359 0.214786
R15567 DVSS.n4210 DVSS.n4209 0.214786
R15568 DVSS.n1357 DVSS.n1356 0.214786
R15569 DVSS.n4216 DVSS.n4215 0.214786
R15570 DVSS.n4217 DVSS.n1355 0.214786
R15571 DVSS.n4219 DVSS.n4218 0.214786
R15572 DVSS.n1353 DVSS.n1352 0.214786
R15573 DVSS.n4224 DVSS.n4223 0.214786
R15574 DVSS.n4225 DVSS.n1351 0.214786
R15575 DVSS.n4227 DVSS.n4226 0.214786
R15576 DVSS.n1349 DVSS.n1348 0.214786
R15577 DVSS.n4232 DVSS.n4231 0.214786
R15578 DVSS.n4233 DVSS.n1347 0.214786
R15579 DVSS.n4235 DVSS.n4234 0.214786
R15580 DVSS.n1345 DVSS.n1344 0.214786
R15581 DVSS.n4241 DVSS.n4240 0.214786
R15582 DVSS.n4242 DVSS.n1343 0.214786
R15583 DVSS.n4244 DVSS.n4243 0.214786
R15584 DVSS.n1341 DVSS.n1340 0.214786
R15585 DVSS.n4249 DVSS.n4248 0.214786
R15586 DVSS.n4250 DVSS.n1339 0.214786
R15587 DVSS.n4252 DVSS.n4251 0.214786
R15588 DVSS.n1337 DVSS.n1336 0.214786
R15589 DVSS.n4257 DVSS.n4256 0.214786
R15590 DVSS.n4258 DVSS.n1335 0.214786
R15591 DVSS.n4260 DVSS.n4259 0.214786
R15592 DVSS.n1333 DVSS.n1332 0.214786
R15593 DVSS.n4265 DVSS.n4264 0.214786
R15594 DVSS.n4266 DVSS.n1331 0.214786
R15595 DVSS.n4268 DVSS.n4267 0.214786
R15596 DVSS.n1329 DVSS.n1328 0.214786
R15597 DVSS.n4273 DVSS.n4272 0.214786
R15598 DVSS.n4274 DVSS.n1327 0.214786
R15599 DVSS.n4276 DVSS.n4275 0.214786
R15600 DVSS.n1325 DVSS.n1324 0.214786
R15601 DVSS.n4281 DVSS.n4280 0.214786
R15602 DVSS.n4282 DVSS.n1323 0.214786
R15603 DVSS.n4284 DVSS.n4283 0.214786
R15604 DVSS.n1321 DVSS.n1320 0.214786
R15605 DVSS.n4289 DVSS.n4288 0.214786
R15606 DVSS.n4290 DVSS.n1319 0.214786
R15607 DVSS.n4421 DVSS.n4291 0.214786
R15608 DVSS.n4202 DVSS.n4201 0.214786
R15609 DVSS.n4938 DVSS.n1174 0.214786
R15610 DVSS.n4940 DVSS.n4939 0.214786
R15611 DVSS.n1175 DVSS.n1173 0.214786
R15612 DVSS.n4342 DVSS.n4341 0.214786
R15613 DVSS.n4343 DVSS.n4330 0.214786
R15614 DVSS.n4345 DVSS.n4344 0.214786
R15615 DVSS.n4346 DVSS.n4329 0.214786
R15616 DVSS.n4348 DVSS.n4347 0.214786
R15617 DVSS.n4349 DVSS.n4324 0.214786
R15618 DVSS.n4351 DVSS.n4350 0.214786
R15619 DVSS.n4352 DVSS.n4323 0.214786
R15620 DVSS.n4354 DVSS.n4353 0.214786
R15621 DVSS.n4355 DVSS.n4318 0.214786
R15622 DVSS.n4357 DVSS.n4356 0.214786
R15623 DVSS.n4358 DVSS.n4317 0.214786
R15624 DVSS.n4360 DVSS.n4359 0.214786
R15625 DVSS.n4361 DVSS.n4312 0.214786
R15626 DVSS.n4363 DVSS.n4362 0.214786
R15627 DVSS.n4364 DVSS.n4311 0.214786
R15628 DVSS.n4366 DVSS.n4365 0.214786
R15629 DVSS.n4368 DVSS.n4367 0.214786
R15630 DVSS.n4369 DVSS.n4306 0.214786
R15631 DVSS.n4371 DVSS.n4370 0.214786
R15632 DVSS.n4372 DVSS.n4301 0.214786
R15633 DVSS.n4374 DVSS.n4373 0.214786
R15634 DVSS.n4375 DVSS.n4300 0.214786
R15635 DVSS.n4420 DVSS.n1318 0.214786
R15636 DVSS.n4419 DVSS.n4418 0.214786
R15637 DVSS.n4417 DVSS.n4294 0.214786
R15638 DVSS.n4416 DVSS.n4415 0.214786
R15639 DVSS.n4414 DVSS.n4295 0.214786
R15640 DVSS.n4413 DVSS.n4412 0.214786
R15641 DVSS.n1367 DVSS.n1366 0.214786
R15642 DVSS.n4194 DVSS.n4193 0.214786
R15643 DVSS.n4195 DVSS.n1365 0.214786
R15644 DVSS.n4197 DVSS.n4196 0.214786
R15645 DVSS.n1363 DVSS.n1362 0.214786
R15646 DVSS.n4204 DVSS.n1361 0.214786
R15647 DVSS.n4206 DVSS.n4205 0.214786
R15648 DVSS.n1359 DVSS.n1358 0.214786
R15649 DVSS.n4211 DVSS.n4210 0.214786
R15650 DVSS.n4212 DVSS.n1357 0.214786
R15651 DVSS.n4215 DVSS.n4214 0.214786
R15652 DVSS.n4213 DVSS.n1355 0.214786
R15653 DVSS.n4220 DVSS.n4219 0.214786
R15654 DVSS.n4221 DVSS.n1353 0.214786
R15655 DVSS.n4223 DVSS.n4222 0.214786
R15656 DVSS.n1351 DVSS.n1350 0.214786
R15657 DVSS.n4228 DVSS.n4227 0.214786
R15658 DVSS.n4229 DVSS.n1349 0.214786
R15659 DVSS.n4231 DVSS.n4230 0.214786
R15660 DVSS.n1347 DVSS.n1346 0.214786
R15661 DVSS.n4236 DVSS.n4235 0.214786
R15662 DVSS.n4237 DVSS.n1345 0.214786
R15663 DVSS.n4240 DVSS.n4239 0.214786
R15664 DVSS.n1343 DVSS.n1342 0.214786
R15665 DVSS.n4245 DVSS.n4244 0.214786
R15666 DVSS.n4246 DVSS.n1341 0.214786
R15667 DVSS.n4248 DVSS.n4247 0.214786
R15668 DVSS.n1339 DVSS.n1338 0.214786
R15669 DVSS.n4253 DVSS.n4252 0.214786
R15670 DVSS.n4254 DVSS.n1337 0.214786
R15671 DVSS.n4256 DVSS.n4255 0.214786
R15672 DVSS.n1335 DVSS.n1334 0.214786
R15673 DVSS.n4261 DVSS.n4260 0.214786
R15674 DVSS.n4262 DVSS.n1333 0.214786
R15675 DVSS.n4264 DVSS.n4263 0.214786
R15676 DVSS.n1331 DVSS.n1330 0.214786
R15677 DVSS.n4269 DVSS.n4268 0.214786
R15678 DVSS.n4270 DVSS.n1329 0.214786
R15679 DVSS.n4272 DVSS.n4271 0.214786
R15680 DVSS.n1327 DVSS.n1326 0.214786
R15681 DVSS.n4277 DVSS.n4276 0.214786
R15682 DVSS.n4278 DVSS.n1325 0.214786
R15683 DVSS.n4280 DVSS.n4279 0.214786
R15684 DVSS.n1323 DVSS.n1322 0.214786
R15685 DVSS.n4285 DVSS.n4284 0.214786
R15686 DVSS.n4286 DVSS.n1321 0.214786
R15687 DVSS.n4288 DVSS.n4287 0.214786
R15688 DVSS.n1319 DVSS.n1317 0.214786
R15689 DVSS.n4422 DVSS.n4421 0.214786
R15690 DVSS.n497 DVSS.n209 0.214786
R15691 DVSS.n828 DVSS.n826 0.214786
R15692 DVSS.n827 DVSS.n825 0.214786
R15693 DVSS.n5565 DVSS.n824 0.214786
R15694 DVSS.n5566 DVSS.n823 0.214786
R15695 DVSS.n5567 DVSS.n822 0.214786
R15696 DVSS.n821 DVSS.n819 0.214786
R15697 DVSS.n5571 DVSS.n818 0.214786
R15698 DVSS.n5572 DVSS.n817 0.214786
R15699 DVSS.n5573 DVSS.n816 0.214786
R15700 DVSS.n815 DVSS.n813 0.214786
R15701 DVSS.n5577 DVSS.n812 0.214786
R15702 DVSS.n5578 DVSS.n811 0.214786
R15703 DVSS.n5579 DVSS.n810 0.214786
R15704 DVSS.n809 DVSS.n807 0.214786
R15705 DVSS.n5583 DVSS.n806 0.214786
R15706 DVSS.n5585 DVSS.n805 0.214786
R15707 DVSS.n753 DVSS.n752 0.214786
R15708 DVSS.n5589 DVSS.n751 0.214786
R15709 DVSS.n5590 DVSS.n750 0.214786
R15710 DVSS.n5591 DVSS.n749 0.214786
R15711 DVSS.n748 DVSS.n746 0.214786
R15712 DVSS.n5595 DVSS.n745 0.214786
R15713 DVSS.n5596 DVSS.n744 0.214786
R15714 DVSS.n5597 DVSS.n743 0.214786
R15715 DVSS.n742 DVSS.n740 0.214786
R15716 DVSS.n5601 DVSS.n739 0.214786
R15717 DVSS.n5602 DVSS.n738 0.214786
R15718 DVSS.n5603 DVSS.n737 0.214786
R15719 DVSS.n736 DVSS.n734 0.214786
R15720 DVSS.n5607 DVSS.n733 0.214786
R15721 DVSS.n5608 DVSS.n732 0.214786
R15722 DVSS.n5609 DVSS.n731 0.214786
R15723 DVSS.n147 DVSS.n145 0.214786
R15724 DVSS.n5614 DVSS.n5613 0.214786
R15725 DVSS.n146 DVSS.n144 0.214786
R15726 DVSS.n727 DVSS.n726 0.214786
R15727 DVSS.n725 DVSS.n149 0.214786
R15728 DVSS.n724 DVSS.n723 0.214786
R15729 DVSS.n151 DVSS.n150 0.214786
R15730 DVSS.n718 DVSS.n717 0.214786
R15731 DVSS.n154 DVSS.n153 0.214786
R15732 DVSS.n541 DVSS.n540 0.214786
R15733 DVSS.n544 DVSS.n539 0.214786
R15734 DVSS.n545 DVSS.n538 0.214786
R15735 DVSS.n546 DVSS.n537 0.214786
R15736 DVSS.n536 DVSS.n534 0.214786
R15737 DVSS.n550 DVSS.n533 0.214786
R15738 DVSS.n551 DVSS.n532 0.214786
R15739 DVSS.n552 DVSS.n531 0.214786
R15740 DVSS.n530 DVSS.n528 0.214786
R15741 DVSS.n556 DVSS.n527 0.214786
R15742 DVSS.n557 DVSS.n526 0.214786
R15743 DVSS.n558 DVSS.n525 0.214786
R15744 DVSS.n524 DVSS.n522 0.214786
R15745 DVSS.n562 DVSS.n521 0.214786
R15746 DVSS.n563 DVSS.n520 0.214786
R15747 DVSS.n564 DVSS.n519 0.214786
R15748 DVSS.n518 DVSS.n516 0.214786
R15749 DVSS.n568 DVSS.n515 0.214786
R15750 DVSS.n569 DVSS.n514 0.214786
R15751 DVSS.n570 DVSS.n513 0.214786
R15752 DVSS.n206 DVSS.n205 0.214786
R15753 DVSS.n575 DVSS.n574 0.214786
R15754 DVSS.n509 DVSS.n204 0.214786
R15755 DVSS.n508 DVSS.n507 0.214786
R15756 DVSS.n506 DVSS.n208 0.214786
R15757 DVSS.n505 DVSS.n504 0.214786
R15758 DVSS.n499 DVSS.n498 0.214786
R15759 DVSS.n496 DVSS.n211 0.214786
R15760 DVSS.n495 DVSS.n494 0.214786
R15761 DVSS.n213 DVSS.n212 0.214786
R15762 DVSS.n490 DVSS.n489 0.214786
R15763 DVSS.n488 DVSS.n215 0.214786
R15764 DVSS.n487 DVSS.n486 0.214786
R15765 DVSS.n217 DVSS.n216 0.214786
R15766 DVSS.n482 DVSS.n481 0.214786
R15767 DVSS.n480 DVSS.n219 0.214786
R15768 DVSS.n479 DVSS.n478 0.214786
R15769 DVSS.n221 DVSS.n220 0.214786
R15770 DVSS.n474 DVSS.n473 0.214786
R15771 DVSS.n472 DVSS.n223 0.214786
R15772 DVSS.n471 DVSS.n470 0.214786
R15773 DVSS.n225 DVSS.n224 0.214786
R15774 DVSS.n466 DVSS.n465 0.214786
R15775 DVSS.n367 DVSS.n366 0.214786
R15776 DVSS.n5563 DVSS.n825 0.214786
R15777 DVSS.n5565 DVSS.n5564 0.214786
R15778 DVSS.n5566 DVSS.n820 0.214786
R15779 DVSS.n5568 DVSS.n5567 0.214786
R15780 DVSS.n5569 DVSS.n819 0.214786
R15781 DVSS.n5571 DVSS.n5570 0.214786
R15782 DVSS.n5572 DVSS.n814 0.214786
R15783 DVSS.n5574 DVSS.n5573 0.214786
R15784 DVSS.n5575 DVSS.n813 0.214786
R15785 DVSS.n5577 DVSS.n5576 0.214786
R15786 DVSS.n5578 DVSS.n808 0.214786
R15787 DVSS.n5580 DVSS.n5579 0.214786
R15788 DVSS.n5581 DVSS.n807 0.214786
R15789 DVSS.n5583 DVSS.n5582 0.214786
R15790 DVSS.n5586 DVSS.n5585 0.214786
R15791 DVSS.n5587 DVSS.n752 0.214786
R15792 DVSS.n5589 DVSS.n5588 0.214786
R15793 DVSS.n5590 DVSS.n747 0.214786
R15794 DVSS.n5592 DVSS.n5591 0.214786
R15795 DVSS.n5593 DVSS.n746 0.214786
R15796 DVSS.n5595 DVSS.n5594 0.214786
R15797 DVSS.n5596 DVSS.n741 0.214786
R15798 DVSS.n5598 DVSS.n5597 0.214786
R15799 DVSS.n5599 DVSS.n740 0.214786
R15800 DVSS.n5601 DVSS.n5600 0.214786
R15801 DVSS.n5602 DVSS.n735 0.214786
R15802 DVSS.n5604 DVSS.n5603 0.214786
R15803 DVSS.n5605 DVSS.n734 0.214786
R15804 DVSS.n5607 DVSS.n5606 0.214786
R15805 DVSS.n5608 DVSS.n730 0.214786
R15806 DVSS.n5610 DVSS.n5609 0.214786
R15807 DVSS.n5611 DVSS.n147 0.214786
R15808 DVSS.n5613 DVSS.n5612 0.214786
R15809 DVSS.n729 DVSS.n146 0.214786
R15810 DVSS.n728 DVSS.n727 0.214786
R15811 DVSS.n149 DVSS.n148 0.214786
R15812 DVSS.n723 DVSS.n722 0.214786
R15813 DVSS.n721 DVSS.n151 0.214786
R15814 DVSS.n719 DVSS.n718 0.214786
R15815 DVSS.n153 DVSS.n152 0.214786
R15816 DVSS.n542 DVSS.n541 0.214786
R15817 DVSS.n544 DVSS.n543 0.214786
R15818 DVSS.n545 DVSS.n535 0.214786
R15819 DVSS.n547 DVSS.n546 0.214786
R15820 DVSS.n548 DVSS.n534 0.214786
R15821 DVSS.n550 DVSS.n549 0.214786
R15822 DVSS.n551 DVSS.n529 0.214786
R15823 DVSS.n553 DVSS.n552 0.214786
R15824 DVSS.n554 DVSS.n528 0.214786
R15825 DVSS.n556 DVSS.n555 0.214786
R15826 DVSS.n557 DVSS.n523 0.214786
R15827 DVSS.n559 DVSS.n558 0.214786
R15828 DVSS.n560 DVSS.n522 0.214786
R15829 DVSS.n562 DVSS.n561 0.214786
R15830 DVSS.n563 DVSS.n517 0.214786
R15831 DVSS.n565 DVSS.n564 0.214786
R15832 DVSS.n566 DVSS.n516 0.214786
R15833 DVSS.n568 DVSS.n567 0.214786
R15834 DVSS.n569 DVSS.n512 0.214786
R15835 DVSS.n571 DVSS.n570 0.214786
R15836 DVSS.n572 DVSS.n206 0.214786
R15837 DVSS.n574 DVSS.n573 0.214786
R15838 DVSS.n510 DVSS.n509 0.214786
R15839 DVSS.n508 DVSS.n207 0.214786
R15840 DVSS.n502 DVSS.n208 0.214786
R15841 DVSS.n504 DVSS.n503 0.214786
R15842 DVSS.n501 DVSS.n209 0.214786
R15843 DVSS.n500 DVSS.n499 0.214786
R15844 DVSS.n211 DVSS.n210 0.214786
R15845 DVSS.n494 DVSS.n493 0.214786
R15846 DVSS.n492 DVSS.n213 0.214786
R15847 DVSS.n491 DVSS.n490 0.214786
R15848 DVSS.n215 DVSS.n214 0.214786
R15849 DVSS.n486 DVSS.n485 0.214786
R15850 DVSS.n484 DVSS.n217 0.214786
R15851 DVSS.n483 DVSS.n482 0.214786
R15852 DVSS.n219 DVSS.n218 0.214786
R15853 DVSS.n478 DVSS.n477 0.214786
R15854 DVSS.n476 DVSS.n221 0.214786
R15855 DVSS.n475 DVSS.n474 0.214786
R15856 DVSS.n223 DVSS.n222 0.214786
R15857 DVSS.n470 DVSS.n469 0.214786
R15858 DVSS.n468 DVSS.n225 0.214786
R15859 DVSS.n467 DVSS.n466 0.214786
R15860 DVSS.n368 DVSS.n367 0.214786
R15861 DVSS.n227 DVSS.n226 0.214786
R15862 DVSS.n228 DVSS.n227 0.214786
R15863 DVSS.n5 DVSS.n3 0.214786
R15864 DVSS.n4 DVSS.n2 0.214786
R15865 DVSS.n5817 DVSS.n1 0.214786
R15866 DVSS.n5756 DVSS.n0 0.214786
R15867 DVSS.n5760 DVSS.n5757 0.214786
R15868 DVSS.n5761 DVSS.n5755 0.214786
R15869 DVSS.n5762 DVSS.n5754 0.214786
R15870 DVSS.n5753 DVSS.n5751 0.214786
R15871 DVSS.n5766 DVSS.n5750 0.214786
R15872 DVSS.n5767 DVSS.n5749 0.214786
R15873 DVSS.n5768 DVSS.n5748 0.214786
R15874 DVSS.n5747 DVSS.n5745 0.214786
R15875 DVSS.n5772 DVSS.n5744 0.214786
R15876 DVSS.n5773 DVSS.n5743 0.214786
R15877 DVSS.n5774 DVSS.n5742 0.214786
R15878 DVSS.n5740 DVSS.n5739 0.214786
R15879 DVSS.n5738 DVSS.n50 0.214786
R15880 DVSS.n54 DVSS.n49 0.214786
R15881 DVSS.n5734 DVSS.n5733 0.214786
R15882 DVSS.n53 DVSS.n52 0.214786
R15883 DVSS.n5637 DVSS.n5636 0.214786
R15884 DVSS.n5635 DVSS.n5634 0.214786
R15885 DVSS.n5641 DVSS.n5633 0.214786
R15886 DVSS.n5642 DVSS.n5632 0.214786
R15887 DVSS.n5643 DVSS.n5631 0.214786
R15888 DVSS.n5630 DVSS.n5628 0.214786
R15889 DVSS.n5647 DVSS.n5627 0.214786
R15890 DVSS.n5648 DVSS.n5626 0.214786
R15891 DVSS.n5649 DVSS.n5625 0.214786
R15892 DVSS.n5624 DVSS.n5622 0.214786
R15893 DVSS.n5653 DVSS.n5621 0.214786
R15894 DVSS.n5654 DVSS.n5620 0.214786
R15895 DVSS.n5655 DVSS.n5619 0.214786
R15896 DVSS.n5618 DVSS.n142 0.214786
R15897 DVSS.n5659 DVSS.n141 0.214786
R15898 DVSS.n5660 DVSS.n140 0.214786
R15899 DVSS.n5661 DVSS.n139 0.214786
R15900 DVSS.n138 DVSS.n136 0.214786
R15901 DVSS.n5665 DVSS.n135 0.214786
R15902 DVSS.n714 DVSS.n134 0.214786
R15903 DVSS.n713 DVSS.n712 0.214786
R15904 DVSS.n157 DVSS.n156 0.214786
R15905 DVSS.n707 DVSS.n706 0.214786
R15906 DVSS.n705 DVSS.n159 0.214786
R15907 DVSS.n704 DVSS.n703 0.214786
R15908 DVSS.n161 DVSS.n160 0.214786
R15909 DVSS.n699 DVSS.n698 0.214786
R15910 DVSS.n697 DVSS.n163 0.214786
R15911 DVSS.n696 DVSS.n695 0.214786
R15912 DVSS.n165 DVSS.n164 0.214786
R15913 DVSS.n691 DVSS.n690 0.214786
R15914 DVSS.n168 DVSS.n167 0.214786
R15915 DVSS.n594 DVSS.n593 0.214786
R15916 DVSS.n592 DVSS.n591 0.214786
R15917 DVSS.n598 DVSS.n590 0.214786
R15918 DVSS.n599 DVSS.n589 0.214786
R15919 DVSS.n600 DVSS.n588 0.214786
R15920 DVSS.n587 DVSS.n585 0.214786
R15921 DVSS.n604 DVSS.n584 0.214786
R15922 DVSS.n605 DVSS.n583 0.214786
R15923 DVSS.n606 DVSS.n582 0.214786
R15924 DVSS.n581 DVSS.n579 0.214786
R15925 DVSS.n610 DVSS.n578 0.214786
R15926 DVSS.n612 DVSS.n202 0.214786
R15927 DVSS.n613 DVSS.n201 0.214786
R15928 DVSS.n198 DVSS.n196 0.214786
R15929 DVSS.n618 DVSS.n617 0.214786
R15930 DVSS.n197 DVSS.n195 0.214786
R15931 DVSS.n396 DVSS.n395 0.214786
R15932 DVSS.n399 DVSS.n394 0.214786
R15933 DVSS.n400 DVSS.n393 0.214786
R15934 DVSS.n401 DVSS.n392 0.214786
R15935 DVSS.n391 DVSS.n389 0.214786
R15936 DVSS.n405 DVSS.n388 0.214786
R15937 DVSS.n406 DVSS.n387 0.214786
R15938 DVSS.n407 DVSS.n386 0.214786
R15939 DVSS.n385 DVSS.n383 0.214786
R15940 DVSS.n411 DVSS.n382 0.214786
R15941 DVSS.n412 DVSS.n381 0.214786
R15942 DVSS.n413 DVSS.n380 0.214786
R15943 DVSS.n379 DVSS.n377 0.214786
R15944 DVSS.n417 DVSS.n376 0.214786
R15945 DVSS.n418 DVSS.n375 0.214786
R15946 DVSS.n419 DVSS.n374 0.214786
R15947 DVSS.n246 DVSS.n244 0.214786
R15948 DVSS.n424 DVSS.n423 0.214786
R15949 DVSS.n245 DVSS.n243 0.214786
R15950 DVSS.n5815 DVSS.n2 0.214786
R15951 DVSS.n5817 DVSS.n5816 0.214786
R15952 DVSS.n5758 DVSS.n0 0.214786
R15953 DVSS.n5760 DVSS.n5759 0.214786
R15954 DVSS.n5761 DVSS.n5752 0.214786
R15955 DVSS.n5763 DVSS.n5762 0.214786
R15956 DVSS.n5764 DVSS.n5751 0.214786
R15957 DVSS.n5766 DVSS.n5765 0.214786
R15958 DVSS.n5767 DVSS.n5746 0.214786
R15959 DVSS.n5769 DVSS.n5768 0.214786
R15960 DVSS.n5770 DVSS.n5745 0.214786
R15961 DVSS.n5772 DVSS.n5771 0.214786
R15962 DVSS.n5773 DVSS.n45 0.214786
R15963 DVSS.n5775 DVSS.n5774 0.214786
R15964 DVSS.n5739 DVSS.n44 0.214786
R15965 DVSS.n5738 DVSS.n5737 0.214786
R15966 DVSS.n5736 DVSS.n49 0.214786
R15967 DVSS.n5735 DVSS.n5734 0.214786
R15968 DVSS.n52 DVSS.n51 0.214786
R15969 DVSS.n5638 DVSS.n5637 0.214786
R15970 DVSS.n5639 DVSS.n5634 0.214786
R15971 DVSS.n5641 DVSS.n5640 0.214786
R15972 DVSS.n5642 DVSS.n5629 0.214786
R15973 DVSS.n5644 DVSS.n5643 0.214786
R15974 DVSS.n5645 DVSS.n5628 0.214786
R15975 DVSS.n5647 DVSS.n5646 0.214786
R15976 DVSS.n5648 DVSS.n5623 0.214786
R15977 DVSS.n5650 DVSS.n5649 0.214786
R15978 DVSS.n5651 DVSS.n5622 0.214786
R15979 DVSS.n5653 DVSS.n5652 0.214786
R15980 DVSS.n5654 DVSS.n143 0.214786
R15981 DVSS.n5656 DVSS.n5655 0.214786
R15982 DVSS.n5657 DVSS.n142 0.214786
R15983 DVSS.n5659 DVSS.n5658 0.214786
R15984 DVSS.n5660 DVSS.n137 0.214786
R15985 DVSS.n5662 DVSS.n5661 0.214786
R15986 DVSS.n5663 DVSS.n136 0.214786
R15987 DVSS.n5665 DVSS.n5664 0.214786
R15988 DVSS.n710 DVSS.n134 0.214786
R15989 DVSS.n712 DVSS.n711 0.214786
R15990 DVSS.n709 DVSS.n157 0.214786
R15991 DVSS.n708 DVSS.n707 0.214786
R15992 DVSS.n159 DVSS.n158 0.214786
R15993 DVSS.n703 DVSS.n702 0.214786
R15994 DVSS.n701 DVSS.n161 0.214786
R15995 DVSS.n700 DVSS.n699 0.214786
R15996 DVSS.n163 DVSS.n162 0.214786
R15997 DVSS.n695 DVSS.n694 0.214786
R15998 DVSS.n693 DVSS.n165 0.214786
R15999 DVSS.n692 DVSS.n691 0.214786
R16000 DVSS.n167 DVSS.n166 0.214786
R16001 DVSS.n595 DVSS.n594 0.214786
R16002 DVSS.n596 DVSS.n591 0.214786
R16003 DVSS.n598 DVSS.n597 0.214786
R16004 DVSS.n599 DVSS.n586 0.214786
R16005 DVSS.n601 DVSS.n600 0.214786
R16006 DVSS.n602 DVSS.n585 0.214786
R16007 DVSS.n604 DVSS.n603 0.214786
R16008 DVSS.n605 DVSS.n580 0.214786
R16009 DVSS.n607 DVSS.n606 0.214786
R16010 DVSS.n608 DVSS.n579 0.214786
R16011 DVSS.n610 DVSS.n609 0.214786
R16012 DVSS.n612 DVSS.n200 0.214786
R16013 DVSS.n614 DVSS.n613 0.214786
R16014 DVSS.n615 DVSS.n198 0.214786
R16015 DVSS.n617 DVSS.n616 0.214786
R16016 DVSS.n199 DVSS.n197 0.214786
R16017 DVSS.n397 DVSS.n396 0.214786
R16018 DVSS.n399 DVSS.n398 0.214786
R16019 DVSS.n400 DVSS.n390 0.214786
R16020 DVSS.n402 DVSS.n401 0.214786
R16021 DVSS.n403 DVSS.n389 0.214786
R16022 DVSS.n405 DVSS.n404 0.214786
R16023 DVSS.n406 DVSS.n384 0.214786
R16024 DVSS.n408 DVSS.n407 0.214786
R16025 DVSS.n409 DVSS.n383 0.214786
R16026 DVSS.n411 DVSS.n410 0.214786
R16027 DVSS.n412 DVSS.n378 0.214786
R16028 DVSS.n414 DVSS.n413 0.214786
R16029 DVSS.n415 DVSS.n377 0.214786
R16030 DVSS.n417 DVSS.n416 0.214786
R16031 DVSS.n418 DVSS.n372 0.214786
R16032 DVSS.n420 DVSS.n419 0.214786
R16033 DVSS.n421 DVSS.n246 0.214786
R16034 DVSS.n423 DVSS.n422 0.214786
R16035 DVSS.n371 DVSS.n245 0.214786
R16036 DVSS.n27 DVSS.n26 0.214786
R16037 DVSS.n5806 DVSS.n5805 0.214786
R16038 DVSS.n5804 DVSS.n29 0.214786
R16039 DVSS.n5803 DVSS.n5802 0.214786
R16040 DVSS.n5799 DVSS.n5798 0.214786
R16041 DVSS.n5797 DVSS.n31 0.214786
R16042 DVSS.n5796 DVSS.n5795 0.214786
R16043 DVSS.n33 DVSS.n32 0.214786
R16044 DVSS.n5791 DVSS.n5790 0.214786
R16045 DVSS.n5789 DVSS.n35 0.214786
R16046 DVSS.n5788 DVSS.n5787 0.214786
R16047 DVSS.n37 DVSS.n36 0.214786
R16048 DVSS.n5783 DVSS.n5782 0.214786
R16049 DVSS.n5781 DVSS.n39 0.214786
R16050 DVSS.n5780 DVSS.n5779 0.214786
R16051 DVSS.n107 DVSS.n106 0.214786
R16052 DVSS.n108 DVSS.n103 0.214786
R16053 DVSS.n5716 DVSS.n5715 0.214786
R16054 DVSS.n104 DVSS.n102 0.214786
R16055 DVSS.n5710 DVSS.n5709 0.214786
R16056 DVSS.n5708 DVSS.n110 0.214786
R16057 DVSS.n5707 DVSS.n5706 0.214786
R16058 DVSS.n112 DVSS.n111 0.214786
R16059 DVSS.n5702 DVSS.n5701 0.214786
R16060 DVSS.n5700 DVSS.n114 0.214786
R16061 DVSS.n5699 DVSS.n5698 0.214786
R16062 DVSS.n116 DVSS.n115 0.214786
R16063 DVSS.n5694 DVSS.n5693 0.214786
R16064 DVSS.n5692 DVSS.n118 0.214786
R16065 DVSS.n5691 DVSS.n5690 0.214786
R16066 DVSS.n120 DVSS.n119 0.214786
R16067 DVSS.n5686 DVSS.n5685 0.214786
R16068 DVSS.n5684 DVSS.n122 0.214786
R16069 DVSS.n5683 DVSS.n5682 0.214786
R16070 DVSS.n5676 DVSS.n124 0.214786
R16071 DVSS.n5678 DVSS.n5677 0.214786
R16072 DVSS.n5675 DVSS.n126 0.214786
R16073 DVSS.n5674 DVSS.n5673 0.214786
R16074 DVSS.n128 DVSS.n127 0.214786
R16075 DVSS.n5668 DVSS.n132 0.214786
R16076 DVSS.n668 DVSS.n131 0.214786
R16077 DVSS.n670 DVSS.n669 0.214786
R16078 DVSS.n673 DVSS.n667 0.214786
R16079 DVSS.n674 DVSS.n666 0.214786
R16080 DVSS.n675 DVSS.n665 0.214786
R16081 DVSS.n664 DVSS.n662 0.214786
R16082 DVSS.n679 DVSS.n661 0.214786
R16083 DVSS.n680 DVSS.n660 0.214786
R16084 DVSS.n681 DVSS.n659 0.214786
R16085 DVSS.n173 DVSS.n171 0.214786
R16086 DVSS.n686 DVSS.n685 0.214786
R16087 DVSS.n172 DVSS.n170 0.214786
R16088 DVSS.n655 DVSS.n654 0.214786
R16089 DVSS.n653 DVSS.n175 0.214786
R16090 DVSS.n652 DVSS.n651 0.214786
R16091 DVSS.n177 DVSS.n176 0.214786
R16092 DVSS.n647 DVSS.n646 0.214786
R16093 DVSS.n645 DVSS.n179 0.214786
R16094 DVSS.n644 DVSS.n643 0.214786
R16095 DVSS.n181 DVSS.n180 0.214786
R16096 DVSS.n639 DVSS.n638 0.214786
R16097 DVSS.n637 DVSS.n183 0.214786
R16098 DVSS.n636 DVSS.n635 0.214786
R16099 DVSS.n631 DVSS.n630 0.214786
R16100 DVSS.n629 DVSS.n188 0.214786
R16101 DVSS.n628 DVSS.n627 0.214786
R16102 DVSS.n190 DVSS.n189 0.214786
R16103 DVSS.n623 DVSS.n622 0.214786
R16104 DVSS.n193 DVSS.n192 0.214786
R16105 DVSS.n333 DVSS.n332 0.214786
R16106 DVSS.n336 DVSS.n331 0.214786
R16107 DVSS.n337 DVSS.n330 0.214786
R16108 DVSS.n338 DVSS.n329 0.214786
R16109 DVSS.n328 DVSS.n326 0.214786
R16110 DVSS.n342 DVSS.n325 0.214786
R16111 DVSS.n343 DVSS.n324 0.214786
R16112 DVSS.n344 DVSS.n323 0.214786
R16113 DVSS.n322 DVSS.n320 0.214786
R16114 DVSS.n348 DVSS.n319 0.214786
R16115 DVSS.n349 DVSS.n318 0.214786
R16116 DVSS.n350 DVSS.n317 0.214786
R16117 DVSS.n316 DVSS.n314 0.214786
R16118 DVSS.n354 DVSS.n313 0.214786
R16119 DVSS.n355 DVSS.n312 0.214786
R16120 DVSS.n356 DVSS.n258 0.214786
R16121 DVSS.n257 DVSS.n255 0.214786
R16122 DVSS.n361 DVSS.n360 0.214786
R16123 DVSS.n5807 DVSS.n5806 0.214786
R16124 DVSS.n29 DVSS.n28 0.214786
R16125 DVSS.n5802 DVSS.n5801 0.214786
R16126 DVSS.n5800 DVSS.n5799 0.214786
R16127 DVSS.n31 DVSS.n30 0.214786
R16128 DVSS.n5795 DVSS.n5794 0.214786
R16129 DVSS.n5793 DVSS.n33 0.214786
R16130 DVSS.n5792 DVSS.n5791 0.214786
R16131 DVSS.n35 DVSS.n34 0.214786
R16132 DVSS.n5787 DVSS.n5786 0.214786
R16133 DVSS.n5785 DVSS.n37 0.214786
R16134 DVSS.n5784 DVSS.n5783 0.214786
R16135 DVSS.n39 DVSS.n38 0.214786
R16136 DVSS.n5779 DVSS.n5778 0.214786
R16137 DVSS.n107 DVSS.n42 0.214786
R16138 DVSS.n5713 DVSS.n108 0.214786
R16139 DVSS.n5715 DVSS.n5714 0.214786
R16140 DVSS.n5712 DVSS.n104 0.214786
R16141 DVSS.n5711 DVSS.n5710 0.214786
R16142 DVSS.n110 DVSS.n109 0.214786
R16143 DVSS.n5706 DVSS.n5705 0.214786
R16144 DVSS.n5704 DVSS.n112 0.214786
R16145 DVSS.n5703 DVSS.n5702 0.214786
R16146 DVSS.n114 DVSS.n113 0.214786
R16147 DVSS.n5698 DVSS.n5697 0.214786
R16148 DVSS.n5696 DVSS.n116 0.214786
R16149 DVSS.n5695 DVSS.n5694 0.214786
R16150 DVSS.n118 DVSS.n117 0.214786
R16151 DVSS.n5690 DVSS.n5689 0.214786
R16152 DVSS.n5688 DVSS.n120 0.214786
R16153 DVSS.n5687 DVSS.n5686 0.214786
R16154 DVSS.n122 DVSS.n121 0.214786
R16155 DVSS.n5682 DVSS.n5681 0.214786
R16156 DVSS.n5680 DVSS.n124 0.214786
R16157 DVSS.n5679 DVSS.n5678 0.214786
R16158 DVSS.n126 DVSS.n125 0.214786
R16159 DVSS.n5673 DVSS.n5672 0.214786
R16160 DVSS.n5671 DVSS.n128 0.214786
R16161 DVSS.n5669 DVSS.n5668 0.214786
R16162 DVSS.n131 DVSS.n130 0.214786
R16163 DVSS.n671 DVSS.n670 0.214786
R16164 DVSS.n673 DVSS.n672 0.214786
R16165 DVSS.n674 DVSS.n663 0.214786
R16166 DVSS.n676 DVSS.n675 0.214786
R16167 DVSS.n677 DVSS.n662 0.214786
R16168 DVSS.n679 DVSS.n678 0.214786
R16169 DVSS.n680 DVSS.n658 0.214786
R16170 DVSS.n682 DVSS.n681 0.214786
R16171 DVSS.n683 DVSS.n173 0.214786
R16172 DVSS.n685 DVSS.n684 0.214786
R16173 DVSS.n657 DVSS.n172 0.214786
R16174 DVSS.n656 DVSS.n655 0.214786
R16175 DVSS.n175 DVSS.n174 0.214786
R16176 DVSS.n651 DVSS.n650 0.214786
R16177 DVSS.n649 DVSS.n177 0.214786
R16178 DVSS.n648 DVSS.n647 0.214786
R16179 DVSS.n179 DVSS.n178 0.214786
R16180 DVSS.n643 DVSS.n642 0.214786
R16181 DVSS.n641 DVSS.n181 0.214786
R16182 DVSS.n640 DVSS.n639 0.214786
R16183 DVSS.n183 DVSS.n182 0.214786
R16184 DVSS.n635 DVSS.n634 0.214786
R16185 DVSS.n632 DVSS.n631 0.214786
R16186 DVSS.n188 DVSS.n187 0.214786
R16187 DVSS.n627 DVSS.n626 0.214786
R16188 DVSS.n625 DVSS.n190 0.214786
R16189 DVSS.n624 DVSS.n623 0.214786
R16190 DVSS.n192 DVSS.n191 0.214786
R16191 DVSS.n334 DVSS.n333 0.214786
R16192 DVSS.n336 DVSS.n335 0.214786
R16193 DVSS.n337 DVSS.n327 0.214786
R16194 DVSS.n339 DVSS.n338 0.214786
R16195 DVSS.n340 DVSS.n326 0.214786
R16196 DVSS.n342 DVSS.n341 0.214786
R16197 DVSS.n343 DVSS.n321 0.214786
R16198 DVSS.n345 DVSS.n344 0.214786
R16199 DVSS.n346 DVSS.n320 0.214786
R16200 DVSS.n348 DVSS.n347 0.214786
R16201 DVSS.n349 DVSS.n315 0.214786
R16202 DVSS.n351 DVSS.n350 0.214786
R16203 DVSS.n352 DVSS.n314 0.214786
R16204 DVSS.n354 DVSS.n353 0.214786
R16205 DVSS.n355 DVSS.n256 0.214786
R16206 DVSS.n357 DVSS.n356 0.214786
R16207 DVSS.n358 DVSS.n255 0.214786
R16208 DVSS.n360 DVSS.n359 0.214786
R16209 DVSS.n4475 DVSS.n1278 0.212265
R16210 DVSS.n1193 DVSS.n1192 0.201836
R16211 DVSS.n3650 DVSS 0.194818
R16212 DVSS.n4484 DVSS.n4483 0.192412
R16213 DVSS.n3576 VSS 0.189765
R16214 VSS DVSS.n3576 0.189765
R16215 DVSS.n3615 DVSS 0.186337
R16216 DVSS.n1476 DVSS.n1475 0.186214
R16217 DVSS.n1477 DVSS.n1476 0.186214
R16218 DVSS.n4381 DVSS.n4376 0.186214
R16219 DVSS.n4383 DVSS.n4381 0.186214
R16220 DVSS.n5359 DVSS.n5358 0.185484
R16221 DVSS.n3947 VSS 0.17855
R16222 DVSS.n3633 DVSS.n1716 0.178408
R16223 DVSS.n3633 DVSS.n3632 0.178408
R16224 DVSS.n3628 DVSS.n3626 0.178408
R16225 DVSS.n3633 DVSS.n3631 0.178408
R16226 DVSS.n3628 DVSS.n3627 0.178408
R16227 DVSS.n3633 DVSS.n3630 0.178408
R16228 DVSS.n3628 DVSS.n1725 0.178408
R16229 DVSS.n1451 DVSS.n1450 0.175807
R16230 DVSS.n1289 DVSS 0.175204
R16231 DVSS.n1294 DVSS 0.175204
R16232 DVSS.n4380 DVSS 0.175204
R16233 DVSS.n1314 DVSS 0.175204
R16234 DVSS.n5718 DVSS.n5717 0.173577
R16235 DVSS.n311 DVSS.n310 0.173577
R16236 VSS DVSS.n3941 0.169912
R16237 DVSS.n5057 DVSS.n5056 0.168658
R16238 DVSS.n5056 DVSS.n1112 0.168658
R16239 DVSS.n5046 DVSS.n1120 0.168658
R16240 DVSS.n5046 DVSS.n5045 0.168658
R16241 DVSS.n1479 DVSS.n1444 0.166289
R16242 DVSS.n5617 DVSS.n5616 0.163909
R16243 DVSS.n689 DVSS.n688 0.163909
R16244 DVSS.n620 DVSS.n619 0.163909
R16245 DVSS.n427 DVSS.n241 0.161214
R16246 DVSS.n765 DVSS.n57 0.161214
R16247 DVSS.n5559 DVSS.n5557 0.149124
R16248 DVSS.n2250 DVSS.n1519 0.145461
R16249 DVSS.n3397 DVSS 0.144526
R16250 DVSS DVSS.n1506 0.1436
R16251 DVSS.n1509 DVSS 0.1436
R16252 DVSS DVSS.n1509 0.1436
R16253 DVSS.n1513 DVSS 0.1436
R16254 DVSS DVSS.n3765 0.143441
R16255 DVSS.n1672 DVSS 0.143441
R16256 DVSS DVSS.n3900 0.143441
R16257 DVSS.n3898 DVSS 0.143441
R16258 DVSS.n802 DVSS.n801 0.141125
R16259 DVSS.n464 DVSS.n463 0.141125
R16260 DVSS.n3765 DVSS.n1660 0.140794
R16261 DVSS.n1672 DVSS.n1660 0.140794
R16262 DVSS.n3900 DVSS.n3899 0.140794
R16263 DVSS.n3899 DVSS.n3898 0.140794
R16264 DVSS.n3577 VSS 0.139932
R16265 DVSS.n2232 DVSS 0.138622
R16266 DVSS.n803 DVSS.n754 0.137596
R16267 DVSS.n461 DVSS.n229 0.137559
R16268 DVSS.n1733 DVSS 0.1355
R16269 DVSS DVSS.n1299 0.1355
R16270 DVSS.n5722 DVSS.n61 0.130943
R16271 DVSS.n2023 DVSS 0.130618
R16272 DVSS.n260 DVSS.n60 0.130587
R16273 DVSS.n4037 DVSS 0.130161
R16274 DVSS.n3728 DVSS 0.130161
R16275 DVSS.n1658 DVSS.n1657 0.129687
R16276 DVSS.n3768 DVSS.n1689 0.129687
R16277 DVSS.n1693 DVSS.n1692 0.129687
R16278 DVSS.n3764 DVSS.n3763 0.129687
R16279 DVSS.n1673 DVSS.n1671 0.129687
R16280 DVSS.n3792 DVSS.n1656 0.129687
R16281 DVSS.n3857 DVSS.n3856 0.129687
R16282 DVSS.n1577 DVSS.n1576 0.129687
R16283 DVSS.n1579 DVSS.n1578 0.129687
R16284 DVSS.n1582 DVSS.n1581 0.129687
R16285 DVSS.n1585 DVSS.n1584 0.129687
R16286 DVSS.n3895 DVSS.n1589 0.129687
R16287 DVSS.n955 DVSS.n954 0.129009
R16288 DVSS.n1925 DVSS.n1813 0.128608
R16289 DVSS.n2152 DVSS.n1925 0.128203
R16290 DVSS DVSS.n856 0.125798
R16291 DVSS.n3652 DVSS.n1703 0.122865
R16292 DVSS.n856 DVSS.n855 0.12265
R16293 DVSS.n2240 DVSS 0.122025
R16294 DVSS DVSS.n3619 0.115647
R16295 DVSS.n1816 DVSS.n1815 0.114824
R16296 DVSS.n2153 DVSS.n1807 0.114824
R16297 DVSS.n5808 DVSS.n5807 0.114699
R16298 DVSS.n5815 DVSS.n5814 0.114699
R16299 DVSS.n5563 DVSS.n5562 0.114699
R16300 DVSS.n4425 DVSS.n4424 0.114184
R16301 DVSS.n1470 DVSS.n1469 0.114184
R16302 DVSS.n4188 DVSS.n4187 0.114184
R16303 DVSS.n4391 DVSS.n4390 0.114184
R16304 DVSS.n4339 DVSS.n4338 0.114184
R16305 DVSS.n2257 VSS 0.113
R16306 DVSS.n3571 VSS 0.113
R16307 VSS DVSS.n1697 0.113
R16308 DVSS.n3397 DVSS 0.111845
R16309 DVSS.n3955 DVSS 0.111373
R16310 DVSS.n4937 DVSS.n1176 0.110634
R16311 DVSS.n3561 VSS 0.110353
R16312 DVSS.n2164 DVSS.n1786 0.109959
R16313 DVSS.n2165 DVSS.n2164 0.109959
R16314 DVSS.n3953 DVSS.n3952 0.109729
R16315 DVSS.n1512 DVSS.n1510 0.109572
R16316 DVSS.n5732 DVSS.n5731 0.107643
R16317 DVSS.n373 DVSS.n242 0.107643
R16318 DVSS.n3955 DVSS 0.107291
R16319 DVSS.n1443 DVSS.n1112 0.107079
R16320 DVSS.n1467 DVSS.n1466 0.105895
R16321 DVSS.n954 DVSS.n949 0.102277
R16322 DVSS.n1509 DVSS 0.102157
R16323 DVSS.n5352 DVSS.n5351 0.101471
R16324 DVSS.n5112 DVSS.n5111 0.101471
R16325 DVSS DVSS.n4037 0.101206
R16326 DVSS DVSS.n3728 0.101206
R16327 DVSS DVSS.n2023 0.10093
R16328 DVSS.n3652 DVSS.n3651 0.100254
R16329 DVSS.n3954 DVSS 0.0991804
R16330 DVSS.n5360 DVSS.n5359 0.0985668
R16331 DVSS.n5359 DVSS.n952 0.0982447
R16332 DVSS.n3746 DVSS.n1705 0.0951262
R16333 DVSS.n1161 DVSS 0.0942039
R16334 DVSS.n1298 DVSS 0.0942039
R16335 DVSS.n4450 DVSS 0.0942039
R16336 DVSS.n4959 DVSS 0.0942039
R16337 DVSS DVSS.n3650 0.0938582
R16338 VSS DVSS.n1444 0.0928684
R16339 DVSS.n2804 DVSS.n2803 0.0923483
R16340 DVSS.n4483 DVSS.n4482 0.0891765
R16341 DVSS.n3981 DVSS.n3980 0.0883604
R16342 DVSS.n3605 DVSS 0.0871834
R16343 DVSS.n3606 DVSS 0.0871834
R16344 DVSS.n3955 DVSS 0.0837012
R16345 DVSS.n1861 DVSS.n1440 0.08175
R16346 DVSS.n3987 DVSS.n3986 0.08175
R16347 DVSS DVSS.n4451 0.0812353
R16348 DVSS DVSS.n4960 0.0812353
R16349 DVSS DVSS.n1162 0.0812353
R16350 DVSS.n2146 DVSS.n1796 0.077375
R16351 DVSS.n2180 DVSS.n1788 0.077375
R16352 DVSS DVSS.n4475 0.0772647
R16353 DVSS.n3604 DVSS.n3602 0.0769706
R16354 DVSS.n3604 DVSS.n3603 0.0769706
R16355 DVSS.n1597 DVSS.n1594 0.0766156
R16356 DVSS.n1868 DVSS.n1811 0.0763777
R16357 DVSS DVSS.n3206 0.0761
R16358 DVSS.n3346 DVSS 0.0761
R16359 DVSS.n3483 DVSS 0.0761
R16360 DVSS.n3247 DVSS 0.0761
R16361 DVSS DVSS.n3250 0.0761
R16362 DVSS.n3251 DVSS 0.0761
R16363 DVSS.n3058 DVSS 0.0761
R16364 DVSS.n3554 DVSS 0.0761
R16365 DVSS.n2991 DVSS 0.0761
R16366 DVSS DVSS.n2709 0.0761
R16367 DVSS DVSS.n2746 0.0761
R16368 DVSS.n2871 DVSS 0.0761
R16369 DVSS DVSS.n2779 0.0761
R16370 DVSS.n2826 DVSS 0.0761
R16371 DVSS.n1880 DVSS.n1868 0.0756596
R16372 DVSS DVSS.n1506 0.0748392
R16373 DVSS DVSS.n1513 0.0746758
R16374 DVSS.n2805 DVSS.n2804 0.07437
R16375 DVSS.n3612 DVSS 0.0743218
R16376 DVSS.n3610 DVSS 0.0743218
R16377 DVSS.n4547 DVSS.n4511 0.0741096
R16378 DVSS.n4183 DVSS.n1370 0.0728571
R16379 DVSS DVSS.n1707 0.0720909
R16380 DVSS DVSS.n3614 0.0720477
R16381 DVSS.n2228 DVSS.n1734 0.0693638
R16382 DVSS.n3940 DVSS.n3939 0.0668158
R16383 DVSS.n3948 DVSS.n3947 0.0656316
R16384 DVSS.n3649 DVSS 0.064306
R16385 DVSS.n4548 DVSS.n4547 0.0624601
R16386 DVSS.n1443 DVSS.n1120 0.0620789
R16387 DVSS.n1598 DVSS.n1597 0.0602043
R16388 DVSS.n5556 DVSS.n847 0.0597445
R16389 DVSS.n846 DVSS.n845 0.0597445
R16390 DVSS.n844 DVSS.n843 0.0597445
R16391 DVSS.n842 DVSS.n841 0.0597445
R16392 DVSS.n840 DVSS.n839 0.0597445
R16393 DVSS.n838 DVSS.n837 0.0597445
R16394 DVSS.n836 DVSS.n835 0.0597445
R16395 DVSS.n834 DVSS.n833 0.0597445
R16396 DVSS.n832 DVSS.n831 0.0597445
R16397 DVSS.n5558 DVSS.n830 0.0597445
R16398 DVSS.n25 DVSS.n24 0.0597445
R16399 DVSS.n23 DVSS.n22 0.0597445
R16400 DVSS.n21 DVSS.n20 0.0597445
R16401 DVSS.n19 DVSS.n18 0.0597445
R16402 DVSS.n17 DVSS.n16 0.0597445
R16403 DVSS.n15 DVSS.n14 0.0597445
R16404 DVSS.n13 DVSS.n12 0.0597445
R16405 DVSS.n11 DVSS.n10 0.0597445
R16406 DVSS.n9 DVSS.n8 0.0597445
R16407 DVSS.n5810 DVSS.n7 0.0597445
R16408 DVSS.n24 DVSS.n23 0.0597445
R16409 DVSS.n22 DVSS.n21 0.0597445
R16410 DVSS.n20 DVSS.n19 0.0597445
R16411 DVSS.n18 DVSS.n17 0.0597445
R16412 DVSS.n16 DVSS.n15 0.0597445
R16413 DVSS.n14 DVSS.n13 0.0597445
R16414 DVSS.n12 DVSS.n11 0.0597445
R16415 DVSS.n10 DVSS.n9 0.0597445
R16416 DVSS.n8 DVSS.n7 0.0597445
R16417 DVSS.n847 DVSS.n846 0.0597445
R16418 DVSS.n845 DVSS.n844 0.0597445
R16419 DVSS.n843 DVSS.n842 0.0597445
R16420 DVSS.n841 DVSS.n840 0.0597445
R16421 DVSS.n839 DVSS.n838 0.0597445
R16422 DVSS.n837 DVSS.n836 0.0597445
R16423 DVSS.n835 DVSS.n834 0.0597445
R16424 DVSS.n833 DVSS.n832 0.0597445
R16425 DVSS.n831 DVSS.n830 0.0597445
R16426 DVSS.n4537 DVSS.n4528 0.0588383
R16427 DVSS.n2151 DVSS.n2150 0.058625
R16428 DVSS.n1879 DVSS.n1878 0.058625
R16429 DVSS.n2224 DVSS.n1734 0.0585457
R16430 DVSS DVSS.n4425 0.0585263
R16431 DVSS DVSS.n1470 0.0585263
R16432 DVSS.n4187 DVSS 0.0585263
R16433 DVSS DVSS.n4391 0.0585263
R16434 DVSS.n4338 DVSS 0.0585263
R16435 DVSS.n1372 DVSS.n1370 0.058308
R16436 DVSS DVSS.n3954 0.0574691
R16437 DVSS DVSS.n1703 0.0569179
R16438 DVSS DVSS.n3747 0.0569179
R16439 DVSS.n4820 DVSS.n1215 0.0562784
R16440 DVSS.n1925 DVSS.n1924 0.0546667
R16441 DVSS.n1924 DVSS.t19 0.0546667
R16442 DVSS.n2163 DVSS.t19 0.0546667
R16443 DVSS.n2164 DVSS.n2163 0.0546667
R16444 DVSS.n2148 DVSS.n2147 0.0544368
R16445 DVSS.n2149 DVSS.n2148 0.0544368
R16446 DVSS.n1876 DVSS.n1875 0.0544368
R16447 DVSS.n1876 DVSS.n1869 0.0544368
R16448 DVSS.n364 DVSS.n249 0.0532401
R16449 DVSS.n2208 DVSS.n1748 0.0532027
R16450 DVSS.n2096 DVSS.n2089 0.0532027
R16451 DVSS.n1215 DVSS.n1214 0.0500653
R16452 DVSS.n1864 DVSS.n1863 0.0495566
R16453 DVSS.n3983 DVSS.n3982 0.0495566
R16454 DVSS.n3988 DVSS.n3987 0.0486793
R16455 DVSS.n369 DVSS.n249 0.0485826
R16456 DVSS DVSS.n1508 0.0479398
R16457 DVSS DVSS.n1505 0.0479398
R16458 DVSS.n4468 DVSS 0.0456808
R16459 DVSS.n4470 DVSS 0.0456808
R16460 DVSS.n4474 DVSS 0.0456808
R16461 DVSS.n1657 DVSS 0.0456808
R16462 DVSS.n1689 DVSS 0.0456808
R16463 DVSS.n1692 DVSS 0.0456808
R16464 DVSS.n3763 DVSS 0.0456808
R16465 DVSS.n1671 DVSS 0.0456808
R16466 DVSS.n1656 DVSS 0.0456808
R16467 DVSS.n3856 DVSS 0.0456808
R16468 DVSS.n1576 DVSS 0.0456808
R16469 DVSS.n1578 DVSS 0.0456808
R16470 DVSS.n1581 DVSS 0.0456808
R16471 DVSS.n1584 DVSS 0.0456808
R16472 DVSS.n1589 DVSS 0.0456808
R16473 DVSS.n2135 DVSS.n1934 0.0450872
R16474 DVSS.n1827 DVSS.n1826 0.0450872
R16475 DVSS.n1919 DVSS.n1835 0.0450872
R16476 DVSS.n1780 DVSS.n1778 0.0450872
R16477 DVSS.n2092 DVSS.n1951 0.0450872
R16478 DVSS.n2206 DVSS.n2205 0.0450718
R16479 DVSS.n2205 DVSS.n2204 0.0450718
R16480 DVSS.n1756 DVSS.n1755 0.0450718
R16481 DVSS.n1757 DVSS.n1756 0.0450718
R16482 DVSS.n1947 DVSS.n1946 0.0450718
R16483 DVSS.n1948 DVSS.n1947 0.0450718
R16484 DVSS.n2108 DVSS.n2099 0.0442838
R16485 DVSS.n2158 DVSS.n1808 0.0442838
R16486 DVSS.n2110 DVSS.n2109 0.0442838
R16487 DVSS.n2109 DVSS.n2100 0.0442838
R16488 DVSS.n2103 DVSS.n2102 0.0442838
R16489 DVSS.n1828 DVSS.n1820 0.0442838
R16490 DVSS.n1829 DVSS.n1828 0.0442838
R16491 DVSS.n1834 DVSS.n1833 0.0442838
R16492 DVSS.n2208 DVSS.n2207 0.0442838
R16493 DVSS.n2203 DVSS.n2202 0.0442838
R16494 DVSS.n2202 DVSS.n1751 0.0442838
R16495 DVSS.n1775 DVSS.n1774 0.0442838
R16496 DVSS.n1776 DVSS.n1775 0.0442838
R16497 DVSS.n1781 DVSS.n1776 0.0442838
R16498 DVSS.n1782 DVSS.n1781 0.0442838
R16499 DVSS.n2185 DVSS.n1782 0.0442838
R16500 DVSS.n2185 DVSS.n2184 0.0442838
R16501 DVSS.n2184 DVSS.n1783 0.0442838
R16502 DVSS.n1935 DVSS.n1802 0.0442838
R16503 DVSS.n1939 DVSS.n1935 0.0442838
R16504 DVSS.n1940 DVSS.n1939 0.0442838
R16505 DVSS.n2134 DVSS.n1940 0.0442838
R16506 DVSS.n2134 DVSS.n2133 0.0442838
R16507 DVSS.n2133 DVSS.n2132 0.0442838
R16508 DVSS.n2132 DVSS.n1941 0.0442838
R16509 DVSS.n2128 DVSS.n1949 0.0442838
R16510 DVSS.n2128 DVSS.n2127 0.0442838
R16511 DVSS.n2127 DVSS.n1950 0.0442838
R16512 DVSS.n2091 DVSS.n1950 0.0442838
R16513 DVSS.n2095 DVSS.n2091 0.0442838
R16514 DVSS.n2096 DVSS.n2095 0.0442838
R16515 DVSS.n1440 DVSS.n1390 0.0432989
R16516 DVSS.n2131 DVSS.n1942 0.0430229
R16517 DVSS.n1777 DVSS.n1753 0.0430229
R16518 DVSS.n1830 DVSS.n1819 0.0426101
R16519 DVSS.n2126 DVSS.n2125 0.0421972
R16520 DVSS.n1965 DVSS.n1959 0.0418677
R16521 DVSS.n2198 DVSS.n1760 0.0418677
R16522 DVSS.n2107 DVSS.n2106 0.0418514
R16523 DVSS.n4927 DVSS.n1215 0.0417698
R16524 DVSS.n4927 DVSS.n4926 0.0417698
R16525 DVSS.n4528 DVSS.n4491 0.0417698
R16526 DVSS.n4491 DVSS.n4490 0.0417698
R16527 DVSS.n1938 DVSS.n1936 0.0405459
R16528 DVSS.n2186 DVSS.n1773 0.0405459
R16529 DVSS.n3556 DVSS.n3555 0.0398939
R16530 DVSS.n3557 DVSS.n3556 0.0398939
R16531 DVSS.n2210 DVSS.n2209 0.0397202
R16532 DVSS.n2795 DVSS 0.0392931
R16533 DVSS.n3651 DVSS 0.0392931
R16534 DVSS DVSS.n2797 0.0392931
R16535 DVSS.n2103 DVSS.n1805 0.0382027
R16536 DVSS.n1833 DVSS.n1818 0.0382027
R16537 DVSS.n1868 DVSS.n1867 0.0381812
R16538 DVSS.n1867 DVSS.t19 0.0381812
R16539 DVSS.n2099 DVSS.n2086 0.0373919
R16540 DVSS.n4191 DVSS.n4190 0.0359178
R16541 DVSS.n1860 DVSS.n1437 0.0357988
R16542 DVSS.n1507 DVSS 0.0351916
R16543 DVSS DVSS.n3953 0.0351916
R16544 DVSS.n1514 DVSS 0.0351154
R16545 DVSS.n1510 DVSS 0.0351154
R16546 DVSS.n3078 DVSS.n1701 0.0349371
R16547 DVSS.n2659 DVSS.n1701 0.0349371
R16548 DVSS.n1448 VSS 0.0348421
R16549 DVSS.n2094 DVSS.n2093 0.0339404
R16550 DVSS.n363 DVSS.n248 0.033707
R16551 DVSS.n362 DVSS.n251 0.033707
R16552 DVSS.n4461 DVSS.n4460 0.0336579
R16553 DVSS.n4408 DVSS.n4407 0.0336579
R16554 DVSS.n4377 DVSS.n1315 0.0336579
R16555 DVSS.n4464 DVSS.n4463 0.0336579
R16556 DVSS.n2136 DVSS.n1933 0.0331147
R16557 DVSS.n1779 DVSS.n1772 0.0331147
R16558 DVSS.n4793 DVSS.n1194 0.033
R16559 DVSS.n4924 DVSS.n1194 0.033
R16560 DVSS.n4922 DVSS.n4921 0.033
R16561 DVSS.n4923 DVSS.n4922 0.033
R16562 DVSS.n4718 DVSS.n1217 0.033
R16563 DVSS.n1217 DVSS.n1216 0.033
R16564 DVSS.n4679 DVSS.n4678 0.033
R16565 DVSS.n4678 DVSS.n4677 0.033
R16566 DVSS.n4600 DVSS.n1272 0.033
R16567 DVSS.n4676 DVSS.n1272 0.033
R16568 DVSS.n4674 DVSS.n4673 0.033
R16569 DVSS.n4675 DVSS.n4674 0.033
R16570 DVSS.n4456 DVSS.n1299 0.0322647
R16571 DVSS DVSS.n1709 0.0320421
R16572 DVSS.n2155 DVSS.n1812 0.031778
R16573 DVSS.n1916 DVSS.n1914 0.031778
R16574 DVSS.n2815 DVSS.n2814 0.0315
R16575 DVSS.n2858 DVSS.n2767 0.0315
R16576 DVSS.n2863 DVSS.n2767 0.0315
R16577 DVSS.n2915 DVSS.n2914 0.0315
R16578 DVSS.n2970 DVSS.n2969 0.0315
R16579 DVSS.n3019 DVSS.n2703 0.0315
R16580 DVSS.n3060 DVSS.n2668 0.0315
R16581 DVSS.n3095 DVSS.n3079 0.0315
R16582 DVSS.n3508 DVSS.n3507 0.0315
R16583 DVSS.n3486 DVSS.n3149 0.0315
R16584 DVSS.n3186 DVSS.n3182 0.0315
R16585 DVSS.n3445 DVSS.n3444 0.0315
R16586 DVSS.n3444 DVSS.n3208 0.0315
R16587 DVSS.n3423 DVSS.n3239 0.0315
R16588 DVSS.n2799 DVSS.n2798 0.0315
R16589 DVSS.n2827 DVSS.n2765 0.0315
R16590 DVSS.n2867 DVSS.n2765 0.0315
R16591 DVSS.n2874 DVSS.n2873 0.0315
R16592 DVSS.n2935 DVSS.n2934 0.0315
R16593 DVSS.n3005 DVSS.n3004 0.0315
R16594 DVSS.n3552 DVSS.n2664 0.0315
R16595 DVSS.n3271 DVSS.n3270 0.0315
R16596 DVSS.n3291 DVSS.n3290 0.0315
R16597 DVSS.n3312 DVSS.n3248 0.0315
R16598 DVSS.n3333 DVSS.n3332 0.0315
R16599 DVSS.n3351 DVSS.n3210 0.0315
R16600 DVSS.n3355 DVSS.n3210 0.0315
R16601 DVSS.n3372 DVSS.n3244 0.0315
R16602 DVSS.n1832 DVSS.n1817 0.0310505
R16603 DVSS.n2813 DVSS.n2789 0.031
R16604 DVSS.n2918 DVSS.n2745 0.031
R16605 DVSS.n3185 DVSS.n3170 0.031
R16606 DVSS.n3419 DVSS.n3242 0.031
R16607 DVSS.n2802 DVSS.n2791 0.031
R16608 DVSS.n2922 DVSS.n2743 0.031
R16609 DVSS.n3328 DVSS.n3246 0.031
R16610 DVSS.n3375 DVSS.n3374 0.031
R16611 DVSS.n2102 DVSS.n1807 0.0309054
R16612 DVSS.n1834 DVSS.n1816 0.0309054
R16613 DVSS.n2098 DVSS.n2097 0.0306376
R16614 DVSS.n2104 DVSS.n2101 0.0305
R16615 DVSS.n2973 DVSS.n2723 0.0305
R16616 DVSS.n3487 DVSS.n3148 0.0305
R16617 DVSS.n2931 DVSS.n2926 0.0305
R16618 DVSS.n3308 DVSS.n3145 0.0305
R16619 DVSS.n370 DVSS.n248 0.0304195
R16620 DVSS.n251 DVSS.n247 0.0304195
R16621 DVSS.n2130 DVSS.n2129 0.0302248
R16622 DVSS.n2201 DVSS.n2200 0.0302248
R16623 DVSS.n5557 DVSS.n25 0.0301222
R16624 DVSS.n5811 DVSS.n5810 0.0301222
R16625 DVSS.n5556 DVSS.n5555 0.0301222
R16626 DVSS.n5559 DVSS.n5558 0.0301222
R16627 DVSS.n3650 DVSS.n3649 0.0300522
R16628 DVSS.n3020 DVSS.n2693 0.03
R16629 DVSS.n3511 DVSS.n3113 0.03
R16630 DVSS.n3001 DVSS.n2702 0.03
R16631 DVSS.n3289 DVSS.n3287 0.03
R16632 DVSS.n4192 DVSS.n4191 0.0298971
R16633 DVSS.n3549 DVSS.n3548 0.0295
R16634 DVSS.n3532 DVSS.n3531 0.0295
R16635 DVSS.n3551 DVSS.n2665 0.0295
R16636 DVSS.n3267 DVSS.n3081 0.0295
R16637 DVSS.n3061 DVSS.n2682 0.029
R16638 DVSS.n3094 DVSS.n3091 0.029
R16639 DVSS.n3046 DVSS.n2681 0.029
R16640 DVSS.n3273 DVSS.n3272 0.029
R16641 DVSS.n1832 DVSS.n1831 0.0285734
R16642 DVSS.n3014 DVSS.n3013 0.0285
R16643 DVSS.n3506 DVSS.n3116 0.0285
R16644 DVSS.n3008 DVSS.n2708 0.0285
R16645 DVSS.n3294 DVSS.n3118 0.0285
R16646 DVSS.n800 DVSS.n799 0.0283304
R16647 DVSS.n799 DVSS.n755 0.0283304
R16648 DVSS.n795 DVSS.n755 0.0283304
R16649 DVSS.n795 DVSS.n794 0.0283304
R16650 DVSS.n794 DVSS.n793 0.0283304
R16651 DVSS.n793 DVSS.n757 0.0283304
R16652 DVSS.n789 DVSS.n757 0.0283304
R16653 DVSS.n789 DVSS.n788 0.0283304
R16654 DVSS.n788 DVSS.n787 0.0283304
R16655 DVSS.n787 DVSS.n759 0.0283304
R16656 DVSS.n783 DVSS.n759 0.0283304
R16657 DVSS.n783 DVSS.n782 0.0283304
R16658 DVSS.n782 DVSS.n781 0.0283304
R16659 DVSS.n781 DVSS.n761 0.0283304
R16660 DVSS.n777 DVSS.n761 0.0283304
R16661 DVSS.n777 DVSS.n776 0.0283304
R16662 DVSS.n776 DVSS.n775 0.0283304
R16663 DVSS.n775 DVSS.n763 0.0283304
R16664 DVSS.n771 DVSS.n763 0.0283304
R16665 DVSS.n771 DVSS.n770 0.0283304
R16666 DVSS.n770 DVSS.n769 0.0283304
R16667 DVSS.n769 DVSS.n766 0.0283304
R16668 DVSS.n5730 DVSS.n56 0.0283304
R16669 DVSS.n72 DVSS.n56 0.0283304
R16670 DVSS.n73 DVSS.n72 0.0283304
R16671 DVSS.n73 DVSS.n71 0.0283304
R16672 DVSS.n77 DVSS.n71 0.0283304
R16673 DVSS.n78 DVSS.n77 0.0283304
R16674 DVSS.n79 DVSS.n78 0.0283304
R16675 DVSS.n79 DVSS.n69 0.0283304
R16676 DVSS.n83 DVSS.n69 0.0283304
R16677 DVSS.n84 DVSS.n83 0.0283304
R16678 DVSS.n85 DVSS.n84 0.0283304
R16679 DVSS.n85 DVSS.n67 0.0283304
R16680 DVSS.n89 DVSS.n67 0.0283304
R16681 DVSS.n90 DVSS.n89 0.0283304
R16682 DVSS.n91 DVSS.n90 0.0283304
R16683 DVSS.n91 DVSS.n65 0.0283304
R16684 DVSS.n95 DVSS.n65 0.0283304
R16685 DVSS.n96 DVSS.n95 0.0283304
R16686 DVSS.n97 DVSS.n96 0.0283304
R16687 DVSS.n97 DVSS.n63 0.0283304
R16688 DVSS.n101 DVSS.n63 0.0283304
R16689 DVSS.n5720 DVSS.n5719 0.0283304
R16690 DVSS.n2129 DVSS.n1945 0.0281606
R16691 DVSS.n2105 DVSS.n2104 0.0280676
R16692 DVSS.n2966 DVSS.n2724 0.028
R16693 DVSS.n3481 DVSS.n3152 0.028
R16694 DVSS.n2937 DVSS.n2936 0.028
R16695 DVSS.n3315 DVSS.n3314 0.028
R16696 DVSS.n2794 DVSS.n2788 0.0279877
R16697 DVSS.n2816 DVSS.n2788 0.0279877
R16698 DVSS.n2818 DVSS.n2816 0.0279877
R16699 DVSS.n2818 DVSS.n2817 0.0279877
R16700 DVSS.n2841 DVSS.n2840 0.0279877
R16701 DVSS.n2841 DVSS.n2768 0.0279877
R16702 DVSS.n2859 DVSS.n2768 0.0279877
R16703 DVSS.n2860 DVSS.n2859 0.0279877
R16704 DVSS.n2862 DVSS.n2860 0.0279877
R16705 DVSS.n2889 DVSS.n2759 0.0279877
R16706 DVSS.n2890 DVSS.n2748 0.0279877
R16707 DVSS.n2912 DVSS.n2748 0.0279877
R16708 DVSS.n2913 DVSS.n2912 0.0279877
R16709 DVSS.n2917 DVSS.n2916 0.0279877
R16710 DVSS.n2917 DVSS.n2737 0.0279877
R16711 DVSS.n2951 DVSS.n2737 0.0279877
R16712 DVSS.n2953 DVSS.n2951 0.0279877
R16713 DVSS.n2953 DVSS.n2952 0.0279877
R16714 DVSS.n2968 DVSS.n2967 0.0279877
R16715 DVSS.n2972 DVSS.n2971 0.0279877
R16716 DVSS.n2972 DVSS.n2713 0.0279877
R16717 DVSS.n2990 DVSS.n2713 0.0279877
R16718 DVSS.n2992 DVSS.n2704 0.0279877
R16719 DVSS.n3015 DVSS.n2704 0.0279877
R16720 DVSS.n3016 DVSS.n3015 0.0279877
R16721 DVSS.n3018 DVSS.n3016 0.0279877
R16722 DVSS.n3018 DVSS.n3017 0.0279877
R16723 DVSS.n3038 DVSS.n3037 0.0279877
R16724 DVSS.n3056 DVSS.n2683 0.0279877
R16725 DVSS.n3057 DVSS.n3056 0.0279877
R16726 DVSS.n3059 DVSS.n3057 0.0279877
R16727 DVSS.n3547 DVSS.n2670 0.0279877
R16728 DVSS.n3547 DVSS.n3546 0.0279877
R16729 DVSS.n3546 DVSS.n2671 0.0279877
R16730 DVSS.n3077 DVSS.n2671 0.0279877
R16731 DVSS.n3535 DVSS.n3077 0.0279877
R16732 DVSS.n3097 DVSS.n3096 0.0279877
R16733 DVSS.n3522 DVSS.n3097 0.0279877
R16734 DVSS.n3522 DVSS.n3521 0.0279877
R16735 DVSS.n3521 DVSS.n3098 0.0279877
R16736 DVSS.n3510 DVSS.n3114 0.0279877
R16737 DVSS.n3510 DVSS.n3509 0.0279877
R16738 DVSS.n3509 DVSS.n3115 0.0279877
R16739 DVSS.n3131 DVSS.n3115 0.0279877
R16740 DVSS.n3132 DVSS.n3131 0.0279877
R16741 DVSS.n3496 DVSS.n3134 0.0279877
R16742 DVSS.n3150 DVSS.n3134 0.0279877
R16743 DVSS.n3485 DVSS.n3150 0.0279877
R16744 DVSS.n3485 DVSS.n3484 0.0279877
R16745 DVSS.n3482 DVSS.n3151 0.0279877
R16746 DVSS.n3168 DVSS.n3151 0.0279877
R16747 DVSS.n3471 DVSS.n3168 0.0279877
R16748 DVSS.n3471 DVSS.n3470 0.0279877
R16749 DVSS.n3470 DVSS.n3169 0.0279877
R16750 DVSS.n3459 DVSS.n3188 0.0279877
R16751 DVSS.n3459 DVSS.n3458 0.0279877
R16752 DVSS.n3458 DVSS.n3189 0.0279877
R16753 DVSS.n3205 DVSS.n3189 0.0279877
R16754 DVSS.n3447 DVSS.n3446 0.0279877
R16755 DVSS.n3446 DVSS.n3207 0.0279877
R16756 DVSS.n3223 DVSS.n3207 0.0279877
R16757 DVSS.n3224 DVSS.n3223 0.0279877
R16758 DVSS.n3435 DVSS.n3224 0.0279877
R16759 DVSS.n3241 DVSS.n3240 0.0279877
R16760 DVSS.n3422 DVSS.n3241 0.0279877
R16761 DVSS.n3422 DVSS.n3421 0.0279877
R16762 DVSS.n3421 DVSS.n3420 0.0279877
R16763 DVSS.n2801 DVSS.n2800 0.0279877
R16764 DVSS.n2800 DVSS.n2784 0.0279877
R16765 DVSS.n2824 DVSS.n2784 0.0279877
R16766 DVSS.n2825 DVSS.n2824 0.0279877
R16767 DVSS.n2833 DVSS.n2832 0.0279877
R16768 DVSS.n2832 DVSS.n2830 0.0279877
R16769 DVSS.n2830 DVSS.n2828 0.0279877
R16770 DVSS.n2828 DVSS.n2764 0.0279877
R16771 DVSS.n2868 DVSS.n2764 0.0279877
R16772 DVSS.n2882 DVSS.n2870 0.0279877
R16773 DVSS.n2881 DVSS.n2879 0.0279877
R16774 DVSS.n2879 DVSS.n2877 0.0279877
R16775 DVSS.n2877 DVSS.n2872 0.0279877
R16776 DVSS.n2923 DVSS.n2742 0.0279877
R16777 DVSS.n2924 DVSS.n2923 0.0279877
R16778 DVSS.n2944 DVSS.n2924 0.0279877
R16779 DVSS.n2944 DVSS.n2943 0.0279877
R16780 DVSS.n2943 DVSS.n2941 0.0279877
R16781 DVSS.n2938 DVSS.n2925 0.0279877
R16782 DVSS.n2933 DVSS.n2932 0.0279877
R16783 DVSS.n2932 DVSS.n2930 0.0279877
R16784 DVSS.n2930 DVSS.n2928 0.0279877
R16785 DVSS.n2999 DVSS.n2998 0.0279877
R16786 DVSS.n3007 DVSS.n2999 0.0279877
R16787 DVSS.n3007 DVSS.n3006 0.0279877
R16788 DVSS.n3006 DVSS.n3003 0.0279877
R16789 DVSS.n3003 DVSS.n3002 0.0279877
R16790 DVSS.n3044 DVSS.n2688 0.0279877
R16791 DVSS.n3048 DVSS.n3045 0.0279877
R16792 DVSS.n3048 DVSS.n3047 0.0279877
R16793 DVSS.n3047 DVSS.n2662 0.0279877
R16794 DVSS.n3553 DVSS.n2663 0.0279877
R16795 DVSS.n3257 DVSS.n2663 0.0279877
R16796 DVSS.n3258 DVSS.n3257 0.0279877
R16797 DVSS.n3262 DVSS.n3258 0.0279877
R16798 DVSS.n3263 DVSS.n3262 0.0279877
R16799 DVSS.n3269 DVSS.n3268 0.0279877
R16800 DVSS.n3274 DVSS.n3252 0.0279877
R16801 DVSS.n3275 DVSS.n3274 0.0279877
R16802 DVSS.n3280 DVSS.n3275 0.0279877
R16803 DVSS.n3281 DVSS.n3280 0.0279877
R16804 DVSS.n3286 DVSS.n3285 0.0279877
R16805 DVSS.n3286 DVSS.n3249 0.0279877
R16806 DVSS.n3292 DVSS.n3249 0.0279877
R16807 DVSS.n3293 DVSS.n3292 0.0279877
R16808 DVSS.n3297 DVSS.n3293 0.0279877
R16809 DVSS.n3305 DVSS.n3304 0.0279877
R16810 DVSS.n3309 DVSS.n3305 0.0279877
R16811 DVSS.n3310 DVSS.n3309 0.0279877
R16812 DVSS.n3311 DVSS.n3310 0.0279877
R16813 DVSS.n3317 DVSS.n3316 0.0279877
R16814 DVSS.n3321 DVSS.n3317 0.0279877
R16815 DVSS.n3322 DVSS.n3321 0.0279877
R16816 DVSS.n3327 DVSS.n3322 0.0279877
R16817 DVSS.n3329 DVSS.n3327 0.0279877
R16818 DVSS.n3335 DVSS.n3334 0.0279877
R16819 DVSS.n3340 DVSS.n3335 0.0279877
R16820 DVSS.n3341 DVSS.n3340 0.0279877
R16821 DVSS.n3345 DVSS.n3341 0.0279877
R16822 DVSS.n3352 DVSS.n3347 0.0279877
R16823 DVSS.n3353 DVSS.n3352 0.0279877
R16824 DVSS.n3354 DVSS.n3353 0.0279877
R16825 DVSS.n3358 DVSS.n3354 0.0279877
R16826 DVSS.n3359 DVSS.n3358 0.0279877
R16827 DVSS.n3369 DVSS.n3365 0.0279877
R16828 DVSS.n3370 DVSS.n3369 0.0279877
R16829 DVSS.n3371 DVSS.n3370 0.0279877
R16830 DVSS.n3371 DVSS.n1704 0.0279877
R16831 DVSS.n3250 DVSS.n3114 0.0275443
R16832 DVSS.n3285 DVSS.n3251 0.0275443
R16833 DVSS.n2819 DVSS.n2787 0.0275
R16834 DVSS.n2911 DVSS.n2747 0.0275
R16835 DVSS.n3461 DVSS.n3460 0.0275
R16836 DVSS.n3424 DVSS.n3238 0.0275
R16837 DVSS.n2823 DVSS.n2785 0.0275
R16838 DVSS.n2876 DVSS.n2875 0.0275
R16839 DVSS.n3336 DVSS.n3180 0.0275
R16840 DVSS.n3368 DVSS.n3235 0.0275
R16841 DVSS.n2150 DVSS.n2149 0.0274684
R16842 DVSS.n2147 DVSS.n2146 0.0274684
R16843 DVSS.n1878 DVSS.n1869 0.0274684
R16844 DVSS.n1875 DVSS.n1788 0.0274684
R16845 DVSS.n5720 DVSS.n61 0.0272082
R16846 DVSS.n3535 DVSS.n3534 0.027101
R16847 DVSS.n3263 DVSS.n3253 0.027101
R16848 DVSS.n2857 DVSS.n2769 0.027
R16849 DVSS.n2864 DVSS.n2760 0.027
R16850 DVSS.n3448 DVSS.n3204 0.027
R16851 DVSS.n3221 DVSS.n3220 0.027
R16852 DVSS.n2829 DVSS.n2771 0.027
R16853 DVSS.n2866 DVSS.n2762 0.027
R16854 DVSS.n3350 DVSS.n3348 0.027
R16855 DVSS.n3357 DVSS.n3356 0.027
R16856 DVSS.n1852 DVSS.n1849 0.026913
R16857 DVSS.n1849 DVSS.n1848 0.026913
R16858 DVSS.n1848 DVSS.n1846 0.026913
R16859 DVSS.n1846 DVSS.n1844 0.026913
R16860 DVSS.n1844 DVSS.n1842 0.026913
R16861 DVSS.n1842 DVSS.n1839 0.026913
R16862 DVSS.n1839 DVSS.n1838 0.026913
R16863 DVSS.n1838 DVSS.n1836 0.026913
R16864 DVSS.n1836 DVSS.n1390 0.026913
R16865 DVSS.n4002 DVSS.n1437 0.026913
R16866 DVSS.n4002 DVSS.n4001 0.026913
R16867 DVSS.n4001 DVSS.n3999 0.026913
R16868 DVSS.n3999 DVSS.n3996 0.026913
R16869 DVSS.n3996 DVSS.n3995 0.026913
R16870 DVSS.n3995 DVSS.n3993 0.026913
R16871 DVSS.n3993 DVSS.n3991 0.026913
R16872 DVSS.n3991 DVSS.n3988 0.026913
R16873 DVSS.n1859 DVSS.n1435 0.026913
R16874 DVSS.n3998 DVSS.n3997 0.026913
R16875 DVSS.n3990 DVSS.n3989 0.026913
R16876 DVSS.n4181 DVSS.n1370 0.0267204
R16877 DVSS.n2226 DVSS.n1734 0.0267108
R16878 DVSS.n1937 DVSS.n1933 0.0265092
R16879 DVSS.n2187 DVSS.n1772 0.0265092
R16880 DVSS.n2919 DVSS.n2738 0.0265
R16881 DVSS.n3469 DVSS.n3468 0.0265
R16882 DVSS.n2921 DVSS.n2740 0.0265
R16883 DVSS.n3326 DVSS.n3172 0.0265
R16884 DVSS.n3533 DVSS.n3078 0.0262143
R16885 DVSS.n3497 DVSS.n3133 0.0262143
R16886 DVSS.n3299 DVSS.n3298 0.0262143
R16887 DVSS.n2420 DVSS.n2277 0.02615
R16888 DVSS.n2974 DVSS.n2714 0.026
R16889 DVSS.n3147 DVSS.n3135 0.026
R16890 DVSS.n2929 DVSS.n2722 0.026
R16891 DVSS.n3307 DVSS.n3306 0.026
R16892 DVSS.n1597 DVSS.n1596 0.0258812
R16893 DVSS.n3059 DVSS.n3058 0.0257709
R16894 DVSS.n462 DVSS.n230 0.0257489
R16895 DVSS.n458 DVSS.n230 0.0257489
R16896 DVSS.n458 DVSS.n457 0.0257489
R16897 DVSS.n457 DVSS.n456 0.0257489
R16898 DVSS.n456 DVSS.n232 0.0257489
R16899 DVSS.n452 DVSS.n232 0.0257489
R16900 DVSS.n452 DVSS.n451 0.0257489
R16901 DVSS.n451 DVSS.n450 0.0257489
R16902 DVSS.n450 DVSS.n234 0.0257489
R16903 DVSS.n446 DVSS.n234 0.0257489
R16904 DVSS.n446 DVSS.n445 0.0257489
R16905 DVSS.n445 DVSS.n444 0.0257489
R16906 DVSS.n444 DVSS.n236 0.0257489
R16907 DVSS.n440 DVSS.n236 0.0257489
R16908 DVSS.n440 DVSS.n439 0.0257489
R16909 DVSS.n439 DVSS.n438 0.0257489
R16910 DVSS.n438 DVSS.n238 0.0257489
R16911 DVSS.n434 DVSS.n238 0.0257489
R16912 DVSS.n434 DVSS.n433 0.0257489
R16913 DVSS.n433 DVSS.n432 0.0257489
R16914 DVSS.n432 DVSS.n240 0.0257489
R16915 DVSS.n428 DVSS.n240 0.0257489
R16916 DVSS.n272 DVSS.n271 0.0257489
R16917 DVSS.n278 DVSS.n271 0.0257489
R16918 DVSS.n279 DVSS.n278 0.0257489
R16919 DVSS.n280 DVSS.n279 0.0257489
R16920 DVSS.n280 DVSS.n269 0.0257489
R16921 DVSS.n284 DVSS.n269 0.0257489
R16922 DVSS.n285 DVSS.n284 0.0257489
R16923 DVSS.n286 DVSS.n285 0.0257489
R16924 DVSS.n286 DVSS.n267 0.0257489
R16925 DVSS.n290 DVSS.n267 0.0257489
R16926 DVSS.n291 DVSS.n290 0.0257489
R16927 DVSS.n292 DVSS.n291 0.0257489
R16928 DVSS.n292 DVSS.n265 0.0257489
R16929 DVSS.n296 DVSS.n265 0.0257489
R16930 DVSS.n297 DVSS.n296 0.0257489
R16931 DVSS.n298 DVSS.n297 0.0257489
R16932 DVSS.n298 DVSS.n263 0.0257489
R16933 DVSS.n302 DVSS.n263 0.0257489
R16934 DVSS.n303 DVSS.n302 0.0257489
R16935 DVSS.n304 DVSS.n303 0.0257489
R16936 DVSS.n304 DVSS.n259 0.0257489
R16937 DVSS.n309 DVSS.n261 0.0257489
R16938 DVSS.n2094 DVSS.n2090 0.0256835
R16939 DVSS.n2890 DVSS 0.0255493
R16940 DVSS DVSS.n2881 0.0255493
R16941 DVSS.n3036 DVSS.n3035 0.0255
R16942 DVSS.n3512 DVSS.n3112 0.0255
R16943 DVSS.n2696 DVSS.n2695 0.0255
R16944 DVSS.n3284 DVSS.n3109 0.0255
R16945 DVSS.n3545 DVSS.n2669 0.025
R16946 DVSS.n3536 DVSS.n3076 0.025
R16947 DVSS.n3256 DVSS.n3255 0.025
R16948 DVSS.n3266 DVSS.n3264 0.025
R16949 DVSS.n5719 DVSS.n5718 0.0249638
R16950 DVSS.n3483 DVSS.n3482 0.0248842
R16951 DVSS.n3316 DVSS.n3247 0.0248842
R16952 DVSS.n4547 DVSS.n4546 0.0248508
R16953 DVSS.n2804 DVSS.n2793 0.0248045
R16954 DVSS.n261 DVSS.n260 0.0247308
R16955 DVSS.n3055 DVSS.n3054 0.0245
R16956 DVSS.n3524 DVSS.n3523 0.0245
R16957 DVSS.n3049 DVSS.n2687 0.0245
R16958 DVSS.n3276 DVSS.n3089 0.0245
R16959 DVSS.n3017 DVSS.n2692 0.0244409
R16960 DVSS.n3002 DVSS.n3000 0.0244409
R16961 DVSS DVSS.n2242 0.0241842
R16962 DVSS.n3012 DVSS.n2705 0.024
R16963 DVSS.n3129 DVSS.n3128 0.024
R16964 DVSS.n3009 DVSS.n2707 0.024
R16965 DVSS.n3296 DVSS.n3295 0.024
R16966 DVSS.n3187 DVSS.n3184 0.0235542
R16967 DVSS.n3331 DVSS.n3330 0.0235542
R16968 DVSS.n2965 DVSS.n2726 0.0235
R16969 DVSS.n3480 DVSS.n3153 0.0235
R16970 DVSS.n2940 DVSS.n2728 0.0235
R16971 DVSS.n3318 DVSS.n3155 0.0235
R16972 DVSS.n2991 DVSS.n2990 0.0231108
R16973 DVSS.n2928 DVSS.n2709 0.0231108
R16974 DVSS.n2820 DVSS.n2780 0.023
R16975 DVSS.n2910 DVSS.n2749 0.023
R16976 DVSS.n3457 DVSS.n3183 0.023
R16977 DVSS.n3237 DVSS.n3225 0.023
R16978 DVSS.n2822 DVSS.n2782 0.023
R16979 DVSS.n2878 DVSS.n2751 0.023
R16980 DVSS.n3339 DVSS.n3338 0.023
R16981 DVSS.n3367 DVSS.n3366 0.023
R16982 DVSS.n2971 DVSS 0.0228892
R16983 DVSS.n2933 DVSS 0.0228892
R16984 DVSS.n1825 DVSS.n1746 0.0227936
R16985 DVSS.n2204 DVSS.n2203 0.0227859
R16986 DVSS.n1774 DVSS.n1757 0.0227859
R16987 DVSS.n1785 DVSS.n1783 0.0227859
R16988 DVSS.n2165 DVSS.n1800 0.0227859
R16989 DVSS.n1949 DVSS.n1948 0.0227859
R16990 DVSS.n1786 DVSS.n1785 0.0227859
R16991 DVSS.n1802 DVSS.n1800 0.0227859
R16992 DVSS.n1946 DVSS.n1941 0.0227859
R16993 DVSS.n1755 DVSS.n1751 0.0227859
R16994 DVSS.n2207 DVSS.n2206 0.0227859
R16995 DVSS.n4000 DVSS.n1432 0.0227554
R16996 DVSS.n3994 DVSS.n1429 0.0227554
R16997 DVSS.n310 DVSS.n309 0.0226946
R16998 DVSS.n250 DVSS.n249 0.0226275
R16999 DVSS.n2843 DVSS.n2842 0.0225
R17000 DVSS.n2888 DVSS.n2887 0.0225
R17001 DVSS.n3449 DVSS.n3203 0.0225
R17002 DVSS.n3437 DVSS.n3436 0.0225
R17003 DVSS.n2831 DVSS.n2777 0.0225
R17004 DVSS.n2884 DVSS.n2883 0.0225
R17005 DVSS.n3344 DVSS.n3200 0.0225
R17006 DVSS.n3360 DVSS.n3218 0.0225
R17007 DVSS.n2114 DVSS.n2098 0.0223919
R17008 DVSS.n2112 DVSS.n2098 0.0223919
R17009 DVSS.n1821 DVSS.n1748 0.0223919
R17010 DVSS.n2111 DVSS.n2089 0.0223919
R17011 DVSS.n2113 DVSS.n2111 0.0223919
R17012 DVSS.n1826 DVSS.n1825 0.0223807
R17013 DVSS.n1825 DVSS.n1824 0.0223807
R17014 DVSS.n3447 DVSS.n3206 0.0222241
R17015 DVSS.n3347 DVSS.n3346 0.0222241
R17016 DVSS.n2950 DVSS.n2949 0.022
R17017 DVSS.n3472 DVSS.n3167 0.022
R17018 DVSS.n2946 DVSS.n2945 0.022
R17019 DVSS.n3325 DVSS.n3323 0.022
R17020 DVSS.n2952 DVSS.n2725 0.0217808
R17021 DVSS.n2941 DVSS.n2939 0.0217808
R17022 DVSS.n4965 DVSS.n1162 0.0216765
R17023 DVSS.n4451 DVSS.n4448 0.0216765
R17024 DVSS.n4960 DVSS.n4957 0.0216765
R17025 DVSS.n2167 DVSS.n1801 0.021555
R17026 DVSS.n2201 DVSS.n1752 0.021555
R17027 DVSS.n5722 DVSS.n5721 0.0215113
R17028 DVSS.n2989 DVSS.n2988 0.0215
R17029 DVSS.n3495 DVSS.n3494 0.0215
R17030 DVSS.n2927 DVSS.n2716 0.0215
R17031 DVSS.n3303 DVSS.n3137 0.0215
R17032 DVSS.n4094 DVSS.n4003 0.021288
R17033 DVSS.n3992 DVSS.n1428 0.021288
R17034 DVSS.n5116 DVSS.n5115 0.021205
R17035 DVSS.n5117 DVSS.n5116 0.021205
R17036 DVSS.n5117 DVSS.n1077 0.021205
R17037 DVSS.n5123 DVSS.n1077 0.021205
R17038 DVSS.n5124 DVSS.n5123 0.021205
R17039 DVSS.n5125 DVSS.n5124 0.021205
R17040 DVSS.n5125 DVSS.n1073 0.021205
R17041 DVSS.n5131 DVSS.n1073 0.021205
R17042 DVSS.n5132 DVSS.n5131 0.021205
R17043 DVSS.n5133 DVSS.n5132 0.021205
R17044 DVSS.n5133 DVSS.n1069 0.021205
R17045 DVSS.n5139 DVSS.n1069 0.021205
R17046 DVSS.n5140 DVSS.n5139 0.021205
R17047 DVSS.n5141 DVSS.n5140 0.021205
R17048 DVSS.n5141 DVSS.n1065 0.021205
R17049 DVSS.n5147 DVSS.n1065 0.021205
R17050 DVSS.n5148 DVSS.n5147 0.021205
R17051 DVSS.n5149 DVSS.n5148 0.021205
R17052 DVSS.n5149 DVSS.n1061 0.021205
R17053 DVSS.n5155 DVSS.n1061 0.021205
R17054 DVSS.n5156 DVSS.n5155 0.021205
R17055 DVSS.n5157 DVSS.n5156 0.021205
R17056 DVSS.n5157 DVSS.n1057 0.021205
R17057 DVSS.n5163 DVSS.n1057 0.021205
R17058 DVSS.n5164 DVSS.n5163 0.021205
R17059 DVSS.n5165 DVSS.n5164 0.021205
R17060 DVSS.n5165 DVSS.n1053 0.021205
R17061 DVSS.n5171 DVSS.n1053 0.021205
R17062 DVSS.n5172 DVSS.n5171 0.021205
R17063 DVSS.n5173 DVSS.n5172 0.021205
R17064 DVSS.n5173 DVSS.n1049 0.021205
R17065 DVSS.n5179 DVSS.n1049 0.021205
R17066 DVSS.n5180 DVSS.n5179 0.021205
R17067 DVSS.n5181 DVSS.n5180 0.021205
R17068 DVSS.n5181 DVSS.n1045 0.021205
R17069 DVSS.n5187 DVSS.n1045 0.021205
R17070 DVSS.n5188 DVSS.n5187 0.021205
R17071 DVSS.n5189 DVSS.n5188 0.021205
R17072 DVSS.n5189 DVSS.n1041 0.021205
R17073 DVSS.n5195 DVSS.n1041 0.021205
R17074 DVSS.n5196 DVSS.n5195 0.021205
R17075 DVSS.n5197 DVSS.n5196 0.021205
R17076 DVSS.n5197 DVSS.n1037 0.021205
R17077 DVSS.n5203 DVSS.n1037 0.021205
R17078 DVSS.n5204 DVSS.n5203 0.021205
R17079 DVSS.n5205 DVSS.n5204 0.021205
R17080 DVSS.n5205 DVSS.n1033 0.021205
R17081 DVSS.n5211 DVSS.n1033 0.021205
R17082 DVSS.n5212 DVSS.n5211 0.021205
R17083 DVSS.n5213 DVSS.n5212 0.021205
R17084 DVSS.n5213 DVSS.n1029 0.021205
R17085 DVSS.n5219 DVSS.n1029 0.021205
R17086 DVSS.n5220 DVSS.n5219 0.021205
R17087 DVSS.n5222 DVSS.n5220 0.021205
R17088 DVSS.n5222 DVSS.n5221 0.021205
R17089 DVSS.n5221 DVSS.n1025 0.021205
R17090 DVSS.n5229 DVSS.n1025 0.021205
R17091 DVSS.n5236 DVSS.n1020 0.021205
R17092 DVSS.n5237 DVSS.n5236 0.021205
R17093 DVSS.n5238 DVSS.n5237 0.021205
R17094 DVSS.n5238 DVSS.n1016 0.021205
R17095 DVSS.n5244 DVSS.n1016 0.021205
R17096 DVSS.n5245 DVSS.n5244 0.021205
R17097 DVSS.n5246 DVSS.n5245 0.021205
R17098 DVSS.n5246 DVSS.n1012 0.021205
R17099 DVSS.n5252 DVSS.n1012 0.021205
R17100 DVSS.n5253 DVSS.n5252 0.021205
R17101 DVSS.n5254 DVSS.n5253 0.021205
R17102 DVSS.n5254 DVSS.n1008 0.021205
R17103 DVSS.n5260 DVSS.n1008 0.021205
R17104 DVSS.n5261 DVSS.n5260 0.021205
R17105 DVSS.n5262 DVSS.n5261 0.021205
R17106 DVSS.n5262 DVSS.n1004 0.021205
R17107 DVSS.n5268 DVSS.n1004 0.021205
R17108 DVSS.n5269 DVSS.n5268 0.021205
R17109 DVSS.n5270 DVSS.n5269 0.021205
R17110 DVSS.n5270 DVSS.n1000 0.021205
R17111 DVSS.n5276 DVSS.n1000 0.021205
R17112 DVSS.n5277 DVSS.n5276 0.021205
R17113 DVSS.n5278 DVSS.n5277 0.021205
R17114 DVSS.n5278 DVSS.n996 0.021205
R17115 DVSS.n5284 DVSS.n996 0.021205
R17116 DVSS.n5285 DVSS.n5284 0.021205
R17117 DVSS.n5286 DVSS.n5285 0.021205
R17118 DVSS.n5286 DVSS.n992 0.021205
R17119 DVSS.n5292 DVSS.n992 0.021205
R17120 DVSS.n5293 DVSS.n5292 0.021205
R17121 DVSS.n5294 DVSS.n5293 0.021205
R17122 DVSS.n5294 DVSS.n988 0.021205
R17123 DVSS.n5300 DVSS.n988 0.021205
R17124 DVSS.n5301 DVSS.n5300 0.021205
R17125 DVSS.n5302 DVSS.n5301 0.021205
R17126 DVSS.n5302 DVSS.n984 0.021205
R17127 DVSS.n5308 DVSS.n984 0.021205
R17128 DVSS.n5309 DVSS.n5308 0.021205
R17129 DVSS.n5310 DVSS.n5309 0.021205
R17130 DVSS.n5310 DVSS.n980 0.021205
R17131 DVSS.n5316 DVSS.n980 0.021205
R17132 DVSS.n5317 DVSS.n5316 0.021205
R17133 DVSS.n5318 DVSS.n5317 0.021205
R17134 DVSS.n5318 DVSS.n976 0.021205
R17135 DVSS.n5324 DVSS.n976 0.021205
R17136 DVSS.n5325 DVSS.n5324 0.021205
R17137 DVSS.n5326 DVSS.n5325 0.021205
R17138 DVSS.n5326 DVSS.n972 0.021205
R17139 DVSS.n5332 DVSS.n972 0.021205
R17140 DVSS.n5333 DVSS.n5332 0.021205
R17141 DVSS.n5334 DVSS.n5333 0.021205
R17142 DVSS.n5334 DVSS.n968 0.021205
R17143 DVSS.n5340 DVSS.n968 0.021205
R17144 DVSS.n5341 DVSS.n5340 0.021205
R17145 DVSS.n5343 DVSS.n5341 0.021205
R17146 DVSS.n5343 DVSS.n5342 0.021205
R17147 DVSS.n5342 DVSS.n964 0.021205
R17148 DVSS.n5350 DVSS.n964 0.021205
R17149 DVSS.n2111 DVSS.n2110 0.0211757
R17150 DVSS.n1821 DVSS.n1820 0.0211757
R17151 DVSS.n2183 DVSS.n2182 0.0211422
R17152 DVSS.n3039 DVSS.n2691 0.021
R17153 DVSS.n3111 DVSS.n3099 0.021
R17154 DVSS.n3043 DVSS.n2689 0.021
R17155 DVSS.n3283 DVSS.n3282 0.021
R17156 DVSS.n3434 DVSS.n3433 0.0208941
R17157 DVSS.n3364 DVSS.n3245 0.0208941
R17158 DVSS.n2168 DVSS.n2167 0.02075
R17159 DVSS.n2167 DVSS.n2166 0.02075
R17160 DVSS.n2182 DVSS.n1784 0.02075
R17161 DVSS.n2182 DVSS.n2181 0.02075
R17162 DVSS.n3555 DVSS.n2662 0.0206724
R17163 DVSS.n307 DVSS.n60 0.0206158
R17164 DVSS.n3544 DVSS.n2672 0.0205
R17165 DVSS.n3537 DVSS.n3075 0.0205
R17166 DVSS.n3259 DVSS.n2674 0.0205
R17167 DVSS.n3261 DVSS.n3072 0.0205
R17168 DVSS.n2913 DVSS.n2746 0.0204507
R17169 DVSS.n2872 DVSS.n2871 0.0204507
R17170 DVSS DVSS.n2683 0.0202291
R17171 DVSS.n3045 DVSS 0.0202291
R17172 DVSS.n5727 DVSS.n5726 0.020197
R17173 DVSS.n3053 DVSS.n2684 0.02
R17174 DVSS.n3520 DVSS.n3092 0.02
R17175 DVSS.n3050 DVSS.n2686 0.02
R17176 DVSS.n3279 DVSS.n3278 0.02
R17177 DVSS.n2097 DVSS.n2090 0.0199037
R17178 DVSS.n2209 DVSS.n1747 0.0199037
R17179 DVSS.n854 DVSS.n852 0.0195912
R17180 DVSS.n854 DVSS.n851 0.0195912
R17181 DVSS.n1191 DVSS.n851 0.0195912
R17182 DVSS.n853 DVSS.n850 0.0195912
R17183 DVSS.n853 DVSS.n849 0.0195912
R17184 DVSS.n849 DVSS.n848 0.0195912
R17185 DVSS.n2994 DVSS.n2993 0.0195
R17186 DVSS.n3499 DVSS.n3498 0.0195
R17187 DVSS.n2997 DVSS.n2996 0.0195
R17188 DVSS.n3300 DVSS.n3126 0.0195
R17189 DVSS.n766 DVSS.n765 0.0191284
R17190 DVSS.n2862 DVSS.n2861 0.0191207
R17191 DVSS.n2869 DVSS.n2868 0.0191207
R17192 DVSS.n1938 DVSS.n1937 0.019078
R17193 DVSS.n2187 DVSS.n2186 0.019078
R17194 DVSS.n2955 DVSS.n2954 0.019
R17195 DVSS.n3166 DVSS.n3165 0.019
R17196 DVSS.n2942 DVSS.n2735 0.019
R17197 DVSS.n3320 DVSS.n3319 0.019
R17198 DVSS.n3433 DVSS 0.018899
R17199 DVSS DVSS.n3364 0.018899
R17200 DVSS.n2839 DVSS.n2838 0.0185
R17201 DVSS.n2892 DVSS.n2891 0.0185
R17202 DVSS.n3456 DVSS.n3190 0.0185
R17203 DVSS.n3432 DVSS.n3431 0.0185
R17204 DVSS.n2835 DVSS.n2834 0.0185
R17205 DVSS.n2880 DVSS.n2757 0.0185
R17206 DVSS.n3342 DVSS.n3192 0.0185
R17207 DVSS.n3363 DVSS.n3227 0.0185
R17208 DVSS.n5551 DVSS.n856 0.018166
R17209 DVSS.n2839 DVSS.n2778 0.018
R17210 DVSS.n2891 DVSS.n2758 0.018
R17211 DVSS.n3202 DVSS.n3190 0.018
R17212 DVSS.n3432 DVSS.n3222 0.018
R17213 DVSS.n2834 DVSS.n2783 0.018
R17214 DVSS.n2880 DVSS.n2763 0.018
R17215 DVSS.n3343 DVSS.n3342 0.018
R17216 DVSS.n3363 DVSS.n3362 0.018
R17217 DVSS.n1752 DVSS.n1747 0.0178394
R17218 DVSS.n2817 DVSS.n2779 0.0177906
R17219 DVSS.n2826 DVSS.n2825 0.0177906
R17220 DVSS.n4822 DVSS.n4821 0.0176
R17221 DVSS.n4538 DVSS.n4527 0.0176
R17222 DVSS.n3096 DVSS 0.017569
R17223 DVSS DVSS.n3252 0.017569
R17224 DVSS.n2954 DVSS.n2736 0.0175
R17225 DVSS.n3473 DVSS.n3166 0.0175
R17226 DVSS.n2942 DVSS.n2741 0.0175
R17227 DVSS.n3320 DVSS.n3163 0.0175
R17228 DVSS.n2126 DVSS.n1945 0.0174266
R17229 DVSS.n428 DVSS.n427 0.0174005
R17230 DVSS.n4537 DVSS.n4529 0.0172066
R17231 DVSS.n2657 DVSS.n2656 0.0171667
R17232 DVSS.n2658 DVSS.n2657 0.0171667
R17233 DVSS.n5231 DVSS.n5230 0.0171667
R17234 DVSS.n5232 DVSS.n5231 0.0171667
R17235 DVSS.n1831 DVSS.n1830 0.0170138
R17236 DVSS.n2993 DVSS.n2712 0.017
R17237 DVSS.n3498 DVSS.n3130 0.017
R17238 DVSS.n2997 DVSS.n2710 0.017
R17239 DVSS.n3302 DVSS.n3300 0.017
R17240 DVSS.n4829 DVSS.n4806 0.0169185
R17241 DVSS.n4834 DVSS.n4806 0.0169185
R17242 DVSS.n4828 DVSS.n4805 0.0169185
R17243 DVSS.n4833 DVSS.n4805 0.0169185
R17244 DVSS.n4827 DVSS.n4804 0.0169185
R17245 DVSS.n4832 DVSS.n4804 0.0169185
R17246 DVSS.n4826 DVSS.n4803 0.0169185
R17247 DVSS.n4873 DVSS.n4803 0.0169185
R17248 DVSS.n4829 DVSS.n4822 0.0169185
R17249 DVSS.n4834 DVSS.n4823 0.0169185
R17250 DVSS.n4828 DVSS.n4823 0.0169185
R17251 DVSS.n4833 DVSS.n4824 0.0169185
R17252 DVSS.n4827 DVSS.n4824 0.0169185
R17253 DVSS.n4832 DVSS.n4825 0.0169185
R17254 DVSS.n4826 DVSS.n4825 0.0169185
R17255 DVSS.n4874 DVSS.n4873 0.0169185
R17256 DVSS.n4524 DVSS.n4523 0.0169185
R17257 DVSS.n4522 DVSS.n4521 0.0169185
R17258 DVSS.n4520 DVSS.n4519 0.0169185
R17259 DVSS.n4518 DVSS.n4517 0.0169185
R17260 DVSS.n4516 DVSS.n4515 0.0169185
R17261 DVSS.n4514 DVSS.n4513 0.0169185
R17262 DVSS.n4541 DVSS.n4512 0.0169185
R17263 DVSS.n4543 DVSS.n4542 0.0169185
R17264 DVSS.n4527 DVSS.n4524 0.0169185
R17265 DVSS.n4523 DVSS.n4522 0.0169185
R17266 DVSS.n4521 DVSS.n4520 0.0169185
R17267 DVSS.n4519 DVSS.n4518 0.0169185
R17268 DVSS.n4517 DVSS.n4516 0.0169185
R17269 DVSS.n4515 DVSS.n4514 0.0169185
R17270 DVSS.n4513 DVSS.n4512 0.0169185
R17271 DVSS.n4542 DVSS.n4541 0.0169185
R17272 DVSS.n3838 DVSS.n1626 0.0169185
R17273 DVSS.n3837 DVSS.n3835 0.0169185
R17274 DVSS.n3836 DVSS.n1627 0.0169185
R17275 DVSS.n3834 DVSS.n3832 0.0169185
R17276 DVSS.n3833 DVSS.n1628 0.0169185
R17277 DVSS.n3831 DVSS.n3829 0.0169185
R17278 DVSS.n3830 DVSS.n1629 0.0169185
R17279 DVSS.n1631 DVSS.n1630 0.0169185
R17280 DVSS.n1890 DVSS.n1632 0.0169185
R17281 DVSS.n1632 DVSS.n1631 0.0169185
R17282 DVSS.n1630 DVSS.n1629 0.0169185
R17283 DVSS.n3831 DVSS.n3830 0.0169185
R17284 DVSS.n3829 DVSS.n1628 0.0169185
R17285 DVSS.n3834 DVSS.n3833 0.0169185
R17286 DVSS.n3832 DVSS.n1627 0.0169185
R17287 DVSS.n3837 DVSS.n3836 0.0169185
R17288 DVSS.n3835 DVSS.n1626 0.0169185
R17289 DVSS.n3839 DVSS.n3838 0.0169185
R17290 DVSS.n2640 DVSS.n2637 0.0169185
R17291 DVSS.n2637 DVSS.n2270 0.0169185
R17292 DVSS.n2641 DVSS.n2638 0.0169185
R17293 DVSS.n2638 DVSS.n2271 0.0169185
R17294 DVSS.n2642 DVSS.n2639 0.0169185
R17295 DVSS.n2639 DVSS.n2272 0.0169185
R17296 DVSS.n2645 DVSS.n2644 0.0169185
R17297 DVSS.n2645 DVSS.n2273 0.0169185
R17298 DVSS.n2647 DVSS.n2274 0.0169185
R17299 DVSS.n2407 DVSS.n2280 0.0169185
R17300 DVSS.n2406 DVSS.n2404 0.0169185
R17301 DVSS.n2405 DVSS.n2281 0.0169185
R17302 DVSS.n2410 DVSS.n2409 0.0169185
R17303 DVSS.n2411 DVSS.n2410 0.0169185
R17304 DVSS.n2414 DVSS.n2413 0.0169185
R17305 DVSS.n2415 DVSS.n2414 0.0169185
R17306 DVSS.n2418 DVSS.n2417 0.0169185
R17307 DVSS.n2408 DVSS.n2407 0.0169185
R17308 DVSS.n2404 DVSS.n2280 0.0169185
R17309 DVSS.n2406 DVSS.n2405 0.0169185
R17310 DVSS.n2409 DVSS.n2281 0.0169185
R17311 DVSS.n2412 DVSS.n2411 0.0169185
R17312 DVSS.n2413 DVSS.n2412 0.0169185
R17313 DVSS.n2416 DVSS.n2415 0.0169185
R17314 DVSS.n2417 DVSS.n2416 0.0169185
R17315 DVSS.n2640 DVSS.n1699 0.0169185
R17316 DVSS.n2425 DVSS.n2270 0.0169185
R17317 DVSS.n2641 DVSS.n2425 0.0169185
R17318 DVSS.n2424 DVSS.n2271 0.0169185
R17319 DVSS.n2642 DVSS.n2424 0.0169185
R17320 DVSS.n2423 DVSS.n2272 0.0169185
R17321 DVSS.n2644 DVSS.n2423 0.0169185
R17322 DVSS.n2422 DVSS.n2273 0.0169185
R17323 DVSS.n2422 DVSS.n2274 0.0169185
R17324 DVSS.n2106 DVSS.n2105 0.0167162
R17325 DVSS.n5724 DVSS.n5723 0.0166994
R17326 DVSS.n5725 DVSS.n5724 0.0166994
R17327 DVSS.n3040 DVSS.n2684 0.0165
R17328 DVSS.n3520 DVSS.n3519 0.0165
R17329 DVSS.n3042 DVSS.n2686 0.0165
R17330 DVSS.n3279 DVSS.n3101 0.0165
R17331 DVSS.n3420 DVSS.n1703 0.0164606
R17332 DVSS.n3747 DVSS.n1704 0.0164606
R17333 DVSS DVSS.n3187 0.0162389
R17334 DVSS.n3331 DVSS 0.0162389
R17335 DVSS.n3074 DVSS.n2672 0.016
R17336 DVSS.n3075 DVSS.n3074 0.016
R17337 DVSS.n3260 DVSS.n3259 0.016
R17338 DVSS.n3261 DVSS.n3260 0.016
R17339 DVSS.n3040 DVSS.n3039 0.0155
R17340 DVSS.n3519 DVSS.n3099 0.0155
R17341 DVSS.n3043 DVSS.n3042 0.0155
R17342 DVSS.n3282 DVSS.n3101 0.0155
R17343 DVSS.n3398 DVSS.n3397 0.0154891
R17344 DVSS.n4821 DVSS.n4807 0.01535
R17345 DVSS.n4539 DVSS.n4538 0.01535
R17346 DVSS.n1979 DVSS.n1976 0.0152819
R17347 DVSS.n1979 DVSS.n1978 0.0152819
R17348 DVSS.n1974 DVSS.n1812 0.0152819
R17349 DVSS.n1976 DVSS.n1965 0.0152819
R17350 DVSS.n1978 DVSS.n1964 0.0152819
R17351 DVSS.n1974 DVSS.n1964 0.0152819
R17352 DVSS.n1912 DVSS.n1910 0.0152819
R17353 DVSS.n1912 DVSS.n1911 0.0152819
R17354 DVSS.n1914 DVSS.n1881 0.0152819
R17355 DVSS.n1910 DVSS.n1760 0.0152819
R17356 DVSS.n1911 DVSS.n1883 0.0152819
R17357 DVSS.n1883 DVSS.n1881 0.0152819
R17358 DVSS.n276 DVSS.n275 0.0152727
R17359 DVSS.n2989 DVSS.n2712 0.015
R17360 DVSS.n3495 DVSS.n3130 0.015
R17361 DVSS.n2927 DVSS.n2710 0.015
R17362 DVSS.n3303 DVSS.n3302 0.015
R17363 DVSS.n2210 DVSS.n1746 0.0149495
R17364 DVSS DVSS.n3496 0.0149089
R17365 DVSS.n3304 DVSS 0.0149089
R17366 DVSS.n4819 DVSS.n4818 0.0149069
R17367 DVSS.n4813 DVSS.n4812 0.0149069
R17368 DVSS.n4816 DVSS.n4812 0.0149069
R17369 DVSS.n4816 DVSS.n4815 0.0149069
R17370 DVSS.n4818 DVSS.n4810 0.0149069
R17371 DVSS.n4813 DVSS.n4810 0.0149069
R17372 DVSS.n4532 DVSS.n4531 0.0149069
R17373 DVSS.n4534 DVSS.n4530 0.0149069
R17374 DVSS.n4533 DVSS.n4525 0.0149069
R17375 DVSS.n4534 DVSS.n4533 0.0149069
R17376 DVSS.n4532 DVSS.n4530 0.0149069
R17377 DVSS.n4536 DVSS.n4531 0.0149069
R17378 DVSS.n1214 DVSS.n1213 0.0145462
R17379 DVSS.n1213 DVSS.n1210 0.0145462
R17380 DVSS.n1210 DVSS.n1209 0.0145462
R17381 DVSS.n1209 DVSS.n1207 0.0145462
R17382 DVSS.n1207 DVSS.n1205 0.0145462
R17383 DVSS.n1205 DVSS.n1202 0.0145462
R17384 DVSS.n1202 DVSS.n1201 0.0145462
R17385 DVSS.n1201 DVSS.n1199 0.0145462
R17386 DVSS.n1199 DVSS.n1197 0.0145462
R17387 DVSS.n1197 DVSS.n1190 0.0145462
R17388 DVSS.n4930 DVSS.n1190 0.0145462
R17389 DVSS.n1835 DVSS.n1817 0.0145367
R17390 DVSS.n2950 DVSS.n2736 0.0145
R17391 DVSS.n3473 DVSS.n3472 0.0145
R17392 DVSS.n2945 DVSS.n2741 0.0145
R17393 DVSS.n3323 DVSS.n3163 0.0145
R17394 DVSS.n4003 DVSS.n1430 0.0144402
R17395 DVSS.n3992 DVSS.n1433 0.0144402
R17396 DVSS.n954 DVSS.n953 0.0144028
R17397 DVSS.n2023 DVSS.n2022 0.0142903
R17398 DVSS.n2101 DVSS.n1808 0.0142838
R17399 DVSS.n3728 DVSS.n3727 0.0142814
R17400 DVSS.n4037 DVSS.n4036 0.0142814
R17401 DVSS.n1857 DVSS.n1853 0.0141679
R17402 DVSS.n1865 DVSS.n1856 0.0141679
R17403 DVSS.n1856 DVSS.n1853 0.0141679
R17404 DVSS.n1857 DVSS.n1854 0.0141679
R17405 DVSS.n2842 DVSS.n2778 0.014
R17406 DVSS.n2888 DVSS.n2758 0.014
R17407 DVSS.n3203 DVSS.n3202 0.014
R17408 DVSS.n3436 DVSS.n3222 0.014
R17409 DVSS.n2831 DVSS.n2783 0.014
R17410 DVSS.n2883 DVSS.n2763 0.014
R17411 DVSS.n3344 DVSS.n3343 0.014
R17412 DVSS.n3362 DVSS.n3360 0.014
R17413 DVSS.n1212 DVSS.n1211 0.0136707
R17414 DVSS.n1204 DVSS.n1203 0.0136707
R17415 DVSS.n1196 DVSS.n1195 0.0136707
R17416 DVSS.n3497 DVSS 0.0135788
R17417 DVSS.n3299 DVSS 0.0135788
R17418 DVSS.n4815 DVSS.n4807 0.01355
R17419 DVSS.n4539 DVSS.n4525 0.01355
R17420 DVSS.n4191 DVSS.n1367 0.0135392
R17421 DVSS.n2838 DVSS.n2780 0.0135
R17422 DVSS.n2892 DVSS.n2749 0.0135
R17423 DVSS.n3457 DVSS.n3456 0.0135
R17424 DVSS.n3431 DVSS.n3225 0.0135
R17425 DVSS.n2835 DVSS.n2782 0.0135
R17426 DVSS.n2878 DVSS.n2757 0.0135
R17427 DVSS.n3339 DVSS.n3192 0.0135
R17428 DVSS.n3366 DVSS.n3227 0.0135
R17429 DVSS.n1920 DVSS.n1816 0.0134255
R17430 DVSS.n1918 DVSS.n1816 0.0134255
R17431 DVSS.n2157 DVSS.n1807 0.0134255
R17432 DVSS.n2159 DVSS.n1807 0.0134255
R17433 DVSS.n1851 DVSS.n1850 0.0133402
R17434 DVSS.n1841 DVSS.n1840 0.0133402
R17435 DVSS.n2955 DVSS.n2726 0.013
R17436 DVSS.n3165 DVSS.n3153 0.013
R17437 DVSS.n2940 DVSS.n2735 0.013
R17438 DVSS.n3319 DVSS.n3318 0.013
R17439 DVSS.n1847 DVSS.n1386 0.0129835
R17440 DVSS.n1843 DVSS.n1380 0.0129835
R17441 DVSS.n4000 DVSS.n1430 0.0129728
R17442 DVSS.n3994 DVSS.n1433 0.0129728
R17443 DVSS.n798 DVSS.n754 0.0129415
R17444 DVSS.n798 DVSS.n797 0.0129415
R17445 DVSS.n797 DVSS.n796 0.0129415
R17446 DVSS.n796 DVSS.n756 0.0129415
R17447 DVSS.n792 DVSS.n756 0.0129415
R17448 DVSS.n792 DVSS.n791 0.0129415
R17449 DVSS.n791 DVSS.n790 0.0129415
R17450 DVSS.n790 DVSS.n758 0.0129415
R17451 DVSS.n786 DVSS.n758 0.0129415
R17452 DVSS.n786 DVSS.n785 0.0129415
R17453 DVSS.n785 DVSS.n784 0.0129415
R17454 DVSS.n784 DVSS.n760 0.0129415
R17455 DVSS.n780 DVSS.n760 0.0129415
R17456 DVSS.n780 DVSS.n779 0.0129415
R17457 DVSS.n779 DVSS.n778 0.0129415
R17458 DVSS.n778 DVSS.n762 0.0129415
R17459 DVSS.n774 DVSS.n762 0.0129415
R17460 DVSS.n774 DVSS.n773 0.0129415
R17461 DVSS.n773 DVSS.n772 0.0129415
R17462 DVSS.n772 DVSS.n764 0.0129415
R17463 DVSS.n768 DVSS.n764 0.0129415
R17464 DVSS.n768 DVSS.n767 0.0129415
R17465 DVSS.n5729 DVSS.n5728 0.0129415
R17466 DVSS.n74 DVSS.n58 0.0129415
R17467 DVSS.n75 DVSS.n74 0.0129415
R17468 DVSS.n76 DVSS.n75 0.0129415
R17469 DVSS.n76 DVSS.n70 0.0129415
R17470 DVSS.n80 DVSS.n70 0.0129415
R17471 DVSS.n81 DVSS.n80 0.0129415
R17472 DVSS.n82 DVSS.n81 0.0129415
R17473 DVSS.n82 DVSS.n68 0.0129415
R17474 DVSS.n86 DVSS.n68 0.0129415
R17475 DVSS.n87 DVSS.n86 0.0129415
R17476 DVSS.n88 DVSS.n87 0.0129415
R17477 DVSS.n88 DVSS.n66 0.0129415
R17478 DVSS.n92 DVSS.n66 0.0129415
R17479 DVSS.n93 DVSS.n92 0.0129415
R17480 DVSS.n94 DVSS.n93 0.0129415
R17481 DVSS.n94 DVSS.n64 0.0129415
R17482 DVSS.n98 DVSS.n64 0.0129415
R17483 DVSS.n99 DVSS.n98 0.0129415
R17484 DVSS.n100 DVSS.n99 0.0129415
R17485 DVSS.n100 DVSS.n62 0.0129415
R17486 DVSS.n5721 DVSS.n62 0.0129415
R17487 DVSS.n253 DVSS.n248 0.0127612
R17488 DVSS.n254 DVSS.n251 0.0127612
R17489 DVSS.n1752 DVSS.n1749 0.01265
R17490 DVSS.n1752 DVSS.n1750 0.01265
R17491 DVSS.n2994 DVSS.n2705 0.0125
R17492 DVSS.n3499 DVSS.n3129 0.0125
R17493 DVSS.n2996 DVSS.n2707 0.0125
R17494 DVSS.n3296 DVSS.n3126 0.0125
R17495 DVSS.n2136 DVSS.n2135 0.0124725
R17496 DVSS.n1780 DVSS.n1779 0.0124725
R17497 DVSS.n461 DVSS.n460 0.0123471
R17498 DVSS.n460 DVSS.n459 0.0123471
R17499 DVSS.n459 DVSS.n231 0.0123471
R17500 DVSS.n455 DVSS.n231 0.0123471
R17501 DVSS.n455 DVSS.n454 0.0123471
R17502 DVSS.n454 DVSS.n453 0.0123471
R17503 DVSS.n453 DVSS.n233 0.0123471
R17504 DVSS.n449 DVSS.n233 0.0123471
R17505 DVSS.n449 DVSS.n448 0.0123471
R17506 DVSS.n448 DVSS.n447 0.0123471
R17507 DVSS.n447 DVSS.n235 0.0123471
R17508 DVSS.n443 DVSS.n235 0.0123471
R17509 DVSS.n443 DVSS.n442 0.0123471
R17510 DVSS.n442 DVSS.n441 0.0123471
R17511 DVSS.n441 DVSS.n237 0.0123471
R17512 DVSS.n437 DVSS.n237 0.0123471
R17513 DVSS.n437 DVSS.n436 0.0123471
R17514 DVSS.n436 DVSS.n435 0.0123471
R17515 DVSS.n435 DVSS.n239 0.0123471
R17516 DVSS.n431 DVSS.n239 0.0123471
R17517 DVSS.n431 DVSS.n430 0.0123471
R17518 DVSS.n430 DVSS.n429 0.0123471
R17519 DVSS.n274 DVSS.n273 0.0123471
R17520 DVSS.n277 DVSS.n270 0.0123471
R17521 DVSS.n281 DVSS.n270 0.0123471
R17522 DVSS.n282 DVSS.n281 0.0123471
R17523 DVSS.n283 DVSS.n282 0.0123471
R17524 DVSS.n283 DVSS.n268 0.0123471
R17525 DVSS.n287 DVSS.n268 0.0123471
R17526 DVSS.n288 DVSS.n287 0.0123471
R17527 DVSS.n289 DVSS.n288 0.0123471
R17528 DVSS.n289 DVSS.n266 0.0123471
R17529 DVSS.n293 DVSS.n266 0.0123471
R17530 DVSS.n294 DVSS.n293 0.0123471
R17531 DVSS.n295 DVSS.n294 0.0123471
R17532 DVSS.n295 DVSS.n264 0.0123471
R17533 DVSS.n299 DVSS.n264 0.0123471
R17534 DVSS.n300 DVSS.n299 0.0123471
R17535 DVSS.n301 DVSS.n300 0.0123471
R17536 DVSS.n301 DVSS.n262 0.0123471
R17537 DVSS.n305 DVSS.n262 0.0123471
R17538 DVSS.n306 DVSS.n305 0.0123471
R17539 DVSS.n308 DVSS.n306 0.0123471
R17540 DVSS.n308 DVSS.n307 0.0123471
R17541 DVSS.n1188 DVSS.n1179 0.0123293
R17542 DVSS.n4931 DVSS.n1185 0.0123293
R17543 DVSS.n1858 DVSS.n1383 0.0122701
R17544 DVSS.n4169 DVSS.n1389 0.0122701
R17545 DVSS.n3188 DVSS 0.0122488
R17546 DVSS.n3334 DVSS 0.0122488
R17547 DVSS.n3055 DVSS.n3053 0.012
R17548 DVSS.n3523 DVSS.n3092 0.012
R17549 DVSS.n3050 DVSS.n3049 0.012
R17550 DVSS.n3278 DVSS.n3276 0.012
R17551 DVSS.n2093 DVSS.n2092 0.0116468
R17552 DVSS.n3620 DVSS.n1724 0.0116
R17553 DVSS.n1206 DVSS.n1189 0.0115976
R17554 DVSS.n1200 DVSS.n1184 0.0115976
R17555 DVSS.n3545 DVSS.n3544 0.0115
R17556 DVSS.n3537 DVSS.n3536 0.0115
R17557 DVSS.n3256 DVSS.n2674 0.0115
R17558 DVSS.n3264 DVSS.n3072 0.0115
R17559 DVSS.n2130 DVSS.n1943 0.0113969
R17560 DVSS.n2130 DVSS.n1944 0.0113969
R17561 DVSS.n2200 DVSS.n1754 0.0113969
R17562 DVSS.n2200 DVSS.n2199 0.0113969
R17563 DVSS.n4898 DVSS.n4777 0.0112561
R17564 DVSS.n4887 DVSS.n4788 0.0112561
R17565 DVSS.n4756 DVSS.n1229 0.0112561
R17566 DVSS.n4768 DVSS.n1221 0.0112561
R17567 DVSS.n4716 DVSS.n4715 0.0112561
R17568 DVSS.n4733 DVSS.n1240 0.0112561
R17569 DVSS.n4618 DVSS.n4615 0.0112561
R17570 DVSS.n4693 DVSS.n1261 0.0112561
R17571 DVSS.n4650 DVSS.n4584 0.0112561
R17572 DVSS.n4639 DVSS.n4595 0.0112561
R17573 DVSS.n4563 DVSS.n4503 0.0112561
R17574 DVSS.n4575 DVSS.n4495 0.0112561
R17575 DVSS.n4970 VSS 0.0110882
R17576 DVSS.n1483 VSS 0.0110882
R17577 VSS DVSS.n1168 0.0110882
R17578 DVSS.n5230 DVSS.n1020 0.0110195
R17579 DVSS.n3036 DVSS.n2691 0.011
R17580 DVSS.n3112 DVSS.n3111 0.011
R17581 DVSS.n2695 DVSS.n2689 0.011
R17582 DVSS.n3284 DVSS.n3283 0.011
R17583 DVSS.n3962 DVSS.n1500 0.0109694
R17584 DVSS.n3963 DVSS.n3962 0.0109694
R17585 DVSS.n3964 DVSS.n3963 0.0109694
R17586 DVSS.n3964 DVSS.n1496 0.0109694
R17587 DVSS.n3971 DVSS.n1496 0.0109694
R17588 DVSS.n3972 DVSS.n3971 0.0109694
R17589 DVSS.n3973 DVSS.n3972 0.0109694
R17590 DVSS.n3973 DVSS.n1441 0.0109694
R17591 DVSS.n3980 DVSS.n1441 0.0109694
R17592 DVSS DVSS.n3093 0.0109187
R17593 DVSS.n3269 DVSS 0.0109187
R17594 DVSS.n3629 DVSS.n1724 0.0109
R17595 DVSS.n3643 DVSS.n3629 0.0109
R17596 DVSS.n3643 DVSS.n3642 0.0109
R17597 DVSS.n3642 DVSS.n3641 0.0109
R17598 DVSS.n3641 DVSS.n3640 0.0109
R17599 DVSS.n3640 DVSS.n3639 0.0109
R17600 DVSS.n3639 DVSS.n3638 0.0109
R17601 DVSS.n3638 DVSS.n3637 0.0109
R17602 DVSS.n3637 DVSS.n3636 0.0109
R17603 DVSS.n3636 DVSS.n3635 0.0109
R17604 DVSS.n3635 DVSS.n3634 0.0109
R17605 DVSS.n1208 DVSS.n1187 0.0108659
R17606 DVSS.n1198 DVSS.n1182 0.0108659
R17607 DVSS.n2840 DVSS.n2779 0.010697
R17608 DVSS.n2833 DVSS.n2826 0.010697
R17609 DVSS.n5230 DVSS.n5229 0.0106855
R17610 DVSS.n2988 DVSS.n2714 0.0105
R17611 DVSS.n3494 DVSS.n3135 0.0105
R17612 DVSS.n2929 DVSS.n2716 0.0105
R17613 DVSS.n3306 DVSS.n3137 0.0105
R17614 DVSS.n2810 DVSS.n2793 0.0105
R17615 DVSS.n2810 DVSS.n2809 0.0105
R17616 DVSS.n2809 DVSS.n2808 0.0105
R17617 DVSS.n2808 DVSS.n2775 0.0105
R17618 DVSS.n2846 DVSS.n2775 0.0105
R17619 DVSS.n2846 DVSS.n2773 0.0105
R17620 DVSS.n2854 DVSS.n2773 0.0105
R17621 DVSS.n2854 DVSS.n2853 0.0105
R17622 DVSS.n2853 DVSS.n2852 0.0105
R17623 DVSS.n2852 DVSS.n2755 0.0105
R17624 DVSS.n2895 DVSS.n2755 0.0105
R17625 DVSS.n2895 DVSS.n2753 0.0105
R17626 DVSS.n2907 DVSS.n2753 0.0105
R17627 DVSS.n2907 DVSS.n2906 0.0105
R17628 DVSS.n2906 DVSS.n2903 0.0105
R17629 DVSS.n2903 DVSS.n2902 0.0105
R17630 DVSS.n2902 DVSS.n2733 0.0105
R17631 DVSS.n2958 DVSS.n2733 0.0105
R17632 DVSS.n2958 DVSS.n2731 0.0105
R17633 DVSS.n2962 DVSS.n2731 0.0105
R17634 DVSS.n2962 DVSS.n2720 0.0105
R17635 DVSS.n2977 DVSS.n2720 0.0105
R17636 DVSS.n2977 DVSS.n2718 0.0105
R17637 DVSS.n2985 DVSS.n2718 0.0105
R17638 DVSS.n2985 DVSS.n2984 0.0105
R17639 DVSS.n2984 DVSS.n2983 0.0105
R17640 DVSS.n2983 DVSS.n2700 0.0105
R17641 DVSS.n3023 DVSS.n2700 0.0105
R17642 DVSS.n3023 DVSS.n2698 0.0105
R17643 DVSS.n3032 DVSS.n2698 0.0105
R17644 DVSS.n3032 DVSS.n3031 0.0105
R17645 DVSS.n3031 DVSS.n3030 0.0105
R17646 DVSS.n3030 DVSS.n2678 0.0105
R17647 DVSS.n3064 DVSS.n2678 0.0105
R17648 DVSS.n3065 DVSS.n3064 0.0105
R17649 DVSS.n3066 DVSS.n3065 0.0105
R17650 DVSS.n3066 DVSS.n2676 0.0105
R17651 DVSS.n3541 DVSS.n2676 0.0105
R17652 DVSS.n3541 DVSS.n3540 0.0105
R17653 DVSS.n3540 DVSS.n3071 0.0105
R17654 DVSS.n3083 DVSS.n3071 0.0105
R17655 DVSS.n3528 DVSS.n3083 0.0105
R17656 DVSS.n3528 DVSS.n3527 0.0105
R17657 DVSS.n3527 DVSS.n3088 0.0105
R17658 DVSS.n3103 DVSS.n3088 0.0105
R17659 DVSS.n3516 DVSS.n3103 0.0105
R17660 DVSS.n3516 DVSS.n3515 0.0105
R17661 DVSS.n3515 DVSS.n3108 0.0105
R17662 DVSS.n3120 DVSS.n3108 0.0105
R17663 DVSS.n3503 DVSS.n3120 0.0105
R17664 DVSS.n3503 DVSS.n3502 0.0105
R17665 DVSS.n3502 DVSS.n3125 0.0105
R17666 DVSS.n3139 DVSS.n3125 0.0105
R17667 DVSS.n3491 DVSS.n3139 0.0105
R17668 DVSS.n3491 DVSS.n3490 0.0105
R17669 DVSS.n3490 DVSS.n3144 0.0105
R17670 DVSS.n3157 DVSS.n3144 0.0105
R17671 DVSS.n3477 DVSS.n3157 0.0105
R17672 DVSS.n3477 DVSS.n3476 0.0105
R17673 DVSS.n3476 DVSS.n3162 0.0105
R17674 DVSS.n3174 DVSS.n3162 0.0105
R17675 DVSS.n3465 DVSS.n3174 0.0105
R17676 DVSS.n3465 DVSS.n3464 0.0105
R17677 DVSS.n3464 DVSS.n3179 0.0105
R17678 DVSS.n3194 DVSS.n3179 0.0105
R17679 DVSS.n3453 DVSS.n3194 0.0105
R17680 DVSS.n3453 DVSS.n3452 0.0105
R17681 DVSS.n3452 DVSS.n3199 0.0105
R17682 DVSS.n3212 DVSS.n3199 0.0105
R17683 DVSS.n3441 DVSS.n3212 0.0105
R17684 DVSS.n3441 DVSS.n3440 0.0105
R17685 DVSS.n3440 DVSS.n3217 0.0105
R17686 DVSS.n3229 DVSS.n3217 0.0105
R17687 DVSS.n3428 DVSS.n3229 0.0105
R17688 DVSS.n3428 DVSS.n3427 0.0105
R17689 DVSS.n3427 DVSS.n3234 0.0105
R17690 DVSS.n3377 DVSS.n3234 0.0105
R17691 DVSS.n3416 DVSS.n3377 0.0105
R17692 DVSS.n3416 DVSS.n3415 0.0105
R17693 DVSS.n3415 DVSS.n3414 0.0105
R17694 DVSS.n3414 DVSS.n3383 0.0105
R17695 DVSS.n3410 DVSS.n3383 0.0105
R17696 DVSS.n3410 DVSS.n3409 0.0105
R17697 DVSS.n3409 DVSS.n3387 0.0105
R17698 DVSS.n3405 DVSS.n3387 0.0105
R17699 DVSS.n3405 DVSS.n3404 0.0105
R17700 DVSS.n3404 DVSS.n3403 0.0105
R17701 DVSS.n3403 DVSS.n3393 0.0105
R17702 DVSS.n3399 DVSS.n3393 0.0105
R17703 DVSS.n3417 DVSS.n3376 0.0105
R17704 DVSS.n3413 DVSS.n3376 0.0105
R17705 DVSS.n3413 DVSS.n3412 0.0105
R17706 DVSS.n3412 DVSS.n3411 0.0105
R17707 DVSS.n3408 DVSS.n3407 0.0105
R17708 DVSS.n3407 DVSS.n3406 0.0105
R17709 DVSS.n3406 DVSS.n3388 0.0105
R17710 DVSS.n3402 DVSS.n3388 0.0105
R17711 DVSS.n3402 DVSS.n3401 0.0105
R17712 DVSS.n3401 DVSS.n3400 0.0105
R17713 DVSS.n3408 DVSS.n1706 0.0104296
R17714 DVSS.n5562 DVSS.n826 0.0103531
R17715 DVSS.n5814 DVSS.n3 0.0103531
R17716 DVSS.n5808 DVSS.n27 0.0103531
R17717 DVSS.n4899 DVSS.n4898 0.0101185
R17718 DVSS.n4885 DVSS.n4788 0.0101185
R17719 DVSS.n4754 DVSS.n1229 0.0101185
R17720 DVSS.n4769 DVSS.n4768 0.0101185
R17721 DVSS.n4715 DVSS.n1251 0.0101185
R17722 DVSS.n4735 DVSS.n1240 0.0101185
R17723 DVSS.n4619 DVSS.n4618 0.0101185
R17724 DVSS.n4695 DVSS.n1261 0.0101185
R17725 DVSS.n4651 DVSS.n4650 0.0101185
R17726 DVSS.n4637 DVSS.n4595 0.0101185
R17727 DVSS.n4561 DVSS.n4503 0.0101185
R17728 DVSS.n4576 DVSS.n4575 0.0101185
R17729 DVSS.n5554 DVSS.n848 0.0100456
R17730 DVSS.n1192 DVSS.n1191 0.0100456
R17731 DVSS.n4932 DVSS.n852 0.0100456
R17732 DVSS.n1192 DVSS.n850 0.0100456
R17733 DVSS.n2949 DVSS.n2738 0.01
R17734 DVSS.n3469 DVSS.n3167 0.01
R17735 DVSS.n2946 DVSS.n2740 0.01
R17736 DVSS.n3326 DVSS.n3325 0.01
R17737 DVSS.n3586 DVSS 0.00997368
R17738 DVSS.n1855 DVSS.n1382 0.00965456
R17739 DVSS.n1837 DVSS.n1388 0.00965456
R17740 DVSS.n953 DVSS.n950 0.00962857
R17741 DVSS.n5364 DVSS.n950 0.00962857
R17742 DVSS.n5364 DVSS.n948 0.00962857
R17743 DVSS.n5368 DVSS.n948 0.00962857
R17744 DVSS.n5368 DVSS.n946 0.00962857
R17745 DVSS.n5372 DVSS.n946 0.00962857
R17746 DVSS.n5372 DVSS.n944 0.00962857
R17747 DVSS.n5376 DVSS.n944 0.00962857
R17748 DVSS.n5376 DVSS.n942 0.00962857
R17749 DVSS.n5380 DVSS.n942 0.00962857
R17750 DVSS.n5380 DVSS.n940 0.00962857
R17751 DVSS.n5384 DVSS.n940 0.00962857
R17752 DVSS.n5384 DVSS.n938 0.00962857
R17753 DVSS.n5388 DVSS.n938 0.00962857
R17754 DVSS.n5388 DVSS.n936 0.00962857
R17755 DVSS.n5392 DVSS.n936 0.00962857
R17756 DVSS.n5392 DVSS.n934 0.00962857
R17757 DVSS.n5396 DVSS.n934 0.00962857
R17758 DVSS.n5396 DVSS.n932 0.00962857
R17759 DVSS.n5400 DVSS.n932 0.00962857
R17760 DVSS.n5400 DVSS.n930 0.00962857
R17761 DVSS.n5404 DVSS.n930 0.00962857
R17762 DVSS.n5404 DVSS.n928 0.00962857
R17763 DVSS.n5408 DVSS.n928 0.00962857
R17764 DVSS.n5408 DVSS.n926 0.00962857
R17765 DVSS.n5412 DVSS.n926 0.00962857
R17766 DVSS.n5412 DVSS.n924 0.00962857
R17767 DVSS.n5416 DVSS.n924 0.00962857
R17768 DVSS.n5416 DVSS.n922 0.00962857
R17769 DVSS.n5420 DVSS.n922 0.00962857
R17770 DVSS.n5420 DVSS.n920 0.00962857
R17771 DVSS.n5424 DVSS.n920 0.00962857
R17772 DVSS.n5424 DVSS.n918 0.00962857
R17773 DVSS.n5428 DVSS.n918 0.00962857
R17774 DVSS.n5428 DVSS.n916 0.00962857
R17775 DVSS.n5432 DVSS.n916 0.00962857
R17776 DVSS.n5432 DVSS.n914 0.00962857
R17777 DVSS.n5436 DVSS.n914 0.00962857
R17778 DVSS.n5436 DVSS.n912 0.00962857
R17779 DVSS.n5440 DVSS.n912 0.00962857
R17780 DVSS.n5440 DVSS.n910 0.00962857
R17781 DVSS.n5444 DVSS.n910 0.00962857
R17782 DVSS.n5444 DVSS.n908 0.00962857
R17783 DVSS.n5448 DVSS.n908 0.00962857
R17784 DVSS.n5448 DVSS.n906 0.00962857
R17785 DVSS.n5452 DVSS.n906 0.00962857
R17786 DVSS.n5452 DVSS.n904 0.00962857
R17787 DVSS.n5456 DVSS.n904 0.00962857
R17788 DVSS.n5456 DVSS.n902 0.00962857
R17789 DVSS.n5460 DVSS.n902 0.00962857
R17790 DVSS.n5460 DVSS.n900 0.00962857
R17791 DVSS.n5464 DVSS.n900 0.00962857
R17792 DVSS.n5464 DVSS.n898 0.00962857
R17793 DVSS.n5468 DVSS.n898 0.00962857
R17794 DVSS.n5468 DVSS.n896 0.00962857
R17795 DVSS.n5472 DVSS.n896 0.00962857
R17796 DVSS.n5472 DVSS.n894 0.00962857
R17797 DVSS.n5476 DVSS.n894 0.00962857
R17798 DVSS.n5476 DVSS.n892 0.00962857
R17799 DVSS.n5480 DVSS.n892 0.00962857
R17800 DVSS.n5480 DVSS.n890 0.00962857
R17801 DVSS.n5484 DVSS.n890 0.00962857
R17802 DVSS.n5484 DVSS.n888 0.00962857
R17803 DVSS.n5488 DVSS.n888 0.00962857
R17804 DVSS.n5488 DVSS.n886 0.00962857
R17805 DVSS.n5492 DVSS.n886 0.00962857
R17806 DVSS.n5492 DVSS.n884 0.00962857
R17807 DVSS.n5496 DVSS.n884 0.00962857
R17808 DVSS.n5496 DVSS.n882 0.00962857
R17809 DVSS.n5500 DVSS.n882 0.00962857
R17810 DVSS.n5500 DVSS.n880 0.00962857
R17811 DVSS.n5504 DVSS.n880 0.00962857
R17812 DVSS.n5504 DVSS.n878 0.00962857
R17813 DVSS.n5508 DVSS.n878 0.00962857
R17814 DVSS.n5508 DVSS.n876 0.00962857
R17815 DVSS.n5512 DVSS.n876 0.00962857
R17816 DVSS.n5512 DVSS.n874 0.00962857
R17817 DVSS.n5516 DVSS.n874 0.00962857
R17818 DVSS.n5516 DVSS.n872 0.00962857
R17819 DVSS.n5520 DVSS.n872 0.00962857
R17820 DVSS.n5520 DVSS.n870 0.00962857
R17821 DVSS.n5524 DVSS.n870 0.00962857
R17822 DVSS.n5524 DVSS.n868 0.00962857
R17823 DVSS.n5528 DVSS.n868 0.00962857
R17824 DVSS.n5528 DVSS.n866 0.00962857
R17825 DVSS.n5532 DVSS.n866 0.00962857
R17826 DVSS.n5532 DVSS.n864 0.00962857
R17827 DVSS.n5536 DVSS.n864 0.00962857
R17828 DVSS.n5536 DVSS.n862 0.00962857
R17829 DVSS.n5540 DVSS.n862 0.00962857
R17830 DVSS.n5540 DVSS.n860 0.00962857
R17831 DVSS.n5544 DVSS.n860 0.00962857
R17832 DVSS.n5544 DVSS.n858 0.00962857
R17833 DVSS.n5548 DVSS.n858 0.00962857
R17834 DVSS.n5363 DVSS.n5362 0.00962857
R17835 DVSS.n5363 DVSS.n947 0.00962857
R17836 DVSS.n5369 DVSS.n947 0.00962857
R17837 DVSS.n5370 DVSS.n5369 0.00962857
R17838 DVSS.n5371 DVSS.n5370 0.00962857
R17839 DVSS.n5371 DVSS.n943 0.00962857
R17840 DVSS.n5377 DVSS.n943 0.00962857
R17841 DVSS.n5378 DVSS.n5377 0.00962857
R17842 DVSS.n5379 DVSS.n5378 0.00962857
R17843 DVSS.n5379 DVSS.n939 0.00962857
R17844 DVSS.n5385 DVSS.n939 0.00962857
R17845 DVSS.n5386 DVSS.n5385 0.00962857
R17846 DVSS.n5387 DVSS.n5386 0.00962857
R17847 DVSS.n5387 DVSS.n935 0.00962857
R17848 DVSS.n5393 DVSS.n935 0.00962857
R17849 DVSS.n5394 DVSS.n5393 0.00962857
R17850 DVSS.n5395 DVSS.n5394 0.00962857
R17851 DVSS.n5395 DVSS.n931 0.00962857
R17852 DVSS.n5401 DVSS.n931 0.00962857
R17853 DVSS.n5402 DVSS.n5401 0.00962857
R17854 DVSS.n5403 DVSS.n5402 0.00962857
R17855 DVSS.n5403 DVSS.n927 0.00962857
R17856 DVSS.n5409 DVSS.n927 0.00962857
R17857 DVSS.n5410 DVSS.n5409 0.00962857
R17858 DVSS.n5411 DVSS.n5410 0.00962857
R17859 DVSS.n5411 DVSS.n923 0.00962857
R17860 DVSS.n5417 DVSS.n923 0.00962857
R17861 DVSS.n5418 DVSS.n5417 0.00962857
R17862 DVSS.n5419 DVSS.n5418 0.00962857
R17863 DVSS.n5419 DVSS.n919 0.00962857
R17864 DVSS.n5425 DVSS.n919 0.00962857
R17865 DVSS.n5426 DVSS.n5425 0.00962857
R17866 DVSS.n5427 DVSS.n5426 0.00962857
R17867 DVSS.n5427 DVSS.n915 0.00962857
R17868 DVSS.n5433 DVSS.n915 0.00962857
R17869 DVSS.n5434 DVSS.n5433 0.00962857
R17870 DVSS.n5435 DVSS.n5434 0.00962857
R17871 DVSS.n5435 DVSS.n911 0.00962857
R17872 DVSS.n5441 DVSS.n911 0.00962857
R17873 DVSS.n5442 DVSS.n5441 0.00962857
R17874 DVSS.n5443 DVSS.n5442 0.00962857
R17875 DVSS.n5443 DVSS.n907 0.00962857
R17876 DVSS.n5449 DVSS.n907 0.00962857
R17877 DVSS.n5450 DVSS.n5449 0.00962857
R17878 DVSS.n5451 DVSS.n5450 0.00962857
R17879 DVSS.n5451 DVSS.n903 0.00962857
R17880 DVSS.n5457 DVSS.n903 0.00962857
R17881 DVSS.n5458 DVSS.n5457 0.00962857
R17882 DVSS.n5459 DVSS.n5458 0.00962857
R17883 DVSS.n5459 DVSS.n899 0.00962857
R17884 DVSS.n5465 DVSS.n899 0.00962857
R17885 DVSS.n5466 DVSS.n5465 0.00962857
R17886 DVSS.n5467 DVSS.n5466 0.00962857
R17887 DVSS.n5467 DVSS.n895 0.00962857
R17888 DVSS.n5473 DVSS.n895 0.00962857
R17889 DVSS.n5474 DVSS.n5473 0.00962857
R17890 DVSS.n5475 DVSS.n5474 0.00962857
R17891 DVSS.n5475 DVSS.n891 0.00962857
R17892 DVSS.n5481 DVSS.n891 0.00962857
R17893 DVSS.n5482 DVSS.n5481 0.00962857
R17894 DVSS.n5483 DVSS.n5482 0.00962857
R17895 DVSS.n5483 DVSS.n887 0.00962857
R17896 DVSS.n5489 DVSS.n887 0.00962857
R17897 DVSS.n5490 DVSS.n5489 0.00962857
R17898 DVSS.n5491 DVSS.n5490 0.00962857
R17899 DVSS.n5491 DVSS.n883 0.00962857
R17900 DVSS.n5497 DVSS.n883 0.00962857
R17901 DVSS.n5498 DVSS.n5497 0.00962857
R17902 DVSS.n5499 DVSS.n5498 0.00962857
R17903 DVSS.n5499 DVSS.n879 0.00962857
R17904 DVSS.n5505 DVSS.n879 0.00962857
R17905 DVSS.n5506 DVSS.n5505 0.00962857
R17906 DVSS.n5507 DVSS.n5506 0.00962857
R17907 DVSS.n5507 DVSS.n875 0.00962857
R17908 DVSS.n5513 DVSS.n875 0.00962857
R17909 DVSS.n5514 DVSS.n5513 0.00962857
R17910 DVSS.n5515 DVSS.n5514 0.00962857
R17911 DVSS.n5515 DVSS.n871 0.00962857
R17912 DVSS.n5521 DVSS.n871 0.00962857
R17913 DVSS.n5522 DVSS.n5521 0.00962857
R17914 DVSS.n5523 DVSS.n5522 0.00962857
R17915 DVSS.n5523 DVSS.n867 0.00962857
R17916 DVSS.n5529 DVSS.n867 0.00962857
R17917 DVSS.n5530 DVSS.n5529 0.00962857
R17918 DVSS.n5531 DVSS.n5530 0.00962857
R17919 DVSS.n5531 DVSS.n863 0.00962857
R17920 DVSS.n5537 DVSS.n863 0.00962857
R17921 DVSS.n5538 DVSS.n5537 0.00962857
R17922 DVSS.n5539 DVSS.n5538 0.00962857
R17923 DVSS.n5539 DVSS.n859 0.00962857
R17924 DVSS.n5545 DVSS.n859 0.00962857
R17925 DVSS.n5546 DVSS.n5545 0.00962857
R17926 DVSS.n5547 DVSS.n5546 0.00962857
R17927 DVSS.n4546 DVSS.n4510 0.00962857
R17928 DVSS.n4550 DVSS.n4510 0.00962857
R17929 DVSS.n4550 DVSS.n4508 0.00962857
R17930 DVSS.n4554 DVSS.n4508 0.00962857
R17931 DVSS.n4554 DVSS.n4506 0.00962857
R17932 DVSS.n4558 DVSS.n4506 0.00962857
R17933 DVSS.n4558 DVSS.n4501 0.00962857
R17934 DVSS.n4569 DVSS.n4501 0.00962857
R17935 DVSS.n4569 DVSS.n4498 0.00962857
R17936 DVSS.n4667 DVSS.n4498 0.00962857
R17937 DVSS.n4667 DVSS.n4499 0.00962857
R17938 DVSS.n4663 DVSS.n4499 0.00962857
R17939 DVSS.n4663 DVSS.n4573 0.00962857
R17940 DVSS.n4659 DVSS.n4573 0.00962857
R17941 DVSS.n4659 DVSS.n4579 0.00962857
R17942 DVSS.n4655 DVSS.n4579 0.00962857
R17943 DVSS.n4655 DVSS.n4581 0.00962857
R17944 DVSS.n4586 DVSS.n4581 0.00962857
R17945 DVSS.n4647 DVSS.n4586 0.00962857
R17946 DVSS.n4647 DVSS.n4587 0.00962857
R17947 DVSS.n4643 DVSS.n4587 0.00962857
R17948 DVSS.n4643 DVSS.n4590 0.00962857
R17949 DVSS.n4605 DVSS.n4590 0.00962857
R17950 DVSS.n4634 DVSS.n4605 0.00962857
R17951 DVSS.n4634 DVSS.n4606 0.00962857
R17952 DVSS.n4630 DVSS.n4606 0.00962857
R17953 DVSS.n4630 DVSS.n4609 0.00962857
R17954 DVSS.n4626 DVSS.n4609 0.00962857
R17955 DVSS.n4626 DVSS.n4611 0.00962857
R17956 DVSS.n4622 DVSS.n4611 0.00962857
R17957 DVSS.n4622 DVSS.n4613 0.00962857
R17958 DVSS.n4613 DVSS.n1268 0.00962857
R17959 DVSS.n4685 DVSS.n1268 0.00962857
R17960 DVSS.n4685 DVSS.n1266 0.00962857
R17961 DVSS.n4689 DVSS.n1266 0.00962857
R17962 DVSS.n4689 DVSS.n1259 0.00962857
R17963 DVSS.n4698 DVSS.n1259 0.00962857
R17964 DVSS.n4698 DVSS.n1257 0.00962857
R17965 DVSS.n4702 DVSS.n1257 0.00962857
R17966 DVSS.n4702 DVSS.n1255 0.00962857
R17967 DVSS.n4707 DVSS.n1255 0.00962857
R17968 DVSS.n4707 DVSS.n1253 0.00962857
R17969 DVSS.n4711 DVSS.n1253 0.00962857
R17970 DVSS.n4711 DVSS.n1248 0.00962857
R17971 DVSS.n4724 DVSS.n1248 0.00962857
R17972 DVSS.n4724 DVSS.n1245 0.00962857
R17973 DVSS.n4729 DVSS.n1245 0.00962857
R17974 DVSS.n4729 DVSS.n1246 0.00962857
R17975 DVSS.n1246 DVSS.n1238 0.00962857
R17976 DVSS.n4739 DVSS.n1238 0.00962857
R17977 DVSS.n4739 DVSS.n1236 0.00962857
R17978 DVSS.n4743 DVSS.n1236 0.00962857
R17979 DVSS.n4743 DVSS.n1234 0.00962857
R17980 DVSS.n4747 DVSS.n1234 0.00962857
R17981 DVSS.n4747 DVSS.n1232 0.00962857
R17982 DVSS.n4751 DVSS.n1232 0.00962857
R17983 DVSS.n4751 DVSS.n1227 0.00962857
R17984 DVSS.n4762 DVSS.n1227 0.00962857
R17985 DVSS.n4762 DVSS.n1224 0.00962857
R17986 DVSS.n4915 DVSS.n1224 0.00962857
R17987 DVSS.n4915 DVSS.n1225 0.00962857
R17988 DVSS.n4911 DVSS.n1225 0.00962857
R17989 DVSS.n4911 DVSS.n4766 0.00962857
R17990 DVSS.n4907 DVSS.n4766 0.00962857
R17991 DVSS.n4907 DVSS.n4772 0.00962857
R17992 DVSS.n4903 DVSS.n4772 0.00962857
R17993 DVSS.n4903 DVSS.n4774 0.00962857
R17994 DVSS.n4779 DVSS.n4774 0.00962857
R17995 DVSS.n4895 DVSS.n4779 0.00962857
R17996 DVSS.n4895 DVSS.n4780 0.00962857
R17997 DVSS.n4891 DVSS.n4780 0.00962857
R17998 DVSS.n4891 DVSS.n4783 0.00962857
R17999 DVSS.n4798 DVSS.n4783 0.00962857
R18000 DVSS.n4882 DVSS.n4798 0.00962857
R18001 DVSS.n4882 DVSS.n4799 0.00962857
R18002 DVSS.n4878 DVSS.n4799 0.00962857
R18003 DVSS.n4878 DVSS.n4802 0.00962857
R18004 DVSS.n4838 DVSS.n4802 0.00962857
R18005 DVSS.n4838 DVSS.n4836 0.00962857
R18006 DVSS.n4870 DVSS.n4836 0.00962857
R18007 DVSS.n4870 DVSS.n4837 0.00962857
R18008 DVSS.n4866 DVSS.n4837 0.00962857
R18009 DVSS.n4866 DVSS.n4842 0.00962857
R18010 DVSS.n4862 DVSS.n4842 0.00962857
R18011 DVSS.n4862 DVSS.n4844 0.00962857
R18012 DVSS.n4858 DVSS.n4844 0.00962857
R18013 DVSS.n4857 DVSS.n4855 0.00962857
R18014 DVSS.n4855 DVSS.n4846 0.00962857
R18015 DVSS.n4851 DVSS.n4846 0.00962857
R18016 DVSS.n4552 DVSS.n4551 0.00962857
R18017 DVSS.n4553 DVSS.n4552 0.00962857
R18018 DVSS.n4553 DVSS.n4504 0.00962857
R18019 DVSS.n4662 DVSS.n4661 0.00962857
R18020 DVSS.n4661 DVSS.n4660 0.00962857
R18021 DVSS.n4660 DVSS.n4578 0.00962857
R18022 DVSS.n4654 DVSS.n4578 0.00962857
R18023 DVSS.n4654 DVSS.n4653 0.00962857
R18024 DVSS.n4635 DVSS.n4604 0.00962857
R18025 DVSS.n4629 DVSS.n4604 0.00962857
R18026 DVSS.n4629 DVSS.n4628 0.00962857
R18027 DVSS.n4628 DVSS.n4627 0.00962857
R18028 DVSS.n4627 DVSS.n4610 0.00962857
R18029 DVSS.n4621 DVSS.n4610 0.00962857
R18030 DVSS.n4697 DVSS.n1256 0.00962857
R18031 DVSS.n4703 DVSS.n1256 0.00962857
R18032 DVSS.n4704 DVSS.n4703 0.00962857
R18033 DVSS.n4706 DVSS.n4704 0.00962857
R18034 DVSS.n4706 DVSS.n4705 0.00962857
R18035 DVSS.n4738 DVSS.n4737 0.00962857
R18036 DVSS.n4738 DVSS.n1235 0.00962857
R18037 DVSS.n4744 DVSS.n1235 0.00962857
R18038 DVSS.n4745 DVSS.n4744 0.00962857
R18039 DVSS.n4746 DVSS.n4745 0.00962857
R18040 DVSS.n4746 DVSS.n1230 0.00962857
R18041 DVSS.n4910 DVSS.n4909 0.00962857
R18042 DVSS.n4909 DVSS.n4908 0.00962857
R18043 DVSS.n4908 DVSS.n4771 0.00962857
R18044 DVSS.n4902 DVSS.n4771 0.00962857
R18045 DVSS.n4902 DVSS.n4901 0.00962857
R18046 DVSS.n4883 DVSS.n4797 0.00962857
R18047 DVSS.n4877 DVSS.n4797 0.00962857
R18048 DVSS.n4877 DVSS.n4876 0.00962857
R18049 DVSS.n4871 DVSS.n4835 0.00962857
R18050 DVSS.n4865 DVSS.n4835 0.00962857
R18051 DVSS.n4865 DVSS.n4864 0.00962857
R18052 DVSS.n4864 DVSS.n4863 0.00962857
R18053 DVSS.n4863 DVSS.n4843 0.00962857
R18054 DVSS.n4843 DVSS.n1181 0.00962857
R18055 DVSS.n4854 DVSS.n4853 0.00962857
R18056 DVSS.n4853 DVSS.n4852 0.00962857
R18057 DVSS.n1536 DVSS.n1533 0.00962857
R18058 DVSS.n1540 DVSS.n1533 0.00962857
R18059 DVSS.n1540 DVSS.n1531 0.00962857
R18060 DVSS.n1544 DVSS.n1531 0.00962857
R18061 DVSS.n1544 DVSS.n1529 0.00962857
R18062 DVSS.n1548 DVSS.n1529 0.00962857
R18063 DVSS.n1548 DVSS.n1527 0.00962857
R18064 DVSS.n1552 DVSS.n1527 0.00962857
R18065 DVSS.n1552 DVSS.n1525 0.00962857
R18066 DVSS.n1556 DVSS.n1525 0.00962857
R18067 DVSS.n1556 DVSS.n1522 0.00962857
R18068 DVSS.n3935 DVSS.n1522 0.00962857
R18069 DVSS.n3935 DVSS.n1523 0.00962857
R18070 DVSS.n3931 DVSS.n1523 0.00962857
R18071 DVSS.n3931 DVSS.n1560 0.00962857
R18072 DVSS.n3927 DVSS.n1560 0.00962857
R18073 DVSS.n3927 DVSS.n1562 0.00962857
R18074 DVSS.n3923 DVSS.n1562 0.00962857
R18075 DVSS.n3923 DVSS.n1564 0.00962857
R18076 DVSS.n3919 DVSS.n1564 0.00962857
R18077 DVSS.n3919 DVSS.n1566 0.00962857
R18078 DVSS.n3915 DVSS.n1566 0.00962857
R18079 DVSS.n3915 DVSS.n1568 0.00962857
R18080 DVSS.n3911 DVSS.n1568 0.00962857
R18081 DVSS.n3911 DVSS.n1570 0.00962857
R18082 DVSS.n3907 DVSS.n1570 0.00962857
R18083 DVSS.n3907 DVSS.n1572 0.00962857
R18084 DVSS.n2494 DVSS.n1572 0.00962857
R18085 DVSS.n2497 DVSS.n2494 0.00962857
R18086 DVSS.n2497 DVSS.n2492 0.00962857
R18087 DVSS.n2501 DVSS.n2492 0.00962857
R18088 DVSS.n2501 DVSS.n2490 0.00962857
R18089 DVSS.n2505 DVSS.n2490 0.00962857
R18090 DVSS.n2505 DVSS.n2488 0.00962857
R18091 DVSS.n2509 DVSS.n2488 0.00962857
R18092 DVSS.n2509 DVSS.n2486 0.00962857
R18093 DVSS.n2513 DVSS.n2486 0.00962857
R18094 DVSS.n2513 DVSS.n2484 0.00962857
R18095 DVSS.n2517 DVSS.n2484 0.00962857
R18096 DVSS.n2517 DVSS.n2482 0.00962857
R18097 DVSS.n2521 DVSS.n2482 0.00962857
R18098 DVSS.n2521 DVSS.n2480 0.00962857
R18099 DVSS.n2525 DVSS.n2480 0.00962857
R18100 DVSS.n2525 DVSS.n2478 0.00962857
R18101 DVSS.n2529 DVSS.n2478 0.00962857
R18102 DVSS.n2529 DVSS.n2476 0.00962857
R18103 DVSS.n2533 DVSS.n2476 0.00962857
R18104 DVSS.n2533 DVSS.n2474 0.00962857
R18105 DVSS.n2537 DVSS.n2474 0.00962857
R18106 DVSS.n2537 DVSS.n2472 0.00962857
R18107 DVSS.n2541 DVSS.n2472 0.00962857
R18108 DVSS.n2541 DVSS.n2470 0.00962857
R18109 DVSS.n2545 DVSS.n2470 0.00962857
R18110 DVSS.n2545 DVSS.n2468 0.00962857
R18111 DVSS.n2549 DVSS.n2468 0.00962857
R18112 DVSS.n2549 DVSS.n2466 0.00962857
R18113 DVSS.n2553 DVSS.n2466 0.00962857
R18114 DVSS.n2553 DVSS.n2464 0.00962857
R18115 DVSS.n2557 DVSS.n2464 0.00962857
R18116 DVSS.n2557 DVSS.n2462 0.00962857
R18117 DVSS.n2561 DVSS.n2462 0.00962857
R18118 DVSS.n2561 DVSS.n2460 0.00962857
R18119 DVSS.n2565 DVSS.n2460 0.00962857
R18120 DVSS.n2565 DVSS.n2458 0.00962857
R18121 DVSS.n2569 DVSS.n2458 0.00962857
R18122 DVSS.n2569 DVSS.n2456 0.00962857
R18123 DVSS.n2573 DVSS.n2456 0.00962857
R18124 DVSS.n2573 DVSS.n2454 0.00962857
R18125 DVSS.n2577 DVSS.n2454 0.00962857
R18126 DVSS.n2577 DVSS.n2452 0.00962857
R18127 DVSS.n2581 DVSS.n2452 0.00962857
R18128 DVSS.n2581 DVSS.n2450 0.00962857
R18129 DVSS.n2585 DVSS.n2450 0.00962857
R18130 DVSS.n2585 DVSS.n2448 0.00962857
R18131 DVSS.n2589 DVSS.n2448 0.00962857
R18132 DVSS.n2589 DVSS.n2446 0.00962857
R18133 DVSS.n2593 DVSS.n2446 0.00962857
R18134 DVSS.n2593 DVSS.n2444 0.00962857
R18135 DVSS.n2597 DVSS.n2444 0.00962857
R18136 DVSS.n2597 DVSS.n2442 0.00962857
R18137 DVSS.n2601 DVSS.n2442 0.00962857
R18138 DVSS.n2601 DVSS.n2440 0.00962857
R18139 DVSS.n2605 DVSS.n2440 0.00962857
R18140 DVSS.n2605 DVSS.n2438 0.00962857
R18141 DVSS.n2609 DVSS.n2438 0.00962857
R18142 DVSS.n2609 DVSS.n2436 0.00962857
R18143 DVSS.n2613 DVSS.n2436 0.00962857
R18144 DVSS.n2613 DVSS.n2434 0.00962857
R18145 DVSS.n2617 DVSS.n2434 0.00962857
R18146 DVSS.n2617 DVSS.n2432 0.00962857
R18147 DVSS.n2621 DVSS.n2432 0.00962857
R18148 DVSS.n2621 DVSS.n2430 0.00962857
R18149 DVSS.n2625 DVSS.n2430 0.00962857
R18150 DVSS.n2625 DVSS.n2428 0.00962857
R18151 DVSS.n2629 DVSS.n2428 0.00962857
R18152 DVSS.n2629 DVSS.n2426 0.00962857
R18153 DVSS.n2635 DVSS.n2426 0.00962857
R18154 DVSS.n2632 DVSS.n2268 0.00962857
R18155 DVSS.n2651 DVSS.n2268 0.00962857
R18156 DVSS.n2651 DVSS.n2266 0.00962857
R18157 DVSS.n1596 DVSS.n1592 0.00962857
R18158 DVSS.n3892 DVSS.n1592 0.00962857
R18159 DVSS.n3892 DVSS.n1593 0.00962857
R18160 DVSS.n3888 DVSS.n1593 0.00962857
R18161 DVSS.n3888 DVSS.n1600 0.00962857
R18162 DVSS.n3883 DVSS.n1600 0.00962857
R18163 DVSS.n3883 DVSS.n1602 0.00962857
R18164 DVSS.n3879 DVSS.n1602 0.00962857
R18165 DVSS.n3879 DVSS.n1604 0.00962857
R18166 DVSS.n3873 DVSS.n1604 0.00962857
R18167 DVSS.n3873 DVSS.n1606 0.00962857
R18168 DVSS.n3869 DVSS.n1606 0.00962857
R18169 DVSS.n3869 DVSS.n1608 0.00962857
R18170 DVSS.n3865 DVSS.n1608 0.00962857
R18171 DVSS.n3865 DVSS.n1611 0.00962857
R18172 DVSS.n3861 DVSS.n1611 0.00962857
R18173 DVSS.n3861 DVSS.n1613 0.00962857
R18174 DVSS.n3854 DVSS.n1613 0.00962857
R18175 DVSS.n3854 DVSS.n1616 0.00962857
R18176 DVSS.n3850 DVSS.n1616 0.00962857
R18177 DVSS.n3850 DVSS.n1618 0.00962857
R18178 DVSS.n3846 DVSS.n1618 0.00962857
R18179 DVSS.n3846 DVSS.n1621 0.00962857
R18180 DVSS.n3842 DVSS.n1621 0.00962857
R18181 DVSS.n3842 DVSS.n1623 0.00962857
R18182 DVSS.n3826 DVSS.n1623 0.00962857
R18183 DVSS.n3826 DVSS.n3825 0.00962857
R18184 DVSS.n3825 DVSS.n1635 0.00962857
R18185 DVSS.n3821 DVSS.n1635 0.00962857
R18186 DVSS.n3821 DVSS.n1637 0.00962857
R18187 DVSS.n3817 DVSS.n1637 0.00962857
R18188 DVSS.n3817 DVSS.n1640 0.00962857
R18189 DVSS.n3813 DVSS.n1640 0.00962857
R18190 DVSS.n3813 DVSS.n1642 0.00962857
R18191 DVSS.n3809 DVSS.n1642 0.00962857
R18192 DVSS.n3809 DVSS.n1644 0.00962857
R18193 DVSS.n3805 DVSS.n1644 0.00962857
R18194 DVSS.n3805 DVSS.n1646 0.00962857
R18195 DVSS.n3800 DVSS.n1646 0.00962857
R18196 DVSS.n3800 DVSS.n1650 0.00962857
R18197 DVSS.n3796 DVSS.n1650 0.00962857
R18198 DVSS.n3796 DVSS.n1652 0.00962857
R18199 DVSS.n1668 DVSS.n1652 0.00962857
R18200 DVSS.n1668 DVSS.n1666 0.00962857
R18201 DVSS.n1676 DVSS.n1666 0.00962857
R18202 DVSS.n1676 DVSS.n1663 0.00962857
R18203 DVSS.n3785 DVSS.n1663 0.00962857
R18204 DVSS.n3785 DVSS.n1664 0.00962857
R18205 DVSS.n3781 DVSS.n1664 0.00962857
R18206 DVSS.n3781 DVSS.n1680 0.00962857
R18207 DVSS.n3777 DVSS.n1680 0.00962857
R18208 DVSS.n3777 DVSS.n1683 0.00962857
R18209 DVSS.n3773 DVSS.n1683 0.00962857
R18210 DVSS.n3773 DVSS.n1685 0.00962857
R18211 DVSS.n3679 DVSS.n1685 0.00962857
R18212 DVSS.n3679 DVSS.n3678 0.00962857
R18213 DVSS.n3683 DVSS.n3678 0.00962857
R18214 DVSS.n3683 DVSS.n3675 0.00962857
R18215 DVSS.n3687 DVSS.n3675 0.00962857
R18216 DVSS.n3687 DVSS.n3673 0.00962857
R18217 DVSS.n3691 DVSS.n3673 0.00962857
R18218 DVSS.n3691 DVSS.n3671 0.00962857
R18219 DVSS.n3695 DVSS.n3671 0.00962857
R18220 DVSS.n3695 DVSS.n3669 0.00962857
R18221 DVSS.n3699 DVSS.n3669 0.00962857
R18222 DVSS.n3699 DVSS.n3667 0.00962857
R18223 DVSS.n3703 DVSS.n3667 0.00962857
R18224 DVSS.n3703 DVSS.n3665 0.00962857
R18225 DVSS.n3707 DVSS.n3665 0.00962857
R18226 DVSS.n3707 DVSS.n3663 0.00962857
R18227 DVSS.n3711 DVSS.n3663 0.00962857
R18228 DVSS.n3711 DVSS.n3661 0.00962857
R18229 DVSS.n3715 DVSS.n3661 0.00962857
R18230 DVSS.n3715 DVSS.n3659 0.00962857
R18231 DVSS.n3719 DVSS.n3659 0.00962857
R18232 DVSS.n3719 DVSS.n3656 0.00962857
R18233 DVSS.n3742 DVSS.n3656 0.00962857
R18234 DVSS.n3742 DVSS.n3657 0.00962857
R18235 DVSS.n3738 DVSS.n3657 0.00962857
R18236 DVSS.n3738 DVSS.n3723 0.00962857
R18237 DVSS.n3734 DVSS.n3723 0.00962857
R18238 DVSS.n3734 DVSS.n3725 0.00962857
R18239 DVSS.n3730 DVSS.n3725 0.00962857
R18240 DVSS.n2226 DVSS.n2225 0.00962857
R18241 DVSS.n2225 DVSS.n1736 0.00962857
R18242 DVSS.n2221 DVSS.n1736 0.00962857
R18243 DVSS.n2221 DVSS.n1738 0.00962857
R18244 DVSS.n2217 DVSS.n1738 0.00962857
R18245 DVSS.n2217 DVSS.n1741 0.00962857
R18246 DVSS.n2213 DVSS.n1741 0.00962857
R18247 DVSS.n2213 DVSS.n1743 0.00962857
R18248 DVSS.n1894 DVSS.n1743 0.00962857
R18249 DVSS.n1897 DVSS.n1894 0.00962857
R18250 DVSS.n1897 DVSS.n1887 0.00962857
R18251 DVSS.n1903 DVSS.n1887 0.00962857
R18252 DVSS.n1903 DVSS.n1885 0.00962857
R18253 DVSS.n1907 DVSS.n1885 0.00962857
R18254 DVSS.n1907 DVSS.n1764 0.00962857
R18255 DVSS.n2194 DVSS.n1764 0.00962857
R18256 DVSS.n2194 DVSS.n1765 0.00962857
R18257 DVSS.n2190 DVSS.n1765 0.00962857
R18258 DVSS.n2190 DVSS.n1768 0.00962857
R18259 DVSS.n1872 DVSS.n1768 0.00962857
R18260 DVSS.n1872 DVSS.n1791 0.00962857
R18261 DVSS.n2176 DVSS.n1791 0.00962857
R18262 DVSS.n2176 DVSS.n1792 0.00962857
R18263 DVSS.n2172 DVSS.n1792 0.00962857
R18264 DVSS.n2172 DVSS.n1795 0.00962857
R18265 DVSS.n2143 DVSS.n1795 0.00962857
R18266 DVSS.n2143 DVSS.n1927 0.00962857
R18267 DVSS.n2139 DVSS.n1927 0.00962857
R18268 DVSS.n2139 DVSS.n1929 0.00962857
R18269 DVSS.n1968 DVSS.n1929 0.00962857
R18270 DVSS.n1968 DVSS.n1967 0.00962857
R18271 DVSS.n1972 DVSS.n1967 0.00962857
R18272 DVSS.n1972 DVSS.n1957 0.00962857
R18273 DVSS.n1986 DVSS.n1957 0.00962857
R18274 DVSS.n1986 DVSS.n1954 0.00962857
R18275 DVSS.n2122 DVSS.n1954 0.00962857
R18276 DVSS.n2122 DVSS.n1955 0.00962857
R18277 DVSS.n2118 DVSS.n1955 0.00962857
R18278 DVSS.n2118 DVSS.n2083 0.00962857
R18279 DVSS.n2083 DVSS.n2082 0.00962857
R18280 DVSS.n2082 DVSS.n1990 0.00962857
R18281 DVSS.n2078 DVSS.n1990 0.00962857
R18282 DVSS.n2078 DVSS.n1993 0.00962857
R18283 DVSS.n2074 DVSS.n1993 0.00962857
R18284 DVSS.n2074 DVSS.n1996 0.00962857
R18285 DVSS.n2070 DVSS.n1996 0.00962857
R18286 DVSS.n2070 DVSS.n1998 0.00962857
R18287 DVSS.n2066 DVSS.n1998 0.00962857
R18288 DVSS.n2066 DVSS.n2000 0.00962857
R18289 DVSS.n2062 DVSS.n2000 0.00962857
R18290 DVSS.n2062 DVSS.n2002 0.00962857
R18291 DVSS.n2058 DVSS.n2002 0.00962857
R18292 DVSS.n2058 DVSS.n2004 0.00962857
R18293 DVSS.n2054 DVSS.n2004 0.00962857
R18294 DVSS.n2054 DVSS.n2006 0.00962857
R18295 DVSS.n2050 DVSS.n2006 0.00962857
R18296 DVSS.n2050 DVSS.n2008 0.00962857
R18297 DVSS.n2046 DVSS.n2008 0.00962857
R18298 DVSS.n2046 DVSS.n2010 0.00962857
R18299 DVSS.n2042 DVSS.n2010 0.00962857
R18300 DVSS.n2042 DVSS.n2012 0.00962857
R18301 DVSS.n2038 DVSS.n2012 0.00962857
R18302 DVSS.n2038 DVSS.n2014 0.00962857
R18303 DVSS.n2034 DVSS.n2014 0.00962857
R18304 DVSS.n2034 DVSS.n2016 0.00962857
R18305 DVSS.n2030 DVSS.n2016 0.00962857
R18306 DVSS.n2030 DVSS.n2018 0.00962857
R18307 DVSS.n2026 DVSS.n2018 0.00962857
R18308 DVSS.n2026 DVSS.n2020 0.00962857
R18309 DVSS.n4181 DVSS.n4180 0.00962857
R18310 DVSS.n4180 DVSS.n1371 0.00962857
R18311 DVSS.n4176 DVSS.n1371 0.00962857
R18312 DVSS.n4176 DVSS.n1374 0.00962857
R18313 DVSS.n4172 DVSS.n1374 0.00962857
R18314 DVSS.n4172 DVSS.n1377 0.00962857
R18315 DVSS.n4166 DVSS.n1377 0.00962857
R18316 DVSS.n4166 DVSS.n1392 0.00962857
R18317 DVSS.n4162 DVSS.n1392 0.00962857
R18318 DVSS.n4162 DVSS.n1394 0.00962857
R18319 DVSS.n4158 DVSS.n1394 0.00962857
R18320 DVSS.n4158 DVSS.n1396 0.00962857
R18321 DVSS.n4154 DVSS.n1396 0.00962857
R18322 DVSS.n4154 DVSS.n1398 0.00962857
R18323 DVSS.n4150 DVSS.n1398 0.00962857
R18324 DVSS.n4150 DVSS.n1400 0.00962857
R18325 DVSS.n4146 DVSS.n1400 0.00962857
R18326 DVSS.n4146 DVSS.n1402 0.00962857
R18327 DVSS.n4142 DVSS.n1402 0.00962857
R18328 DVSS.n4142 DVSS.n1404 0.00962857
R18329 DVSS.n4138 DVSS.n1404 0.00962857
R18330 DVSS.n4138 DVSS.n1406 0.00962857
R18331 DVSS.n4134 DVSS.n1406 0.00962857
R18332 DVSS.n4134 DVSS.n1408 0.00962857
R18333 DVSS.n4130 DVSS.n1408 0.00962857
R18334 DVSS.n4130 DVSS.n1410 0.00962857
R18335 DVSS.n4126 DVSS.n1410 0.00962857
R18336 DVSS.n4126 DVSS.n1412 0.00962857
R18337 DVSS.n4122 DVSS.n1412 0.00962857
R18338 DVSS.n4122 DVSS.n1414 0.00962857
R18339 DVSS.n4118 DVSS.n1414 0.00962857
R18340 DVSS.n4118 DVSS.n1416 0.00962857
R18341 DVSS.n4114 DVSS.n1416 0.00962857
R18342 DVSS.n4114 DVSS.n1418 0.00962857
R18343 DVSS.n4110 DVSS.n1418 0.00962857
R18344 DVSS.n4110 DVSS.n1420 0.00962857
R18345 DVSS.n4106 DVSS.n1420 0.00962857
R18346 DVSS.n4106 DVSS.n1422 0.00962857
R18347 DVSS.n4102 DVSS.n1422 0.00962857
R18348 DVSS.n4102 DVSS.n1424 0.00962857
R18349 DVSS.n4098 DVSS.n1424 0.00962857
R18350 DVSS.n4098 DVSS.n1426 0.00962857
R18351 DVSS.n4008 DVSS.n1426 0.00962857
R18352 DVSS.n4008 DVSS.n4006 0.00962857
R18353 DVSS.n4091 DVSS.n4006 0.00962857
R18354 DVSS.n4091 DVSS.n4007 0.00962857
R18355 DVSS.n4087 DVSS.n4007 0.00962857
R18356 DVSS.n4087 DVSS.n4012 0.00962857
R18357 DVSS.n4083 DVSS.n4012 0.00962857
R18358 DVSS.n4083 DVSS.n4014 0.00962857
R18359 DVSS.n4079 DVSS.n4014 0.00962857
R18360 DVSS.n4079 DVSS.n4016 0.00962857
R18361 DVSS.n4075 DVSS.n4016 0.00962857
R18362 DVSS.n4075 DVSS.n4018 0.00962857
R18363 DVSS.n4071 DVSS.n4018 0.00962857
R18364 DVSS.n4071 DVSS.n4020 0.00962857
R18365 DVSS.n4067 DVSS.n4020 0.00962857
R18366 DVSS.n4067 DVSS.n4022 0.00962857
R18367 DVSS.n4063 DVSS.n4022 0.00962857
R18368 DVSS.n4063 DVSS.n4024 0.00962857
R18369 DVSS.n4059 DVSS.n4024 0.00962857
R18370 DVSS.n4059 DVSS.n4026 0.00962857
R18371 DVSS.n4055 DVSS.n4026 0.00962857
R18372 DVSS.n4055 DVSS.n4028 0.00962857
R18373 DVSS.n4051 DVSS.n4028 0.00962857
R18374 DVSS.n4051 DVSS.n4030 0.00962857
R18375 DVSS.n4047 DVSS.n4030 0.00962857
R18376 DVSS.n4047 DVSS.n4032 0.00962857
R18377 DVSS.n4043 DVSS.n4032 0.00962857
R18378 DVSS.n4043 DVSS.n4034 0.00962857
R18379 DVSS.n4039 DVSS.n4034 0.00962857
R18380 DVSS.n4179 DVSS.n4178 0.00962857
R18381 DVSS.n4178 DVSS.n4177 0.00962857
R18382 DVSS.n4177 DVSS.n1373 0.00962857
R18383 DVSS.n4167 DVSS.n1391 0.00962857
R18384 DVSS.n4161 DVSS.n1391 0.00962857
R18385 DVSS.n4161 DVSS.n4160 0.00962857
R18386 DVSS.n4160 DVSS.n4159 0.00962857
R18387 DVSS.n4159 DVSS.n1395 0.00962857
R18388 DVSS.n4153 DVSS.n1395 0.00962857
R18389 DVSS.n4153 DVSS.n4152 0.00962857
R18390 DVSS.n4152 DVSS.n4151 0.00962857
R18391 DVSS.n4151 DVSS.n1399 0.00962857
R18392 DVSS.n4145 DVSS.n1399 0.00962857
R18393 DVSS.n4145 DVSS.n4144 0.00962857
R18394 DVSS.n4144 DVSS.n4143 0.00962857
R18395 DVSS.n4143 DVSS.n1403 0.00962857
R18396 DVSS.n4137 DVSS.n1403 0.00962857
R18397 DVSS.n4137 DVSS.n4136 0.00962857
R18398 DVSS.n4136 DVSS.n4135 0.00962857
R18399 DVSS.n4135 DVSS.n1407 0.00962857
R18400 DVSS.n4129 DVSS.n1407 0.00962857
R18401 DVSS.n4129 DVSS.n4128 0.00962857
R18402 DVSS.n4128 DVSS.n4127 0.00962857
R18403 DVSS.n4127 DVSS.n1411 0.00962857
R18404 DVSS.n4121 DVSS.n1411 0.00962857
R18405 DVSS.n4121 DVSS.n4120 0.00962857
R18406 DVSS.n4120 DVSS.n4119 0.00962857
R18407 DVSS.n4119 DVSS.n1415 0.00962857
R18408 DVSS.n4113 DVSS.n1415 0.00962857
R18409 DVSS.n4113 DVSS.n4112 0.00962857
R18410 DVSS.n4112 DVSS.n4111 0.00962857
R18411 DVSS.n4111 DVSS.n1419 0.00962857
R18412 DVSS.n4105 DVSS.n1419 0.00962857
R18413 DVSS.n4105 DVSS.n4104 0.00962857
R18414 DVSS.n4104 DVSS.n4103 0.00962857
R18415 DVSS.n4103 DVSS.n1423 0.00962857
R18416 DVSS.n4097 DVSS.n1423 0.00962857
R18417 DVSS.n4097 DVSS.n4096 0.00962857
R18418 DVSS.n4092 DVSS.n4005 0.00962857
R18419 DVSS.n4086 DVSS.n4005 0.00962857
R18420 DVSS.n4086 DVSS.n4085 0.00962857
R18421 DVSS.n4085 DVSS.n4084 0.00962857
R18422 DVSS.n4084 DVSS.n4013 0.00962857
R18423 DVSS.n4078 DVSS.n4013 0.00962857
R18424 DVSS.n4078 DVSS.n4077 0.00962857
R18425 DVSS.n4077 DVSS.n4076 0.00962857
R18426 DVSS.n4076 DVSS.n4017 0.00962857
R18427 DVSS.n4070 DVSS.n4017 0.00962857
R18428 DVSS.n4070 DVSS.n4069 0.00962857
R18429 DVSS.n4069 DVSS.n4068 0.00962857
R18430 DVSS.n4068 DVSS.n4021 0.00962857
R18431 DVSS.n4062 DVSS.n4021 0.00962857
R18432 DVSS.n4062 DVSS.n4061 0.00962857
R18433 DVSS.n4061 DVSS.n4060 0.00962857
R18434 DVSS.n4060 DVSS.n4025 0.00962857
R18435 DVSS.n4054 DVSS.n4025 0.00962857
R18436 DVSS.n4054 DVSS.n4053 0.00962857
R18437 DVSS.n4053 DVSS.n4052 0.00962857
R18438 DVSS.n4052 DVSS.n4029 0.00962857
R18439 DVSS.n4046 DVSS.n4029 0.00962857
R18440 DVSS.n4046 DVSS.n4045 0.00962857
R18441 DVSS.n4045 DVSS.n4044 0.00962857
R18442 DVSS.n4044 DVSS.n4033 0.00962857
R18443 DVSS.n4038 DVSS.n4033 0.00962857
R18444 DVSS.n2227 DVSS.n1735 0.00962857
R18445 DVSS.n2220 DVSS.n1739 0.00962857
R18446 DVSS.n2220 DVSS.n2219 0.00962857
R18447 DVSS.n2219 DVSS.n2218 0.00962857
R18448 DVSS.n2177 DVSS.n1790 0.00962857
R18449 DVSS.n2171 DVSS.n1790 0.00962857
R18450 DVSS.n2081 DVSS.n2080 0.00962857
R18451 DVSS.n2080 DVSS.n2079 0.00962857
R18452 DVSS.n2079 DVSS.n1992 0.00962857
R18453 DVSS.n2073 DVSS.n1992 0.00962857
R18454 DVSS.n2073 DVSS.n2072 0.00962857
R18455 DVSS.n2072 DVSS.n2071 0.00962857
R18456 DVSS.n2071 DVSS.n1997 0.00962857
R18457 DVSS.n2065 DVSS.n1997 0.00962857
R18458 DVSS.n2065 DVSS.n2064 0.00962857
R18459 DVSS.n2064 DVSS.n2063 0.00962857
R18460 DVSS.n2063 DVSS.n2001 0.00962857
R18461 DVSS.n2057 DVSS.n2001 0.00962857
R18462 DVSS.n2057 DVSS.n2056 0.00962857
R18463 DVSS.n2056 DVSS.n2055 0.00962857
R18464 DVSS.n2055 DVSS.n2005 0.00962857
R18465 DVSS.n2049 DVSS.n2005 0.00962857
R18466 DVSS.n2049 DVSS.n2048 0.00962857
R18467 DVSS.n2048 DVSS.n2047 0.00962857
R18468 DVSS.n2047 DVSS.n2009 0.00962857
R18469 DVSS.n2041 DVSS.n2009 0.00962857
R18470 DVSS.n2041 DVSS.n2040 0.00962857
R18471 DVSS.n2040 DVSS.n2039 0.00962857
R18472 DVSS.n2039 DVSS.n2013 0.00962857
R18473 DVSS.n2033 DVSS.n2013 0.00962857
R18474 DVSS.n2033 DVSS.n2032 0.00962857
R18475 DVSS.n2032 DVSS.n2031 0.00962857
R18476 DVSS.n2031 DVSS.n2017 0.00962857
R18477 DVSS.n2025 DVSS.n2017 0.00962857
R18478 DVSS.n2025 DVSS.n2024 0.00962857
R18479 DVSS.n1595 DVSS.n1590 0.00962857
R18480 DVSS.n3893 DVSS.n1591 0.00962857
R18481 DVSS.n3887 DVSS.n1591 0.00962857
R18482 DVSS.n3885 DVSS.n3884 0.00962857
R18483 DVSS.n3884 DVSS.n1601 0.00962857
R18484 DVSS.n3878 DVSS.n1601 0.00962857
R18485 DVSS.n3868 DVSS.n1609 0.00962857
R18486 DVSS.n3868 DVSS.n3867 0.00962857
R18487 DVSS.n3867 DVSS.n3866 0.00962857
R18488 DVSS.n3860 DVSS.n1614 0.00962857
R18489 DVSS.n3860 DVSS.n3859 0.00962857
R18490 DVSS.n3849 DVSS.n1619 0.00962857
R18491 DVSS.n3849 DVSS.n3848 0.00962857
R18492 DVSS.n3848 DVSS.n3847 0.00962857
R18493 DVSS.n3828 DVSS.n3827 0.00962857
R18494 DVSS.n3827 DVSS.n1633 0.00962857
R18495 DVSS.n1638 DVSS.n1633 0.00962857
R18496 DVSS.n3820 DVSS.n1638 0.00962857
R18497 DVSS.n3820 DVSS.n3819 0.00962857
R18498 DVSS.n3819 DVSS.n3818 0.00962857
R18499 DVSS.n3818 DVSS.n1639 0.00962857
R18500 DVSS.n3812 DVSS.n1639 0.00962857
R18501 DVSS.n3812 DVSS.n3811 0.00962857
R18502 DVSS.n3811 DVSS.n3810 0.00962857
R18503 DVSS.n3810 DVSS.n1643 0.00962857
R18504 DVSS.n3804 DVSS.n3803 0.00962857
R18505 DVSS.n3801 DVSS.n1649 0.00962857
R18506 DVSS.n3795 DVSS.n1649 0.00962857
R18507 DVSS.n1669 DVSS.n1653 0.00962857
R18508 DVSS.n1670 DVSS.n1669 0.00962857
R18509 DVSS.n1675 DVSS.n1670 0.00962857
R18510 DVSS.n3780 DVSS.n1681 0.00962857
R18511 DVSS.n3780 DVSS.n3779 0.00962857
R18512 DVSS.n3779 DVSS.n3778 0.00962857
R18513 DVSS.n3772 DVSS.n1686 0.00962857
R18514 DVSS.n3772 DVSS.n3771 0.00962857
R18515 DVSS.n3684 DVSS.n3677 0.00962857
R18516 DVSS.n3685 DVSS.n3684 0.00962857
R18517 DVSS.n3686 DVSS.n3685 0.00962857
R18518 DVSS.n3686 DVSS.n3672 0.00962857
R18519 DVSS.n3692 DVSS.n3672 0.00962857
R18520 DVSS.n3693 DVSS.n3692 0.00962857
R18521 DVSS.n3694 DVSS.n3693 0.00962857
R18522 DVSS.n3694 DVSS.n3668 0.00962857
R18523 DVSS.n3700 DVSS.n3668 0.00962857
R18524 DVSS.n3701 DVSS.n3700 0.00962857
R18525 DVSS.n3702 DVSS.n3701 0.00962857
R18526 DVSS.n3702 DVSS.n3664 0.00962857
R18527 DVSS.n3708 DVSS.n3664 0.00962857
R18528 DVSS.n3709 DVSS.n3708 0.00962857
R18529 DVSS.n3710 DVSS.n3709 0.00962857
R18530 DVSS.n3710 DVSS.n3660 0.00962857
R18531 DVSS.n3716 DVSS.n3660 0.00962857
R18532 DVSS.n3717 DVSS.n3716 0.00962857
R18533 DVSS.n3718 DVSS.n3717 0.00962857
R18534 DVSS.n3718 DVSS.n3654 0.00962857
R18535 DVSS.n3743 DVSS.n3655 0.00962857
R18536 DVSS.n3737 DVSS.n3655 0.00962857
R18537 DVSS.n3737 DVSS.n3736 0.00962857
R18538 DVSS.n3736 DVSS.n3735 0.00962857
R18539 DVSS.n3735 DVSS.n3724 0.00962857
R18540 DVSS.n3729 DVSS.n3724 0.00962857
R18541 DVSS.n5106 DVSS.n5105 0.00962857
R18542 DVSS.n5105 DVSS.n1084 0.00962857
R18543 DVSS.n5101 DVSS.n1084 0.00962857
R18544 DVSS.n5101 DVSS.n1086 0.00962857
R18545 DVSS.n5097 DVSS.n1086 0.00962857
R18546 DVSS.n5097 DVSS.n1089 0.00962857
R18547 DVSS.n5093 DVSS.n1089 0.00962857
R18548 DVSS.n5093 DVSS.n1091 0.00962857
R18549 DVSS.n5089 DVSS.n1091 0.00962857
R18550 DVSS.n5089 DVSS.n1093 0.00962857
R18551 DVSS.n5085 DVSS.n1093 0.00962857
R18552 DVSS.n5085 DVSS.n1095 0.00962857
R18553 DVSS.n5081 DVSS.n1095 0.00962857
R18554 DVSS.n5081 DVSS.n1097 0.00962857
R18555 DVSS.n5077 DVSS.n1097 0.00962857
R18556 DVSS.n5077 DVSS.n1099 0.00962857
R18557 DVSS.n5072 DVSS.n1099 0.00962857
R18558 DVSS.n5072 DVSS.n1103 0.00962857
R18559 DVSS.n5068 DVSS.n1103 0.00962857
R18560 DVSS.n5068 DVSS.n1105 0.00962857
R18561 DVSS.n5064 DVSS.n1105 0.00962857
R18562 DVSS.n5064 DVSS.n1107 0.00962857
R18563 DVSS.n5060 DVSS.n1107 0.00962857
R18564 DVSS.n5060 DVSS.n1109 0.00962857
R18565 DVSS.n5053 DVSS.n1109 0.00962857
R18566 DVSS.n5053 DVSS.n1114 0.00962857
R18567 DVSS.n5049 DVSS.n1114 0.00962857
R18568 DVSS.n5049 DVSS.n1116 0.00962857
R18569 DVSS.n5042 DVSS.n1116 0.00962857
R18570 DVSS.n5042 DVSS.n1122 0.00962857
R18571 DVSS.n5038 DVSS.n1122 0.00962857
R18572 DVSS.n5038 DVSS.n1124 0.00962857
R18573 DVSS.n5034 DVSS.n1124 0.00962857
R18574 DVSS.n5034 DVSS.n1127 0.00962857
R18575 DVSS.n5030 DVSS.n1127 0.00962857
R18576 DVSS.n5030 DVSS.n1129 0.00962857
R18577 DVSS.n5026 DVSS.n1129 0.00962857
R18578 DVSS.n5026 DVSS.n1131 0.00962857
R18579 DVSS.n5022 DVSS.n1131 0.00962857
R18580 DVSS.n5022 DVSS.n1133 0.00962857
R18581 DVSS.n5018 DVSS.n1133 0.00962857
R18582 DVSS.n5018 DVSS.n1135 0.00962857
R18583 DVSS.n5014 DVSS.n1135 0.00962857
R18584 DVSS.n5014 DVSS.n1137 0.00962857
R18585 DVSS.n5010 DVSS.n1137 0.00962857
R18586 DVSS.n5010 DVSS.n1139 0.00962857
R18587 DVSS.n5006 DVSS.n1139 0.00962857
R18588 DVSS.n5006 DVSS.n1141 0.00962857
R18589 DVSS.n5002 DVSS.n1141 0.00962857
R18590 DVSS.n5002 DVSS.n1143 0.00962857
R18591 DVSS.n4998 DVSS.n1143 0.00962857
R18592 DVSS.n4998 DVSS.n1145 0.00962857
R18593 DVSS.n4994 DVSS.n1145 0.00962857
R18594 DVSS.n4994 DVSS.n1147 0.00962857
R18595 DVSS.n4990 DVSS.n1147 0.00962857
R18596 DVSS.n4990 DVSS.n1149 0.00962857
R18597 DVSS.n4986 DVSS.n1149 0.00962857
R18598 DVSS.n4986 DVSS.n1151 0.00962857
R18599 DVSS.n4982 DVSS.n1151 0.00962857
R18600 DVSS.n4982 DVSS.n1153 0.00962857
R18601 DVSS.n2319 DVSS.n1153 0.00962857
R18602 DVSS.n2322 DVSS.n2319 0.00962857
R18603 DVSS.n2322 DVSS.n2318 0.00962857
R18604 DVSS.n2326 DVSS.n2318 0.00962857
R18605 DVSS.n2326 DVSS.n2316 0.00962857
R18606 DVSS.n2330 DVSS.n2316 0.00962857
R18607 DVSS.n2330 DVSS.n2314 0.00962857
R18608 DVSS.n2334 DVSS.n2314 0.00962857
R18609 DVSS.n2334 DVSS.n2312 0.00962857
R18610 DVSS.n2338 DVSS.n2312 0.00962857
R18611 DVSS.n2338 DVSS.n2310 0.00962857
R18612 DVSS.n2342 DVSS.n2310 0.00962857
R18613 DVSS.n2342 DVSS.n2308 0.00962857
R18614 DVSS.n2346 DVSS.n2308 0.00962857
R18615 DVSS.n2346 DVSS.n2306 0.00962857
R18616 DVSS.n2350 DVSS.n2306 0.00962857
R18617 DVSS.n2350 DVSS.n2304 0.00962857
R18618 DVSS.n2354 DVSS.n2304 0.00962857
R18619 DVSS.n2354 DVSS.n2302 0.00962857
R18620 DVSS.n2358 DVSS.n2302 0.00962857
R18621 DVSS.n2358 DVSS.n2300 0.00962857
R18622 DVSS.n2362 DVSS.n2300 0.00962857
R18623 DVSS.n2362 DVSS.n2298 0.00962857
R18624 DVSS.n2366 DVSS.n2298 0.00962857
R18625 DVSS.n2366 DVSS.n2296 0.00962857
R18626 DVSS.n2370 DVSS.n2296 0.00962857
R18627 DVSS.n2370 DVSS.n2294 0.00962857
R18628 DVSS.n2374 DVSS.n2294 0.00962857
R18629 DVSS.n2374 DVSS.n2292 0.00962857
R18630 DVSS.n2378 DVSS.n2292 0.00962857
R18631 DVSS.n2378 DVSS.n2290 0.00962857
R18632 DVSS.n2382 DVSS.n2290 0.00962857
R18633 DVSS.n2382 DVSS.n2288 0.00962857
R18634 DVSS.n2387 DVSS.n2288 0.00962857
R18635 DVSS.n2387 DVSS.n2286 0.00962857
R18636 DVSS.n2391 DVSS.n2286 0.00962857
R18637 DVSS.n2393 DVSS.n2391 0.00962857
R18638 DVSS.n2402 DVSS.n2283 0.00962857
R18639 DVSS.n2402 DVSS.n2284 0.00962857
R18640 DVSS.n2398 DVSS.n2284 0.00962857
R18641 DVSS.n5108 DVSS.n5107 0.00962857
R18642 DVSS.n5107 DVSS.n1083 0.00962857
R18643 DVSS.n1087 DVSS.n1083 0.00962857
R18644 DVSS.n5100 DVSS.n1087 0.00962857
R18645 DVSS.n5100 DVSS.n5099 0.00962857
R18646 DVSS.n5099 DVSS.n5098 0.00962857
R18647 DVSS.n5098 DVSS.n1088 0.00962857
R18648 DVSS.n5092 DVSS.n1088 0.00962857
R18649 DVSS.n5092 DVSS.n5091 0.00962857
R18650 DVSS.n5091 DVSS.n5090 0.00962857
R18651 DVSS.n5090 DVSS.n1092 0.00962857
R18652 DVSS.n5084 DVSS.n1092 0.00962857
R18653 DVSS.n5084 DVSS.n5083 0.00962857
R18654 DVSS.n5083 DVSS.n5082 0.00962857
R18655 DVSS.n5082 DVSS.n1096 0.00962857
R18656 DVSS.n5074 DVSS.n5073 0.00962857
R18657 DVSS.n5073 DVSS.n1102 0.00962857
R18658 DVSS.n5067 DVSS.n1102 0.00962857
R18659 DVSS.n5067 DVSS.n5066 0.00962857
R18660 DVSS.n5066 DVSS.n5065 0.00962857
R18661 DVSS.n5065 DVSS.n1106 0.00962857
R18662 DVSS.n5037 DVSS.n1125 0.00962857
R18663 DVSS.n5037 DVSS.n5036 0.00962857
R18664 DVSS.n5036 DVSS.n5035 0.00962857
R18665 DVSS.n5035 DVSS.n1126 0.00962857
R18666 DVSS.n5029 DVSS.n1126 0.00962857
R18667 DVSS.n5029 DVSS.n5028 0.00962857
R18668 DVSS.n5028 DVSS.n5027 0.00962857
R18669 DVSS.n5027 DVSS.n1130 0.00962857
R18670 DVSS.n5021 DVSS.n1130 0.00962857
R18671 DVSS.n5021 DVSS.n5020 0.00962857
R18672 DVSS.n5020 DVSS.n5019 0.00962857
R18673 DVSS.n5019 DVSS.n1134 0.00962857
R18674 DVSS.n5013 DVSS.n1134 0.00962857
R18675 DVSS.n5013 DVSS.n5012 0.00962857
R18676 DVSS.n5012 DVSS.n5011 0.00962857
R18677 DVSS.n5011 DVSS.n1138 0.00962857
R18678 DVSS.n5005 DVSS.n1138 0.00962857
R18679 DVSS.n5005 DVSS.n5004 0.00962857
R18680 DVSS.n5004 DVSS.n5003 0.00962857
R18681 DVSS.n5003 DVSS.n1142 0.00962857
R18682 DVSS.n4997 DVSS.n1142 0.00962857
R18683 DVSS.n4997 DVSS.n4996 0.00962857
R18684 DVSS.n4996 DVSS.n4995 0.00962857
R18685 DVSS.n4995 DVSS.n1146 0.00962857
R18686 DVSS.n4989 DVSS.n1146 0.00962857
R18687 DVSS.n4989 DVSS.n4988 0.00962857
R18688 DVSS.n4988 DVSS.n4987 0.00962857
R18689 DVSS.n4987 DVSS.n1150 0.00962857
R18690 DVSS.n4981 DVSS.n1150 0.00962857
R18691 DVSS.n4981 DVSS.n4980 0.00962857
R18692 DVSS.n2323 DVSS.n1154 0.00962857
R18693 DVSS.n2324 DVSS.n2323 0.00962857
R18694 DVSS.n2325 DVSS.n2324 0.00962857
R18695 DVSS.n2325 DVSS.n2315 0.00962857
R18696 DVSS.n2331 DVSS.n2315 0.00962857
R18697 DVSS.n2332 DVSS.n2331 0.00962857
R18698 DVSS.n2333 DVSS.n2332 0.00962857
R18699 DVSS.n2333 DVSS.n2311 0.00962857
R18700 DVSS.n2339 DVSS.n2311 0.00962857
R18701 DVSS.n2340 DVSS.n2339 0.00962857
R18702 DVSS.n2341 DVSS.n2340 0.00962857
R18703 DVSS.n2341 DVSS.n2307 0.00962857
R18704 DVSS.n2347 DVSS.n2307 0.00962857
R18705 DVSS.n2348 DVSS.n2347 0.00962857
R18706 DVSS.n2349 DVSS.n2348 0.00962857
R18707 DVSS.n2349 DVSS.n2303 0.00962857
R18708 DVSS.n2355 DVSS.n2303 0.00962857
R18709 DVSS.n2356 DVSS.n2355 0.00962857
R18710 DVSS.n2357 DVSS.n2356 0.00962857
R18711 DVSS.n2357 DVSS.n2299 0.00962857
R18712 DVSS.n2363 DVSS.n2299 0.00962857
R18713 DVSS.n2364 DVSS.n2363 0.00962857
R18714 DVSS.n2365 DVSS.n2364 0.00962857
R18715 DVSS.n2365 DVSS.n2295 0.00962857
R18716 DVSS.n2371 DVSS.n2295 0.00962857
R18717 DVSS.n2372 DVSS.n2371 0.00962857
R18718 DVSS.n2373 DVSS.n2372 0.00962857
R18719 DVSS.n2373 DVSS.n2291 0.00962857
R18720 DVSS.n2379 DVSS.n2291 0.00962857
R18721 DVSS.n2380 DVSS.n2379 0.00962857
R18722 DVSS.n2381 DVSS.n2380 0.00962857
R18723 DVSS.n2381 DVSS.n2287 0.00962857
R18724 DVSS.n2388 DVSS.n2287 0.00962857
R18725 DVSS.n2389 DVSS.n2388 0.00962857
R18726 DVSS.n2390 DVSS.n2389 0.00962857
R18727 DVSS.n2403 DVSS.n2282 0.00962857
R18728 DVSS.n2397 DVSS.n2282 0.00962857
R18729 DVSS.n2397 DVSS.n2396 0.00962857
R18730 DVSS.n1537 DVSS.n1534 0.00962857
R18731 DVSS.n1538 DVSS.n1537 0.00962857
R18732 DVSS.n1539 DVSS.n1538 0.00962857
R18733 DVSS.n1539 DVSS.n1530 0.00962857
R18734 DVSS.n1545 DVSS.n1530 0.00962857
R18735 DVSS.n1546 DVSS.n1545 0.00962857
R18736 DVSS.n1547 DVSS.n1546 0.00962857
R18737 DVSS.n1547 DVSS.n1526 0.00962857
R18738 DVSS.n1553 DVSS.n1526 0.00962857
R18739 DVSS.n1554 DVSS.n1553 0.00962857
R18740 DVSS.n1555 DVSS.n1554 0.00962857
R18741 DVSS.n1555 DVSS.n1520 0.00962857
R18742 DVSS.n3936 DVSS.n1521 0.00962857
R18743 DVSS.n3930 DVSS.n1521 0.00962857
R18744 DVSS.n3930 DVSS.n3929 0.00962857
R18745 DVSS.n3929 DVSS.n3928 0.00962857
R18746 DVSS.n3928 DVSS.n1561 0.00962857
R18747 DVSS.n3922 DVSS.n1561 0.00962857
R18748 DVSS.n3922 DVSS.n3921 0.00962857
R18749 DVSS.n3921 DVSS.n3920 0.00962857
R18750 DVSS.n3920 DVSS.n1565 0.00962857
R18751 DVSS.n3914 DVSS.n1565 0.00962857
R18752 DVSS.n3914 DVSS.n3913 0.00962857
R18753 DVSS.n3913 DVSS.n3912 0.00962857
R18754 DVSS.n3912 DVSS.n1569 0.00962857
R18755 DVSS.n3906 DVSS.n1569 0.00962857
R18756 DVSS.n2493 DVSS.n1573 0.00962857
R18757 DVSS.n2498 DVSS.n2493 0.00962857
R18758 DVSS.n2499 DVSS.n2498 0.00962857
R18759 DVSS.n2500 DVSS.n2499 0.00962857
R18760 DVSS.n2500 DVSS.n2489 0.00962857
R18761 DVSS.n2506 DVSS.n2489 0.00962857
R18762 DVSS.n2507 DVSS.n2506 0.00962857
R18763 DVSS.n2508 DVSS.n2507 0.00962857
R18764 DVSS.n2508 DVSS.n2485 0.00962857
R18765 DVSS.n2514 DVSS.n2485 0.00962857
R18766 DVSS.n2515 DVSS.n2514 0.00962857
R18767 DVSS.n2516 DVSS.n2515 0.00962857
R18768 DVSS.n2516 DVSS.n2481 0.00962857
R18769 DVSS.n2522 DVSS.n2481 0.00962857
R18770 DVSS.n2523 DVSS.n2522 0.00962857
R18771 DVSS.n2524 DVSS.n2523 0.00962857
R18772 DVSS.n2524 DVSS.n2477 0.00962857
R18773 DVSS.n2530 DVSS.n2477 0.00962857
R18774 DVSS.n2531 DVSS.n2530 0.00962857
R18775 DVSS.n2532 DVSS.n2531 0.00962857
R18776 DVSS.n2532 DVSS.n2473 0.00962857
R18777 DVSS.n2538 DVSS.n2473 0.00962857
R18778 DVSS.n2539 DVSS.n2538 0.00962857
R18779 DVSS.n2540 DVSS.n2539 0.00962857
R18780 DVSS.n2540 DVSS.n2469 0.00962857
R18781 DVSS.n2546 DVSS.n2469 0.00962857
R18782 DVSS.n2547 DVSS.n2546 0.00962857
R18783 DVSS.n2548 DVSS.n2547 0.00962857
R18784 DVSS.n2548 DVSS.n2465 0.00962857
R18785 DVSS.n2554 DVSS.n2465 0.00962857
R18786 DVSS.n2555 DVSS.n2554 0.00962857
R18787 DVSS.n2556 DVSS.n2555 0.00962857
R18788 DVSS.n2556 DVSS.n2461 0.00962857
R18789 DVSS.n2562 DVSS.n2461 0.00962857
R18790 DVSS.n2563 DVSS.n2562 0.00962857
R18791 DVSS.n2564 DVSS.n2563 0.00962857
R18792 DVSS.n2564 DVSS.n2457 0.00962857
R18793 DVSS.n2570 DVSS.n2457 0.00962857
R18794 DVSS.n2571 DVSS.n2570 0.00962857
R18795 DVSS.n2572 DVSS.n2571 0.00962857
R18796 DVSS.n2572 DVSS.n2453 0.00962857
R18797 DVSS.n2578 DVSS.n2453 0.00962857
R18798 DVSS.n2579 DVSS.n2578 0.00962857
R18799 DVSS.n2580 DVSS.n2579 0.00962857
R18800 DVSS.n2580 DVSS.n2449 0.00962857
R18801 DVSS.n2586 DVSS.n2449 0.00962857
R18802 DVSS.n2587 DVSS.n2586 0.00962857
R18803 DVSS.n2588 DVSS.n2587 0.00962857
R18804 DVSS.n2588 DVSS.n2445 0.00962857
R18805 DVSS.n2594 DVSS.n2445 0.00962857
R18806 DVSS.n2595 DVSS.n2594 0.00962857
R18807 DVSS.n2596 DVSS.n2595 0.00962857
R18808 DVSS.n2596 DVSS.n2441 0.00962857
R18809 DVSS.n2602 DVSS.n2441 0.00962857
R18810 DVSS.n2603 DVSS.n2602 0.00962857
R18811 DVSS.n2604 DVSS.n2603 0.00962857
R18812 DVSS.n2604 DVSS.n2437 0.00962857
R18813 DVSS.n2610 DVSS.n2437 0.00962857
R18814 DVSS.n2611 DVSS.n2610 0.00962857
R18815 DVSS.n2612 DVSS.n2611 0.00962857
R18816 DVSS.n2612 DVSS.n2433 0.00962857
R18817 DVSS.n2618 DVSS.n2433 0.00962857
R18818 DVSS.n2619 DVSS.n2618 0.00962857
R18819 DVSS.n2620 DVSS.n2619 0.00962857
R18820 DVSS.n2620 DVSS.n2429 0.00962857
R18821 DVSS.n2626 DVSS.n2429 0.00962857
R18822 DVSS.n2627 DVSS.n2626 0.00962857
R18823 DVSS.n2628 DVSS.n2627 0.00962857
R18824 DVSS.n2628 DVSS.n2421 0.00962857
R18825 DVSS.n2650 DVSS.n2649 0.00962857
R18826 DVSS.n2650 DVSS.n2265 0.00962857
R18827 DVSS.n2654 DVSS.n2265 0.00962857
R18828 DVSS.n3240 DVSS 0.00958867
R18829 DVSS.n3365 DVSS 0.00958867
R18830 DVSS.n2131 DVSS.n2130 0.00958257
R18831 DVSS.n2200 DVSS.n1753 0.00958257
R18832 DVSS.n3744 DVSS.n3743 0.00956429
R18833 DVSS.n5727 DVSS.n58 0.0095301
R18834 DVSS.n2211 DVSS.n1745 0.0095
R18835 DVSS.n1893 DVSS.n1892 0.0095
R18836 DVSS.n1899 DVSS.n1898 0.0095
R18837 DVSS.n1891 DVSS.n1888 0.0095
R18838 DVSS.n1902 DVSS.n1901 0.0095
R18839 DVSS.n2197 DVSS.n2195 0.0095
R18840 DVSS.n1769 DVSS.n1763 0.0095
R18841 DVSS.n2189 DVSS.n1770 0.0095
R18842 DVSS.n2188 DVSS.n1771 0.0095
R18843 DVSS.n2179 DVSS.n2177 0.0095
R18844 DVSS.n1930 DVSS.n1926 0.0095
R18845 DVSS.n2138 DVSS.n1931 0.0095
R18846 DVSS.n2137 DVSS.n1932 0.0095
R18847 DVSS.n1963 DVSS.n1962 0.0095
R18848 DVSS.n1985 DVSS.n1983 0.0095
R18849 DVSS.n1984 DVSS.n1952 0.0095
R18850 DVSS.n2124 DVSS.n2123 0.0095
R18851 DVSS.n2084 DVSS.n1953 0.0095
R18852 DVSS.n2117 DVSS.n2085 0.0095
R18853 DVSS.n2843 DVSS.n2769 0.0095
R18854 DVSS.n2887 DVSS.n2760 0.0095
R18855 DVSS.n3449 DVSS.n3448 0.0095
R18856 DVSS.n3437 DVSS.n3221 0.0095
R18857 DVSS.n2829 DVSS.n2777 0.0095
R18858 DVSS.n2884 DVSS.n2762 0.0095
R18859 DVSS.n3348 DVSS.n3200 0.0095
R18860 DVSS.n3357 DVSS.n3218 0.0095
R18861 DVSS.n2861 DVSS.n2759 0.00936699
R18862 DVSS.n2870 DVSS.n2869 0.00936699
R18863 DVSS.n959 DVSS.n957 0.00934354
R18864 DVSS.n5354 DVSS.n959 0.00934354
R18865 DVSS.n4817 DVSS.n4809 0.00933782
R18866 DVSS.n4814 DVSS.n4811 0.00933782
R18867 DVSS.n4814 DVSS.n4809 0.00933782
R18868 DVSS.n4820 DVSS.n4811 0.00933782
R18869 DVSS.n4535 DVSS.n4526 0.00933782
R18870 DVSS.n4529 DVSS.n4526 0.00933782
R18871 DVSS.n4791 DVSS.n4789 0.00928049
R18872 DVSS.n4888 DVSS.n4787 0.00928049
R18873 DVSS.n4758 DVSS.n4757 0.00928049
R18874 DVSS.n4919 DVSS.n4918 0.00928049
R18875 DVSS.n4720 DVSS.n1250 0.00928049
R18876 DVSS.n4732 DVSS.n1242 0.00928049
R18877 DVSS.n4681 DVSS.n1270 0.00928049
R18878 DVSS.n4692 DVSS.n1263 0.00928049
R18879 DVSS.n4598 DVSS.n4596 0.00928049
R18880 DVSS.n4640 DVSS.n4594 0.00928049
R18881 DVSS.n4565 DVSS.n4564 0.00928049
R18882 DVSS.n4671 DVSS.n4670 0.00928049
R18883 DVSS.n5552 DVSS.n855 0.00924286
R18884 DVSS.n5110 DVSS.n1023 0.00910927
R18885 DVSS.n1024 DVSS.n963 0.00910927
R18886 DVSS.n277 DVSS.n276 0.00909873
R18887 DVSS.n2820 DVSS.n2819 0.009
R18888 DVSS.n2911 DVSS.n2910 0.009
R18889 DVSS.n3460 DVSS.n3183 0.009
R18890 DVSS.n3238 DVSS.n3237 0.009
R18891 DVSS.n2823 DVSS.n2822 0.009
R18892 DVSS.n2876 DVSS.n2751 0.009
R18893 DVSS.n3338 DVSS.n3336 0.009
R18894 DVSS.n3368 DVSS.n3367 0.009
R18895 DVSS.n1845 DVSS.n1381 0.00894122
R18896 DVSS.n1845 DVSS.n1387 0.00894122
R18897 DVSS.n1674 DVSS.n1661 0.00892143
R18898 DVSS.n1686 DVSS.n1682 0.00892143
R18899 DVSS.n1100 DVSS.n1096 0.00892143
R18900 DVSS.n5076 DVSS.n5075 0.00892143
R18901 DVSS.n767 DVSS.n57 0.00882776
R18902 DVSS.n4096 DVSS.n4095 0.00879286
R18903 DVSS.n1436 DVSS.n1431 0.00879286
R18904 DVSS.n4093 DVSS.n4004 0.00879286
R18905 DVSS.n3855 DVSS.n1615 0.00879286
R18906 DVSS.n2218 DVSS.n1740 0.0086
R18907 DVSS.n4753 DVSS.n4752 0.00853571
R18908 DVSS.n1231 DVSS.n1228 0.00853571
R18909 DVSS.n4761 DVSS.n4759 0.00853571
R18910 DVSS.n4760 DVSS.n1222 0.00853571
R18911 DVSS.n4917 DVSS.n4916 0.00853571
R18912 DVSS.n4767 DVSS.n1223 0.00853571
R18913 DVSS.n4910 DVSS.n4770 0.00853571
R18914 DVSS.n4171 DVSS.n1378 0.00853571
R18915 DVSS.n4170 DVSS.n1384 0.00853571
R18916 DVSS.n4168 DVSS.n4167 0.00853571
R18917 DVSS.n1647 DVSS.n1643 0.00853571
R18918 DVSS.n3399 DVSS 0.00852817
R18919 DVSS.n3400 DVSS 0.00852817
R18920 DVSS.n2966 DVSS.n2965 0.0085
R18921 DVSS.n3481 DVSS.n3480 0.0085
R18922 DVSS.n2937 DVSS.n2728 0.0085
R18923 DVSS.n3315 DVSS.n3155 0.0085
R18924 DVSS.n4848 DVSS.n1178 0.00847143
R18925 DVSS.n1823 DVSS.n1744 0.00847143
R18926 DVSS.n1110 DVSS.n1106 0.00847143
R18927 DVSS.n5059 DVSS.n5058 0.00847143
R18928 DVSS.n5055 DVSS.n1111 0.00847143
R18929 DVSS.n5054 DVSS.n1113 0.00847143
R18930 DVSS.n1118 DVSS.n1117 0.00847143
R18931 DVSS.n5048 DVSS.n5047 0.00847143
R18932 DVSS.n5044 DVSS.n1119 0.00847143
R18933 DVSS.n5043 DVSS.n1121 0.00847143
R18934 DVSS.n429 DVSS.n241 0.00842994
R18935 DVSS.n2087 DVSS.n1810 0.00834286
R18936 DVSS.n2081 DVSS.n1809 0.00834286
R18937 DVSS.n3877 DVSS.n3876 0.00827857
R18938 DVSS.n1614 DVSS.n1610 0.00827857
R18939 DVSS.n3038 DVSS 0.00825862
R18940 DVSS DVSS.n3044 0.00825862
R18941 DVSS.n3952 DVSS.n1506 0.00823128
R18942 DVSS.n1855 DVSS.n1385 0.00822787
R18943 DVSS.n1837 DVSS.n1379 0.00822787
R18944 DVSS.n1513 DVSS.n1512 0.00821429
R18945 DVSS.n3676 DVSS.n1687 0.00815
R18946 DVSS.n2916 DVSS.n2746 0.00803695
R18947 DVSS.n2871 DVSS.n2742 0.00803695
R18948 DVSS.n2812 DVSS.n2790 0.00803521
R18949 DVSS.n2811 DVSS.n2792 0.00803521
R18950 DVSS.n2821 DVSS.n2786 0.00803521
R18951 DVSS.n2837 DVSS.n2781 0.00803521
R18952 DVSS.n2836 DVSS.n2776 0.00803521
R18953 DVSS.n2845 DVSS.n2844 0.00803521
R18954 DVSS.n2856 DVSS.n2770 0.00803521
R18955 DVSS.n2855 DVSS.n2772 0.00803521
R18956 DVSS.n2865 DVSS.n2766 0.00803521
R18957 DVSS.n2886 DVSS.n2761 0.00803521
R18958 DVSS.n2885 DVSS.n2756 0.00803521
R18959 DVSS.n2894 DVSS.n2893 0.00803521
R18960 DVSS.n2909 DVSS.n2750 0.00803521
R18961 DVSS.n2908 DVSS.n2752 0.00803521
R18962 DVSS.n2905 DVSS.n2904 0.00803521
R18963 DVSS.n2920 DVSS.n2744 0.00803521
R18964 DVSS.n2948 DVSS.n2739 0.00803521
R18965 DVSS.n2947 DVSS.n2734 0.00803521
R18966 DVSS.n2957 DVSS.n2956 0.00803521
R18967 DVSS.n2964 DVSS.n2727 0.00803521
R18968 DVSS.n2963 DVSS.n2730 0.00803521
R18969 DVSS.n2729 DVSS.n2721 0.00803521
R18970 DVSS.n2976 DVSS.n2975 0.00803521
R18971 DVSS.n2987 DVSS.n2715 0.00803521
R18972 DVSS.n2986 DVSS.n2717 0.00803521
R18973 DVSS.n2995 DVSS.n2711 0.00803521
R18974 DVSS.n3011 DVSS.n2706 0.00803521
R18975 DVSS.n3010 DVSS.n2701 0.00803521
R18976 DVSS.n3022 DVSS.n3021 0.00803521
R18977 DVSS.n3034 DVSS.n2694 0.00803521
R18978 DVSS.n3033 DVSS.n2697 0.00803521
R18979 DVSS.n3041 DVSS.n2690 0.00803521
R18980 DVSS.n3052 DVSS.n2685 0.00803521
R18981 DVSS.n3051 DVSS.n2680 0.00803521
R18982 DVSS.n3063 DVSS.n3062 0.00803521
R18983 DVSS.n3550 DVSS.n2666 0.00803521
R18984 DVSS.n3254 DVSS.n2667 0.00803521
R18985 DVSS.n3543 DVSS.n2673 0.00803521
R18986 DVSS.n3542 DVSS.n2675 0.00803521
R18987 DVSS.n3539 DVSS.n3538 0.00803521
R18988 DVSS.n3265 DVSS.n3073 0.00803521
R18989 DVSS.n3530 DVSS.n3080 0.00803521
R18990 DVSS.n3529 DVSS.n3082 0.00803521
R18991 DVSS.n3526 DVSS.n3525 0.00803521
R18992 DVSS.n3277 DVSS.n3090 0.00803521
R18993 DVSS.n3518 DVSS.n3100 0.00803521
R18994 DVSS.n3517 DVSS.n3102 0.00803521
R18995 DVSS.n3514 DVSS.n3513 0.00803521
R18996 DVSS.n3288 DVSS.n3110 0.00803521
R18997 DVSS.n3505 DVSS.n3117 0.00803521
R18998 DVSS.n3504 DVSS.n3119 0.00803521
R18999 DVSS.n3501 DVSS.n3500 0.00803521
R19000 DVSS.n3301 DVSS.n3127 0.00803521
R19001 DVSS.n3493 DVSS.n3136 0.00803521
R19002 DVSS.n3492 DVSS.n3138 0.00803521
R19003 DVSS.n3489 DVSS.n3488 0.00803521
R19004 DVSS.n3313 DVSS.n3146 0.00803521
R19005 DVSS.n3479 DVSS.n3154 0.00803521
R19006 DVSS.n3478 DVSS.n3156 0.00803521
R19007 DVSS.n3475 DVSS.n3474 0.00803521
R19008 DVSS.n3324 DVSS.n3164 0.00803521
R19009 DVSS.n3467 DVSS.n3171 0.00803521
R19010 DVSS.n3466 DVSS.n3173 0.00803521
R19011 DVSS.n3463 DVSS.n3462 0.00803521
R19012 DVSS.n3337 DVSS.n3181 0.00803521
R19013 DVSS.n3455 DVSS.n3191 0.00803521
R19014 DVSS.n3454 DVSS.n3193 0.00803521
R19015 DVSS.n3451 DVSS.n3450 0.00803521
R19016 DVSS.n3349 DVSS.n3201 0.00803521
R19017 DVSS.n3443 DVSS.n3209 0.00803521
R19018 DVSS.n3442 DVSS.n3211 0.00803521
R19019 DVSS.n3439 DVSS.n3438 0.00803521
R19020 DVSS.n3361 DVSS.n3219 0.00803521
R19021 DVSS.n3430 DVSS.n3226 0.00803521
R19022 DVSS.n3429 DVSS.n3228 0.00803521
R19023 DVSS.n3426 DVSS.n3425 0.00803521
R19024 DVSS.n3373 DVSS.n3236 0.00803521
R19025 DVSS.n3418 DVSS.n3243 0.00803521
R19026 DVSS.n3014 DVSS.n3012 0.008
R19027 DVSS.n3128 DVSS.n3116 0.008
R19028 DVSS.n3009 DVSS.n3008 0.008
R19029 DVSS.n3295 DVSS.n3294 0.008
R19030 DVSS.n2392 DVSS.n2275 0.00789286
R19031 DVSS.n2419 DVSS.n2403 0.00789286
R19032 DVSS.n2646 DVSS.n2636 0.00789286
R19033 DVSS.n2649 DVSS.n2648 0.00789286
R19034 DVSS.n5548 DVSS 0.00782857
R19035 DVSS.n5547 DVSS 0.00782857
R19036 DVSS.n4858 DVSS 0.00782857
R19037 DVSS.n2635 VSS 0.00782857
R19038 DVSS.n3730 DVSS 0.00782857
R19039 DVSS DVSS.n2020 0.00782857
R19040 DVSS.n4039 DVSS 0.00782857
R19041 DVSS.n4038 DVSS 0.00782857
R19042 DVSS.n2024 DVSS 0.00782857
R19043 DVSS.n3729 DVSS 0.00782857
R19044 DVSS.n2393 VSS 0.00782857
R19045 DVSS.n3802 DVSS.n3801 0.00776429
R19046 DVSS.n4792 DVSS.n4776 0.00761735
R19047 DVSS.n4886 DVSS.n4794 0.00761735
R19048 DVSS.n4755 DVSS.n1218 0.00761735
R19049 DVSS.n4920 DVSS.n1219 0.00761735
R19050 DVSS.n4719 DVSS.n4717 0.00761735
R19051 DVSS.n4734 DVSS.n1241 0.00761735
R19052 DVSS.n4680 DVSS.n1271 0.00761735
R19053 DVSS.n4694 DVSS.n1262 0.00761735
R19054 DVSS.n4599 DVSS.n4583 0.00761735
R19055 DVSS.n4638 DVSS.n4601 0.00761735
R19056 DVSS.n4562 DVSS.n4492 0.00761735
R19057 DVSS.n4672 DVSS.n4493 0.00761735
R19058 DVSS.n3435 DVSS.n3434 0.0075936
R19059 DVSS.n3359 DVSS.n3245 0.0075936
R19060 DVSS.n4653 DVSS.n4652 0.00757143
R19061 DVSS.n4649 DVSS.n4582 0.00757143
R19062 DVSS.n4648 DVSS.n4585 0.00757143
R19063 DVSS.n4592 DVSS.n4591 0.00757143
R19064 DVSS.n4642 DVSS.n4641 0.00757143
R19065 DVSS.n4602 DVSS.n4593 0.00757143
R19066 DVSS.n4636 DVSS.n4603 0.00757143
R19067 DVSS.n1877 DVSS.n1870 0.00757143
R19068 DVSS.n1874 DVSS.n1787 0.00757143
R19069 DVSS.n4620 DVSS.n4614 0.00750714
R19070 DVSS.n4617 DVSS.n4616 0.00750714
R19071 DVSS.n4684 DVSS.n1269 0.00750714
R19072 DVSS.n4683 DVSS.n1264 0.00750714
R19073 DVSS.n4691 DVSS.n4690 0.00750714
R19074 DVSS.n1265 DVSS.n1260 0.00750714
R19075 DVSS.n4697 DVSS.n4696 0.00750714
R19076 DVSS.n4876 DVSS.n4875 0.00750714
R19077 DVSS.n4830 DVSS.n4808 0.00750714
R19078 DVSS.n4872 DVSS.n4831 0.00750714
R19079 DVSS.n1798 DVSS.n1797 0.00750714
R19080 DVSS.n2145 DVSS.n2144 0.00750714
R19081 DVSS.n3054 DVSS.n2682 0.0075
R19082 DVSS.n3524 DVSS.n3091 0.0075
R19083 DVSS.n3046 DVSS.n2687 0.0075
R19084 DVSS.n3273 DVSS.n3089 0.0075
R19085 DVSS.n1208 DVSS.n1183 0.00745122
R19086 DVSS.n1198 DVSS.n1186 0.00745122
R19087 DVSS.n2115 DVSS.n2114 0.00739189
R19088 DVSS.n2112 DVSS.n2086 0.00739189
R19089 DVSS.n4791 DVSS.n4790 0.00730488
R19090 DVSS.n4790 DVSS.n4787 0.00730488
R19091 DVSS.n4757 DVSS.n1220 0.00730488
R19092 DVSS.n4919 DVSS.n1220 0.00730488
R19093 DVSS.n4721 DVSS.n4720 0.00730488
R19094 DVSS.n4721 DVSS.n1242 0.00730488
R19095 DVSS.n4682 DVSS.n4681 0.00730488
R19096 DVSS.n4682 DVSS.n1263 0.00730488
R19097 DVSS.n4598 DVSS.n4597 0.00730488
R19098 DVSS.n4597 DVSS.n4594 0.00730488
R19099 DVSS.n4564 DVSS.n4494 0.00730488
R19100 DVSS.n4671 DVSS.n4494 0.00730488
R19101 DVSS.n2806 DVSS.n2805 0.00716667
R19102 DVSS.n2807 DVSS.n2806 0.00716667
R19103 DVSS.n2807 DVSS.n2774 0.00716667
R19104 DVSS.n2847 DVSS.n2774 0.00716667
R19105 DVSS.n2848 DVSS.n2847 0.00716667
R19106 DVSS.n2849 DVSS.n2848 0.00716667
R19107 DVSS.n2850 DVSS.n2849 0.00716667
R19108 DVSS.n2851 DVSS.n2850 0.00716667
R19109 DVSS.n2851 DVSS.n2754 0.00716667
R19110 DVSS.n2896 DVSS.n2754 0.00716667
R19111 DVSS.n2897 DVSS.n2896 0.00716667
R19112 DVSS.n2898 DVSS.n2897 0.00716667
R19113 DVSS.n2899 DVSS.n2898 0.00716667
R19114 DVSS.n2900 DVSS.n2899 0.00716667
R19115 DVSS.n2901 DVSS.n2900 0.00716667
R19116 DVSS.n2901 DVSS.n2732 0.00716667
R19117 DVSS.n2959 DVSS.n2732 0.00716667
R19118 DVSS.n2960 DVSS.n2959 0.00716667
R19119 DVSS.n2961 DVSS.n2960 0.00716667
R19120 DVSS.n2961 DVSS.n2719 0.00716667
R19121 DVSS.n2978 DVSS.n2719 0.00716667
R19122 DVSS.n2979 DVSS.n2978 0.00716667
R19123 DVSS.n2980 DVSS.n2979 0.00716667
R19124 DVSS.n2981 DVSS.n2980 0.00716667
R19125 DVSS.n2982 DVSS.n2981 0.00716667
R19126 DVSS.n2982 DVSS.n2699 0.00716667
R19127 DVSS.n3024 DVSS.n2699 0.00716667
R19128 DVSS.n3025 DVSS.n3024 0.00716667
R19129 DVSS.n3026 DVSS.n3025 0.00716667
R19130 DVSS.n3027 DVSS.n3026 0.00716667
R19131 DVSS.n3029 DVSS.n3027 0.00716667
R19132 DVSS.n3029 DVSS.n3028 0.00716667
R19133 DVSS.n3028 DVSS.n2679 0.00716667
R19134 DVSS.n2679 DVSS.n2677 0.00716667
R19135 DVSS.n3067 DVSS.n2677 0.00716667
R19136 DVSS.n3068 DVSS.n3067 0.00716667
R19137 DVSS.n3069 DVSS.n3068 0.00716667
R19138 DVSS.n3070 DVSS.n3069 0.00716667
R19139 DVSS.n3084 DVSS.n3070 0.00716667
R19140 DVSS.n3085 DVSS.n3084 0.00716667
R19141 DVSS.n3086 DVSS.n3085 0.00716667
R19142 DVSS.n3087 DVSS.n3086 0.00716667
R19143 DVSS.n3104 DVSS.n3087 0.00716667
R19144 DVSS.n3105 DVSS.n3104 0.00716667
R19145 DVSS.n3106 DVSS.n3105 0.00716667
R19146 DVSS.n3107 DVSS.n3106 0.00716667
R19147 DVSS.n3121 DVSS.n3107 0.00716667
R19148 DVSS.n3122 DVSS.n3121 0.00716667
R19149 DVSS.n3123 DVSS.n3122 0.00716667
R19150 DVSS.n3124 DVSS.n3123 0.00716667
R19151 DVSS.n3140 DVSS.n3124 0.00716667
R19152 DVSS.n3141 DVSS.n3140 0.00716667
R19153 DVSS.n3142 DVSS.n3141 0.00716667
R19154 DVSS.n3143 DVSS.n3142 0.00716667
R19155 DVSS.n3158 DVSS.n3143 0.00716667
R19156 DVSS.n3159 DVSS.n3158 0.00716667
R19157 DVSS.n3160 DVSS.n3159 0.00716667
R19158 DVSS.n3161 DVSS.n3160 0.00716667
R19159 DVSS.n3175 DVSS.n3161 0.00716667
R19160 DVSS.n3176 DVSS.n3175 0.00716667
R19161 DVSS.n3177 DVSS.n3176 0.00716667
R19162 DVSS.n3178 DVSS.n3177 0.00716667
R19163 DVSS.n3195 DVSS.n3178 0.00716667
R19164 DVSS.n3196 DVSS.n3195 0.00716667
R19165 DVSS.n3197 DVSS.n3196 0.00716667
R19166 DVSS.n3198 DVSS.n3197 0.00716667
R19167 DVSS.n3213 DVSS.n3198 0.00716667
R19168 DVSS.n3214 DVSS.n3213 0.00716667
R19169 DVSS.n3215 DVSS.n3214 0.00716667
R19170 DVSS.n3216 DVSS.n3215 0.00716667
R19171 DVSS.n3230 DVSS.n3216 0.00716667
R19172 DVSS.n3231 DVSS.n3230 0.00716667
R19173 DVSS.n3232 DVSS.n3231 0.00716667
R19174 DVSS.n3233 DVSS.n3232 0.00716667
R19175 DVSS.n3378 DVSS.n3233 0.00716667
R19176 DVSS.n3379 DVSS.n3378 0.00716667
R19177 DVSS.n3380 DVSS.n3379 0.00716667
R19178 DVSS.n3381 DVSS.n3380 0.00716667
R19179 DVSS.n3382 DVSS.n3381 0.00716667
R19180 DVSS.n3384 DVSS.n3382 0.00716667
R19181 DVSS.n3385 DVSS.n3384 0.00716667
R19182 DVSS.n3386 DVSS.n3385 0.00716667
R19183 DVSS.n3389 DVSS.n3386 0.00716667
R19184 DVSS.n3390 DVSS.n3389 0.00716667
R19185 DVSS.n3391 DVSS.n3390 0.00716667
R19186 DVSS.n3392 DVSS.n3391 0.00716667
R19187 DVSS.n3394 DVSS.n3392 0.00716667
R19188 DVSS.n3395 DVSS.n3394 0.00716667
R19189 DVSS.n955 DVSS.n951 0.00712143
R19190 DVSS.n5362 DVSS.n5361 0.00712143
R19191 DVSS.n4934 DVSS.n1181 0.00712143
R19192 DVSS.n4856 DVSS.n1177 0.00712143
R19193 DVSS.n3894 DVSS.n3893 0.00712143
R19194 DVSS.n3847 DVSS.n1620 0.00705714
R19195 DVSS.n1625 DVSS.n1624 0.00705714
R19196 DVSS.n3841 DVSS.n3840 0.00705714
R19197 DVSS.n802 DVSS.n800 0.00700873
R19198 DVSS.n3548 DVSS.n2669 0.007
R19199 DVSS.n3532 DVSS.n3076 0.007
R19200 DVSS.n3255 DVSS.n2665 0.007
R19201 DVSS.n3267 DVSS.n3266 0.007
R19202 DVSS.n3887 DVSS.n3886 0.00699286
R19203 DVSS.n3874 DVSS.n1605 0.00699286
R19204 DVSS.n3906 DVSS.n3905 0.00692857
R19205 DVSS.n2169 DVSS.n2168 0.006875
R19206 DVSS.n2166 DVSS.n1796 0.006875
R19207 DVSS.n2178 DVSS.n1784 0.006875
R19208 DVSS.n2181 DVSS.n2180 0.006875
R19209 DVSS.n4705 DVSS.n1252 0.0068
R19210 DVSS.n4714 DVSS.n4712 0.0068
R19211 DVSS.n4713 DVSS.n1249 0.0068
R19212 DVSS.n4723 DVSS.n4722 0.0068
R19213 DVSS.n4731 DVSS.n1243 0.0068
R19214 DVSS.n4730 DVSS.n1244 0.0068
R19215 DVSS.n4736 DVSS.n1239 0.0068
R19216 DVSS.n4980 DVSS.n4979 0.0068
R19217 DVSS.n2408 DVSS.n2277 0.0068
R19218 DVSS.n1206 DVSS.n1183 0.00671951
R19219 DVSS.n1200 DVSS.n1186 0.00671951
R19220 DVSS.n2967 DVSS.n2725 0.0067069
R19221 DVSS.n2939 DVSS.n2938 0.0067069
R19222 DVSS.n5365 DVSS.n949 0.00658571
R19223 DVSS.n5366 DVSS.n5365 0.00658571
R19224 DVSS.n5367 DVSS.n5366 0.00658571
R19225 DVSS.n5367 DVSS.n945 0.00658571
R19226 DVSS.n5373 DVSS.n945 0.00658571
R19227 DVSS.n5374 DVSS.n5373 0.00658571
R19228 DVSS.n5375 DVSS.n5374 0.00658571
R19229 DVSS.n5375 DVSS.n941 0.00658571
R19230 DVSS.n5381 DVSS.n941 0.00658571
R19231 DVSS.n5382 DVSS.n5381 0.00658571
R19232 DVSS.n5383 DVSS.n5382 0.00658571
R19233 DVSS.n5383 DVSS.n937 0.00658571
R19234 DVSS.n5389 DVSS.n937 0.00658571
R19235 DVSS.n5390 DVSS.n5389 0.00658571
R19236 DVSS.n5391 DVSS.n5390 0.00658571
R19237 DVSS.n5391 DVSS.n933 0.00658571
R19238 DVSS.n5397 DVSS.n933 0.00658571
R19239 DVSS.n5398 DVSS.n5397 0.00658571
R19240 DVSS.n5399 DVSS.n5398 0.00658571
R19241 DVSS.n5399 DVSS.n929 0.00658571
R19242 DVSS.n5405 DVSS.n929 0.00658571
R19243 DVSS.n5406 DVSS.n5405 0.00658571
R19244 DVSS.n5407 DVSS.n5406 0.00658571
R19245 DVSS.n5407 DVSS.n925 0.00658571
R19246 DVSS.n5413 DVSS.n925 0.00658571
R19247 DVSS.n5414 DVSS.n5413 0.00658571
R19248 DVSS.n5415 DVSS.n5414 0.00658571
R19249 DVSS.n5415 DVSS.n921 0.00658571
R19250 DVSS.n5421 DVSS.n921 0.00658571
R19251 DVSS.n5422 DVSS.n5421 0.00658571
R19252 DVSS.n5423 DVSS.n5422 0.00658571
R19253 DVSS.n5423 DVSS.n917 0.00658571
R19254 DVSS.n5429 DVSS.n917 0.00658571
R19255 DVSS.n5430 DVSS.n5429 0.00658571
R19256 DVSS.n5431 DVSS.n5430 0.00658571
R19257 DVSS.n5431 DVSS.n913 0.00658571
R19258 DVSS.n5437 DVSS.n913 0.00658571
R19259 DVSS.n5438 DVSS.n5437 0.00658571
R19260 DVSS.n5439 DVSS.n5438 0.00658571
R19261 DVSS.n5439 DVSS.n909 0.00658571
R19262 DVSS.n5445 DVSS.n909 0.00658571
R19263 DVSS.n5446 DVSS.n5445 0.00658571
R19264 DVSS.n5447 DVSS.n5446 0.00658571
R19265 DVSS.n5447 DVSS.n905 0.00658571
R19266 DVSS.n5453 DVSS.n905 0.00658571
R19267 DVSS.n5454 DVSS.n5453 0.00658571
R19268 DVSS.n5455 DVSS.n5454 0.00658571
R19269 DVSS.n5455 DVSS.n901 0.00658571
R19270 DVSS.n5461 DVSS.n901 0.00658571
R19271 DVSS.n5462 DVSS.n5461 0.00658571
R19272 DVSS.n5463 DVSS.n5462 0.00658571
R19273 DVSS.n5463 DVSS.n897 0.00658571
R19274 DVSS.n5469 DVSS.n897 0.00658571
R19275 DVSS.n5470 DVSS.n5469 0.00658571
R19276 DVSS.n5471 DVSS.n5470 0.00658571
R19277 DVSS.n5471 DVSS.n893 0.00658571
R19278 DVSS.n5477 DVSS.n893 0.00658571
R19279 DVSS.n5478 DVSS.n5477 0.00658571
R19280 DVSS.n5479 DVSS.n5478 0.00658571
R19281 DVSS.n5479 DVSS.n889 0.00658571
R19282 DVSS.n5485 DVSS.n889 0.00658571
R19283 DVSS.n5486 DVSS.n5485 0.00658571
R19284 DVSS.n5487 DVSS.n5486 0.00658571
R19285 DVSS.n5487 DVSS.n885 0.00658571
R19286 DVSS.n5493 DVSS.n885 0.00658571
R19287 DVSS.n5494 DVSS.n5493 0.00658571
R19288 DVSS.n5495 DVSS.n5494 0.00658571
R19289 DVSS.n5495 DVSS.n881 0.00658571
R19290 DVSS.n5501 DVSS.n881 0.00658571
R19291 DVSS.n5502 DVSS.n5501 0.00658571
R19292 DVSS.n5503 DVSS.n5502 0.00658571
R19293 DVSS.n5503 DVSS.n877 0.00658571
R19294 DVSS.n5509 DVSS.n877 0.00658571
R19295 DVSS.n5510 DVSS.n5509 0.00658571
R19296 DVSS.n5511 DVSS.n5510 0.00658571
R19297 DVSS.n5511 DVSS.n873 0.00658571
R19298 DVSS.n5517 DVSS.n873 0.00658571
R19299 DVSS.n5518 DVSS.n5517 0.00658571
R19300 DVSS.n5519 DVSS.n5518 0.00658571
R19301 DVSS.n5519 DVSS.n869 0.00658571
R19302 DVSS.n5525 DVSS.n869 0.00658571
R19303 DVSS.n5526 DVSS.n5525 0.00658571
R19304 DVSS.n5527 DVSS.n5526 0.00658571
R19305 DVSS.n5527 DVSS.n865 0.00658571
R19306 DVSS.n5533 DVSS.n865 0.00658571
R19307 DVSS.n5534 DVSS.n5533 0.00658571
R19308 DVSS.n5535 DVSS.n5534 0.00658571
R19309 DVSS.n5535 DVSS.n861 0.00658571
R19310 DVSS.n5541 DVSS.n861 0.00658571
R19311 DVSS.n5542 DVSS.n5541 0.00658571
R19312 DVSS.n5543 DVSS.n5542 0.00658571
R19313 DVSS.n5543 DVSS.n857 0.00658571
R19314 DVSS.n5549 DVSS.n857 0.00658571
R19315 DVSS.n5550 DVSS.n5549 0.00658571
R19316 DVSS.n4549 DVSS.n4548 0.00658571
R19317 DVSS.n4549 DVSS.n4507 0.00658571
R19318 DVSS.n4555 DVSS.n4507 0.00658571
R19319 DVSS.n4556 DVSS.n4555 0.00658571
R19320 DVSS.n4557 DVSS.n4556 0.00658571
R19321 DVSS.n4557 DVSS.n4500 0.00658571
R19322 DVSS.n4570 DVSS.n4500 0.00658571
R19323 DVSS.n4571 DVSS.n4570 0.00658571
R19324 DVSS.n4666 DVSS.n4571 0.00658571
R19325 DVSS.n4666 DVSS.n4665 0.00658571
R19326 DVSS.n4665 DVSS.n4664 0.00658571
R19327 DVSS.n4664 DVSS.n4572 0.00658571
R19328 DVSS.n4658 DVSS.n4572 0.00658571
R19329 DVSS.n4658 DVSS.n4657 0.00658571
R19330 DVSS.n4657 DVSS.n4656 0.00658571
R19331 DVSS.n4656 DVSS.n4580 0.00658571
R19332 DVSS.n4588 DVSS.n4580 0.00658571
R19333 DVSS.n4646 DVSS.n4588 0.00658571
R19334 DVSS.n4646 DVSS.n4645 0.00658571
R19335 DVSS.n4645 DVSS.n4644 0.00658571
R19336 DVSS.n4644 DVSS.n4589 0.00658571
R19337 DVSS.n4607 DVSS.n4589 0.00658571
R19338 DVSS.n4633 DVSS.n4607 0.00658571
R19339 DVSS.n4633 DVSS.n4632 0.00658571
R19340 DVSS.n4632 DVSS.n4631 0.00658571
R19341 DVSS.n4631 DVSS.n4608 0.00658571
R19342 DVSS.n4625 DVSS.n4608 0.00658571
R19343 DVSS.n4625 DVSS.n4624 0.00658571
R19344 DVSS.n4624 DVSS.n4623 0.00658571
R19345 DVSS.n4623 DVSS.n4612 0.00658571
R19346 DVSS.n4612 DVSS.n1267 0.00658571
R19347 DVSS.n4686 DVSS.n1267 0.00658571
R19348 DVSS.n4687 DVSS.n4686 0.00658571
R19349 DVSS.n4688 DVSS.n4687 0.00658571
R19350 DVSS.n4688 DVSS.n1258 0.00658571
R19351 DVSS.n4699 DVSS.n1258 0.00658571
R19352 DVSS.n4700 DVSS.n4699 0.00658571
R19353 DVSS.n4701 DVSS.n4700 0.00658571
R19354 DVSS.n4701 DVSS.n1254 0.00658571
R19355 DVSS.n4708 DVSS.n1254 0.00658571
R19356 DVSS.n4709 DVSS.n4708 0.00658571
R19357 DVSS.n4710 DVSS.n4709 0.00658571
R19358 DVSS.n4710 DVSS.n1247 0.00658571
R19359 DVSS.n4725 DVSS.n1247 0.00658571
R19360 DVSS.n4726 DVSS.n4725 0.00658571
R19361 DVSS.n4728 DVSS.n4726 0.00658571
R19362 DVSS.n4728 DVSS.n4727 0.00658571
R19363 DVSS.n4727 DVSS.n1237 0.00658571
R19364 DVSS.n4740 DVSS.n1237 0.00658571
R19365 DVSS.n4741 DVSS.n4740 0.00658571
R19366 DVSS.n4742 DVSS.n4741 0.00658571
R19367 DVSS.n4742 DVSS.n1233 0.00658571
R19368 DVSS.n4748 DVSS.n1233 0.00658571
R19369 DVSS.n4749 DVSS.n4748 0.00658571
R19370 DVSS.n4750 DVSS.n4749 0.00658571
R19371 DVSS.n4750 DVSS.n1226 0.00658571
R19372 DVSS.n4763 DVSS.n1226 0.00658571
R19373 DVSS.n4764 DVSS.n4763 0.00658571
R19374 DVSS.n4914 DVSS.n4764 0.00658571
R19375 DVSS.n4914 DVSS.n4913 0.00658571
R19376 DVSS.n4913 DVSS.n4912 0.00658571
R19377 DVSS.n4912 DVSS.n4765 0.00658571
R19378 DVSS.n4906 DVSS.n4765 0.00658571
R19379 DVSS.n4906 DVSS.n4905 0.00658571
R19380 DVSS.n4905 DVSS.n4904 0.00658571
R19381 DVSS.n4904 DVSS.n4773 0.00658571
R19382 DVSS.n4781 DVSS.n4773 0.00658571
R19383 DVSS.n4894 DVSS.n4781 0.00658571
R19384 DVSS.n4894 DVSS.n4893 0.00658571
R19385 DVSS.n4893 DVSS.n4892 0.00658571
R19386 DVSS.n4892 DVSS.n4782 0.00658571
R19387 DVSS.n4800 DVSS.n4782 0.00658571
R19388 DVSS.n4881 DVSS.n4800 0.00658571
R19389 DVSS.n4881 DVSS.n4880 0.00658571
R19390 DVSS.n4880 DVSS.n4879 0.00658571
R19391 DVSS.n4879 DVSS.n4801 0.00658571
R19392 DVSS.n4839 DVSS.n4801 0.00658571
R19393 DVSS.n4840 DVSS.n4839 0.00658571
R19394 DVSS.n4869 DVSS.n4840 0.00658571
R19395 DVSS.n4869 DVSS.n4868 0.00658571
R19396 DVSS.n4868 DVSS.n4867 0.00658571
R19397 DVSS.n4867 DVSS.n4841 0.00658571
R19398 DVSS.n4861 DVSS.n4841 0.00658571
R19399 DVSS.n4861 DVSS.n4860 0.00658571
R19400 DVSS.n4860 DVSS.n4859 0.00658571
R19401 DVSS.n4859 DVSS.n4845 0.00658571
R19402 DVSS.n4849 DVSS.n4847 0.00658571
R19403 DVSS.n1541 DVSS.n1532 0.00658571
R19404 DVSS.n1542 DVSS.n1541 0.00658571
R19405 DVSS.n1543 DVSS.n1542 0.00658571
R19406 DVSS.n1543 DVSS.n1528 0.00658571
R19407 DVSS.n1549 DVSS.n1528 0.00658571
R19408 DVSS.n1550 DVSS.n1549 0.00658571
R19409 DVSS.n1551 DVSS.n1550 0.00658571
R19410 DVSS.n1551 DVSS.n1524 0.00658571
R19411 DVSS.n1557 DVSS.n1524 0.00658571
R19412 DVSS.n1558 DVSS.n1557 0.00658571
R19413 DVSS.n3934 DVSS.n1558 0.00658571
R19414 DVSS.n3934 DVSS.n3933 0.00658571
R19415 DVSS.n3933 DVSS.n3932 0.00658571
R19416 DVSS.n3932 DVSS.n1559 0.00658571
R19417 DVSS.n3926 DVSS.n1559 0.00658571
R19418 DVSS.n3926 DVSS.n3925 0.00658571
R19419 DVSS.n3925 DVSS.n3924 0.00658571
R19420 DVSS.n3924 DVSS.n1563 0.00658571
R19421 DVSS.n3918 DVSS.n1563 0.00658571
R19422 DVSS.n3918 DVSS.n3917 0.00658571
R19423 DVSS.n3917 DVSS.n3916 0.00658571
R19424 DVSS.n3916 DVSS.n1567 0.00658571
R19425 DVSS.n3910 DVSS.n1567 0.00658571
R19426 DVSS.n3910 DVSS.n3909 0.00658571
R19427 DVSS.n3909 DVSS.n3908 0.00658571
R19428 DVSS.n3908 DVSS.n1571 0.00658571
R19429 DVSS.n2495 DVSS.n1571 0.00658571
R19430 DVSS.n2496 DVSS.n2495 0.00658571
R19431 DVSS.n2496 DVSS.n2491 0.00658571
R19432 DVSS.n2502 DVSS.n2491 0.00658571
R19433 DVSS.n2503 DVSS.n2502 0.00658571
R19434 DVSS.n2504 DVSS.n2503 0.00658571
R19435 DVSS.n2504 DVSS.n2487 0.00658571
R19436 DVSS.n2510 DVSS.n2487 0.00658571
R19437 DVSS.n2511 DVSS.n2510 0.00658571
R19438 DVSS.n2512 DVSS.n2511 0.00658571
R19439 DVSS.n2512 DVSS.n2483 0.00658571
R19440 DVSS.n2518 DVSS.n2483 0.00658571
R19441 DVSS.n2519 DVSS.n2518 0.00658571
R19442 DVSS.n2520 DVSS.n2519 0.00658571
R19443 DVSS.n2520 DVSS.n2479 0.00658571
R19444 DVSS.n2526 DVSS.n2479 0.00658571
R19445 DVSS.n2527 DVSS.n2526 0.00658571
R19446 DVSS.n2528 DVSS.n2527 0.00658571
R19447 DVSS.n2528 DVSS.n2475 0.00658571
R19448 DVSS.n2534 DVSS.n2475 0.00658571
R19449 DVSS.n2535 DVSS.n2534 0.00658571
R19450 DVSS.n2536 DVSS.n2535 0.00658571
R19451 DVSS.n2536 DVSS.n2471 0.00658571
R19452 DVSS.n2542 DVSS.n2471 0.00658571
R19453 DVSS.n2543 DVSS.n2542 0.00658571
R19454 DVSS.n2544 DVSS.n2543 0.00658571
R19455 DVSS.n2544 DVSS.n2467 0.00658571
R19456 DVSS.n2550 DVSS.n2467 0.00658571
R19457 DVSS.n2551 DVSS.n2550 0.00658571
R19458 DVSS.n2552 DVSS.n2551 0.00658571
R19459 DVSS.n2552 DVSS.n2463 0.00658571
R19460 DVSS.n2558 DVSS.n2463 0.00658571
R19461 DVSS.n2559 DVSS.n2558 0.00658571
R19462 DVSS.n2560 DVSS.n2559 0.00658571
R19463 DVSS.n2560 DVSS.n2459 0.00658571
R19464 DVSS.n2566 DVSS.n2459 0.00658571
R19465 DVSS.n2567 DVSS.n2566 0.00658571
R19466 DVSS.n2568 DVSS.n2567 0.00658571
R19467 DVSS.n2568 DVSS.n2455 0.00658571
R19468 DVSS.n2574 DVSS.n2455 0.00658571
R19469 DVSS.n2575 DVSS.n2574 0.00658571
R19470 DVSS.n2576 DVSS.n2575 0.00658571
R19471 DVSS.n2576 DVSS.n2451 0.00658571
R19472 DVSS.n2582 DVSS.n2451 0.00658571
R19473 DVSS.n2583 DVSS.n2582 0.00658571
R19474 DVSS.n2584 DVSS.n2583 0.00658571
R19475 DVSS.n2584 DVSS.n2447 0.00658571
R19476 DVSS.n2590 DVSS.n2447 0.00658571
R19477 DVSS.n2591 DVSS.n2590 0.00658571
R19478 DVSS.n2592 DVSS.n2591 0.00658571
R19479 DVSS.n2592 DVSS.n2443 0.00658571
R19480 DVSS.n2598 DVSS.n2443 0.00658571
R19481 DVSS.n2599 DVSS.n2598 0.00658571
R19482 DVSS.n2600 DVSS.n2599 0.00658571
R19483 DVSS.n2600 DVSS.n2439 0.00658571
R19484 DVSS.n2606 DVSS.n2439 0.00658571
R19485 DVSS.n2607 DVSS.n2606 0.00658571
R19486 DVSS.n2608 DVSS.n2607 0.00658571
R19487 DVSS.n2608 DVSS.n2435 0.00658571
R19488 DVSS.n2614 DVSS.n2435 0.00658571
R19489 DVSS.n2615 DVSS.n2614 0.00658571
R19490 DVSS.n2616 DVSS.n2615 0.00658571
R19491 DVSS.n2616 DVSS.n2431 0.00658571
R19492 DVSS.n2622 DVSS.n2431 0.00658571
R19493 DVSS.n2623 DVSS.n2622 0.00658571
R19494 DVSS.n2624 DVSS.n2623 0.00658571
R19495 DVSS.n2624 DVSS.n2427 0.00658571
R19496 DVSS.n2630 DVSS.n2427 0.00658571
R19497 DVSS.n2631 DVSS.n2630 0.00658571
R19498 DVSS.n2634 DVSS.n2631 0.00658571
R19499 DVSS.n2634 DVSS.n2633 0.00658571
R19500 DVSS.n2652 DVSS.n2267 0.00658571
R19501 DVSS.n3891 DVSS.n1598 0.00658571
R19502 DVSS.n3891 DVSS.n3890 0.00658571
R19503 DVSS.n3890 DVSS.n3889 0.00658571
R19504 DVSS.n3889 DVSS.n1599 0.00658571
R19505 DVSS.n3882 DVSS.n1599 0.00658571
R19506 DVSS.n3882 DVSS.n3881 0.00658571
R19507 DVSS.n3881 DVSS.n3880 0.00658571
R19508 DVSS.n3880 DVSS.n1603 0.00658571
R19509 DVSS.n3872 DVSS.n1603 0.00658571
R19510 DVSS.n3872 DVSS.n3871 0.00658571
R19511 DVSS.n3871 DVSS.n3870 0.00658571
R19512 DVSS.n3870 DVSS.n1607 0.00658571
R19513 DVSS.n3864 DVSS.n1607 0.00658571
R19514 DVSS.n3864 DVSS.n3863 0.00658571
R19515 DVSS.n3863 DVSS.n3862 0.00658571
R19516 DVSS.n3862 DVSS.n1612 0.00658571
R19517 DVSS.n3853 DVSS.n1612 0.00658571
R19518 DVSS.n3853 DVSS.n3852 0.00658571
R19519 DVSS.n3852 DVSS.n3851 0.00658571
R19520 DVSS.n3851 DVSS.n1617 0.00658571
R19521 DVSS.n3845 DVSS.n1617 0.00658571
R19522 DVSS.n3845 DVSS.n3844 0.00658571
R19523 DVSS.n3844 DVSS.n3843 0.00658571
R19524 DVSS.n3843 DVSS.n1622 0.00658571
R19525 DVSS.n1634 DVSS.n1622 0.00658571
R19526 DVSS.n3824 DVSS.n1634 0.00658571
R19527 DVSS.n3824 DVSS.n3823 0.00658571
R19528 DVSS.n3823 DVSS.n3822 0.00658571
R19529 DVSS.n3822 DVSS.n1636 0.00658571
R19530 DVSS.n3816 DVSS.n1636 0.00658571
R19531 DVSS.n3816 DVSS.n3815 0.00658571
R19532 DVSS.n3815 DVSS.n3814 0.00658571
R19533 DVSS.n3814 DVSS.n1641 0.00658571
R19534 DVSS.n3808 DVSS.n1641 0.00658571
R19535 DVSS.n3808 DVSS.n3807 0.00658571
R19536 DVSS.n3807 DVSS.n3806 0.00658571
R19537 DVSS.n3806 DVSS.n1645 0.00658571
R19538 DVSS.n3799 DVSS.n1645 0.00658571
R19539 DVSS.n3799 DVSS.n3798 0.00658571
R19540 DVSS.n3798 DVSS.n3797 0.00658571
R19541 DVSS.n3797 DVSS.n1651 0.00658571
R19542 DVSS.n1667 DVSS.n1651 0.00658571
R19543 DVSS.n1667 DVSS.n1665 0.00658571
R19544 DVSS.n1677 DVSS.n1665 0.00658571
R19545 DVSS.n1678 DVSS.n1677 0.00658571
R19546 DVSS.n3784 DVSS.n1678 0.00658571
R19547 DVSS.n3784 DVSS.n3783 0.00658571
R19548 DVSS.n3783 DVSS.n3782 0.00658571
R19549 DVSS.n3782 DVSS.n1679 0.00658571
R19550 DVSS.n3776 DVSS.n1679 0.00658571
R19551 DVSS.n3776 DVSS.n3775 0.00658571
R19552 DVSS.n3775 DVSS.n3774 0.00658571
R19553 DVSS.n3774 DVSS.n1684 0.00658571
R19554 DVSS.n3680 DVSS.n1684 0.00658571
R19555 DVSS.n3681 DVSS.n3680 0.00658571
R19556 DVSS.n3682 DVSS.n3681 0.00658571
R19557 DVSS.n3682 DVSS.n3674 0.00658571
R19558 DVSS.n3688 DVSS.n3674 0.00658571
R19559 DVSS.n3689 DVSS.n3688 0.00658571
R19560 DVSS.n3690 DVSS.n3689 0.00658571
R19561 DVSS.n3690 DVSS.n3670 0.00658571
R19562 DVSS.n3696 DVSS.n3670 0.00658571
R19563 DVSS.n3697 DVSS.n3696 0.00658571
R19564 DVSS.n3698 DVSS.n3697 0.00658571
R19565 DVSS.n3698 DVSS.n3666 0.00658571
R19566 DVSS.n3704 DVSS.n3666 0.00658571
R19567 DVSS.n3705 DVSS.n3704 0.00658571
R19568 DVSS.n3706 DVSS.n3705 0.00658571
R19569 DVSS.n3706 DVSS.n3662 0.00658571
R19570 DVSS.n3712 DVSS.n3662 0.00658571
R19571 DVSS.n3713 DVSS.n3712 0.00658571
R19572 DVSS.n3714 DVSS.n3713 0.00658571
R19573 DVSS.n3714 DVSS.n3658 0.00658571
R19574 DVSS.n3720 DVSS.n3658 0.00658571
R19575 DVSS.n3721 DVSS.n3720 0.00658571
R19576 DVSS.n3741 DVSS.n3721 0.00658571
R19577 DVSS.n3741 DVSS.n3740 0.00658571
R19578 DVSS.n3740 DVSS.n3739 0.00658571
R19579 DVSS.n3739 DVSS.n3722 0.00658571
R19580 DVSS.n3733 DVSS.n3722 0.00658571
R19581 DVSS.n3733 DVSS.n3732 0.00658571
R19582 DVSS.n3732 DVSS.n3731 0.00658571
R19583 DVSS.n3731 DVSS.n3726 0.00658571
R19584 DVSS.n2224 DVSS.n2223 0.00658571
R19585 DVSS.n2223 DVSS.n2222 0.00658571
R19586 DVSS.n2222 DVSS.n1737 0.00658571
R19587 DVSS.n2216 DVSS.n1737 0.00658571
R19588 DVSS.n2216 DVSS.n2215 0.00658571
R19589 DVSS.n2215 DVSS.n2214 0.00658571
R19590 DVSS.n2214 DVSS.n1742 0.00658571
R19591 DVSS.n1895 DVSS.n1742 0.00658571
R19592 DVSS.n1896 DVSS.n1895 0.00658571
R19593 DVSS.n1896 DVSS.n1886 0.00658571
R19594 DVSS.n1904 DVSS.n1886 0.00658571
R19595 DVSS.n1905 DVSS.n1904 0.00658571
R19596 DVSS.n1906 DVSS.n1905 0.00658571
R19597 DVSS.n1906 DVSS.n1766 0.00658571
R19598 DVSS.n2193 DVSS.n1766 0.00658571
R19599 DVSS.n2193 DVSS.n2192 0.00658571
R19600 DVSS.n2192 DVSS.n2191 0.00658571
R19601 DVSS.n2191 DVSS.n1767 0.00658571
R19602 DVSS.n1871 DVSS.n1767 0.00658571
R19603 DVSS.n1871 DVSS.n1793 0.00658571
R19604 DVSS.n2175 DVSS.n1793 0.00658571
R19605 DVSS.n2175 DVSS.n2174 0.00658571
R19606 DVSS.n2174 DVSS.n2173 0.00658571
R19607 DVSS.n2173 DVSS.n1794 0.00658571
R19608 DVSS.n2142 DVSS.n1794 0.00658571
R19609 DVSS.n2142 DVSS.n2141 0.00658571
R19610 DVSS.n2141 DVSS.n2140 0.00658571
R19611 DVSS.n2140 DVSS.n1928 0.00658571
R19612 DVSS.n1969 DVSS.n1928 0.00658571
R19613 DVSS.n1970 DVSS.n1969 0.00658571
R19614 DVSS.n1971 DVSS.n1970 0.00658571
R19615 DVSS.n1971 DVSS.n1956 0.00658571
R19616 DVSS.n1987 DVSS.n1956 0.00658571
R19617 DVSS.n1988 DVSS.n1987 0.00658571
R19618 DVSS.n2121 DVSS.n1988 0.00658571
R19619 DVSS.n2121 DVSS.n2120 0.00658571
R19620 DVSS.n2120 DVSS.n2119 0.00658571
R19621 DVSS.n2119 DVSS.n1989 0.00658571
R19622 DVSS.n1991 DVSS.n1989 0.00658571
R19623 DVSS.n1994 DVSS.n1991 0.00658571
R19624 DVSS.n2077 DVSS.n1994 0.00658571
R19625 DVSS.n2077 DVSS.n2076 0.00658571
R19626 DVSS.n2076 DVSS.n2075 0.00658571
R19627 DVSS.n2075 DVSS.n1995 0.00658571
R19628 DVSS.n2069 DVSS.n1995 0.00658571
R19629 DVSS.n2069 DVSS.n2068 0.00658571
R19630 DVSS.n2068 DVSS.n2067 0.00658571
R19631 DVSS.n2067 DVSS.n1999 0.00658571
R19632 DVSS.n2061 DVSS.n1999 0.00658571
R19633 DVSS.n2061 DVSS.n2060 0.00658571
R19634 DVSS.n2060 DVSS.n2059 0.00658571
R19635 DVSS.n2059 DVSS.n2003 0.00658571
R19636 DVSS.n2053 DVSS.n2003 0.00658571
R19637 DVSS.n2053 DVSS.n2052 0.00658571
R19638 DVSS.n2052 DVSS.n2051 0.00658571
R19639 DVSS.n2051 DVSS.n2007 0.00658571
R19640 DVSS.n2045 DVSS.n2007 0.00658571
R19641 DVSS.n2045 DVSS.n2044 0.00658571
R19642 DVSS.n2044 DVSS.n2043 0.00658571
R19643 DVSS.n2043 DVSS.n2011 0.00658571
R19644 DVSS.n2037 DVSS.n2011 0.00658571
R19645 DVSS.n2037 DVSS.n2036 0.00658571
R19646 DVSS.n2036 DVSS.n2035 0.00658571
R19647 DVSS.n2035 DVSS.n2015 0.00658571
R19648 DVSS.n2029 DVSS.n2015 0.00658571
R19649 DVSS.n2029 DVSS.n2028 0.00658571
R19650 DVSS.n2028 DVSS.n2027 0.00658571
R19651 DVSS.n2027 DVSS.n2019 0.00658571
R19652 DVSS.n2021 DVSS.n2019 0.00658571
R19653 DVSS.n1375 DVSS.n1372 0.00658571
R19654 DVSS.n4175 DVSS.n1375 0.00658571
R19655 DVSS.n4175 DVSS.n4174 0.00658571
R19656 DVSS.n4174 DVSS.n4173 0.00658571
R19657 DVSS.n4173 DVSS.n1376 0.00658571
R19658 DVSS.n4165 DVSS.n1376 0.00658571
R19659 DVSS.n4165 DVSS.n4164 0.00658571
R19660 DVSS.n4164 DVSS.n4163 0.00658571
R19661 DVSS.n4163 DVSS.n1393 0.00658571
R19662 DVSS.n4157 DVSS.n1393 0.00658571
R19663 DVSS.n4157 DVSS.n4156 0.00658571
R19664 DVSS.n4156 DVSS.n4155 0.00658571
R19665 DVSS.n4155 DVSS.n1397 0.00658571
R19666 DVSS.n4149 DVSS.n1397 0.00658571
R19667 DVSS.n4149 DVSS.n4148 0.00658571
R19668 DVSS.n4148 DVSS.n4147 0.00658571
R19669 DVSS.n4147 DVSS.n1401 0.00658571
R19670 DVSS.n4141 DVSS.n1401 0.00658571
R19671 DVSS.n4141 DVSS.n4140 0.00658571
R19672 DVSS.n4140 DVSS.n4139 0.00658571
R19673 DVSS.n4139 DVSS.n1405 0.00658571
R19674 DVSS.n4133 DVSS.n1405 0.00658571
R19675 DVSS.n4133 DVSS.n4132 0.00658571
R19676 DVSS.n4132 DVSS.n4131 0.00658571
R19677 DVSS.n4131 DVSS.n1409 0.00658571
R19678 DVSS.n4125 DVSS.n1409 0.00658571
R19679 DVSS.n4125 DVSS.n4124 0.00658571
R19680 DVSS.n4124 DVSS.n4123 0.00658571
R19681 DVSS.n4123 DVSS.n1413 0.00658571
R19682 DVSS.n4117 DVSS.n1413 0.00658571
R19683 DVSS.n4117 DVSS.n4116 0.00658571
R19684 DVSS.n4116 DVSS.n4115 0.00658571
R19685 DVSS.n4115 DVSS.n1417 0.00658571
R19686 DVSS.n4109 DVSS.n1417 0.00658571
R19687 DVSS.n4109 DVSS.n4108 0.00658571
R19688 DVSS.n4108 DVSS.n4107 0.00658571
R19689 DVSS.n4107 DVSS.n1421 0.00658571
R19690 DVSS.n4101 DVSS.n1421 0.00658571
R19691 DVSS.n4101 DVSS.n4100 0.00658571
R19692 DVSS.n4100 DVSS.n4099 0.00658571
R19693 DVSS.n4099 DVSS.n1425 0.00658571
R19694 DVSS.n4009 DVSS.n1425 0.00658571
R19695 DVSS.n4010 DVSS.n4009 0.00658571
R19696 DVSS.n4090 DVSS.n4010 0.00658571
R19697 DVSS.n4090 DVSS.n4089 0.00658571
R19698 DVSS.n4089 DVSS.n4088 0.00658571
R19699 DVSS.n4088 DVSS.n4011 0.00658571
R19700 DVSS.n4082 DVSS.n4011 0.00658571
R19701 DVSS.n4082 DVSS.n4081 0.00658571
R19702 DVSS.n4081 DVSS.n4080 0.00658571
R19703 DVSS.n4080 DVSS.n4015 0.00658571
R19704 DVSS.n4074 DVSS.n4015 0.00658571
R19705 DVSS.n4074 DVSS.n4073 0.00658571
R19706 DVSS.n4073 DVSS.n4072 0.00658571
R19707 DVSS.n4072 DVSS.n4019 0.00658571
R19708 DVSS.n4066 DVSS.n4019 0.00658571
R19709 DVSS.n4066 DVSS.n4065 0.00658571
R19710 DVSS.n4065 DVSS.n4064 0.00658571
R19711 DVSS.n4064 DVSS.n4023 0.00658571
R19712 DVSS.n4058 DVSS.n4023 0.00658571
R19713 DVSS.n4058 DVSS.n4057 0.00658571
R19714 DVSS.n4057 DVSS.n4056 0.00658571
R19715 DVSS.n4056 DVSS.n4027 0.00658571
R19716 DVSS.n4050 DVSS.n4027 0.00658571
R19717 DVSS.n4050 DVSS.n4049 0.00658571
R19718 DVSS.n4049 DVSS.n4048 0.00658571
R19719 DVSS.n4048 DVSS.n4031 0.00658571
R19720 DVSS.n4042 DVSS.n4031 0.00658571
R19721 DVSS.n4042 DVSS.n4041 0.00658571
R19722 DVSS.n4041 DVSS.n4040 0.00658571
R19723 DVSS.n4040 DVSS.n4035 0.00658571
R19724 DVSS.n5104 DVSS.n5103 0.00658571
R19725 DVSS.n5103 DVSS.n5102 0.00658571
R19726 DVSS.n5102 DVSS.n1085 0.00658571
R19727 DVSS.n5096 DVSS.n1085 0.00658571
R19728 DVSS.n5096 DVSS.n5095 0.00658571
R19729 DVSS.n5095 DVSS.n5094 0.00658571
R19730 DVSS.n5094 DVSS.n1090 0.00658571
R19731 DVSS.n5088 DVSS.n1090 0.00658571
R19732 DVSS.n5088 DVSS.n5087 0.00658571
R19733 DVSS.n5087 DVSS.n5086 0.00658571
R19734 DVSS.n5086 DVSS.n1094 0.00658571
R19735 DVSS.n5080 DVSS.n1094 0.00658571
R19736 DVSS.n5080 DVSS.n5079 0.00658571
R19737 DVSS.n5079 DVSS.n5078 0.00658571
R19738 DVSS.n5078 DVSS.n1098 0.00658571
R19739 DVSS.n5071 DVSS.n1098 0.00658571
R19740 DVSS.n5071 DVSS.n5070 0.00658571
R19741 DVSS.n5070 DVSS.n5069 0.00658571
R19742 DVSS.n5069 DVSS.n1104 0.00658571
R19743 DVSS.n5063 DVSS.n1104 0.00658571
R19744 DVSS.n5063 DVSS.n5062 0.00658571
R19745 DVSS.n5062 DVSS.n5061 0.00658571
R19746 DVSS.n5061 DVSS.n1108 0.00658571
R19747 DVSS.n5052 DVSS.n1108 0.00658571
R19748 DVSS.n5052 DVSS.n5051 0.00658571
R19749 DVSS.n5051 DVSS.n5050 0.00658571
R19750 DVSS.n5050 DVSS.n1115 0.00658571
R19751 DVSS.n5041 DVSS.n1115 0.00658571
R19752 DVSS.n5041 DVSS.n5040 0.00658571
R19753 DVSS.n5040 DVSS.n5039 0.00658571
R19754 DVSS.n5039 DVSS.n1123 0.00658571
R19755 DVSS.n5033 DVSS.n1123 0.00658571
R19756 DVSS.n5033 DVSS.n5032 0.00658571
R19757 DVSS.n5032 DVSS.n5031 0.00658571
R19758 DVSS.n5031 DVSS.n1128 0.00658571
R19759 DVSS.n5025 DVSS.n1128 0.00658571
R19760 DVSS.n5025 DVSS.n5024 0.00658571
R19761 DVSS.n5024 DVSS.n5023 0.00658571
R19762 DVSS.n5023 DVSS.n1132 0.00658571
R19763 DVSS.n5017 DVSS.n1132 0.00658571
R19764 DVSS.n5017 DVSS.n5016 0.00658571
R19765 DVSS.n5016 DVSS.n5015 0.00658571
R19766 DVSS.n5015 DVSS.n1136 0.00658571
R19767 DVSS.n5009 DVSS.n1136 0.00658571
R19768 DVSS.n5009 DVSS.n5008 0.00658571
R19769 DVSS.n5008 DVSS.n5007 0.00658571
R19770 DVSS.n5007 DVSS.n1140 0.00658571
R19771 DVSS.n5001 DVSS.n1140 0.00658571
R19772 DVSS.n5001 DVSS.n5000 0.00658571
R19773 DVSS.n5000 DVSS.n4999 0.00658571
R19774 DVSS.n4999 DVSS.n1144 0.00658571
R19775 DVSS.n4993 DVSS.n1144 0.00658571
R19776 DVSS.n4993 DVSS.n4992 0.00658571
R19777 DVSS.n4992 DVSS.n4991 0.00658571
R19778 DVSS.n4991 DVSS.n1148 0.00658571
R19779 DVSS.n4985 DVSS.n1148 0.00658571
R19780 DVSS.n4985 DVSS.n4984 0.00658571
R19781 DVSS.n4984 DVSS.n4983 0.00658571
R19782 DVSS.n4983 DVSS.n1152 0.00658571
R19783 DVSS.n2320 DVSS.n1152 0.00658571
R19784 DVSS.n2321 DVSS.n2320 0.00658571
R19785 DVSS.n2321 DVSS.n2317 0.00658571
R19786 DVSS.n2327 DVSS.n2317 0.00658571
R19787 DVSS.n2328 DVSS.n2327 0.00658571
R19788 DVSS.n2329 DVSS.n2328 0.00658571
R19789 DVSS.n2329 DVSS.n2313 0.00658571
R19790 DVSS.n2335 DVSS.n2313 0.00658571
R19791 DVSS.n2336 DVSS.n2335 0.00658571
R19792 DVSS.n2337 DVSS.n2336 0.00658571
R19793 DVSS.n2337 DVSS.n2309 0.00658571
R19794 DVSS.n2343 DVSS.n2309 0.00658571
R19795 DVSS.n2344 DVSS.n2343 0.00658571
R19796 DVSS.n2345 DVSS.n2344 0.00658571
R19797 DVSS.n2345 DVSS.n2305 0.00658571
R19798 DVSS.n2351 DVSS.n2305 0.00658571
R19799 DVSS.n2352 DVSS.n2351 0.00658571
R19800 DVSS.n2353 DVSS.n2352 0.00658571
R19801 DVSS.n2353 DVSS.n2301 0.00658571
R19802 DVSS.n2359 DVSS.n2301 0.00658571
R19803 DVSS.n2360 DVSS.n2359 0.00658571
R19804 DVSS.n2361 DVSS.n2360 0.00658571
R19805 DVSS.n2361 DVSS.n2297 0.00658571
R19806 DVSS.n2367 DVSS.n2297 0.00658571
R19807 DVSS.n2368 DVSS.n2367 0.00658571
R19808 DVSS.n2369 DVSS.n2368 0.00658571
R19809 DVSS.n2369 DVSS.n2293 0.00658571
R19810 DVSS.n2375 DVSS.n2293 0.00658571
R19811 DVSS.n2376 DVSS.n2375 0.00658571
R19812 DVSS.n2377 DVSS.n2376 0.00658571
R19813 DVSS.n2377 DVSS.n2289 0.00658571
R19814 DVSS.n2383 DVSS.n2289 0.00658571
R19815 DVSS.n2384 DVSS.n2383 0.00658571
R19816 DVSS.n2386 DVSS.n2384 0.00658571
R19817 DVSS.n2386 DVSS.n2385 0.00658571
R19818 DVSS.n2385 DVSS.n2285 0.00658571
R19819 DVSS.n2394 DVSS.n2285 0.00658571
R19820 DVSS.n2401 DVSS.n2400 0.00658571
R19821 DVSS.n2100 DVSS.n1805 0.00658108
R19822 DVSS.n1829 DVSS.n1818 0.00658108
R19823 DVSS.n4560 DVSS.n4559 0.00654286
R19824 DVSS.n4505 DVSS.n4502 0.00654286
R19825 DVSS.n4568 DVSS.n4566 0.00654286
R19826 DVSS.n4567 DVSS.n4496 0.00654286
R19827 DVSS.n4669 DVSS.n4668 0.00654286
R19828 DVSS.n4574 DVSS.n4497 0.00654286
R19829 DVSS.n4662 DVSS.n4577 0.00654286
R19830 DVSS.n254 DVSS.n253 0.0065
R19831 DVSS.n611 DVSS.n185 0.0065
R19832 DVSS.n577 DVSS.n576 0.0065
R19833 DVSS.n716 DVSS.n715 0.0065
R19834 DVSS.n3035 DVSS.n2693 0.0065
R19835 DVSS.n3512 DVSS.n3511 0.0065
R19836 DVSS.n3001 DVSS.n2696 0.0065
R19837 DVSS.n3287 DVSS.n3109 0.0065
R19838 DVSS.n363 DVSS.n362 0.0065
R19839 DVSS.n577 DVSS.n184 0.0065
R19840 DVSS.n715 DVSS.n155 0.0065
R19841 DVSS.n5741 DVSS.n47 0.0065
R19842 DVSS.n5741 DVSS.n40 0.0065
R19843 DVSS.n364 DVSS.n363 0.0065
R19844 DVSS.n5584 DVSS.n46 0.0065
R19845 DVSS.n611 DVSS.n203 0.0065
R19846 DVSS.n253 DVSS.n250 0.0065
R19847 DVSS.n5666 DVSS.n133 0.0065
R19848 DVSS.n5667 DVSS.n5666 0.0065
R19849 DVSS.n46 DVSS.n41 0.0065
R19850 DVSS.n4847 DVSS 0.00641429
R19851 VSS DVSS.n2267 0.00641429
R19852 DVSS.n2401 VSS 0.00641429
R19853 DVSS.n463 DVSS.n462 0.00640498
R19854 DVSS.n2228 DVSS.n2227 0.00635
R19855 DVSS.n3795 DVSS.n3794 0.00635
R19856 DVSS.n3787 DVSS.n3786 0.00635
R19857 DVSS.n3786 DVSS.n1662 0.00635
R19858 DVSS.n3206 DVSS.n3205 0.00626355
R19859 DVSS.n3346 DVSS.n3345 0.00626355
R19860 DVSS.n4094 DVSS.n1435 0.006125
R19861 DVSS.n3990 DVSS.n1428 0.006125
R19862 DVSS.n4182 DVSS.n1369 0.00609286
R19863 VSS DVSS.n2278 0.00609286
R19864 DVSS.n2643 VSS 0.00609286
R19865 DVSS.n4545 DVSS.n4511 0.00602857
R19866 DVSS.n4544 DVSS.n4540 0.00602857
R19867 DVSS.n4551 DVSS.n4509 0.00602857
R19868 DVSS.n2974 DVSS.n2973 0.006
R19869 DVSS.n3148 DVSS.n3147 0.006
R19870 DVSS.n2931 DVSS.n2722 0.006
R19871 DVSS.n3308 DVSS.n3307 0.006
R19872 DVSS.n4935 DVSS.n1179 0.0059878
R19873 DVSS.n4933 DVSS.n4931 0.0059878
R19874 DVSS.n4901 DVSS.n4900 0.00596429
R19875 DVSS.n4897 DVSS.n4775 0.00596429
R19876 DVSS.n4896 DVSS.n4778 0.00596429
R19877 DVSS.n4785 DVSS.n4784 0.00596429
R19878 DVSS.n4890 DVSS.n4889 0.00596429
R19879 DVSS.n4795 DVSS.n4786 0.00596429
R19880 DVSS.n4884 DVSS.n4796 0.00596429
R19881 DVSS DVSS.n3395 0.00585211
R19882 DVSS.n3859 DVSS.n3858 0.00583571
R19883 DVSS.n1709 DVSS.n1705 0.00575701
R19884 DVSS.n3875 DVSS.n3874 0.00570714
R19885 DVSS.n1858 DVSS.n1385 0.00561229
R19886 DVSS.n1389 DVSS.n1379 0.00561229
R19887 DVSS.n2968 DVSS 0.00559852
R19888 DVSS DVSS.n2925 0.00559852
R19889 DVSS.n3555 DVSS.n3554 0.00559852
R19890 DVSS.n5356 DVSS.n959 0.00559091
R19891 DVSS.n1913 DVSS.n1759 0.00551429
R19892 DVSS.n1909 DVSS.n1761 0.00551429
R19893 DVSS.n1882 DVSS.n1758 0.00551429
R19894 DVSS.n2919 DVSS.n2918 0.0055
R19895 DVSS.n3468 DVSS.n3170 0.0055
R19896 DVSS.n2922 DVSS.n2921 0.0055
R19897 DVSS.n3328 DVSS.n3172 0.0055
R19898 DVSS.n4851 DVSS.n4850 0.00548841
R19899 DVSS.n2653 DVSS.n2266 0.00548841
R19900 DVSS.n1536 DVSS.n1535 0.00548841
R19901 DVSS.n2399 DVSS.n2398 0.00548841
R19902 DVSS.n5106 DVSS.n1082 0.00548841
R19903 DVSS.n1980 DVSS.n1966 0.00538571
R19904 DVSS.n1975 DVSS.n1973 0.00538571
R19905 DVSS.n1977 DVSS.n1958 0.00538571
R19906 VSS DVSS.n2394 0.00538571
R19907 DVSS.n2992 DVSS.n2991 0.00537685
R19908 DVSS.n2998 DVSS.n2709 0.00537685
R19909 DVSS.n4789 DVSS.n4777 0.00532927
R19910 DVSS.n4888 DVSS.n4887 0.00532927
R19911 DVSS.n4758 DVSS.n4756 0.00532927
R19912 DVSS.n4918 DVSS.n1221 0.00532927
R19913 DVSS.n4716 DVSS.n1250 0.00532927
R19914 DVSS.n4733 DVSS.n4732 0.00532927
R19915 DVSS.n4615 DVSS.n1270 0.00532927
R19916 DVSS.n4693 DVSS.n4692 0.00532927
R19917 DVSS.n4596 DVSS.n4584 0.00532927
R19918 DVSS.n4640 DVSS.n4639 0.00532927
R19919 DVSS.n4565 DVSS.n4563 0.00532927
R19920 DVSS.n4670 DVSS.n4495 0.00532927
R19921 DVSS.n1735 DVSS.n1368 0.00519286
R19922 DVSS.n3771 DVSS.n3770 0.00519286
R19923 DVSS.n3937 DVSS.n3936 0.00519286
R19924 DVSS.n1853 DVSS.n1852 0.00514674
R19925 DVSS.n4929 DVSS.n4928 0.00505741
R19926 DVSS.n4928 DVSS.n961 0.00505741
R19927 DVSS.n958 DVSS.n956 0.00505741
R19928 DVSS.n1273 DVSS.n958 0.00505741
R19929 DVSS.n1936 DVSS.n1801 0.00504128
R19930 DVSS.n2183 DVSS.n1773 0.00504128
R19931 DVSS.n2858 DVSS.n2857 0.005
R19932 DVSS.n2864 DVSS.n2863 0.005
R19933 DVSS.n3445 DVSS.n3204 0.005
R19934 DVSS.n3220 DVSS.n3208 0.005
R19935 DVSS.n2827 DVSS.n2771 0.005
R19936 DVSS.n2867 DVSS.n2866 0.005
R19937 DVSS.n3351 DVSS.n3350 0.005
R19938 DVSS.n3356 DVSS.n3355 0.005
R19939 DVSS.n5731 DVSS.n5730 0.00498878
R19940 DVSS.n5357 DVSS.n5356 0.0049789
R19941 DVSS.n5356 DVSS.n5355 0.0049789
R19942 DVSS.n1739 DVSS.n1368 0.00493571
R19943 DVSS.n3770 DVSS.n1687 0.00493571
R19944 DVSS.n3937 DVSS.n1520 0.00493571
R19945 DVSS.n3184 DVSS.n3169 0.0049335
R19946 DVSS.n3330 DVSS.n3329 0.0049335
R19947 DVSS.n1847 DVSS.n1381 0.00489894
R19948 DVSS.n1843 DVSS.n1387 0.00489894
R19949 DVSS.n4193 DVSS.n1367 0.00476
R19950 DVSS.n4193 DVSS.n1365 0.00476
R19951 DVSS.n4197 DVSS.n1365 0.00476
R19952 DVSS.n4197 DVSS.n1363 0.00476
R19953 DVSS.n4201 DVSS.n1363 0.00476
R19954 DVSS.n4201 DVSS.n1361 0.00476
R19955 DVSS.n4206 DVSS.n1361 0.00476
R19956 DVSS.n4206 DVSS.n1359 0.00476
R19957 DVSS.n4210 DVSS.n1359 0.00476
R19958 DVSS.n4210 DVSS.n1357 0.00476
R19959 DVSS.n4215 DVSS.n1357 0.00476
R19960 DVSS.n4215 DVSS.n1355 0.00476
R19961 DVSS.n4219 DVSS.n1355 0.00476
R19962 DVSS.n4219 DVSS.n1353 0.00476
R19963 DVSS.n4223 DVSS.n1353 0.00476
R19964 DVSS.n4223 DVSS.n1351 0.00476
R19965 DVSS.n4227 DVSS.n1351 0.00476
R19966 DVSS.n4227 DVSS.n1349 0.00476
R19967 DVSS.n4231 DVSS.n1349 0.00476
R19968 DVSS.n4231 DVSS.n1347 0.00476
R19969 DVSS.n4235 DVSS.n1347 0.00476
R19970 DVSS.n4235 DVSS.n1345 0.00476
R19971 DVSS.n4240 DVSS.n1345 0.00476
R19972 DVSS.n4240 DVSS.n1343 0.00476
R19973 DVSS.n4244 DVSS.n1343 0.00476
R19974 DVSS.n4244 DVSS.n1341 0.00476
R19975 DVSS.n4248 DVSS.n1341 0.00476
R19976 DVSS.n4248 DVSS.n1339 0.00476
R19977 DVSS.n4252 DVSS.n1339 0.00476
R19978 DVSS.n4252 DVSS.n1337 0.00476
R19979 DVSS.n4256 DVSS.n1337 0.00476
R19980 DVSS.n4256 DVSS.n1335 0.00476
R19981 DVSS.n4260 DVSS.n1335 0.00476
R19982 DVSS.n4260 DVSS.n1333 0.00476
R19983 DVSS.n4264 DVSS.n1333 0.00476
R19984 DVSS.n4264 DVSS.n1331 0.00476
R19985 DVSS.n4268 DVSS.n1331 0.00476
R19986 DVSS.n4268 DVSS.n1329 0.00476
R19987 DVSS.n4272 DVSS.n1329 0.00476
R19988 DVSS.n4272 DVSS.n1327 0.00476
R19989 DVSS.n4276 DVSS.n1327 0.00476
R19990 DVSS.n4276 DVSS.n1325 0.00476
R19991 DVSS.n4280 DVSS.n1325 0.00476
R19992 DVSS.n4280 DVSS.n1323 0.00476
R19993 DVSS.n4284 DVSS.n1323 0.00476
R19994 DVSS.n4284 DVSS.n1321 0.00476
R19995 DVSS.n4288 DVSS.n1321 0.00476
R19996 DVSS.n4288 DVSS.n1319 0.00476
R19997 DVSS.n4421 DVSS.n1319 0.00476
R19998 DVSS.n4421 DVSS.n4420 0.00476
R19999 DVSS.n4420 DVSS.n4419 0.00476
R20000 DVSS.n4419 DVSS.n4294 0.00476
R20001 DVSS.n4415 DVSS.n4294 0.00476
R20002 DVSS.n4415 DVSS.n4414 0.00476
R20003 DVSS.n4414 DVSS.n4413 0.00476
R20004 DVSS.n4413 DVSS.n4300 0.00476
R20005 DVSS.n4373 DVSS.n4300 0.00476
R20006 DVSS.n4373 DVSS.n4372 0.00476
R20007 DVSS.n4372 DVSS.n4371 0.00476
R20008 DVSS.n4371 DVSS.n4306 0.00476
R20009 DVSS.n4367 DVSS.n4306 0.00476
R20010 DVSS.n4367 DVSS.n4366 0.00476
R20011 DVSS.n4366 DVSS.n4311 0.00476
R20012 DVSS.n4362 DVSS.n4311 0.00476
R20013 DVSS.n4362 DVSS.n4361 0.00476
R20014 DVSS.n4361 DVSS.n4360 0.00476
R20015 DVSS.n4360 DVSS.n4317 0.00476
R20016 DVSS.n4356 DVSS.n4317 0.00476
R20017 DVSS.n4356 DVSS.n4355 0.00476
R20018 DVSS.n4355 DVSS.n4354 0.00476
R20019 DVSS.n4354 DVSS.n4323 0.00476
R20020 DVSS.n4350 DVSS.n4323 0.00476
R20021 DVSS.n4350 DVSS.n4349 0.00476
R20022 DVSS.n4349 DVSS.n4348 0.00476
R20023 DVSS.n4348 DVSS.n4329 0.00476
R20024 DVSS.n4344 DVSS.n4329 0.00476
R20025 DVSS.n4344 DVSS.n4343 0.00476
R20026 DVSS.n4342 DVSS.n1175 0.00476
R20027 DVSS.n4939 DVSS.n1175 0.00476
R20028 DVSS.n4939 DVSS.n4938 0.00476
R20029 DVSS.n4194 DVSS.n1366 0.00476
R20030 DVSS.n4195 DVSS.n4194 0.00476
R20031 DVSS.n4196 DVSS.n4195 0.00476
R20032 DVSS.n4196 DVSS.n1362 0.00476
R20033 DVSS.n4202 DVSS.n1362 0.00476
R20034 DVSS.n4205 DVSS.n4204 0.00476
R20035 DVSS.n4205 DVSS.n1358 0.00476
R20036 DVSS.n4211 DVSS.n1358 0.00476
R20037 DVSS.n4212 DVSS.n4211 0.00476
R20038 DVSS.n4214 DVSS.n4212 0.00476
R20039 DVSS.n4214 DVSS.n4213 0.00476
R20040 DVSS.n4221 DVSS.n4220 0.00476
R20041 DVSS.n4222 DVSS.n4221 0.00476
R20042 DVSS.n4222 DVSS.n1350 0.00476
R20043 DVSS.n4228 DVSS.n1350 0.00476
R20044 DVSS.n4229 DVSS.n4228 0.00476
R20045 DVSS.n4230 DVSS.n4229 0.00476
R20046 DVSS.n4230 DVSS.n1346 0.00476
R20047 DVSS.n4236 DVSS.n1346 0.00476
R20048 DVSS.n4237 DVSS.n4236 0.00476
R20049 DVSS.n4239 DVSS.n1342 0.00476
R20050 DVSS.n4245 DVSS.n1342 0.00476
R20051 DVSS.n4246 DVSS.n4245 0.00476
R20052 DVSS.n4247 DVSS.n4246 0.00476
R20053 DVSS.n4247 DVSS.n1338 0.00476
R20054 DVSS.n4253 DVSS.n1338 0.00476
R20055 DVSS.n4254 DVSS.n4253 0.00476
R20056 DVSS.n4255 DVSS.n4254 0.00476
R20057 DVSS.n4255 DVSS.n1334 0.00476
R20058 DVSS.n4261 DVSS.n1334 0.00476
R20059 DVSS.n4262 DVSS.n4261 0.00476
R20060 DVSS.n4263 DVSS.n4262 0.00476
R20061 DVSS.n4263 DVSS.n1330 0.00476
R20062 DVSS.n4269 DVSS.n1330 0.00476
R20063 DVSS.n4270 DVSS.n4269 0.00476
R20064 DVSS.n4271 DVSS.n4270 0.00476
R20065 DVSS.n4271 DVSS.n1326 0.00476
R20066 DVSS.n4277 DVSS.n1326 0.00476
R20067 DVSS.n4278 DVSS.n4277 0.00476
R20068 DVSS.n4279 DVSS.n4278 0.00476
R20069 DVSS.n4279 DVSS.n1322 0.00476
R20070 DVSS.n4285 DVSS.n1322 0.00476
R20071 DVSS.n4286 DVSS.n4285 0.00476
R20072 DVSS.n4287 DVSS.n4286 0.00476
R20073 DVSS.n4287 DVSS.n1317 0.00476
R20074 DVSS.n4422 DVSS.n1318 0.00476
R20075 DVSS.n4418 DVSS.n1318 0.00476
R20076 DVSS.n4418 DVSS.n4417 0.00476
R20077 DVSS.n4417 DVSS.n4416 0.00476
R20078 DVSS.n4416 DVSS.n4295 0.00476
R20079 DVSS.n4412 DVSS.n4295 0.00476
R20080 DVSS.n4375 DVSS.n4374 0.00476
R20081 DVSS.n4374 DVSS.n4301 0.00476
R20082 DVSS.n4370 DVSS.n4301 0.00476
R20083 DVSS.n4370 DVSS.n4369 0.00476
R20084 DVSS.n4369 DVSS.n4368 0.00476
R20085 DVSS.n4365 DVSS.n4364 0.00476
R20086 DVSS.n4364 DVSS.n4363 0.00476
R20087 DVSS.n4363 DVSS.n4312 0.00476
R20088 DVSS.n4359 DVSS.n4312 0.00476
R20089 DVSS.n4359 DVSS.n4358 0.00476
R20090 DVSS.n4358 DVSS.n4357 0.00476
R20091 DVSS.n4357 DVSS.n4318 0.00476
R20092 DVSS.n4353 DVSS.n4318 0.00476
R20093 DVSS.n4353 DVSS.n4352 0.00476
R20094 DVSS.n4352 DVSS.n4351 0.00476
R20095 DVSS.n4351 DVSS.n4324 0.00476
R20096 DVSS.n4347 DVSS.n4324 0.00476
R20097 DVSS.n4347 DVSS.n4346 0.00476
R20098 DVSS.n4346 DVSS.n4345 0.00476
R20099 DVSS.n4345 DVSS.n4330 0.00476
R20100 DVSS.n4940 DVSS.n1174 0.00476
R20101 DVSS.n258 DVSS.n257 0.00476
R20102 DVSS.n313 DVSS.n312 0.00476
R20103 DVSS.n316 DVSS.n313 0.00476
R20104 DVSS.n317 DVSS.n316 0.00476
R20105 DVSS.n318 DVSS.n317 0.00476
R20106 DVSS.n319 DVSS.n318 0.00476
R20107 DVSS.n322 DVSS.n319 0.00476
R20108 DVSS.n323 DVSS.n322 0.00476
R20109 DVSS.n324 DVSS.n323 0.00476
R20110 DVSS.n325 DVSS.n324 0.00476
R20111 DVSS.n328 DVSS.n325 0.00476
R20112 DVSS.n329 DVSS.n328 0.00476
R20113 DVSS.n330 DVSS.n329 0.00476
R20114 DVSS.n331 DVSS.n330 0.00476
R20115 DVSS.n332 DVSS.n331 0.00476
R20116 DVSS.n332 DVSS.n193 0.00476
R20117 DVSS.n622 DVSS.n193 0.00476
R20118 DVSS.n628 DVSS.n189 0.00476
R20119 DVSS.n629 DVSS.n628 0.00476
R20120 DVSS.n630 DVSS.n629 0.00476
R20121 DVSS.n637 DVSS.n636 0.00476
R20122 DVSS.n638 DVSS.n637 0.00476
R20123 DVSS.n638 DVSS.n180 0.00476
R20124 DVSS.n644 DVSS.n180 0.00476
R20125 DVSS.n645 DVSS.n644 0.00476
R20126 DVSS.n646 DVSS.n645 0.00476
R20127 DVSS.n646 DVSS.n176 0.00476
R20128 DVSS.n652 DVSS.n176 0.00476
R20129 DVSS.n653 DVSS.n652 0.00476
R20130 DVSS.n654 DVSS.n653 0.00476
R20131 DVSS.n654 DVSS.n170 0.00476
R20132 DVSS.n686 DVSS.n171 0.00476
R20133 DVSS.n659 DVSS.n171 0.00476
R20134 DVSS.n660 DVSS.n659 0.00476
R20135 DVSS.n661 DVSS.n660 0.00476
R20136 DVSS.n664 DVSS.n661 0.00476
R20137 DVSS.n665 DVSS.n664 0.00476
R20138 DVSS.n666 DVSS.n665 0.00476
R20139 DVSS.n667 DVSS.n666 0.00476
R20140 DVSS.n669 DVSS.n667 0.00476
R20141 DVSS.n669 DVSS.n668 0.00476
R20142 DVSS.n668 DVSS.n132 0.00476
R20143 DVSS.n5674 DVSS.n127 0.00476
R20144 DVSS.n5675 DVSS.n5674 0.00476
R20145 DVSS.n5677 DVSS.n5675 0.00476
R20146 DVSS.n5677 DVSS.n5676 0.00476
R20147 DVSS.n5684 DVSS.n5683 0.00476
R20148 DVSS.n5685 DVSS.n5684 0.00476
R20149 DVSS.n5685 DVSS.n119 0.00476
R20150 DVSS.n5691 DVSS.n119 0.00476
R20151 DVSS.n5692 DVSS.n5691 0.00476
R20152 DVSS.n5693 DVSS.n5692 0.00476
R20153 DVSS.n5693 DVSS.n115 0.00476
R20154 DVSS.n5699 DVSS.n115 0.00476
R20155 DVSS.n5700 DVSS.n5699 0.00476
R20156 DVSS.n5701 DVSS.n5700 0.00476
R20157 DVSS.n5701 DVSS.n111 0.00476
R20158 DVSS.n5707 DVSS.n111 0.00476
R20159 DVSS.n5708 DVSS.n5707 0.00476
R20160 DVSS.n5709 DVSS.n5708 0.00476
R20161 DVSS.n5709 DVSS.n102 0.00476
R20162 DVSS.n5716 DVSS.n103 0.00476
R20163 DVSS.n5781 DVSS.n5780 0.00476
R20164 DVSS.n5782 DVSS.n5781 0.00476
R20165 DVSS.n5782 DVSS.n36 0.00476
R20166 DVSS.n5788 DVSS.n36 0.00476
R20167 DVSS.n5789 DVSS.n5788 0.00476
R20168 DVSS.n5790 DVSS.n5789 0.00476
R20169 DVSS.n5790 DVSS.n32 0.00476
R20170 DVSS.n5796 DVSS.n32 0.00476
R20171 DVSS.n5797 DVSS.n5796 0.00476
R20172 DVSS.n5798 DVSS.n5797 0.00476
R20173 DVSS.n5804 DVSS.n5803 0.00476
R20174 DVSS.n5805 DVSS.n5804 0.00476
R20175 DVSS.n5805 DVSS.n26 0.00476
R20176 DVSS.n424 DVSS.n244 0.00476
R20177 DVSS.n375 DVSS.n374 0.00476
R20178 DVSS.n376 DVSS.n375 0.00476
R20179 DVSS.n379 DVSS.n376 0.00476
R20180 DVSS.n380 DVSS.n379 0.00476
R20181 DVSS.n381 DVSS.n380 0.00476
R20182 DVSS.n382 DVSS.n381 0.00476
R20183 DVSS.n385 DVSS.n382 0.00476
R20184 DVSS.n386 DVSS.n385 0.00476
R20185 DVSS.n387 DVSS.n386 0.00476
R20186 DVSS.n388 DVSS.n387 0.00476
R20187 DVSS.n391 DVSS.n388 0.00476
R20188 DVSS.n392 DVSS.n391 0.00476
R20189 DVSS.n393 DVSS.n392 0.00476
R20190 DVSS.n394 DVSS.n393 0.00476
R20191 DVSS.n395 DVSS.n394 0.00476
R20192 DVSS.n395 DVSS.n195 0.00476
R20193 DVSS.n618 DVSS.n196 0.00476
R20194 DVSS.n201 DVSS.n196 0.00476
R20195 DVSS.n202 DVSS.n201 0.00476
R20196 DVSS.n581 DVSS.n578 0.00476
R20197 DVSS.n582 DVSS.n581 0.00476
R20198 DVSS.n583 DVSS.n582 0.00476
R20199 DVSS.n584 DVSS.n583 0.00476
R20200 DVSS.n587 DVSS.n584 0.00476
R20201 DVSS.n588 DVSS.n587 0.00476
R20202 DVSS.n589 DVSS.n588 0.00476
R20203 DVSS.n590 DVSS.n589 0.00476
R20204 DVSS.n592 DVSS.n590 0.00476
R20205 DVSS.n593 DVSS.n592 0.00476
R20206 DVSS.n593 DVSS.n168 0.00476
R20207 DVSS.n690 DVSS.n164 0.00476
R20208 DVSS.n696 DVSS.n164 0.00476
R20209 DVSS.n697 DVSS.n696 0.00476
R20210 DVSS.n698 DVSS.n697 0.00476
R20211 DVSS.n698 DVSS.n160 0.00476
R20212 DVSS.n704 DVSS.n160 0.00476
R20213 DVSS.n705 DVSS.n704 0.00476
R20214 DVSS.n706 DVSS.n705 0.00476
R20215 DVSS.n706 DVSS.n156 0.00476
R20216 DVSS.n713 DVSS.n156 0.00476
R20217 DVSS.n714 DVSS.n713 0.00476
R20218 DVSS.n138 DVSS.n135 0.00476
R20219 DVSS.n139 DVSS.n138 0.00476
R20220 DVSS.n140 DVSS.n139 0.00476
R20221 DVSS.n141 DVSS.n140 0.00476
R20222 DVSS.n5619 DVSS.n5618 0.00476
R20223 DVSS.n5620 DVSS.n5619 0.00476
R20224 DVSS.n5621 DVSS.n5620 0.00476
R20225 DVSS.n5624 DVSS.n5621 0.00476
R20226 DVSS.n5625 DVSS.n5624 0.00476
R20227 DVSS.n5626 DVSS.n5625 0.00476
R20228 DVSS.n5627 DVSS.n5626 0.00476
R20229 DVSS.n5630 DVSS.n5627 0.00476
R20230 DVSS.n5631 DVSS.n5630 0.00476
R20231 DVSS.n5632 DVSS.n5631 0.00476
R20232 DVSS.n5633 DVSS.n5632 0.00476
R20233 DVSS.n5635 DVSS.n5633 0.00476
R20234 DVSS.n5636 DVSS.n5635 0.00476
R20235 DVSS.n5636 DVSS.n53 0.00476
R20236 DVSS.n5733 DVSS.n53 0.00476
R20237 DVSS.n54 DVSS.n50 0.00476
R20238 DVSS.n5743 DVSS.n5742 0.00476
R20239 DVSS.n5744 DVSS.n5743 0.00476
R20240 DVSS.n5747 DVSS.n5744 0.00476
R20241 DVSS.n5748 DVSS.n5747 0.00476
R20242 DVSS.n5749 DVSS.n5748 0.00476
R20243 DVSS.n5750 DVSS.n5749 0.00476
R20244 DVSS.n5753 DVSS.n5750 0.00476
R20245 DVSS.n5754 DVSS.n5753 0.00476
R20246 DVSS.n5755 DVSS.n5754 0.00476
R20247 DVSS.n5757 DVSS.n5755 0.00476
R20248 DVSS.n5757 DVSS.n5756 0.00476
R20249 DVSS.n4 DVSS.n1 0.00476
R20250 DVSS.n5 DVSS.n4 0.00476
R20251 DVSS.n465 DVSS.n228 0.00476
R20252 DVSS.n471 DVSS.n224 0.00476
R20253 DVSS.n472 DVSS.n471 0.00476
R20254 DVSS.n473 DVSS.n472 0.00476
R20255 DVSS.n473 DVSS.n220 0.00476
R20256 DVSS.n479 DVSS.n220 0.00476
R20257 DVSS.n480 DVSS.n479 0.00476
R20258 DVSS.n481 DVSS.n480 0.00476
R20259 DVSS.n481 DVSS.n216 0.00476
R20260 DVSS.n487 DVSS.n216 0.00476
R20261 DVSS.n488 DVSS.n487 0.00476
R20262 DVSS.n489 DVSS.n488 0.00476
R20263 DVSS.n489 DVSS.n212 0.00476
R20264 DVSS.n495 DVSS.n212 0.00476
R20265 DVSS.n496 DVSS.n495 0.00476
R20266 DVSS.n498 DVSS.n496 0.00476
R20267 DVSS.n498 DVSS.n497 0.00476
R20268 DVSS.n506 DVSS.n505 0.00476
R20269 DVSS.n507 DVSS.n506 0.00476
R20270 DVSS.n507 DVSS.n204 0.00476
R20271 DVSS.n575 DVSS.n205 0.00476
R20272 DVSS.n513 DVSS.n205 0.00476
R20273 DVSS.n514 DVSS.n513 0.00476
R20274 DVSS.n515 DVSS.n514 0.00476
R20275 DVSS.n518 DVSS.n515 0.00476
R20276 DVSS.n519 DVSS.n518 0.00476
R20277 DVSS.n520 DVSS.n519 0.00476
R20278 DVSS.n521 DVSS.n520 0.00476
R20279 DVSS.n524 DVSS.n521 0.00476
R20280 DVSS.n525 DVSS.n524 0.00476
R20281 DVSS.n526 DVSS.n525 0.00476
R20282 DVSS.n530 DVSS.n527 0.00476
R20283 DVSS.n531 DVSS.n530 0.00476
R20284 DVSS.n532 DVSS.n531 0.00476
R20285 DVSS.n533 DVSS.n532 0.00476
R20286 DVSS.n536 DVSS.n533 0.00476
R20287 DVSS.n537 DVSS.n536 0.00476
R20288 DVSS.n538 DVSS.n537 0.00476
R20289 DVSS.n539 DVSS.n538 0.00476
R20290 DVSS.n540 DVSS.n539 0.00476
R20291 DVSS.n540 DVSS.n154 0.00476
R20292 DVSS.n717 DVSS.n154 0.00476
R20293 DVSS.n724 DVSS.n150 0.00476
R20294 DVSS.n725 DVSS.n724 0.00476
R20295 DVSS.n726 DVSS.n725 0.00476
R20296 DVSS.n726 DVSS.n144 0.00476
R20297 DVSS.n5614 DVSS.n145 0.00476
R20298 DVSS.n731 DVSS.n145 0.00476
R20299 DVSS.n732 DVSS.n731 0.00476
R20300 DVSS.n733 DVSS.n732 0.00476
R20301 DVSS.n736 DVSS.n733 0.00476
R20302 DVSS.n737 DVSS.n736 0.00476
R20303 DVSS.n738 DVSS.n737 0.00476
R20304 DVSS.n739 DVSS.n738 0.00476
R20305 DVSS.n742 DVSS.n739 0.00476
R20306 DVSS.n743 DVSS.n742 0.00476
R20307 DVSS.n744 DVSS.n743 0.00476
R20308 DVSS.n745 DVSS.n744 0.00476
R20309 DVSS.n748 DVSS.n745 0.00476
R20310 DVSS.n749 DVSS.n748 0.00476
R20311 DVSS.n750 DVSS.n749 0.00476
R20312 DVSS.n753 DVSS.n751 0.00476
R20313 DVSS.n809 DVSS.n806 0.00476
R20314 DVSS.n810 DVSS.n809 0.00476
R20315 DVSS.n811 DVSS.n810 0.00476
R20316 DVSS.n812 DVSS.n811 0.00476
R20317 DVSS.n815 DVSS.n812 0.00476
R20318 DVSS.n816 DVSS.n815 0.00476
R20319 DVSS.n817 DVSS.n816 0.00476
R20320 DVSS.n818 DVSS.n817 0.00476
R20321 DVSS.n821 DVSS.n818 0.00476
R20322 DVSS.n822 DVSS.n821 0.00476
R20323 DVSS.n824 DVSS.n823 0.00476
R20324 DVSS.n827 DVSS.n824 0.00476
R20325 DVSS.n828 DVSS.n827 0.00476
R20326 DVSS.n367 DVSS.n227 0.00476
R20327 DVSS.n466 DVSS.n227 0.00476
R20328 DVSS.n466 DVSS.n225 0.00476
R20329 DVSS.n470 DVSS.n225 0.00476
R20330 DVSS.n470 DVSS.n223 0.00476
R20331 DVSS.n474 DVSS.n223 0.00476
R20332 DVSS.n474 DVSS.n221 0.00476
R20333 DVSS.n478 DVSS.n221 0.00476
R20334 DVSS.n478 DVSS.n219 0.00476
R20335 DVSS.n482 DVSS.n219 0.00476
R20336 DVSS.n482 DVSS.n217 0.00476
R20337 DVSS.n486 DVSS.n217 0.00476
R20338 DVSS.n486 DVSS.n215 0.00476
R20339 DVSS.n490 DVSS.n215 0.00476
R20340 DVSS.n490 DVSS.n213 0.00476
R20341 DVSS.n494 DVSS.n213 0.00476
R20342 DVSS.n494 DVSS.n211 0.00476
R20343 DVSS.n499 DVSS.n211 0.00476
R20344 DVSS.n499 DVSS.n209 0.00476
R20345 DVSS.n504 DVSS.n209 0.00476
R20346 DVSS.n504 DVSS.n208 0.00476
R20347 DVSS.n508 DVSS.n208 0.00476
R20348 DVSS.n509 DVSS.n508 0.00476
R20349 DVSS.n574 DVSS.n206 0.00476
R20350 DVSS.n570 DVSS.n206 0.00476
R20351 DVSS.n570 DVSS.n569 0.00476
R20352 DVSS.n569 DVSS.n568 0.00476
R20353 DVSS.n568 DVSS.n516 0.00476
R20354 DVSS.n564 DVSS.n516 0.00476
R20355 DVSS.n564 DVSS.n563 0.00476
R20356 DVSS.n563 DVSS.n562 0.00476
R20357 DVSS.n562 DVSS.n522 0.00476
R20358 DVSS.n558 DVSS.n522 0.00476
R20359 DVSS.n558 DVSS.n557 0.00476
R20360 DVSS.n557 DVSS.n556 0.00476
R20361 DVSS.n556 DVSS.n528 0.00476
R20362 DVSS.n552 DVSS.n528 0.00476
R20363 DVSS.n552 DVSS.n551 0.00476
R20364 DVSS.n551 DVSS.n550 0.00476
R20365 DVSS.n550 DVSS.n534 0.00476
R20366 DVSS.n546 DVSS.n534 0.00476
R20367 DVSS.n546 DVSS.n545 0.00476
R20368 DVSS.n545 DVSS.n544 0.00476
R20369 DVSS.n544 DVSS.n541 0.00476
R20370 DVSS.n541 DVSS.n153 0.00476
R20371 DVSS.n718 DVSS.n153 0.00476
R20372 DVSS.n723 DVSS.n151 0.00476
R20373 DVSS.n723 DVSS.n149 0.00476
R20374 DVSS.n727 DVSS.n149 0.00476
R20375 DVSS.n727 DVSS.n146 0.00476
R20376 DVSS.n5613 DVSS.n146 0.00476
R20377 DVSS.n5613 DVSS.n147 0.00476
R20378 DVSS.n5609 DVSS.n147 0.00476
R20379 DVSS.n5609 DVSS.n5608 0.00476
R20380 DVSS.n5608 DVSS.n5607 0.00476
R20381 DVSS.n5607 DVSS.n734 0.00476
R20382 DVSS.n5603 DVSS.n734 0.00476
R20383 DVSS.n5603 DVSS.n5602 0.00476
R20384 DVSS.n5602 DVSS.n5601 0.00476
R20385 DVSS.n5601 DVSS.n740 0.00476
R20386 DVSS.n5597 DVSS.n740 0.00476
R20387 DVSS.n5597 DVSS.n5596 0.00476
R20388 DVSS.n5596 DVSS.n5595 0.00476
R20389 DVSS.n5595 DVSS.n746 0.00476
R20390 DVSS.n5591 DVSS.n746 0.00476
R20391 DVSS.n5591 DVSS.n5590 0.00476
R20392 DVSS.n5590 DVSS.n5589 0.00476
R20393 DVSS.n5589 DVSS.n752 0.00476
R20394 DVSS.n5585 DVSS.n752 0.00476
R20395 DVSS.n5583 DVSS.n807 0.00476
R20396 DVSS.n5579 DVSS.n807 0.00476
R20397 DVSS.n5579 DVSS.n5578 0.00476
R20398 DVSS.n5578 DVSS.n5577 0.00476
R20399 DVSS.n5577 DVSS.n813 0.00476
R20400 DVSS.n5573 DVSS.n813 0.00476
R20401 DVSS.n5573 DVSS.n5572 0.00476
R20402 DVSS.n5572 DVSS.n5571 0.00476
R20403 DVSS.n5571 DVSS.n819 0.00476
R20404 DVSS.n5567 DVSS.n819 0.00476
R20405 DVSS.n5566 DVSS.n5565 0.00476
R20406 DVSS.n5565 DVSS.n825 0.00476
R20407 DVSS.n826 DVSS.n825 0.00476
R20408 DVSS.n423 DVSS.n245 0.00476
R20409 DVSS.n423 DVSS.n246 0.00476
R20410 DVSS.n419 DVSS.n246 0.00476
R20411 DVSS.n419 DVSS.n418 0.00476
R20412 DVSS.n418 DVSS.n417 0.00476
R20413 DVSS.n417 DVSS.n377 0.00476
R20414 DVSS.n413 DVSS.n377 0.00476
R20415 DVSS.n413 DVSS.n412 0.00476
R20416 DVSS.n412 DVSS.n411 0.00476
R20417 DVSS.n411 DVSS.n383 0.00476
R20418 DVSS.n407 DVSS.n383 0.00476
R20419 DVSS.n407 DVSS.n406 0.00476
R20420 DVSS.n406 DVSS.n405 0.00476
R20421 DVSS.n405 DVSS.n389 0.00476
R20422 DVSS.n401 DVSS.n389 0.00476
R20423 DVSS.n401 DVSS.n400 0.00476
R20424 DVSS.n400 DVSS.n399 0.00476
R20425 DVSS.n399 DVSS.n396 0.00476
R20426 DVSS.n396 DVSS.n197 0.00476
R20427 DVSS.n617 DVSS.n197 0.00476
R20428 DVSS.n617 DVSS.n198 0.00476
R20429 DVSS.n613 DVSS.n198 0.00476
R20430 DVSS.n613 DVSS.n612 0.00476
R20431 DVSS.n610 DVSS.n579 0.00476
R20432 DVSS.n606 DVSS.n579 0.00476
R20433 DVSS.n606 DVSS.n605 0.00476
R20434 DVSS.n605 DVSS.n604 0.00476
R20435 DVSS.n604 DVSS.n585 0.00476
R20436 DVSS.n600 DVSS.n585 0.00476
R20437 DVSS.n600 DVSS.n599 0.00476
R20438 DVSS.n599 DVSS.n598 0.00476
R20439 DVSS.n598 DVSS.n591 0.00476
R20440 DVSS.n594 DVSS.n591 0.00476
R20441 DVSS.n594 DVSS.n167 0.00476
R20442 DVSS.n691 DVSS.n167 0.00476
R20443 DVSS.n691 DVSS.n165 0.00476
R20444 DVSS.n695 DVSS.n165 0.00476
R20445 DVSS.n695 DVSS.n163 0.00476
R20446 DVSS.n699 DVSS.n163 0.00476
R20447 DVSS.n699 DVSS.n161 0.00476
R20448 DVSS.n703 DVSS.n161 0.00476
R20449 DVSS.n703 DVSS.n159 0.00476
R20450 DVSS.n707 DVSS.n159 0.00476
R20451 DVSS.n707 DVSS.n157 0.00476
R20452 DVSS.n712 DVSS.n157 0.00476
R20453 DVSS.n712 DVSS.n134 0.00476
R20454 DVSS.n5665 DVSS.n136 0.00476
R20455 DVSS.n5661 DVSS.n136 0.00476
R20456 DVSS.n5661 DVSS.n5660 0.00476
R20457 DVSS.n5660 DVSS.n5659 0.00476
R20458 DVSS.n5659 DVSS.n142 0.00476
R20459 DVSS.n5655 DVSS.n142 0.00476
R20460 DVSS.n5655 DVSS.n5654 0.00476
R20461 DVSS.n5654 DVSS.n5653 0.00476
R20462 DVSS.n5653 DVSS.n5622 0.00476
R20463 DVSS.n5649 DVSS.n5622 0.00476
R20464 DVSS.n5649 DVSS.n5648 0.00476
R20465 DVSS.n5648 DVSS.n5647 0.00476
R20466 DVSS.n5647 DVSS.n5628 0.00476
R20467 DVSS.n5643 DVSS.n5628 0.00476
R20468 DVSS.n5643 DVSS.n5642 0.00476
R20469 DVSS.n5642 DVSS.n5641 0.00476
R20470 DVSS.n5641 DVSS.n5634 0.00476
R20471 DVSS.n5637 DVSS.n5634 0.00476
R20472 DVSS.n5637 DVSS.n52 0.00476
R20473 DVSS.n5734 DVSS.n52 0.00476
R20474 DVSS.n5734 DVSS.n49 0.00476
R20475 DVSS.n5738 DVSS.n49 0.00476
R20476 DVSS.n5739 DVSS.n5738 0.00476
R20477 DVSS.n5774 DVSS.n5773 0.00476
R20478 DVSS.n5773 DVSS.n5772 0.00476
R20479 DVSS.n5772 DVSS.n5745 0.00476
R20480 DVSS.n5768 DVSS.n5745 0.00476
R20481 DVSS.n5768 DVSS.n5767 0.00476
R20482 DVSS.n5767 DVSS.n5766 0.00476
R20483 DVSS.n5766 DVSS.n5751 0.00476
R20484 DVSS.n5762 DVSS.n5751 0.00476
R20485 DVSS.n5762 DVSS.n5761 0.00476
R20486 DVSS.n5761 DVSS.n5760 0.00476
R20487 DVSS.n5760 DVSS.n0 0.00476
R20488 DVSS.n5817 DVSS.n2 0.00476
R20489 DVSS.n3 DVSS.n2 0.00476
R20490 DVSS.n360 DVSS.n255 0.00476
R20491 DVSS.n356 DVSS.n255 0.00476
R20492 DVSS.n356 DVSS.n355 0.00476
R20493 DVSS.n355 DVSS.n354 0.00476
R20494 DVSS.n354 DVSS.n314 0.00476
R20495 DVSS.n350 DVSS.n314 0.00476
R20496 DVSS.n350 DVSS.n349 0.00476
R20497 DVSS.n349 DVSS.n348 0.00476
R20498 DVSS.n348 DVSS.n320 0.00476
R20499 DVSS.n344 DVSS.n320 0.00476
R20500 DVSS.n344 DVSS.n343 0.00476
R20501 DVSS.n343 DVSS.n342 0.00476
R20502 DVSS.n342 DVSS.n326 0.00476
R20503 DVSS.n338 DVSS.n326 0.00476
R20504 DVSS.n338 DVSS.n337 0.00476
R20505 DVSS.n337 DVSS.n336 0.00476
R20506 DVSS.n336 DVSS.n333 0.00476
R20507 DVSS.n333 DVSS.n192 0.00476
R20508 DVSS.n623 DVSS.n192 0.00476
R20509 DVSS.n623 DVSS.n190 0.00476
R20510 DVSS.n627 DVSS.n190 0.00476
R20511 DVSS.n627 DVSS.n188 0.00476
R20512 DVSS.n631 DVSS.n188 0.00476
R20513 DVSS.n635 DVSS.n183 0.00476
R20514 DVSS.n639 DVSS.n183 0.00476
R20515 DVSS.n639 DVSS.n181 0.00476
R20516 DVSS.n643 DVSS.n181 0.00476
R20517 DVSS.n643 DVSS.n179 0.00476
R20518 DVSS.n647 DVSS.n179 0.00476
R20519 DVSS.n647 DVSS.n177 0.00476
R20520 DVSS.n651 DVSS.n177 0.00476
R20521 DVSS.n651 DVSS.n175 0.00476
R20522 DVSS.n655 DVSS.n175 0.00476
R20523 DVSS.n655 DVSS.n172 0.00476
R20524 DVSS.n685 DVSS.n172 0.00476
R20525 DVSS.n685 DVSS.n173 0.00476
R20526 DVSS.n681 DVSS.n173 0.00476
R20527 DVSS.n681 DVSS.n680 0.00476
R20528 DVSS.n680 DVSS.n679 0.00476
R20529 DVSS.n679 DVSS.n662 0.00476
R20530 DVSS.n675 DVSS.n662 0.00476
R20531 DVSS.n675 DVSS.n674 0.00476
R20532 DVSS.n674 DVSS.n673 0.00476
R20533 DVSS.n673 DVSS.n670 0.00476
R20534 DVSS.n670 DVSS.n131 0.00476
R20535 DVSS.n5668 DVSS.n131 0.00476
R20536 DVSS.n5673 DVSS.n128 0.00476
R20537 DVSS.n5673 DVSS.n126 0.00476
R20538 DVSS.n5678 DVSS.n126 0.00476
R20539 DVSS.n5678 DVSS.n124 0.00476
R20540 DVSS.n5682 DVSS.n124 0.00476
R20541 DVSS.n5682 DVSS.n122 0.00476
R20542 DVSS.n5686 DVSS.n122 0.00476
R20543 DVSS.n5686 DVSS.n120 0.00476
R20544 DVSS.n5690 DVSS.n120 0.00476
R20545 DVSS.n5690 DVSS.n118 0.00476
R20546 DVSS.n5694 DVSS.n118 0.00476
R20547 DVSS.n5694 DVSS.n116 0.00476
R20548 DVSS.n5698 DVSS.n116 0.00476
R20549 DVSS.n5698 DVSS.n114 0.00476
R20550 DVSS.n5702 DVSS.n114 0.00476
R20551 DVSS.n5702 DVSS.n112 0.00476
R20552 DVSS.n5706 DVSS.n112 0.00476
R20553 DVSS.n5706 DVSS.n110 0.00476
R20554 DVSS.n5710 DVSS.n110 0.00476
R20555 DVSS.n5710 DVSS.n104 0.00476
R20556 DVSS.n5715 DVSS.n104 0.00476
R20557 DVSS.n5715 DVSS.n108 0.00476
R20558 DVSS.n108 DVSS.n107 0.00476
R20559 DVSS.n5779 DVSS.n39 0.00476
R20560 DVSS.n5783 DVSS.n39 0.00476
R20561 DVSS.n5783 DVSS.n37 0.00476
R20562 DVSS.n5787 DVSS.n37 0.00476
R20563 DVSS.n5787 DVSS.n35 0.00476
R20564 DVSS.n5791 DVSS.n35 0.00476
R20565 DVSS.n5791 DVSS.n33 0.00476
R20566 DVSS.n5795 DVSS.n33 0.00476
R20567 DVSS.n5795 DVSS.n31 0.00476
R20568 DVSS.n5799 DVSS.n31 0.00476
R20569 DVSS.n5802 DVSS.n29 0.00476
R20570 DVSS.n5806 DVSS.n29 0.00476
R20571 DVSS.n5806 DVSS.n27 0.00476
R20572 DVSS.n3998 DVSS.n1432 0.00465761
R20573 DVSS.n3997 DVSS.n1429 0.00465761
R20574 DVSS.n1981 DVSS.n1980 0.00461429
R20575 DVSS.n1975 DVSS.n1960 0.00461429
R20576 DVSS.n1977 DVSS.n1961 0.00461429
R20577 DVSS.n5729 DVSS.n57 0.00461371
R20578 DVSS.n5798 DVSS 0.00458
R20579 DVSS.n5799 DVSS 0.00458
R20580 DVSS.n272 DVSS.n242 0.0045724
R20581 DVSS.n511 DVSS.n186 0.0045
R20582 DVSS.n720 DVSS.n129 0.0045
R20583 DVSS.n370 DVSS.n247 0.0045
R20584 DVSS.n633 DVSS.n186 0.0045
R20585 DVSS.n5670 DVSS.n129 0.0045
R20586 DVSS.n5776 DVSS.n43 0.0045
R20587 DVSS.n5777 DVSS.n5776 0.0045
R20588 DVSS.n370 DVSS.n369 0.0045
R20589 DVSS.n2815 DVSS.n2787 0.0045
R20590 DVSS.n2914 DVSS.n2747 0.0045
R20591 DVSS.n3461 DVSS.n3182 0.0045
R20592 DVSS.n3424 DVSS.n3423 0.0045
R20593 DVSS.n2798 DVSS.n2785 0.0045
R20594 DVSS.n2875 DVSS.n2874 0.0045
R20595 DVSS.n3333 DVSS.n3180 0.0045
R20596 DVSS.n3244 DVSS.n3235 0.0045
R20597 DVSS.n1913 DVSS.n1884 0.00448571
R20598 DVSS.n1909 DVSS.n1908 0.00448571
R20599 DVSS.n1882 DVSS.n1762 0.00448571
R20600 DVSS.n3876 DVSS.n3875 0.00442143
R20601 DVSS.n273 DVSS.n241 0.0044172
R20602 DVSS.n361 DVSS.n252 0.00434
R20603 DVSS.n425 DVSS.n243 0.00434
R20604 DVSS.n366 DVSS.n365 0.00434
R20605 DVSS.n1900 DVSS.n1749 0.004325
R20606 DVSS.n1889 DVSS.n1750 0.004325
R20607 DVSS.n3858 DVSS.n3855 0.00429286
R20608 DVSS.n4793 DVSS.n4792 0.00428827
R20609 DVSS.n4921 DVSS.n1218 0.00428827
R20610 DVSS.n4719 DVSS.n4718 0.00428827
R20611 DVSS.n4680 DVSS.n4679 0.00428827
R20612 DVSS.n4600 DVSS.n4599 0.00428827
R20613 DVSS.n4673 DVSS.n4492 0.00428827
R20614 DVSS.n621 DVSS.n189 0.00425
R20615 DVSS.n619 DVSS.n618 0.00425
R20616 DVSS.n505 DVSS.n194 0.00425
R20617 DVSS.n5813 DVSS.n6 0.00422
R20618 DVSS.n5561 DVSS.n829 0.00422
R20619 DVSS.n4423 DVSS.n1317 0.00419
R20620 DVSS.n4941 DVSS.n1173 0.00419
R20621 DVSS.n1851 DVSS.n1382 0.0041856
R20622 DVSS.n1840 DVSS.n1388 0.0041856
R20623 DVSS.n4900 DVSS.n4775 0.00416429
R20624 DVSS.n4897 DVSS.n4896 0.00416429
R20625 DVSS.n4784 DVSS.n4778 0.00416429
R20626 DVSS.n4890 DVSS.n4785 0.00416429
R20627 DVSS.n4889 DVSS.n4786 0.00416429
R20628 DVSS.n4796 DVSS.n4795 0.00416429
R20629 DVSS.n4884 DVSS.n4883 0.00416429
R20630 DVSS.n4545 DVSS.n4544 0.0041
R20631 DVSS.n4540 DVSS.n4509 0.0041
R20632 DVSS.n4203 DVSS.n4202 0.00407
R20633 DVSS.n4220 DVSS.n1354 0.00407
R20634 DVSS.n3037 DVSS.n2692 0.0040468
R20635 DVSS.n3000 DVSS.n2688 0.0040468
R20636 DVSS.n5780 DVSS.n40 0.00404
R20637 DVSS.n5742 DVSS.n5741 0.00404
R20638 DVSS.n806 DVSS.n47 0.00404
R20639 DVSS.n5584 DVSS.n5583 0.00404
R20640 DVSS.n5774 DVSS.n46 0.00404
R20641 DVSS.n5779 DVSS.n41 0.00404
R20642 DVSS.n4179 DVSS.n1369 0.00403571
R20643 DVSS.n2969 DVSS.n2724 0.004
R20644 DVSS.n3152 DVSS.n3149 0.004
R20645 DVSS.n2936 DVSS.n2935 0.004
R20646 DVSS.n3314 DVSS.n3312 0.004
R20647 DVSS.n4411 DVSS.n4375 0.00395
R20648 DVSS.n4340 DVSS.n1173 0.00395
R20649 DVSS.n5683 DVSS.n123 0.00395
R20650 DVSS.n5618 DVSS.n5617 0.00395
R20651 DVSS.n5615 DVSS.n5614 0.00395
R20652 DVSS.n1982 DVSS.n1943 0.00393049
R20653 DVSS.n1959 DVSS.n1944 0.00393049
R20654 DVSS.n2196 DVSS.n1754 0.00393049
R20655 DVSS.n2199 DVSS.n2198 0.00393049
R20656 DVSS.n4343 DVSS 0.00392
R20657 DVSS DVSS.n4330 0.00392
R20658 DVSS DVSS.n822 0.00392
R20659 DVSS.n5567 DVSS 0.00392
R20660 DVSS.n5728 DVSS.n5727 0.00391137
R20661 DVSS.n5718 DVSS.n101 0.00386658
R20662 DVSS.n4794 DVSS.n4793 0.00382908
R20663 DVSS.n4921 DVSS.n4920 0.00382908
R20664 DVSS.n4718 DVSS.n1241 0.00382908
R20665 DVSS.n4679 DVSS.n1262 0.00382908
R20666 DVSS.n4601 DVSS.n4600 0.00382908
R20667 DVSS.n4673 DVSS.n4672 0.00382908
R20668 DVSS.n4239 DVSS.n4238 0.0038
R20669 DVSS.n155 DVSS.n127 0.0038
R20670 DVSS.n715 DVSS.n135 0.0038
R20671 DVSS.n716 DVSS.n150 0.0038
R20672 DVSS.n151 DVSS.n133 0.0038
R20673 DVSS.n5666 DVSS.n5665 0.0038
R20674 DVSS.n5667 DVSS.n128 0.0038
R20675 DVSS.n3794 DVSS.n1653 0.00377857
R20676 DVSS.n3787 DVSS.n1661 0.00377857
R20677 DVSS.n1681 DVSS.n1662 0.00377857
R20678 DVSS.n276 DVSS.n274 0.00374841
R20679 DVSS.n3954 DVSS.n1500 0.00362245
R20680 DVSS.n3484 DVSS.n3483 0.00360345
R20681 DVSS.n3311 DVSS.n3247 0.00360345
R20682 DVSS.n5717 DVSS.n102 0.00359
R20683 DVSS.n5733 DVSS.n5732 0.00359
R20684 DVSS.n801 DVSS.n750 0.00359
R20685 DVSS.n4560 DVSS.n4504 0.00358571
R20686 DVSS.n4559 DVSS.n4505 0.00358571
R20687 DVSS.n4566 DVSS.n4502 0.00358571
R20688 DVSS.n4568 DVSS.n4567 0.00358571
R20689 DVSS.n4669 DVSS.n4496 0.00358571
R20690 DVSS.n4668 DVSS.n4497 0.00358571
R20691 DVSS.n4577 DVSS.n4574 0.00358571
R20692 DVSS.n636 DVSS.n184 0.00356
R20693 DVSS.n578 DVSS.n577 0.00356
R20694 DVSS.n576 DVSS.n575 0.00356
R20695 DVSS.n574 DVSS.n203 0.00356
R20696 DVSS.n611 DVSS.n610 0.00356
R20697 DVSS.n635 DVSS.n185 0.00356
R20698 DVSS.n310 DVSS.n259 0.0035543
R20699 DVSS DVSS.n1 0.00353
R20700 DVSS DVSS.n5817 0.00353
R20701 DVSS.n3013 DVSS.n2703 0.0035
R20702 DVSS.n3507 DVSS.n3506 0.0035
R20703 DVSS.n3005 DVSS.n2708 0.0035
R20704 DVSS.n3291 DVSS.n3118 0.0035
R20705 DVSS.n803 DVSS.n802 0.00341771
R20706 DVSS.n2125 DVSS.n1951 0.00338991
R20707 DVSS.n5809 DVSS.n26 0.0033824
R20708 DVSS.n4936 DVSS.n1174 0.00338166
R20709 DVSS.n359 DVSS.n358 0.00334
R20710 DVSS.n358 DVSS.n357 0.00334
R20711 DVSS.n357 DVSS.n256 0.00334
R20712 DVSS.n353 DVSS.n256 0.00334
R20713 DVSS.n353 DVSS.n352 0.00334
R20714 DVSS.n352 DVSS.n351 0.00334
R20715 DVSS.n351 DVSS.n315 0.00334
R20716 DVSS.n347 DVSS.n315 0.00334
R20717 DVSS.n347 DVSS.n346 0.00334
R20718 DVSS.n346 DVSS.n345 0.00334
R20719 DVSS.n345 DVSS.n321 0.00334
R20720 DVSS.n341 DVSS.n321 0.00334
R20721 DVSS.n341 DVSS.n340 0.00334
R20722 DVSS.n340 DVSS.n339 0.00334
R20723 DVSS.n339 DVSS.n327 0.00334
R20724 DVSS.n335 DVSS.n327 0.00334
R20725 DVSS.n335 DVSS.n334 0.00334
R20726 DVSS.n334 DVSS.n191 0.00334
R20727 DVSS.n624 DVSS.n191 0.00334
R20728 DVSS.n625 DVSS.n624 0.00334
R20729 DVSS.n626 DVSS.n625 0.00334
R20730 DVSS.n626 DVSS.n187 0.00334
R20731 DVSS.n632 DVSS.n187 0.00334
R20732 DVSS.n634 DVSS.n182 0.00334
R20733 DVSS.n640 DVSS.n182 0.00334
R20734 DVSS.n641 DVSS.n640 0.00334
R20735 DVSS.n642 DVSS.n641 0.00334
R20736 DVSS.n642 DVSS.n178 0.00334
R20737 DVSS.n648 DVSS.n178 0.00334
R20738 DVSS.n649 DVSS.n648 0.00334
R20739 DVSS.n650 DVSS.n649 0.00334
R20740 DVSS.n650 DVSS.n174 0.00334
R20741 DVSS.n656 DVSS.n174 0.00334
R20742 DVSS.n657 DVSS.n656 0.00334
R20743 DVSS.n684 DVSS.n657 0.00334
R20744 DVSS.n684 DVSS.n683 0.00334
R20745 DVSS.n683 DVSS.n682 0.00334
R20746 DVSS.n682 DVSS.n658 0.00334
R20747 DVSS.n678 DVSS.n658 0.00334
R20748 DVSS.n678 DVSS.n677 0.00334
R20749 DVSS.n677 DVSS.n676 0.00334
R20750 DVSS.n676 DVSS.n663 0.00334
R20751 DVSS.n672 DVSS.n663 0.00334
R20752 DVSS.n672 DVSS.n671 0.00334
R20753 DVSS.n671 DVSS.n130 0.00334
R20754 DVSS.n5669 DVSS.n130 0.00334
R20755 DVSS.n5672 DVSS.n5671 0.00334
R20756 DVSS.n5672 DVSS.n125 0.00334
R20757 DVSS.n5679 DVSS.n125 0.00334
R20758 DVSS.n5680 DVSS.n5679 0.00334
R20759 DVSS.n5681 DVSS.n5680 0.00334
R20760 DVSS.n5681 DVSS.n121 0.00334
R20761 DVSS.n5687 DVSS.n121 0.00334
R20762 DVSS.n5688 DVSS.n5687 0.00334
R20763 DVSS.n5689 DVSS.n5688 0.00334
R20764 DVSS.n5689 DVSS.n117 0.00334
R20765 DVSS.n5695 DVSS.n117 0.00334
R20766 DVSS.n5696 DVSS.n5695 0.00334
R20767 DVSS.n5697 DVSS.n5696 0.00334
R20768 DVSS.n5697 DVSS.n113 0.00334
R20769 DVSS.n5703 DVSS.n113 0.00334
R20770 DVSS.n5704 DVSS.n5703 0.00334
R20771 DVSS.n5705 DVSS.n5704 0.00334
R20772 DVSS.n5705 DVSS.n109 0.00334
R20773 DVSS.n5711 DVSS.n109 0.00334
R20774 DVSS.n5712 DVSS.n5711 0.00334
R20775 DVSS.n5714 DVSS.n5712 0.00334
R20776 DVSS.n5714 DVSS.n5713 0.00334
R20777 DVSS.n5713 DVSS.n42 0.00334
R20778 DVSS.n5778 DVSS.n38 0.00334
R20779 DVSS.n5784 DVSS.n38 0.00334
R20780 DVSS.n5785 DVSS.n5784 0.00334
R20781 DVSS.n5786 DVSS.n5785 0.00334
R20782 DVSS.n5786 DVSS.n34 0.00334
R20783 DVSS.n5792 DVSS.n34 0.00334
R20784 DVSS.n5793 DVSS.n5792 0.00334
R20785 DVSS.n5794 DVSS.n5793 0.00334
R20786 DVSS.n5794 DVSS.n30 0.00334
R20787 DVSS.n5800 DVSS.n30 0.00334
R20788 DVSS.n5801 DVSS.n5800 0.00334
R20789 DVSS.n5807 DVSS.n28 0.00334
R20790 DVSS.n422 DVSS.n371 0.00334
R20791 DVSS.n422 DVSS.n421 0.00334
R20792 DVSS.n421 DVSS.n420 0.00334
R20793 DVSS.n420 DVSS.n372 0.00334
R20794 DVSS.n416 DVSS.n372 0.00334
R20795 DVSS.n416 DVSS.n415 0.00334
R20796 DVSS.n415 DVSS.n414 0.00334
R20797 DVSS.n414 DVSS.n378 0.00334
R20798 DVSS.n410 DVSS.n378 0.00334
R20799 DVSS.n410 DVSS.n409 0.00334
R20800 DVSS.n409 DVSS.n408 0.00334
R20801 DVSS.n408 DVSS.n384 0.00334
R20802 DVSS.n404 DVSS.n384 0.00334
R20803 DVSS.n404 DVSS.n403 0.00334
R20804 DVSS.n403 DVSS.n402 0.00334
R20805 DVSS.n402 DVSS.n390 0.00334
R20806 DVSS.n398 DVSS.n390 0.00334
R20807 DVSS.n398 DVSS.n397 0.00334
R20808 DVSS.n397 DVSS.n199 0.00334
R20809 DVSS.n616 DVSS.n199 0.00334
R20810 DVSS.n616 DVSS.n615 0.00334
R20811 DVSS.n615 DVSS.n614 0.00334
R20812 DVSS.n614 DVSS.n200 0.00334
R20813 DVSS.n609 DVSS.n608 0.00334
R20814 DVSS.n608 DVSS.n607 0.00334
R20815 DVSS.n607 DVSS.n580 0.00334
R20816 DVSS.n603 DVSS.n580 0.00334
R20817 DVSS.n603 DVSS.n602 0.00334
R20818 DVSS.n602 DVSS.n601 0.00334
R20819 DVSS.n601 DVSS.n586 0.00334
R20820 DVSS.n597 DVSS.n586 0.00334
R20821 DVSS.n597 DVSS.n596 0.00334
R20822 DVSS.n596 DVSS.n595 0.00334
R20823 DVSS.n595 DVSS.n166 0.00334
R20824 DVSS.n692 DVSS.n166 0.00334
R20825 DVSS.n693 DVSS.n692 0.00334
R20826 DVSS.n694 DVSS.n693 0.00334
R20827 DVSS.n694 DVSS.n162 0.00334
R20828 DVSS.n700 DVSS.n162 0.00334
R20829 DVSS.n701 DVSS.n700 0.00334
R20830 DVSS.n702 DVSS.n701 0.00334
R20831 DVSS.n702 DVSS.n158 0.00334
R20832 DVSS.n708 DVSS.n158 0.00334
R20833 DVSS.n709 DVSS.n708 0.00334
R20834 DVSS.n711 DVSS.n709 0.00334
R20835 DVSS.n711 DVSS.n710 0.00334
R20836 DVSS.n5664 DVSS.n5663 0.00334
R20837 DVSS.n5663 DVSS.n5662 0.00334
R20838 DVSS.n5662 DVSS.n137 0.00334
R20839 DVSS.n5658 DVSS.n137 0.00334
R20840 DVSS.n5658 DVSS.n5657 0.00334
R20841 DVSS.n5657 DVSS.n5656 0.00334
R20842 DVSS.n5656 DVSS.n143 0.00334
R20843 DVSS.n5652 DVSS.n143 0.00334
R20844 DVSS.n5652 DVSS.n5651 0.00334
R20845 DVSS.n5651 DVSS.n5650 0.00334
R20846 DVSS.n5650 DVSS.n5623 0.00334
R20847 DVSS.n5646 DVSS.n5623 0.00334
R20848 DVSS.n5646 DVSS.n5645 0.00334
R20849 DVSS.n5645 DVSS.n5644 0.00334
R20850 DVSS.n5644 DVSS.n5629 0.00334
R20851 DVSS.n5640 DVSS.n5629 0.00334
R20852 DVSS.n5640 DVSS.n5639 0.00334
R20853 DVSS.n5639 DVSS.n5638 0.00334
R20854 DVSS.n5638 DVSS.n51 0.00334
R20855 DVSS.n5735 DVSS.n51 0.00334
R20856 DVSS.n5736 DVSS.n5735 0.00334
R20857 DVSS.n5737 DVSS.n5736 0.00334
R20858 DVSS.n5737 DVSS.n44 0.00334
R20859 DVSS.n5775 DVSS.n45 0.00334
R20860 DVSS.n5771 DVSS.n45 0.00334
R20861 DVSS.n5771 DVSS.n5770 0.00334
R20862 DVSS.n5770 DVSS.n5769 0.00334
R20863 DVSS.n5769 DVSS.n5746 0.00334
R20864 DVSS.n5765 DVSS.n5746 0.00334
R20865 DVSS.n5765 DVSS.n5764 0.00334
R20866 DVSS.n5764 DVSS.n5763 0.00334
R20867 DVSS.n5763 DVSS.n5752 0.00334
R20868 DVSS.n5759 DVSS.n5752 0.00334
R20869 DVSS.n5759 DVSS.n5758 0.00334
R20870 DVSS.n5816 DVSS.n5815 0.00334
R20871 DVSS.n368 DVSS.n226 0.00334
R20872 DVSS.n467 DVSS.n226 0.00334
R20873 DVSS.n468 DVSS.n467 0.00334
R20874 DVSS.n469 DVSS.n468 0.00334
R20875 DVSS.n469 DVSS.n222 0.00334
R20876 DVSS.n475 DVSS.n222 0.00334
R20877 DVSS.n476 DVSS.n475 0.00334
R20878 DVSS.n477 DVSS.n476 0.00334
R20879 DVSS.n477 DVSS.n218 0.00334
R20880 DVSS.n483 DVSS.n218 0.00334
R20881 DVSS.n484 DVSS.n483 0.00334
R20882 DVSS.n485 DVSS.n484 0.00334
R20883 DVSS.n485 DVSS.n214 0.00334
R20884 DVSS.n491 DVSS.n214 0.00334
R20885 DVSS.n492 DVSS.n491 0.00334
R20886 DVSS.n493 DVSS.n492 0.00334
R20887 DVSS.n493 DVSS.n210 0.00334
R20888 DVSS.n500 DVSS.n210 0.00334
R20889 DVSS.n501 DVSS.n500 0.00334
R20890 DVSS.n503 DVSS.n501 0.00334
R20891 DVSS.n503 DVSS.n502 0.00334
R20892 DVSS.n502 DVSS.n207 0.00334
R20893 DVSS.n510 DVSS.n207 0.00334
R20894 DVSS.n573 DVSS.n572 0.00334
R20895 DVSS.n572 DVSS.n571 0.00334
R20896 DVSS.n571 DVSS.n512 0.00334
R20897 DVSS.n567 DVSS.n512 0.00334
R20898 DVSS.n567 DVSS.n566 0.00334
R20899 DVSS.n566 DVSS.n565 0.00334
R20900 DVSS.n565 DVSS.n517 0.00334
R20901 DVSS.n561 DVSS.n517 0.00334
R20902 DVSS.n561 DVSS.n560 0.00334
R20903 DVSS.n560 DVSS.n559 0.00334
R20904 DVSS.n559 DVSS.n523 0.00334
R20905 DVSS.n555 DVSS.n523 0.00334
R20906 DVSS.n555 DVSS.n554 0.00334
R20907 DVSS.n554 DVSS.n553 0.00334
R20908 DVSS.n553 DVSS.n529 0.00334
R20909 DVSS.n549 DVSS.n529 0.00334
R20910 DVSS.n549 DVSS.n548 0.00334
R20911 DVSS.n548 DVSS.n547 0.00334
R20912 DVSS.n547 DVSS.n535 0.00334
R20913 DVSS.n543 DVSS.n535 0.00334
R20914 DVSS.n543 DVSS.n542 0.00334
R20915 DVSS.n542 DVSS.n152 0.00334
R20916 DVSS.n719 DVSS.n152 0.00334
R20917 DVSS.n722 DVSS.n721 0.00334
R20918 DVSS.n722 DVSS.n148 0.00334
R20919 DVSS.n728 DVSS.n148 0.00334
R20920 DVSS.n729 DVSS.n728 0.00334
R20921 DVSS.n5612 DVSS.n729 0.00334
R20922 DVSS.n5612 DVSS.n5611 0.00334
R20923 DVSS.n5611 DVSS.n5610 0.00334
R20924 DVSS.n5610 DVSS.n730 0.00334
R20925 DVSS.n5606 DVSS.n730 0.00334
R20926 DVSS.n5606 DVSS.n5605 0.00334
R20927 DVSS.n5605 DVSS.n5604 0.00334
R20928 DVSS.n5604 DVSS.n735 0.00334
R20929 DVSS.n5600 DVSS.n735 0.00334
R20930 DVSS.n5600 DVSS.n5599 0.00334
R20931 DVSS.n5599 DVSS.n5598 0.00334
R20932 DVSS.n5598 DVSS.n741 0.00334
R20933 DVSS.n5594 DVSS.n741 0.00334
R20934 DVSS.n5594 DVSS.n5593 0.00334
R20935 DVSS.n5593 DVSS.n5592 0.00334
R20936 DVSS.n5592 DVSS.n747 0.00334
R20937 DVSS.n5588 DVSS.n747 0.00334
R20938 DVSS.n5588 DVSS.n5587 0.00334
R20939 DVSS.n5587 DVSS.n5586 0.00334
R20940 DVSS.n5582 DVSS.n5581 0.00334
R20941 DVSS.n5581 DVSS.n5580 0.00334
R20942 DVSS.n5580 DVSS.n808 0.00334
R20943 DVSS.n5576 DVSS.n808 0.00334
R20944 DVSS.n5576 DVSS.n5575 0.00334
R20945 DVSS.n5575 DVSS.n5574 0.00334
R20946 DVSS.n5574 DVSS.n814 0.00334
R20947 DVSS.n5570 DVSS.n814 0.00334
R20948 DVSS.n5570 DVSS.n5569 0.00334
R20949 DVSS.n5569 DVSS.n5568 0.00334
R20950 DVSS.n5568 DVSS.n820 0.00334
R20951 DVSS.n5564 DVSS.n5563 0.00334
R20952 DVSS.n4192 DVSS.n1364 0.00334
R20953 DVSS.n4198 DVSS.n1364 0.00334
R20954 DVSS.n4199 DVSS.n4198 0.00334
R20955 DVSS.n4200 DVSS.n4199 0.00334
R20956 DVSS.n4200 DVSS.n1360 0.00334
R20957 DVSS.n4207 DVSS.n1360 0.00334
R20958 DVSS.n4208 DVSS.n4207 0.00334
R20959 DVSS.n4209 DVSS.n4208 0.00334
R20960 DVSS.n4209 DVSS.n1356 0.00334
R20961 DVSS.n4216 DVSS.n1356 0.00334
R20962 DVSS.n4217 DVSS.n4216 0.00334
R20963 DVSS.n4218 DVSS.n4217 0.00334
R20964 DVSS.n4218 DVSS.n1352 0.00334
R20965 DVSS.n4224 DVSS.n1352 0.00334
R20966 DVSS.n4225 DVSS.n4224 0.00334
R20967 DVSS.n4226 DVSS.n4225 0.00334
R20968 DVSS.n4226 DVSS.n1348 0.00334
R20969 DVSS.n4232 DVSS.n1348 0.00334
R20970 DVSS.n4233 DVSS.n4232 0.00334
R20971 DVSS.n4234 DVSS.n4233 0.00334
R20972 DVSS.n4234 DVSS.n1344 0.00334
R20973 DVSS.n4241 DVSS.n1344 0.00334
R20974 DVSS.n4242 DVSS.n4241 0.00334
R20975 DVSS.n4243 DVSS.n4242 0.00334
R20976 DVSS.n4243 DVSS.n1340 0.00334
R20977 DVSS.n4249 DVSS.n1340 0.00334
R20978 DVSS.n4250 DVSS.n4249 0.00334
R20979 DVSS.n4251 DVSS.n4250 0.00334
R20980 DVSS.n4251 DVSS.n1336 0.00334
R20981 DVSS.n4257 DVSS.n1336 0.00334
R20982 DVSS.n4258 DVSS.n4257 0.00334
R20983 DVSS.n4259 DVSS.n4258 0.00334
R20984 DVSS.n4259 DVSS.n1332 0.00334
R20985 DVSS.n4265 DVSS.n1332 0.00334
R20986 DVSS.n4266 DVSS.n4265 0.00334
R20987 DVSS.n4267 DVSS.n4266 0.00334
R20988 DVSS.n4267 DVSS.n1328 0.00334
R20989 DVSS.n4273 DVSS.n1328 0.00334
R20990 DVSS.n4274 DVSS.n4273 0.00334
R20991 DVSS.n4275 DVSS.n4274 0.00334
R20992 DVSS.n4275 DVSS.n1324 0.00334
R20993 DVSS.n4281 DVSS.n1324 0.00334
R20994 DVSS.n4282 DVSS.n4281 0.00334
R20995 DVSS.n4283 DVSS.n4282 0.00334
R20996 DVSS.n4283 DVSS.n1320 0.00334
R20997 DVSS.n4289 DVSS.n1320 0.00334
R20998 DVSS.n4290 DVSS.n4289 0.00334
R20999 DVSS.n4291 DVSS.n4290 0.00334
R21000 DVSS.n4292 DVSS.n4291 0.00334
R21001 DVSS.n4293 DVSS.n4292 0.00334
R21002 DVSS.n4296 DVSS.n4293 0.00334
R21003 DVSS.n4297 DVSS.n4296 0.00334
R21004 DVSS.n4298 DVSS.n4297 0.00334
R21005 DVSS.n4299 DVSS.n4298 0.00334
R21006 DVSS.n4302 DVSS.n4299 0.00334
R21007 DVSS.n4303 DVSS.n4302 0.00334
R21008 DVSS.n4304 DVSS.n4303 0.00334
R21009 DVSS.n4305 DVSS.n4304 0.00334
R21010 DVSS.n4308 DVSS.n4305 0.00334
R21011 DVSS.n4309 DVSS.n4308 0.00334
R21012 DVSS.n4310 DVSS.n4309 0.00334
R21013 DVSS.n4313 DVSS.n4310 0.00334
R21014 DVSS.n4314 DVSS.n4313 0.00334
R21015 DVSS.n4315 DVSS.n4314 0.00334
R21016 DVSS.n4316 DVSS.n4315 0.00334
R21017 DVSS.n4319 DVSS.n4316 0.00334
R21018 DVSS.n4320 DVSS.n4319 0.00334
R21019 DVSS.n4321 DVSS.n4320 0.00334
R21020 DVSS.n4322 DVSS.n4321 0.00334
R21021 DVSS.n4325 DVSS.n4322 0.00334
R21022 DVSS.n4326 DVSS.n4325 0.00334
R21023 DVSS.n4327 DVSS.n4326 0.00334
R21024 DVSS.n4328 DVSS.n4327 0.00334
R21025 DVSS.n4331 DVSS.n4328 0.00334
R21026 DVSS.n4332 DVSS.n4331 0.00334
R21027 DVSS.n4333 DVSS.n4332 0.00334
R21028 DVSS.n4334 DVSS.n1176 0.00334
R21029 DVSS.n4712 DVSS.n1252 0.00332857
R21030 DVSS.n4714 DVSS.n4713 0.00332857
R21031 DVSS.n4723 DVSS.n1249 0.00332857
R21032 DVSS.n4722 DVSS.n1243 0.00332857
R21033 DVSS.n4731 DVSS.n4730 0.00332857
R21034 DVSS.n1244 DVSS.n1239 0.00332857
R21035 DVSS.n4737 DVSS.n4736 0.00332857
R21036 DVSS.n4979 DVSS.n1154 0.00332857
R21037 DVSS.n362 DVSS.n361 0.00332
R21038 DVSS.n363 DVSS.n243 0.00332
R21039 DVSS.n366 DVSS.n364 0.00332
R21040 DVSS.n367 DVSS.n250 0.00332
R21041 DVSS.n253 DVSS.n245 0.00332
R21042 DVSS.n360 DVSS.n254 0.00332
R21043 DVSS.n1211 DVSS.n1187 0.00330488
R21044 DVSS.n1196 DVSS.n1182 0.00330488
R21045 DVSS.n687 DVSS.n170 0.00329
R21046 DVSS.n689 DVSS.n168 0.00329
R21047 DVSS.n526 DVSS.n169 0.00329
R21048 DVSS.n5564 DVSS 0.00326
R21049 DVSS DVSS.n4334 0.00326
R21050 DVSS.n4183 DVSS.n4182 0.0032
R21051 DVSS.n3905 DVSS.n1573 0.0032
R21052 DVSS.n5731 DVSS.n55 0.00319327
R21053 DVSS.n1859 DVSS.n1427 0.00319022
R21054 DVSS.n3989 DVSS.n1434 0.00319022
R21055 VSS DVSS.n1503 0.00314706
R21056 DVSS.n3946 VSS 0.00314706
R21057 DVSS.n463 DVSS.n229 0.00314706
R21058 DVSS.n3886 DVSS.n3885 0.00313571
R21059 DVSS.n1609 DVSS.n1605 0.00313571
R21060 DVSS.n311 DVSS.n258 0.00311
R21061 DVSS.n373 DVSS.n244 0.00311
R21062 DVSS.n465 DVSS.n464 0.00311
R21063 DVSS.n4938 DVSS.n4937 0.00309529
R21064 DVSS.n1624 DVSS.n1620 0.00307143
R21065 DVSS.n3841 DVSS.n1625 0.00307143
R21066 DVSS.n3840 DVSS.n3828 0.00307143
R21067 DVSS.n5361 DVSS.n951 0.00300714
R21068 DVSS.n4854 DVSS.n1177 0.00300714
R21069 DVSS.n3894 DVSS.n1590 0.00300714
R21070 DVSS.n3061 DVSS.n3060 0.003
R21071 DVSS.n3095 DVSS.n3094 0.003
R21072 DVSS.n2681 DVSS.n2664 0.003
R21073 DVSS.n3272 DVSS.n3271 0.003
R21074 DVSS.n1827 DVSS.n1819 0.00297706
R21075 DVSS.n2803 DVSS.n2790 0.00296479
R21076 DVSS.n2812 DVSS.n2811 0.00296479
R21077 DVSS.n2792 DVSS.n2786 0.00296479
R21078 DVSS.n2821 DVSS.n2781 0.00296479
R21079 DVSS.n2837 DVSS.n2836 0.00296479
R21080 DVSS.n2845 DVSS.n2776 0.00296479
R21081 DVSS.n2844 DVSS.n2770 0.00296479
R21082 DVSS.n2856 DVSS.n2855 0.00296479
R21083 DVSS.n2772 DVSS.n2766 0.00296479
R21084 DVSS.n2865 DVSS.n2761 0.00296479
R21085 DVSS.n2886 DVSS.n2885 0.00296479
R21086 DVSS.n2894 DVSS.n2756 0.00296479
R21087 DVSS.n2893 DVSS.n2750 0.00296479
R21088 DVSS.n2909 DVSS.n2908 0.00296479
R21089 DVSS.n2905 DVSS.n2752 0.00296479
R21090 DVSS.n2904 DVSS.n2744 0.00296479
R21091 DVSS.n2920 DVSS.n2739 0.00296479
R21092 DVSS.n2948 DVSS.n2947 0.00296479
R21093 DVSS.n2957 DVSS.n2734 0.00296479
R21094 DVSS.n2956 DVSS.n2727 0.00296479
R21095 DVSS.n2964 DVSS.n2963 0.00296479
R21096 DVSS.n2730 DVSS.n2729 0.00296479
R21097 DVSS.n2976 DVSS.n2721 0.00296479
R21098 DVSS.n2975 DVSS.n2715 0.00296479
R21099 DVSS.n2987 DVSS.n2986 0.00296479
R21100 DVSS.n2717 DVSS.n2711 0.00296479
R21101 DVSS.n2995 DVSS.n2706 0.00296479
R21102 DVSS.n3011 DVSS.n3010 0.00296479
R21103 DVSS.n3022 DVSS.n2701 0.00296479
R21104 DVSS.n3021 DVSS.n2694 0.00296479
R21105 DVSS.n3034 DVSS.n3033 0.00296479
R21106 DVSS.n2697 DVSS.n2690 0.00296479
R21107 DVSS.n3041 DVSS.n2685 0.00296479
R21108 DVSS.n3052 DVSS.n3051 0.00296479
R21109 DVSS.n3063 DVSS.n2680 0.00296479
R21110 DVSS.n3062 DVSS.n2666 0.00296479
R21111 DVSS.n3550 DVSS.n2667 0.00296479
R21112 DVSS.n3254 DVSS.n2673 0.00296479
R21113 DVSS.n3543 DVSS.n3542 0.00296479
R21114 DVSS.n3539 DVSS.n2675 0.00296479
R21115 DVSS.n3538 DVSS.n3073 0.00296479
R21116 DVSS.n3265 DVSS.n3080 0.00296479
R21117 DVSS.n3530 DVSS.n3529 0.00296479
R21118 DVSS.n3526 DVSS.n3082 0.00296479
R21119 DVSS.n3525 DVSS.n3090 0.00296479
R21120 DVSS.n3277 DVSS.n3100 0.00296479
R21121 DVSS.n3518 DVSS.n3517 0.00296479
R21122 DVSS.n3514 DVSS.n3102 0.00296479
R21123 DVSS.n3513 DVSS.n3110 0.00296479
R21124 DVSS.n3288 DVSS.n3117 0.00296479
R21125 DVSS.n3505 DVSS.n3504 0.00296479
R21126 DVSS.n3501 DVSS.n3119 0.00296479
R21127 DVSS.n3500 DVSS.n3127 0.00296479
R21128 DVSS.n3301 DVSS.n3136 0.00296479
R21129 DVSS.n3493 DVSS.n3492 0.00296479
R21130 DVSS.n3489 DVSS.n3138 0.00296479
R21131 DVSS.n3488 DVSS.n3146 0.00296479
R21132 DVSS.n3313 DVSS.n3154 0.00296479
R21133 DVSS.n3479 DVSS.n3478 0.00296479
R21134 DVSS.n3475 DVSS.n3156 0.00296479
R21135 DVSS.n3474 DVSS.n3164 0.00296479
R21136 DVSS.n3324 DVSS.n3171 0.00296479
R21137 DVSS.n3467 DVSS.n3466 0.00296479
R21138 DVSS.n3463 DVSS.n3173 0.00296479
R21139 DVSS.n3462 DVSS.n3181 0.00296479
R21140 DVSS.n3337 DVSS.n3191 0.00296479
R21141 DVSS.n3455 DVSS.n3454 0.00296479
R21142 DVSS.n3451 DVSS.n3193 0.00296479
R21143 DVSS.n3450 DVSS.n3201 0.00296479
R21144 DVSS.n3349 DVSS.n3209 0.00296479
R21145 DVSS.n3443 DVSS.n3442 0.00296479
R21146 DVSS.n3439 DVSS.n3211 0.00296479
R21147 DVSS.n3438 DVSS.n3219 0.00296479
R21148 DVSS.n3361 DVSS.n3226 0.00296479
R21149 DVSS.n3430 DVSS.n3429 0.00296479
R21150 DVSS.n3426 DVSS.n3228 0.00296479
R21151 DVSS.n3425 DVSS.n3236 0.00296479
R21152 DVSS.n3373 DVSS.n3243 0.00296479
R21153 DVSS.n3418 DVSS.n3417 0.00296479
R21154 DVSS.n426 DVSS.n242 0.00294344
R21155 DVSS DVSS.n2889 0.00293842
R21156 DVSS.n2882 DVSS 0.00293842
R21157 DVSS.n2108 DVSS.n2107 0.00293243
R21158 DVSS.n106 DVSS.n105 0.0029
R21159 DVSS.n5740 DVSS.n48 0.0029
R21160 DVSS.n805 DVSS.n804 0.0029
R21161 DVSS.n4484 DVSS 0.00286842
R21162 DVSS.n4442 DVSS 0.00286842
R21163 DVSS.n1308 DVSS 0.00286842
R21164 DVSS.n1450 VSS 0.00286842
R21165 DVSS DVSS.n1172 0.00286842
R21166 DVSS.n5778 DVSS.n5777 0.00286
R21167 DVSS.n5776 DVSS.n5775 0.00286
R21168 DVSS.n5582 DVSS.n43 0.00286
R21169 DVSS DVSS.n28 0.00282
R21170 DVSS DVSS.n4333 0.00278
R21171 DVSS.n3058 DVSS.n2670 0.00271675
R21172 DVSS.n3554 DVSS.n3553 0.00271675
R21173 DVSS.n5671 DVSS.n5670 0.0027
R21174 DVSS.n5664 DVSS.n129 0.0027
R21175 DVSS.n721 DVSS.n720 0.0027
R21176 DVSS.n4368 DVSS.n4307 0.00269
R21177 DVSS.n4621 DVSS.n4620 0.00262143
R21178 DVSS.n4617 DVSS.n4614 0.00262143
R21179 DVSS.n4616 DVSS.n1269 0.00262143
R21180 DVSS.n4684 DVSS.n4683 0.00262143
R21181 DVSS.n4691 DVSS.n1264 0.00262143
R21182 DVSS.n4690 DVSS.n1265 0.00262143
R21183 DVSS.n4696 DVSS.n1260 0.00262143
R21184 DVSS.n4875 DVSS.n4808 0.00262143
R21185 DVSS.n4831 DVSS.n4830 0.00262143
R21186 DVSS.n4872 DVSS.n4871 0.00262143
R21187 DVSS.n1204 DVSS.n1189 0.00257317
R21188 DVSS.n1203 DVSS.n1184 0.00257317
R21189 DVSS.n4190 DVSS.n1366 0.00257
R21190 DVSS.n4365 DVSS.n4307 0.00257
R21191 DVSS.n1942 DVSS.n1934 0.00256422
R21192 DVSS.n1778 DVSS.n1777 0.00256422
R21193 DVSS.n4652 DVSS.n4582 0.00255714
R21194 DVSS.n4649 DVSS.n4648 0.00255714
R21195 DVSS.n4591 DVSS.n4585 0.00255714
R21196 DVSS.n4642 DVSS.n4592 0.00255714
R21197 DVSS.n4641 DVSS.n4593 0.00255714
R21198 DVSS.n4603 DVSS.n4602 0.00255714
R21199 DVSS.n4636 DVSS.n4635 0.00255714
R21200 DVSS.n634 DVSS.n633 0.00254
R21201 DVSS.n609 DVSS.n186 0.00254
R21202 DVSS.n573 DVSS.n511 0.00254
R21203 DVSS.n765 DVSS.n55 0.00251995
R21204 DVSS.n3549 DVSS.n2668 0.0025
R21205 DVSS.n3531 DVSS.n3079 0.0025
R21206 DVSS.n3552 DVSS.n3551 0.0025
R21207 DVSS.n3270 DVSS.n3081 0.0025
R21208 DVSS.n2170 DVSS.n1797 0.00249286
R21209 DVSS.n2145 DVSS.n1799 0.00249286
R21210 DVSS DVSS.n3398 0.00247183
R21211 DVSS.n1877 DVSS.n1873 0.00242857
R21212 DVSS.n1874 DVSS.n1789 0.00242857
R21213 DVSS.n359 DVSS.n247 0.00238
R21214 DVSS.n371 DVSS.n370 0.00238
R21215 DVSS.n369 DVSS.n368 0.00238
R21216 DVSS.n3803 DVSS.n3802 0.00236429
R21217 DVSS.n105 DVSS.n103 0.00236
R21218 DVSS.n50 DVSS.n48 0.00236
R21219 DVSS.n804 DVSS.n753 0.00236
R21220 DVSS.n427 DVSS.n426 0.00233258
R21221 DVSS.n5551 DVSS 0.0023
R21222 DVSS DVSS.n4857 0.0023
R21223 DVSS.n4856 DVSS 0.0023
R21224 DVSS.n2632 VSS 0.0023
R21225 DVSS.n3727 DVSS 0.0023
R21226 DVSS.n2022 DVSS 0.0023
R21227 DVSS.n4036 DVSS 0.0023
R21228 VSS DVSS.n2283 0.0023
R21229 DVSS.n2279 VSS 0.0023
R21230 VSS DVSS.n2269 0.0023
R21231 DVSS.n3093 DVSS.n3078 0.0022734
R21232 DVSS.n3133 DVSS.n3132 0.0022734
R21233 DVSS.n3298 DVSS.n3297 0.0022734
R21234 DVSS.n2390 DVSS.n2275 0.00223571
R21235 DVSS.n2392 DVSS.n2278 0.00223571
R21236 DVSS.n2419 DVSS.n2279 0.00223571
R21237 DVSS.n2646 DVSS.n2421 0.00223571
R21238 DVSS.n2643 DVSS.n2636 0.00223571
R21239 DVSS.n2648 DVSS.n2269 0.00223571
R21240 DVSS.n312 DVSS.n311 0.00215
R21241 DVSS.n374 DVSS.n373 0.00215
R21242 DVSS.n464 DVSS.n224 0.00215
R21243 DVSS.n3020 DVSS.n3019 0.002
R21244 DVSS.n3508 DVSS.n3113 0.002
R21245 DVSS.n3004 DVSS.n2702 0.002
R21246 DVSS.n3290 DVSS.n3289 0.002
R21247 DVSS.n3677 DVSS.n3676 0.00197857
R21248 DVSS.n687 DVSS.n686 0.00197
R21249 DVSS.n690 DVSS.n689 0.00197
R21250 DVSS.n527 DVSS.n169 0.00197
R21251 DVSS.n5758 DVSS 0.00196
R21252 DVSS.n5553 DVSS 0.00191429
R21253 DVSS.n5816 DVSS 0.00188
R21254 DVSS.n3878 DVSS.n3877 0.00185
R21255 DVSS.n3866 DVSS.n1610 0.00185
R21256 DVSS.n1212 DVSS.n1188 0.00184146
R21257 DVSS.n1195 DVSS.n1185 0.00184146
R21258 DVSS.n3396 DVSS 0.00181455
R21259 DVSS.n5756 DVSS 0.00173
R21260 DVSS DVSS.n0 0.00173
R21261 DVSS.n2395 VSS 0.0017
R21262 DVSS.n630 DVSS.n184 0.0017
R21263 DVSS.n577 DVSS.n202 0.0017
R21264 DVSS.n576 DVSS.n204 0.0017
R21265 DVSS.n509 DVSS.n203 0.0017
R21266 DVSS.n612 DVSS.n611 0.0017
R21267 DVSS.n631 DVSS.n185 0.0017
R21268 DVSS.n5717 DVSS.n5716 0.00167
R21269 DVSS.n5732 DVSS.n54 0.00167
R21270 DVSS.n801 DVSS.n751 0.00167
R21271 DVSS.n4852 DVSS.n1178 0.00165714
R21272 DVSS.n4848 DVSS.n1180 0.00165714
R21273 DVSS.n2116 DVSS.n1810 0.00165714
R21274 DVSS.n2088 DVSS.n1809 0.00165714
R21275 DVSS.n5059 DVSS.n1110 0.00165714
R21276 DVSS.n5058 DVSS.n1111 0.00165714
R21277 DVSS.n5055 DVSS.n5054 0.00165714
R21278 DVSS.n1117 DVSS.n1113 0.00165714
R21279 DVSS.n5048 DVSS.n1118 0.00165714
R21280 DVSS.n5047 DVSS.n1119 0.00165714
R21281 DVSS.n5044 DVSS.n5043 0.00165714
R21282 DVSS.n1125 DVSS.n1121 0.00165714
R21283 DVSS.n4753 DVSS.n1230 0.00159286
R21284 DVSS.n4752 DVSS.n1231 0.00159286
R21285 DVSS.n4759 DVSS.n1228 0.00159286
R21286 DVSS.n4761 DVSS.n4760 0.00159286
R21287 DVSS.n4917 DVSS.n1222 0.00159286
R21288 DVSS.n4916 DVSS.n1223 0.00159286
R21289 DVSS.n4770 DVSS.n4767 0.00159286
R21290 DVSS.n1378 DVSS.n1373 0.00159286
R21291 DVSS.n4171 DVSS.n4170 0.00159286
R21292 DVSS.n4168 DVSS.n1384 0.00159286
R21293 DVSS.n3804 DVSS.n1647 0.00159286
R21294 DVSS.n1866 DVSS.n1383 0.00157001
R21295 DVSS.n1822 DVSS.n1740 0.00152857
R21296 DVSS.n2212 DVSS.n1744 0.00152857
R21297 DVSS.n2970 DVSS.n2723 0.0015
R21298 DVSS.n3487 DVSS.n3486 0.0015
R21299 DVSS.n2934 DVSS.n2926 0.0015
R21300 DVSS.n3248 DVSS.n3145 0.0015
R21301 DVSS.n4238 DVSS.n4237 0.00146
R21302 DVSS.n155 DVSS.n132 0.00146
R21303 DVSS.n715 DVSS.n714 0.00146
R21304 DVSS.n717 DVSS.n716 0.00146
R21305 DVSS.n718 DVSS.n133 0.00146
R21306 DVSS.n5666 DVSS.n134 0.00146
R21307 DVSS.n5668 DVSS.n5667 0.00146
R21308 DVSS.n3534 DVSS.n3533 0.0013867
R21309 DVSS.n3268 DVSS.n3253 0.0013867
R21310 DVSS DVSS.n4342 0.00134
R21311 DVSS.n4341 DVSS 0.00134
R21312 DVSS.n823 DVSS 0.00134
R21313 DVSS DVSS.n5566 0.00134
R21314 DVSS.n4095 DVSS.n1431 0.00133571
R21315 DVSS.n4004 DVSS.n1436 0.00133571
R21316 DVSS.n4093 DVSS.n4092 0.00133571
R21317 DVSS.n1619 DVSS.n1615 0.00133571
R21318 DVSS.n4412 DVSS.n4411 0.00131
R21319 DVSS.n4341 DVSS.n4340 0.00131
R21320 DVSS.n5676 DVSS.n123 0.00131
R21321 DVSS.n5617 DVSS.n141 0.00131
R21322 DVSS.n5615 DVSS.n144 0.00131
R21323 DVSS.n633 DVSS.n632 0.0013
R21324 DVSS.n200 DVSS.n186 0.0013
R21325 DVSS.n511 DVSS.n510 0.0013
R21326 DVSS.n106 DVSS.n40 0.00122
R21327 DVSS.n5741 DVSS.n5740 0.00122
R21328 DVSS.n805 DVSS.n47 0.00122
R21329 DVSS.n5585 DVSS.n5584 0.00122
R21330 DVSS.n5739 DVSS.n46 0.00122
R21331 DVSS.n107 DVSS.n41 0.00122
R21332 DVSS.n4934 DVSS 0.00120714
R21333 DVSS.n1675 DVSS.n1674 0.00120714
R21334 DVSS.n3778 DVSS.n1682 0.00120714
R21335 DVSS.n5076 DVSS.n1100 0.00120714
R21336 DVSS.n5075 DVSS.n5074 0.00120714
R21337 DVSS.n4204 DVSS.n4203 0.00119
R21338 DVSS.n4213 DVSS.n1354 0.00119
R21339 DVSS.n5670 DVSS.n5669 0.00114
R21340 DVSS.n710 DVSS.n129 0.00114
R21341 DVSS.n720 DVSS.n719 0.00114
R21342 DVSS.n4423 DVSS.n4422 0.00107
R21343 DVSS.n4941 DVSS.n4940 0.00107
R21344 DVSS.n4335 DVSS 0.00106
R21345 DVSS.n6 DVSS.n5 0.00104
R21346 DVSS.n5813 DVSS.n5812 0.00104
R21347 DVSS.n829 DVSS.n828 0.00104
R21348 DVSS.n5561 DVSS.n5560 0.00104
R21349 DVSS.n5801 DVSS 0.00102
R21350 DVSS.n622 DVSS.n621 0.00101
R21351 DVSS.n619 DVSS.n195 0.00101
R21352 DVSS.n497 DVSS.n194 0.00101
R21353 DVSS.n2814 DVSS.n2813 0.001
R21354 DVSS.n2915 DVSS.n2745 0.001
R21355 DVSS.n3186 DVSS.n3185 0.001
R21356 DVSS.n3242 DVSS.n3239 0.001
R21357 DVSS.n2799 DVSS.n2791 0.001
R21358 DVSS.n2873 DVSS.n2743 0.001
R21359 DVSS.n3332 DVSS.n3246 0.001
R21360 DVSS.n3374 DVSS.n3372 0.001
R21361 DVSS.n5777 DVSS.n42 0.00098
R21362 DVSS.n5776 DVSS.n44 0.00098
R21363 DVSS.n5586 DVSS.n43 0.00098
R21364 DVSS.n1595 DVSS.n1594 0.00095
R21365 DVSS.n3250 DVSS.n3098 0.00094335
R21366 DVSS.n3281 DVSS.n3251 0.00094335
R21367 DVSS.n257 DVSS.n252 0.00092
R21368 DVSS.n425 DVSS.n424 0.00092
R21369 DVSS.n365 DVSS.n228 0.00092
R21370 DVSS.n5553 DVSS.n5552 0.000885714
R21371 DVSS.n1850 DVSS.n1386 0.000856671
R21372 DVSS.n1841 DVSS.n1380 0.000856671
R21373 DVSS DVSS.n2794 0.000721675
R21374 DVSS.n2801 DVSS 0.000721675
R21375 DVSS DVSS.n3396 0.000687793
R21376 DVSS.n5803 DVSS 0.00068
R21377 DVSS.n5802 DVSS 0.00068
R21378 DVSS.n5550 DVSS 0.000671429
R21379 DVSS DVSS.n4845 0.000671429
R21380 DVSS.n2633 VSS 0.000671429
R21381 DVSS DVSS.n3726 0.000671429
R21382 DVSS.n2021 DVSS 0.000671429
R21383 DVSS DVSS.n4035 0.000671429
R21384 VSS DVSS.n2395 0.000671429
R21385 DVSS.n1823 DVSS.n1822 0.000628571
R21386 DVSS.n2212 DVSS.n2211 0.000628571
R21387 DVSS.n1892 DVSS.n1745 0.000628571
R21388 DVSS.n1899 DVSS.n1893 0.000628571
R21389 DVSS.n1898 DVSS.n1891 0.000628571
R21390 DVSS.n1901 DVSS.n1888 0.000628571
R21391 DVSS.n1902 DVSS.n1759 0.000628571
R21392 DVSS.n1884 DVSS.n1761 0.000628571
R21393 DVSS.n1908 DVSS.n1758 0.000628571
R21394 DVSS.n2197 DVSS.n1762 0.000628571
R21395 DVSS.n2195 DVSS.n1763 0.000628571
R21396 DVSS.n1770 DVSS.n1769 0.000628571
R21397 DVSS.n2189 DVSS.n2188 0.000628571
R21398 DVSS.n1870 DVSS.n1771 0.000628571
R21399 DVSS.n1873 DVSS.n1787 0.000628571
R21400 DVSS.n2179 DVSS.n1789 0.000628571
R21401 DVSS.n2171 DVSS.n2170 0.000628571
R21402 DVSS.n1799 DVSS.n1798 0.000628571
R21403 DVSS.n2144 DVSS.n1926 0.000628571
R21404 DVSS.n1931 DVSS.n1930 0.000628571
R21405 DVSS.n2138 DVSS.n2137 0.000628571
R21406 DVSS.n1962 DVSS.n1932 0.000628571
R21407 DVSS.n1981 DVSS.n1963 0.000628571
R21408 DVSS.n1966 DVSS.n1960 0.000628571
R21409 DVSS.n1973 DVSS.n1961 0.000628571
R21410 DVSS.n1983 DVSS.n1958 0.000628571
R21411 DVSS.n1985 DVSS.n1984 0.000628571
R21412 DVSS.n2124 DVSS.n1952 0.000628571
R21413 DVSS.n2123 DVSS.n1953 0.000628571
R21414 DVSS.n2085 DVSS.n2084 0.000628571
R21415 DVSS.n2117 DVSS.n2116 0.000628571
R21416 DVSS.n2088 DVSS.n2087 0.000628571
R21417 DVSS DVSS.n820 0.00058
R21418 DVSS.n4335 DVSS 0.00058
R21419 DVSS.n3411 DVSS.n1706 0.000570422
R21420 DVSS.n5357 DVSS.n957 0.000566519
R21421 DVSS.n3744 DVSS.n3654 0.000564286
R21422 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t7 40.5676
R21423 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t12 40.5676
R21424 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t2 37.5434
R21425 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t9 37.5434
R21426 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t10 25.3941
R21427 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t5 25.3941
R21428 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t6 24.8726
R21429 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t11 24.8726
R21430 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t4 22.3127
R21431 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t1 21.9898
R21432 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t8 20.6262
R21433 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t3 20.1126
R21434 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n4 8.44221
R21435 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n1 6.88071
R21436 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n0 6.22439
R21437 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n5 4.40816
R21438 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n3 4.09994
R21439 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n2 4.03661
R21440 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t0 2.75597
R21441 DVDD.n1327 DVDD.n1326 13303.9
R21442 DVDD.n1377 DVDD.n1327 13198.6
R21443 DVDD.n1378 DVDD.n1326 10692.2
R21444 DVDD.n1378 DVDD.n1377 10540.9
R21445 DVDD.t61 DVDD.n3446 926.309
R21446 DVDD.n4237 DVDD.t184 902.129
R21447 DVDD.n4237 DVDD.t183 902.129
R21448 DVDD.t57 DVDD.t47 746.523
R21449 DVDD.t18 DVDD.t204 596.601
R21450 DVDD.n1884 DVDD.t185 502.392
R21451 DVDD.n4201 DVDD.t186 502.392
R21452 DVDD.t10 DVDD.t3 482.226
R21453 DVDD.t26 DVDD.t61 425.889
R21454 DVDD.n3448 DVDD.n2685 359.661
R21455 DVDD.t23 DVDD.t191 357.033
R21456 DVDD.t141 DVDD.n2523 353.346
R21457 DVDD.t8 DVDD.t53 349.305
R21458 DVDD.t51 DVDD.n2595 309.892
R21459 DVDD.t204 DVDD.t141 299.846
R21460 DVDD.t2 DVDD.t17 299.846
R21461 DVDD.n2597 DVDD.n2519 261.661
R21462 DVDD.n2290 DVDD.t168 237.623
R21463 DVDD.t77 DVDD.n2260 237.623
R21464 DVDD.n2365 DVDD.t129 237.623
R21465 DVDD.t133 DVDD.n2335 237.623
R21466 DVDD.t49 DVDD.n2288 234.93
R21467 DVDD.n2288 DVDD.t193 234.93
R21468 DVDD.t113 DVDD.n2363 234.93
R21469 DVDD.n2363 DVDD.t67 234.93
R21470 DVDD.t4 DVDD.n3694 210.464
R21471 DVDD.t187 DVDD.n1961 208.482
R21472 DVDD.n1934 DVDD.t139 208.482
R21473 DVDD.t117 DVDD.n1934 208.482
R21474 DVDD.t158 DVDD.n3695 208.102
R21475 DVDD.n1961 DVDD.t148 203.769
R21476 DVDD.t168 DVDD.t146 188.564
R21477 DVDD.t55 DVDD.t49 188.564
R21478 DVDD.t62 DVDD.t193 188.564
R21479 DVDD.t59 DVDD.t77 188.564
R21480 DVDD.t129 DVDD.t172 188.564
R21481 DVDD.t111 DVDD.t113 188.564
R21482 DVDD.t162 DVDD.t67 188.564
R21483 DVDD.t166 DVDD.t133 188.564
R21484 DVDD.t17 DVDD.t18 188.564
R21485 DVDD.t3 DVDD.t2 188.564
R21486 DVDD.t191 DVDD.t12 188.564
R21487 DVDD.t12 DVDD.t8 188.564
R21488 DVDD.t53 DVDD.t57 188.564
R21489 DVDD.t47 DVDD.t51 188.564
R21490 DVDD.n2596 DVDD.t10 145.286
R21491 DVDD.t15 DVDD.t4 143.698
R21492 DVDD.t160 DVDD.t158 143.698
R21493 DVDD.t0 DVDD.t93 139.505
R21494 DVDD.t150 DVDD.t31 139.505
R21495 DVDD.t39 DVDD.t156 139.505
R21496 DVDD.t75 DVDD.t19 139.505
R21497 DVDD.t20 DVDD.t76 139.505
R21498 DVDD.t154 DVDD.t135 139.505
R21499 DVDD.t152 DVDD.t69 139.505
R21500 DVDD.t25 DVDD.t198 139.505
R21501 DVDD.n2595 DVDD.n2594 122.816
R21502 DVDD.n1885 DVDD.t96 121.04
R21503 DVDD.n4202 DVDD.t115 121.04
R21504 DVDD.n4238 DVDD.t29 120.725
R21505 DVDD.n4238 DVDD.t37 120.725
R21506 DVDD.t43 DVDD.n4237 120.725
R21507 DVDD.n4237 DVDD.t202 120.725
R21508 DVDD.t123 DVDD.n4236 120.725
R21509 DVDD.n4236 DVDD.t170 120.725
R21510 DVDD.n1372 DVDD.n1328 114.094
R21511 DVDD.n1376 DVDD.n1328 113.204
R21512 DVDD.t148 DVDD.n1960 108.52
R21513 DVDD.t139 DVDD.n1933 103.829
R21514 DVDD.n1935 DVDD.t117 103.829
R21515 DVDD.n1963 DVDD.t187 103.829
R21516 DVDD.n2575 DVDD.n2569 96.2887
R21517 DVDD.n5487 DVDD.n260 96.0189
R21518 DVDD.n5661 DVDD.n5502 95.6467
R21519 DVDD.n2594 DVDD.n2524 95.5887
R21520 DVDD.n2590 DVDD.n2524 95.5887
R21521 DVDD.n2590 DVDD.n2589 95.5887
R21522 DVDD.n2589 DVDD.n2584 95.5887
R21523 DVDD.n2584 DVDD.n2583 95.5887
R21524 DVDD.n2583 DVDD.n2547 95.5887
R21525 DVDD.n2579 DVDD.n2547 95.5887
R21526 DVDD.n2579 DVDD.n2578 95.5887
R21527 DVDD.n2578 DVDD.n2577 95.5887
R21528 DVDD.n2577 DVDD.n2576 95.5887
R21529 DVDD.n2576 DVDD.n2575 95.5887
R21530 DVDD.n2289 DVDD.t55 95.0546
R21531 DVDD.n2261 DVDD.t62 95.0546
R21532 DVDD.n2364 DVDD.t111 95.0546
R21533 DVDD.n2336 DVDD.t162 95.0546
R21534 DVDD.t146 DVDD.n2289 93.509
R21535 DVDD.n2261 DVDD.t59 93.509
R21536 DVDD.t172 DVDD.n2364 93.509
R21537 DVDD.n2336 DVDD.t166 93.509
R21538 DVDD.n3148 DVDD.n3111 87.5869
R21539 DVDD.n3149 DVDD.n3148 87.546
R21540 DVDD.t142 DVDD.t21 81.8248
R21541 DVDD.t21 DVDD.t0 81.8248
R21542 DVDD.t93 DVDD.t189 81.8248
R21543 DVDD.t189 DVDD.t150 81.8248
R21544 DVDD.t31 DVDD.t33 81.8248
R21545 DVDD.t33 DVDD.t27 81.8248
R21546 DVDD.t27 DVDD.t29 81.8248
R21547 DVDD.t37 DVDD.t35 81.8248
R21548 DVDD.t35 DVDD.t41 81.8248
R21549 DVDD.t41 DVDD.t39 81.8248
R21550 DVDD.t156 DVDD.t119 81.8248
R21551 DVDD.t119 DVDD.t75 81.8248
R21552 DVDD.t19 DVDD.t14 81.8248
R21553 DVDD.t14 DVDD.t45 81.8248
R21554 DVDD.t45 DVDD.t43 81.8248
R21555 DVDD.t202 DVDD.t98 81.8248
R21556 DVDD.t98 DVDD.t1 81.8248
R21557 DVDD.t1 DVDD.t20 81.8248
R21558 DVDD.t76 DVDD.t127 81.8248
R21559 DVDD.t127 DVDD.t154 81.8248
R21560 DVDD.t135 DVDD.t137 81.8248
R21561 DVDD.t137 DVDD.t121 81.8248
R21562 DVDD.t121 DVDD.t123 81.8248
R21563 DVDD.t71 DVDD.t170 81.8248
R21564 DVDD.t73 DVDD.t71 81.8248
R21565 DVDD.t69 DVDD.t73 81.8248
R21566 DVDD.t144 DVDD.t152 81.8248
R21567 DVDD.t198 DVDD.t144 81.8248
R21568 DVDD.t22 DVDD.t25 81.8248
R21569 DVDD.t125 DVDD.t22 81.8248
R21570 DVDD.n3696 DVDD.t160 73.0276
R21571 DVDD.n3696 DVDD.t15 70.6719
R21572 DVDD.n3215 DVDD.n3116 66.4038
R21573 DVDD.n3216 DVDD.n3215 66.4007
R21574 DVDD.n3224 DVDD.n3109 66.1618
R21575 DVDD.n3224 DVDD.n3223 66.1584
R21576 DVDD.n3148 DVDD.n3112 55.0525
R21577 DVDD.n3148 DVDD.n3147 54.9859
R21578 DVDD.n5492 DVDD.t179 52.7139
R21579 DVDD.n5496 DVDD.t82 52.7139
R21580 DVDD.n5494 DVDD.t100 52.4178
R21581 DVDD.t85 DVDD.n5500 52.4178
R21582 DVDD.n5493 DVDD.t64 51.3813
R21583 DVDD.n5497 DVDD.t195 51.3813
R21584 DVDD.t199 DVDD.n5493 51.0851
R21585 DVDD.n5497 DVDD.t106 51.0851
R21586 DVDD.n5494 DVDD.t103 50.0486
R21587 DVDD.n5500 DVDD.t88 50.0486
R21588 DVDD.t176 DVDD.n5492 49.7525
R21589 DVDD.t79 DVDD.n5496 49.7525
R21590 DVDD.t96 DVDD.n1884 46.6135
R21591 DVDD.t115 DVDD.n4201 46.6135
R21592 DVDD.n2430 DVDD 46.0855
R21593 DVDD.n2596 DVDD.t23 43.2772
R21594 DVDD.n2522 DVDD.n2520 39.6905
R21595 DVDD.n3447 DVDD.t26 39.5713
R21596 DVDD.n1884 DVDD.t142 35.2118
R21597 DVDD.n4201 DVDD.t125 35.2118
R21598 DVDD.n1963 DVDD.t164 34.7933
R21599 DVDD.n1935 DVDD.t174 34.7929
R21600 DVDD.n1933 DVDD.t91 34.7928
R21601 DVDD.n1960 DVDD.t131 31.2268
R21602 DVDD.t64 DVDD.t176 28.4302
R21603 DVDD.t103 DVDD.t199 28.4302
R21604 DVDD.t106 DVDD.t88 28.4302
R21605 DVDD.t195 DVDD.t79 28.4302
R21606 DVDD.n5489 DVDD.t179 25.0246
R21607 DVDD.n5663 DVDD.t82 25.0246
R21608 DVDD.n4149 DVDD.t210 21.0793
R21609 DVDD.n1873 DVDD.t213 21.0793
R21610 DVDD.n3961 DVDD.t217 21.0793
R21611 DVDD.n4139 DVDD.t205 21.0793
R21612 DVDD.n3150 DVDD.n3116 20.9305
R21613 DVDD.n3216 DVDD.n3115 20.9305
R21614 DVDD.n3146 DVDD.n3109 20.7205
R21615 DVDD.n3223 DVDD.n3221 20.7205
R21616 DVDD.n3062 DVDD 19.7447
R21617 DVDD.n3041 DVDD 19.7447
R21618 DVDD.n2997 DVDD 19.7447
R21619 DVDD.n3016 DVDD 19.7447
R21620 DVDD.n5663 DVDD.n5662 19.6523
R21621 DVDD.n5489 DVDD.n5488 19.5041
R21622 DVDD DVDD.t222 19.104
R21623 DVDD.t222 DVDD 19.104
R21624 DVDD DVDD.t209 19.104
R21625 DVDD.t209 DVDD 19.104
R21626 DVDD DVDD.t219 19.104
R21627 DVDD.t219 DVDD 19.104
R21628 DVDD DVDD.t207 19.104
R21629 DVDD.t207 DVDD 19.104
R21630 DVDD DVDD.t218 19.104
R21631 DVDD.t218 DVDD 19.104
R21632 DVDD DVDD.t211 19.104
R21633 DVDD.t211 DVDD 19.104
R21634 DVDD DVDD.t221 19.104
R21635 DVDD.t221 DVDD 19.104
R21636 DVDD.t208 DVDD 19.104
R21637 DVDD DVDD.t208 19.104
R21638 DVDD DVDD.t206 19.104
R21639 DVDD.t206 DVDD 19.104
R21640 DVDD DVDD.t212 19.104
R21641 DVDD.t212 DVDD 19.104
R21642 DVDD.n3217 DVDD.n3216 14.6999
R21643 DVDD.n3152 DVDD.n3116 14.6999
R21644 DVDD.n3223 DVDD.n3110 14.6413
R21645 DVDD.n3143 DVDD.n3109 14.6413
R21646 DVDD.n3063 DVDD 14.3168
R21647 DVDD.n3042 DVDD 14.3168
R21648 DVDD.n2998 DVDD 14.3168
R21649 DVDD.n3017 DVDD 14.3168
R21650 DVDD.n5501 DVDD.t85 14.2154
R21651 DVDD.t100 DVDD.n261 12.8827
R21652 DVDD.n5488 DVDD.n5487 12.4047
R21653 DVDD.n5662 DVDD.n5661 12.3937
R21654 DVDD.n2687 DVDD.n2685 9.73503
R21655 DVDD DVDD.t220 7.42907
R21656 DVDD DVDD.t215 7.42907
R21657 DVDD DVDD.t216 7.42907
R21658 DVDD DVDD.t214 7.42907
R21659 DVDD.n3446 DVDD.n2687 7.19237
R21660 DVDD.n2512 DVDD.t182 6.5562
R21661 DVDD.n2574 DVDD.n2573 6.3005
R21662 DVDD.n2580 DVDD.n2551 6.3005
R21663 DVDD.n2582 DVDD.n2551 6.3005
R21664 DVDD.n2588 DVDD.n2528 6.3005
R21665 DVDD.n2591 DVDD.n2528 6.3005
R21666 DVDD.n2593 DVDD.n2528 6.3005
R21667 DVDD.n2574 DVDD.n2553 6.3005
R21668 DVDD.n2557 DVDD.n2553 6.3005
R21669 DVDD.n2560 DVDD.n2553 6.3005
R21670 DVDD.n2556 DVDD.n2553 6.3005
R21671 DVDD.n2580 DVDD.n2553 6.3005
R21672 DVDD.n2582 DVDD.n2553 6.3005
R21673 DVDD.n2542 DVDD.n2530 6.3005
R21674 DVDD.n2591 DVDD.n2530 6.3005
R21675 DVDD.n2593 DVDD.n2530 6.3005
R21676 DVDD.n2574 DVDD.n2550 6.3005
R21677 DVDD.n2557 DVDD.n2550 6.3005
R21678 DVDD.n2560 DVDD.n2550 6.3005
R21679 DVDD.n2556 DVDD.n2550 6.3005
R21680 DVDD.n2580 DVDD.n2550 6.3005
R21681 DVDD.n2582 DVDD.n2550 6.3005
R21682 DVDD.n2542 DVDD.n2527 6.3005
R21683 DVDD.n2593 DVDD.n2527 6.3005
R21684 DVDD.n2574 DVDD.n2532 6.3005
R21685 DVDD.n2557 DVDD.n2532 6.3005
R21686 DVDD.n2560 DVDD.n2532 6.3005
R21687 DVDD.n2556 DVDD.n2532 6.3005
R21688 DVDD.n2580 DVDD.n2532 6.3005
R21689 DVDD.n2582 DVDD.n2532 6.3005
R21690 DVDD.n2591 DVDD.n2532 6.3005
R21691 DVDD.n2593 DVDD.n2532 6.3005
R21692 DVDD.n2574 DVDD.n2549 6.3005
R21693 DVDD.n2557 DVDD.n2549 6.3005
R21694 DVDD.n2560 DVDD.n2549 6.3005
R21695 DVDD.n2556 DVDD.n2549 6.3005
R21696 DVDD.n2580 DVDD.n2549 6.3005
R21697 DVDD.n2582 DVDD.n2549 6.3005
R21698 DVDD.n2542 DVDD.n2526 6.3005
R21699 DVDD.n2591 DVDD.n2526 6.3005
R21700 DVDD.n2593 DVDD.n2526 6.3005
R21701 DVDD.n2574 DVDD.n2554 6.3005
R21702 DVDD.n2557 DVDD.n2554 6.3005
R21703 DVDD.n2560 DVDD.n2554 6.3005
R21704 DVDD.n2556 DVDD.n2554 6.3005
R21705 DVDD.n2580 DVDD.n2554 6.3005
R21706 DVDD.n2582 DVDD.n2554 6.3005
R21707 DVDD.n2542 DVDD.n2533 6.3005
R21708 DVDD.n2591 DVDD.n2533 6.3005
R21709 DVDD.n2593 DVDD.n2533 6.3005
R21710 DVDD.n2574 DVDD.n2548 6.3005
R21711 DVDD.n2557 DVDD.n2548 6.3005
R21712 DVDD.n2560 DVDD.n2548 6.3005
R21713 DVDD.n2556 DVDD.n2548 6.3005
R21714 DVDD.n2580 DVDD.n2548 6.3005
R21715 DVDD.n2582 DVDD.n2548 6.3005
R21716 DVDD.n2542 DVDD.n2525 6.3005
R21717 DVDD.n2591 DVDD.n2525 6.3005
R21718 DVDD.n2593 DVDD.n2525 6.3005
R21719 DVDD.n2581 DVDD.n2557 6.3005
R21720 DVDD.n2581 DVDD.n2560 6.3005
R21721 DVDD.n2581 DVDD.n2556 6.3005
R21722 DVDD.n2581 DVDD.n2580 6.3005
R21723 DVDD.n2582 DVDD.n2581 6.3005
R21724 DVDD.n2592 DVDD.n2542 6.3005
R21725 DVDD.n2592 DVDD.n2591 6.3005
R21726 DVDD.n2592 DVDD.n2538 6.3005
R21727 DVDD.n2593 DVDD.n2592 6.3005
R21728 DVDD.n5499 DVDD.n5495 5.57024
R21729 DVDD.n3145 DVDD.n3143 5.56181
R21730 DVDD.n3220 DVDD.n3110 5.56181
R21731 DVDD.n5491 DVDD.n262 5.41553
R21732 DVDD.n5495 DVDD.n262 5.41553
R21733 DVDD.n5499 DVDD.n5498 5.41553
R21734 DVDD.n5498 DVDD.n256 5.41553
R21735 DVDD.n3217 DVDD.n3113 5.21853
R21736 DVDD.n3152 DVDD.n3151 5.21853
R21737 DVDD.n3153 DVDD.n3144 4.9705
R21738 DVDD.n3219 DVDD.n3218 4.9005
R21739 DVDD.n3398 DVDD.n3397 4.66866
R21740 DVDD.n3407 DVDD.n2725 4.66866
R21741 DVDD.n3434 DVDD.n3433 4.66866
R21742 DVDD.n1682 DVDD.n1675 4.66866
R21743 DVDD.n3817 DVDD.n1836 4.66866
R21744 DVDD.n4067 DVDD.n4054 4.66866
R21745 DVDD.n1761 DVDD.n1730 4.66866
R21746 DVDD.n2521 DVDD.t95 4.51467
R21747 DVDD.n2950 DVDD.n2949 4.5005
R21748 DVDD.n2950 DVDD.n2934 4.5005
R21749 DVDD.n2952 DVDD.n2934 4.5005
R21750 DVDD.n2951 DVDD.n2950 4.5005
R21751 DVDD.n2952 DVDD.n2951 4.5005
R21752 DVDD.n3274 DVDD.n2953 4.5005
R21753 DVDD.n2956 DVDD.n2953 4.5005
R21754 DVDD.n2956 DVDD.n2955 4.5005
R21755 DVDD.n2957 DVDD.n2953 4.5005
R21756 DVDD.n2957 DVDD.n2955 4.5005
R21757 DVDD.n3123 DVDD.n3122 4.5005
R21758 DVDD.n3252 DVDD.n3251 4.5005
R21759 DVDD.n3205 DVDD.n3122 4.5005
R21760 DVDD.n3250 DVDD.n3085 4.5005
R21761 DVDD.n3251 DVDD.n3250 4.5005
R21762 DVDD.n3206 DVDD.n3123 4.5005
R21763 DVDD.n3206 DVDD.n3205 4.5005
R21764 DVDD.n3252 DVDD.n3085 4.5005
R21765 DVDD.n3114 DVDD.n3096 4.5005
R21766 DVDD.n3163 DVDD.n3154 4.5005
R21767 DVDD.n3163 DVDD.n3155 4.5005
R21768 DVDD.n3229 DVDD.n3096 4.5005
R21769 DVDD.n2609 DVDD.n2507 4.5005
R21770 DVDD.n2609 DVDD.n2608 4.5005
R21771 DVDD.n2608 DVDD.n2509 4.5005
R21772 DVDD.n2607 DVDD.n2605 4.5005
R21773 DVDD.n2608 DVDD.n2607 4.5005
R21774 DVDD.n2647 DVDD.n2646 4.5005
R21775 DVDD.n2647 DVDD.n2626 4.5005
R21776 DVDD.n2645 DVDD.n2626 4.5005
R21777 DVDD.n2650 DVDD.n2626 4.5005
R21778 DVDD.n2650 DVDD.n2649 4.5005
R21779 DVDD.n2447 DVDD.n2442 4.5005
R21780 DVDD.n3603 DVDD.n2447 4.5005
R21781 DVDD.n3601 DVDD.n2447 4.5005
R21782 DVDD.n3601 DVDD.n2449 4.5005
R21783 DVDD.n3603 DVDD.n2449 4.5005
R21784 DVDD.n2449 DVDD.n2442 4.5005
R21785 DVDD.n2446 DVDD.n2442 4.5005
R21786 DVDD.n3603 DVDD.n2446 4.5005
R21787 DVDD.n3601 DVDD.n2446 4.5005
R21788 DVDD.n2450 DVDD.n2442 4.5005
R21789 DVDD.n3603 DVDD.n2450 4.5005
R21790 DVDD.n3601 DVDD.n2450 4.5005
R21791 DVDD.n3601 DVDD.n2445 4.5005
R21792 DVDD.n3603 DVDD.n2445 4.5005
R21793 DVDD.n2445 DVDD.n2442 4.5005
R21794 DVDD.n2451 DVDD.n2442 4.5005
R21795 DVDD.n3603 DVDD.n2451 4.5005
R21796 DVDD.n3601 DVDD.n2451 4.5005
R21797 DVDD.n2444 DVDD.n2442 4.5005
R21798 DVDD.n3603 DVDD.n2444 4.5005
R21799 DVDD.n3601 DVDD.n2444 4.5005
R21800 DVDD.n3601 DVDD.n2452 4.5005
R21801 DVDD.n3603 DVDD.n2452 4.5005
R21802 DVDD.n2452 DVDD.n2442 4.5005
R21803 DVDD.n3601 DVDD.n2443 4.5005
R21804 DVDD.n3603 DVDD.n2443 4.5005
R21805 DVDD.n2443 DVDD.n2442 4.5005
R21806 DVDD.n3602 DVDD.n2442 4.5005
R21807 DVDD.n3603 DVDD.n3602 4.5005
R21808 DVDD.n3602 DVDD.n3601 4.5005
R21809 DVDD.n3526 DVDD.n2494 4.5005
R21810 DVDD.n2500 DVDD.n2494 4.5005
R21811 DVDD.n3528 DVDD.n2494 4.5005
R21812 DVDD.n3526 DVDD.n2496 4.5005
R21813 DVDD.n2500 DVDD.n2496 4.5005
R21814 DVDD.n3528 DVDD.n2496 4.5005
R21815 DVDD.n3528 DVDD.n2493 4.5005
R21816 DVDD.n2500 DVDD.n2493 4.5005
R21817 DVDD.n3526 DVDD.n2493 4.5005
R21818 DVDD.n3526 DVDD.n2497 4.5005
R21819 DVDD.n2500 DVDD.n2497 4.5005
R21820 DVDD.n3528 DVDD.n2497 4.5005
R21821 DVDD.n3526 DVDD.n2492 4.5005
R21822 DVDD.n2500 DVDD.n2492 4.5005
R21823 DVDD.n3528 DVDD.n2492 4.5005
R21824 DVDD.n3528 DVDD.n2498 4.5005
R21825 DVDD.n2500 DVDD.n2498 4.5005
R21826 DVDD.n3526 DVDD.n2498 4.5005
R21827 DVDD.n3526 DVDD.n2491 4.5005
R21828 DVDD.n2500 DVDD.n2491 4.5005
R21829 DVDD.n3528 DVDD.n2491 4.5005
R21830 DVDD.n3528 DVDD.n3527 4.5005
R21831 DVDD.n3527 DVDD.n2500 4.5005
R21832 DVDD.n3527 DVDD.n3526 4.5005
R21833 DVDD.n3433 DVDD.n3432 4.5005
R21834 DVDD.n2698 DVDD.n2697 4.5005
R21835 DVDD.n3423 DVDD.n3422 4.5005
R21836 DVDD.n3421 DVDD.n2703 4.5005
R21837 DVDD.n3419 DVDD.n3418 4.5005
R21838 DVDD.n3410 DVDD.n2705 4.5005
R21839 DVDD.n3409 DVDD.n3408 4.5005
R21840 DVDD.n3407 DVDD.n3406 4.5005
R21841 DVDD.n3397 DVDD.n2729 4.5005
R21842 DVDD.n3396 DVDD.n3395 4.5005
R21843 DVDD.n2732 DVDD.n2731 4.5005
R21844 DVDD.n2985 DVDD.n2984 4.5005
R21845 DVDD.n2982 DVDD.n2981 4.5005
R21846 DVDD.n2967 DVDD.n2966 4.5005
R21847 DVDD.n2973 DVDD.n2972 4.5005
R21848 DVDD.n3210 DVDD.n3209 4.5005
R21849 DVDD.n3135 DVDD.n3134 4.5005
R21850 DVDD.n3187 DVDD.n3182 4.5005
R21851 DVDD.n3183 DVDD.n3130 4.5005
R21852 DVDD.n3197 DVDD.n3196 4.5005
R21853 DVDD.n3131 DVDD.n2986 4.5005
R21854 DVDD.n3211 DVDD.n3210 4.5005
R21855 DVDD.n3134 DVDD.n3098 4.5005
R21856 DVDD.n3187 DVDD.n3186 4.5005
R21857 DVDD.n3183 DVDD.n3093 4.5005
R21858 DVDD.n3196 DVDD.n3090 4.5005
R21859 DVDD.n3082 DVDD.n2986 4.5005
R21860 DVDD.n2870 DVDD.n2861 4.5005
R21861 DVDD.n2873 DVDD.n2861 4.5005
R21862 DVDD.n2863 DVDD.n2861 4.5005
R21863 DVDD.n2879 DVDD.n2861 4.5005
R21864 DVDD.n2864 DVDD.n2861 4.5005
R21865 DVDD.n2878 DVDD.n2861 4.5005
R21866 DVDD.n2865 DVDD.n2861 4.5005
R21867 DVDD.n2877 DVDD.n2861 4.5005
R21868 DVDD.n2866 DVDD.n2861 4.5005
R21869 DVDD.n2876 DVDD.n2861 4.5005
R21870 DVDD.n2867 DVDD.n2861 4.5005
R21871 DVDD.n2875 DVDD.n2861 4.5005
R21872 DVDD.n2868 DVDD.n2861 4.5005
R21873 DVDD.n2874 DVDD.n2861 4.5005
R21874 DVDD.n2869 DVDD.n2861 4.5005
R21875 DVDD.n3342 DVDD.n2861 4.5005
R21876 DVDD.n3341 DVDD.n2871 4.5005
R21877 DVDD.n3341 DVDD.n2873 4.5005
R21878 DVDD.n3341 DVDD.n2870 4.5005
R21879 DVDD.n3342 DVDD.n2859 4.5005
R21880 DVDD.n2869 DVDD.n2859 4.5005
R21881 DVDD.n2874 DVDD.n2859 4.5005
R21882 DVDD.n2868 DVDD.n2859 4.5005
R21883 DVDD.n2875 DVDD.n2859 4.5005
R21884 DVDD.n2867 DVDD.n2859 4.5005
R21885 DVDD.n2876 DVDD.n2859 4.5005
R21886 DVDD.n2866 DVDD.n2859 4.5005
R21887 DVDD.n2877 DVDD.n2859 4.5005
R21888 DVDD.n2865 DVDD.n2859 4.5005
R21889 DVDD.n2878 DVDD.n2859 4.5005
R21890 DVDD.n2864 DVDD.n2859 4.5005
R21891 DVDD.n2879 DVDD.n2859 4.5005
R21892 DVDD.n2863 DVDD.n2859 4.5005
R21893 DVDD.n3340 DVDD.n2859 4.5005
R21894 DVDD.n2871 DVDD.n2859 4.5005
R21895 DVDD.n2873 DVDD.n2859 4.5005
R21896 DVDD.n2870 DVDD.n2859 4.5005
R21897 DVDD.n3342 DVDD.n3341 4.5005
R21898 DVDD.n3341 DVDD.n2869 4.5005
R21899 DVDD.n3341 DVDD.n2874 4.5005
R21900 DVDD.n3341 DVDD.n2868 4.5005
R21901 DVDD.n3341 DVDD.n2875 4.5005
R21902 DVDD.n3341 DVDD.n2867 4.5005
R21903 DVDD.n3341 DVDD.n2876 4.5005
R21904 DVDD.n3341 DVDD.n2866 4.5005
R21905 DVDD.n3341 DVDD.n2877 4.5005
R21906 DVDD.n3341 DVDD.n2865 4.5005
R21907 DVDD.n3341 DVDD.n2878 4.5005
R21908 DVDD.n3341 DVDD.n2864 4.5005
R21909 DVDD.n3341 DVDD.n2879 4.5005
R21910 DVDD.n3341 DVDD.n2863 4.5005
R21911 DVDD.n3341 DVDD.n3340 4.5005
R21912 DVDD.n3347 DVDD.n3346 4.5005
R21913 DVDD.n3346 DVDD.n2781 4.5005
R21914 DVDD.n3346 DVDD.n2797 4.5005
R21915 DVDD.n3346 DVDD.n2782 4.5005
R21916 DVDD.n3346 DVDD.n2796 4.5005
R21917 DVDD.n3346 DVDD.n2783 4.5005
R21918 DVDD.n3346 DVDD.n2795 4.5005
R21919 DVDD.n3346 DVDD.n2784 4.5005
R21920 DVDD.n3346 DVDD.n2794 4.5005
R21921 DVDD.n3346 DVDD.n2785 4.5005
R21922 DVDD.n3346 DVDD.n2793 4.5005
R21923 DVDD.n3346 DVDD.n2786 4.5005
R21924 DVDD.n3346 DVDD.n2792 4.5005
R21925 DVDD.n3346 DVDD.n2787 4.5005
R21926 DVDD.n3346 DVDD.n2790 4.5005
R21927 DVDD.n3346 DVDD.n2789 4.5005
R21928 DVDD.n3347 DVDD.n2799 4.5005
R21929 DVDD.n2799 DVDD.n2781 4.5005
R21930 DVDD.n2799 DVDD.n2797 4.5005
R21931 DVDD.n2799 DVDD.n2782 4.5005
R21932 DVDD.n2799 DVDD.n2796 4.5005
R21933 DVDD.n2799 DVDD.n2783 4.5005
R21934 DVDD.n2799 DVDD.n2795 4.5005
R21935 DVDD.n2799 DVDD.n2784 4.5005
R21936 DVDD.n2799 DVDD.n2794 4.5005
R21937 DVDD.n2799 DVDD.n2785 4.5005
R21938 DVDD.n2799 DVDD.n2793 4.5005
R21939 DVDD.n2799 DVDD.n2786 4.5005
R21940 DVDD.n2799 DVDD.n2792 4.5005
R21941 DVDD.n2799 DVDD.n2787 4.5005
R21942 DVDD.n2799 DVDD.n2791 4.5005
R21943 DVDD.n2799 DVDD.n2788 4.5005
R21944 DVDD.n2799 DVDD.n2790 4.5005
R21945 DVDD.n2799 DVDD.n2789 4.5005
R21946 DVDD.n3348 DVDD.n2789 4.5005
R21947 DVDD.n3348 DVDD.n2790 4.5005
R21948 DVDD.n3348 DVDD.n2788 4.5005
R21949 DVDD.n3348 DVDD.n2791 4.5005
R21950 DVDD.n3348 DVDD.n2787 4.5005
R21951 DVDD.n3348 DVDD.n2792 4.5005
R21952 DVDD.n3348 DVDD.n2786 4.5005
R21953 DVDD.n3348 DVDD.n2793 4.5005
R21954 DVDD.n3348 DVDD.n2785 4.5005
R21955 DVDD.n3348 DVDD.n2794 4.5005
R21956 DVDD.n3348 DVDD.n2784 4.5005
R21957 DVDD.n3348 DVDD.n2795 4.5005
R21958 DVDD.n3348 DVDD.n2783 4.5005
R21959 DVDD.n3348 DVDD.n2796 4.5005
R21960 DVDD.n3348 DVDD.n2782 4.5005
R21961 DVDD.n3348 DVDD.n2797 4.5005
R21962 DVDD.n3348 DVDD.n2781 4.5005
R21963 DVDD.n3348 DVDD.n3347 4.5005
R21964 DVDD.n4068 DVDD.n4067 4.5005
R21965 DVDD.n4066 DVDD.n4065 4.5005
R21966 DVDD.n4057 DVDD.n4056 4.5005
R21967 DVDD.n4058 DVDD.n1719 4.5005
R21968 DVDD.n4228 DVDD.n4227 4.5005
R21969 DVDD.n1728 DVDD.n1720 4.5005
R21970 DVDD.n1763 DVDD.n1762 4.5005
R21971 DVDD.n1761 DVDD.n1760 4.5005
R21972 DVDD.n1682 DVDD.n1680 4.5005
R21973 DVDD.n4267 DVDD.n4266 4.5005
R21974 DVDD.n4265 DVDD.n4264 4.5005
R21975 DVDD.n1684 DVDD.n1683 4.5005
R21976 DVDD.n1843 DVDD.n1842 4.5005
R21977 DVDD.n3815 DVDD.n3814 4.5005
R21978 DVDD.n3816 DVDD.n1840 4.5005
R21979 DVDD.n3818 DVDD.n3817 4.5005
R21980 DVDD.n3779 DVDD.n1887 4.5005
R21981 DVDD.n3779 DVDD.n1861 4.5005
R21982 DVDD.n3779 DVDD.n3778 4.5005
R21983 DVDD.n3675 DVDD.n1982 4.5005
R21984 DVDD.n3675 DVDD.n3674 4.5005
R21985 DVDD.n3674 DVDD.n1990 4.5005
R21986 DVDD.n3674 DVDD.n1987 4.5005
R21987 DVDD.n3674 DVDD.n1992 4.5005
R21988 DVDD.n3674 DVDD.n1986 4.5005
R21989 DVDD.n3674 DVDD.n1994 4.5005
R21990 DVDD.n3674 DVDD.n1985 4.5005
R21991 DVDD.n3674 DVDD.n1996 4.5005
R21992 DVDD.n3674 DVDD.n1984 4.5005
R21993 DVDD.n3673 DVDD.n1982 4.5005
R21994 DVDD.n3674 DVDD.n3673 4.5005
R21995 DVDD.n2405 DVDD.n1997 4.5005
R21996 DVDD.n2405 DVDD.n2404 4.5005
R21997 DVDD.n2404 DVDD.n2006 4.5005
R21998 DVDD.n2404 DVDD.n2003 4.5005
R21999 DVDD.n2404 DVDD.n2008 4.5005
R22000 DVDD.n2404 DVDD.n2002 4.5005
R22001 DVDD.n2404 DVDD.n2010 4.5005
R22002 DVDD.n2404 DVDD.n2001 4.5005
R22003 DVDD.n2404 DVDD.n2012 4.5005
R22004 DVDD.n2404 DVDD.n2000 4.5005
R22005 DVDD.n2403 DVDD.n1997 4.5005
R22006 DVDD.n2404 DVDD.n2403 4.5005
R22007 DVDD.n3778 DVDD.n3777 4.5005
R22008 DVDD.n3777 DVDD.n3732 4.5005
R22009 DVDD.n3777 DVDD.n3737 4.5005
R22010 DVDD.n3777 DVDD.n3731 4.5005
R22011 DVDD.n3777 DVDD.n3738 4.5005
R22012 DVDD.n3777 DVDD.n3730 4.5005
R22013 DVDD.n3777 DVDD.n3739 4.5005
R22014 DVDD.n3777 DVDD.n3729 4.5005
R22015 DVDD.n3777 DVDD.n3740 4.5005
R22016 DVDD.n3777 DVDD.n1861 4.5005
R22017 DVDD.n3777 DVDD.n1887 4.5005
R22018 DVDD.n3777 DVDD.n3728 4.5005
R22019 DVDD.n3777 DVDD.n3741 4.5005
R22020 DVDD.n3777 DVDD.n3727 4.5005
R22021 DVDD.n3777 DVDD.n3742 4.5005
R22022 DVDD.n3777 DVDD.n3726 4.5005
R22023 DVDD.n3777 DVDD.n3743 4.5005
R22024 DVDD.n3777 DVDD.n3725 4.5005
R22025 DVDD.n3777 DVDD.n3744 4.5005
R22026 DVDD.n3777 DVDD.n3724 4.5005
R22027 DVDD.n3776 DVDD.n3754 4.5005
R22028 DVDD.n3777 DVDD.n3776 4.5005
R22029 DVDD.n1323 DVDD.n1321 4.5005
R22030 DVDD.n1388 DVDD.n1383 4.5005
R22031 DVDD.n1388 DVDD.n1385 4.5005
R22032 DVDD.n1323 DVDD.n1322 4.5005
R22033 DVDD.n1388 DVDD.n1382 4.5005
R22034 DVDD.n1382 DVDD.n1380 4.5005
R22035 DVDD.n1325 DVDD.n1318 4.5005
R22036 DVDD.n1323 DVDD.n1318 4.5005
R22037 DVDD.n1388 DVDD.n1386 4.5005
R22038 DVDD.n1386 DVDD.n1380 4.5005
R22039 DVDD.n1325 DVDD.n1320 4.5005
R22040 DVDD.n1323 DVDD.n1320 4.5005
R22041 DVDD.n1325 DVDD.n1317 4.5005
R22042 DVDD.n1323 DVDD.n1317 4.5005
R22043 DVDD.n1381 DVDD.n1380 4.5005
R22044 DVDD.n1388 DVDD.n1381 4.5005
R22045 DVDD.n1325 DVDD.n1324 4.5005
R22046 DVDD.n1324 DVDD.n1323 4.5005
R22047 DVDD.n1387 DVDD.n1380 4.5005
R22048 DVDD.n1388 DVDD.n1387 4.5005
R22049 DVDD.n1365 DVDD.n1331 4.5005
R22050 DVDD.n1332 DVDD.n1331 4.5005
R22051 DVDD.n1369 DVDD.n1331 4.5005
R22052 DVDD.n1394 DVDD.n1309 4.5005
R22053 DVDD.n1394 DVDD.n1311 4.5005
R22054 DVDD.n1394 DVDD.n1308 4.5005
R22055 DVDD.n1312 DVDD.n1305 4.5005
R22056 DVDD.n1394 DVDD.n1312 4.5005
R22057 DVDD.n1307 DVDD.n1305 4.5005
R22058 DVDD.n1394 DVDD.n1307 4.5005
R22059 DVDD.n1313 DVDD.n1305 4.5005
R22060 DVDD.n1394 DVDD.n1313 4.5005
R22061 DVDD.n1306 DVDD.n1305 4.5005
R22062 DVDD.n1394 DVDD.n1306 4.5005
R22063 DVDD.n1308 DVDD.n1305 4.5005
R22064 DVDD.n1311 DVDD.n1305 4.5005
R22065 DVDD.n1309 DVDD.n1305 4.5005
R22066 DVDD.n1393 DVDD.n1305 4.5005
R22067 DVDD.n1394 DVDD.n1393 4.5005
R22068 DVDD.n1554 DVDD.n1214 4.5005
R22069 DVDD.n1554 DVDD.n1221 4.5005
R22070 DVDD.n1554 DVDD.n1215 4.5005
R22071 DVDD.n1556 DVDD.n1217 4.5005
R22072 DVDD.n1554 DVDD.n1217 4.5005
R22073 DVDD.n1556 DVDD.n1219 4.5005
R22074 DVDD.n1554 DVDD.n1219 4.5005
R22075 DVDD.n1556 DVDD.n1216 4.5005
R22076 DVDD.n1554 DVDD.n1216 4.5005
R22077 DVDD.n1556 DVDD.n1220 4.5005
R22078 DVDD.n1554 DVDD.n1220 4.5005
R22079 DVDD.n1556 DVDD.n1215 4.5005
R22080 DVDD.n1556 DVDD.n1221 4.5005
R22081 DVDD.n1556 DVDD.n1214 4.5005
R22082 DVDD.n1556 DVDD.n1555 4.5005
R22083 DVDD.n1555 DVDD.n1554 4.5005
R22084 DVDD.n1364 DVDD.n1329 4.5005
R22085 DVDD.n1364 DVDD.n1336 4.5005
R22086 DVDD.n1368 DVDD.n1336 4.5005
R22087 DVDD.n1368 DVDD.n1339 4.5005
R22088 DVDD.n1368 DVDD.n1335 4.5005
R22089 DVDD.n1368 DVDD.n1329 4.5005
R22090 DVDD.n1369 DVDD.n1368 4.5005
R22091 DVDD.n1368 DVDD.n1367 4.5005
R22092 DVDD.n1367 DVDD.n1331 4.5005
R22093 DVDD.n1195 DVDD.n1192 4.5005
R22094 DVDD.n1200 DVDD.n1192 4.5005
R22095 DVDD.n1577 DVDD.n1192 4.5005
R22096 DVDD.n1577 DVDD.n1576 4.5005
R22097 DVDD.n1576 DVDD.n1199 4.5005
R22098 DVDD.n1576 DVDD.n1196 4.5005
R22099 DVDD.n1576 DVDD.n1200 4.5005
R22100 DVDD.n1576 DVDD.n1195 4.5005
R22101 DVDD.n1576 DVDD.n1202 4.5005
R22102 DVDD.n1576 DVDD.n1194 4.5005
R22103 DVDD.n1576 DVDD.n1575 4.5005
R22104 DVDD.n1575 DVDD.n1192 4.5005
R22105 DVDD.n5424 DVDD.n341 4.5005
R22106 DVDD.n5917 DVDD.n5916 4.5005
R22107 DVDD.n5422 DVDD.n5419 4.5005
R22108 DVDD.n5919 DVDD.n94 4.5005
R22109 DVDD.n5424 DVDD.n342 4.5005
R22110 DVDD.n350 DVDD.n342 4.5005
R22111 DVDD.n5422 DVDD.n342 4.5005
R22112 DVDD.n5917 DVDD.n95 4.5005
R22113 DVDD.n105 DVDD.n95 4.5005
R22114 DVDD.n5919 DVDD.n95 4.5005
R22115 DVDD.n350 DVDD.n347 4.5005
R22116 DVDD.n5422 DVDD.n347 4.5005
R22117 DVDD.n5917 DVDD.n93 4.5005
R22118 DVDD.n350 DVDD.n335 4.5005
R22119 DVDD.n5422 DVDD.n335 4.5005
R22120 DVDD.n5917 DVDD.n96 4.5005
R22121 DVDD.n350 DVDD.n346 4.5005
R22122 DVDD.n5422 DVDD.n346 4.5005
R22123 DVDD.n5917 DVDD.n92 4.5005
R22124 DVDD.n350 DVDD.n336 4.5005
R22125 DVDD.n5422 DVDD.n336 4.5005
R22126 DVDD.n5917 DVDD.n97 4.5005
R22127 DVDD.n350 DVDD.n345 4.5005
R22128 DVDD.n5422 DVDD.n345 4.5005
R22129 DVDD.n5917 DVDD.n91 4.5005
R22130 DVDD.n350 DVDD.n337 4.5005
R22131 DVDD.n5917 DVDD.n98 4.5005
R22132 DVDD.n350 DVDD.n344 4.5005
R22133 DVDD.n5917 DVDD.n90 4.5005
R22134 DVDD.n350 DVDD.n338 4.5005
R22135 DVDD.n5422 DVDD.n338 4.5005
R22136 DVDD.n5917 DVDD.n99 4.5005
R22137 DVDD.n350 DVDD.n343 4.5005
R22138 DVDD.n5422 DVDD.n343 4.5005
R22139 DVDD.n5917 DVDD.n89 4.5005
R22140 DVDD.n350 DVDD.n339 4.5005
R22141 DVDD.n5422 DVDD.n339 4.5005
R22142 DVDD.n5917 DVDD.n100 4.5005
R22143 DVDD.n5424 DVDD.n339 4.5005
R22144 DVDD.n5424 DVDD.n343 4.5005
R22145 DVDD.n5424 DVDD.n338 4.5005
R22146 DVDD.n5424 DVDD.n344 4.5005
R22147 DVDD.n5424 DVDD.n337 4.5005
R22148 DVDD.n5424 DVDD.n345 4.5005
R22149 DVDD.n5424 DVDD.n336 4.5005
R22150 DVDD.n5424 DVDD.n346 4.5005
R22151 DVDD.n5424 DVDD.n335 4.5005
R22152 DVDD.n5424 DVDD.n347 4.5005
R22153 DVDD.n105 DVDD.n93 4.5005
R22154 DVDD.n5919 DVDD.n93 4.5005
R22155 DVDD.n105 DVDD.n96 4.5005
R22156 DVDD.n5919 DVDD.n96 4.5005
R22157 DVDD.n105 DVDD.n92 4.5005
R22158 DVDD.n5919 DVDD.n92 4.5005
R22159 DVDD.n105 DVDD.n97 4.5005
R22160 DVDD.n5919 DVDD.n97 4.5005
R22161 DVDD.n105 DVDD.n91 4.5005
R22162 DVDD.n5919 DVDD.n91 4.5005
R22163 DVDD.n5919 DVDD.n98 4.5005
R22164 DVDD.n5919 DVDD.n90 4.5005
R22165 DVDD.n105 DVDD.n99 4.5005
R22166 DVDD.n5919 DVDD.n99 4.5005
R22167 DVDD.n105 DVDD.n89 4.5005
R22168 DVDD.n5919 DVDD.n89 4.5005
R22169 DVDD.n105 DVDD.n100 4.5005
R22170 DVDD.n5919 DVDD.n100 4.5005
R22171 DVDD.n5919 DVDD.n88 4.5005
R22172 DVDD.n5917 DVDD.n88 4.5005
R22173 DVDD.n5422 DVDD.n334 4.5005
R22174 DVDD.n5424 DVDD.n334 4.5005
R22175 DVDD.n5919 DVDD.n5918 4.5005
R22176 DVDD.n5918 DVDD.n5917 4.5005
R22177 DVDD.n5423 DVDD.n5422 4.5005
R22178 DVDD.n5424 DVDD.n5423 4.5005
R22179 DVDD.n5429 DVDD.n327 4.5005
R22180 DVDD.n327 DVDD.n321 4.5005
R22181 DVDD.n5429 DVDD.n5428 4.5005
R22182 DVDD.n5428 DVDD.n321 4.5005
R22183 DVDD.n5429 DVDD.n326 4.5005
R22184 DVDD.n326 DVDD.n321 4.5005
R22185 DVDD.n5921 DVDD.n77 4.5005
R22186 DVDD.n5921 DVDD.n79 4.5005
R22187 DVDD.n81 DVDD.n77 4.5005
R22188 DVDD.n81 DVDD.n79 4.5005
R22189 DVDD.n5923 DVDD.n77 4.5005
R22190 DVDD.n5923 DVDD.n79 4.5005
R22191 DVDD.n1578 DVDD.n1120 4.5005
R22192 DVDD.n1579 DVDD.n1578 4.5005
R22193 DVDD.n1189 DVDD.n1120 4.5005
R22194 DVDD.n1582 DVDD.n1134 4.5005
R22195 DVDD.n1582 DVDD.n1130 4.5005
R22196 DVDD.n1582 DVDD.n1136 4.5005
R22197 DVDD.n1582 DVDD.n1129 4.5005
R22198 DVDD.n1582 DVDD.n1138 4.5005
R22199 DVDD.n1582 DVDD.n1128 4.5005
R22200 DVDD.n1582 DVDD.n1140 4.5005
R22201 DVDD.n1582 DVDD.n1127 4.5005
R22202 DVDD.n1582 DVDD.n1142 4.5005
R22203 DVDD.n1582 DVDD.n1126 4.5005
R22204 DVDD.n1582 DVDD.n1144 4.5005
R22205 DVDD.n1582 DVDD.n1125 4.5005
R22206 DVDD.n1582 DVDD.n1146 4.5005
R22207 DVDD.n1582 DVDD.n1124 4.5005
R22208 DVDD.n1582 DVDD.n1148 4.5005
R22209 DVDD.n1582 DVDD.n1123 4.5005
R22210 DVDD.n1582 DVDD.n1581 4.5005
R22211 DVDD.n1582 DVDD.n1122 4.5005
R22212 DVDD.n1583 DVDD.n1120 4.5005
R22213 DVDD.n1583 DVDD.n1582 4.5005
R22214 DVDD.n5381 DVDD.n378 4.5005
R22215 DVDD.n5383 DVDD.n378 4.5005
R22216 DVDD.n5381 DVDD.n380 4.5005
R22217 DVDD.n5383 DVDD.n380 4.5005
R22218 DVDD.n5381 DVDD.n377 4.5005
R22219 DVDD.n5383 DVDD.n377 4.5005
R22220 DVDD.n5382 DVDD.n5381 4.5005
R22221 DVDD.n5383 DVDD.n5382 4.5005
R22222 DVDD.n5361 DVDD.n401 4.5005
R22223 DVDD.n5363 DVDD.n401 4.5005
R22224 DVDD.n5361 DVDD.n403 4.5005
R22225 DVDD.n5363 DVDD.n403 4.5005
R22226 DVDD.n5361 DVDD.n400 4.5005
R22227 DVDD.n5363 DVDD.n400 4.5005
R22228 DVDD.n5362 DVDD.n5361 4.5005
R22229 DVDD.n5363 DVDD.n5362 4.5005
R22230 DVDD.n5340 DVDD.n425 4.5005
R22231 DVDD.n5342 DVDD.n425 4.5005
R22232 DVDD.n5340 DVDD.n427 4.5005
R22233 DVDD.n5342 DVDD.n427 4.5005
R22234 DVDD.n5340 DVDD.n424 4.5005
R22235 DVDD.n5342 DVDD.n424 4.5005
R22236 DVDD.n5341 DVDD.n5340 4.5005
R22237 DVDD.n5342 DVDD.n5341 4.5005
R22238 DVDD.n5136 DVDD.n5104 4.5005
R22239 DVDD.n5104 DVDD.n449 4.5005
R22240 DVDD.n5141 DVDD.n5136 4.5005
R22241 DVDD.n5141 DVDD.n449 4.5005
R22242 DVDD.n5139 DVDD.n5136 4.5005
R22243 DVDD.n5139 DVDD.n449 4.5005
R22244 DVDD.n5137 DVDD.n5136 4.5005
R22245 DVDD.n5137 DVDD.n449 4.5005
R22246 DVDD.n136 DVDD.n130 4.5005
R22247 DVDD.n5851 DVDD.n136 4.5005
R22248 DVDD.n138 DVDD.n130 4.5005
R22249 DVDD.n5851 DVDD.n138 4.5005
R22250 DVDD.n135 DVDD.n130 4.5005
R22251 DVDD.n5851 DVDD.n135 4.5005
R22252 DVDD.n5850 DVDD.n130 4.5005
R22253 DVDD.n5851 DVDD.n5850 4.5005
R22254 DVDD.n79 DVDD.n74 4.5005
R22255 DVDD.n77 DVDD.n74 4.5005
R22256 DVDD.n76 DVDD.n74 4.5005
R22257 DVDD.n5922 DVDD.n74 4.5005
R22258 DVDD.n5923 DVDD.n76 4.5005
R22259 DVDD.n5923 DVDD.n5922 4.5005
R22260 DVDD.n81 DVDD.n76 4.5005
R22261 DVDD.n5922 DVDD.n81 4.5005
R22262 DVDD.n5921 DVDD.n76 4.5005
R22263 DVDD.n5922 DVDD.n5921 4.5005
R22264 DVDD.n5430 DVDD.n322 4.5005
R22265 DVDD.n5430 DVDD.n324 4.5005
R22266 DVDD.n5430 DVDD.n321 4.5005
R22267 DVDD.n5430 DVDD.n5429 4.5005
R22268 DVDD.n327 DVDD.n322 4.5005
R22269 DVDD.n5428 DVDD.n322 4.5005
R22270 DVDD.n326 DVDD.n322 4.5005
R22271 DVDD.n326 DVDD.n324 4.5005
R22272 DVDD.n5428 DVDD.n324 4.5005
R22273 DVDD.n327 DVDD.n324 4.5005
R22274 DVDD.n5914 DVDD.n114 4.5005
R22275 DVDD.n5914 DVDD.n5910 4.5005
R22276 DVDD.n5914 DVDD.n113 4.5005
R22277 DVDD.n5911 DVDD.n108 4.5005
R22278 DVDD.n5911 DVDD.n107 4.5005
R22279 DVDD.n5914 DVDD.n5911 4.5005
R22280 DVDD.n112 DVDD.n108 4.5005
R22281 DVDD.n112 DVDD.n107 4.5005
R22282 DVDD.n5914 DVDD.n112 4.5005
R22283 DVDD.n5912 DVDD.n108 4.5005
R22284 DVDD.n5912 DVDD.n107 4.5005
R22285 DVDD.n5914 DVDD.n5912 4.5005
R22286 DVDD.n111 DVDD.n108 4.5005
R22287 DVDD.n111 DVDD.n107 4.5005
R22288 DVDD.n5914 DVDD.n111 4.5005
R22289 DVDD.n5914 DVDD.n5913 4.5005
R22290 DVDD.n5914 DVDD.n110 4.5005
R22291 DVDD.n110 DVDD.n107 4.5005
R22292 DVDD.n110 DVDD.n108 4.5005
R22293 DVDD.n5913 DVDD.n107 4.5005
R22294 DVDD.n5913 DVDD.n108 4.5005
R22295 DVDD.n113 DVDD.n107 4.5005
R22296 DVDD.n113 DVDD.n108 4.5005
R22297 DVDD.n5910 DVDD.n107 4.5005
R22298 DVDD.n5910 DVDD.n108 4.5005
R22299 DVDD.n114 DVDD.n107 4.5005
R22300 DVDD.n114 DVDD.n108 4.5005
R22301 DVDD.n5914 DVDD.n102 4.5005
R22302 DVDD.n109 DVDD.n108 4.5005
R22303 DVDD.n109 DVDD.n107 4.5005
R22304 DVDD.n5914 DVDD.n109 4.5005
R22305 DVDD.n5915 DVDD.n108 4.5005
R22306 DVDD.n5915 DVDD.n107 4.5005
R22307 DVDD.n5915 DVDD.n5914 4.5005
R22308 DVDD.n108 DVDD.n102 4.5005
R22309 DVDD.n107 DVDD.n102 4.5005
R22310 DVDD.n5417 DVDD.n5412 4.5005
R22311 DVDD.n5417 DVDD.n5413 4.5005
R22312 DVDD.n5417 DVDD.n5411 4.5005
R22313 DVDD.n5414 DVDD.n325 4.5005
R22314 DVDD.n5414 DVDD.n353 4.5005
R22315 DVDD.n5417 DVDD.n5414 4.5005
R22316 DVDD.n5410 DVDD.n325 4.5005
R22317 DVDD.n5410 DVDD.n353 4.5005
R22318 DVDD.n5417 DVDD.n5410 4.5005
R22319 DVDD.n5415 DVDD.n325 4.5005
R22320 DVDD.n5415 DVDD.n353 4.5005
R22321 DVDD.n5417 DVDD.n5415 4.5005
R22322 DVDD.n5409 DVDD.n325 4.5005
R22323 DVDD.n5409 DVDD.n353 4.5005
R22324 DVDD.n5417 DVDD.n5409 4.5005
R22325 DVDD.n5417 DVDD.n5416 4.5005
R22326 DVDD.n5417 DVDD.n5408 4.5005
R22327 DVDD.n5408 DVDD.n353 4.5005
R22328 DVDD.n5408 DVDD.n325 4.5005
R22329 DVDD.n5416 DVDD.n353 4.5005
R22330 DVDD.n5416 DVDD.n325 4.5005
R22331 DVDD.n5411 DVDD.n353 4.5005
R22332 DVDD.n5411 DVDD.n325 4.5005
R22333 DVDD.n5413 DVDD.n353 4.5005
R22334 DVDD.n5413 DVDD.n325 4.5005
R22335 DVDD.n5412 DVDD.n353 4.5005
R22336 DVDD.n5412 DVDD.n325 4.5005
R22337 DVDD.n5417 DVDD.n349 4.5005
R22338 DVDD.n352 DVDD.n325 4.5005
R22339 DVDD.n353 DVDD.n352 4.5005
R22340 DVDD.n5417 DVDD.n352 4.5005
R22341 DVDD.n5418 DVDD.n325 4.5005
R22342 DVDD.n5418 DVDD.n353 4.5005
R22343 DVDD.n5418 DVDD.n5417 4.5005
R22344 DVDD.n349 DVDD.n325 4.5005
R22345 DVDD.n353 DVDD.n349 4.5005
R22346 DVDD.n285 DVDD.n271 4.5005
R22347 DVDD.n5477 DVDD.n285 4.5005
R22348 DVDD.n283 DVDD.n271 4.5005
R22349 DVDD.n5477 DVDD.n283 4.5005
R22350 DVDD.n286 DVDD.n271 4.5005
R22351 DVDD.n5477 DVDD.n286 4.5005
R22352 DVDD.n282 DVDD.n271 4.5005
R22353 DVDD.n5477 DVDD.n282 4.5005
R22354 DVDD.n287 DVDD.n271 4.5005
R22355 DVDD.n5477 DVDD.n287 4.5005
R22356 DVDD.n281 DVDD.n271 4.5005
R22357 DVDD.n5477 DVDD.n281 4.5005
R22358 DVDD.n288 DVDD.n271 4.5005
R22359 DVDD.n5477 DVDD.n288 4.5005
R22360 DVDD.n280 DVDD.n271 4.5005
R22361 DVDD.n5477 DVDD.n280 4.5005
R22362 DVDD.n289 DVDD.n271 4.5005
R22363 DVDD.n5477 DVDD.n289 4.5005
R22364 DVDD.n279 DVDD.n271 4.5005
R22365 DVDD.n5477 DVDD.n279 4.5005
R22366 DVDD.n290 DVDD.n271 4.5005
R22367 DVDD.n5477 DVDD.n290 4.5005
R22368 DVDD.n278 DVDD.n271 4.5005
R22369 DVDD.n5477 DVDD.n278 4.5005
R22370 DVDD.n291 DVDD.n271 4.5005
R22371 DVDD.n5477 DVDD.n291 4.5005
R22372 DVDD.n277 DVDD.n271 4.5005
R22373 DVDD.n5477 DVDD.n277 4.5005
R22374 DVDD.n292 DVDD.n271 4.5005
R22375 DVDD.n5477 DVDD.n292 4.5005
R22376 DVDD.n276 DVDD.n271 4.5005
R22377 DVDD.n5477 DVDD.n276 4.5005
R22378 DVDD.n293 DVDD.n271 4.5005
R22379 DVDD.n5477 DVDD.n293 4.5005
R22380 DVDD.n275 DVDD.n271 4.5005
R22381 DVDD.n5477 DVDD.n275 4.5005
R22382 DVDD.n5478 DVDD.n271 4.5005
R22383 DVDD.n5478 DVDD.n5477 4.5005
R22384 DVDD.n5565 DVDD.n69 4.5005
R22385 DVDD.n5651 DVDD.n69 4.5005
R22386 DVDD.n5576 DVDD.n5565 4.5005
R22387 DVDD.n5651 DVDD.n5576 4.5005
R22388 DVDD.n5604 DVDD.n5565 4.5005
R22389 DVDD.n5651 DVDD.n5604 4.5005
R22390 DVDD.n5575 DVDD.n5565 4.5005
R22391 DVDD.n5651 DVDD.n5575 4.5005
R22392 DVDD.n5605 DVDD.n5565 4.5005
R22393 DVDD.n5651 DVDD.n5605 4.5005
R22394 DVDD.n5574 DVDD.n5565 4.5005
R22395 DVDD.n5651 DVDD.n5574 4.5005
R22396 DVDD.n5606 DVDD.n5565 4.5005
R22397 DVDD.n5651 DVDD.n5606 4.5005
R22398 DVDD.n5573 DVDD.n5565 4.5005
R22399 DVDD.n5651 DVDD.n5573 4.5005
R22400 DVDD.n5607 DVDD.n5565 4.5005
R22401 DVDD.n5651 DVDD.n5607 4.5005
R22402 DVDD.n5572 DVDD.n5565 4.5005
R22403 DVDD.n5651 DVDD.n5572 4.5005
R22404 DVDD.n5608 DVDD.n5565 4.5005
R22405 DVDD.n5651 DVDD.n5608 4.5005
R22406 DVDD.n5571 DVDD.n5565 4.5005
R22407 DVDD.n5651 DVDD.n5571 4.5005
R22408 DVDD.n5609 DVDD.n5565 4.5005
R22409 DVDD.n5651 DVDD.n5609 4.5005
R22410 DVDD.n5570 DVDD.n5565 4.5005
R22411 DVDD.n5651 DVDD.n5570 4.5005
R22412 DVDD.n5610 DVDD.n5565 4.5005
R22413 DVDD.n5651 DVDD.n5610 4.5005
R22414 DVDD.n5569 DVDD.n5565 4.5005
R22415 DVDD.n5651 DVDD.n5569 4.5005
R22416 DVDD.n5650 DVDD.n5565 4.5005
R22417 DVDD.n5651 DVDD.n5650 4.5005
R22418 DVDD.n5568 DVDD.n5565 4.5005
R22419 DVDD.n5651 DVDD.n5568 4.5005
R22420 DVDD.n5652 DVDD.n5565 4.5005
R22421 DVDD.n5652 DVDD.n5651 4.5005
R22422 DVDD.n4413 DVDD.n1584 4.5005
R22423 DVDD.n4416 DVDD.n1584 4.5005
R22424 DVDD.n4416 DVDD.n1118 4.5005
R22425 DVDD.n4416 DVDD.n1585 4.5005
R22426 DVDD.n4416 DVDD.n1117 4.5005
R22427 DVDD.n4416 DVDD.n1586 4.5005
R22428 DVDD.n4416 DVDD.n1116 4.5005
R22429 DVDD.n4416 DVDD.n1587 4.5005
R22430 DVDD.n4416 DVDD.n1115 4.5005
R22431 DVDD.n4416 DVDD.n1588 4.5005
R22432 DVDD.n4416 DVDD.n1114 4.5005
R22433 DVDD.n4416 DVDD.n1589 4.5005
R22434 DVDD.n4416 DVDD.n1113 4.5005
R22435 DVDD.n4416 DVDD.n1590 4.5005
R22436 DVDD.n4416 DVDD.n1112 4.5005
R22437 DVDD.n4416 DVDD.n1591 4.5005
R22438 DVDD.n4416 DVDD.n1111 4.5005
R22439 DVDD.n4416 DVDD.n1592 4.5005
R22440 DVDD.n4416 DVDD.n1110 4.5005
R22441 DVDD.n4416 DVDD.n1593 4.5005
R22442 DVDD.n4416 DVDD.n1109 4.5005
R22443 DVDD.n4415 DVDD.n4400 4.5005
R22444 DVDD.n4416 DVDD.n4415 4.5005
R22445 DVDD.n4500 DVDD.n1073 4.5005
R22446 DVDD.n4562 DVDD.n4500 4.5005
R22447 DVDD.n4562 DVDD.n1084 4.5005
R22448 DVDD.n1084 DVDD.n1073 4.5005
R22449 DVDD.n4562 DVDD.n4501 4.5005
R22450 DVDD.n4501 DVDD.n1073 4.5005
R22451 DVDD.n1076 DVDD.n1073 4.5005
R22452 DVDD.n4508 DVDD.n1073 4.5005
R22453 DVDD.n1077 DVDD.n1073 4.5005
R22454 DVDD.n4562 DVDD.n1083 4.5005
R22455 DVDD.n1083 DVDD.n1073 4.5005
R22456 DVDD.n4562 DVDD.n4502 4.5005
R22457 DVDD.n4502 DVDD.n1073 4.5005
R22458 DVDD.n4562 DVDD.n1082 4.5005
R22459 DVDD.n1082 DVDD.n1073 4.5005
R22460 DVDD.n4562 DVDD.n4503 4.5005
R22461 DVDD.n4503 DVDD.n1073 4.5005
R22462 DVDD.n4507 DVDD.n1073 4.5005
R22463 DVDD.n1078 DVDD.n1073 4.5005
R22464 DVDD.n4506 DVDD.n1073 4.5005
R22465 DVDD.n4562 DVDD.n1081 4.5005
R22466 DVDD.n1081 DVDD.n1073 4.5005
R22467 DVDD.n4562 DVDD.n4504 4.5005
R22468 DVDD.n4504 DVDD.n1073 4.5005
R22469 DVDD.n4562 DVDD.n1080 4.5005
R22470 DVDD.n1080 DVDD.n1073 4.5005
R22471 DVDD.n4562 DVDD.n4505 4.5005
R22472 DVDD.n4505 DVDD.n1073 4.5005
R22473 DVDD.n1079 DVDD.n1073 4.5005
R22474 DVDD.n4563 DVDD.n1073 4.5005
R22475 DVDD.n1073 DVDD.n1071 4.5005
R22476 DVDD.n4562 DVDD.n1071 4.5005
R22477 DVDD.n4563 DVDD.n4562 4.5005
R22478 DVDD.n4562 DVDD.n1079 4.5005
R22479 DVDD.n4562 DVDD.n4506 4.5005
R22480 DVDD.n4562 DVDD.n1078 4.5005
R22481 DVDD.n4562 DVDD.n4507 4.5005
R22482 DVDD.n4562 DVDD.n1077 4.5005
R22483 DVDD.n4562 DVDD.n4508 4.5005
R22484 DVDD.n4562 DVDD.n1076 4.5005
R22485 DVDD.n4562 DVDD.n4561 4.5005
R22486 DVDD.n4561 DVDD.n1073 4.5005
R22487 DVDD.n756 DVDD.n695 4.5005
R22488 DVDD.n756 DVDD.n702 4.5005
R22489 DVDD.n771 DVDD.n702 4.5005
R22490 DVDD.n771 DVDD.n695 4.5005
R22491 DVDD.n755 DVDD.n702 4.5005
R22492 DVDD.n755 DVDD.n695 4.5005
R22493 DVDD.n777 DVDD.n695 4.5005
R22494 DVDD.n779 DVDD.n695 4.5005
R22495 DVDD.n751 DVDD.n695 4.5005
R22496 DVDD.n784 DVDD.n702 4.5005
R22497 DVDD.n784 DVDD.n695 4.5005
R22498 DVDD.n786 DVDD.n702 4.5005
R22499 DVDD.n786 DVDD.n695 4.5005
R22500 DVDD.n749 DVDD.n702 4.5005
R22501 DVDD.n749 DVDD.n695 4.5005
R22502 DVDD.n791 DVDD.n702 4.5005
R22503 DVDD.n791 DVDD.n695 4.5005
R22504 DVDD.n747 DVDD.n695 4.5005
R22505 DVDD.n797 DVDD.n695 4.5005
R22506 DVDD.n799 DVDD.n695 4.5005
R22507 DVDD.n745 DVDD.n702 4.5005
R22508 DVDD.n745 DVDD.n695 4.5005
R22509 DVDD.n804 DVDD.n702 4.5005
R22510 DVDD.n804 DVDD.n695 4.5005
R22511 DVDD.n806 DVDD.n702 4.5005
R22512 DVDD.n806 DVDD.n695 4.5005
R22513 DVDD.n744 DVDD.n702 4.5005
R22514 DVDD.n744 DVDD.n695 4.5005
R22515 DVDD.n812 DVDD.n695 4.5005
R22516 DVDD.n814 DVDD.n695 4.5005
R22517 DVDD.n740 DVDD.n695 4.5005
R22518 DVDD.n740 DVDD.n702 4.5005
R22519 DVDD.n814 DVDD.n702 4.5005
R22520 DVDD.n812 DVDD.n702 4.5005
R22521 DVDD.n799 DVDD.n702 4.5005
R22522 DVDD.n797 DVDD.n702 4.5005
R22523 DVDD.n747 DVDD.n702 4.5005
R22524 DVDD.n751 DVDD.n702 4.5005
R22525 DVDD.n779 DVDD.n702 4.5005
R22526 DVDD.n777 DVDD.n702 4.5005
R22527 DVDD.n769 DVDD.n702 4.5005
R22528 DVDD.n769 DVDD.n695 4.5005
R22529 DVDD.n4941 DVDD.n672 4.5005
R22530 DVDD.n5006 DVDD.n4941 4.5005
R22531 DVDD.n5006 DVDD.n683 4.5005
R22532 DVDD.n683 DVDD.n672 4.5005
R22533 DVDD.n5006 DVDD.n4942 4.5005
R22534 DVDD.n4942 DVDD.n672 4.5005
R22535 DVDD.n675 DVDD.n672 4.5005
R22536 DVDD.n4950 DVDD.n672 4.5005
R22537 DVDD.n676 DVDD.n672 4.5005
R22538 DVDD.n5006 DVDD.n682 4.5005
R22539 DVDD.n682 DVDD.n672 4.5005
R22540 DVDD.n5006 DVDD.n4943 4.5005
R22541 DVDD.n4943 DVDD.n672 4.5005
R22542 DVDD.n5006 DVDD.n681 4.5005
R22543 DVDD.n681 DVDD.n672 4.5005
R22544 DVDD.n5006 DVDD.n4944 4.5005
R22545 DVDD.n4944 DVDD.n672 4.5005
R22546 DVDD.n4949 DVDD.n672 4.5005
R22547 DVDD.n677 DVDD.n672 4.5005
R22548 DVDD.n4948 DVDD.n672 4.5005
R22549 DVDD.n5006 DVDD.n680 4.5005
R22550 DVDD.n680 DVDD.n672 4.5005
R22551 DVDD.n5006 DVDD.n4945 4.5005
R22552 DVDD.n4945 DVDD.n672 4.5005
R22553 DVDD.n5006 DVDD.n679 4.5005
R22554 DVDD.n679 DVDD.n672 4.5005
R22555 DVDD.n5006 DVDD.n4946 4.5005
R22556 DVDD.n4946 DVDD.n672 4.5005
R22557 DVDD.n678 DVDD.n672 4.5005
R22558 DVDD.n4947 DVDD.n672 4.5005
R22559 DVDD.n5007 DVDD.n672 4.5005
R22560 DVDD.n5007 DVDD.n5006 4.5005
R22561 DVDD.n5006 DVDD.n4947 4.5005
R22562 DVDD.n5006 DVDD.n678 4.5005
R22563 DVDD.n5006 DVDD.n4948 4.5005
R22564 DVDD.n5006 DVDD.n677 4.5005
R22565 DVDD.n5006 DVDD.n4949 4.5005
R22566 DVDD.n5006 DVDD.n676 4.5005
R22567 DVDD.n5006 DVDD.n4950 4.5005
R22568 DVDD.n5006 DVDD.n675 4.5005
R22569 DVDD.n5006 DVDD.n5005 4.5005
R22570 DVDD.n5005 DVDD.n672 4.5005
R22571 DVDD.n5318 DVDD.n463 4.5005
R22572 DVDD.n5320 DVDD.n463 4.5005
R22573 DVDD.n5320 DVDD.n461 4.5005
R22574 DVDD.n5318 DVDD.n461 4.5005
R22575 DVDD.n5320 DVDD.n464 4.5005
R22576 DVDD.n5318 DVDD.n464 4.5005
R22577 DVDD.n5318 DVDD.n452 4.5005
R22578 DVDD.n5318 DVDD.n472 4.5005
R22579 DVDD.n5318 DVDD.n453 4.5005
R22580 DVDD.n5320 DVDD.n460 4.5005
R22581 DVDD.n5318 DVDD.n460 4.5005
R22582 DVDD.n5320 DVDD.n465 4.5005
R22583 DVDD.n5318 DVDD.n465 4.5005
R22584 DVDD.n5320 DVDD.n459 4.5005
R22585 DVDD.n5318 DVDD.n459 4.5005
R22586 DVDD.n5320 DVDD.n466 4.5005
R22587 DVDD.n5318 DVDD.n466 4.5005
R22588 DVDD.n5318 DVDD.n471 4.5005
R22589 DVDD.n5318 DVDD.n454 4.5005
R22590 DVDD.n5318 DVDD.n470 4.5005
R22591 DVDD.n5320 DVDD.n458 4.5005
R22592 DVDD.n5318 DVDD.n458 4.5005
R22593 DVDD.n5320 DVDD.n467 4.5005
R22594 DVDD.n5318 DVDD.n467 4.5005
R22595 DVDD.n5320 DVDD.n457 4.5005
R22596 DVDD.n5318 DVDD.n457 4.5005
R22597 DVDD.n5320 DVDD.n468 4.5005
R22598 DVDD.n5318 DVDD.n468 4.5005
R22599 DVDD.n5318 DVDD.n455 4.5005
R22600 DVDD.n5318 DVDD.n469 4.5005
R22601 DVDD.n5318 DVDD.n456 4.5005
R22602 DVDD.n5320 DVDD.n456 4.5005
R22603 DVDD.n5320 DVDD.n469 4.5005
R22604 DVDD.n5320 DVDD.n455 4.5005
R22605 DVDD.n5320 DVDD.n470 4.5005
R22606 DVDD.n5320 DVDD.n454 4.5005
R22607 DVDD.n5320 DVDD.n471 4.5005
R22608 DVDD.n5320 DVDD.n453 4.5005
R22609 DVDD.n5320 DVDD.n472 4.5005
R22610 DVDD.n5320 DVDD.n452 4.5005
R22611 DVDD.n5320 DVDD.n5319 4.5005
R22612 DVDD.n5319 DVDD.n5318 4.5005
R22613 DVDD.n5836 DVDD.n140 4.5005
R22614 DVDD.n143 DVDD.n140 4.5005
R22615 DVDD.n154 DVDD.n143 4.5005
R22616 DVDD.n5836 DVDD.n154 4.5005
R22617 DVDD.n156 DVDD.n143 4.5005
R22618 DVDD.n5836 DVDD.n156 4.5005
R22619 DVDD.n5836 DVDD.n153 4.5005
R22620 DVDD.n5836 DVDD.n157 4.5005
R22621 DVDD.n5836 DVDD.n152 4.5005
R22622 DVDD.n158 DVDD.n143 4.5005
R22623 DVDD.n5836 DVDD.n158 4.5005
R22624 DVDD.n151 DVDD.n143 4.5005
R22625 DVDD.n5836 DVDD.n151 4.5005
R22626 DVDD.n159 DVDD.n143 4.5005
R22627 DVDD.n5836 DVDD.n159 4.5005
R22628 DVDD.n150 DVDD.n143 4.5005
R22629 DVDD.n5836 DVDD.n150 4.5005
R22630 DVDD.n5836 DVDD.n160 4.5005
R22631 DVDD.n5836 DVDD.n149 4.5005
R22632 DVDD.n5836 DVDD.n161 4.5005
R22633 DVDD.n148 DVDD.n143 4.5005
R22634 DVDD.n5836 DVDD.n148 4.5005
R22635 DVDD.n162 DVDD.n143 4.5005
R22636 DVDD.n5836 DVDD.n162 4.5005
R22637 DVDD.n147 DVDD.n143 4.5005
R22638 DVDD.n5836 DVDD.n147 4.5005
R22639 DVDD.n163 DVDD.n143 4.5005
R22640 DVDD.n5836 DVDD.n163 4.5005
R22641 DVDD.n5836 DVDD.n146 4.5005
R22642 DVDD.n5836 DVDD.n5835 4.5005
R22643 DVDD.n5836 DVDD.n145 4.5005
R22644 DVDD.n145 DVDD.n143 4.5005
R22645 DVDD.n5835 DVDD.n143 4.5005
R22646 DVDD.n146 DVDD.n143 4.5005
R22647 DVDD.n161 DVDD.n143 4.5005
R22648 DVDD.n149 DVDD.n143 4.5005
R22649 DVDD.n160 DVDD.n143 4.5005
R22650 DVDD.n152 DVDD.n143 4.5005
R22651 DVDD.n157 DVDD.n143 4.5005
R22652 DVDD.n153 DVDD.n143 4.5005
R22653 DVDD.n5837 DVDD.n143 4.5005
R22654 DVDD.n5837 DVDD.n5836 4.5005
R22655 DVDD.n59 DVDD.n43 4.5005
R22656 DVDD.n5934 DVDD.n59 4.5005
R22657 DVDD.n57 DVDD.n43 4.5005
R22658 DVDD.n5934 DVDD.n57 4.5005
R22659 DVDD.n5934 DVDD.n60 4.5005
R22660 DVDD.n5934 DVDD.n56 4.5005
R22661 DVDD.n5934 DVDD.n61 4.5005
R22662 DVDD.n55 DVDD.n43 4.5005
R22663 DVDD.n5934 DVDD.n55 4.5005
R22664 DVDD.n62 DVDD.n43 4.5005
R22665 DVDD.n5934 DVDD.n62 4.5005
R22666 DVDD.n54 DVDD.n43 4.5005
R22667 DVDD.n5934 DVDD.n54 4.5005
R22668 DVDD.n63 DVDD.n43 4.5005
R22669 DVDD.n5934 DVDD.n63 4.5005
R22670 DVDD.n5934 DVDD.n53 4.5005
R22671 DVDD.n5934 DVDD.n64 4.5005
R22672 DVDD.n5934 DVDD.n52 4.5005
R22673 DVDD.n65 DVDD.n43 4.5005
R22674 DVDD.n5934 DVDD.n65 4.5005
R22675 DVDD.n51 DVDD.n43 4.5005
R22676 DVDD.n5934 DVDD.n51 4.5005
R22677 DVDD.n66 DVDD.n43 4.5005
R22678 DVDD.n5934 DVDD.n66 4.5005
R22679 DVDD.n50 DVDD.n43 4.5005
R22680 DVDD.n5934 DVDD.n50 4.5005
R22681 DVDD.n5934 DVDD.n67 4.5005
R22682 DVDD.n5934 DVDD.n49 4.5005
R22683 DVDD.n5934 DVDD.n68 4.5005
R22684 DVDD.n5565 DVDD.n5563 4.5005
R22685 DVDD.n5651 DVDD.n5563 4.5005
R22686 DVDD.n68 DVDD.n43 4.5005
R22687 DVDD.n5651 DVDD.n70 4.5005
R22688 DVDD.n5565 DVDD.n70 4.5005
R22689 DVDD.n5934 DVDD.n48 4.5005
R22690 DVDD.n48 DVDD.n43 4.5005
R22691 DVDD.n49 DVDD.n43 4.5005
R22692 DVDD.n67 DVDD.n43 4.5005
R22693 DVDD.n52 DVDD.n43 4.5005
R22694 DVDD.n64 DVDD.n43 4.5005
R22695 DVDD.n53 DVDD.n43 4.5005
R22696 DVDD.n61 DVDD.n43 4.5005
R22697 DVDD.n56 DVDD.n43 4.5005
R22698 DVDD.n60 DVDD.n43 4.5005
R22699 DVDD.n5933 DVDD.n43 4.5005
R22700 DVDD.n5934 DVDD.n5933 4.5005
R22701 DVDD.n5477 DVDD.n268 4.5005
R22702 DVDD.n271 DVDD.n268 4.5005
R22703 DVDD.n295 DVDD.n270 4.5005
R22704 DVDD.n308 DVDD.n295 4.5005
R22705 DVDD.n5474 DVDD.n308 4.5005
R22706 DVDD.n306 DVDD.n295 4.5005
R22707 DVDD.n5474 DVDD.n306 4.5005
R22708 DVDD.n309 DVDD.n295 4.5005
R22709 DVDD.n5474 DVDD.n309 4.5005
R22710 DVDD.n5474 DVDD.n305 4.5005
R22711 DVDD.n5474 DVDD.n310 4.5005
R22712 DVDD.n5474 DVDD.n304 4.5005
R22713 DVDD.n311 DVDD.n295 4.5005
R22714 DVDD.n5474 DVDD.n311 4.5005
R22715 DVDD.n303 DVDD.n295 4.5005
R22716 DVDD.n5474 DVDD.n303 4.5005
R22717 DVDD.n312 DVDD.n295 4.5005
R22718 DVDD.n5474 DVDD.n312 4.5005
R22719 DVDD.n302 DVDD.n295 4.5005
R22720 DVDD.n5474 DVDD.n302 4.5005
R22721 DVDD.n5474 DVDD.n313 4.5005
R22722 DVDD.n5474 DVDD.n301 4.5005
R22723 DVDD.n5474 DVDD.n314 4.5005
R22724 DVDD.n300 DVDD.n295 4.5005
R22725 DVDD.n5474 DVDD.n300 4.5005
R22726 DVDD.n315 DVDD.n295 4.5005
R22727 DVDD.n5474 DVDD.n315 4.5005
R22728 DVDD.n299 DVDD.n295 4.5005
R22729 DVDD.n5474 DVDD.n299 4.5005
R22730 DVDD.n5473 DVDD.n295 4.5005
R22731 DVDD.n5474 DVDD.n5473 4.5005
R22732 DVDD.n5474 DVDD.n298 4.5005
R22733 DVDD.n5474 DVDD.n272 4.5005
R22734 DVDD.n5474 DVDD.n270 4.5005
R22735 DVDD.n295 DVDD.n272 4.5005
R22736 DVDD.n298 DVDD.n295 4.5005
R22737 DVDD.n314 DVDD.n295 4.5005
R22738 DVDD.n301 DVDD.n295 4.5005
R22739 DVDD.n313 DVDD.n295 4.5005
R22740 DVDD.n304 DVDD.n295 4.5005
R22741 DVDD.n310 DVDD.n295 4.5005
R22742 DVDD.n305 DVDD.n295 4.5005
R22743 DVDD.n5477 DVDD.n5476 4.5005
R22744 DVDD.n5476 DVDD.n271 4.5005
R22745 DVDD.n5475 DVDD.n295 4.5005
R22746 DVDD.n5475 DVDD.n5474 4.5005
R22747 DVDD.n4700 DVDD.n4647 4.5005
R22748 DVDD.n4647 DVDD.n971 4.5005
R22749 DVDD.n4700 DVDD.n984 4.5005
R22750 DVDD.n984 DVDD.n971 4.5005
R22751 DVDD.n4700 DVDD.n4648 4.5005
R22752 DVDD.n4648 DVDD.n971 4.5005
R22753 DVDD.n4700 DVDD.n983 4.5005
R22754 DVDD.n983 DVDD.n971 4.5005
R22755 DVDD.n4700 DVDD.n4649 4.5005
R22756 DVDD.n4649 DVDD.n971 4.5005
R22757 DVDD.n4700 DVDD.n982 4.5005
R22758 DVDD.n982 DVDD.n971 4.5005
R22759 DVDD.n4700 DVDD.n4650 4.5005
R22760 DVDD.n4650 DVDD.n971 4.5005
R22761 DVDD.n4700 DVDD.n981 4.5005
R22762 DVDD.n981 DVDD.n971 4.5005
R22763 DVDD.n4700 DVDD.n4651 4.5005
R22764 DVDD.n4651 DVDD.n971 4.5005
R22765 DVDD.n4700 DVDD.n980 4.5005
R22766 DVDD.n980 DVDD.n971 4.5005
R22767 DVDD.n4700 DVDD.n4652 4.5005
R22768 DVDD.n4652 DVDD.n971 4.5005
R22769 DVDD.n4700 DVDD.n979 4.5005
R22770 DVDD.n979 DVDD.n971 4.5005
R22771 DVDD.n4700 DVDD.n4653 4.5005
R22772 DVDD.n4653 DVDD.n971 4.5005
R22773 DVDD.n4700 DVDD.n978 4.5005
R22774 DVDD.n978 DVDD.n971 4.5005
R22775 DVDD.n4700 DVDD.n4654 4.5005
R22776 DVDD.n4654 DVDD.n971 4.5005
R22777 DVDD.n4700 DVDD.n977 4.5005
R22778 DVDD.n977 DVDD.n971 4.5005
R22779 DVDD.n4700 DVDD.n4655 4.5005
R22780 DVDD.n4655 DVDD.n971 4.5005
R22781 DVDD.n4700 DVDD.n976 4.5005
R22782 DVDD.n976 DVDD.n971 4.5005
R22783 DVDD.n4700 DVDD.n4699 4.5005
R22784 DVDD.n4699 DVDD.n971 4.5005
R22785 DVDD.n31 DVDD.n18 4.5005
R22786 DVDD.n5956 DVDD.n18 4.5005
R22787 DVDD.n31 DVDD.n17 4.5005
R22788 DVDD.n5956 DVDD.n17 4.5005
R22789 DVDD.n31 DVDD.n19 4.5005
R22790 DVDD.n5956 DVDD.n19 4.5005
R22791 DVDD.n31 DVDD.n16 4.5005
R22792 DVDD.n5956 DVDD.n16 4.5005
R22793 DVDD.n31 DVDD.n20 4.5005
R22794 DVDD.n5956 DVDD.n20 4.5005
R22795 DVDD.n31 DVDD.n15 4.5005
R22796 DVDD.n5956 DVDD.n15 4.5005
R22797 DVDD.n31 DVDD.n21 4.5005
R22798 DVDD.n5956 DVDD.n21 4.5005
R22799 DVDD.n31 DVDD.n14 4.5005
R22800 DVDD.n5956 DVDD.n14 4.5005
R22801 DVDD.n31 DVDD.n22 4.5005
R22802 DVDD.n5956 DVDD.n22 4.5005
R22803 DVDD.n31 DVDD.n13 4.5005
R22804 DVDD.n5956 DVDD.n13 4.5005
R22805 DVDD.n31 DVDD.n23 4.5005
R22806 DVDD.n5956 DVDD.n23 4.5005
R22807 DVDD.n31 DVDD.n12 4.5005
R22808 DVDD.n5956 DVDD.n12 4.5005
R22809 DVDD.n31 DVDD.n24 4.5005
R22810 DVDD.n5956 DVDD.n24 4.5005
R22811 DVDD.n31 DVDD.n11 4.5005
R22812 DVDD.n5956 DVDD.n11 4.5005
R22813 DVDD.n31 DVDD.n25 4.5005
R22814 DVDD.n5956 DVDD.n25 4.5005
R22815 DVDD.n31 DVDD.n10 4.5005
R22816 DVDD.n5956 DVDD.n10 4.5005
R22817 DVDD.n31 DVDD.n26 4.5005
R22818 DVDD.n5956 DVDD.n26 4.5005
R22819 DVDD.n31 DVDD.n9 4.5005
R22820 DVDD.n5956 DVDD.n9 4.5005
R22821 DVDD.n31 DVDD.n27 4.5005
R22822 DVDD.n5956 DVDD.n27 4.5005
R22823 DVDD.n4389 DVDD.n1595 4.5005
R22824 DVDD.n4389 DVDD.n4388 4.5005
R22825 DVDD.n4388 DVDD.n1606 4.5005
R22826 DVDD.n4388 DVDD.n1609 4.5005
R22827 DVDD.n4388 DVDD.n1605 4.5005
R22828 DVDD.n4388 DVDD.n1611 4.5005
R22829 DVDD.n4388 DVDD.n1604 4.5005
R22830 DVDD.n4388 DVDD.n1613 4.5005
R22831 DVDD.n4388 DVDD.n1603 4.5005
R22832 DVDD.n4388 DVDD.n1615 4.5005
R22833 DVDD.n4388 DVDD.n1602 4.5005
R22834 DVDD.n4388 DVDD.n1617 4.5005
R22835 DVDD.n4388 DVDD.n1601 4.5005
R22836 DVDD.n4388 DVDD.n1619 4.5005
R22837 DVDD.n4388 DVDD.n1600 4.5005
R22838 DVDD.n4388 DVDD.n1621 4.5005
R22839 DVDD.n4388 DVDD.n1599 4.5005
R22840 DVDD.n4388 DVDD.n1623 4.5005
R22841 DVDD.n4388 DVDD.n1598 4.5005
R22842 DVDD.n4388 DVDD.n1625 4.5005
R22843 DVDD.n4388 DVDD.n1597 4.5005
R22844 DVDD.n4387 DVDD.n4385 4.5005
R22845 DVDD.n4388 DVDD.n4387 4.5005
R22846 DVDD.n4617 DVDD.n1047 4.5005
R22847 DVDD.n4617 DVDD.n1019 4.5005
R22848 DVDD.n1048 DVDD.n1005 4.5005
R22849 DVDD.n4617 DVDD.n1048 4.5005
R22850 DVDD.n1018 DVDD.n1005 4.5005
R22851 DVDD.n4617 DVDD.n1018 4.5005
R22852 DVDD.n1049 DVDD.n1005 4.5005
R22853 DVDD.n4617 DVDD.n1049 4.5005
R22854 DVDD.n1017 DVDD.n1005 4.5005
R22855 DVDD.n4617 DVDD.n1017 4.5005
R22856 DVDD.n4617 DVDD.n1050 4.5005
R22857 DVDD.n4617 DVDD.n1016 4.5005
R22858 DVDD.n4617 DVDD.n1051 4.5005
R22859 DVDD.n1015 DVDD.n1005 4.5005
R22860 DVDD.n4617 DVDD.n1015 4.5005
R22861 DVDD.n1052 DVDD.n1005 4.5005
R22862 DVDD.n4617 DVDD.n1052 4.5005
R22863 DVDD.n1014 DVDD.n1005 4.5005
R22864 DVDD.n4617 DVDD.n1014 4.5005
R22865 DVDD.n1053 DVDD.n1005 4.5005
R22866 DVDD.n4617 DVDD.n1053 4.5005
R22867 DVDD.n4617 DVDD.n1013 4.5005
R22868 DVDD.n4617 DVDD.n1054 4.5005
R22869 DVDD.n4617 DVDD.n1012 4.5005
R22870 DVDD.n1055 DVDD.n1005 4.5005
R22871 DVDD.n4617 DVDD.n1055 4.5005
R22872 DVDD.n1011 DVDD.n1005 4.5005
R22873 DVDD.n4617 DVDD.n1011 4.5005
R22874 DVDD.n1056 DVDD.n1005 4.5005
R22875 DVDD.n4617 DVDD.n1056 4.5005
R22876 DVDD.n1010 DVDD.n1005 4.5005
R22877 DVDD.n4617 DVDD.n1010 4.5005
R22878 DVDD.n4617 DVDD.n4616 4.5005
R22879 DVDD.n4616 DVDD.n1005 4.5005
R22880 DVDD.n1012 DVDD.n1005 4.5005
R22881 DVDD.n1054 DVDD.n1005 4.5005
R22882 DVDD.n1013 DVDD.n1005 4.5005
R22883 DVDD.n1051 DVDD.n1005 4.5005
R22884 DVDD.n1016 DVDD.n1005 4.5005
R22885 DVDD.n1050 DVDD.n1005 4.5005
R22886 DVDD.n1019 DVDD.n1005 4.5005
R22887 DVDD.n1047 DVDD.n1005 4.5005
R22888 DVDD.n4879 DVDD.n716 4.5005
R22889 DVDD.n4879 DVDD.n714 4.5005
R22890 DVDD.n4877 DVDD.n717 4.5005
R22891 DVDD.n4879 DVDD.n717 4.5005
R22892 DVDD.n4877 DVDD.n713 4.5005
R22893 DVDD.n4879 DVDD.n713 4.5005
R22894 DVDD.n4877 DVDD.n718 4.5005
R22895 DVDD.n4879 DVDD.n718 4.5005
R22896 DVDD.n4877 DVDD.n712 4.5005
R22897 DVDD.n4879 DVDD.n712 4.5005
R22898 DVDD.n4879 DVDD.n719 4.5005
R22899 DVDD.n4879 DVDD.n711 4.5005
R22900 DVDD.n4879 DVDD.n720 4.5005
R22901 DVDD.n4877 DVDD.n710 4.5005
R22902 DVDD.n4879 DVDD.n710 4.5005
R22903 DVDD.n4877 DVDD.n721 4.5005
R22904 DVDD.n4879 DVDD.n721 4.5005
R22905 DVDD.n4877 DVDD.n709 4.5005
R22906 DVDD.n4879 DVDD.n709 4.5005
R22907 DVDD.n4877 DVDD.n722 4.5005
R22908 DVDD.n4879 DVDD.n722 4.5005
R22909 DVDD.n4879 DVDD.n708 4.5005
R22910 DVDD.n4879 DVDD.n723 4.5005
R22911 DVDD.n4879 DVDD.n707 4.5005
R22912 DVDD.n4877 DVDD.n724 4.5005
R22913 DVDD.n4879 DVDD.n724 4.5005
R22914 DVDD.n4877 DVDD.n706 4.5005
R22915 DVDD.n4879 DVDD.n706 4.5005
R22916 DVDD.n4877 DVDD.n725 4.5005
R22917 DVDD.n4879 DVDD.n725 4.5005
R22918 DVDD.n4877 DVDD.n705 4.5005
R22919 DVDD.n4879 DVDD.n705 4.5005
R22920 DVDD.n4879 DVDD.n4878 4.5005
R22921 DVDD.n4878 DVDD.n4877 4.5005
R22922 DVDD.n4877 DVDD.n707 4.5005
R22923 DVDD.n4877 DVDD.n723 4.5005
R22924 DVDD.n4877 DVDD.n708 4.5005
R22925 DVDD.n4877 DVDD.n720 4.5005
R22926 DVDD.n4877 DVDD.n711 4.5005
R22927 DVDD.n4877 DVDD.n719 4.5005
R22928 DVDD.n4877 DVDD.n714 4.5005
R22929 DVDD.n4877 DVDD.n716 4.5005
R22930 DVDD.n5013 DVDD.n603 4.5005
R22931 DVDD.n606 DVDD.n603 4.5005
R22932 DVDD.n5014 DVDD.n617 4.5005
R22933 DVDD.n617 DVDD.n603 4.5005
R22934 DVDD.n5014 DVDD.n615 4.5005
R22935 DVDD.n615 DVDD.n603 4.5005
R22936 DVDD.n5014 DVDD.n618 4.5005
R22937 DVDD.n618 DVDD.n603 4.5005
R22938 DVDD.n5014 DVDD.n614 4.5005
R22939 DVDD.n614 DVDD.n603 4.5005
R22940 DVDD.n625 DVDD.n603 4.5005
R22941 DVDD.n607 DVDD.n603 4.5005
R22942 DVDD.n624 DVDD.n603 4.5005
R22943 DVDD.n5014 DVDD.n619 4.5005
R22944 DVDD.n619 DVDD.n603 4.5005
R22945 DVDD.n5014 DVDD.n613 4.5005
R22946 DVDD.n613 DVDD.n603 4.5005
R22947 DVDD.n5014 DVDD.n620 4.5005
R22948 DVDD.n620 DVDD.n603 4.5005
R22949 DVDD.n5014 DVDD.n612 4.5005
R22950 DVDD.n612 DVDD.n603 4.5005
R22951 DVDD.n608 DVDD.n603 4.5005
R22952 DVDD.n623 DVDD.n603 4.5005
R22953 DVDD.n609 DVDD.n603 4.5005
R22954 DVDD.n5014 DVDD.n621 4.5005
R22955 DVDD.n621 DVDD.n603 4.5005
R22956 DVDD.n5014 DVDD.n611 4.5005
R22957 DVDD.n611 DVDD.n603 4.5005
R22958 DVDD.n5014 DVDD.n622 4.5005
R22959 DVDD.n622 DVDD.n603 4.5005
R22960 DVDD.n5014 DVDD.n610 4.5005
R22961 DVDD.n610 DVDD.n603 4.5005
R22962 DVDD.n5015 DVDD.n603 4.5005
R22963 DVDD.n5015 DVDD.n5014 4.5005
R22964 DVDD.n5014 DVDD.n609 4.5005
R22965 DVDD.n5014 DVDD.n623 4.5005
R22966 DVDD.n5014 DVDD.n608 4.5005
R22967 DVDD.n5014 DVDD.n624 4.5005
R22968 DVDD.n5014 DVDD.n607 4.5005
R22969 DVDD.n5014 DVDD.n625 4.5005
R22970 DVDD.n5014 DVDD.n606 4.5005
R22971 DVDD.n5014 DVDD.n5013 4.5005
R22972 DVDD.n5244 DVDD.n556 4.5005
R22973 DVDD.n5244 DVDD.n495 4.5005
R22974 DVDD.n557 DVDD.n485 4.5005
R22975 DVDD.n5244 DVDD.n557 4.5005
R22976 DVDD.n494 DVDD.n485 4.5005
R22977 DVDD.n5244 DVDD.n494 4.5005
R22978 DVDD.n558 DVDD.n485 4.5005
R22979 DVDD.n5244 DVDD.n558 4.5005
R22980 DVDD.n493 DVDD.n485 4.5005
R22981 DVDD.n5244 DVDD.n493 4.5005
R22982 DVDD.n5244 DVDD.n559 4.5005
R22983 DVDD.n5244 DVDD.n492 4.5005
R22984 DVDD.n5244 DVDD.n560 4.5005
R22985 DVDD.n491 DVDD.n485 4.5005
R22986 DVDD.n5244 DVDD.n491 4.5005
R22987 DVDD.n561 DVDD.n485 4.5005
R22988 DVDD.n5244 DVDD.n561 4.5005
R22989 DVDD.n490 DVDD.n485 4.5005
R22990 DVDD.n5244 DVDD.n490 4.5005
R22991 DVDD.n562 DVDD.n485 4.5005
R22992 DVDD.n5244 DVDD.n562 4.5005
R22993 DVDD.n5244 DVDD.n489 4.5005
R22994 DVDD.n5244 DVDD.n563 4.5005
R22995 DVDD.n5244 DVDD.n488 4.5005
R22996 DVDD.n564 DVDD.n485 4.5005
R22997 DVDD.n5244 DVDD.n564 4.5005
R22998 DVDD.n487 DVDD.n485 4.5005
R22999 DVDD.n5244 DVDD.n487 4.5005
R23000 DVDD.n565 DVDD.n485 4.5005
R23001 DVDD.n5244 DVDD.n565 4.5005
R23002 DVDD.n486 DVDD.n485 4.5005
R23003 DVDD.n5244 DVDD.n486 4.5005
R23004 DVDD.n5244 DVDD.n5243 4.5005
R23005 DVDD.n5243 DVDD.n485 4.5005
R23006 DVDD.n488 DVDD.n485 4.5005
R23007 DVDD.n563 DVDD.n485 4.5005
R23008 DVDD.n489 DVDD.n485 4.5005
R23009 DVDD.n560 DVDD.n485 4.5005
R23010 DVDD.n492 DVDD.n485 4.5005
R23011 DVDD.n559 DVDD.n485 4.5005
R23012 DVDD.n495 DVDD.n485 4.5005
R23013 DVDD.n556 DVDD.n485 4.5005
R23014 DVDD.n169 DVDD.n166 4.5005
R23015 DVDD.n5786 DVDD.n169 4.5005
R23016 DVDD.n5785 DVDD.n181 4.5005
R23017 DVDD.n181 DVDD.n169 4.5005
R23018 DVDD.n5785 DVDD.n179 4.5005
R23019 DVDD.n179 DVDD.n169 4.5005
R23020 DVDD.n5785 DVDD.n182 4.5005
R23021 DVDD.n182 DVDD.n169 4.5005
R23022 DVDD.n5785 DVDD.n178 4.5005
R23023 DVDD.n178 DVDD.n169 4.5005
R23024 DVDD.n5784 DVDD.n169 4.5005
R23025 DVDD.n171 DVDD.n169 4.5005
R23026 DVDD.n189 DVDD.n169 4.5005
R23027 DVDD.n5785 DVDD.n183 4.5005
R23028 DVDD.n183 DVDD.n169 4.5005
R23029 DVDD.n5785 DVDD.n177 4.5005
R23030 DVDD.n177 DVDD.n169 4.5005
R23031 DVDD.n5785 DVDD.n184 4.5005
R23032 DVDD.n184 DVDD.n169 4.5005
R23033 DVDD.n5785 DVDD.n176 4.5005
R23034 DVDD.n176 DVDD.n169 4.5005
R23035 DVDD.n172 DVDD.n169 4.5005
R23036 DVDD.n188 DVDD.n169 4.5005
R23037 DVDD.n173 DVDD.n169 4.5005
R23038 DVDD.n5785 DVDD.n185 4.5005
R23039 DVDD.n185 DVDD.n169 4.5005
R23040 DVDD.n5785 DVDD.n175 4.5005
R23041 DVDD.n175 DVDD.n169 4.5005
R23042 DVDD.n5785 DVDD.n186 4.5005
R23043 DVDD.n186 DVDD.n169 4.5005
R23044 DVDD.n5785 DVDD.n174 4.5005
R23045 DVDD.n174 DVDD.n169 4.5005
R23046 DVDD.n187 DVDD.n169 4.5005
R23047 DVDD.n5785 DVDD.n187 4.5005
R23048 DVDD.n5785 DVDD.n173 4.5005
R23049 DVDD.n5785 DVDD.n188 4.5005
R23050 DVDD.n5785 DVDD.n172 4.5005
R23051 DVDD.n5785 DVDD.n189 4.5005
R23052 DVDD.n5785 DVDD.n171 4.5005
R23053 DVDD.n5785 DVDD.n5784 4.5005
R23054 DVDD.n5786 DVDD.n5785 4.5005
R23055 DVDD.n5785 DVDD.n166 4.5005
R23056 DVDD.n29 DVDD.n8 4.5005
R23057 DVDD.n31 DVDD.n8 4.5005
R23058 DVDD.n5956 DVDD.n8 4.5005
R23059 DVDD.n5955 DVDD.n29 4.5005
R23060 DVDD.n5955 DVDD.n31 4.5005
R23061 DVDD.n5956 DVDD.n5955 4.5005
R23062 DVDD.n5955 DVDD.n5954 4.5005
R23063 DVDD.n5954 DVDD.n27 4.5005
R23064 DVDD.n29 DVDD.n27 4.5005
R23065 DVDD.n5954 DVDD.n9 4.5005
R23066 DVDD.n29 DVDD.n9 4.5005
R23067 DVDD.n5954 DVDD.n26 4.5005
R23068 DVDD.n29 DVDD.n26 4.5005
R23069 DVDD.n29 DVDD.n10 4.5005
R23070 DVDD.n5954 DVDD.n10 4.5005
R23071 DVDD.n29 DVDD.n25 4.5005
R23072 DVDD.n5954 DVDD.n25 4.5005
R23073 DVDD.n29 DVDD.n11 4.5005
R23074 DVDD.n5954 DVDD.n11 4.5005
R23075 DVDD.n29 DVDD.n24 4.5005
R23076 DVDD.n5954 DVDD.n24 4.5005
R23077 DVDD.n5954 DVDD.n12 4.5005
R23078 DVDD.n29 DVDD.n12 4.5005
R23079 DVDD.n5954 DVDD.n23 4.5005
R23080 DVDD.n29 DVDD.n23 4.5005
R23081 DVDD.n5954 DVDD.n13 4.5005
R23082 DVDD.n29 DVDD.n13 4.5005
R23083 DVDD.n29 DVDD.n22 4.5005
R23084 DVDD.n5954 DVDD.n22 4.5005
R23085 DVDD.n29 DVDD.n14 4.5005
R23086 DVDD.n5954 DVDD.n14 4.5005
R23087 DVDD.n29 DVDD.n21 4.5005
R23088 DVDD.n5954 DVDD.n21 4.5005
R23089 DVDD.n29 DVDD.n15 4.5005
R23090 DVDD.n5954 DVDD.n15 4.5005
R23091 DVDD.n5954 DVDD.n20 4.5005
R23092 DVDD.n29 DVDD.n20 4.5005
R23093 DVDD.n5954 DVDD.n16 4.5005
R23094 DVDD.n29 DVDD.n16 4.5005
R23095 DVDD.n5954 DVDD.n19 4.5005
R23096 DVDD.n29 DVDD.n19 4.5005
R23097 DVDD.n29 DVDD.n17 4.5005
R23098 DVDD.n5954 DVDD.n17 4.5005
R23099 DVDD.n29 DVDD.n18 4.5005
R23100 DVDD.n5954 DVDD.n18 4.5005
R23101 DVDD.n5954 DVDD.n8 4.5005
R23102 DVDD.n4701 DVDD.n972 4.5005
R23103 DVDD.n4701 DVDD.n974 4.5005
R23104 DVDD.n4701 DVDD.n971 4.5005
R23105 DVDD.n4701 DVDD.n4700 4.5005
R23106 DVDD.n4647 DVDD.n972 4.5005
R23107 DVDD.n984 DVDD.n974 4.5005
R23108 DVDD.n984 DVDD.n972 4.5005
R23109 DVDD.n4648 DVDD.n974 4.5005
R23110 DVDD.n4648 DVDD.n972 4.5005
R23111 DVDD.n983 DVDD.n974 4.5005
R23112 DVDD.n983 DVDD.n972 4.5005
R23113 DVDD.n4649 DVDD.n974 4.5005
R23114 DVDD.n4649 DVDD.n972 4.5005
R23115 DVDD.n982 DVDD.n972 4.5005
R23116 DVDD.n4650 DVDD.n972 4.5005
R23117 DVDD.n981 DVDD.n972 4.5005
R23118 DVDD.n4651 DVDD.n974 4.5005
R23119 DVDD.n4651 DVDD.n972 4.5005
R23120 DVDD.n980 DVDD.n974 4.5005
R23121 DVDD.n980 DVDD.n972 4.5005
R23122 DVDD.n4652 DVDD.n974 4.5005
R23123 DVDD.n4652 DVDD.n972 4.5005
R23124 DVDD.n979 DVDD.n974 4.5005
R23125 DVDD.n979 DVDD.n972 4.5005
R23126 DVDD.n4653 DVDD.n972 4.5005
R23127 DVDD.n978 DVDD.n972 4.5005
R23128 DVDD.n4654 DVDD.n972 4.5005
R23129 DVDD.n977 DVDD.n974 4.5005
R23130 DVDD.n977 DVDD.n972 4.5005
R23131 DVDD.n4655 DVDD.n974 4.5005
R23132 DVDD.n4655 DVDD.n972 4.5005
R23133 DVDD.n976 DVDD.n974 4.5005
R23134 DVDD.n976 DVDD.n972 4.5005
R23135 DVDD.n4699 DVDD.n974 4.5005
R23136 DVDD.n4699 DVDD.n972 4.5005
R23137 DVDD.n4654 DVDD.n974 4.5005
R23138 DVDD.n978 DVDD.n974 4.5005
R23139 DVDD.n4653 DVDD.n974 4.5005
R23140 DVDD.n981 DVDD.n974 4.5005
R23141 DVDD.n4650 DVDD.n974 4.5005
R23142 DVDD.n982 DVDD.n974 4.5005
R23143 DVDD.n4647 DVDD.n974 4.5005
R23144 DVDD.n972 DVDD.n267 4.5005
R23145 DVDD.n974 DVDD.n267 4.5005
R23146 DVDD.n971 DVDD.n267 4.5005
R23147 DVDD.n4700 DVDD.n267 4.5005
R23148 DVDD.n4708 DVDD.n946 4.5005
R23149 DVDD.n946 DVDD.n914 4.5005
R23150 DVDD.n4708 DVDD.n945 4.5005
R23151 DVDD.n945 DVDD.n914 4.5005
R23152 DVDD.n4708 DVDD.n947 4.5005
R23153 DVDD.n947 DVDD.n914 4.5005
R23154 DVDD.n224 DVDD.n222 4.5005
R23155 DVDD.n5707 DVDD.n222 4.5005
R23156 DVDD.n224 DVDD.n219 4.5005
R23157 DVDD.n5707 DVDD.n219 4.5005
R23158 DVDD.n224 DVDD.n221 4.5005
R23159 DVDD.n5707 DVDD.n221 4.5005
R23160 DVDD.n4346 DVDD.n1627 4.5005
R23161 DVDD.n4346 DVDD.n4345 4.5005
R23162 DVDD.n4345 DVDD.n1638 4.5005
R23163 DVDD.n4345 DVDD.n1641 4.5005
R23164 DVDD.n4345 DVDD.n1637 4.5005
R23165 DVDD.n4345 DVDD.n1643 4.5005
R23166 DVDD.n4345 DVDD.n1636 4.5005
R23167 DVDD.n4345 DVDD.n1645 4.5005
R23168 DVDD.n4345 DVDD.n1635 4.5005
R23169 DVDD.n4345 DVDD.n1647 4.5005
R23170 DVDD.n4345 DVDD.n1634 4.5005
R23171 DVDD.n4345 DVDD.n1649 4.5005
R23172 DVDD.n4345 DVDD.n1633 4.5005
R23173 DVDD.n4345 DVDD.n1651 4.5005
R23174 DVDD.n4345 DVDD.n1632 4.5005
R23175 DVDD.n4345 DVDD.n1653 4.5005
R23176 DVDD.n4345 DVDD.n1631 4.5005
R23177 DVDD.n4345 DVDD.n1655 4.5005
R23178 DVDD.n4345 DVDD.n1630 4.5005
R23179 DVDD.n4345 DVDD.n1657 4.5005
R23180 DVDD.n4345 DVDD.n1629 4.5005
R23181 DVDD.n4344 DVDD.n4342 4.5005
R23182 DVDD.n4345 DVDD.n4344 4.5005
R23183 DVDD.n4746 DVDD.n894 4.5005
R23184 DVDD.n4744 DVDD.n893 4.5005
R23185 DVDD.n4746 DVDD.n893 4.5005
R23186 DVDD.n4744 DVDD.n895 4.5005
R23187 DVDD.n4746 DVDD.n895 4.5005
R23188 DVDD.n4744 DVDD.n892 4.5005
R23189 DVDD.n4746 DVDD.n892 4.5005
R23190 DVDD.n4745 DVDD.n4744 4.5005
R23191 DVDD.n4746 DVDD.n4745 4.5005
R23192 DVDD.n4744 DVDD.n894 4.5005
R23193 DVDD.n4775 DVDD.n737 4.5005
R23194 DVDD.n4773 DVDD.n736 4.5005
R23195 DVDD.n4775 DVDD.n736 4.5005
R23196 DVDD.n4773 DVDD.n738 4.5005
R23197 DVDD.n4775 DVDD.n738 4.5005
R23198 DVDD.n4773 DVDD.n735 4.5005
R23199 DVDD.n4775 DVDD.n735 4.5005
R23200 DVDD.n4774 DVDD.n4773 4.5005
R23201 DVDD.n4775 DVDD.n4774 4.5005
R23202 DVDD.n4773 DVDD.n737 4.5005
R23203 DVDD.n5021 DVDD.n584 4.5005
R23204 DVDD.n5022 DVDD.n592 4.5005
R23205 DVDD.n592 DVDD.n584 4.5005
R23206 DVDD.n5022 DVDD.n590 4.5005
R23207 DVDD.n590 DVDD.n584 4.5005
R23208 DVDD.n5022 DVDD.n593 4.5005
R23209 DVDD.n593 DVDD.n584 4.5005
R23210 DVDD.n5022 DVDD.n589 4.5005
R23211 DVDD.n589 DVDD.n584 4.5005
R23212 DVDD.n5022 DVDD.n5021 4.5005
R23213 DVDD.n5097 DVDD.n570 4.5005
R23214 DVDD.n5096 DVDD.n5088 4.5005
R23215 DVDD.n5088 DVDD.n570 4.5005
R23216 DVDD.n5096 DVDD.n573 4.5005
R23217 DVDD.n573 DVDD.n570 4.5005
R23218 DVDD.n5096 DVDD.n5095 4.5005
R23219 DVDD.n5095 DVDD.n570 4.5005
R23220 DVDD.n5096 DVDD.n572 4.5005
R23221 DVDD.n572 DVDD.n570 4.5005
R23222 DVDD.n5097 DVDD.n5096 4.5005
R23223 DVDD.n5735 DVDD.n193 4.5005
R23224 DVDD.n5736 DVDD.n196 4.5005
R23225 DVDD.n5736 DVDD.n5735 4.5005
R23226 DVDD.n5730 DVDD.n196 4.5005
R23227 DVDD.n5735 DVDD.n5730 4.5005
R23228 DVDD.n198 DVDD.n196 4.5005
R23229 DVDD.n5735 DVDD.n198 4.5005
R23230 DVDD.n5734 DVDD.n196 4.5005
R23231 DVDD.n5735 DVDD.n5734 4.5005
R23232 DVDD.n196 DVDD.n193 4.5005
R23233 DVDD.n5706 DVDD.n233 4.5005
R23234 DVDD.n5706 DVDD.n235 4.5005
R23235 DVDD.n241 DVDD.n235 4.5005
R23236 DVDD.n5704 DVDD.n235 4.5005
R23237 DVDD.n241 DVDD.n233 4.5005
R23238 DVDD.n5704 DVDD.n233 4.5005
R23239 DVDD.n5704 DVDD.n232 4.5005
R23240 DVDD.n241 DVDD.n232 4.5005
R23241 DVDD.n5706 DVDD.n232 4.5005
R23242 DVDD.n5704 DVDD.n236 4.5005
R23243 DVDD.n241 DVDD.n236 4.5005
R23244 DVDD.n5706 DVDD.n236 4.5005
R23245 DVDD.n5704 DVDD.n231 4.5005
R23246 DVDD.n241 DVDD.n231 4.5005
R23247 DVDD.n5706 DVDD.n231 4.5005
R23248 DVDD.n5706 DVDD.n237 4.5005
R23249 DVDD.n241 DVDD.n237 4.5005
R23250 DVDD.n5704 DVDD.n237 4.5005
R23251 DVDD.n5706 DVDD.n230 4.5005
R23252 DVDD.n241 DVDD.n230 4.5005
R23253 DVDD.n5704 DVDD.n230 4.5005
R23254 DVDD.n5706 DVDD.n238 4.5005
R23255 DVDD.n241 DVDD.n238 4.5005
R23256 DVDD.n5704 DVDD.n238 4.5005
R23257 DVDD.n5706 DVDD.n229 4.5005
R23258 DVDD.n241 DVDD.n229 4.5005
R23259 DVDD.n5704 DVDD.n229 4.5005
R23260 DVDD.n5704 DVDD.n239 4.5005
R23261 DVDD.n241 DVDD.n239 4.5005
R23262 DVDD.n5706 DVDD.n239 4.5005
R23263 DVDD.n5704 DVDD.n228 4.5005
R23264 DVDD.n241 DVDD.n228 4.5005
R23265 DVDD.n5706 DVDD.n228 4.5005
R23266 DVDD.n5705 DVDD.n5704 4.5005
R23267 DVDD.n5705 DVDD.n241 4.5005
R23268 DVDD.n5706 DVDD.n5705 4.5005
R23269 DVDD.n226 DVDD.n218 4.5005
R23270 DVDD.n224 DVDD.n218 4.5005
R23271 DVDD.n5707 DVDD.n218 4.5005
R23272 DVDD.n5709 DVDD.n221 4.5005
R23273 DVDD.n226 DVDD.n221 4.5005
R23274 DVDD.n5709 DVDD.n219 4.5005
R23275 DVDD.n226 DVDD.n219 4.5005
R23276 DVDD.n226 DVDD.n222 4.5005
R23277 DVDD.n5709 DVDD.n222 4.5005
R23278 DVDD.n5709 DVDD.n218 4.5005
R23279 DVDD.n5709 DVDD.n5708 4.5005
R23280 DVDD.n5708 DVDD.n226 4.5005
R23281 DVDD.n5708 DVDD.n224 4.5005
R23282 DVDD.n5708 DVDD.n5707 4.5005
R23283 DVDD.n943 DVDD.n920 4.5005
R23284 DVDD.n4710 DVDD.n920 4.5005
R23285 DVDD.n4712 DVDD.n920 4.5005
R23286 DVDD.n943 DVDD.n923 4.5005
R23287 DVDD.n4710 DVDD.n923 4.5005
R23288 DVDD.n4712 DVDD.n923 4.5005
R23289 DVDD.n4712 DVDD.n919 4.5005
R23290 DVDD.n4712 DVDD.n924 4.5005
R23291 DVDD.n4712 DVDD.n918 4.5005
R23292 DVDD.n943 DVDD.n925 4.5005
R23293 DVDD.n4710 DVDD.n925 4.5005
R23294 DVDD.n4712 DVDD.n925 4.5005
R23295 DVDD.n943 DVDD.n917 4.5005
R23296 DVDD.n4710 DVDD.n917 4.5005
R23297 DVDD.n4712 DVDD.n917 4.5005
R23298 DVDD.n943 DVDD.n926 4.5005
R23299 DVDD.n4710 DVDD.n926 4.5005
R23300 DVDD.n4712 DVDD.n926 4.5005
R23301 DVDD.n943 DVDD.n916 4.5005
R23302 DVDD.n4710 DVDD.n916 4.5005
R23303 DVDD.n4712 DVDD.n916 4.5005
R23304 DVDD.n4712 DVDD.n941 4.5005
R23305 DVDD.n4712 DVDD.n915 4.5005
R23306 DVDD.n4710 DVDD.n915 4.5005
R23307 DVDD.n943 DVDD.n915 4.5005
R23308 DVDD.n4710 DVDD.n941 4.5005
R23309 DVDD.n943 DVDD.n941 4.5005
R23310 DVDD.n4710 DVDD.n918 4.5005
R23311 DVDD.n943 DVDD.n918 4.5005
R23312 DVDD.n4710 DVDD.n924 4.5005
R23313 DVDD.n943 DVDD.n924 4.5005
R23314 DVDD.n4710 DVDD.n919 4.5005
R23315 DVDD.n943 DVDD.n919 4.5005
R23316 DVDD.n4712 DVDD.n4711 4.5005
R23317 DVDD.n4711 DVDD.n943 4.5005
R23318 DVDD.n4711 DVDD.n4710 4.5005
R23319 DVDD.n944 DVDD.n922 4.5005
R23320 DVDD.n944 DVDD.n910 4.5005
R23321 DVDD.n944 DVDD.n914 4.5005
R23322 DVDD.n4708 DVDD.n944 4.5005
R23323 DVDD.n4708 DVDD.n4707 4.5005
R23324 DVDD.n4707 DVDD.n914 4.5005
R23325 DVDD.n4707 DVDD.n922 4.5005
R23326 DVDD.n4707 DVDD.n910 4.5005
R23327 DVDD.n946 DVDD.n922 4.5005
R23328 DVDD.n946 DVDD.n910 4.5005
R23329 DVDD.n945 DVDD.n922 4.5005
R23330 DVDD.n945 DVDD.n910 4.5005
R23331 DVDD.n947 DVDD.n922 4.5005
R23332 DVDD.n947 DVDD.n910 4.5005
R23333 DVDD.n2601 DVDD.n2512 4.39376
R23334 DVDD.n3450 DVDD.n2685 4.29432
R23335 DVDD.n3115 DVDD.n3112 4.03391
R23336 DVDD.n2516 DVDD.t9 3.97738
R23337 DVDD.n3147 DVDD.n3146 3.90569
R23338 DVDD.n2517 DVDD.t54 3.75601
R23339 DVDD.n2539 DVDD.t58 3.75601
R23340 DVDD.t220 DVDD.n3063 3.6505
R23341 DVDD.t215 DVDD.n3042 3.6505
R23342 DVDD.t216 DVDD.n2998 3.6505
R23343 DVDD.t214 DVDD.n3017 3.6505
R23344 DVDD.n5491 DVDD.n5490 3.24952
R23345 DVDD.n5664 DVDD.n256 3.24952
R23346 DVDD.n3150 DVDD.n3149 3.1505
R23347 DVDD.n2572 DVDD.n2569 3.148
R23348 DVDD.n2564 DVDD.n2561 3.148
R23349 DVDD.n2569 DVDD.n2568 3.148
R23350 DVDD.n2564 DVDD.n2562 3.148
R23351 DVDD.n2569 DVDD.n2567 3.148
R23352 DVDD.n2564 DVDD.n2563 3.148
R23353 DVDD.n2569 DVDD.n2566 3.148
R23354 DVDD.n2564 DVDD.n2555 3.148
R23355 DVDD.n2544 DVDD.n2542 3.14761
R23356 DVDD.n2538 DVDD.n2537 3.14761
R23357 DVDD.n2588 DVDD.n2585 3.14761
R23358 DVDD.n2538 DVDD.n2536 3.14761
R23359 DVDD.n2588 DVDD.n2587 3.14761
R23360 DVDD.n2538 DVDD.n2535 3.14761
R23361 DVDD.n2588 DVDD.n2534 3.14761
R23362 DVDD.n2573 DVDD.n2571 2.98283
R23363 DVDD.n2573 DVDD.n2565 2.98283
R23364 DVDD.n2573 DVDD.n2552 2.98283
R23365 DVDD.n2546 DVDD.n2545 2.98283
R23366 DVDD.n2545 DVDD.n2529 2.98283
R23367 DVDD.n2570 DVDD.n2551 2.98283
R23368 DVDD.n2559 DVDD.n2551 2.98283
R23369 DVDD.n2543 DVDD.n2527 2.98283
R23370 DVDD.n2586 DVDD.n2532 2.98283
R23371 DVDD.n2581 DVDD.n2558 2.98283
R23372 DVDD.n3219 DVDD.n3111 2.94507
R23373 DVDD.n3063 DVDD.n3062 2.85774
R23374 DVDD.n3042 DVDD.n3041 2.85774
R23375 DVDD.n2998 DVDD.n2997 2.85774
R23376 DVDD.n3017 DVDD.n3016 2.85774
R23377 DVDD.n2516 DVDD.n2515 2.76877
R23378 DVDD.n3149 DVDD.n3144 2.76479
R23379 DVDD.n3221 DVDD.n3111 2.74405
R23380 DVDD.n4237 DVDD.n1710 2.69653
R23381 DVDD.n3450 DVDD.n3449 2.63997
R23382 DVDD.n3062 DVDD 2.57263
R23383 DVDD.n3041 DVDD 2.57263
R23384 DVDD.n2997 DVDD 2.57263
R23385 DVDD.n3016 DVDD 2.57263
R23386 DVDD.n3445 DVDD.n2688 2.56264
R23387 DVDD.n1948 DVDD.n1947 2.54396
R23388 DVDD.n2600 DVDD.n2599 2.52684
R23389 DVDD DVDD.n4202 2.51792
R23390 DVDD.n1885 DVDD 2.51792
R23391 DVDD.n2972 DVDD.n2970 2.45964
R23392 DVDD.n3218 DVDD.n3217 2.42304
R23393 DVDD.n3153 DVDD.n3152 2.42304
R23394 DVDD.n3218 DVDD.n3110 2.38608
R23395 DVDD.n3153 DVDD.n3143 2.38608
R23396 DVDD.n3695 DVDD.t159 2.32044
R23397 DVDD.n3694 DVDD.t5 2.32044
R23398 DVDD.n5708 DVDD.n223 2.25251
R23399 DVDD.n961 DVDD.n944 2.25251
R23400 DVDD.n5921 DVDD.n5920 2.25174
R23401 DVDD.n5425 DVDD.n327 2.25174
R23402 DVDD.n5732 DVDD.n5731 2.2505
R23403 DVDD.n195 DVDD.n194 2.2505
R23404 DVDD.n5738 DVDD.n5737 2.2505
R23405 DVDD.n5740 DVDD.n5739 2.2505
R23406 DVDD.n5741 DVDD.n192 2.2505
R23407 DVDD.n5743 DVDD.n5742 2.2505
R23408 DVDD.n5745 DVDD.n5744 2.2505
R23409 DVDD.n5747 DVDD.n5746 2.2505
R23410 DVDD.n5749 DVDD.n5748 2.2505
R23411 DVDD.n5751 DVDD.n5750 2.2505
R23412 DVDD.n5753 DVDD.n5752 2.2505
R23413 DVDD.n5755 DVDD.n5754 2.2505
R23414 DVDD.n5757 DVDD.n5756 2.2505
R23415 DVDD.n5759 DVDD.n5758 2.2505
R23416 DVDD.n5761 DVDD.n5760 2.2505
R23417 DVDD.n5763 DVDD.n5762 2.2505
R23418 DVDD.n5765 DVDD.n5764 2.2505
R23419 DVDD.n5767 DVDD.n5766 2.2505
R23420 DVDD.n5769 DVDD.n5768 2.2505
R23421 DVDD.n5771 DVDD.n5770 2.2505
R23422 DVDD.n5773 DVDD.n5772 2.2505
R23423 DVDD.n5774 DVDD.n190 2.2505
R23424 DVDD.n5783 DVDD.n5782 2.2505
R23425 DVDD.n5781 DVDD.n191 2.2505
R23426 DVDD.n5780 DVDD.n5779 2.2505
R23427 DVDD.n5778 DVDD.n5777 2.2505
R23428 DVDD.n5776 DVDD.n5775 2.2505
R23429 DVDD.n168 DVDD.n167 2.2505
R23430 DVDD.n5788 DVDD.n5787 2.2505
R23431 DVDD.n5790 DVDD.n5789 2.2505
R23432 DVDD.n5791 DVDD.n165 2.2505
R23433 DVDD.n5793 DVDD.n5792 2.2505
R23434 DVDD.n5794 DVDD.n164 2.2505
R23435 DVDD.n5834 DVDD.n5833 2.2505
R23436 DVDD.n5832 DVDD.n5831 2.2505
R23437 DVDD.n5830 DVDD.n5829 2.2505
R23438 DVDD.n5828 DVDD.n5827 2.2505
R23439 DVDD.n5826 DVDD.n5825 2.2505
R23440 DVDD.n5824 DVDD.n5823 2.2505
R23441 DVDD.n5822 DVDD.n5821 2.2505
R23442 DVDD.n5820 DVDD.n5819 2.2505
R23443 DVDD.n5818 DVDD.n5817 2.2505
R23444 DVDD.n5816 DVDD.n5815 2.2505
R23445 DVDD.n5814 DVDD.n5813 2.2505
R23446 DVDD.n5812 DVDD.n5811 2.2505
R23447 DVDD.n5810 DVDD.n5809 2.2505
R23448 DVDD.n5808 DVDD.n5807 2.2505
R23449 DVDD.n5806 DVDD.n5805 2.2505
R23450 DVDD.n5804 DVDD.n5803 2.2505
R23451 DVDD.n5802 DVDD.n5801 2.2505
R23452 DVDD.n5800 DVDD.n5799 2.2505
R23453 DVDD.n5798 DVDD.n5797 2.2505
R23454 DVDD.n5796 DVDD.n5795 2.2505
R23455 DVDD.n142 DVDD.n141 2.2505
R23456 DVDD.n5839 DVDD.n5838 2.2505
R23457 DVDD.n5841 DVDD.n5840 2.2505
R23458 DVDD.n5842 DVDD.n139 2.2505
R23459 DVDD.n5844 DVDD.n5843 2.2505
R23460 DVDD.n5846 DVDD.n5845 2.2505
R23461 DVDD.n5848 DVDD.n5847 2.2505
R23462 DVDD.n5094 DVDD.n5093 2.2505
R23463 DVDD.n5092 DVDD.n5091 2.2505
R23464 DVDD.n5090 DVDD.n569 2.2505
R23465 DVDD.n5098 DVDD.n568 2.2505
R23466 DVDD.n5100 DVDD.n5099 2.2505
R23467 DVDD.n5101 DVDD.n566 2.2505
R23468 DVDD.n5242 DVDD.n5241 2.2505
R23469 DVDD.n5240 DVDD.n567 2.2505
R23470 DVDD.n5239 DVDD.n5238 2.2505
R23471 DVDD.n5237 DVDD.n5236 2.2505
R23472 DVDD.n5235 DVDD.n5234 2.2505
R23473 DVDD.n5233 DVDD.n5232 2.2505
R23474 DVDD.n5231 DVDD.n5230 2.2505
R23475 DVDD.n5229 DVDD.n5228 2.2505
R23476 DVDD.n5227 DVDD.n5226 2.2505
R23477 DVDD.n5225 DVDD.n5224 2.2505
R23478 DVDD.n5223 DVDD.n5222 2.2505
R23479 DVDD.n5221 DVDD.n5220 2.2505
R23480 DVDD.n5219 DVDD.n5218 2.2505
R23481 DVDD.n5217 DVDD.n5216 2.2505
R23482 DVDD.n5215 DVDD.n5214 2.2505
R23483 DVDD.n5213 DVDD.n5212 2.2505
R23484 DVDD.n5211 DVDD.n5210 2.2505
R23485 DVDD.n5209 DVDD.n5208 2.2505
R23486 DVDD.n5207 DVDD.n5206 2.2505
R23487 DVDD.n5205 DVDD.n5204 2.2505
R23488 DVDD.n5203 DVDD.n5202 2.2505
R23489 DVDD.n5201 DVDD.n5200 2.2505
R23490 DVDD.n5199 DVDD.n5198 2.2505
R23491 DVDD.n5197 DVDD.n5196 2.2505
R23492 DVDD.n5195 DVDD.n5102 2.2505
R23493 DVDD.n5194 DVDD.n5193 2.2505
R23494 DVDD.n5192 DVDD.n5191 2.2505
R23495 DVDD.n5190 DVDD.n5189 2.2505
R23496 DVDD.n5188 DVDD.n5187 2.2505
R23497 DVDD.n5186 DVDD.n5185 2.2505
R23498 DVDD.n5184 DVDD.n5183 2.2505
R23499 DVDD.n5182 DVDD.n5181 2.2505
R23500 DVDD.n5180 DVDD.n5179 2.2505
R23501 DVDD.n5178 DVDD.n5177 2.2505
R23502 DVDD.n5176 DVDD.n5175 2.2505
R23503 DVDD.n5174 DVDD.n5173 2.2505
R23504 DVDD.n5172 DVDD.n5171 2.2505
R23505 DVDD.n5170 DVDD.n5169 2.2505
R23506 DVDD.n5168 DVDD.n5167 2.2505
R23507 DVDD.n5166 DVDD.n5165 2.2505
R23508 DVDD.n5164 DVDD.n5163 2.2505
R23509 DVDD.n5162 DVDD.n5161 2.2505
R23510 DVDD.n5160 DVDD.n5159 2.2505
R23511 DVDD.n5158 DVDD.n5157 2.2505
R23512 DVDD.n5156 DVDD.n5155 2.2505
R23513 DVDD.n5154 DVDD.n5153 2.2505
R23514 DVDD.n5152 DVDD.n5151 2.2505
R23515 DVDD.n5150 DVDD.n473 2.2505
R23516 DVDD.n5149 DVDD.n474 2.2505
R23517 DVDD.n5148 DVDD.n5147 2.2505
R23518 DVDD.n5146 DVDD.n5103 2.2505
R23519 DVDD.n5145 DVDD.n5144 2.2505
R23520 DVDD.n5143 DVDD.n5142 2.2505
R23521 DVDD.n5140 DVDD.n5105 2.2505
R23522 DVDD.n598 DVDD.n597 2.2505
R23523 DVDD.n600 DVDD.n599 2.2505
R23524 DVDD.n601 DVDD.n594 2.2505
R23525 DVDD.n5020 DVDD.n5019 2.2505
R23526 DVDD.n5018 DVDD.n595 2.2505
R23527 DVDD.n5017 DVDD.n5016 2.2505
R23528 DVDD.n604 DVDD.n602 2.2505
R23529 DVDD.n629 DVDD.n628 2.2505
R23530 DVDD.n631 DVDD.n630 2.2505
R23531 DVDD.n633 DVDD.n632 2.2505
R23532 DVDD.n635 DVDD.n634 2.2505
R23533 DVDD.n637 DVDD.n636 2.2505
R23534 DVDD.n639 DVDD.n638 2.2505
R23535 DVDD.n641 DVDD.n640 2.2505
R23536 DVDD.n643 DVDD.n642 2.2505
R23537 DVDD.n645 DVDD.n644 2.2505
R23538 DVDD.n647 DVDD.n646 2.2505
R23539 DVDD.n649 DVDD.n648 2.2505
R23540 DVDD.n651 DVDD.n650 2.2505
R23541 DVDD.n653 DVDD.n652 2.2505
R23542 DVDD.n655 DVDD.n654 2.2505
R23543 DVDD.n657 DVDD.n656 2.2505
R23544 DVDD.n659 DVDD.n658 2.2505
R23545 DVDD.n661 DVDD.n660 2.2505
R23546 DVDD.n663 DVDD.n662 2.2505
R23547 DVDD.n665 DVDD.n664 2.2505
R23548 DVDD.n667 DVDD.n666 2.2505
R23549 DVDD.n669 DVDD.n668 2.2505
R23550 DVDD.n670 DVDD.n626 2.2505
R23551 DVDD.n5012 DVDD.n5011 2.2505
R23552 DVDD.n5010 DVDD.n627 2.2505
R23553 DVDD.n5009 DVDD.n5008 2.2505
R23554 DVDD.n673 DVDD.n671 2.2505
R23555 DVDD.n4953 DVDD.n4952 2.2505
R23556 DVDD.n4955 DVDD.n4954 2.2505
R23557 DVDD.n4957 DVDD.n4956 2.2505
R23558 DVDD.n4959 DVDD.n4958 2.2505
R23559 DVDD.n4961 DVDD.n4960 2.2505
R23560 DVDD.n4963 DVDD.n4962 2.2505
R23561 DVDD.n4965 DVDD.n4964 2.2505
R23562 DVDD.n4967 DVDD.n4966 2.2505
R23563 DVDD.n4969 DVDD.n4968 2.2505
R23564 DVDD.n4971 DVDD.n4970 2.2505
R23565 DVDD.n4973 DVDD.n4972 2.2505
R23566 DVDD.n4975 DVDD.n4974 2.2505
R23567 DVDD.n4977 DVDD.n4976 2.2505
R23568 DVDD.n4979 DVDD.n4978 2.2505
R23569 DVDD.n4981 DVDD.n4980 2.2505
R23570 DVDD.n4983 DVDD.n4982 2.2505
R23571 DVDD.n4985 DVDD.n4984 2.2505
R23572 DVDD.n4987 DVDD.n4986 2.2505
R23573 DVDD.n4989 DVDD.n4988 2.2505
R23574 DVDD.n4991 DVDD.n4990 2.2505
R23575 DVDD.n4992 DVDD.n4951 2.2505
R23576 DVDD.n5004 DVDD.n5003 2.2505
R23577 DVDD.n5002 DVDD.n5001 2.2505
R23578 DVDD.n5000 DVDD.n4993 2.2505
R23579 DVDD.n4999 DVDD.n4998 2.2505
R23580 DVDD.n4997 DVDD.n4996 2.2505
R23581 DVDD.n4995 DVDD.n4994 2.2505
R23582 DVDD.n877 DVDD.n876 2.2505
R23583 DVDD.n875 DVDD.n874 2.2505
R23584 DVDD.n873 DVDD.n872 2.2505
R23585 DVDD.n871 DVDD.n870 2.2505
R23586 DVDD.n869 DVDD.n868 2.2505
R23587 DVDD.n867 DVDD.n726 2.2505
R23588 DVDD.n866 DVDD.n727 2.2505
R23589 DVDD.n865 DVDD.n864 2.2505
R23590 DVDD.n863 DVDD.n862 2.2505
R23591 DVDD.n861 DVDD.n860 2.2505
R23592 DVDD.n859 DVDD.n858 2.2505
R23593 DVDD.n857 DVDD.n856 2.2505
R23594 DVDD.n855 DVDD.n854 2.2505
R23595 DVDD.n853 DVDD.n852 2.2505
R23596 DVDD.n851 DVDD.n850 2.2505
R23597 DVDD.n849 DVDD.n848 2.2505
R23598 DVDD.n847 DVDD.n846 2.2505
R23599 DVDD.n845 DVDD.n844 2.2505
R23600 DVDD.n843 DVDD.n842 2.2505
R23601 DVDD.n841 DVDD.n840 2.2505
R23602 DVDD.n839 DVDD.n838 2.2505
R23603 DVDD.n837 DVDD.n836 2.2505
R23604 DVDD.n835 DVDD.n834 2.2505
R23605 DVDD.n833 DVDD.n832 2.2505
R23606 DVDD.n831 DVDD.n830 2.2505
R23607 DVDD.n829 DVDD.n828 2.2505
R23608 DVDD.n827 DVDD.n826 2.2505
R23609 DVDD.n825 DVDD.n824 2.2505
R23610 DVDD.n823 DVDD.n822 2.2505
R23611 DVDD.n821 DVDD.n820 2.2505
R23612 DVDD.n819 DVDD.n739 2.2505
R23613 DVDD.n818 DVDD.n817 2.2505
R23614 DVDD.n816 DVDD.n815 2.2505
R23615 DVDD.n813 DVDD.n741 2.2505
R23616 DVDD.n811 DVDD.n810 2.2505
R23617 DVDD.n809 DVDD.n742 2.2505
R23618 DVDD.n808 DVDD.n807 2.2505
R23619 DVDD.n805 DVDD.n743 2.2505
R23620 DVDD.n803 DVDD.n802 2.2505
R23621 DVDD.n801 DVDD.n800 2.2505
R23622 DVDD.n798 DVDD.n746 2.2505
R23623 DVDD.n796 DVDD.n795 2.2505
R23624 DVDD.n794 DVDD.n793 2.2505
R23625 DVDD.n792 DVDD.n748 2.2505
R23626 DVDD.n790 DVDD.n789 2.2505
R23627 DVDD.n788 DVDD.n787 2.2505
R23628 DVDD.n785 DVDD.n750 2.2505
R23629 DVDD.n783 DVDD.n782 2.2505
R23630 DVDD.n781 DVDD.n780 2.2505
R23631 DVDD.n778 DVDD.n752 2.2505
R23632 DVDD.n776 DVDD.n775 2.2505
R23633 DVDD.n774 DVDD.n753 2.2505
R23634 DVDD.n773 DVDD.n772 2.2505
R23635 DVDD.n770 DVDD.n754 2.2505
R23636 DVDD.n768 DVDD.n767 2.2505
R23637 DVDD.n766 DVDD.n765 2.2505
R23638 DVDD.n764 DVDD.n757 2.2505
R23639 DVDD.n763 DVDD.n762 2.2505
R23640 DVDD.n761 DVDD.n760 2.2505
R23641 DVDD.n759 DVDD.n758 2.2505
R23642 DVDD.n1060 DVDD.n1059 2.2505
R23643 DVDD.n1062 DVDD.n1061 2.2505
R23644 DVDD.n1064 DVDD.n1063 2.2505
R23645 DVDD.n1066 DVDD.n1065 2.2505
R23646 DVDD.n1068 DVDD.n1067 2.2505
R23647 DVDD.n1069 DVDD.n1057 2.2505
R23648 DVDD.n4615 DVDD.n4614 2.2505
R23649 DVDD.n4613 DVDD.n1058 2.2505
R23650 DVDD.n4612 DVDD.n4611 2.2505
R23651 DVDD.n4610 DVDD.n4609 2.2505
R23652 DVDD.n4608 DVDD.n4607 2.2505
R23653 DVDD.n4606 DVDD.n4605 2.2505
R23654 DVDD.n4604 DVDD.n4603 2.2505
R23655 DVDD.n4602 DVDD.n4601 2.2505
R23656 DVDD.n4600 DVDD.n4599 2.2505
R23657 DVDD.n4598 DVDD.n4597 2.2505
R23658 DVDD.n4596 DVDD.n4595 2.2505
R23659 DVDD.n4594 DVDD.n4593 2.2505
R23660 DVDD.n4592 DVDD.n4591 2.2505
R23661 DVDD.n4590 DVDD.n4589 2.2505
R23662 DVDD.n4588 DVDD.n4587 2.2505
R23663 DVDD.n4586 DVDD.n4585 2.2505
R23664 DVDD.n4584 DVDD.n4583 2.2505
R23665 DVDD.n4582 DVDD.n4581 2.2505
R23666 DVDD.n4580 DVDD.n4579 2.2505
R23667 DVDD.n4578 DVDD.n4577 2.2505
R23668 DVDD.n4576 DVDD.n4575 2.2505
R23669 DVDD.n4574 DVDD.n4573 2.2505
R23670 DVDD.n4572 DVDD.n4571 2.2505
R23671 DVDD.n4570 DVDD.n4569 2.2505
R23672 DVDD.n4568 DVDD.n1070 2.2505
R23673 DVDD.n4567 DVDD.n4566 2.2505
R23674 DVDD.n4565 DVDD.n4564 2.2505
R23675 DVDD.n1074 DVDD.n1072 2.2505
R23676 DVDD.n4511 DVDD.n4510 2.2505
R23677 DVDD.n4513 DVDD.n4512 2.2505
R23678 DVDD.n4515 DVDD.n4514 2.2505
R23679 DVDD.n4517 DVDD.n4516 2.2505
R23680 DVDD.n4519 DVDD.n4518 2.2505
R23681 DVDD.n4521 DVDD.n4520 2.2505
R23682 DVDD.n4523 DVDD.n4522 2.2505
R23683 DVDD.n4525 DVDD.n4524 2.2505
R23684 DVDD.n4527 DVDD.n4526 2.2505
R23685 DVDD.n4529 DVDD.n4528 2.2505
R23686 DVDD.n4531 DVDD.n4530 2.2505
R23687 DVDD.n4533 DVDD.n4532 2.2505
R23688 DVDD.n4535 DVDD.n4534 2.2505
R23689 DVDD.n4537 DVDD.n4536 2.2505
R23690 DVDD.n4539 DVDD.n4538 2.2505
R23691 DVDD.n4541 DVDD.n4540 2.2505
R23692 DVDD.n4543 DVDD.n4542 2.2505
R23693 DVDD.n4545 DVDD.n4544 2.2505
R23694 DVDD.n4547 DVDD.n4546 2.2505
R23695 DVDD.n4548 DVDD.n4509 2.2505
R23696 DVDD.n4560 DVDD.n4559 2.2505
R23697 DVDD.n4558 DVDD.n4557 2.2505
R23698 DVDD.n4556 DVDD.n4549 2.2505
R23699 DVDD.n4555 DVDD.n4554 2.2505
R23700 DVDD.n4553 DVDD.n4552 2.2505
R23701 DVDD.n4551 DVDD.n4550 2.2505
R23702 DVDD.n3044 DVDD.n3018 2.2505
R23703 DVDD.n3065 DVDD.n2999 2.2505
R23704 DVDD.n3044 DVDD.n3043 2.2505
R23705 DVDD.n3065 DVDD.n3064 2.2505
R23706 DVDD.n3174 DVDD.n3139 2.2505
R23707 DVDD.n3202 DVDD.n3201 2.2505
R23708 DVDD.n3125 DVDD.n3124 2.2505
R23709 DVDD.n3177 DVDD.n3176 2.2505
R23710 DVDD.n3179 DVDD.n3178 2.2505
R23711 DVDD.n3248 DVDD.n3084 2.2505
R23712 DVDD.n3247 DVDD.n3246 2.2505
R23713 DVDD.n3237 DVDD.n3088 2.2505
R23714 DVDD.n3239 DVDD.n3238 2.2505
R23715 DVDD.n3236 DVDD.n3235 2.2505
R23716 DVDD.n3211 DVDD.n2962 2.2505
R23717 DVDD.n3233 DVDD.n3098 2.2505
R23718 DVDD.n3186 DVDD.n3185 2.2505
R23719 DVDD.n3241 DVDD.n3093 2.2505
R23720 DVDD.n3244 DVDD.n3090 2.2505
R23721 DVDD.n3254 DVDD.n3082 2.2505
R23722 DVDD.n3086 DVDD.n2962 2.2505
R23723 DVDD.n3245 DVDD.n3244 2.2505
R23724 DVDD.n3234 DVDD.n3233 2.2505
R23725 DVDD.n3185 DVDD.n3094 2.2505
R23726 DVDD.n3241 DVDD.n3240 2.2505
R23727 DVDD.n3254 DVDD.n3253 2.2505
R23728 DVDD.n3209 DVDD.n3208 2.2505
R23729 DVDD.n3165 DVDD.n3135 2.2505
R23730 DVDD.n3182 DVDD.n3181 2.2505
R23731 DVDD.n3141 DVDD.n3130 2.2505
R23732 DVDD.n3198 DVDD.n3197 2.2505
R23733 DVDD.n3131 DVDD.n3078 2.2505
R23734 DVDD.n3181 DVDD.n3180 2.2505
R23735 DVDD.n3142 DVDD.n3141 2.2505
R23736 DVDD.n3199 DVDD.n3198 2.2505
R23737 DVDD.n3200 DVDD.n3078 2.2505
R23738 DVDD.n3208 DVDD.n3207 2.2505
R23739 DVDD.n3165 DVDD.n3164 2.2505
R23740 DVDD.n1391 DVDD.n1390 2.2505
R23741 DVDD.n1315 DVDD.n1314 2.2505
R23742 DVDD.n5503 DVDD.n225 2.2505
R23743 DVDD.n5505 DVDD.n5504 2.2505
R23744 DVDD.n5508 DVDD.n5507 2.2505
R23745 DVDD.n5510 DVDD.n5509 2.2505
R23746 DVDD.n5512 DVDD.n5511 2.2505
R23747 DVDD.n5514 DVDD.n5513 2.2505
R23748 DVDD.n5515 DVDD.n28 2.2505
R23749 DVDD.n5516 DVDD.n30 2.2505
R23750 DVDD.n5518 DVDD.n5517 2.2505
R23751 DVDD.n5520 DVDD.n5519 2.2505
R23752 DVDD.n5522 DVDD.n5521 2.2505
R23753 DVDD.n5524 DVDD.n5523 2.2505
R23754 DVDD.n5526 DVDD.n5525 2.2505
R23755 DVDD.n5528 DVDD.n5527 2.2505
R23756 DVDD.n5530 DVDD.n5529 2.2505
R23757 DVDD.n5532 DVDD.n5531 2.2505
R23758 DVDD.n5534 DVDD.n5533 2.2505
R23759 DVDD.n5536 DVDD.n5535 2.2505
R23760 DVDD.n5538 DVDD.n5537 2.2505
R23761 DVDD.n5541 DVDD.n5540 2.2505
R23762 DVDD.n5543 DVDD.n5542 2.2505
R23763 DVDD.n5545 DVDD.n5544 2.2505
R23764 DVDD.n5547 DVDD.n5546 2.2505
R23765 DVDD.n5549 DVDD.n5548 2.2505
R23766 DVDD.n5551 DVDD.n5550 2.2505
R23767 DVDD.n5553 DVDD.n5552 2.2505
R23768 DVDD.n5555 DVDD.n5554 2.2505
R23769 DVDD.n5557 DVDD.n5556 2.2505
R23770 DVDD.n5559 DVDD.n5558 2.2505
R23771 DVDD.n5561 DVDD.n5560 2.2505
R23772 DVDD.n5659 DVDD.n5658 2.2505
R23773 DVDD.n5657 DVDD.n5562 2.2505
R23774 DVDD.n5656 DVDD.n5655 2.2505
R23775 DVDD.n5654 DVDD.n5653 2.2505
R23776 DVDD.n5567 DVDD.n5564 2.2505
R23777 DVDD.n5612 DVDD.n5611 2.2505
R23778 DVDD.n5649 DVDD.n5648 2.2505
R23779 DVDD.n5647 DVDD.n5646 2.2505
R23780 DVDD.n5645 DVDD.n5644 2.2505
R23781 DVDD.n5643 DVDD.n5642 2.2505
R23782 DVDD.n5641 DVDD.n5640 2.2505
R23783 DVDD.n5639 DVDD.n5638 2.2505
R23784 DVDD.n5637 DVDD.n5636 2.2505
R23785 DVDD.n5635 DVDD.n5634 2.2505
R23786 DVDD.n5631 DVDD.n5572 2.2505
R23787 DVDD.n5630 DVDD.n5629 2.2505
R23788 DVDD.n5628 DVDD.n5627 2.2505
R23789 DVDD.n5626 DVDD.n5625 2.2505
R23790 DVDD.n5624 DVDD.n5623 2.2505
R23791 DVDD.n5622 DVDD.n5621 2.2505
R23792 DVDD.n5620 DVDD.n5619 2.2505
R23793 DVDD.n5618 DVDD.n5617 2.2505
R23794 DVDD.n5616 DVDD.n5615 2.2505
R23795 DVDD.n5614 DVDD.n5613 2.2505
R23796 DVDD.n72 DVDD.n71 2.2505
R23797 DVDD.n5932 DVDD.n5931 2.2505
R23798 DVDD.n5930 DVDD.n5929 2.2505
R23799 DVDD.n5928 DVDD.n73 2.2505
R23800 DVDD.n5927 DVDD.n5926 2.2505
R23801 DVDD.n5925 DVDD.n5924 2.2505
R23802 DVDD.n78 DVDD.n75 2.2505
R23803 DVDD.n86 DVDD.n83 2.2505
R23804 DVDD.n4706 DVDD.n4705 2.2505
R23805 DVDD.n969 DVDD.n948 2.2505
R23806 DVDD.n968 DVDD.n967 2.2505
R23807 DVDD.n965 DVDD.n964 2.2505
R23808 DVDD.n963 DVDD.n962 2.2505
R23809 DVDD.n4704 DVDD.n949 2.2505
R23810 DVDD.n4703 DVDD.n4702 2.2505
R23811 DVDD.n973 DVDD.n970 2.2505
R23812 DVDD.n5485 DVDD.n5484 2.2505
R23813 DVDD.n4646 DVDD.n265 2.2505
R23814 DVDD.n4659 DVDD.n4658 2.2505
R23815 DVDD.n4661 DVDD.n4660 2.2505
R23816 DVDD.n4663 DVDD.n4662 2.2505
R23817 DVDD.n4665 DVDD.n4664 2.2505
R23818 DVDD.n4667 DVDD.n4666 2.2505
R23819 DVDD.n4669 DVDD.n4668 2.2505
R23820 DVDD.n4671 DVDD.n4670 2.2505
R23821 DVDD.n4673 DVDD.n4672 2.2505
R23822 DVDD.n4675 DVDD.n4674 2.2505
R23823 DVDD.n4677 DVDD.n4676 2.2505
R23824 DVDD.n4680 DVDD.n4679 2.2505
R23825 DVDD.n4682 DVDD.n4681 2.2505
R23826 DVDD.n4684 DVDD.n4683 2.2505
R23827 DVDD.n4686 DVDD.n4685 2.2505
R23828 DVDD.n4688 DVDD.n4687 2.2505
R23829 DVDD.n4690 DVDD.n4689 2.2505
R23830 DVDD.n4692 DVDD.n4691 2.2505
R23831 DVDD.n4694 DVDD.n4693 2.2505
R23832 DVDD.n4696 DVDD.n4695 2.2505
R23833 DVDD.n4698 DVDD.n4697 2.2505
R23834 DVDD.n4657 DVDD.n4656 2.2505
R23835 DVDD.n5483 DVDD.n266 2.2505
R23836 DVDD.n5482 DVDD.n5481 2.2505
R23837 DVDD.n5480 DVDD.n5479 2.2505
R23838 DVDD.n5435 DVDD.n294 2.2505
R23839 DVDD.n5434 DVDD.n296 2.2505
R23840 DVDD.n5437 DVDD.n5436 2.2505
R23841 DVDD.n5439 DVDD.n5438 2.2505
R23842 DVDD.n5441 DVDD.n5440 2.2505
R23843 DVDD.n5443 DVDD.n5442 2.2505
R23844 DVDD.n5445 DVDD.n5444 2.2505
R23845 DVDD.n5447 DVDD.n5446 2.2505
R23846 DVDD.n5449 DVDD.n5448 2.2505
R23847 DVDD.n5451 DVDD.n5450 2.2505
R23848 DVDD.n5453 DVDD.n5452 2.2505
R23849 DVDD.n5455 DVDD.n5454 2.2505
R23850 DVDD.n5456 DVDD.n279 2.2505
R23851 DVDD.n5460 DVDD.n5459 2.2505
R23852 DVDD.n5462 DVDD.n5461 2.2505
R23853 DVDD.n5464 DVDD.n5463 2.2505
R23854 DVDD.n5466 DVDD.n5465 2.2505
R23855 DVDD.n5468 DVDD.n5467 2.2505
R23856 DVDD.n5470 DVDD.n5469 2.2505
R23857 DVDD.n5472 DVDD.n5471 2.2505
R23858 DVDD.n319 DVDD.n316 2.2505
R23859 DVDD.n318 DVDD.n317 2.2505
R23860 DVDD.n274 DVDD.n269 2.2505
R23861 DVDD.n5433 DVDD.n5432 2.2505
R23862 DVDD.n5431 DVDD.n320 2.2505
R23863 DVDD.n5427 DVDD.n5426 2.2505
R23864 DVDD.n332 DVDD.n331 2.2505
R23865 DVDD.n330 DVDD.n323 2.2505
R23866 DVDD.n351 DVDD.n341 2.24971
R23867 DVDD.n5916 DVDD.n87 2.24971
R23868 DVDD.n5419 DVDD.n340 2.24971
R23869 DVDD.n106 DVDD.n94 2.24971
R23870 DVDD.n1573 DVDD.n1204 2.24621
R23871 DVDD.n1573 DVDD.n1203 2.24621
R23872 DVDD.n1573 DVDD.n1191 2.24621
R23873 DVDD.n1574 DVDD.n1573 2.24621
R23874 DVDD.n1201 DVDD.n1192 2.24621
R23875 DVDD.n1198 DVDD.n1192 2.24621
R23876 DVDD.n2949 DVDD.n2933 2.24442
R23877 DVDD.n2937 DVDD.n2936 2.24442
R23878 DVDD.n3275 DVDD.n3274 2.24442
R23879 DVDD.n3276 DVDD.n2954 2.24442
R23880 DVDD.n2646 DVDD.n2627 2.24442
R23881 DVDD.n2649 DVDD.n2648 2.24442
R23882 DVDD.n2605 DVDD.n2506 2.24405
R23883 DVDD.n2606 DVDD.n2507 2.24405
R23884 DVDD.n1582 DVDD.n1132 2.24398
R23885 DVDD.n1579 DVDD.n1190 2.24398
R23886 DVDD.n1133 DVDD.n1120 2.24398
R23887 DVDD.n1579 DVDD.n1188 2.24398
R23888 DVDD.n1135 DVDD.n1120 2.24398
R23889 DVDD.n1579 DVDD.n1187 2.24398
R23890 DVDD.n1137 DVDD.n1120 2.24398
R23891 DVDD.n1579 DVDD.n1186 2.24398
R23892 DVDD.n1139 DVDD.n1120 2.24398
R23893 DVDD.n1579 DVDD.n1185 2.24398
R23894 DVDD.n1141 DVDD.n1120 2.24398
R23895 DVDD.n1579 DVDD.n1184 2.24398
R23896 DVDD.n1143 DVDD.n1120 2.24398
R23897 DVDD.n1579 DVDD.n1183 2.24398
R23898 DVDD.n1145 DVDD.n1120 2.24398
R23899 DVDD.n1579 DVDD.n1182 2.24398
R23900 DVDD.n1147 DVDD.n1120 2.24398
R23901 DVDD.n1580 DVDD.n1579 2.24398
R23902 DVDD.n1149 DVDD.n1120 2.24398
R23903 DVDD.n1579 DVDD.n1119 2.24398
R23904 DVDD.n5422 DVDD.n5421 2.24383
R23905 DVDD.n105 DVDD.n104 2.24383
R23906 DVDD.n105 DVDD.n101 2.24383
R23907 DVDD.n350 DVDD.n348 2.24383
R23908 DVDD.n3779 DVDD.n1866 2.24304
R23909 DVDD.n3779 DVDD.n1865 2.24304
R23910 DVDD.n3779 DVDD.n1864 2.24304
R23911 DVDD.n3779 DVDD.n1863 2.24304
R23912 DVDD.n3779 DVDD.n1862 2.24304
R23913 DVDD.n3779 DVDD.n1860 2.24304
R23914 DVDD.n3779 DVDD.n1859 2.24304
R23915 DVDD.n3779 DVDD.n1858 2.24304
R23916 DVDD.n3779 DVDD.n1857 2.24304
R23917 DVDD.n3671 DVDD.n1981 2.24304
R23918 DVDD.n1989 DVDD.n1982 2.24304
R23919 DVDD.n3671 DVDD.n3670 2.24304
R23920 DVDD.n1991 DVDD.n1982 2.24304
R23921 DVDD.n3671 DVDD.n3669 2.24304
R23922 DVDD.n1993 DVDD.n1982 2.24304
R23923 DVDD.n3671 DVDD.n3668 2.24304
R23924 DVDD.n1995 DVDD.n1982 2.24304
R23925 DVDD.n3672 DVDD.n3671 2.24304
R23926 DVDD.n2401 DVDD.n1998 2.24304
R23927 DVDD.n2005 DVDD.n1997 2.24304
R23928 DVDD.n2401 DVDD.n2042 2.24304
R23929 DVDD.n2007 DVDD.n1997 2.24304
R23930 DVDD.n2401 DVDD.n2041 2.24304
R23931 DVDD.n2009 DVDD.n1997 2.24304
R23932 DVDD.n2401 DVDD.n2040 2.24304
R23933 DVDD.n2011 DVDD.n1997 2.24304
R23934 DVDD.n2402 DVDD.n2401 2.24304
R23935 DVDD.n3754 DVDD.n3722 2.24304
R23936 DVDD.n3754 DVDD.n3753 2.24304
R23937 DVDD.n3754 DVDD.n3752 2.24304
R23938 DVDD.n3754 DVDD.n3751 2.24304
R23939 DVDD.n3754 DVDD.n3750 2.24304
R23940 DVDD.n3754 DVDD.n3749 2.24304
R23941 DVDD.n3754 DVDD.n3748 2.24304
R23942 DVDD.n3754 DVDD.n3747 2.24304
R23943 DVDD.n3754 DVDD.n3746 2.24304
R23944 DVDD.n3754 DVDD.n3745 2.24304
R23945 DVDD.n4400 DVDD.n4390 2.24304
R23946 DVDD.n4413 DVDD.n4410 2.24304
R23947 DVDD.n4400 DVDD.n4391 2.24304
R23948 DVDD.n4413 DVDD.n4409 2.24304
R23949 DVDD.n4400 DVDD.n4392 2.24304
R23950 DVDD.n4413 DVDD.n4408 2.24304
R23951 DVDD.n4400 DVDD.n4393 2.24304
R23952 DVDD.n4413 DVDD.n4407 2.24304
R23953 DVDD.n4400 DVDD.n4394 2.24304
R23954 DVDD.n4413 DVDD.n4406 2.24304
R23955 DVDD.n4400 DVDD.n4395 2.24304
R23956 DVDD.n4413 DVDD.n4405 2.24304
R23957 DVDD.n4400 DVDD.n4396 2.24304
R23958 DVDD.n4413 DVDD.n4404 2.24304
R23959 DVDD.n4400 DVDD.n4397 2.24304
R23960 DVDD.n4413 DVDD.n4403 2.24304
R23961 DVDD.n4400 DVDD.n4398 2.24304
R23962 DVDD.n4413 DVDD.n4402 2.24304
R23963 DVDD.n4400 DVDD.n4399 2.24304
R23964 DVDD.n4414 DVDD.n4413 2.24304
R23965 DVDD.n4385 DVDD.n1594 2.24304
R23966 DVDD.n1608 DVDD.n1595 2.24304
R23967 DVDD.n4385 DVDD.n4376 2.24304
R23968 DVDD.n1610 DVDD.n1595 2.24304
R23969 DVDD.n4385 DVDD.n4377 2.24304
R23970 DVDD.n1612 DVDD.n1595 2.24304
R23971 DVDD.n4385 DVDD.n4378 2.24304
R23972 DVDD.n1614 DVDD.n1595 2.24304
R23973 DVDD.n4385 DVDD.n4379 2.24304
R23974 DVDD.n1616 DVDD.n1595 2.24304
R23975 DVDD.n4385 DVDD.n4380 2.24304
R23976 DVDD.n1618 DVDD.n1595 2.24304
R23977 DVDD.n4385 DVDD.n4381 2.24304
R23978 DVDD.n1620 DVDD.n1595 2.24304
R23979 DVDD.n4385 DVDD.n4382 2.24304
R23980 DVDD.n1622 DVDD.n1595 2.24304
R23981 DVDD.n4385 DVDD.n4383 2.24304
R23982 DVDD.n1624 DVDD.n1595 2.24304
R23983 DVDD.n4385 DVDD.n4384 2.24304
R23984 DVDD.n4386 DVDD.n1595 2.24304
R23985 DVDD.n4342 DVDD.n1626 2.24304
R23986 DVDD.n1640 DVDD.n1627 2.24304
R23987 DVDD.n4342 DVDD.n4333 2.24304
R23988 DVDD.n1642 DVDD.n1627 2.24304
R23989 DVDD.n4342 DVDD.n4334 2.24304
R23990 DVDD.n1644 DVDD.n1627 2.24304
R23991 DVDD.n4342 DVDD.n4335 2.24304
R23992 DVDD.n1646 DVDD.n1627 2.24304
R23993 DVDD.n4342 DVDD.n4336 2.24304
R23994 DVDD.n1648 DVDD.n1627 2.24304
R23995 DVDD.n4342 DVDD.n4337 2.24304
R23996 DVDD.n1650 DVDD.n1627 2.24304
R23997 DVDD.n4342 DVDD.n4338 2.24304
R23998 DVDD.n1652 DVDD.n1627 2.24304
R23999 DVDD.n4342 DVDD.n4339 2.24304
R24000 DVDD.n1654 DVDD.n1627 2.24304
R24001 DVDD.n4342 DVDD.n4340 2.24304
R24002 DVDD.n1656 DVDD.n1627 2.24304
R24003 DVDD.n4342 DVDD.n4341 2.24304
R24004 DVDD.n4343 DVDD.n1627 2.24304
R24005 DVDD.n3339 DVDD.n2861 2.24235
R24006 DVDD.n3346 DVDD.n3345 2.24235
R24007 DVDD.n1334 DVDD.n1331 2.24216
R24008 DVDD.n1338 DVDD.n1331 2.24216
R24009 DVDD.n1364 DVDD.n1330 2.24216
R24010 DVDD.n1364 DVDD.n1341 2.24216
R24011 DVDD.n1368 DVDD.n1333 2.24216
R24012 DVDD.n1366 DVDD.n1364 2.24216
R24013 DVDD.n1384 DVDD.n1380 2.23827
R24014 DVDD.n1325 DVDD.n1319 2.23827
R24015 DVDD.n1947 DVDD.n1928 2.20973
R24016 DVDD.n3146 DVDD.n3145 2.1705
R24017 DVDD.n3221 DVDD.n3220 2.1705
R24018 DVDD.n2540 DVDD.t48 2.09436
R24019 DVDD.n2541 DVDD.t52 2.09436
R24020 DVDD.n3145 DVDD.n3144 2.05485
R24021 DVDD.n3220 DVDD.n3219 1.98637
R24022 DVDD.n3151 DVDD.n3150 1.9605
R24023 DVDD.n3115 DVDD.n3113 1.9605
R24024 DVDD.n2520 DVDD.t94 1.95886
R24025 DVDD.n2688 DVDD.n2686 1.93369
R24026 DVDD.n3151 DVDD.n3144 1.92907
R24027 DVDD.n3219 DVDD.n3113 1.86479
R24028 DVDD.n3147 DVDD.n3144 1.8504
R24029 DVDD.n2599 DVDD.n2514 1.81438
R24030 DVDD.n2430 DVDD.t109 1.75468
R24031 DVDD.n2433 DVDD.n2432 1.74881
R24032 DVDD.n3219 DVDD.n3112 1.73846
R24033 DVDD.n2513 DVDD.n2511 1.71988
R24034 DVDD.n1375 DVDD.n1374 1.7146
R24035 DVDD.n3693 DVDD.n3692 1.71444
R24036 DVDD.n1374 DVDD.n1373 1.71412
R24037 DVDD.n2431 DVDD.n2430 1.70307
R24038 DVDD.n4239 DVDD.n1708 1.6972
R24039 DVDD.n4235 DVDD.n4234 1.6972
R24040 DVDD.n4205 DVDD.n4203 1.688
R24041 DVDD.n4138 DVDD.n1713 1.688
R24042 DVDD.n4128 DVDD.n4126 1.688
R24043 DVDD.n4125 DVDD.n1785 1.688
R24044 DVDD.n4124 DVDD.n4123 1.688
R24045 DVDD.n4015 DVDD.n4013 1.688
R24046 DVDD.n3996 DVDD.n3994 1.688
R24047 DVDD.n3932 DVDD.n3931 1.688
R24048 DVDD.n3966 DVDD.n3965 1.688
R24049 DVDD.n3964 DVDD.n3934 1.688
R24050 DVDD.n3963 DVDD.n3962 1.688
R24051 DVDD.n1875 DVDD.n1874 1.688
R24052 DVDD.n1878 DVDD.n1877 1.688
R24053 DVDD.n1869 DVDD.n1868 1.688
R24054 DVDD.n4233 DVDD.n1714 1.688
R24055 DVDD.n1965 DVDD.n1961 1.67609
R24056 DVDD.n1934 DVDD.n1929 1.67609
R24057 DVDD.n1882 DVDD.n1871 1.63826
R24058 DVDD.n1879 DVDD.n1872 1.63826
R24059 DVDD.n4232 DVDD.n1716 1.63826
R24060 DVDD.n4231 DVDD.n1717 1.63826
R24061 DVDD.n4176 DVDD.n1718 1.63826
R24062 DVDD.n4013 DVDD.n1711 1.63109
R24063 DVDD.n3994 DVDD.n1709 1.63109
R24064 DVDD.n3449 DVDD.n2686 1.62357
R24065 DVDD.n4203 DVDD.n4190 1.59264
R24066 DVDD.n2521 DVDD.n2520 1.58954
R24067 DVDD.n1883 DVDD.n1869 1.56519
R24068 DVDD.n2432 DVDD.t110 1.54008
R24069 DVDD.n3066 DVDD.n2991 1.52019
R24070 DVDD.n3347 DVDD.n3344 1.51933
R24071 DVDD.n3343 DVDD.n3342 1.51933
R24072 DVDD.n3673 DVDD.n2405 1.51793
R24073 DVDD.n3190 DVDD.n3134 1.51782
R24074 DVDD.n3778 DVDD.n3721 1.51565
R24075 DVDD.n2651 DVDD.n2491 1.50841
R24076 DVDD.n3044 DVDD.n3040 1.50806
R24077 DVDD.n2151 DVDD.t50 1.50625
R24078 DVDD.n2264 DVDD.t194 1.50625
R24079 DVDD.n2292 DVDD.t169 1.50625
R24080 DVDD.n2085 DVDD.t114 1.50625
R24081 DVDD.n2343 DVDD.t134 1.50625
R24082 DVDD.n2339 DVDD.t68 1.50625
R24083 DVDD.n2367 DVDD.t130 1.50625
R24084 DVDD.n2958 DVDD.n2957 1.50588
R24085 DVDD.n2951 DVDD.n2935 1.50588
R24086 DVDD.n3118 DVDD.n2962 1.50474
R24087 DVDD.n3208 DVDD.n3121 1.50474
R24088 DVDD.n3602 DVDD.n2453 1.50441
R24089 DVDD.n3775 DVDD.n3774 1.50405
R24090 DVDD.n3677 DVDD.n3676 1.50248
R24091 DVDD.n3332 DVDD.n3331 1.5005
R24092 DVDD.n3330 DVDD.n2914 1.5005
R24093 DVDD.n3329 DVDD.n3328 1.5005
R24094 DVDD.n3327 DVDD.n3326 1.5005
R24095 DVDD.n2917 DVDD.n2916 1.5005
R24096 DVDD.n3301 DVDD.n3300 1.5005
R24097 DVDD.n3299 DVDD.n2924 1.5005
R24098 DVDD.n3298 DVDD.n3297 1.5005
R24099 DVDD.n3292 DVDD.n2925 1.5005
R24100 DVDD.n3278 DVDD.n2926 1.5005
R24101 DVDD.n3280 DVDD.n3279 1.5005
R24102 DVDD.n3277 DVDD.n2932 1.5005
R24103 DVDD.n2816 DVDD.n2815 1.5005
R24104 DVDD.n2814 DVDD.n2800 1.5005
R24105 DVDD.n2813 DVDD.n2812 1.5005
R24106 DVDD.n2811 DVDD.n2810 1.5005
R24107 DVDD.n2806 DVDD.n2803 1.5005
R24108 DVDD.n2805 DVDD.n2804 1.5005
R24109 DVDD.n2767 DVDD.n2766 1.5005
R24110 DVDD.n3368 DVDD.n3367 1.5005
R24111 DVDD.n3370 DVDD.n3369 1.5005
R24112 DVDD.n2765 DVDD.n2763 1.5005
R24113 DVDD.n2943 DVDD.n2942 1.5005
R24114 DVDD.n2941 DVDD.n2940 1.5005
R24115 DVDD.n2820 DVDD.n2819 1.5005
R24116 DVDD.n2824 DVDD.n2823 1.5005
R24117 DVDD.n2826 DVDD.n2825 1.5005
R24118 DVDD.n2828 DVDD.n2827 1.5005
R24119 DVDD.n2830 DVDD.n2829 1.5005
R24120 DVDD.n2832 DVDD.n2831 1.5005
R24121 DVDD.n2834 DVDD.n2833 1.5005
R24122 DVDD.n2836 DVDD.n2835 1.5005
R24123 DVDD.n2838 DVDD.n2837 1.5005
R24124 DVDD.n2840 DVDD.n2839 1.5005
R24125 DVDD.n2842 DVDD.n2841 1.5005
R24126 DVDD.n2844 DVDD.n2843 1.5005
R24127 DVDD.n2846 DVDD.n2845 1.5005
R24128 DVDD.n2848 DVDD.n2847 1.5005
R24129 DVDD.n2850 DVDD.n2849 1.5005
R24130 DVDD.n2852 DVDD.n2851 1.5005
R24131 DVDD.n2854 DVDD.n2853 1.5005
R24132 DVDD.n2856 DVDD.n2855 1.5005
R24133 DVDD.n2857 DVDD.n2798 1.5005
R24134 DVDD.n2822 DVDD.n2821 1.5005
R24135 DVDD.n2860 DVDD.n2858 1.5005
R24136 DVDD.n2882 DVDD.n2881 1.5005
R24137 DVDD.n2884 DVDD.n2883 1.5005
R24138 DVDD.n2886 DVDD.n2885 1.5005
R24139 DVDD.n2888 DVDD.n2887 1.5005
R24140 DVDD.n2890 DVDD.n2889 1.5005
R24141 DVDD.n2892 DVDD.n2891 1.5005
R24142 DVDD.n2894 DVDD.n2893 1.5005
R24143 DVDD.n2896 DVDD.n2895 1.5005
R24144 DVDD.n2898 DVDD.n2897 1.5005
R24145 DVDD.n2900 DVDD.n2899 1.5005
R24146 DVDD.n2902 DVDD.n2901 1.5005
R24147 DVDD.n2904 DVDD.n2903 1.5005
R24148 DVDD.n2906 DVDD.n2905 1.5005
R24149 DVDD.n2908 DVDD.n2907 1.5005
R24150 DVDD.n2910 DVDD.n2909 1.5005
R24151 DVDD.n2912 DVDD.n2911 1.5005
R24152 DVDD.n2913 DVDD.n2880 1.5005
R24153 DVDD.n3336 DVDD.n3335 1.5005
R24154 DVDD.n3338 DVDD.n3337 1.5005
R24155 DVDD.n2653 DVDD.n2652 1.5005
R24156 DVDD.n2655 DVDD.n2654 1.5005
R24157 DVDD.n2657 DVDD.n2656 1.5005
R24158 DVDD.n2659 DVDD.n2658 1.5005
R24159 DVDD.n2661 DVDD.n2660 1.5005
R24160 DVDD.n2663 DVDD.n2662 1.5005
R24161 DVDD.n2665 DVDD.n2664 1.5005
R24162 DVDD.n2667 DVDD.n2666 1.5005
R24163 DVDD.n2669 DVDD.n2668 1.5005
R24164 DVDD.n2625 DVDD.n2499 1.5005
R24165 DVDD.n2624 DVDD.n2623 1.5005
R24166 DVDD.n2622 DVDD.n2501 1.5005
R24167 DVDD.n2621 DVDD.n2620 1.5005
R24168 DVDD.n2619 DVDD.n2502 1.5005
R24169 DVDD.n2618 DVDD.n2617 1.5005
R24170 DVDD.n2616 DVDD.n2503 1.5005
R24171 DVDD.n2615 DVDD.n2614 1.5005
R24172 DVDD.n2613 DVDD.n2504 1.5005
R24173 DVDD.n2612 DVDD.n2611 1.5005
R24174 DVDD.n2610 DVDD.n2505 1.5005
R24175 DVDD.n2644 DVDD.n2643 1.5005
R24176 DVDD.n2642 DVDD.n2641 1.5005
R24177 DVDD.n2640 DVDD.n2639 1.5005
R24178 DVDD.n2638 DVDD.n2637 1.5005
R24179 DVDD.n2636 DVDD.n2635 1.5005
R24180 DVDD.n2634 DVDD.n2633 1.5005
R24181 DVDD.n2632 DVDD.n2631 1.5005
R24182 DVDD.n2630 DVDD.n2629 1.5005
R24183 DVDD.n2628 DVDD.n2454 1.5005
R24184 DVDD.n1923 DVDD.n1901 1.5005
R24185 DVDD.n1925 DVDD.n1922 1.5005
R24186 DVDD.n3194 DVDD.n2738 1.5005
R24187 DVDD.n3193 DVDD.n3192 1.5005
R24188 DVDD.n3191 DVDD.n3133 1.5005
R24189 DVDD.n1923 DVDD.n1916 1.5005
R24190 DVDD.n1925 DVDD.n1924 1.5005
R24191 DVDD.n1926 DVDD.n1921 1.5005
R24192 DVDD.n3189 DVDD.n3188 1.5005
R24193 DVDD.n3184 DVDD.n3133 1.5005
R24194 DVDD.n3193 DVDD.n3132 1.5005
R24195 DVDD.n3195 DVDD.n3194 1.5005
R24196 DVDD.n3080 DVDD.n3079 1.5005
R24197 DVDD.n3233 DVDD.n3232 1.5005
R24198 DVDD.n3185 DVDD.n3091 1.5005
R24199 DVDD.n3242 DVDD.n3241 1.5005
R24200 DVDD.n3244 DVDD.n3243 1.5005
R24201 DVDD.n3254 DVDD.n3083 1.5005
R24202 DVDD.n3325 DVDD.n3324 1.5005
R24203 DVDD.n3302 DVDD.n3301 1.5005
R24204 DVDD.n3295 DVDD.n3294 1.5005
R24205 DVDD.n3291 DVDD.n3290 1.5005
R24206 DVDD.n3273 DVDD.n2931 1.5005
R24207 DVDD.n3272 DVDD.n3271 1.5005
R24208 DVDD.n3282 DVDD.n3281 1.5005
R24209 DVDD.n3296 DVDD.n2923 1.5005
R24210 DVDD.n2919 DVDD.n2915 1.5005
R24211 DVDD.n3166 DVDD.n3165 1.5005
R24212 DVDD.n3181 DVDD.n3138 1.5005
R24213 DVDD.n3141 DVDD.n3140 1.5005
R24214 DVDD.n3198 DVDD.n3129 1.5005
R24215 DVDD.n3128 DVDD.n3078 1.5005
R24216 DVDD.n2948 DVDD.n2947 1.5005
R24217 DVDD.n2945 DVDD.n2944 1.5005
R24218 DVDD.n3372 DVDD.n3371 1.5005
R24219 DVDD.n2768 DVDD.n2764 1.5005
R24220 DVDD.n3366 DVDD.n3365 1.5005
R24221 DVDD.n2805 DVDD.n2770 1.5005
R24222 DVDD.n2809 DVDD.n2808 1.5005
R24223 DVDD.n2802 DVDD.n2801 1.5005
R24224 DVDD.n2939 DVDD.n2938 1.5005
R24225 DVDD.n3061 DVDD.n3060 1.5005
R24226 DVDD.n3067 DVDD.n3066 1.5005
R24227 DVDD.n3001 DVDD.n3000 1.5005
R24228 DVDD.n3009 DVDD.n3007 1.5005
R24229 DVDD.n3055 DVDD.n3054 1.5005
R24230 DVDD.n3053 DVDD.n3052 1.5005
R24231 DVDD.n3011 DVDD.n3010 1.5005
R24232 DVDD.n3047 DVDD.n3046 1.5005
R24233 DVDD.n3045 DVDD.n3015 1.5005
R24234 DVDD.n4301 DVDD.n4300 1.5005
R24235 DVDD.n4295 DVDD.n1658 1.5005
R24236 DVDD.n4294 DVDD.n4293 1.5005
R24237 DVDD.n4292 DVDD.n4291 1.5005
R24238 DVDD.n1665 DVDD.n1664 1.5005
R24239 DVDD.n3767 DVDD.n3766 1.5005
R24240 DVDD.n3769 DVDD.n3768 1.5005
R24241 DVDD.n3763 DVDD.n3761 1.5005
R24242 DVDD.n3756 DVDD.n3755 1.5005
R24243 DVDD.n3721 DVDD.n3720 1.5005
R24244 DVDD.n3715 DVDD.n1888 1.5005
R24245 DVDD.n3714 DVDD.n3713 1.5005
R24246 DVDD.n3712 DVDD.n3711 1.5005
R24247 DVDD.n1895 DVDD.n1894 1.5005
R24248 DVDD.n3684 DVDD.n1975 1.5005
R24249 DVDD.n3686 DVDD.n3685 1.5005
R24250 DVDD.n3683 DVDD.n3682 1.5005
R24251 DVDD.n1980 DVDD.n1979 1.5005
R24252 DVDD.n960 DVDD.n942 1.5005
R24253 DVDD.n928 DVDD.n927 1.5005
R24254 DVDD.n940 DVDD.n939 1.5005
R24255 DVDD.n938 DVDD.n937 1.5005
R24256 DVDD.n936 DVDD.n935 1.5005
R24257 DVDD.n934 DVDD.n933 1.5005
R24258 DVDD.n932 DVDD.n931 1.5005
R24259 DVDD.n930 DVDD.n929 1.5005
R24260 DVDD.n951 DVDD.n950 1.5005
R24261 DVDD.n953 DVDD.n952 1.5005
R24262 DVDD.n955 DVDD.n954 1.5005
R24263 DVDD.n957 DVDD.n956 1.5005
R24264 DVDD.n959 DVDD.n958 1.5005
R24265 DVDD.n245 DVDD.n244 1.5005
R24266 DVDD.n258 DVDD.n257 1.5005
R24267 DVDD.n247 DVDD.n246 1.5005
R24268 DVDD.n249 DVDD.n248 1.5005
R24269 DVDD.n251 DVDD.n250 1.5005
R24270 DVDD.n253 DVDD.n252 1.5005
R24271 DVDD.n255 DVDD.n254 1.5005
R24272 DVDD.n5667 DVDD.n5666 1.5005
R24273 DVDD.n5669 DVDD.n5668 1.5005
R24274 DVDD.n5671 DVDD.n5670 1.5005
R24275 DVDD.n5672 DVDD.n242 1.5005
R24276 DVDD.n5674 DVDD.n5673 1.5005
R24277 DVDD.n243 DVDD.n240 1.5005
R24278 DVDD.n2268 DVDD.t78 1.49967
R24279 DVDD.n2269 DVDD.n2268 1.45483
R24280 DVDD.n2075 DVDD.n2074 1.4515
R24281 DVDD.n2338 DVDD.n2094 1.4515
R24282 DVDD.n2141 DVDD.n2140 1.4515
R24283 DVDD.n2263 DVDD.n2160 1.4515
R24284 DVDD.n2368 DVDD.n2367 1.45148
R24285 DVDD.n2086 DVDD.n2085 1.45148
R24286 DVDD.n2339 DVDD.n2063 1.45148
R24287 DVDD.n2344 DVDD.n2343 1.45148
R24288 DVDD.n2293 DVDD.n2292 1.45148
R24289 DVDD.n2152 DVDD.n2151 1.45148
R24290 DVDD.n2264 DVDD.n2127 1.45148
R24291 DVDD.n2403 DVDD 1.39329
R24292 DVDD.n2202 DVDD.n2200 1.3472
R24293 DVDD.n2038 DVDD.n2037 1.33383
R24294 DVDD.n5501 DVDD.n261 1.33314
R24295 DVDD.n2598 DVDD.n2518 1.33037
R24296 DVDD.n4240 DVDD.n4239 1.3141
R24297 DVDD.n4235 DVDD.n1712 1.3141
R24298 DVDD.n2651 DVDD.n2650 1.31276
R24299 DVDD.n1960 DVDD.n1959 1.31159
R24300 DVDD.n2287 DVDD.n2286 1.2972
R24301 DVDD.n2260 DVDD.n2259 1.2972
R24302 DVDD.n2290 DVDD.n2122 1.2972
R24303 DVDD.n2362 DVDD.n2361 1.2972
R24304 DVDD.n2335 DVDD.n2334 1.2972
R24305 DVDD.n2365 DVDD.n2054 1.2972
R24306 DVDD.n2953 DVDD.n2952 1.29474
R24307 DVDD.n1964 DVDD.n1963 1.28124
R24308 DVDD.n1936 DVDD.n1935 1.28123
R24309 DVDD.n1933 DVDD.n1932 1.28123
R24310 DVDD.n4159 DVDD.n1716 1.26907
R24311 DVDD.n1877 DVDD.n1695 1.26907
R24312 DVDD.n3954 DVDD.n3934 1.26907
R24313 DVDD.n3967 DVDD.n3966 1.26907
R24314 DVDD.n3931 DVDD.n3925 1.26907
R24315 DVDD.n4123 DVDD.n4121 1.26907
R24316 DVDD.n4115 DVDD.n1785 1.26907
R24317 DVDD.n4129 DVDD.n4128 1.26907
R24318 DVDD.n1392 DVDD.n1391 1.18293
R24319 DVDD.n1315 DVDD.n1222 1.18293
R24320 DVDD.n5733 DVDD.n5732 1.17409
R24321 DVDD.n5093 DVDD.n5089 1.17409
R24322 DVDD.n598 DVDD.n596 1.17409
R24323 DVDD.n878 DVDD.n877 1.17409
R24324 DVDD.n1060 DVDD.n896 1.17409
R24325 DVDD.n5849 DVDD.n5848 1.17318
R24326 DVDD.n5138 DVDD.n5105 1.17318
R24327 DVDD.n4995 DVDD.n428 1.17318
R24328 DVDD.n759 DVDD.n404 1.17318
R24329 DVDD.n4551 DVDD.n381 1.17318
R24330 DVDD.n3676 DVDD.n3675 1.15295
R24331 DVDD.n2288 DVDD.n2287 1.14595
R24332 DVDD.n2363 DVDD.n2362 1.14595
R24333 DVDD.n3699 DVDD.n3698 1.1282
R24334 DVDD.n2035 DVDD.n2034 1.1255
R24335 DVDD.n2037 DVDD.n2036 1.1255
R24336 DVDD.n2031 DVDD.n2030 1.1255
R24337 DVDD.n2033 DVDD.n2032 1.1255
R24338 DVDD.n2027 DVDD.n2026 1.1255
R24339 DVDD.n2029 DVDD.n2028 1.1255
R24340 DVDD.n2023 DVDD.n2022 1.1255
R24341 DVDD.n2025 DVDD.n2024 1.1255
R24342 DVDD.n2019 DVDD.n2018 1.1255
R24343 DVDD.n2021 DVDD.n2020 1.1255
R24344 DVDD.n2015 DVDD.n2014 1.1255
R24345 DVDD.n2017 DVDD.n2016 1.1255
R24346 DVDD.n2202 DVDD.n2201 1.1255
R24347 DVDD.n2601 DVDD.n2600 1.1255
R24348 DVDD.n1964 DVDD.n1962 1.11867
R24349 DVDD.n1959 DVDD.n1958 1.11867
R24350 DVDD.n1936 DVDD.n1930 1.11867
R24351 DVDD.n1932 DVDD.n1931 1.11867
R24352 DVDD.n3451 DVDD.n3450 1.08635
R24353 DVDD.n2266 DVDD.n2261 1.0505
R24354 DVDD.n2289 DVDD.n2124 1.0505
R24355 DVDD.n2341 DVDD.n2336 1.0505
R24356 DVDD.n2364 DVDD.n2060 1.0505
R24357 DVDD.n3697 DVDD.n3696 0.969731
R24358 DVDD.n1578 DVDD.n1577 0.969652
R24359 DVDD.n2604 DVDD.n2603 0.968342
R24360 DVDD.n2514 DVDD.t11 0.958395
R24361 DVDD.n2514 DVDD.t24 0.958395
R24362 DVDD.n4300 DVDD.n4299 0.91193
R24363 DVDD.n2515 DVDD.t192 0.9105
R24364 DVDD.n2515 DVDD.t13 0.9105
R24365 DVDD.n3720 DVDD.n3719 0.910366
R24366 DVDD.n3679 DVDD.n3677 0.908384
R24367 DVDD.n3774 DVDD.n3773 0.908384
R24368 DVDD.n4139 DVDD.n4138 0.904312
R24369 DVDD.n3962 DVDD.n3961 0.904312
R24370 DVDD.n1874 DVDD.n1873 0.904312
R24371 DVDD.n4149 DVDD.n1714 0.904312
R24372 DVDD.n3175 DVDD.n3116 0.9005
R24373 DVDD.n3223 DVDD.n3222 0.9005
R24374 DVDD.n3216 DVDD.n3087 0.9005
R24375 DVDD.n3172 DVDD.n3109 0.9005
R24376 DVDD.n3678 DVDD.n1976 0.9005
R24377 DVDD.n3688 DVDD.n1977 0.9005
R24378 DVDD.n3689 DVDD.n1910 0.9005
R24379 DVDD.n3709 DVDD.n3708 0.9005
R24380 DVDD.n1892 DVDD.n1891 0.9005
R24381 DVDD.n3718 DVDD.n3717 0.9005
R24382 DVDD.n3681 DVDD.n3680 0.9005
R24383 DVDD.n1978 DVDD.n1976 0.9005
R24384 DVDD.n3688 DVDD.n3687 0.9005
R24385 DVDD.n3690 DVDD.n3689 0.9005
R24386 DVDD.n3710 DVDD.n3709 0.9005
R24387 DVDD.n1893 DVDD.n1892 0.9005
R24388 DVDD.n3717 DVDD.n3716 0.9005
R24389 DVDD.n1890 DVDD.n1889 0.9005
R24390 DVDD.n3772 DVDD.n3771 0.9005
R24391 DVDD.n3759 DVDD.n3758 0.9005
R24392 DVDD.n3764 DVDD.n1667 0.9005
R24393 DVDD.n4289 DVDD.n4288 0.9005
R24394 DVDD.n1662 DVDD.n1661 0.9005
R24395 DVDD.n4298 DVDD.n4297 0.9005
R24396 DVDD.n3760 DVDD.n3757 0.9005
R24397 DVDD.n3771 DVDD.n3770 0.9005
R24398 DVDD.n3762 DVDD.n3759 0.9005
R24399 DVDD.n3765 DVDD.n3764 0.9005
R24400 DVDD.n4290 DVDD.n4289 0.9005
R24401 DVDD.n1663 DVDD.n1662 0.9005
R24402 DVDD.n4297 DVDD.n4296 0.9005
R24403 DVDD.n1660 DVDD.n1659 0.9005
R24404 DVDD.n2263 DVDD.n2262 0.899883
R24405 DVDD.n2140 DVDD.n2139 0.899883
R24406 DVDD.n2338 DVDD.n2337 0.899883
R24407 DVDD.n2074 DVDD.n2073 0.899883
R24408 DVDD.n1375 DVDD.n1370 0.886656
R24409 DVDD.n2600 DVDD.n2513 0.875562
R24410 DVDD.n1373 DVDD.n1371 0.87516
R24411 DVDD.n2540 DVDD.n2539 0.8555
R24412 DVDD.n5664 DVDD.n259 0.82049
R24413 DVDD.n5490 DVDD.n263 0.814302
R24414 DVDD.n1928 DVDD.n1927 0.797897
R24415 DVDD.n1868 DVDD.n1852 0.773058
R24416 DVDD.n1871 DVDD.n1690 0.773058
R24417 DVDD.n1872 DVDD.n1691 0.773058
R24418 DVDD.n3997 DVDD.n3996 0.773058
R24419 DVDD.n4016 DVDD.n4015 0.773058
R24420 DVDD.n1769 DVDD.n1717 0.773058
R24421 DVDD.n4177 DVDD.n4176 0.773058
R24422 DVDD.n4206 DVDD.n4205 0.773058
R24423 DVDD.n2014 DVDD.n2013 0.771833
R24424 DVDD.n1967 DVDD.n1966 0.769687
R24425 DVDD.n3191 DVDD.n3190 0.769684
R24426 DVDD.n3445 DVDD.n3444 0.755277
R24427 DVDD.n2818 DVDD.n2817 0.751
R24428 DVDD.n3334 DVDD.n3333 0.751
R24429 DVDD.n2719 DVDD.n2718 0.7505
R24430 DVDD.n2718 DVDD.n2717 0.7505
R24431 DVDD.n3231 DVDD.n3106 0.735937
R24432 DVDD.n3227 DVDD.n3226 0.735937
R24433 DVDD.n3171 DVDD.n3170 0.735937
R24434 DVDD.n3167 DVDD.n3108 0.735937
R24435 DVDD.n2511 DVDD.n2453 0.734685
R24436 DVDD.n2267 DVDD.n2260 0.714509
R24437 DVDD.n2291 DVDD.n2290 0.714509
R24438 DVDD.n2342 DVDD.n2335 0.714509
R24439 DVDD.n2366 DVDD.n2365 0.714509
R24440 DVDD.n2582 DVDD.n2542 0.711129
R24441 DVDD.n2580 DVDD.n2564 0.711129
R24442 DVDD.n2575 DVDD.n2574 0.7005
R24443 DVDD.n2576 DVDD.n2557 0.7005
R24444 DVDD.n2577 DVDD.n2560 0.7005
R24445 DVDD.n2578 DVDD.n2556 0.7005
R24446 DVDD.n2580 DVDD.n2579 0.7005
R24447 DVDD.n2564 DVDD.n2547 0.7005
R24448 DVDD.n2583 DVDD.n2582 0.7005
R24449 DVDD.n2584 DVDD.n2542 0.7005
R24450 DVDD.n2589 DVDD.n2588 0.7005
R24451 DVDD.n2591 DVDD.n2590 0.7005
R24452 DVDD.n2538 DVDD.n2524 0.7005
R24453 DVDD.n2594 DVDD.n2593 0.7005
R24454 DVDD.n2523 DVDD.n2522 0.668882
R24455 DVDD.n2518 DVDD.n2516 0.666798
R24456 DVDD.n3695 DVDD.n3693 0.646382
R24457 DVDD.n2523 DVDD.n2513 0.645825
R24458 DVDD.n4202 DVDD.n4200 0.634998
R24459 DVDD.n1947 DVDD.n1946 0.634532
R24460 DVDD.n1379 DVDD.n1325 0.634344
R24461 DVDD.n1380 DVDD.n1379 0.632309
R24462 DVDD.n2262 DVDD.t63 0.607167
R24463 DVDD.n2262 DVDD.t60 0.607167
R24464 DVDD.n2139 DVDD.t147 0.607167
R24465 DVDD.n2139 DVDD.t56 0.607167
R24466 DVDD.n2337 DVDD.t163 0.607167
R24467 DVDD.n2337 DVDD.t167 0.607167
R24468 DVDD.n2073 DVDD.t173 0.607167
R24469 DVDD.n2073 DVDD.t112 0.607167
R24470 DVDD.n3692 DVDD.t16 0.607167
R24471 DVDD.n3692 DVDD.t161 0.607167
R24472 DVDD.n2602 DVDD.n2601 0.594875
R24473 DVDD.n4233 DVDD.n4232 0.590794
R24474 DVDD.n4232 DVDD.n4231 0.578395
R24475 DVDD.n2531 DVDD.n2519 0.573227
R24476 DVDD.n2595 DVDD.n2519 0.573227
R24477 DVDD.n2203 DVDD.n2202 0.571463
R24478 DVDD.n2541 DVDD 0.565368
R24479 DVDD.n3204 DVDD.n3121 0.563
R24480 DVDD.n3213 DVDD.n3212 0.563
R24481 DVDD.n3119 DVDD.n3118 0.563
R24482 DVDD.n3120 DVDD.n3117 0.563
R24483 DVDD.n3446 DVDD.n3445 0.563
R24484 DVDD.n2287 DVDD.n2125 0.557079
R24485 DVDD.n2362 DVDD.n2061 0.557079
R24486 DVDD.n1879 DVDD.n1878 0.552481
R24487 DVDD.n2267 DVDD.n2266 0.545794
R24488 DVDD.n2291 DVDD.n2124 0.545794
R24489 DVDD.n2342 DVDD.n2341 0.545794
R24490 DVDD.n2366 DVDD.n2060 0.545794
R24491 DVDD.n4126 DVDD.n1713 0.545794
R24492 DVDD.n4126 DVDD.n4125 0.545794
R24493 DVDD.n3965 DVDD.n3964 0.545794
R24494 DVDD.n3964 DVDD.n3963 0.545794
R24495 DVDD.n1878 DVDD.n1875 0.545794
R24496 DVDD.n3222 DVDD.n3106 0.527932
R24497 DVDD.n3172 DVDD.n3171 0.527932
R24498 DVDD.n1927 DVDD.n1922 0.525612
R24499 DVDD.n3698 DVDD 0.471676
R24500 DVDD.n2268 DVDD.n2267 0.463605
R24501 DVDD.n2401 DVDD.n2039 0.463585
R24502 DVDD.n3665 DVDD.n1982 0.463585
R24503 DVDD.n3679 DVDD.n3678 0.459655
R24504 DVDD.n3719 DVDD.n3718 0.459655
R24505 DVDD.n3773 DVDD.n3772 0.459655
R24506 DVDD.n4299 DVDD.n4298 0.459655
R24507 DVDD.n2151 DVDD.n2150 0.457026
R24508 DVDD.n2265 DVDD.n2264 0.457026
R24509 DVDD.n2292 DVDD.n2291 0.457026
R24510 DVDD.n2085 DVDD.n2084 0.457026
R24511 DVDD.n2343 DVDD.n2342 0.457026
R24512 DVDD.n2340 DVDD.n2339 0.457026
R24513 DVDD.n2367 DVDD.n2366 0.457026
R24514 DVDD.n2266 DVDD.n2263 0.457011
R24515 DVDD.n2140 DVDD.n2124 0.457011
R24516 DVDD.n2341 DVDD.n2338 0.457011
R24517 DVDD.n2074 DVDD.n2060 0.457011
R24518 DVDD.n1965 DVDD 0.455237
R24519 DVDD DVDD.n1929 0.455237
R24520 DVDD.n2197 DVDD.n2196 0.4505
R24521 DVDD.n2195 DVDD.n2194 0.4505
R24522 DVDD.n2206 DVDD.n2205 0.4505
R24523 DVDD.n2207 DVDD.n2193 0.4505
R24524 DVDD.n2209 DVDD.n2208 0.4505
R24525 DVDD.n2191 DVDD.n2190 0.4505
R24526 DVDD.n2214 DVDD.n2213 0.4505
R24527 DVDD.n2215 DVDD.n2189 0.4505
R24528 DVDD.n2217 DVDD.n2216 0.4505
R24529 DVDD.n2187 DVDD.n2186 0.4505
R24530 DVDD.n2222 DVDD.n2221 0.4505
R24531 DVDD.n2223 DVDD.n2185 0.4505
R24532 DVDD.n2225 DVDD.n2224 0.4505
R24533 DVDD.n2183 DVDD.n2182 0.4505
R24534 DVDD.n2230 DVDD.n2229 0.4505
R24535 DVDD.n2231 DVDD.n2181 0.4505
R24536 DVDD.n2233 DVDD.n2232 0.4505
R24537 DVDD.n2179 DVDD.n2178 0.4505
R24538 DVDD.n2238 DVDD.n2237 0.4505
R24539 DVDD.n2239 DVDD.n2177 0.4505
R24540 DVDD.n2241 DVDD.n2240 0.4505
R24541 DVDD.n2175 DVDD.n2174 0.4505
R24542 DVDD.n2246 DVDD.n2245 0.4505
R24543 DVDD.n2247 DVDD.n2173 0.4505
R24544 DVDD.n2249 DVDD.n2248 0.4505
R24545 DVDD.n2171 DVDD.n2170 0.4505
R24546 DVDD.n2254 DVDD.n2253 0.4505
R24547 DVDD.n2255 DVDD.n2168 0.4505
R24548 DVDD.n2257 DVDD.n2256 0.4505
R24549 DVDD.n2169 DVDD.n2167 0.4505
R24550 DVDD.n2163 DVDD.n2162 0.4505
R24551 DVDD.n2273 DVDD.n2272 0.4505
R24552 DVDD.n2274 DVDD.n2161 0.4505
R24553 DVDD.n2276 DVDD.n2275 0.4505
R24554 DVDD.n2158 DVDD.n2157 0.4505
R24555 DVDD.n2281 DVDD.n2280 0.4505
R24556 DVDD.n2282 DVDD.n2129 0.4505
R24557 DVDD.n2284 DVDD.n2283 0.4505
R24558 DVDD.n2156 DVDD.n2128 0.4505
R24559 DVDD.n2155 DVDD.n2154 0.4505
R24560 DVDD.n2131 DVDD.n2130 0.4505
R24561 DVDD.n2147 DVDD.n2146 0.4505
R24562 DVDD.n2145 DVDD.n2133 0.4505
R24563 DVDD.n2144 DVDD.n2143 0.4505
R24564 DVDD.n2137 DVDD.n2134 0.4505
R24565 DVDD.n2136 DVDD.n2135 0.4505
R24566 DVDD.n2121 DVDD.n2120 0.4505
R24567 DVDD.n2398 DVDD.n2397 0.4505
R24568 DVDD.n2396 DVDD.n2043 0.4505
R24569 DVDD.n2395 DVDD.n2394 0.4505
R24570 DVDD.n2045 DVDD.n2044 0.4505
R24571 DVDD.n2390 DVDD.n2389 0.4505
R24572 DVDD.n2388 DVDD.n2047 0.4505
R24573 DVDD.n2387 DVDD.n2386 0.4505
R24574 DVDD.n2049 DVDD.n2048 0.4505
R24575 DVDD.n2382 DVDD.n2381 0.4505
R24576 DVDD.n2380 DVDD.n2051 0.4505
R24577 DVDD.n2379 DVDD.n2378 0.4505
R24578 DVDD.n2053 DVDD.n2052 0.4505
R24579 DVDD.n2374 DVDD.n2373 0.4505
R24580 DVDD.n2372 DVDD.n2055 0.4505
R24581 DVDD.n2371 DVDD.n2370 0.4505
R24582 DVDD.n2057 DVDD.n2056 0.4505
R24583 DVDD.n2071 DVDD.n2070 0.4505
R24584 DVDD.n2078 DVDD.n2077 0.4505
R24585 DVDD.n2079 DVDD.n2069 0.4505
R24586 DVDD.n2081 DVDD.n2080 0.4505
R24587 DVDD.n2067 DVDD.n2066 0.4505
R24588 DVDD.n2089 DVDD.n2088 0.4505
R24589 DVDD.n2090 DVDD.n2064 0.4505
R24590 DVDD.n2359 DVDD.n2358 0.4505
R24591 DVDD.n2357 DVDD.n2065 0.4505
R24592 DVDD.n2356 DVDD.n2355 0.4505
R24593 DVDD.n2092 DVDD.n2091 0.4505
R24594 DVDD.n2351 DVDD.n2350 0.4505
R24595 DVDD.n2349 DVDD.n2095 0.4505
R24596 DVDD.n2348 DVDD.n2347 0.4505
R24597 DVDD.n2097 DVDD.n2096 0.4505
R24598 DVDD.n2103 DVDD.n2101 0.4505
R24599 DVDD.n2332 DVDD.n2331 0.4505
R24600 DVDD.n2330 DVDD.n2102 0.4505
R24601 DVDD.n2329 DVDD.n2328 0.4505
R24602 DVDD.n2105 DVDD.n2104 0.4505
R24603 DVDD.n2324 DVDD.n2323 0.4505
R24604 DVDD.n2322 DVDD.n2107 0.4505
R24605 DVDD.n2321 DVDD.n2320 0.4505
R24606 DVDD.n2109 DVDD.n2108 0.4505
R24607 DVDD.n2316 DVDD.n2315 0.4505
R24608 DVDD.n2314 DVDD.n2111 0.4505
R24609 DVDD.n2313 DVDD.n2312 0.4505
R24610 DVDD.n2113 DVDD.n2112 0.4505
R24611 DVDD.n2308 DVDD.n2307 0.4505
R24612 DVDD.n2306 DVDD.n2115 0.4505
R24613 DVDD.n2305 DVDD.n2304 0.4505
R24614 DVDD.n2117 DVDD.n2116 0.4505
R24615 DVDD.n2300 DVDD.n2299 0.4505
R24616 DVDD.n2298 DVDD.n2119 0.4505
R24617 DVDD.n2297 DVDD.n2296 0.4505
R24618 DVDD.n2205 DVDD.n2204 0.4505
R24619 DVDD.n2400 DVDD.n2399 0.4505
R24620 DVDD.n2398 DVDD.n1999 0.4505
R24621 DVDD.n2043 DVDD.n2004 0.4505
R24622 DVDD.n2394 DVDD.n2393 0.4505
R24623 DVDD.n2392 DVDD.n2045 0.4505
R24624 DVDD.n2391 DVDD.n2390 0.4505
R24625 DVDD.n2047 DVDD.n2046 0.4505
R24626 DVDD.n2386 DVDD.n2385 0.4505
R24627 DVDD.n2384 DVDD.n2049 0.4505
R24628 DVDD.n2383 DVDD.n2382 0.4505
R24629 DVDD.n2051 DVDD.n2050 0.4505
R24630 DVDD.n2378 DVDD.n2377 0.4505
R24631 DVDD.n2376 DVDD.n2053 0.4505
R24632 DVDD.n2375 DVDD.n2374 0.4505
R24633 DVDD.n2058 DVDD.n2055 0.4505
R24634 DVDD.n2370 DVDD.n2369 0.4505
R24635 DVDD.n2059 DVDD.n2057 0.4505
R24636 DVDD.n2072 DVDD.n2071 0.4505
R24637 DVDD.n2077 DVDD.n2076 0.4505
R24638 DVDD.n2069 DVDD.n2068 0.4505
R24639 DVDD.n2082 DVDD.n2081 0.4505
R24640 DVDD.n2083 DVDD.n2067 0.4505
R24641 DVDD.n2088 DVDD.n2087 0.4505
R24642 DVDD.n2064 DVDD.n2062 0.4505
R24643 DVDD.n2360 DVDD.n2359 0.4505
R24644 DVDD.n2093 DVDD.n2065 0.4505
R24645 DVDD.n2355 DVDD.n2354 0.4505
R24646 DVDD.n2353 DVDD.n2092 0.4505
R24647 DVDD.n2352 DVDD.n2351 0.4505
R24648 DVDD.n2098 DVDD.n2095 0.4505
R24649 DVDD.n2347 DVDD.n2346 0.4505
R24650 DVDD.n2345 DVDD.n2097 0.4505
R24651 DVDD.n2101 DVDD.n2099 0.4505
R24652 DVDD.n2333 DVDD.n2332 0.4505
R24653 DVDD.n2102 DVDD.n2100 0.4505
R24654 DVDD.n2328 DVDD.n2327 0.4505
R24655 DVDD.n2326 DVDD.n2105 0.4505
R24656 DVDD.n2325 DVDD.n2324 0.4505
R24657 DVDD.n2107 DVDD.n2106 0.4505
R24658 DVDD.n2320 DVDD.n2319 0.4505
R24659 DVDD.n2318 DVDD.n2109 0.4505
R24660 DVDD.n2317 DVDD.n2316 0.4505
R24661 DVDD.n2111 DVDD.n2110 0.4505
R24662 DVDD.n2312 DVDD.n2311 0.4505
R24663 DVDD.n2310 DVDD.n2113 0.4505
R24664 DVDD.n2309 DVDD.n2308 0.4505
R24665 DVDD.n2115 DVDD.n2114 0.4505
R24666 DVDD.n2304 DVDD.n2303 0.4505
R24667 DVDD.n2302 DVDD.n2117 0.4505
R24668 DVDD.n2301 DVDD.n2300 0.4505
R24669 DVDD.n2119 DVDD.n2118 0.4505
R24670 DVDD.n2294 DVDD.n2121 0.4505
R24671 DVDD.n2136 DVDD.n2123 0.4505
R24672 DVDD.n2138 DVDD.n2137 0.4505
R24673 DVDD.n2143 DVDD.n2142 0.4505
R24674 DVDD.n2133 DVDD.n2132 0.4505
R24675 DVDD.n2148 DVDD.n2147 0.4505
R24676 DVDD.n2149 DVDD.n2131 0.4505
R24677 DVDD.n2154 DVDD.n2153 0.4505
R24678 DVDD.n2128 DVDD.n2126 0.4505
R24679 DVDD.n2285 DVDD.n2284 0.4505
R24680 DVDD.n2159 DVDD.n2129 0.4505
R24681 DVDD.n2280 DVDD.n2279 0.4505
R24682 DVDD.n2278 DVDD.n2158 0.4505
R24683 DVDD.n2277 DVDD.n2276 0.4505
R24684 DVDD.n2164 DVDD.n2161 0.4505
R24685 DVDD.n2272 DVDD.n2271 0.4505
R24686 DVDD.n2270 DVDD.n2163 0.4505
R24687 DVDD.n2167 DVDD.n2165 0.4505
R24688 DVDD.n2258 DVDD.n2257 0.4505
R24689 DVDD.n2168 DVDD.n2166 0.4505
R24690 DVDD.n2253 DVDD.n2252 0.4505
R24691 DVDD.n2251 DVDD.n2171 0.4505
R24692 DVDD.n2250 DVDD.n2249 0.4505
R24693 DVDD.n2173 DVDD.n2172 0.4505
R24694 DVDD.n2245 DVDD.n2244 0.4505
R24695 DVDD.n2243 DVDD.n2175 0.4505
R24696 DVDD.n2242 DVDD.n2241 0.4505
R24697 DVDD.n2177 DVDD.n2176 0.4505
R24698 DVDD.n2237 DVDD.n2236 0.4505
R24699 DVDD.n2235 DVDD.n2179 0.4505
R24700 DVDD.n2234 DVDD.n2233 0.4505
R24701 DVDD.n2181 DVDD.n2180 0.4505
R24702 DVDD.n2229 DVDD.n2228 0.4505
R24703 DVDD.n2227 DVDD.n2183 0.4505
R24704 DVDD.n2226 DVDD.n2225 0.4505
R24705 DVDD.n2185 DVDD.n2184 0.4505
R24706 DVDD.n2221 DVDD.n2220 0.4505
R24707 DVDD.n2219 DVDD.n2187 0.4505
R24708 DVDD.n2218 DVDD.n2217 0.4505
R24709 DVDD.n2189 DVDD.n2188 0.4505
R24710 DVDD.n2213 DVDD.n2212 0.4505
R24711 DVDD.n2211 DVDD.n2191 0.4505
R24712 DVDD.n2210 DVDD.n2209 0.4505
R24713 DVDD.n2193 DVDD.n2192 0.4505
R24714 DVDD.n2199 DVDD.n2195 0.4505
R24715 DVDD.n2296 DVDD.n2295 0.4505
R24716 DVDD.n3472 DVDD.n3471 0.4505
R24717 DVDD.n3473 DVDD.n3469 0.4505
R24718 DVDD.n3475 DVDD.n3474 0.4505
R24719 DVDD.n3467 DVDD.n3466 0.4505
R24720 DVDD.n3480 DVDD.n3479 0.4505
R24721 DVDD.n3481 DVDD.n3465 0.4505
R24722 DVDD.n3483 DVDD.n3482 0.4505
R24723 DVDD.n3463 DVDD.n3462 0.4505
R24724 DVDD.n3488 DVDD.n3487 0.4505
R24725 DVDD.n3489 DVDD.n3461 0.4505
R24726 DVDD.n3491 DVDD.n3490 0.4505
R24727 DVDD.n3459 DVDD.n3458 0.4505
R24728 DVDD.n3496 DVDD.n3495 0.4505
R24729 DVDD.n3497 DVDD.n3457 0.4505
R24730 DVDD.n3499 DVDD.n3498 0.4505
R24731 DVDD.n3455 DVDD.n3454 0.4505
R24732 DVDD.n3504 DVDD.n3503 0.4505
R24733 DVDD.n3505 DVDD.n3453 0.4505
R24734 DVDD.n3507 DVDD.n3506 0.4505
R24735 DVDD.n2684 DVDD.n2683 0.4505
R24736 DVDD.n3512 DVDD.n3511 0.4505
R24737 DVDD.n3513 DVDD.n2682 0.4505
R24738 DVDD.n3515 DVDD.n3514 0.4505
R24739 DVDD.n2680 DVDD.n2679 0.4505
R24740 DVDD.n3520 DVDD.n3519 0.4505
R24741 DVDD.n3521 DVDD.n2673 0.4505
R24742 DVDD.n3523 DVDD.n3522 0.4505
R24743 DVDD.n2678 DVDD.n2671 0.4505
R24744 DVDD.n2677 DVDD.n2676 0.4505
R24745 DVDD.n2675 DVDD.n2674 0.4505
R24746 DVDD.n2490 DVDD.n2489 0.4505
R24747 DVDD.n3532 DVDD.n3531 0.4505
R24748 DVDD.n3533 DVDD.n2488 0.4505
R24749 DVDD.n3535 DVDD.n3534 0.4505
R24750 DVDD.n2486 DVDD.n2485 0.4505
R24751 DVDD.n3540 DVDD.n3539 0.4505
R24752 DVDD.n3541 DVDD.n2484 0.4505
R24753 DVDD.n3543 DVDD.n3542 0.4505
R24754 DVDD.n2482 DVDD.n2481 0.4505
R24755 DVDD.n3548 DVDD.n3547 0.4505
R24756 DVDD.n3549 DVDD.n2480 0.4505
R24757 DVDD.n3551 DVDD.n3550 0.4505
R24758 DVDD.n2478 DVDD.n2477 0.4505
R24759 DVDD.n3556 DVDD.n3555 0.4505
R24760 DVDD.n3557 DVDD.n2476 0.4505
R24761 DVDD.n3559 DVDD.n3558 0.4505
R24762 DVDD.n2474 DVDD.n2473 0.4505
R24763 DVDD.n3564 DVDD.n3563 0.4505
R24764 DVDD.n3565 DVDD.n2472 0.4505
R24765 DVDD.n3567 DVDD.n3566 0.4505
R24766 DVDD.n2470 DVDD.n2469 0.4505
R24767 DVDD.n3572 DVDD.n3571 0.4505
R24768 DVDD.n3573 DVDD.n2468 0.4505
R24769 DVDD.n3575 DVDD.n3574 0.4505
R24770 DVDD.n2466 DVDD.n2465 0.4505
R24771 DVDD.n3580 DVDD.n3579 0.4505
R24772 DVDD.n3581 DVDD.n2464 0.4505
R24773 DVDD.n3583 DVDD.n3582 0.4505
R24774 DVDD.n2462 DVDD.n2461 0.4505
R24775 DVDD.n3588 DVDD.n3587 0.4505
R24776 DVDD.n3589 DVDD.n2460 0.4505
R24777 DVDD.n3591 DVDD.n3590 0.4505
R24778 DVDD.n2458 DVDD.n2457 0.4505
R24779 DVDD.n3596 DVDD.n3595 0.4505
R24780 DVDD.n3597 DVDD.n2456 0.4505
R24781 DVDD.n3599 DVDD.n3598 0.4505
R24782 DVDD.n2441 DVDD.n2440 0.4505
R24783 DVDD.n3606 DVDD.n3605 0.4505
R24784 DVDD.n3607 DVDD.n2439 0.4505
R24785 DVDD.n3609 DVDD.n3608 0.4505
R24786 DVDD.n2436 DVDD.n2435 0.4505
R24787 DVDD.n3614 DVDD.n3613 0.4505
R24788 DVDD.n3664 DVDD.n2406 0.4505
R24789 DVDD.n3663 DVDD.n3662 0.4505
R24790 DVDD.n3661 DVDD.n2407 0.4505
R24791 DVDD.n2411 DVDD.n2408 0.4505
R24792 DVDD.n3657 DVDD.n3656 0.4505
R24793 DVDD.n3655 DVDD.n2410 0.4505
R24794 DVDD.n3654 DVDD.n3653 0.4505
R24795 DVDD.n2413 DVDD.n2412 0.4505
R24796 DVDD.n3649 DVDD.n3648 0.4505
R24797 DVDD.n3647 DVDD.n2415 0.4505
R24798 DVDD.n3646 DVDD.n3645 0.4505
R24799 DVDD.n2417 DVDD.n2416 0.4505
R24800 DVDD.n3641 DVDD.n3640 0.4505
R24801 DVDD.n3639 DVDD.n2419 0.4505
R24802 DVDD.n3638 DVDD.n3637 0.4505
R24803 DVDD.n2421 DVDD.n2420 0.4505
R24804 DVDD.n3633 DVDD.n3632 0.4505
R24805 DVDD.n3631 DVDD.n2423 0.4505
R24806 DVDD.n3630 DVDD.n3629 0.4505
R24807 DVDD.n2425 DVDD.n2424 0.4505
R24808 DVDD.n3625 DVDD.n3624 0.4505
R24809 DVDD.n3623 DVDD.n2427 0.4505
R24810 DVDD.n3622 DVDD.n3621 0.4505
R24811 DVDD.n2429 DVDD.n2428 0.4505
R24812 DVDD.n3617 DVDD.n3616 0.4505
R24813 DVDD.n3615 DVDD.n2434 0.4505
R24814 DVDD.n3525 DVDD.n2671 0.4505
R24815 DVDD.n2676 DVDD.n2670 0.4505
R24816 DVDD.n3524 DVDD.n3523 0.4505
R24817 DVDD.n2673 DVDD.n2672 0.4505
R24818 DVDD.n3519 DVDD.n3518 0.4505
R24819 DVDD.n3517 DVDD.n2680 0.4505
R24820 DVDD.n3516 DVDD.n3515 0.4505
R24821 DVDD.n2682 DVDD.n2681 0.4505
R24822 DVDD.n3511 DVDD.n3510 0.4505
R24823 DVDD.n3509 DVDD.n2684 0.4505
R24824 DVDD.n3508 DVDD.n3507 0.4505
R24825 DVDD.n3453 DVDD.n3452 0.4505
R24826 DVDD.n3503 DVDD.n3502 0.4505
R24827 DVDD.n3501 DVDD.n3455 0.4505
R24828 DVDD.n3500 DVDD.n3499 0.4505
R24829 DVDD.n3457 DVDD.n3456 0.4505
R24830 DVDD.n3495 DVDD.n3494 0.4505
R24831 DVDD.n3493 DVDD.n3459 0.4505
R24832 DVDD.n3492 DVDD.n3491 0.4505
R24833 DVDD.n3461 DVDD.n3460 0.4505
R24834 DVDD.n3487 DVDD.n3486 0.4505
R24835 DVDD.n3485 DVDD.n3463 0.4505
R24836 DVDD.n3484 DVDD.n3483 0.4505
R24837 DVDD.n3465 DVDD.n3464 0.4505
R24838 DVDD.n3479 DVDD.n3478 0.4505
R24839 DVDD.n3477 DVDD.n3467 0.4505
R24840 DVDD.n3476 DVDD.n3475 0.4505
R24841 DVDD.n3469 DVDD.n3468 0.4505
R24842 DVDD.n2675 DVDD.n2495 0.4505
R24843 DVDD.n3529 DVDD.n2490 0.4505
R24844 DVDD.n3531 DVDD.n3530 0.4505
R24845 DVDD.n2488 DVDD.n2487 0.4505
R24846 DVDD.n3536 DVDD.n3535 0.4505
R24847 DVDD.n3537 DVDD.n2486 0.4505
R24848 DVDD.n3539 DVDD.n3538 0.4505
R24849 DVDD.n2484 DVDD.n2483 0.4505
R24850 DVDD.n3544 DVDD.n3543 0.4505
R24851 DVDD.n3545 DVDD.n2482 0.4505
R24852 DVDD.n3547 DVDD.n3546 0.4505
R24853 DVDD.n2480 DVDD.n2479 0.4505
R24854 DVDD.n3552 DVDD.n3551 0.4505
R24855 DVDD.n3553 DVDD.n2478 0.4505
R24856 DVDD.n3555 DVDD.n3554 0.4505
R24857 DVDD.n2476 DVDD.n2475 0.4505
R24858 DVDD.n3560 DVDD.n3559 0.4505
R24859 DVDD.n3561 DVDD.n2474 0.4505
R24860 DVDD.n3563 DVDD.n3562 0.4505
R24861 DVDD.n2472 DVDD.n2471 0.4505
R24862 DVDD.n3568 DVDD.n3567 0.4505
R24863 DVDD.n3569 DVDD.n2470 0.4505
R24864 DVDD.n3571 DVDD.n3570 0.4505
R24865 DVDD.n2468 DVDD.n2467 0.4505
R24866 DVDD.n3576 DVDD.n3575 0.4505
R24867 DVDD.n3577 DVDD.n2466 0.4505
R24868 DVDD.n3579 DVDD.n3578 0.4505
R24869 DVDD.n2464 DVDD.n2463 0.4505
R24870 DVDD.n3584 DVDD.n3583 0.4505
R24871 DVDD.n3585 DVDD.n2462 0.4505
R24872 DVDD.n3587 DVDD.n3586 0.4505
R24873 DVDD.n2460 DVDD.n2459 0.4505
R24874 DVDD.n3592 DVDD.n3591 0.4505
R24875 DVDD.n3593 DVDD.n2458 0.4505
R24876 DVDD.n3595 DVDD.n3594 0.4505
R24877 DVDD.n2456 DVDD.n2455 0.4505
R24878 DVDD.n3600 DVDD.n3599 0.4505
R24879 DVDD.n2448 DVDD.n2441 0.4505
R24880 DVDD.n3605 DVDD.n3604 0.4505
R24881 DVDD.n3613 DVDD.n3612 0.4505
R24882 DVDD.n3611 DVDD.n2436 0.4505
R24883 DVDD.n3610 DVDD.n3609 0.4505
R24884 DVDD.n2439 DVDD.n2438 0.4505
R24885 DVDD.n3667 DVDD.n3666 0.4505
R24886 DVDD.n2406 DVDD.n1983 0.4505
R24887 DVDD.n3662 DVDD.n1988 0.4505
R24888 DVDD.n3661 DVDD.n3660 0.4505
R24889 DVDD.n3659 DVDD.n2408 0.4505
R24890 DVDD.n3658 DVDD.n3657 0.4505
R24891 DVDD.n2410 DVDD.n2409 0.4505
R24892 DVDD.n3653 DVDD.n3652 0.4505
R24893 DVDD.n3651 DVDD.n2413 0.4505
R24894 DVDD.n3650 DVDD.n3649 0.4505
R24895 DVDD.n2415 DVDD.n2414 0.4505
R24896 DVDD.n3645 DVDD.n3644 0.4505
R24897 DVDD.n3643 DVDD.n2417 0.4505
R24898 DVDD.n3642 DVDD.n3641 0.4505
R24899 DVDD.n2419 DVDD.n2418 0.4505
R24900 DVDD.n3637 DVDD.n3636 0.4505
R24901 DVDD.n3635 DVDD.n2421 0.4505
R24902 DVDD.n3634 DVDD.n3633 0.4505
R24903 DVDD.n2423 DVDD.n2422 0.4505
R24904 DVDD.n3629 DVDD.n3628 0.4505
R24905 DVDD.n3627 DVDD.n2425 0.4505
R24906 DVDD.n3626 DVDD.n3625 0.4505
R24907 DVDD.n2427 DVDD.n2426 0.4505
R24908 DVDD.n3621 DVDD.n3620 0.4505
R24909 DVDD.n3619 DVDD.n2429 0.4505
R24910 DVDD.n3618 DVDD.n3617 0.4505
R24911 DVDD.n2437 DVDD.n2434 0.4505
R24912 DVDD.n4125 DVDD.n4124 0.4505
R24913 DVDD.n3965 DVDD.n3932 0.4505
R24914 DVDD.n4079 DVDD.n4044 0.4505
R24915 DVDD.n4078 DVDD.n4077 0.4505
R24916 DVDD.n4076 DVDD.n4048 0.4505
R24917 DVDD.n4075 DVDD.n4074 0.4505
R24918 DVDD.n4050 DVDD.n4049 0.4505
R24919 DVDD.n4070 DVDD.n4069 0.4505
R24920 DVDD.n4055 DVDD.n4053 0.4505
R24921 DVDD.n4064 DVDD.n4063 0.4505
R24922 DVDD.n4060 DVDD.n4059 0.4505
R24923 DVDD.n1723 DVDD.n1721 0.4505
R24924 DVDD.n4226 DVDD.n4225 0.4505
R24925 DVDD.n1765 DVDD.n1764 0.4505
R24926 DVDD.n1729 DVDD.n1727 0.4505
R24927 DVDD.n1759 DVDD.n1758 0.4505
R24928 DVDD.n1734 DVDD.n1731 0.4505
R24929 DVDD.n1754 DVDD.n1753 0.4505
R24930 DVDD.n1752 DVDD.n1733 0.4505
R24931 DVDD.n1751 DVDD.n1750 0.4505
R24932 DVDD.n1736 DVDD.n1735 0.4505
R24933 DVDD.n1746 DVDD.n1745 0.4505
R24934 DVDD.n1744 DVDD.n1738 0.4505
R24935 DVDD.n1738 DVDD.n1737 0.4505
R24936 DVDD.n1747 DVDD.n1746 0.4505
R24937 DVDD.n1748 DVDD.n1736 0.4505
R24938 DVDD.n1750 DVDD.n1749 0.4505
R24939 DVDD.n1733 DVDD.n1732 0.4505
R24940 DVDD.n1755 DVDD.n1754 0.4505
R24941 DVDD.n1756 DVDD.n1731 0.4505
R24942 DVDD.n1758 DVDD.n1757 0.4505
R24943 DVDD.n1727 DVDD.n1726 0.4505
R24944 DVDD.n1766 DVDD.n1765 0.4505
R24945 DVDD.n4225 DVDD.n4224 0.4505
R24946 DVDD.n1725 DVDD.n1723 0.4505
R24947 DVDD.n4061 DVDD.n4060 0.4505
R24948 DVDD.n4063 DVDD.n4062 0.4505
R24949 DVDD.n4053 DVDD.n4052 0.4505
R24950 DVDD.n4071 DVDD.n4070 0.4505
R24951 DVDD.n4072 DVDD.n4050 0.4505
R24952 DVDD.n4074 DVDD.n4073 0.4505
R24953 DVDD.n4051 DVDD.n4048 0.4505
R24954 DVDD.n4078 DVDD.n4047 0.4505
R24955 DVDD.n4080 DVDD.n4079 0.4505
R24956 DVDD.n3901 DVDD.n3900 0.4505
R24957 DVDD.n3899 DVDD.n3872 0.4505
R24958 DVDD.n3898 DVDD.n3897 0.4505
R24959 DVDD.n3874 DVDD.n3873 0.4505
R24960 DVDD.n3893 DVDD.n3892 0.4505
R24961 DVDD.n3891 DVDD.n3877 0.4505
R24962 DVDD.n3890 DVDD.n3889 0.4505
R24963 DVDD.n3879 DVDD.n3878 0.4505
R24964 DVDD.n3885 DVDD.n3884 0.4505
R24965 DVDD.n3883 DVDD.n3882 0.4505
R24966 DVDD.n3881 DVDD.n1794 0.4505
R24967 DVDD.n4102 DVDD.n4101 0.4505
R24968 DVDD.n4100 DVDD.n1793 0.4505
R24969 DVDD.n4099 DVDD.n4098 0.4505
R24970 DVDD.n4037 DVDD.n4036 0.4505
R24971 DVDD.n4094 DVDD.n4093 0.4505
R24972 DVDD.n4092 DVDD.n4039 0.4505
R24973 DVDD.n4091 DVDD.n4090 0.4505
R24974 DVDD.n4041 DVDD.n4040 0.4505
R24975 DVDD.n4086 DVDD.n4085 0.4505
R24976 DVDD.n4084 DVDD.n4043 0.4505
R24977 DVDD.n4043 DVDD.n4042 0.4505
R24978 DVDD.n4087 DVDD.n4086 0.4505
R24979 DVDD.n4088 DVDD.n4041 0.4505
R24980 DVDD.n4090 DVDD.n4089 0.4505
R24981 DVDD.n4039 DVDD.n4038 0.4505
R24982 DVDD.n4095 DVDD.n4094 0.4505
R24983 DVDD.n4096 DVDD.n4037 0.4505
R24984 DVDD.n4098 DVDD.n4097 0.4505
R24985 DVDD.n1793 DVDD.n1791 0.4505
R24986 DVDD.n4103 DVDD.n4102 0.4505
R24987 DVDD.n3881 DVDD.n1790 0.4505
R24988 DVDD.n3882 DVDD.n3880 0.4505
R24989 DVDD.n3886 DVDD.n3885 0.4505
R24990 DVDD.n3887 DVDD.n3879 0.4505
R24991 DVDD.n3889 DVDD.n3888 0.4505
R24992 DVDD.n3877 DVDD.n3876 0.4505
R24993 DVDD.n3894 DVDD.n3893 0.4505
R24994 DVDD.n3895 DVDD.n3874 0.4505
R24995 DVDD.n3897 DVDD.n3896 0.4505
R24996 DVDD.n3875 DVDD.n3872 0.4505
R24997 DVDD.n3901 DVDD.n3869 0.4505
R24998 DVDD.n3905 DVDD.n3868 0.4505
R24999 DVDD.n3907 DVDD.n3906 0.4505
R25000 DVDD.n3866 DVDD.n3865 0.4505
R25001 DVDD.n3912 DVDD.n3911 0.4505
R25002 DVDD.n3913 DVDD.n3864 0.4505
R25003 DVDD.n3915 DVDD.n3914 0.4505
R25004 DVDD.n3862 DVDD.n3861 0.4505
R25005 DVDD.n3920 DVDD.n3919 0.4505
R25006 DVDD.n3921 DVDD.n3860 0.4505
R25007 DVDD.n3923 DVDD.n3922 0.4505
R25008 DVDD.n3857 DVDD.n3856 0.4505
R25009 DVDD.n3855 DVDD.n1820 0.4505
R25010 DVDD.n3854 DVDD.n3853 0.4505
R25011 DVDD.n1822 DVDD.n1821 0.4505
R25012 DVDD.n3849 DVDD.n3848 0.4505
R25013 DVDD.n3847 DVDD.n1824 0.4505
R25014 DVDD.n3846 DVDD.n3845 0.4505
R25015 DVDD.n1826 DVDD.n1825 0.4505
R25016 DVDD.n3841 DVDD.n3840 0.4505
R25017 DVDD.n3839 DVDD.n1828 0.4505
R25018 DVDD.n3838 DVDD.n3837 0.4505
R25019 DVDD.n3832 DVDD.n3831 0.4505
R25020 DVDD.n3830 DVDD.n1833 0.4505
R25021 DVDD.n3829 DVDD.n3828 0.4505
R25022 DVDD.n1835 DVDD.n1834 0.4505
R25023 DVDD.n3824 DVDD.n3823 0.4505
R25024 DVDD.n3822 DVDD.n1837 0.4505
R25025 DVDD.n3821 DVDD.n3820 0.4505
R25026 DVDD.n1839 DVDD.n1838 0.4505
R25027 DVDD.n3811 DVDD.n3810 0.4505
R25028 DVDD.n3809 DVDD.n1686 0.4505
R25029 DVDD.n4262 DVDD.n4261 0.4505
R25030 DVDD.n1678 DVDD.n1677 0.4505
R25031 DVDD.n4270 DVDD.n4269 0.4505
R25032 DVDD.n4271 DVDD.n1676 0.4505
R25033 DVDD.n4273 DVDD.n4272 0.4505
R25034 DVDD.n1674 DVDD.n1673 0.4505
R25035 DVDD.n4278 DVDD.n4277 0.4505
R25036 DVDD.n4279 DVDD.n1672 0.4505
R25037 DVDD.n4281 DVDD.n4280 0.4505
R25038 DVDD.n1669 DVDD.n1668 0.4505
R25039 DVDD.n4286 DVDD.n4285 0.4505
R25040 DVDD.n3837 DVDD.n3836 0.4505
R25041 DVDD.n1828 DVDD.n1827 0.4505
R25042 DVDD.n3842 DVDD.n3841 0.4505
R25043 DVDD.n3843 DVDD.n1826 0.4505
R25044 DVDD.n3845 DVDD.n3844 0.4505
R25045 DVDD.n1824 DVDD.n1823 0.4505
R25046 DVDD.n3850 DVDD.n3849 0.4505
R25047 DVDD.n3851 DVDD.n1822 0.4505
R25048 DVDD.n3853 DVDD.n3852 0.4505
R25049 DVDD.n1820 DVDD.n1819 0.4505
R25050 DVDD.n3858 DVDD.n3857 0.4505
R25051 DVDD.n3924 DVDD.n3923 0.4505
R25052 DVDD.n3860 DVDD.n3859 0.4505
R25053 DVDD.n3919 DVDD.n3918 0.4505
R25054 DVDD.n3917 DVDD.n3862 0.4505
R25055 DVDD.n3916 DVDD.n3915 0.4505
R25056 DVDD.n3864 DVDD.n3863 0.4505
R25057 DVDD.n3911 DVDD.n3910 0.4505
R25058 DVDD.n3909 DVDD.n3866 0.4505
R25059 DVDD.n3908 DVDD.n3907 0.4505
R25060 DVDD.n3868 DVDD.n3867 0.4505
R25061 DVDD.n4285 DVDD.n4284 0.4505
R25062 DVDD.n4283 DVDD.n1669 0.4505
R25063 DVDD.n4282 DVDD.n4281 0.4505
R25064 DVDD.n1672 DVDD.n1671 0.4505
R25065 DVDD.n4277 DVDD.n4276 0.4505
R25066 DVDD.n4275 DVDD.n1674 0.4505
R25067 DVDD.n4274 DVDD.n4273 0.4505
R25068 DVDD.n1679 DVDD.n1676 0.4505
R25069 DVDD.n4269 DVDD.n4268 0.4505
R25070 DVDD.n1681 DVDD.n1678 0.4505
R25071 DVDD.n4263 DVDD.n4262 0.4505
R25072 DVDD.n3809 DVDD.n3808 0.4505
R25073 DVDD.n3812 DVDD.n3811 0.4505
R25074 DVDD.n3813 DVDD.n1839 0.4505
R25075 DVDD.n3820 DVDD.n3819 0.4505
R25076 DVDD.n1841 DVDD.n1837 0.4505
R25077 DVDD.n3825 DVDD.n3824 0.4505
R25078 DVDD.n3826 DVDD.n1835 0.4505
R25079 DVDD.n3828 DVDD.n3827 0.4505
R25080 DVDD.n1833 DVDD.n1832 0.4505
R25081 DVDD.n3833 DVDD.n3832 0.4505
R25082 DVDD.n1571 DVDD.n1570 0.4505
R25083 DVDD.n1569 DVDD.n1206 0.4505
R25084 DVDD.n1568 DVDD.n1567 0.4505
R25085 DVDD.n1208 DVDD.n1207 0.4505
R25086 DVDD.n1563 DVDD.n1562 0.4505
R25087 DVDD.n1561 DVDD.n1211 0.4505
R25088 DVDD.n1560 DVDD.n1559 0.4505
R25089 DVDD.n1213 DVDD.n1212 0.4505
R25090 DVDD.n1226 DVDD.n1224 0.4505
R25091 DVDD.n1552 DVDD.n1551 0.4505
R25092 DVDD.n1550 DVDD.n1225 0.4505
R25093 DVDD.n1549 DVDD.n1548 0.4505
R25094 DVDD.n1228 DVDD.n1227 0.4505
R25095 DVDD.n1544 DVDD.n1543 0.4505
R25096 DVDD.n1542 DVDD.n1230 0.4505
R25097 DVDD.n1541 DVDD.n1540 0.4505
R25098 DVDD.n1232 DVDD.n1231 0.4505
R25099 DVDD.n1536 DVDD.n1535 0.4505
R25100 DVDD.n1534 DVDD.n1234 0.4505
R25101 DVDD.n1533 DVDD.n1532 0.4505
R25102 DVDD.n1236 DVDD.n1235 0.4505
R25103 DVDD.n1528 DVDD.n1527 0.4505
R25104 DVDD.n1526 DVDD.n1238 0.4505
R25105 DVDD.n1525 DVDD.n1524 0.4505
R25106 DVDD.n1240 DVDD.n1239 0.4505
R25107 DVDD.n1520 DVDD.n1519 0.4505
R25108 DVDD.n1518 DVDD.n1242 0.4505
R25109 DVDD.n1517 DVDD.n1516 0.4505
R25110 DVDD.n1244 DVDD.n1243 0.4505
R25111 DVDD.n1512 DVDD.n1511 0.4505
R25112 DVDD.n1510 DVDD.n1246 0.4505
R25113 DVDD.n1509 DVDD.n1508 0.4505
R25114 DVDD.n1248 DVDD.n1247 0.4505
R25115 DVDD.n1504 DVDD.n1503 0.4505
R25116 DVDD.n1502 DVDD.n1250 0.4505
R25117 DVDD.n1501 DVDD.n1500 0.4505
R25118 DVDD.n1252 DVDD.n1251 0.4505
R25119 DVDD.n1496 DVDD.n1495 0.4505
R25120 DVDD.n1494 DVDD.n1254 0.4505
R25121 DVDD.n1493 DVDD.n1492 0.4505
R25122 DVDD.n1256 DVDD.n1255 0.4505
R25123 DVDD.n1488 DVDD.n1487 0.4505
R25124 DVDD.n1486 DVDD.n1258 0.4505
R25125 DVDD.n1485 DVDD.n1484 0.4505
R25126 DVDD.n1260 DVDD.n1259 0.4505
R25127 DVDD.n1480 DVDD.n1479 0.4505
R25128 DVDD.n1478 DVDD.n1262 0.4505
R25129 DVDD.n1477 DVDD.n1476 0.4505
R25130 DVDD.n1264 DVDD.n1263 0.4505
R25131 DVDD.n1472 DVDD.n1471 0.4505
R25132 DVDD.n1470 DVDD.n1266 0.4505
R25133 DVDD.n1469 DVDD.n1468 0.4505
R25134 DVDD.n1268 DVDD.n1267 0.4505
R25135 DVDD.n1464 DVDD.n1463 0.4505
R25136 DVDD.n1462 DVDD.n1270 0.4505
R25137 DVDD.n1461 DVDD.n1460 0.4505
R25138 DVDD.n1272 DVDD.n1271 0.4505
R25139 DVDD.n1456 DVDD.n1455 0.4505
R25140 DVDD.n1454 DVDD.n1274 0.4505
R25141 DVDD.n1453 DVDD.n1452 0.4505
R25142 DVDD.n1276 DVDD.n1275 0.4505
R25143 DVDD.n1448 DVDD.n1447 0.4505
R25144 DVDD.n1446 DVDD.n1278 0.4505
R25145 DVDD.n1445 DVDD.n1444 0.4505
R25146 DVDD.n1280 DVDD.n1279 0.4505
R25147 DVDD.n1440 DVDD.n1439 0.4505
R25148 DVDD.n1438 DVDD.n1282 0.4505
R25149 DVDD.n1437 DVDD.n1436 0.4505
R25150 DVDD.n1284 DVDD.n1283 0.4505
R25151 DVDD.n1432 DVDD.n1431 0.4505
R25152 DVDD.n1430 DVDD.n1286 0.4505
R25153 DVDD.n1429 DVDD.n1428 0.4505
R25154 DVDD.n1288 DVDD.n1287 0.4505
R25155 DVDD.n1424 DVDD.n1423 0.4505
R25156 DVDD.n1422 DVDD.n1290 0.4505
R25157 DVDD.n1421 DVDD.n1420 0.4505
R25158 DVDD.n1292 DVDD.n1291 0.4505
R25159 DVDD.n1416 DVDD.n1415 0.4505
R25160 DVDD.n1414 DVDD.n1294 0.4505
R25161 DVDD.n1413 DVDD.n1412 0.4505
R25162 DVDD.n1296 DVDD.n1295 0.4505
R25163 DVDD.n1408 DVDD.n1407 0.4505
R25164 DVDD.n1406 DVDD.n1298 0.4505
R25165 DVDD.n1405 DVDD.n1404 0.4505
R25166 DVDD.n1300 DVDD.n1299 0.4505
R25167 DVDD.n1400 DVDD.n1399 0.4505
R25168 DVDD.n1398 DVDD.n1302 0.4505
R25169 DVDD.n1397 DVDD.n1396 0.4505
R25170 DVDD.n1304 DVDD.n1303 0.4505
R25171 DVDD.n1347 DVDD.n1346 0.4505
R25172 DVDD.n1351 DVDD.n1350 0.4505
R25173 DVDD.n1352 DVDD.n1345 0.4505
R25174 DVDD.n1354 DVDD.n1353 0.4505
R25175 DVDD.n1343 DVDD.n1342 0.4505
R25176 DVDD.n1359 DVDD.n1358 0.4505
R25177 DVDD.n1361 DVDD.n1360 0.4505
R25178 DVDD.n1205 DVDD.n1197 0.4505
R25179 DVDD.n1572 DVDD.n1571 0.4505
R25180 DVDD.n1209 DVDD.n1206 0.4505
R25181 DVDD.n1567 DVDD.n1566 0.4505
R25182 DVDD.n1565 DVDD.n1208 0.4505
R25183 DVDD.n1564 DVDD.n1563 0.4505
R25184 DVDD.n1211 DVDD.n1210 0.4505
R25185 DVDD.n1559 DVDD.n1558 0.4505
R25186 DVDD.n1557 DVDD.n1213 0.4505
R25187 DVDD.n1224 DVDD.n1218 0.4505
R25188 DVDD.n1553 DVDD.n1552 0.4505
R25189 DVDD.n1225 DVDD.n1223 0.4505
R25190 DVDD.n1548 DVDD.n1547 0.4505
R25191 DVDD.n1546 DVDD.n1228 0.4505
R25192 DVDD.n1545 DVDD.n1544 0.4505
R25193 DVDD.n1230 DVDD.n1229 0.4505
R25194 DVDD.n1540 DVDD.n1539 0.4505
R25195 DVDD.n1538 DVDD.n1232 0.4505
R25196 DVDD.n1537 DVDD.n1536 0.4505
R25197 DVDD.n1234 DVDD.n1233 0.4505
R25198 DVDD.n1532 DVDD.n1531 0.4505
R25199 DVDD.n1530 DVDD.n1236 0.4505
R25200 DVDD.n1529 DVDD.n1528 0.4505
R25201 DVDD.n1238 DVDD.n1237 0.4505
R25202 DVDD.n1524 DVDD.n1523 0.4505
R25203 DVDD.n1522 DVDD.n1240 0.4505
R25204 DVDD.n1521 DVDD.n1520 0.4505
R25205 DVDD.n1242 DVDD.n1241 0.4505
R25206 DVDD.n1516 DVDD.n1515 0.4505
R25207 DVDD.n1514 DVDD.n1244 0.4505
R25208 DVDD.n1513 DVDD.n1512 0.4505
R25209 DVDD.n1246 DVDD.n1245 0.4505
R25210 DVDD.n1508 DVDD.n1507 0.4505
R25211 DVDD.n1506 DVDD.n1248 0.4505
R25212 DVDD.n1505 DVDD.n1504 0.4505
R25213 DVDD.n1250 DVDD.n1249 0.4505
R25214 DVDD.n1500 DVDD.n1499 0.4505
R25215 DVDD.n1498 DVDD.n1252 0.4505
R25216 DVDD.n1497 DVDD.n1496 0.4505
R25217 DVDD.n1254 DVDD.n1253 0.4505
R25218 DVDD.n1492 DVDD.n1491 0.4505
R25219 DVDD.n1490 DVDD.n1256 0.4505
R25220 DVDD.n1489 DVDD.n1488 0.4505
R25221 DVDD.n1258 DVDD.n1257 0.4505
R25222 DVDD.n1484 DVDD.n1483 0.4505
R25223 DVDD.n1482 DVDD.n1260 0.4505
R25224 DVDD.n1481 DVDD.n1480 0.4505
R25225 DVDD.n1262 DVDD.n1261 0.4505
R25226 DVDD.n1476 DVDD.n1475 0.4505
R25227 DVDD.n1474 DVDD.n1264 0.4505
R25228 DVDD.n1473 DVDD.n1472 0.4505
R25229 DVDD.n1266 DVDD.n1265 0.4505
R25230 DVDD.n1468 DVDD.n1467 0.4505
R25231 DVDD.n1466 DVDD.n1268 0.4505
R25232 DVDD.n1465 DVDD.n1464 0.4505
R25233 DVDD.n1270 DVDD.n1269 0.4505
R25234 DVDD.n1460 DVDD.n1459 0.4505
R25235 DVDD.n1458 DVDD.n1272 0.4505
R25236 DVDD.n1457 DVDD.n1456 0.4505
R25237 DVDD.n1274 DVDD.n1273 0.4505
R25238 DVDD.n1452 DVDD.n1451 0.4505
R25239 DVDD.n1450 DVDD.n1276 0.4505
R25240 DVDD.n1449 DVDD.n1448 0.4505
R25241 DVDD.n1278 DVDD.n1277 0.4505
R25242 DVDD.n1444 DVDD.n1443 0.4505
R25243 DVDD.n1442 DVDD.n1280 0.4505
R25244 DVDD.n1441 DVDD.n1440 0.4505
R25245 DVDD.n1282 DVDD.n1281 0.4505
R25246 DVDD.n1436 DVDD.n1435 0.4505
R25247 DVDD.n1434 DVDD.n1284 0.4505
R25248 DVDD.n1433 DVDD.n1432 0.4505
R25249 DVDD.n1286 DVDD.n1285 0.4505
R25250 DVDD.n1428 DVDD.n1427 0.4505
R25251 DVDD.n1426 DVDD.n1288 0.4505
R25252 DVDD.n1425 DVDD.n1424 0.4505
R25253 DVDD.n1290 DVDD.n1289 0.4505
R25254 DVDD.n1420 DVDD.n1419 0.4505
R25255 DVDD.n1418 DVDD.n1292 0.4505
R25256 DVDD.n1417 DVDD.n1416 0.4505
R25257 DVDD.n1294 DVDD.n1293 0.4505
R25258 DVDD.n1412 DVDD.n1411 0.4505
R25259 DVDD.n1410 DVDD.n1296 0.4505
R25260 DVDD.n1409 DVDD.n1408 0.4505
R25261 DVDD.n1298 DVDD.n1297 0.4505
R25262 DVDD.n1404 DVDD.n1403 0.4505
R25263 DVDD.n1402 DVDD.n1300 0.4505
R25264 DVDD.n1401 DVDD.n1400 0.4505
R25265 DVDD.n1302 DVDD.n1301 0.4505
R25266 DVDD.n1396 DVDD.n1395 0.4505
R25267 DVDD.n1310 DVDD.n1304 0.4505
R25268 DVDD.n1348 DVDD.n1347 0.4505
R25269 DVDD.n1350 DVDD.n1349 0.4505
R25270 DVDD.n1345 DVDD.n1344 0.4505
R25271 DVDD.n1355 DVDD.n1354 0.4505
R25272 DVDD.n1356 DVDD.n1343 0.4505
R25273 DVDD.n1358 DVDD.n1357 0.4505
R25274 DVDD.n1361 DVDD.n1337 0.4505
R25275 DVDD.n1362 DVDD.n1340 0.4505
R25276 DVDD.n2603 DVDD.n2602 0.449506
R25277 DVDD.n1937 DVDD 0.448132
R25278 DVDD.n3210 DVDD.n2745 0.447304
R25279 DVDD DVDD.n2038 0.4405
R25280 DVDD.n4344 DVDD.n4301 0.437225
R25281 DVDD.n1946 DVDD.n1945 0.427206
R25282 DVDD.n2432 DVDD.n2431 0.423396
R25283 DVDD.n4239 DVDD.n4238 0.4205
R25284 DVDD.n4236 DVDD.n4235 0.4205
R25285 DVDD.n2200 DVDD 0.418417
R25286 DVDD.n2201 DVDD 0.418417
R25287 DVDD.n2016 DVDD.n2015 0.417167
R25288 DVDD.n2020 DVDD.n2019 0.417167
R25289 DVDD.n2024 DVDD.n2023 0.417167
R25290 DVDD.n2028 DVDD.n2027 0.417167
R25291 DVDD.n2032 DVDD.n2031 0.417167
R25292 DVDD.n2036 DVDD.n2035 0.417167
R25293 DVDD.n2037 DVDD.n2034 0.417167
R25294 DVDD.n2033 DVDD.n2030 0.417167
R25295 DVDD.n2029 DVDD.n2026 0.417167
R25296 DVDD.n2025 DVDD.n2022 0.417167
R25297 DVDD.n2021 DVDD.n2018 0.417167
R25298 DVDD.n2017 DVDD.n2014 0.417167
R25299 DVDD DVDD.n2124 0.414765
R25300 DVDD.n2266 DVDD 0.414765
R25301 DVDD DVDD.n2060 0.414765
R25302 DVDD.n2341 DVDD 0.414765
R25303 DVDD.n1881 DVDD.n1879 0.413789
R25304 DVDD.n3204 DVDD.n3117 0.41077
R25305 DVDD.n3213 DVDD.n3119 0.41077
R25306 DVDD.n3171 DVDD.n3108 0.41077
R25307 DVDD.n3226 DVDD.n3106 0.41077
R25308 DVDD.n2604 DVDD.n2510 0.402145
R25309 DVDD.n2539 DVDD.n2510 0.399579
R25310 DVDD DVDD.n1710 0.397559
R25311 DVDD DVDD.n1710 0.397559
R25312 DVDD.n3205 DVDD.n3204 0.391716
R25313 DVDD.n3119 DVDD.n3085 0.391716
R25314 DVDD.n3154 DVDD.n3153 0.376594
R25315 DVDD.n3218 DVDD.n3114 0.376594
R25316 DVDD.n3170 DVDD.n3169 0.3755
R25317 DVDD.n3228 DVDD.n3227 0.3755
R25318 DVDD.n3231 DVDD.n3230 0.3755
R25319 DVDD.n3168 DVDD.n3167 0.3755
R25320 DVDD.n1946 DVDD.n1937 0.36126
R25321 DVDD.t189 DVDD.n1883 0.3605
R25322 DVDD.t119 DVDD.n1709 0.3605
R25323 DVDD.t127 DVDD.n1711 0.3605
R25324 DVDD.t144 DVDD.n4190 0.3605
R25325 DVDD.n4138 DVDD.t124 0.360167
R25326 DVDD.n1785 DVDD.t136 0.360167
R25327 DVDD.n3966 DVDD.t40 0.360167
R25328 DVDD.n3962 DVDD.t38 0.360167
R25329 DVDD.n1874 DVDD.t30 0.360167
R25330 DVDD.n1872 DVDD.t32 0.360167
R25331 DVDD.n1714 DVDD.t171 0.360167
R25332 DVDD.n1717 DVDD.t70 0.360167
R25333 DVDD.n3691 DVDD.n1902 0.356801
R25334 DVDD.n3691 DVDD.n1906 0.356801
R25335 DVDD.n2720 DVDD.n2710 0.35585
R25336 DVDD.n2720 DVDD.n2714 0.35585
R25337 DVDD.n2720 DVDD.n2712 0.35585
R25338 DVDD.n4083 DVDD.n4082 0.35585
R25339 DVDD.n3903 DVDD.n3871 0.35585
R25340 DVDD.n3255 DVDD.n2741 0.355594
R25341 DVDD.n4083 DVDD.n4045 0.355001
R25342 DVDD.n3691 DVDD.n1897 0.35492
R25343 DVDD.n3255 DVDD.n2746 0.35492
R25344 DVDD.n3835 DVDD.n3834 0.35492
R25345 DVDD.n2720 DVDD.n2707 0.354416
R25346 DVDD.n2720 DVDD.n2711 0.354416
R25347 DVDD.n2720 DVDD.n2713 0.354416
R25348 DVDD.n3871 DVDD.n3870 0.354416
R25349 DVDD.n3691 DVDD.n1905 0.35405
R25350 DVDD.n3691 DVDD.n1909 0.35405
R25351 DVDD.n3255 DVDD.n2740 0.35312
R25352 DVDD.n3255 DVDD.n2747 0.35312
R25353 DVDD.n3835 DVDD.n1831 0.35312
R25354 DVDD.n2983 DVDD.n2686 0.346654
R25355 DVDD.n3420 DVDD.n2688 0.346654
R25356 DVDD.n1881 DVDD.n1880 0.346654
R25357 DVDD.n4230 DVDD.n4229 0.346654
R25358 DVDD.n3707 DVDD.n1902 0.340118
R25359 DVDD.n3707 DVDD.n1906 0.340118
R25360 DVDD.n3707 DVDD.n1897 0.339393
R25361 DVDD.n3389 DVDD.n2746 0.339393
R25362 DVDD.n3834 DVDD.n1829 0.339393
R25363 DVDD.n4081 DVDD.n4045 0.338918
R25364 DVDD.n3389 DVDD.n2741 0.33872
R25365 DVDD.n2711 DVDD.n2701 0.33857
R25366 DVDD.n2713 DVDD.n2701 0.33857
R25367 DVDD.n2707 DVDD.n2701 0.33857
R25368 DVDD.n3904 DVDD.n3870 0.33857
R25369 DVDD.n2710 DVDD.n2701 0.338454
R25370 DVDD.n2714 DVDD.n2701 0.338454
R25371 DVDD.n2712 DVDD.n2701 0.338454
R25372 DVDD.n4082 DVDD.n4081 0.338454
R25373 DVDD.n3904 DVDD.n3903 0.338454
R25374 DVDD.n1831 DVDD.n1829 0.338193
R25375 DVDD.n3389 DVDD.n2747 0.338193
R25376 DVDD.n3389 DVDD.n2740 0.338193
R25377 DVDD.n2593 DVDD.n2529 0.337345
R25378 DVDD.n2543 DVDD.n2538 0.337345
R25379 DVDD.n2591 DVDD.n2546 0.337345
R25380 DVDD.n2588 DVDD.n2586 0.337345
R25381 DVDD.n2582 DVDD.n2552 0.337345
R25382 DVDD.n2580 DVDD.n2565 0.337345
R25383 DVDD.n2559 DVDD.n2556 0.337345
R25384 DVDD.n2571 DVDD.n2560 0.337345
R25385 DVDD.n2570 DVDD.n2557 0.337345
R25386 DVDD.n2569 DVDD.n2558 0.337345
R25387 DVDD.n2571 DVDD.n2557 0.337345
R25388 DVDD.n2565 DVDD.n2556 0.337345
R25389 DVDD.n2564 DVDD.n2552 0.337345
R25390 DVDD.n2588 DVDD.n2546 0.337345
R25391 DVDD.n2538 DVDD.n2529 0.337345
R25392 DVDD.n2574 DVDD.n2570 0.337345
R25393 DVDD.n2560 DVDD.n2559 0.337345
R25394 DVDD.n2591 DVDD.n2543 0.337345
R25395 DVDD.n2586 DVDD.n2542 0.337345
R25396 DVDD.n2574 DVDD.n2558 0.337345
R25397 DVDD.n3707 DVDD.n1905 0.337254
R25398 DVDD.n3707 DVDD.n1909 0.337254
R25399 DVDD.n3389 DVDD.n2745 0.327632
R25400 DVDD.n4230 DVDD.n1718 0.313132
R25401 DVDD.n4150 DVDD.n4149 0.306049
R25402 DVDD.n1873 DVDD.n1706 0.306049
R25403 DVDD.n3961 DVDD.n3960 0.306049
R25404 DVDD.n4140 DVDD.n4139 0.306049
R25405 DVDD.n1962 DVDD.t188 0.303833
R25406 DVDD.n1962 DVDD.t165 0.303833
R25407 DVDD.n1958 DVDD.t132 0.303833
R25408 DVDD.n1958 DVDD.t149 0.303833
R25409 DVDD.n1930 DVDD.t118 0.303833
R25410 DVDD.n1930 DVDD.t175 0.303833
R25411 DVDD.n1931 DVDD.t92 0.303833
R25412 DVDD.n1931 DVDD.t140 0.303833
R25413 DVDD.n85 DVDD.n84 0.3005
R25414 DVDD.n333 DVDD.n329 0.3005
R25415 DVDD.n2592 DVDD.n2541 0.291153
R25416 DVDD.n1875 DVDD.n1708 0.265206
R25417 DVDD.n3963 DVDD.n1708 0.265206
R25418 DVDD.n4234 DVDD.n1713 0.265206
R25419 DVDD.n4234 DVDD.n4233 0.265206
R25420 DVDD.n2603 DVDD.n2507 0.260889
R25421 DVDD.n1966 DVDD 0.258658
R25422 DVDD.n2518 DVDD.n2517 0.252737
R25423 DVDD.n5506 DVDD.n219 0.2505
R25424 DVDD.n966 DVDD.n945 0.2505
R25425 DVDD.n3169 DVDD.n3168 0.242734
R25426 DVDD.n3230 DVDD.n3228 0.242734
R25427 DVDD.n2013 DVDD 0.232667
R25428 DVDD.n3169 DVDD.n3155 0.231484
R25429 DVDD.n3230 DVDD.n3229 0.231484
R25430 DVDD.n2397 DVDD.n2039 0.231338
R25431 DVDD.n3665 DVDD.n3664 0.231338
R25432 DVDD.n5917 DVDD.n103 0.22706
R25433 DVDD.n5422 DVDD.n5420 0.225937
R25434 DVDD.n928 DVDD.n263 0.224497
R25435 DVDD.n259 DVDD.n258 0.224242
R25436 DVDD.n2431 DVDD 0.224176
R25437 DVDD.n3777 DVDD.n3723 0.221159
R25438 DVDD.n1150 DVDD.n1120 0.221159
R25439 DVDD.n4413 DVDD.n4401 0.221159
R25440 DVDD.n4347 DVDD.n1595 0.221159
R25441 DVDD.n4302 DVDD.n1627 0.221159
R25442 DVDD.n2976 DVDD.n2970 0.219787
R25443 DVDD.n3233 DVDD.n3097 0.217529
R25444 DVDD.n3165 DVDD.n3162 0.217529
R25445 DVDD.n4330 DVDD.n4303 0.214786
R25446 DVDD.n4329 DVDD.n4304 0.214786
R25447 DVDD.n4328 DVDD.n4305 0.214786
R25448 DVDD.n4308 DVDD.n4306 0.214786
R25449 DVDD.n4324 DVDD.n4309 0.214786
R25450 DVDD.n4323 DVDD.n4310 0.214786
R25451 DVDD.n4322 DVDD.n4311 0.214786
R25452 DVDD.n4314 DVDD.n4312 0.214786
R25453 DVDD.n4318 DVDD.n4315 0.214786
R25454 DVDD.n4317 DVDD.n4316 0.214786
R25455 DVDD.n913 DVDD.n912 0.214786
R25456 DVDD.n4715 DVDD.n4714 0.214786
R25457 DVDD.n4716 DVDD.n911 0.214786
R25458 DVDD.n4718 DVDD.n4717 0.214786
R25459 DVDD.n4723 DVDD.n4722 0.214786
R25460 DVDD.n4724 DVDD.n906 0.214786
R25461 DVDD.n4726 DVDD.n4725 0.214786
R25462 DVDD.n904 DVDD.n903 0.214786
R25463 DVDD.n4731 DVDD.n4730 0.214786
R25464 DVDD.n4732 DVDD.n902 0.214786
R25465 DVDD.n4734 DVDD.n4733 0.214786
R25466 DVDD.n900 DVDD.n899 0.214786
R25467 DVDD.n4739 DVDD.n4738 0.214786
R25468 DVDD.n4740 DVDD.n898 0.214786
R25469 DVDD.n4742 DVDD.n4741 0.214786
R25470 DVDD.n890 DVDD.n889 0.214786
R25471 DVDD.n4749 DVDD.n4748 0.214786
R25472 DVDD.n4750 DVDD.n888 0.214786
R25473 DVDD.n4752 DVDD.n4751 0.214786
R25474 DVDD.n886 DVDD.n885 0.214786
R25475 DVDD.n4757 DVDD.n4756 0.214786
R25476 DVDD.n4758 DVDD.n884 0.214786
R25477 DVDD.n4760 DVDD.n4759 0.214786
R25478 DVDD.n882 DVDD.n881 0.214786
R25479 DVDD.n4765 DVDD.n4764 0.214786
R25480 DVDD.n4766 DVDD.n880 0.214786
R25481 DVDD.n4770 DVDD.n4769 0.214786
R25482 DVDD.n4768 DVDD.n732 0.214786
R25483 DVDD.n4803 DVDD.n733 0.214786
R25484 DVDD.n4777 DVDD.n734 0.214786
R25485 DVDD.n4799 DVDD.n4778 0.214786
R25486 DVDD.n4798 DVDD.n4779 0.214786
R25487 DVDD.n4797 DVDD.n4780 0.214786
R25488 DVDD.n4783 DVDD.n4781 0.214786
R25489 DVDD.n4793 DVDD.n4784 0.214786
R25490 DVDD.n4792 DVDD.n4785 0.214786
R25491 DVDD.n4791 DVDD.n4786 0.214786
R25492 DVDD.n4788 DVDD.n4787 0.214786
R25493 DVDD.n587 DVDD.n586 0.214786
R25494 DVDD.n5025 DVDD.n5024 0.214786
R25495 DVDD.n5026 DVDD.n585 0.214786
R25496 DVDD.n5028 DVDD.n5027 0.214786
R25497 DVDD.n583 DVDD.n582 0.214786
R25498 DVDD.n5033 DVDD.n5032 0.214786
R25499 DVDD.n5034 DVDD.n581 0.214786
R25500 DVDD.n5036 DVDD.n5035 0.214786
R25501 DVDD.n579 DVDD.n578 0.214786
R25502 DVDD.n5041 DVDD.n5040 0.214786
R25503 DVDD.n5042 DVDD.n577 0.214786
R25504 DVDD.n5044 DVDD.n5043 0.214786
R25505 DVDD.n575 DVDD.n574 0.214786
R25506 DVDD.n5049 DVDD.n5048 0.214786
R25507 DVDD.n5086 DVDD.n5051 0.214786
R25508 DVDD.n5085 DVDD.n5052 0.214786
R25509 DVDD.n5055 DVDD.n5053 0.214786
R25510 DVDD.n5081 DVDD.n5056 0.214786
R25511 DVDD.n5080 DVDD.n5057 0.214786
R25512 DVDD.n5079 DVDD.n5058 0.214786
R25513 DVDD.n5061 DVDD.n5059 0.214786
R25514 DVDD.n5075 DVDD.n5062 0.214786
R25515 DVDD.n5074 DVDD.n5063 0.214786
R25516 DVDD.n5073 DVDD.n5064 0.214786
R25517 DVDD.n5066 DVDD.n5065 0.214786
R25518 DVDD.n5069 DVDD.n5068 0.214786
R25519 DVDD.n5067 DVDD.n200 0.214786
R25520 DVDD.n5728 DVDD.n201 0.214786
R25521 DVDD.n5727 DVDD.n202 0.214786
R25522 DVDD.n5726 DVDD.n203 0.214786
R25523 DVDD.n206 DVDD.n204 0.214786
R25524 DVDD.n5722 DVDD.n207 0.214786
R25525 DVDD.n5721 DVDD.n208 0.214786
R25526 DVDD.n5720 DVDD.n209 0.214786
R25527 DVDD.n212 DVDD.n210 0.214786
R25528 DVDD.n5716 DVDD.n213 0.214786
R25529 DVDD.n5715 DVDD.n214 0.214786
R25530 DVDD.n5714 DVDD.n215 0.214786
R25531 DVDD.n5711 DVDD.n216 0.214786
R25532 DVDD.n5675 DVDD.n217 0.214786
R25533 DVDD.n5702 DVDD.n5676 0.214786
R25534 DVDD.n5701 DVDD.n5677 0.214786
R25535 DVDD.n5700 DVDD.n5678 0.214786
R25536 DVDD.n5699 DVDD.n5679 0.214786
R25537 DVDD.n5682 DVDD.n5680 0.214786
R25538 DVDD.n5695 DVDD.n5683 0.214786
R25539 DVDD.n5694 DVDD.n5684 0.214786
R25540 DVDD.n5693 DVDD.n5685 0.214786
R25541 DVDD.n5687 DVDD.n5686 0.214786
R25542 DVDD.n5689 DVDD.n5688 0.214786
R25543 DVDD.n4373 DVDD.n4348 0.214786
R25544 DVDD.n4372 DVDD.n4349 0.214786
R25545 DVDD.n4371 DVDD.n4350 0.214786
R25546 DVDD.n4353 DVDD.n4351 0.214786
R25547 DVDD.n4367 DVDD.n4354 0.214786
R25548 DVDD.n4366 DVDD.n4355 0.214786
R25549 DVDD.n4365 DVDD.n4356 0.214786
R25550 DVDD.n4358 DVDD.n4357 0.214786
R25551 DVDD.n4361 DVDD.n4360 0.214786
R25552 DVDD.n4359 DVDD.n985 0.214786
R25553 DVDD.n4644 DVDD.n986 0.214786
R25554 DVDD.n4643 DVDD.n987 0.214786
R25555 DVDD.n4641 DVDD.n988 0.214786
R25556 DVDD.n4639 DVDD.n989 0.214786
R25557 DVDD.n4636 DVDD.n991 0.214786
R25558 DVDD.n994 DVDD.n992 0.214786
R25559 DVDD.n4632 DVDD.n995 0.214786
R25560 DVDD.n4631 DVDD.n996 0.214786
R25561 DVDD.n4630 DVDD.n997 0.214786
R25562 DVDD.n1000 DVDD.n998 0.214786
R25563 DVDD.n4626 DVDD.n1001 0.214786
R25564 DVDD.n4625 DVDD.n1002 0.214786
R25565 DVDD.n4624 DVDD.n1003 0.214786
R25566 DVDD.n1006 DVDD.n1004 0.214786
R25567 DVDD.n4620 DVDD.n1007 0.214786
R25568 DVDD.n4619 DVDD.n1008 0.214786
R25569 DVDD.n1021 DVDD.n1009 0.214786
R25570 DVDD.n1044 DVDD.n1022 0.214786
R25571 DVDD.n1043 DVDD.n1023 0.214786
R25572 DVDD.n1042 DVDD.n1024 0.214786
R25573 DVDD.n1027 DVDD.n1025 0.214786
R25574 DVDD.n1038 DVDD.n1028 0.214786
R25575 DVDD.n1037 DVDD.n1029 0.214786
R25576 DVDD.n1036 DVDD.n1030 0.214786
R25577 DVDD.n1033 DVDD.n1032 0.214786
R25578 DVDD.n1031 DVDD.n729 0.214786
R25579 DVDD.n4875 DVDD.n730 0.214786
R25580 DVDD.n4874 DVDD.n731 0.214786
R25581 DVDD.n4872 DVDD.n4805 0.214786
R25582 DVDD.n4871 DVDD.n4806 0.214786
R25583 DVDD.n4809 DVDD.n4807 0.214786
R25584 DVDD.n4867 DVDD.n4810 0.214786
R25585 DVDD.n4866 DVDD.n4811 0.214786
R25586 DVDD.n4865 DVDD.n4812 0.214786
R25587 DVDD.n4815 DVDD.n4813 0.214786
R25588 DVDD.n4861 DVDD.n4816 0.214786
R25589 DVDD.n4860 DVDD.n4817 0.214786
R25590 DVDD.n4859 DVDD.n4818 0.214786
R25591 DVDD.n4856 DVDD.n4819 0.214786
R25592 DVDD.n4855 DVDD.n4820 0.214786
R25593 DVDD.n4854 DVDD.n4821 0.214786
R25594 DVDD.n4853 DVDD.n4822 0.214786
R25595 DVDD.n4825 DVDD.n4823 0.214786
R25596 DVDD.n4849 DVDD.n4826 0.214786
R25597 DVDD.n4848 DVDD.n4827 0.214786
R25598 DVDD.n4847 DVDD.n4828 0.214786
R25599 DVDD.n4831 DVDD.n4829 0.214786
R25600 DVDD.n4843 DVDD.n4832 0.214786
R25601 DVDD.n4842 DVDD.n4833 0.214786
R25602 DVDD.n4841 DVDD.n4834 0.214786
R25603 DVDD.n4837 DVDD.n4836 0.214786
R25604 DVDD.n4835 DVDD.n482 0.214786
R25605 DVDD.n5246 DVDD.n483 0.214786
R25606 DVDD.n497 DVDD.n484 0.214786
R25607 DVDD.n553 DVDD.n498 0.214786
R25608 DVDD.n552 DVDD.n499 0.214786
R25609 DVDD.n551 DVDD.n500 0.214786
R25610 DVDD.n503 DVDD.n501 0.214786
R25611 DVDD.n547 DVDD.n504 0.214786
R25612 DVDD.n546 DVDD.n505 0.214786
R25613 DVDD.n545 DVDD.n506 0.214786
R25614 DVDD.n508 DVDD.n507 0.214786
R25615 DVDD.n541 DVDD.n509 0.214786
R25616 DVDD.n540 DVDD.n510 0.214786
R25617 DVDD.n539 DVDD.n511 0.214786
R25618 DVDD.n538 DVDD.n512 0.214786
R25619 DVDD.n515 DVDD.n513 0.214786
R25620 DVDD.n534 DVDD.n516 0.214786
R25621 DVDD.n533 DVDD.n517 0.214786
R25622 DVDD.n532 DVDD.n518 0.214786
R25623 DVDD.n521 DVDD.n519 0.214786
R25624 DVDD.n528 DVDD.n522 0.214786
R25625 DVDD.n527 DVDD.n523 0.214786
R25626 DVDD.n526 DVDD.n524 0.214786
R25627 DVDD.n37 DVDD.n36 0.214786
R25628 DVDD.n5943 DVDD.n5942 0.214786
R25629 DVDD.n5945 DVDD.n33 0.214786
R25630 DVDD.n5952 DVDD.n5946 0.214786
R25631 DVDD.n5951 DVDD.n5947 0.214786
R25632 DVDD.n5949 DVDD.n5948 0.214786
R25633 DVDD.n6 DVDD.n5 0.214786
R25634 DVDD.n5960 DVDD.n5959 0.214786
R25635 DVDD.n5961 DVDD.n4 0.214786
R25636 DVDD.n5964 DVDD.n5963 0.214786
R25637 DVDD.n5962 DVDD.n2 0.214786
R25638 DVDD.n5968 DVDD.n1 0.214786
R25639 DVDD.n5970 DVDD.n5969 0.214786
R25640 DVDD.n5972 DVDD.n5971 0.214786
R25641 DVDD.n1107 DVDD.n1106 0.214786
R25642 DVDD.n4419 DVDD.n4418 0.214786
R25643 DVDD.n4420 DVDD.n1105 0.214786
R25644 DVDD.n4422 DVDD.n4421 0.214786
R25645 DVDD.n1103 DVDD.n1102 0.214786
R25646 DVDD.n4427 DVDD.n4426 0.214786
R25647 DVDD.n4428 DVDD.n1101 0.214786
R25648 DVDD.n4430 DVDD.n4429 0.214786
R25649 DVDD.n1099 DVDD.n1098 0.214786
R25650 DVDD.n4435 DVDD.n4434 0.214786
R25651 DVDD.n4436 DVDD.n1097 0.214786
R25652 DVDD.n4438 DVDD.n4437 0.214786
R25653 DVDD.n4439 DVDD.n1096 0.214786
R25654 DVDD.n4441 DVDD.n4440 0.214786
R25655 DVDD.n4444 DVDD.n4443 0.214786
R25656 DVDD.n4448 DVDD.n4447 0.214786
R25657 DVDD.n4449 DVDD.n1093 0.214786
R25658 DVDD.n4451 DVDD.n4450 0.214786
R25659 DVDD.n1091 DVDD.n1090 0.214786
R25660 DVDD.n4456 DVDD.n4455 0.214786
R25661 DVDD.n4457 DVDD.n1089 0.214786
R25662 DVDD.n4459 DVDD.n4458 0.214786
R25663 DVDD.n1087 DVDD.n1086 0.214786
R25664 DVDD.n4464 DVDD.n4463 0.214786
R25665 DVDD.n4465 DVDD.n1085 0.214786
R25666 DVDD.n4498 DVDD.n4466 0.214786
R25667 DVDD.n4497 DVDD.n4467 0.214786
R25668 DVDD.n4470 DVDD.n4468 0.214786
R25669 DVDD.n4493 DVDD.n4471 0.214786
R25670 DVDD.n4492 DVDD.n4472 0.214786
R25671 DVDD.n4491 DVDD.n4473 0.214786
R25672 DVDD.n4476 DVDD.n4474 0.214786
R25673 DVDD.n4487 DVDD.n4477 0.214786
R25674 DVDD.n4486 DVDD.n4478 0.214786
R25675 DVDD.n4485 DVDD.n4479 0.214786
R25676 DVDD.n4481 DVDD.n4480 0.214786
R25677 DVDD.n701 DVDD.n700 0.214786
R25678 DVDD.n4884 DVDD.n4883 0.214786
R25679 DVDD.n4887 DVDD.n4886 0.214786
R25680 DVDD.n694 DVDD.n693 0.214786
R25681 DVDD.n4892 DVDD.n4891 0.214786
R25682 DVDD.n4893 DVDD.n692 0.214786
R25683 DVDD.n4895 DVDD.n4894 0.214786
R25684 DVDD.n690 DVDD.n689 0.214786
R25685 DVDD.n4900 DVDD.n4899 0.214786
R25686 DVDD.n4901 DVDD.n688 0.214786
R25687 DVDD.n4903 DVDD.n4902 0.214786
R25688 DVDD.n686 DVDD.n685 0.214786
R25689 DVDD.n4908 DVDD.n4907 0.214786
R25690 DVDD.n4909 DVDD.n684 0.214786
R25691 DVDD.n4939 DVDD.n4910 0.214786
R25692 DVDD.n4938 DVDD.n4911 0.214786
R25693 DVDD.n4914 DVDD.n4912 0.214786
R25694 DVDD.n4934 DVDD.n4915 0.214786
R25695 DVDD.n4933 DVDD.n4916 0.214786
R25696 DVDD.n4932 DVDD.n4917 0.214786
R25697 DVDD.n4920 DVDD.n4918 0.214786
R25698 DVDD.n4928 DVDD.n4921 0.214786
R25699 DVDD.n4927 DVDD.n4922 0.214786
R25700 DVDD.n4926 DVDD.n4923 0.214786
R25701 DVDD.n480 DVDD.n479 0.214786
R25702 DVDD.n5250 DVDD.n5249 0.214786
R25703 DVDD.n5252 DVDD.n476 0.214786
R25704 DVDD.n5316 DVDD.n5253 0.214786
R25705 DVDD.n5315 DVDD.n5254 0.214786
R25706 DVDD.n5314 DVDD.n5255 0.214786
R25707 DVDD.n5258 DVDD.n5256 0.214786
R25708 DVDD.n5310 DVDD.n5259 0.214786
R25709 DVDD.n5309 DVDD.n5260 0.214786
R25710 DVDD.n5308 DVDD.n5261 0.214786
R25711 DVDD.n5264 DVDD.n5262 0.214786
R25712 DVDD.n5304 DVDD.n5265 0.214786
R25713 DVDD.n5303 DVDD.n5266 0.214786
R25714 DVDD.n5302 DVDD.n5267 0.214786
R25715 DVDD.n5300 DVDD.n5268 0.214786
R25716 DVDD.n5299 DVDD.n5269 0.214786
R25717 DVDD.n5298 DVDD.n5270 0.214786
R25718 DVDD.n5273 DVDD.n5271 0.214786
R25719 DVDD.n5294 DVDD.n5274 0.214786
R25720 DVDD.n5293 DVDD.n5275 0.214786
R25721 DVDD.n5292 DVDD.n5276 0.214786
R25722 DVDD.n5279 DVDD.n5277 0.214786
R25723 DVDD.n5288 DVDD.n5280 0.214786
R25724 DVDD.n5287 DVDD.n5281 0.214786
R25725 DVDD.n5286 DVDD.n5282 0.214786
R25726 DVDD.n5284 DVDD.n5283 0.214786
R25727 DVDD.n5937 DVDD.n45 0.214786
R25728 DVDD.n5936 DVDD.n46 0.214786
R25729 DVDD.n5579 DVDD.n47 0.214786
R25730 DVDD.n5580 DVDD.n5578 0.214786
R25731 DVDD.n5602 DVDD.n5581 0.214786
R25732 DVDD.n5601 DVDD.n5582 0.214786
R25733 DVDD.n5600 DVDD.n5583 0.214786
R25734 DVDD.n5586 DVDD.n5584 0.214786
R25735 DVDD.n5596 DVDD.n5587 0.214786
R25736 DVDD.n5595 DVDD.n5588 0.214786
R25737 DVDD.n5594 DVDD.n5589 0.214786
R25738 DVDD.n5591 DVDD.n5590 0.214786
R25739 DVDD.n5897 DVDD.n5896 0.214786
R25740 DVDD.n5900 DVDD.n5895 0.214786
R25741 DVDD.n5901 DVDD.n5894 0.214786
R25742 DVDD.n5902 DVDD.n5893 0.214786
R25743 DVDD.n5892 DVDD.n5890 0.214786
R25744 DVDD.n5906 DVDD.n5889 0.214786
R25745 DVDD.n5907 DVDD.n5888 0.214786
R25746 DVDD.n5908 DVDD.n5887 0.214786
R25747 DVDD.n5886 DVDD.n117 0.214786
R25748 DVDD.n5885 DVDD.n5884 0.214786
R25749 DVDD.n5882 DVDD.n118 0.214786
R25750 DVDD.n5881 DVDD.n5880 0.214786
R25751 DVDD.n5878 DVDD.n5877 0.214786
R25752 DVDD.n121 DVDD.n120 0.214786
R25753 DVDD.n5873 DVDD.n5872 0.214786
R25754 DVDD.n5871 DVDD.n123 0.214786
R25755 DVDD.n5870 DVDD.n5869 0.214786
R25756 DVDD.n125 DVDD.n124 0.214786
R25757 DVDD.n5865 DVDD.n5864 0.214786
R25758 DVDD.n5863 DVDD.n127 0.214786
R25759 DVDD.n5862 DVDD.n5861 0.214786
R25760 DVDD.n129 DVDD.n128 0.214786
R25761 DVDD.n5857 DVDD.n5856 0.214786
R25762 DVDD.n5855 DVDD.n131 0.214786
R25763 DVDD.n5854 DVDD.n5853 0.214786
R25764 DVDD.n133 DVDD.n132 0.214786
R25765 DVDD.n5122 DVDD.n5121 0.214786
R25766 DVDD.n5120 DVDD.n5119 0.214786
R25767 DVDD.n5126 DVDD.n5118 0.214786
R25768 DVDD.n5127 DVDD.n5117 0.214786
R25769 DVDD.n5128 DVDD.n5116 0.214786
R25770 DVDD.n5115 DVDD.n5113 0.214786
R25771 DVDD.n5132 DVDD.n5112 0.214786
R25772 DVDD.n5133 DVDD.n5111 0.214786
R25773 DVDD.n5134 DVDD.n5110 0.214786
R25774 DVDD.n5109 DVDD.n5108 0.214786
R25775 DVDD.n5324 DVDD.n447 0.214786
R25776 DVDD.n5325 DVDD.n446 0.214786
R25777 DVDD.n5326 DVDD.n445 0.214786
R25778 DVDD.n444 DVDD.n442 0.214786
R25779 DVDD.n5330 DVDD.n441 0.214786
R25780 DVDD.n5331 DVDD.n440 0.214786
R25781 DVDD.n5332 DVDD.n439 0.214786
R25782 DVDD.n438 DVDD.n436 0.214786
R25783 DVDD.n5336 DVDD.n435 0.214786
R25784 DVDD.n5337 DVDD.n434 0.214786
R25785 DVDD.n5338 DVDD.n433 0.214786
R25786 DVDD.n432 DVDD.n430 0.214786
R25787 DVDD.n431 DVDD.n423 0.214786
R25788 DVDD.n5345 DVDD.n422 0.214786
R25789 DVDD.n5346 DVDD.n421 0.214786
R25790 DVDD.n5347 DVDD.n420 0.214786
R25791 DVDD.n419 DVDD.n417 0.214786
R25792 DVDD.n5351 DVDD.n416 0.214786
R25793 DVDD.n5352 DVDD.n415 0.214786
R25794 DVDD.n5353 DVDD.n414 0.214786
R25795 DVDD.n413 DVDD.n411 0.214786
R25796 DVDD.n5357 DVDD.n410 0.214786
R25797 DVDD.n5358 DVDD.n409 0.214786
R25798 DVDD.n5359 DVDD.n408 0.214786
R25799 DVDD.n698 DVDD.n399 0.214786
R25800 DVDD.n5365 DVDD.n398 0.214786
R25801 DVDD.n5366 DVDD.n397 0.214786
R25802 DVDD.n5367 DVDD.n396 0.214786
R25803 DVDD.n395 DVDD.n393 0.214786
R25804 DVDD.n5371 DVDD.n392 0.214786
R25805 DVDD.n5372 DVDD.n391 0.214786
R25806 DVDD.n5373 DVDD.n390 0.214786
R25807 DVDD.n389 DVDD.n387 0.214786
R25808 DVDD.n5377 DVDD.n386 0.214786
R25809 DVDD.n5378 DVDD.n385 0.214786
R25810 DVDD.n5379 DVDD.n384 0.214786
R25811 DVDD.n383 DVDD.n376 0.214786
R25812 DVDD.n5385 DVDD.n375 0.214786
R25813 DVDD.n5386 DVDD.n374 0.214786
R25814 DVDD.n5387 DVDD.n373 0.214786
R25815 DVDD.n372 DVDD.n370 0.214786
R25816 DVDD.n5391 DVDD.n369 0.214786
R25817 DVDD.n5392 DVDD.n368 0.214786
R25818 DVDD.n5393 DVDD.n367 0.214786
R25819 DVDD.n366 DVDD.n364 0.214786
R25820 DVDD.n5397 DVDD.n363 0.214786
R25821 DVDD.n5398 DVDD.n362 0.214786
R25822 DVDD.n5399 DVDD.n361 0.214786
R25823 DVDD.n5403 DVDD.n357 0.214786
R25824 DVDD.n1179 DVDD.n1151 0.214786
R25825 DVDD.n1178 DVDD.n1152 0.214786
R25826 DVDD.n1177 DVDD.n1153 0.214786
R25827 DVDD.n1156 DVDD.n1154 0.214786
R25828 DVDD.n1173 DVDD.n1157 0.214786
R25829 DVDD.n1172 DVDD.n1158 0.214786
R25830 DVDD.n1171 DVDD.n1159 0.214786
R25831 DVDD.n1162 DVDD.n1160 0.214786
R25832 DVDD.n1167 DVDD.n1163 0.214786
R25833 DVDD.n1166 DVDD.n1165 0.214786
R25834 DVDD.n1164 DVDD.n354 0.214786
R25835 DVDD.n5406 DVDD.n355 0.214786
R25836 DVDD.n5405 DVDD.n356 0.214786
R25837 DVDD.n3405 DVDD.n3404 0.214786
R25838 DVDD.n2724 DVDD.n2723 0.214786
R25839 DVDD.n3412 DVDD.n3411 0.214786
R25840 DVDD.n2721 DVDD.n2706 0.214786
R25841 DVDD.n3417 DVDD.n3416 0.214786
R25842 DVDD.n3425 DVDD.n3424 0.214786
R25843 DVDD.n2704 DVDD.n2699 0.214786
R25844 DVDD.n3431 DVDD.n3430 0.214786
R25845 DVDD.n2700 DVDD.n2696 0.214786
R25846 DVDD.n3435 DVDD.n2695 0.214786
R25847 DVDD.n3437 DVDD.n3436 0.214786
R25848 DVDD.n2691 DVDD.n2689 0.214786
R25849 DVDD.n3443 DVDD.n3442 0.214786
R25850 DVDD.n2693 DVDD.n2690 0.214786
R25851 DVDD.n2692 DVDD.n1915 0.214786
R25852 DVDD.n1940 DVDD.n1914 0.214786
R25853 DVDD.n1942 DVDD.n1941 0.214786
R25854 DVDD.n1943 DVDD.n1938 0.214786
R25855 DVDD.n3400 DVDD.n3399 0.214786
R25856 DVDD.n3394 DVDD.n2728 0.214786
R25857 DVDD.n3393 DVDD.n3392 0.214786
R25858 DVDD.n2965 DVDD.n2733 0.214786
R25859 DVDD.n2969 DVDD.n2964 0.214786
R25860 DVDD.n2980 DVDD.n2979 0.214786
R25861 DVDD.n2971 DVDD.n2968 0.214786
R25862 DVDD.n2975 DVDD.n2974 0.214786
R25863 DVDD.n3401 DVDD.n3400 0.214786
R25864 DVDD.n2728 DVDD.n2727 0.214786
R25865 DVDD.n3392 DVDD.n3391 0.214786
R25866 DVDD.n3390 DVDD.n2733 0.214786
R25867 DVDD.n2969 DVDD.n2739 0.214786
R25868 DVDD.n2979 DVDD.n2978 0.214786
R25869 DVDD.n2977 DVDD.n2968 0.214786
R25870 DVDD.n3404 DVDD.n3403 0.214786
R25871 DVDD.n2723 DVDD.n2722 0.214786
R25872 DVDD.n3413 DVDD.n3412 0.214786
R25873 DVDD.n3414 DVDD.n2721 0.214786
R25874 DVDD.n3416 DVDD.n3415 0.214786
R25875 DVDD.n3426 DVDD.n3425 0.214786
R25876 DVDD.n3427 DVDD.n2699 0.214786
R25877 DVDD.n3430 DVDD.n3429 0.214786
R25878 DVDD.n3428 DVDD.n2700 0.214786
R25879 DVDD.n2695 DVDD.n2694 0.214786
R25880 DVDD.n3438 DVDD.n3437 0.214786
R25881 DVDD.n3439 DVDD.n2691 0.214786
R25882 DVDD.n3442 DVDD.n3441 0.214786
R25883 DVDD.n3440 DVDD.n2693 0.214786
R25884 DVDD.n2692 DVDD.n1900 0.214786
R25885 DVDD.n1940 DVDD.n1899 0.214786
R25886 DVDD.n1942 DVDD.n1939 0.214786
R25887 DVDD.n3402 DVDD.n2726 0.214786
R25888 DVDD.n2730 DVDD.n2726 0.214786
R25889 DVDD.n3265 DVDD.n3264 0.214786
R25890 DVDD.n2961 DVDD.n2960 0.214786
R25891 DVDD.n3259 DVDD.n3258 0.214786
R25892 DVDD.n3257 DVDD.n2743 0.214786
R25893 DVDD.n3101 DVDD.n2744 0.214786
R25894 DVDD.n3102 DVDD.n3100 0.214786
R25895 DVDD.n3103 DVDD.n3099 0.214786
R25896 DVDD.n3268 DVDD.n3267 0.214786
R25897 DVDD.n2930 DVDD.n2929 0.214786
R25898 DVDD.n3285 DVDD.n3284 0.214786
R25899 DVDD.n3286 DVDD.n2928 0.214786
R25900 DVDD.n3288 DVDD.n3287 0.214786
R25901 DVDD.n2922 DVDD.n2921 0.214786
R25902 DVDD.n3305 DVDD.n3304 0.214786
R25903 DVDD.n3306 DVDD.n2920 0.214786
R25904 DVDD.n3322 DVDD.n3307 0.214786
R25905 DVDD.n3321 DVDD.n3308 0.214786
R25906 DVDD.n3319 DVDD.n3309 0.214786
R25907 DVDD.n3318 DVDD.n3310 0.214786
R25908 DVDD.n3317 DVDD.n3311 0.214786
R25909 DVDD.n3314 DVDD.n3312 0.214786
R25910 DVDD.n3313 DVDD.n1904 0.214786
R25911 DVDD.n1952 DVDD.n1903 0.214786
R25912 DVDD.n1951 DVDD.n1919 0.214786
R25913 DVDD.n3266 DVDD.n2959 0.214786
R25914 DVDD.n3269 DVDD.n3268 0.214786
R25915 DVDD.n3270 DVDD.n2930 0.214786
R25916 DVDD.n3284 DVDD.n3283 0.214786
R25917 DVDD.n2928 DVDD.n2927 0.214786
R25918 DVDD.n3289 DVDD.n3288 0.214786
R25919 DVDD.n3293 DVDD.n2922 0.214786
R25920 DVDD.n3304 DVDD.n3303 0.214786
R25921 DVDD.n2920 DVDD.n2918 0.214786
R25922 DVDD.n3323 DVDD.n3322 0.214786
R25923 DVDD.n3321 DVDD.n3320 0.214786
R25924 DVDD.n3319 DVDD.n2862 0.214786
R25925 DVDD.n3318 DVDD.n2872 0.214786
R25926 DVDD.n3317 DVDD.n3316 0.214786
R25927 DVDD.n3315 DVDD.n3314 0.214786
R25928 DVDD.n3313 DVDD.n1917 0.214786
R25929 DVDD.n1953 DVDD.n1952 0.214786
R25930 DVDD.n1951 DVDD.n1918 0.214786
R25931 DVDD.n1950 DVDD.n1949 0.214786
R25932 DVDD.n3264 DVDD.n3263 0.214786
R25933 DVDD.n3261 DVDD.n2961 0.214786
R25934 DVDD.n3260 DVDD.n3259 0.214786
R25935 DVDD.n3105 DVDD.n3104 0.214786
R25936 DVDD.n3103 DVDD.n3092 0.214786
R25937 DVDD.n3102 DVDD.n3089 0.214786
R25938 DVDD.n3101 DVDD.n3081 0.214786
R25939 DVDD.n3257 DVDD.n3256 0.214786
R25940 DVDD.n3262 DVDD.n2959 0.214786
R25941 DVDD.n3380 DVDD.n2758 0.214786
R25942 DVDD.n3379 DVDD.n2759 0.214786
R25943 DVDD.n2946 DVDD.n2760 0.214786
R25944 DVDD.n3375 DVDD.n2762 0.214786
R25945 DVDD.n3374 DVDD.n3373 0.214786
R25946 DVDD.n2771 DVDD.n2769 0.214786
R25947 DVDD.n3364 DVDD.n3363 0.214786
R25948 DVDD.n2807 DVDD.n2772 0.214786
R25949 DVDD.n3359 DVDD.n2775 0.214786
R25950 DVDD.n3358 DVDD.n2776 0.214786
R25951 DVDD.n3357 DVDD.n2777 0.214786
R25952 DVDD.n2780 DVDD.n2778 0.214786
R25953 DVDD.n3353 DVDD.n3349 0.214786
R25954 DVDD.n3352 DVDD.n3350 0.214786
R25955 DVDD.n3351 DVDD.n1973 0.214786
R25956 DVDD.n1972 DVDD.n1971 0.214786
R25957 DVDD.n1970 DVDD.n1955 0.214786
R25958 DVDD.n1957 DVDD.n1956 0.214786
R25959 DVDD.n2756 DVDD.n2754 0.214786
R25960 DVDD.n3385 DVDD.n2753 0.214786
R25961 DVDD.n3386 DVDD.n2752 0.214786
R25962 DVDD.n3156 DVDD.n3136 0.214786
R25963 DVDD.n3160 DVDD.n3137 0.214786
R25964 DVDD.n3159 DVDD.n3126 0.214786
R25965 DVDD.n3158 DVDD.n3127 0.214786
R25966 DVDD.n3387 DVDD.n2751 0.214786
R25967 DVDD.n3381 DVDD.n2757 0.214786
R25968 DVDD.n3383 DVDD.n2754 0.214786
R25969 DVDD.n3385 DVDD.n3384 0.214786
R25970 DVDD.n3386 DVDD.n2749 0.214786
R25971 DVDD.n3388 DVDD.n3387 0.214786
R25972 DVDD.n3158 DVDD.n2748 0.214786
R25973 DVDD.n3159 DVDD.n3157 0.214786
R25974 DVDD.n3161 DVDD.n3160 0.214786
R25975 DVDD.n3380 DVDD.n2755 0.214786
R25976 DVDD.n3379 DVDD.n3378 0.214786
R25977 DVDD.n3377 DVDD.n2760 0.214786
R25978 DVDD.n3376 DVDD.n3375 0.214786
R25979 DVDD.n3374 DVDD.n2761 0.214786
R25980 DVDD.n2773 DVDD.n2771 0.214786
R25981 DVDD.n3363 DVDD.n3362 0.214786
R25982 DVDD.n3361 DVDD.n2772 0.214786
R25983 DVDD.n3360 DVDD.n3359 0.214786
R25984 DVDD.n3358 DVDD.n2774 0.214786
R25985 DVDD.n3357 DVDD.n3356 0.214786
R25986 DVDD.n3355 DVDD.n2778 0.214786
R25987 DVDD.n3354 DVDD.n3353 0.214786
R25988 DVDD.n3352 DVDD.n2779 0.214786
R25989 DVDD.n3351 DVDD.n1908 0.214786
R25990 DVDD.n1971 DVDD.n1907 0.214786
R25991 DVDD.n1970 DVDD.n1969 0.214786
R25992 DVDD.n3382 DVDD.n3381 0.214786
R25993 DVDD.n2992 DVDD.n2990 0.214786
R25994 DVDD.n3074 DVDD.n2989 0.214786
R25995 DVDD.n3075 DVDD.n2988 0.214786
R25996 DVDD.n3076 DVDD.n2737 0.214786
R25997 DVDD.n3069 DVDD.n2994 0.214786
R25998 DVDD.n3002 DVDD.n2995 0.214786
R25999 DVDD.n3058 DVDD.n3003 0.214786
R26000 DVDD.n3057 DVDD.n3004 0.214786
R26001 DVDD.n3006 DVDD.n3005 0.214786
R26002 DVDD.n3050 DVDD.n3012 0.214786
R26003 DVDD.n3049 DVDD.n3013 0.214786
R26004 DVDD.n3021 DVDD.n3014 0.214786
R26005 DVDD.n3038 DVDD.n3022 0.214786
R26006 DVDD.n3037 DVDD.n3023 0.214786
R26007 DVDD.n3036 DVDD.n3024 0.214786
R26008 DVDD.n3027 DVDD.n3025 0.214786
R26009 DVDD.n3032 DVDD.n3028 0.214786
R26010 DVDD.n3031 DVDD.n3029 0.214786
R26011 DVDD.n3030 DVDD.n1911 0.214786
R26012 DVDD.n3706 DVDD.n3705 0.214786
R26013 DVDD.n1913 DVDD.n1912 0.214786
R26014 DVDD.n3070 DVDD.n2993 0.214786
R26015 DVDD.n3069 DVDD.n3068 0.214786
R26016 DVDD.n2996 DVDD.n2995 0.214786
R26017 DVDD.n3059 DVDD.n3058 0.214786
R26018 DVDD.n3057 DVDD.n3056 0.214786
R26019 DVDD.n3008 DVDD.n3006 0.214786
R26020 DVDD.n3051 DVDD.n3050 0.214786
R26021 DVDD.n3049 DVDD.n3048 0.214786
R26022 DVDD.n3019 DVDD.n3014 0.214786
R26023 DVDD.n3039 DVDD.n3038 0.214786
R26024 DVDD.n3037 DVDD.n3020 0.214786
R26025 DVDD.n3036 DVDD.n3035 0.214786
R26026 DVDD.n3034 DVDD.n3025 0.214786
R26027 DVDD.n3033 DVDD.n3032 0.214786
R26028 DVDD.n3031 DVDD.n3026 0.214786
R26029 DVDD.n3030 DVDD.n1974 0.214786
R26030 DVDD.n3705 DVDD.n3704 0.214786
R26031 DVDD.n3703 DVDD.n1913 0.214786
R26032 DVDD.n3702 DVDD.n3701 0.214786
R26033 DVDD.n3072 DVDD.n2990 0.214786
R26034 DVDD.n3074 DVDD.n3073 0.214786
R26035 DVDD.n3075 DVDD.n2987 0.214786
R26036 DVDD.n3077 DVDD.n3076 0.214786
R26037 DVDD.n3071 DVDD.n3070 0.214786
R26038 DVDD.n4197 DVDD.n4195 0.214786
R26039 DVDD.n4194 DVDD.n4193 0.214786
R26040 DVDD.n4192 DVDD.n4188 0.214786
R26041 DVDD.n4209 DVDD.n4187 0.214786
R26042 DVDD.n4210 DVDD.n4186 0.214786
R26043 DVDD.n4211 DVDD.n4185 0.214786
R26044 DVDD.n4184 DVDD.n4182 0.214786
R26045 DVDD.n4215 DVDD.n4181 0.214786
R26046 DVDD.n4216 DVDD.n4180 0.214786
R26047 DVDD.n4217 DVDD.n4179 0.214786
R26048 DVDD.n4174 DVDD.n4173 0.214786
R26049 DVDD.n4222 DVDD.n4221 0.214786
R26050 DVDD.n4172 DVDD.n4171 0.214786
R26051 DVDD.n1768 DVDD.n1767 0.214786
R26052 DVDD.n4167 DVDD.n4166 0.214786
R26053 DVDD.n4165 DVDD.n1770 0.214786
R26054 DVDD.n4164 DVDD.n4163 0.214786
R26055 DVDD.n1772 DVDD.n1771 0.214786
R26056 DVDD.n4157 DVDD.n4156 0.214786
R26057 DVDD.n4155 DVDD.n1774 0.214786
R26058 DVDD.n4154 DVDD.n4153 0.214786
R26059 DVDD.n1776 DVDD.n1775 0.214786
R26060 DVDD.n4147 DVDD.n4146 0.214786
R26061 DVDD.n4145 DVDD.n1777 0.214786
R26062 DVDD.n4144 DVDD.n4143 0.214786
R26063 DVDD.n1779 DVDD.n1778 0.214786
R26064 DVDD.n4135 DVDD.n4134 0.214786
R26065 DVDD.n4133 DVDD.n1781 0.214786
R26066 DVDD.n4132 DVDD.n4131 0.214786
R26067 DVDD.n1783 DVDD.n1782 0.214786
R26068 DVDD.n4112 DVDD.n4111 0.214786
R26069 DVDD.n4110 DVDD.n4109 0.214786
R26070 DVDD.n4117 DVDD.n4108 0.214786
R26071 DVDD.n4118 DVDD.n4107 0.214786
R26072 DVDD.n4119 DVDD.n4106 0.214786
R26073 DVDD.n4105 DVDD.n1788 0.214786
R26074 DVDD.n4033 DVDD.n1789 0.214786
R26075 DVDD.n4032 DVDD.n4031 0.214786
R26076 DVDD.n4030 DVDD.n1796 0.214786
R26077 DVDD.n4029 DVDD.n4028 0.214786
R26078 DVDD.n1798 DVDD.n1797 0.214786
R26079 DVDD.n4023 DVDD.n4022 0.214786
R26080 DVDD.n4021 DVDD.n1800 0.214786
R26081 DVDD.n4020 DVDD.n4019 0.214786
R26082 DVDD.n1802 DVDD.n1801 0.214786
R26083 DVDD.n4011 DVDD.n4010 0.214786
R26084 DVDD.n4009 DVDD.n1804 0.214786
R26085 DVDD.n4008 DVDD.n4007 0.214786
R26086 DVDD.n1806 DVDD.n1805 0.214786
R26087 DVDD.n4003 DVDD.n4002 0.214786
R26088 DVDD.n4001 DVDD.n1808 0.214786
R26089 DVDD.n4000 DVDD.n3999 0.214786
R26090 DVDD.n1810 DVDD.n1809 0.214786
R26091 DVDD.n3991 DVDD.n3990 0.214786
R26092 DVDD.n3989 DVDD.n1812 0.214786
R26093 DVDD.n3988 DVDD.n3987 0.214786
R26094 DVDD.n1814 DVDD.n1813 0.214786
R26095 DVDD.n3983 DVDD.n3982 0.214786
R26096 DVDD.n3981 DVDD.n1816 0.214786
R26097 DVDD.n3980 DVDD.n3979 0.214786
R26098 DVDD.n3975 DVDD.n3974 0.214786
R26099 DVDD.n3973 DVDD.n3926 0.214786
R26100 DVDD.n3972 DVDD.n3971 0.214786
R26101 DVDD.n3928 DVDD.n3927 0.214786
R26102 DVDD.n3949 DVDD.n3948 0.214786
R26103 DVDD.n3950 DVDD.n3947 0.214786
R26104 DVDD.n3951 DVDD.n3946 0.214786
R26105 DVDD.n3945 DVDD.n3943 0.214786
R26106 DVDD.n3956 DVDD.n3942 0.214786
R26107 DVDD.n3957 DVDD.n3941 0.214786
R26108 DVDD.n3958 DVDD.n3940 0.214786
R26109 DVDD.n3939 DVDD.n3937 0.214786
R26110 DVDD.n3734 DVDD.n3733 0.214786
R26111 DVDD.n1855 DVDD.n1854 0.214786
R26112 DVDD.n3784 DVDD.n3783 0.214786
R26113 DVDD.n3785 DVDD.n1853 0.214786
R26114 DVDD.n3787 DVDD.n3786 0.214786
R26115 DVDD.n1851 DVDD.n1850 0.214786
R26116 DVDD.n3792 DVDD.n3791 0.214786
R26117 DVDD.n3793 DVDD.n1849 0.214786
R26118 DVDD.n3795 DVDD.n3794 0.214786
R26119 DVDD.n1847 DVDD.n1846 0.214786
R26120 DVDD.n3801 DVDD.n3800 0.214786
R26121 DVDD.n3802 DVDD.n1845 0.214786
R26122 DVDD.n3804 DVDD.n3803 0.214786
R26123 DVDD.n3805 DVDD.n1687 0.214786
R26124 DVDD.n4259 DVDD.n4258 0.214786
R26125 DVDD.n1689 DVDD.n1688 0.214786
R26126 DVDD.n4254 DVDD.n1692 0.214786
R26127 DVDD.n4253 DVDD.n1693 0.214786
R26128 DVDD.n1696 DVDD.n1694 0.214786
R26129 DVDD.n4249 DVDD.n1697 0.214786
R26130 DVDD.n4248 DVDD.n1698 0.214786
R26131 DVDD.n1701 DVDD.n1699 0.214786
R26132 DVDD.n4244 DVDD.n1702 0.214786
R26133 DVDD.n4243 DVDD.n1703 0.214786
R26134 DVDD.n4242 DVDD.n1704 0.214786
R26135 DVDD.n3938 DVDD.n1705 0.214786
R26136 DVDD.n4193 DVDD.n4189 0.214786
R26137 DVDD.n4197 DVDD.n4196 0.214786
R26138 DVDD.n4198 DVDD.n4191 0.214786
R26139 DVDD.n4207 DVDD.n4188 0.214786
R26140 DVDD.n4209 DVDD.n4208 0.214786
R26141 DVDD.n4210 DVDD.n4183 0.214786
R26142 DVDD.n4212 DVDD.n4211 0.214786
R26143 DVDD.n4213 DVDD.n4182 0.214786
R26144 DVDD.n4215 DVDD.n4214 0.214786
R26145 DVDD.n4216 DVDD.n4178 0.214786
R26146 DVDD.n4218 DVDD.n4217 0.214786
R26147 DVDD.n4219 DVDD.n4174 0.214786
R26148 DVDD.n4221 DVDD.n4220 0.214786
R26149 DVDD.n4171 DVDD.n4170 0.214786
R26150 DVDD.n4169 DVDD.n1768 0.214786
R26151 DVDD.n4168 DVDD.n4167 0.214786
R26152 DVDD.n4161 DVDD.n1770 0.214786
R26153 DVDD.n4163 DVDD.n4162 0.214786
R26154 DVDD.n4160 DVDD.n1772 0.214786
R26155 DVDD.n4158 DVDD.n4157 0.214786
R26156 DVDD.n1774 DVDD.n1773 0.214786
R26157 DVDD.n4153 DVDD.n4152 0.214786
R26158 DVDD.n4151 DVDD.n1776 0.214786
R26159 DVDD.n4148 DVDD.n4147 0.214786
R26160 DVDD.n4141 DVDD.n1777 0.214786
R26161 DVDD.n4143 DVDD.n4142 0.214786
R26162 DVDD.n4137 DVDD.n1779 0.214786
R26163 DVDD.n4136 DVDD.n4135 0.214786
R26164 DVDD.n1781 DVDD.n1780 0.214786
R26165 DVDD.n4131 DVDD.n4130 0.214786
R26166 DVDD.n1784 DVDD.n1783 0.214786
R26167 DVDD.n4113 DVDD.n4112 0.214786
R26168 DVDD.n4114 DVDD.n4109 0.214786
R26169 DVDD.n4117 DVDD.n4116 0.214786
R26170 DVDD.n4118 DVDD.n1787 0.214786
R26171 DVDD.n4120 DVDD.n4119 0.214786
R26172 DVDD.n1788 DVDD.n1786 0.214786
R26173 DVDD.n4034 DVDD.n4033 0.214786
R26174 DVDD.n4032 DVDD.n1795 0.214786
R26175 DVDD.n4026 DVDD.n1796 0.214786
R26176 DVDD.n4028 DVDD.n4027 0.214786
R26177 DVDD.n4025 DVDD.n1798 0.214786
R26178 DVDD.n4024 DVDD.n4023 0.214786
R26179 DVDD.n1800 DVDD.n1799 0.214786
R26180 DVDD.n4019 DVDD.n4018 0.214786
R26181 DVDD.n4017 DVDD.n1802 0.214786
R26182 DVDD.n4012 DVDD.n4011 0.214786
R26183 DVDD.n1804 DVDD.n1803 0.214786
R26184 DVDD.n4007 DVDD.n4006 0.214786
R26185 DVDD.n4005 DVDD.n1806 0.214786
R26186 DVDD.n4004 DVDD.n4003 0.214786
R26187 DVDD.n1808 DVDD.n1807 0.214786
R26188 DVDD.n3999 DVDD.n3998 0.214786
R26189 DVDD.n3993 DVDD.n1810 0.214786
R26190 DVDD.n3992 DVDD.n3991 0.214786
R26191 DVDD.n1812 DVDD.n1811 0.214786
R26192 DVDD.n3987 DVDD.n3986 0.214786
R26193 DVDD.n3985 DVDD.n1814 0.214786
R26194 DVDD.n3984 DVDD.n3983 0.214786
R26195 DVDD.n1816 DVDD.n1815 0.214786
R26196 DVDD.n3979 DVDD.n3978 0.214786
R26197 DVDD.n3976 DVDD.n3975 0.214786
R26198 DVDD.n3969 DVDD.n3926 0.214786
R26199 DVDD.n3971 DVDD.n3970 0.214786
R26200 DVDD.n3968 DVDD.n3928 0.214786
R26201 DVDD.n3949 DVDD.n3929 0.214786
R26202 DVDD.n3950 DVDD.n3944 0.214786
R26203 DVDD.n3952 DVDD.n3951 0.214786
R26204 DVDD.n3953 DVDD.n3943 0.214786
R26205 DVDD.n3956 DVDD.n3955 0.214786
R26206 DVDD.n3957 DVDD.n3936 0.214786
R26207 DVDD.n3959 DVDD.n3958 0.214786
R26208 DVDD.n3937 DVDD.n3935 0.214786
R26209 DVDD.n3736 DVDD.n3735 0.214786
R26210 DVDD.n3734 DVDD.n1856 0.214786
R26211 DVDD.n3780 DVDD.n1855 0.214786
R26212 DVDD.n3783 DVDD.n3782 0.214786
R26213 DVDD.n3781 DVDD.n1853 0.214786
R26214 DVDD.n3788 DVDD.n3787 0.214786
R26215 DVDD.n3789 DVDD.n1851 0.214786
R26216 DVDD.n3791 DVDD.n3790 0.214786
R26217 DVDD.n1849 DVDD.n1848 0.214786
R26218 DVDD.n3796 DVDD.n3795 0.214786
R26219 DVDD.n3797 DVDD.n1847 0.214786
R26220 DVDD.n3800 DVDD.n3799 0.214786
R26221 DVDD.n3798 DVDD.n1845 0.214786
R26222 DVDD.n3804 DVDD.n1844 0.214786
R26223 DVDD.n3806 DVDD.n3805 0.214786
R26224 DVDD.n4258 DVDD.n4257 0.214786
R26225 DVDD.n4256 DVDD.n1689 0.214786
R26226 DVDD.n4255 DVDD.n4254 0.214786
R26227 DVDD.n4253 DVDD.n4252 0.214786
R26228 DVDD.n4251 DVDD.n1694 0.214786
R26229 DVDD.n4250 DVDD.n4249 0.214786
R26230 DVDD.n4248 DVDD.n4247 0.214786
R26231 DVDD.n4246 DVDD.n1699 0.214786
R26232 DVDD.n4245 DVDD.n4244 0.214786
R26233 DVDD.n4243 DVDD.n1700 0.214786
R26234 DVDD.n4242 DVDD.n4241 0.214786
R26235 DVDD.n1707 DVDD.n1705 0.214786
R26236 DVDD.n5900 DVDD.n5899 0.214786
R26237 DVDD.n5901 DVDD.n5891 0.214786
R26238 DVDD.n5903 DVDD.n5902 0.214786
R26239 DVDD.n5904 DVDD.n5890 0.214786
R26240 DVDD.n5906 DVDD.n5905 0.214786
R26241 DVDD.n5907 DVDD.n115 0.214786
R26242 DVDD.n5909 DVDD.n5908 0.214786
R26243 DVDD.n117 DVDD.n116 0.214786
R26244 DVDD.n5884 DVDD.n5883 0.214786
R26245 DVDD.n5882 DVDD.n82 0.214786
R26246 DVDD.n5881 DVDD.n80 0.214786
R26247 DVDD.n5877 DVDD.n5876 0.214786
R26248 DVDD.n5875 DVDD.n121 0.214786
R26249 DVDD.n5874 DVDD.n5873 0.214786
R26250 DVDD.n123 DVDD.n122 0.214786
R26251 DVDD.n5869 DVDD.n5868 0.214786
R26252 DVDD.n5867 DVDD.n125 0.214786
R26253 DVDD.n5866 DVDD.n5865 0.214786
R26254 DVDD.n127 DVDD.n126 0.214786
R26255 DVDD.n5861 DVDD.n5860 0.214786
R26256 DVDD.n5859 DVDD.n129 0.214786
R26257 DVDD.n5858 DVDD.n5857 0.214786
R26258 DVDD.n137 DVDD.n131 0.214786
R26259 DVDD.n5853 DVDD.n5852 0.214786
R26260 DVDD.n134 DVDD.n133 0.214786
R26261 DVDD.n5123 DVDD.n5122 0.214786
R26262 DVDD.n5124 DVDD.n5119 0.214786
R26263 DVDD.n5126 DVDD.n5125 0.214786
R26264 DVDD.n5127 DVDD.n5114 0.214786
R26265 DVDD.n5129 DVDD.n5128 0.214786
R26266 DVDD.n5130 DVDD.n5113 0.214786
R26267 DVDD.n5132 DVDD.n5131 0.214786
R26268 DVDD.n5133 DVDD.n5107 0.214786
R26269 DVDD.n5135 DVDD.n5134 0.214786
R26270 DVDD.n5108 DVDD.n5106 0.214786
R26271 DVDD.n5324 DVDD.n5323 0.214786
R26272 DVDD.n5325 DVDD.n443 0.214786
R26273 DVDD.n5327 DVDD.n5326 0.214786
R26274 DVDD.n5328 DVDD.n442 0.214786
R26275 DVDD.n5330 DVDD.n5329 0.214786
R26276 DVDD.n5331 DVDD.n437 0.214786
R26277 DVDD.n5333 DVDD.n5332 0.214786
R26278 DVDD.n5334 DVDD.n436 0.214786
R26279 DVDD.n5336 DVDD.n5335 0.214786
R26280 DVDD.n5337 DVDD.n429 0.214786
R26281 DVDD.n5339 DVDD.n5338 0.214786
R26282 DVDD.n430 DVDD.n426 0.214786
R26283 DVDD.n5343 DVDD.n423 0.214786
R26284 DVDD.n5345 DVDD.n5344 0.214786
R26285 DVDD.n5346 DVDD.n418 0.214786
R26286 DVDD.n5348 DVDD.n5347 0.214786
R26287 DVDD.n5349 DVDD.n417 0.214786
R26288 DVDD.n5351 DVDD.n5350 0.214786
R26289 DVDD.n5352 DVDD.n412 0.214786
R26290 DVDD.n5354 DVDD.n5353 0.214786
R26291 DVDD.n5355 DVDD.n411 0.214786
R26292 DVDD.n5357 DVDD.n5356 0.214786
R26293 DVDD.n5358 DVDD.n406 0.214786
R26294 DVDD.n5360 DVDD.n5359 0.214786
R26295 DVDD.n402 DVDD.n399 0.214786
R26296 DVDD.n5365 DVDD.n5364 0.214786
R26297 DVDD.n5366 DVDD.n394 0.214786
R26298 DVDD.n5368 DVDD.n5367 0.214786
R26299 DVDD.n5369 DVDD.n393 0.214786
R26300 DVDD.n5371 DVDD.n5370 0.214786
R26301 DVDD.n5372 DVDD.n388 0.214786
R26302 DVDD.n5374 DVDD.n5373 0.214786
R26303 DVDD.n5375 DVDD.n387 0.214786
R26304 DVDD.n5377 DVDD.n5376 0.214786
R26305 DVDD.n5378 DVDD.n382 0.214786
R26306 DVDD.n5380 DVDD.n5379 0.214786
R26307 DVDD.n379 DVDD.n376 0.214786
R26308 DVDD.n5385 DVDD.n5384 0.214786
R26309 DVDD.n5386 DVDD.n371 0.214786
R26310 DVDD.n5388 DVDD.n5387 0.214786
R26311 DVDD.n5389 DVDD.n370 0.214786
R26312 DVDD.n5391 DVDD.n5390 0.214786
R26313 DVDD.n5392 DVDD.n365 0.214786
R26314 DVDD.n5394 DVDD.n5393 0.214786
R26315 DVDD.n5395 DVDD.n364 0.214786
R26316 DVDD.n5397 DVDD.n5396 0.214786
R26317 DVDD.n5398 DVDD.n360 0.214786
R26318 DVDD.n5400 DVDD.n5399 0.214786
R26319 DVDD.n5403 DVDD.n5402 0.214786
R26320 DVDD.n1181 DVDD.n1180 0.214786
R26321 DVDD.n1179 DVDD.n1121 0.214786
R26322 DVDD.n1178 DVDD.n1131 0.214786
R26323 DVDD.n1177 DVDD.n1176 0.214786
R26324 DVDD.n1175 DVDD.n1154 0.214786
R26325 DVDD.n1174 DVDD.n1173 0.214786
R26326 DVDD.n1172 DVDD.n1155 0.214786
R26327 DVDD.n1171 DVDD.n1170 0.214786
R26328 DVDD.n1169 DVDD.n1160 0.214786
R26329 DVDD.n1168 DVDD.n1167 0.214786
R26330 DVDD.n1166 DVDD.n1161 0.214786
R26331 DVDD.n354 DVDD.n328 0.214786
R26332 DVDD.n5407 DVDD.n5406 0.214786
R26333 DVDD.n5405 DVDD.n5404 0.214786
R26334 DVDD.n4412 DVDD.n4411 0.214786
R26335 DVDD.n1108 DVDD.n1107 0.214786
R26336 DVDD.n4418 DVDD.n4417 0.214786
R26337 DVDD.n1105 DVDD.n1104 0.214786
R26338 DVDD.n4423 DVDD.n4422 0.214786
R26339 DVDD.n4424 DVDD.n1103 0.214786
R26340 DVDD.n4426 DVDD.n4425 0.214786
R26341 DVDD.n1101 DVDD.n1100 0.214786
R26342 DVDD.n4431 DVDD.n4430 0.214786
R26343 DVDD.n4432 DVDD.n1099 0.214786
R26344 DVDD.n4434 DVDD.n4433 0.214786
R26345 DVDD.n1097 DVDD.n273 0.214786
R26346 DVDD.n4438 DVDD.n284 0.214786
R26347 DVDD.n4439 DVDD.n297 0.214786
R26348 DVDD.n4440 DVDD.n307 0.214786
R26349 DVDD.n4445 DVDD.n4444 0.214786
R26350 DVDD.n4447 DVDD.n4446 0.214786
R26351 DVDD.n1093 DVDD.n1092 0.214786
R26352 DVDD.n4452 DVDD.n4451 0.214786
R26353 DVDD.n4453 DVDD.n1091 0.214786
R26354 DVDD.n4455 DVDD.n4454 0.214786
R26355 DVDD.n1089 DVDD.n1088 0.214786
R26356 DVDD.n4460 DVDD.n4459 0.214786
R26357 DVDD.n4461 DVDD.n1087 0.214786
R26358 DVDD.n4463 DVDD.n4462 0.214786
R26359 DVDD.n1085 DVDD.n1075 0.214786
R26360 DVDD.n4499 DVDD.n4498 0.214786
R26361 DVDD.n4497 DVDD.n4496 0.214786
R26362 DVDD.n4495 DVDD.n4468 0.214786
R26363 DVDD.n4494 DVDD.n4493 0.214786
R26364 DVDD.n4492 DVDD.n4469 0.214786
R26365 DVDD.n4491 DVDD.n4490 0.214786
R26366 DVDD.n4489 DVDD.n4474 0.214786
R26367 DVDD.n4488 DVDD.n4487 0.214786
R26368 DVDD.n4486 DVDD.n4475 0.214786
R26369 DVDD.n4485 DVDD.n4484 0.214786
R26370 DVDD.n4483 DVDD.n4481 0.214786
R26371 DVDD.n4482 DVDD.n701 0.214786
R26372 DVDD.n4883 DVDD.n4882 0.214786
R26373 DVDD.n4888 DVDD.n4887 0.214786
R26374 DVDD.n4889 DVDD.n694 0.214786
R26375 DVDD.n4891 DVDD.n4890 0.214786
R26376 DVDD.n692 DVDD.n691 0.214786
R26377 DVDD.n4896 DVDD.n4895 0.214786
R26378 DVDD.n4897 DVDD.n690 0.214786
R26379 DVDD.n4899 DVDD.n4898 0.214786
R26380 DVDD.n688 DVDD.n687 0.214786
R26381 DVDD.n4904 DVDD.n4903 0.214786
R26382 DVDD.n4905 DVDD.n686 0.214786
R26383 DVDD.n4907 DVDD.n4906 0.214786
R26384 DVDD.n684 DVDD.n674 0.214786
R26385 DVDD.n4940 DVDD.n4939 0.214786
R26386 DVDD.n4938 DVDD.n4937 0.214786
R26387 DVDD.n4936 DVDD.n4912 0.214786
R26388 DVDD.n4935 DVDD.n4934 0.214786
R26389 DVDD.n4933 DVDD.n4913 0.214786
R26390 DVDD.n4932 DVDD.n4931 0.214786
R26391 DVDD.n4930 DVDD.n4918 0.214786
R26392 DVDD.n4929 DVDD.n4928 0.214786
R26393 DVDD.n4927 DVDD.n4919 0.214786
R26394 DVDD.n4926 DVDD.n4925 0.214786
R26395 DVDD.n4924 DVDD.n480 0.214786
R26396 DVDD.n5249 DVDD.n451 0.214786
R26397 DVDD.n476 DVDD.n462 0.214786
R26398 DVDD.n5317 DVDD.n5316 0.214786
R26399 DVDD.n5315 DVDD.n475 0.214786
R26400 DVDD.n5314 DVDD.n5313 0.214786
R26401 DVDD.n5312 DVDD.n5256 0.214786
R26402 DVDD.n5311 DVDD.n5310 0.214786
R26403 DVDD.n5309 DVDD.n5257 0.214786
R26404 DVDD.n5308 DVDD.n5307 0.214786
R26405 DVDD.n5306 DVDD.n5262 0.214786
R26406 DVDD.n5305 DVDD.n5304 0.214786
R26407 DVDD.n5303 DVDD.n5263 0.214786
R26408 DVDD.n5302 DVDD.n5301 0.214786
R26409 DVDD.n5300 DVDD.n144 0.214786
R26410 DVDD.n5299 DVDD.n155 0.214786
R26411 DVDD.n5298 DVDD.n5297 0.214786
R26412 DVDD.n5296 DVDD.n5271 0.214786
R26413 DVDD.n5295 DVDD.n5294 0.214786
R26414 DVDD.n5293 DVDD.n5272 0.214786
R26415 DVDD.n5292 DVDD.n5291 0.214786
R26416 DVDD.n5290 DVDD.n5277 0.214786
R26417 DVDD.n5289 DVDD.n5288 0.214786
R26418 DVDD.n5287 DVDD.n5278 0.214786
R26419 DVDD.n5286 DVDD.n5285 0.214786
R26420 DVDD.n5284 DVDD.n42 0.214786
R26421 DVDD.n5938 DVDD.n5937 0.214786
R26422 DVDD.n5936 DVDD.n5935 0.214786
R26423 DVDD.n58 DVDD.n47 0.214786
R26424 DVDD.n5578 DVDD.n5566 0.214786
R26425 DVDD.n5603 DVDD.n5602 0.214786
R26426 DVDD.n5601 DVDD.n5577 0.214786
R26427 DVDD.n5600 DVDD.n5599 0.214786
R26428 DVDD.n5598 DVDD.n5584 0.214786
R26429 DVDD.n5597 DVDD.n5596 0.214786
R26430 DVDD.n5595 DVDD.n5585 0.214786
R26431 DVDD.n5594 DVDD.n5593 0.214786
R26432 DVDD.n4375 DVDD.n4374 0.214786
R26433 DVDD.n4373 DVDD.n1596 0.214786
R26434 DVDD.n4372 DVDD.n1607 0.214786
R26435 DVDD.n4371 DVDD.n4370 0.214786
R26436 DVDD.n4369 DVDD.n4351 0.214786
R26437 DVDD.n4368 DVDD.n4367 0.214786
R26438 DVDD.n4366 DVDD.n4352 0.214786
R26439 DVDD.n4365 DVDD.n4364 0.214786
R26440 DVDD.n4363 DVDD.n4357 0.214786
R26441 DVDD.n4362 DVDD.n4361 0.214786
R26442 DVDD.n985 DVDD.n975 0.214786
R26443 DVDD.n4645 DVDD.n4644 0.214786
R26444 DVDD.n4643 DVDD.n4642 0.214786
R26445 DVDD.n4641 DVDD.n4640 0.214786
R26446 DVDD.n4639 DVDD.n4638 0.214786
R26447 DVDD.n4636 DVDD.n4635 0.214786
R26448 DVDD.n4634 DVDD.n992 0.214786
R26449 DVDD.n4633 DVDD.n4632 0.214786
R26450 DVDD.n4631 DVDD.n993 0.214786
R26451 DVDD.n4630 DVDD.n4629 0.214786
R26452 DVDD.n4628 DVDD.n998 0.214786
R26453 DVDD.n4627 DVDD.n4626 0.214786
R26454 DVDD.n4625 DVDD.n999 0.214786
R26455 DVDD.n4624 DVDD.n4623 0.214786
R26456 DVDD.n4622 DVDD.n1004 0.214786
R26457 DVDD.n4621 DVDD.n4620 0.214786
R26458 DVDD.n4619 DVDD.n4618 0.214786
R26459 DVDD.n1046 DVDD.n1009 0.214786
R26460 DVDD.n1045 DVDD.n1044 0.214786
R26461 DVDD.n1043 DVDD.n1020 0.214786
R26462 DVDD.n1042 DVDD.n1041 0.214786
R26463 DVDD.n1040 DVDD.n1025 0.214786
R26464 DVDD.n1039 DVDD.n1038 0.214786
R26465 DVDD.n1037 DVDD.n1026 0.214786
R26466 DVDD.n1036 DVDD.n1035 0.214786
R26467 DVDD.n1034 DVDD.n1033 0.214786
R26468 DVDD.n729 DVDD.n728 0.214786
R26469 DVDD.n4876 DVDD.n4875 0.214786
R26470 DVDD.n4874 DVDD.n704 0.214786
R26471 DVDD.n4872 DVDD.n715 0.214786
R26472 DVDD.n4871 DVDD.n4870 0.214786
R26473 DVDD.n4869 DVDD.n4807 0.214786
R26474 DVDD.n4868 DVDD.n4867 0.214786
R26475 DVDD.n4866 DVDD.n4808 0.214786
R26476 DVDD.n4865 DVDD.n4864 0.214786
R26477 DVDD.n4863 DVDD.n4813 0.214786
R26478 DVDD.n4862 DVDD.n4861 0.214786
R26479 DVDD.n4860 DVDD.n4814 0.214786
R26480 DVDD.n4859 DVDD.n4858 0.214786
R26481 DVDD.n4857 DVDD.n4856 0.214786
R26482 DVDD.n4855 DVDD.n605 0.214786
R26483 DVDD.n4854 DVDD.n616 0.214786
R26484 DVDD.n4853 DVDD.n4852 0.214786
R26485 DVDD.n4851 DVDD.n4823 0.214786
R26486 DVDD.n4850 DVDD.n4849 0.214786
R26487 DVDD.n4848 DVDD.n4824 0.214786
R26488 DVDD.n4847 DVDD.n4846 0.214786
R26489 DVDD.n4845 DVDD.n4829 0.214786
R26490 DVDD.n4844 DVDD.n4843 0.214786
R26491 DVDD.n4842 DVDD.n4830 0.214786
R26492 DVDD.n4841 DVDD.n4840 0.214786
R26493 DVDD.n4839 DVDD.n4837 0.214786
R26494 DVDD.n4838 DVDD.n482 0.214786
R26495 DVDD.n5246 DVDD.n5245 0.214786
R26496 DVDD.n555 DVDD.n484 0.214786
R26497 DVDD.n554 DVDD.n553 0.214786
R26498 DVDD.n552 DVDD.n496 0.214786
R26499 DVDD.n551 DVDD.n550 0.214786
R26500 DVDD.n549 DVDD.n501 0.214786
R26501 DVDD.n548 DVDD.n547 0.214786
R26502 DVDD.n546 DVDD.n502 0.214786
R26503 DVDD.n545 DVDD.n544 0.214786
R26504 DVDD.n543 DVDD.n507 0.214786
R26505 DVDD.n542 DVDD.n541 0.214786
R26506 DVDD.n540 DVDD.n170 0.214786
R26507 DVDD.n539 DVDD.n180 0.214786
R26508 DVDD.n538 DVDD.n537 0.214786
R26509 DVDD.n536 DVDD.n513 0.214786
R26510 DVDD.n535 DVDD.n534 0.214786
R26511 DVDD.n533 DVDD.n514 0.214786
R26512 DVDD.n532 DVDD.n531 0.214786
R26513 DVDD.n530 DVDD.n519 0.214786
R26514 DVDD.n529 DVDD.n528 0.214786
R26515 DVDD.n527 DVDD.n520 0.214786
R26516 DVDD.n526 DVDD.n525 0.214786
R26517 DVDD.n39 DVDD.n37 0.214786
R26518 DVDD.n5942 DVDD.n5941 0.214786
R26519 DVDD.n33 DVDD.n32 0.214786
R26520 DVDD.n5953 DVDD.n5952 0.214786
R26521 DVDD.n5951 DVDD.n5950 0.214786
R26522 DVDD.n5949 DVDD.n7 0.214786
R26523 DVDD.n5957 DVDD.n6 0.214786
R26524 DVDD.n5959 DVDD.n5958 0.214786
R26525 DVDD.n4 DVDD.n3 0.214786
R26526 DVDD.n5965 DVDD.n5964 0.214786
R26527 DVDD.n5966 DVDD.n2 0.214786
R26528 DVDD.n5968 DVDD.n5967 0.214786
R26529 DVDD.n5969 DVDD.n0 0.214786
R26530 DVDD.n4332 DVDD.n4331 0.214786
R26531 DVDD.n4330 DVDD.n1628 0.214786
R26532 DVDD.n4329 DVDD.n1639 0.214786
R26533 DVDD.n4328 DVDD.n4327 0.214786
R26534 DVDD.n4326 DVDD.n4306 0.214786
R26535 DVDD.n4325 DVDD.n4324 0.214786
R26536 DVDD.n4323 DVDD.n4307 0.214786
R26537 DVDD.n4322 DVDD.n4321 0.214786
R26538 DVDD.n4320 DVDD.n4312 0.214786
R26539 DVDD.n4319 DVDD.n4318 0.214786
R26540 DVDD.n4317 DVDD.n4313 0.214786
R26541 DVDD.n4709 DVDD.n913 0.214786
R26542 DVDD.n4714 DVDD.n4713 0.214786
R26543 DVDD.n921 DVDD.n911 0.214786
R26544 DVDD.n4719 DVDD.n4718 0.214786
R26545 DVDD.n4722 DVDD.n4721 0.214786
R26546 DVDD.n906 DVDD.n905 0.214786
R26547 DVDD.n4727 DVDD.n4726 0.214786
R26548 DVDD.n4728 DVDD.n904 0.214786
R26549 DVDD.n4730 DVDD.n4729 0.214786
R26550 DVDD.n902 DVDD.n901 0.214786
R26551 DVDD.n4735 DVDD.n4734 0.214786
R26552 DVDD.n4736 DVDD.n900 0.214786
R26553 DVDD.n4738 DVDD.n4737 0.214786
R26554 DVDD.n898 DVDD.n897 0.214786
R26555 DVDD.n4743 DVDD.n4742 0.214786
R26556 DVDD.n891 DVDD.n890 0.214786
R26557 DVDD.n4748 DVDD.n4747 0.214786
R26558 DVDD.n888 DVDD.n887 0.214786
R26559 DVDD.n4753 DVDD.n4752 0.214786
R26560 DVDD.n4754 DVDD.n886 0.214786
R26561 DVDD.n4756 DVDD.n4755 0.214786
R26562 DVDD.n884 DVDD.n883 0.214786
R26563 DVDD.n4761 DVDD.n4760 0.214786
R26564 DVDD.n4762 DVDD.n882 0.214786
R26565 DVDD.n4764 DVDD.n4763 0.214786
R26566 DVDD.n880 DVDD.n879 0.214786
R26567 DVDD.n4771 DVDD.n4770 0.214786
R26568 DVDD.n4772 DVDD.n732 0.214786
R26569 DVDD.n4803 DVDD.n4802 0.214786
R26570 DVDD.n4801 DVDD.n734 0.214786
R26571 DVDD.n4800 DVDD.n4799 0.214786
R26572 DVDD.n4798 DVDD.n4776 0.214786
R26573 DVDD.n4797 DVDD.n4796 0.214786
R26574 DVDD.n4795 DVDD.n4781 0.214786
R26575 DVDD.n4794 DVDD.n4793 0.214786
R26576 DVDD.n4792 DVDD.n4782 0.214786
R26577 DVDD.n4791 DVDD.n4790 0.214786
R26578 DVDD.n4789 DVDD.n4788 0.214786
R26579 DVDD.n588 DVDD.n587 0.214786
R26580 DVDD.n5024 DVDD.n5023 0.214786
R26581 DVDD.n591 DVDD.n585 0.214786
R26582 DVDD.n5029 DVDD.n5028 0.214786
R26583 DVDD.n5030 DVDD.n583 0.214786
R26584 DVDD.n5032 DVDD.n5031 0.214786
R26585 DVDD.n581 DVDD.n580 0.214786
R26586 DVDD.n5037 DVDD.n5036 0.214786
R26587 DVDD.n5038 DVDD.n579 0.214786
R26588 DVDD.n5040 DVDD.n5039 0.214786
R26589 DVDD.n577 DVDD.n576 0.214786
R26590 DVDD.n5045 DVDD.n5044 0.214786
R26591 DVDD.n5046 DVDD.n575 0.214786
R26592 DVDD.n5048 DVDD.n5047 0.214786
R26593 DVDD.n5087 DVDD.n5086 0.214786
R26594 DVDD.n5085 DVDD.n5084 0.214786
R26595 DVDD.n5083 DVDD.n5053 0.214786
R26596 DVDD.n5082 DVDD.n5081 0.214786
R26597 DVDD.n5080 DVDD.n5054 0.214786
R26598 DVDD.n5079 DVDD.n5078 0.214786
R26599 DVDD.n5077 DVDD.n5059 0.214786
R26600 DVDD.n5076 DVDD.n5075 0.214786
R26601 DVDD.n5074 DVDD.n5060 0.214786
R26602 DVDD.n5073 DVDD.n5072 0.214786
R26603 DVDD.n5071 DVDD.n5065 0.214786
R26604 DVDD.n5070 DVDD.n5069 0.214786
R26605 DVDD.n200 DVDD.n197 0.214786
R26606 DVDD.n5729 DVDD.n5728 0.214786
R26607 DVDD.n5727 DVDD.n199 0.214786
R26608 DVDD.n5726 DVDD.n5725 0.214786
R26609 DVDD.n5724 DVDD.n204 0.214786
R26610 DVDD.n5723 DVDD.n5722 0.214786
R26611 DVDD.n5721 DVDD.n205 0.214786
R26612 DVDD.n5720 DVDD.n5719 0.214786
R26613 DVDD.n5718 DVDD.n210 0.214786
R26614 DVDD.n5717 DVDD.n5716 0.214786
R26615 DVDD.n5715 DVDD.n211 0.214786
R26616 DVDD.n5714 DVDD.n5713 0.214786
R26617 DVDD.n5711 DVDD.n5710 0.214786
R26618 DVDD.n220 DVDD.n217 0.214786
R26619 DVDD.n5703 DVDD.n5702 0.214786
R26620 DVDD.n5701 DVDD.n227 0.214786
R26621 DVDD.n5700 DVDD.n234 0.214786
R26622 DVDD.n5699 DVDD.n5698 0.214786
R26623 DVDD.n5697 DVDD.n5680 0.214786
R26624 DVDD.n5696 DVDD.n5695 0.214786
R26625 DVDD.n5694 DVDD.n5681 0.214786
R26626 DVDD.n5693 DVDD.n5692 0.214786
R26627 DVDD.n5691 DVDD.n5686 0.214786
R26628 DVDD.n2716 DVDD 0.209356
R26629 DVDD.n2720 DVDD.n2709 0.209134
R26630 DVDD.n961 DVDD.n960 0.208983
R26631 DVDD.n245 DVDD.n223 0.208899
R26632 DVDD.n2034 DVDD.n2033 0.208833
R26633 DVDD.n2030 DVDD.n2029 0.208833
R26634 DVDD.n2026 DVDD.n2025 0.208833
R26635 DVDD.n2022 DVDD.n2021 0.208833
R26636 DVDD.n2018 DVDD.n2017 0.208833
R26637 DVDD.n4205 DVDD.n4204 0.2085
R26638 DVDD.n4128 DVDD.n4127 0.2085
R26639 DVDD.n4123 DVDD.n4122 0.2085
R26640 DVDD.n4015 DVDD.n4014 0.2085
R26641 DVDD.n3996 DVDD.n3995 0.2085
R26642 DVDD.n3931 DVDD.n3930 0.2085
R26643 DVDD.n3934 DVDD.n3933 0.2085
R26644 DVDD.n1877 DVDD.n1876 0.2085
R26645 DVDD.n1868 DVDD.n1867 0.2085
R26646 DVDD.n1871 DVDD.n1870 0.2085
R26647 DVDD.n1716 DVDD.n1715 0.2085
R26648 DVDD.n4176 DVDD.n4175 0.2085
R26649 DVDD.n2720 DVDD.n2708 0.207634
R26650 DVDD.n3255 DVDD.n2734 0.2067
R26651 DVDD.n3255 DVDD.n2735 0.205865
R26652 DVDD.n5425 DVDD.n5424 0.204558
R26653 DVDD.n5920 DVDD.n5919 0.204245
R26654 DVDD DVDD.n2716 0.203019
R26655 DVDD.n2709 DVDD.n2701 0.201269
R26656 DVDD.n3389 DVDD.n2734 0.19985
R26657 DVDD.n3389 DVDD.n2735 0.199294
R26658 DVDD.n2708 DVDD.n2701 0.198908
R26659 DVDD.n3344 DVDD.n3343 0.198598
R26660 DVDD.n4203 DVDD 0.191088
R26661 DVDD.n3994 DVDD 0.191088
R26662 DVDD.n4013 DVDD 0.191088
R26663 DVDD.n1869 DVDD 0.191088
R26664 DVDD.n2607 DVDD.n2604 0.190625
R26665 DVDD.n4231 DVDD.n4230 0.1805
R26666 DVDD.n2517 DVDD.n2510 0.179316
R26667 DVDD.n1959 DVDD 0.176947
R26668 DVDD.n2013 DVDD 0.17636
R26669 DVDD.n3255 DVDD.n2742 0.174559
R26670 DVDD.n2720 DVDD.n2715 0.174401
R26671 DVDD.n3691 DVDD.n1898 0.174162
R26672 DVDD.n1743 DVDD.n1739 0.174048
R26673 DVDD DVDD.n1742 0.173778
R26674 DVDD.n1886 DVDD.n1885 0.173043
R26675 DVDD.n2602 DVDD.n2511 0.172185
R26676 DVDD DVDD.n2963 0.172062
R26677 DVDD DVDD.n1954 0.171551
R26678 DVDD.n2972 DVDD.n2966 0.168658
R26679 DVDD.n2982 DVDD.n2966 0.168658
R26680 DVDD.n2984 DVDD.n2731 0.168658
R26681 DVDD.n3396 DVDD.n2731 0.168658
R26682 DVDD.n3397 DVDD.n3396 0.168658
R26683 DVDD.n3408 DVDD.n3407 0.168658
R26684 DVDD.n3408 DVDD.n2705 0.168658
R26685 DVDD.n3419 DVDD.n2705 0.168658
R26686 DVDD.n3422 DVDD.n3421 0.168658
R26687 DVDD.n3422 DVDD.n2697 0.168658
R26688 DVDD.n3433 DVDD.n2697 0.168658
R26689 DVDD.n4266 DVDD.n1682 0.168658
R26690 DVDD.n4266 DVDD.n4265 0.168658
R26691 DVDD.n4265 DVDD.n1683 0.168658
R26692 DVDD.n3815 DVDD.n1842 0.168658
R26693 DVDD.n3816 DVDD.n3815 0.168658
R26694 DVDD.n3817 DVDD.n3816 0.168658
R26695 DVDD.n4067 DVDD.n4066 0.168658
R26696 DVDD.n4066 DVDD.n4056 0.168658
R26697 DVDD.n4056 DVDD.n1719 0.168658
R26698 DVDD.n4228 DVDD.n1720 0.168658
R26699 DVDD.n1762 DVDD.n1720 0.168658
R26700 DVDD.n1762 DVDD.n1761 0.168658
R26701 DVDD.n1740 DVDD.n1739 0.16842
R26702 DVDD.n2715 DVDD.n2701 0.168052
R26703 DVDD.n3707 DVDD.n1898 0.16771
R26704 DVDD.n1742 DVDD 0.167454
R26705 DVDD.n3389 DVDD.n2742 0.16731
R26706 DVDD.n1954 DVDD 0.166755
R26707 DVDD.n5488 DVDD.n263 0.165735
R26708 DVDD.n2963 DVDD 0.165645
R26709 DVDD.n5662 DVDD.n259 0.165589
R26710 DVDD.n1364 DVDD.n1363 0.164191
R26711 DVDD.n1576 DVDD.n1193 0.163126
R26712 DVDD.n2522 DVDD 0.160647
R26713 DVDD.n4204 DVDD.t126 0.152167
R26714 DVDD.n4204 DVDD.t116 0.152167
R26715 DVDD.n4127 DVDD.t138 0.152167
R26716 DVDD.n4127 DVDD.t122 0.152167
R26717 DVDD.n4122 DVDD.t128 0.152167
R26718 DVDD.n4122 DVDD.t155 0.152167
R26719 DVDD.n4014 DVDD.t203 0.152167
R26720 DVDD.n4014 DVDD.t99 0.152167
R26721 DVDD.n3995 DVDD.t46 0.152167
R26722 DVDD.n3995 DVDD.t44 0.152167
R26723 DVDD.n3930 DVDD.t157 0.152167
R26724 DVDD.n3930 DVDD.t120 0.152167
R26725 DVDD.n3933 DVDD.t36 0.152167
R26726 DVDD.n3933 DVDD.t42 0.152167
R26727 DVDD.n1876 DVDD.t34 0.152167
R26728 DVDD.n1876 DVDD.t28 0.152167
R26729 DVDD.n1867 DVDD.t97 0.152167
R26730 DVDD.n1867 DVDD.t143 0.152167
R26731 DVDD.n1870 DVDD.t190 0.152167
R26732 DVDD.n1870 DVDD.t151 0.152167
R26733 DVDD.n1715 DVDD.t72 0.152167
R26734 DVDD.n1715 DVDD.t74 0.152167
R26735 DVDD.n4175 DVDD.t153 0.152167
R26736 DVDD.n4175 DVDD.t145 0.152167
R26737 DVDD.n3447 DVDD.n2687 0.145128
R26738 DVDD.n1883 DVDD.n1882 0.144974
R26739 DVDD.n4190 DVDD.n1718 0.144974
R26740 DVDD.n2265 DVDD.n2125 0.140794
R26741 DVDD.n2150 DVDD.n2125 0.140794
R26742 DVDD.n2340 DVDD.n2061 0.140794
R26743 DVDD.n2084 DVDD.n2061 0.140794
R26744 DVDD.n5490 DVDD.n264 0.1405
R26745 DVDD.n5490 DVDD.n5489 0.1405
R26746 DVDD.n5665 DVDD.n5664 0.1405
R26747 DVDD.n5664 DVDD.n5663 0.1405
R26748 DVDD.n2150 DVDD 0.131529
R26749 DVDD DVDD.n2265 0.131529
R26750 DVDD.n2084 DVDD 0.131529
R26751 DVDD DVDD.n2340 0.131529
R26752 DVDD.n2198 DVDD 0.130161
R26753 DVDD.n3470 DVDD 0.130161
R26754 DVDD.n1363 DVDD 0.124869
R26755 DVDD.n3064 DVDD 0.123988
R26756 DVDD.n3043 DVDD 0.123988
R26757 DVDD.n2999 DVDD 0.123988
R26758 DVDD.n3018 DVDD 0.123988
R26759 DVDD.n1570 DVDD.n1193 0.122916
R26760 DVDD.n1966 DVDD.n1965 0.120105
R26761 DVDD.n1968 DVDD.n1967 0.115798
R26762 DVDD.n1945 DVDD.n1944 0.115798
R26763 DVDD.n3694 DVDD 0.115647
R26764 DVDD.n1948 DVDD.n1920 0.115053
R26765 DVDD.n3700 DVDD.n3699 0.115053
R26766 DVDD.n3222 DVDD.n3095 0.112392
R26767 DVDD.n3173 DVDD.n3172 0.112392
R26768 DVDD.n4124 DVDD.n1711 0.111676
R26769 DVDD.n3932 DVDD.n1709 0.111676
R26770 DVDD.n1151 DVDD.n1150 0.110634
R26771 DVDD.n4401 DVDD.n1106 0.110634
R26772 DVDD.n4348 DVDD.n4347 0.110634
R26773 DVDD.n4303 DVDD.n4302 0.110634
R26774 DVDD.n3162 DVDD.n3161 0.110634
R26775 DVDD.n3099 DVDD.n3097 0.110634
R26776 DVDD.n2977 DVDD.n2976 0.110634
R26777 DVDD.n3733 DVDD.n3723 0.110634
R26778 DVDD DVDD.n1964 0.109447
R26779 DVDD.n1932 DVDD 0.109447
R26780 DVDD DVDD.n1936 0.109447
R26781 DVDD.n3214 DVDD.n3117 0.1055
R26782 DVDD.n3214 DVDD.n3213 0.1055
R26783 DVDD.n3225 DVDD.n3108 0.1055
R26784 DVDD.n3226 DVDD.n3225 0.1055
R26785 DVDD DVDD.n2198 0.101206
R26786 DVDD.n3470 DVDD 0.101206
R26787 DVDD.n2598 DVDD.n2597 0.0931471
R26788 DVDD.n2597 DVDD.n2596 0.0931471
R26789 DVDD.n2983 DVDD.n2982 0.084579
R26790 DVDD.n2984 DVDD.n2983 0.084579
R26791 DVDD.n3420 DVDD.n3419 0.084579
R26792 DVDD.n3421 DVDD.n3420 0.084579
R26793 DVDD.n1880 DVDD.n1683 0.084579
R26794 DVDD.n1880 DVDD.n1842 0.084579
R26795 DVDD.n4229 DVDD.n1719 0.084579
R26796 DVDD.n4229 DVDD.n4228 0.084579
R26797 DVDD.n4387 DVDD.n4346 0.0815
R26798 DVDD.n4415 DVDD.n4389 0.0815
R26799 DVDD DVDD.n2521 0.0799118
R26800 DVDD.n1882 DVDD.n1881 0.0798421
R26801 DVDD.n1584 DVDD.n1583 0.079359
R26802 DVDD.n2599 DVDD.n2598 0.0786579
R26803 DVDD.n4200 DVDD.n4199 0.0780879
R26804 DVDD.n3776 DVDD.n3775 0.077225
R26805 DVDD.n3700 DVDD.n1912 0.0760366
R26806 DVDD.n1920 DVDD.n1919 0.0760366
R26807 DVDD.n1969 DVDD.n1968 0.0757132
R26808 DVDD.n1944 DVDD.n1939 0.0757132
R26809 DVDD.n3449 DVDD.n3448 0.0737558
R26810 DVDD.n3448 DVDD.n3447 0.0737558
R26811 DVDD.n3215 DVDD.n3214 0.066125
R26812 DVDD.n3225 DVDD.n3224 0.066125
R26813 DVDD.n5592 DVDD 0.0638222
R26814 DVDD.n5973 DVDD 0.0638222
R26815 DVDD.n5690 DVDD 0.0638222
R26816 DVDD.n5898 DVDD 0.0638222
R26817 DVDD.n3168 DVDD.n3107 0.0624947
R26818 DVDD.n3228 DVDD.n3107 0.0624947
R26819 DVDD.n4199 DVDD 0.0592637
R26820 DVDD.n3698 DVDD.n3697 0.0574118
R26821 DVDD.n5633 DVDD.n5632 0.0560556
R26822 DVDD.n5539 DVDD.n13 0.0560556
R26823 DVDD.n4678 DVDD.n980 0.0560556
R26824 DVDD.n5458 DVDD.n5457 0.0560556
R26825 DVDD.n1902 DVDD.n1896 0.0527336
R26826 DVDD.n1906 DVDD.n1896 0.0527336
R26827 DVDD.n5502 DVDD.n260 0.0523993
R26828 DVDD.n3255 DVDD.n2736 0.0518309
R26829 DVDD.n2714 DVDD.n2702 0.0515891
R26830 DVDD.n2712 DVDD.n2702 0.0515891
R26831 DVDD.n2710 DVDD.n2702 0.0515891
R26832 DVDD.n4082 DVDD.n4046 0.0515891
R26833 DVDD.n3903 DVDD.n3902 0.0515891
R26834 DVDD.n2750 DVDD.n2741 0.0515881
R26835 DVDD.n1897 DVDD.n1896 0.0515834
R26836 DVDD.n2750 DVDD.n2746 0.0515834
R26837 DVDD.n3834 DVDD.n1830 0.0515834
R26838 DVDD.n4046 DVDD.n4045 0.0509336
R26839 DVDD.n3389 DVDD.n2736 0.0505959
R26840 DVDD.n2711 DVDD.n2702 0.0503876
R26841 DVDD.n2713 DVDD.n2702 0.0503876
R26842 DVDD.n2707 DVDD.n2702 0.0503876
R26843 DVDD.n3902 DVDD.n3870 0.0503876
R26844 DVDD.n1905 DVDD.n1896 0.0497891
R26845 DVDD.n1909 DVDD.n1896 0.0497891
R26846 DVDD.n1831 DVDD.n1830 0.0497834
R26847 DVDD.n2750 DVDD.n2740 0.0497834
R26848 DVDD.n2750 DVDD.n2747 0.0497834
R26849 DVDD DVDD.n5898 0.0487259
R26850 DVDD DVDD.n5592 0.0487259
R26851 DVDD DVDD.n5973 0.0487259
R26852 DVDD DVDD.n5690 0.0487259
R26853 DVDD.n2821 DVDD.n2820 0.0467228
R26854 DVDD.n3337 DVDD.n3336 0.0467228
R26855 DVDD.n5732 DVDD.n194 0.0462377
R26856 DVDD.n5738 DVDD.n194 0.0462377
R26857 DVDD.n5739 DVDD.n5738 0.0462377
R26858 DVDD.n5739 DVDD.n192 0.0462377
R26859 DVDD.n5743 DVDD.n192 0.0462377
R26860 DVDD.n5744 DVDD.n5743 0.0462377
R26861 DVDD.n5747 DVDD.n5744 0.0462377
R26862 DVDD.n5749 DVDD.n5747 0.0462377
R26863 DVDD.n5751 DVDD.n5749 0.0462377
R26864 DVDD.n5753 DVDD.n5751 0.0462377
R26865 DVDD.n5755 DVDD.n5753 0.0462377
R26866 DVDD.n5757 DVDD.n5755 0.0462377
R26867 DVDD.n5759 DVDD.n5757 0.0462377
R26868 DVDD.n5760 DVDD.n5759 0.0462377
R26869 DVDD.n5763 DVDD.n5760 0.0462377
R26870 DVDD.n5765 DVDD.n5763 0.0462377
R26871 DVDD.n5767 DVDD.n5765 0.0462377
R26872 DVDD.n5769 DVDD.n5767 0.0462377
R26873 DVDD.n5771 DVDD.n5769 0.0462377
R26874 DVDD.n5773 DVDD.n5771 0.0462377
R26875 DVDD.n5774 DVDD.n5773 0.0462377
R26876 DVDD.n5782 DVDD.n5774 0.0462377
R26877 DVDD.n5782 DVDD.n5781 0.0462377
R26878 DVDD.n5781 DVDD.n5780 0.0462377
R26879 DVDD.n5780 DVDD.n5778 0.0462377
R26880 DVDD.n5778 DVDD.n5776 0.0462377
R26881 DVDD.n5776 DVDD.n167 0.0462377
R26882 DVDD.n5788 DVDD.n167 0.0462377
R26883 DVDD.n5789 DVDD.n5788 0.0462377
R26884 DVDD.n5793 DVDD.n165 0.0462377
R26885 DVDD.n5794 DVDD.n5793 0.0462377
R26886 DVDD.n5833 DVDD.n5794 0.0462377
R26887 DVDD.n5833 DVDD.n5832 0.0462377
R26888 DVDD.n5832 DVDD.n5829 0.0462377
R26889 DVDD.n5829 DVDD.n5828 0.0462377
R26890 DVDD.n5828 DVDD.n5826 0.0462377
R26891 DVDD.n5826 DVDD.n5824 0.0462377
R26892 DVDD.n5824 DVDD.n5822 0.0462377
R26893 DVDD.n5822 DVDD.n5820 0.0462377
R26894 DVDD.n5820 DVDD.n5818 0.0462377
R26895 DVDD.n5818 DVDD.n5816 0.0462377
R26896 DVDD.n5816 DVDD.n5813 0.0462377
R26897 DVDD.n5813 DVDD.n5812 0.0462377
R26898 DVDD.n5812 DVDD.n5810 0.0462377
R26899 DVDD.n5810 DVDD.n5808 0.0462377
R26900 DVDD.n5808 DVDD.n5806 0.0462377
R26901 DVDD.n5806 DVDD.n5804 0.0462377
R26902 DVDD.n5804 DVDD.n5802 0.0462377
R26903 DVDD.n5802 DVDD.n5800 0.0462377
R26904 DVDD.n5800 DVDD.n5797 0.0462377
R26905 DVDD.n5797 DVDD.n5796 0.0462377
R26906 DVDD.n5796 DVDD.n141 0.0462377
R26907 DVDD.n5839 DVDD.n141 0.0462377
R26908 DVDD.n5840 DVDD.n5839 0.0462377
R26909 DVDD.n5840 DVDD.n139 0.0462377
R26910 DVDD.n5844 DVDD.n139 0.0462377
R26911 DVDD.n5846 DVDD.n5844 0.0462377
R26912 DVDD.n5848 DVDD.n5846 0.0462377
R26913 DVDD.n5741 DVDD.n5740 0.0462377
R26914 DVDD.n5742 DVDD.n5741 0.0462377
R26915 DVDD.n5746 DVDD.n5745 0.0462377
R26916 DVDD.n5762 DVDD.n5761 0.0462377
R26917 DVDD.n5783 DVDD.n191 0.0462377
R26918 DVDD.n5791 DVDD.n5790 0.0462377
R26919 DVDD.n5792 DVDD.n5791 0.0462377
R26920 DVDD.n5831 DVDD.n5830 0.0462377
R26921 DVDD.n5815 DVDD.n5814 0.0462377
R26922 DVDD.n5799 DVDD.n5798 0.0462377
R26923 DVDD.n5842 DVDD.n5841 0.0462377
R26924 DVDD.n5843 DVDD.n5842 0.0462377
R26925 DVDD.n5093 DVDD.n5092 0.0462377
R26926 DVDD.n5092 DVDD.n5090 0.0462377
R26927 DVDD.n5090 DVDD.n568 0.0462377
R26928 DVDD.n5100 DVDD.n568 0.0462377
R26929 DVDD.n5101 DVDD.n5100 0.0462377
R26930 DVDD.n5241 DVDD.n5101 0.0462377
R26931 DVDD.n5241 DVDD.n5240 0.0462377
R26932 DVDD.n5240 DVDD.n5239 0.0462377
R26933 DVDD.n5239 DVDD.n5237 0.0462377
R26934 DVDD.n5237 DVDD.n5235 0.0462377
R26935 DVDD.n5235 DVDD.n5233 0.0462377
R26936 DVDD.n5233 DVDD.n5231 0.0462377
R26937 DVDD.n5231 DVDD.n5229 0.0462377
R26938 DVDD.n5229 DVDD.n5227 0.0462377
R26939 DVDD.n5227 DVDD.n5224 0.0462377
R26940 DVDD.n5224 DVDD.n5223 0.0462377
R26941 DVDD.n5223 DVDD.n5221 0.0462377
R26942 DVDD.n5221 DVDD.n5219 0.0462377
R26943 DVDD.n5219 DVDD.n5217 0.0462377
R26944 DVDD.n5217 DVDD.n5215 0.0462377
R26945 DVDD.n5215 DVDD.n5213 0.0462377
R26946 DVDD.n5213 DVDD.n5211 0.0462377
R26947 DVDD.n5211 DVDD.n5208 0.0462377
R26948 DVDD.n5208 DVDD.n5207 0.0462377
R26949 DVDD.n5207 DVDD.n5205 0.0462377
R26950 DVDD.n5205 DVDD.n5203 0.0462377
R26951 DVDD.n5203 DVDD.n5201 0.0462377
R26952 DVDD.n5201 DVDD.n5199 0.0462377
R26953 DVDD.n5199 DVDD.n5197 0.0462377
R26954 DVDD.n5193 DVDD.n5102 0.0462377
R26955 DVDD.n5193 DVDD.n5192 0.0462377
R26956 DVDD.n5192 DVDD.n5190 0.0462377
R26957 DVDD.n5190 DVDD.n5188 0.0462377
R26958 DVDD.n5188 DVDD.n5185 0.0462377
R26959 DVDD.n5185 DVDD.n5184 0.0462377
R26960 DVDD.n5184 DVDD.n5182 0.0462377
R26961 DVDD.n5182 DVDD.n5180 0.0462377
R26962 DVDD.n5180 DVDD.n5178 0.0462377
R26963 DVDD.n5178 DVDD.n5176 0.0462377
R26964 DVDD.n5176 DVDD.n5174 0.0462377
R26965 DVDD.n5174 DVDD.n5172 0.0462377
R26966 DVDD.n5172 DVDD.n5169 0.0462377
R26967 DVDD.n5169 DVDD.n5168 0.0462377
R26968 DVDD.n5168 DVDD.n5166 0.0462377
R26969 DVDD.n5166 DVDD.n5164 0.0462377
R26970 DVDD.n5164 DVDD.n5162 0.0462377
R26971 DVDD.n5162 DVDD.n5160 0.0462377
R26972 DVDD.n5160 DVDD.n5158 0.0462377
R26973 DVDD.n5158 DVDD.n5156 0.0462377
R26974 DVDD.n5156 DVDD.n5153 0.0462377
R26975 DVDD.n5153 DVDD.n5152 0.0462377
R26976 DVDD.n5152 DVDD.n5150 0.0462377
R26977 DVDD.n5150 DVDD.n5149 0.0462377
R26978 DVDD.n5149 DVDD.n5148 0.0462377
R26979 DVDD.n5148 DVDD.n5103 0.0462377
R26980 DVDD.n5144 DVDD.n5103 0.0462377
R26981 DVDD.n5144 DVDD.n5143 0.0462377
R26982 DVDD.n5143 DVDD.n5105 0.0462377
R26983 DVDD.n5099 DVDD.n5098 0.0462377
R26984 DVDD.n5099 DVDD.n566 0.0462377
R26985 DVDD.n5242 DVDD.n567 0.0462377
R26986 DVDD.n5226 DVDD.n5225 0.0462377
R26987 DVDD.n5210 DVDD.n5209 0.0462377
R26988 DVDD.n5196 DVDD.n5195 0.0462377
R26989 DVDD.n5195 DVDD.n5194 0.0462377
R26990 DVDD.n5187 DVDD.n5186 0.0462377
R26991 DVDD.n5171 DVDD.n5170 0.0462377
R26992 DVDD.n5155 DVDD.n5154 0.0462377
R26993 DVDD.n5147 DVDD.n5146 0.0462377
R26994 DVDD.n5146 DVDD.n5145 0.0462377
R26995 DVDD.n600 DVDD.n598 0.0462377
R26996 DVDD.n601 DVDD.n600 0.0462377
R26997 DVDD.n5019 DVDD.n601 0.0462377
R26998 DVDD.n5019 DVDD.n5018 0.0462377
R26999 DVDD.n5018 DVDD.n5017 0.0462377
R27000 DVDD.n5017 DVDD.n602 0.0462377
R27001 DVDD.n629 DVDD.n602 0.0462377
R27002 DVDD.n631 DVDD.n629 0.0462377
R27003 DVDD.n633 DVDD.n631 0.0462377
R27004 DVDD.n635 DVDD.n633 0.0462377
R27005 DVDD.n637 DVDD.n635 0.0462377
R27006 DVDD.n639 DVDD.n637 0.0462377
R27007 DVDD.n641 DVDD.n639 0.0462377
R27008 DVDD.n642 DVDD.n641 0.0462377
R27009 DVDD.n645 DVDD.n642 0.0462377
R27010 DVDD.n647 DVDD.n645 0.0462377
R27011 DVDD.n649 DVDD.n647 0.0462377
R27012 DVDD.n651 DVDD.n649 0.0462377
R27013 DVDD.n653 DVDD.n651 0.0462377
R27014 DVDD.n655 DVDD.n653 0.0462377
R27015 DVDD.n657 DVDD.n655 0.0462377
R27016 DVDD.n658 DVDD.n657 0.0462377
R27017 DVDD.n661 DVDD.n658 0.0462377
R27018 DVDD.n663 DVDD.n661 0.0462377
R27019 DVDD.n665 DVDD.n663 0.0462377
R27020 DVDD.n667 DVDD.n665 0.0462377
R27021 DVDD.n669 DVDD.n667 0.0462377
R27022 DVDD.n670 DVDD.n669 0.0462377
R27023 DVDD.n5011 DVDD.n670 0.0462377
R27024 DVDD.n5010 DVDD.n5009 0.0462377
R27025 DVDD.n5009 DVDD.n671 0.0462377
R27026 DVDD.n4953 DVDD.n671 0.0462377
R27027 DVDD.n4954 DVDD.n4953 0.0462377
R27028 DVDD.n4957 DVDD.n4954 0.0462377
R27029 DVDD.n4959 DVDD.n4957 0.0462377
R27030 DVDD.n4961 DVDD.n4959 0.0462377
R27031 DVDD.n4963 DVDD.n4961 0.0462377
R27032 DVDD.n4965 DVDD.n4963 0.0462377
R27033 DVDD.n4967 DVDD.n4965 0.0462377
R27034 DVDD.n4969 DVDD.n4967 0.0462377
R27035 DVDD.n4970 DVDD.n4969 0.0462377
R27036 DVDD.n4973 DVDD.n4970 0.0462377
R27037 DVDD.n4975 DVDD.n4973 0.0462377
R27038 DVDD.n4977 DVDD.n4975 0.0462377
R27039 DVDD.n4979 DVDD.n4977 0.0462377
R27040 DVDD.n4981 DVDD.n4979 0.0462377
R27041 DVDD.n4983 DVDD.n4981 0.0462377
R27042 DVDD.n4985 DVDD.n4983 0.0462377
R27043 DVDD.n4986 DVDD.n4985 0.0462377
R27044 DVDD.n4989 DVDD.n4986 0.0462377
R27045 DVDD.n4991 DVDD.n4989 0.0462377
R27046 DVDD.n4992 DVDD.n4991 0.0462377
R27047 DVDD.n5003 DVDD.n4992 0.0462377
R27048 DVDD.n5003 DVDD.n5002 0.0462377
R27049 DVDD.n5002 DVDD.n4993 0.0462377
R27050 DVDD.n4998 DVDD.n4993 0.0462377
R27051 DVDD.n4998 DVDD.n4997 0.0462377
R27052 DVDD.n4997 DVDD.n4995 0.0462377
R27053 DVDD.n5020 DVDD.n595 0.0462377
R27054 DVDD.n5016 DVDD.n595 0.0462377
R27055 DVDD.n628 DVDD.n604 0.0462377
R27056 DVDD.n644 DVDD.n643 0.0462377
R27057 DVDD.n660 DVDD.n659 0.0462377
R27058 DVDD.n5012 DVDD.n627 0.0462377
R27059 DVDD.n5008 DVDD.n627 0.0462377
R27060 DVDD.n4956 DVDD.n4955 0.0462377
R27061 DVDD.n4972 DVDD.n4971 0.0462377
R27062 DVDD.n4988 DVDD.n4987 0.0462377
R27063 DVDD.n5001 DVDD.n5000 0.0462377
R27064 DVDD.n5000 DVDD.n4999 0.0462377
R27065 DVDD.n877 DVDD.n875 0.0462377
R27066 DVDD.n875 DVDD.n873 0.0462377
R27067 DVDD.n873 DVDD.n871 0.0462377
R27068 DVDD.n871 DVDD.n868 0.0462377
R27069 DVDD.n868 DVDD.n867 0.0462377
R27070 DVDD.n867 DVDD.n866 0.0462377
R27071 DVDD.n866 DVDD.n865 0.0462377
R27072 DVDD.n865 DVDD.n863 0.0462377
R27073 DVDD.n863 DVDD.n861 0.0462377
R27074 DVDD.n861 DVDD.n859 0.0462377
R27075 DVDD.n859 DVDD.n857 0.0462377
R27076 DVDD.n857 DVDD.n855 0.0462377
R27077 DVDD.n855 DVDD.n853 0.0462377
R27078 DVDD.n853 DVDD.n851 0.0462377
R27079 DVDD.n851 DVDD.n848 0.0462377
R27080 DVDD.n848 DVDD.n847 0.0462377
R27081 DVDD.n847 DVDD.n845 0.0462377
R27082 DVDD.n845 DVDD.n843 0.0462377
R27083 DVDD.n843 DVDD.n841 0.0462377
R27084 DVDD.n841 DVDD.n839 0.0462377
R27085 DVDD.n839 DVDD.n837 0.0462377
R27086 DVDD.n837 DVDD.n835 0.0462377
R27087 DVDD.n835 DVDD.n832 0.0462377
R27088 DVDD.n832 DVDD.n831 0.0462377
R27089 DVDD.n831 DVDD.n829 0.0462377
R27090 DVDD.n829 DVDD.n827 0.0462377
R27091 DVDD.n827 DVDD.n825 0.0462377
R27092 DVDD.n825 DVDD.n823 0.0462377
R27093 DVDD.n823 DVDD.n821 0.0462377
R27094 DVDD.n817 DVDD.n739 0.0462377
R27095 DVDD.n817 DVDD.n816 0.0462377
R27096 DVDD.n816 DVDD.n741 0.0462377
R27097 DVDD.n810 DVDD.n741 0.0462377
R27098 DVDD.n810 DVDD.n809 0.0462377
R27099 DVDD.n809 DVDD.n808 0.0462377
R27100 DVDD.n808 DVDD.n743 0.0462377
R27101 DVDD.n802 DVDD.n743 0.0462377
R27102 DVDD.n802 DVDD.n801 0.0462377
R27103 DVDD.n801 DVDD.n746 0.0462377
R27104 DVDD.n795 DVDD.n746 0.0462377
R27105 DVDD.n795 DVDD.n794 0.0462377
R27106 DVDD.n794 DVDD.n748 0.0462377
R27107 DVDD.n789 DVDD.n748 0.0462377
R27108 DVDD.n789 DVDD.n788 0.0462377
R27109 DVDD.n788 DVDD.n750 0.0462377
R27110 DVDD.n782 DVDD.n750 0.0462377
R27111 DVDD.n782 DVDD.n781 0.0462377
R27112 DVDD.n781 DVDD.n752 0.0462377
R27113 DVDD.n775 DVDD.n752 0.0462377
R27114 DVDD.n775 DVDD.n774 0.0462377
R27115 DVDD.n774 DVDD.n773 0.0462377
R27116 DVDD.n773 DVDD.n754 0.0462377
R27117 DVDD.n767 DVDD.n754 0.0462377
R27118 DVDD.n767 DVDD.n766 0.0462377
R27119 DVDD.n766 DVDD.n757 0.0462377
R27120 DVDD.n762 DVDD.n757 0.0462377
R27121 DVDD.n762 DVDD.n761 0.0462377
R27122 DVDD.n761 DVDD.n759 0.0462377
R27123 DVDD.n870 DVDD.n869 0.0462377
R27124 DVDD.n869 DVDD.n726 0.0462377
R27125 DVDD.n864 DVDD.n727 0.0462377
R27126 DVDD.n850 DVDD.n849 0.0462377
R27127 DVDD.n834 DVDD.n833 0.0462377
R27128 DVDD.n820 DVDD.n819 0.0462377
R27129 DVDD.n819 DVDD.n818 0.0462377
R27130 DVDD.n811 DVDD.n742 0.0462377
R27131 DVDD.n793 DVDD.n792 0.0462377
R27132 DVDD.n776 DVDD.n753 0.0462377
R27133 DVDD.n765 DVDD.n764 0.0462377
R27134 DVDD.n764 DVDD.n763 0.0462377
R27135 DVDD.n1062 DVDD.n1060 0.0462377
R27136 DVDD.n1064 DVDD.n1062 0.0462377
R27137 DVDD.n1065 DVDD.n1064 0.0462377
R27138 DVDD.n1068 DVDD.n1065 0.0462377
R27139 DVDD.n1069 DVDD.n1068 0.0462377
R27140 DVDD.n4614 DVDD.n1069 0.0462377
R27141 DVDD.n4614 DVDD.n4613 0.0462377
R27142 DVDD.n4613 DVDD.n4612 0.0462377
R27143 DVDD.n4612 DVDD.n4610 0.0462377
R27144 DVDD.n4610 DVDD.n4608 0.0462377
R27145 DVDD.n4608 DVDD.n4606 0.0462377
R27146 DVDD.n4606 DVDD.n4604 0.0462377
R27147 DVDD.n4604 DVDD.n4602 0.0462377
R27148 DVDD.n4602 DVDD.n4600 0.0462377
R27149 DVDD.n4600 DVDD.n4597 0.0462377
R27150 DVDD.n4597 DVDD.n4596 0.0462377
R27151 DVDD.n4596 DVDD.n4594 0.0462377
R27152 DVDD.n4594 DVDD.n4592 0.0462377
R27153 DVDD.n4592 DVDD.n4590 0.0462377
R27154 DVDD.n4590 DVDD.n4588 0.0462377
R27155 DVDD.n4588 DVDD.n4586 0.0462377
R27156 DVDD.n4586 DVDD.n4584 0.0462377
R27157 DVDD.n4584 DVDD.n4581 0.0462377
R27158 DVDD.n4581 DVDD.n4580 0.0462377
R27159 DVDD.n4580 DVDD.n4578 0.0462377
R27160 DVDD.n4578 DVDD.n4576 0.0462377
R27161 DVDD.n4576 DVDD.n4574 0.0462377
R27162 DVDD.n4574 DVDD.n4572 0.0462377
R27163 DVDD.n4572 DVDD.n4570 0.0462377
R27164 DVDD.n4566 DVDD.n1070 0.0462377
R27165 DVDD.n4566 DVDD.n4565 0.0462377
R27166 DVDD.n4565 DVDD.n1072 0.0462377
R27167 DVDD.n4510 DVDD.n1072 0.0462377
R27168 DVDD.n4513 DVDD.n4510 0.0462377
R27169 DVDD.n4515 DVDD.n4513 0.0462377
R27170 DVDD.n4517 DVDD.n4515 0.0462377
R27171 DVDD.n4519 DVDD.n4517 0.0462377
R27172 DVDD.n4521 DVDD.n4519 0.0462377
R27173 DVDD.n4523 DVDD.n4521 0.0462377
R27174 DVDD.n4525 DVDD.n4523 0.0462377
R27175 DVDD.n4526 DVDD.n4525 0.0462377
R27176 DVDD.n4529 DVDD.n4526 0.0462377
R27177 DVDD.n4531 DVDD.n4529 0.0462377
R27178 DVDD.n4533 DVDD.n4531 0.0462377
R27179 DVDD.n4535 DVDD.n4533 0.0462377
R27180 DVDD.n4537 DVDD.n4535 0.0462377
R27181 DVDD.n4539 DVDD.n4537 0.0462377
R27182 DVDD.n4541 DVDD.n4539 0.0462377
R27183 DVDD.n4542 DVDD.n4541 0.0462377
R27184 DVDD.n4545 DVDD.n4542 0.0462377
R27185 DVDD.n4547 DVDD.n4545 0.0462377
R27186 DVDD.n4548 DVDD.n4547 0.0462377
R27187 DVDD.n4559 DVDD.n4548 0.0462377
R27188 DVDD.n4559 DVDD.n4558 0.0462377
R27189 DVDD.n4558 DVDD.n4549 0.0462377
R27190 DVDD.n4554 DVDD.n4549 0.0462377
R27191 DVDD.n4554 DVDD.n4553 0.0462377
R27192 DVDD.n4553 DVDD.n4551 0.0462377
R27193 DVDD.n1067 DVDD.n1066 0.0462377
R27194 DVDD.n1067 DVDD.n1057 0.0462377
R27195 DVDD.n4615 DVDD.n1058 0.0462377
R27196 DVDD.n4599 DVDD.n4598 0.0462377
R27197 DVDD.n4583 DVDD.n4582 0.0462377
R27198 DVDD.n4569 DVDD.n4568 0.0462377
R27199 DVDD.n4568 DVDD.n4567 0.0462377
R27200 DVDD.n4512 DVDD.n4511 0.0462377
R27201 DVDD.n4528 DVDD.n4527 0.0462377
R27202 DVDD.n4544 DVDD.n4543 0.0462377
R27203 DVDD.n4557 DVDD.n4556 0.0462377
R27204 DVDD.n4556 DVDD.n4555 0.0462377
R27205 DVDD.n5513 DVDD.n28 0.0462377
R27206 DVDD.n4702 DVDD.n949 0.0462377
R27207 DVDD.n5789 DVDD.n165 0.0462377
R27208 DVDD.n5197 DVDD.n5102 0.0462377
R27209 DVDD.n5011 DVDD.n5010 0.0462377
R27210 DVDD.n821 DVDD.n739 0.0462377
R27211 DVDD.n4570 DVDD.n1070 0.0462377
R27212 DVDD.n3148 DVDD.n3107 0.0461522
R27213 DVDD.n2200 DVDD 0.0459167
R27214 DVDD.n2201 DVDD 0.0459167
R27215 DVDD.n3079 DVDD.n2745 0.0452755
R27216 DVDD.n5827 DVDD.n163 0.0451311
R27217 DVDD.n5183 DVDD.n468 0.0451311
R27218 DVDD.n4958 DVDD.n4946 0.0451311
R27219 DVDD.n807 DVDD.n744 0.0451311
R27220 DVDD.n4514 DVDD.n4505 0.0451311
R27221 DVDD.n5748 DVDD.n174 0.0447623
R27222 DVDD.n5238 DVDD.n486 0.0447623
R27223 DVDD.n630 DVDD.n610 0.0447623
R27224 DVDD.n862 DVDD.n705 0.0447623
R27225 DVDD.n4611 DVDD.n1010 0.0447623
R27226 DVDD.n1382 DVDD.n1313 0.0446743
R27227 DVDD.n1390 DVDD.n1309 0.0446743
R27228 DVDD.n1318 DVDD.n1216 0.0446743
R27229 DVDD.n1314 DVDD.n1214 0.0446743
R27230 DVDD.n5657 DVDD.n5656 0.0445261
R27231 DVDD.n5483 DVDD.n5482 0.0445261
R27232 DVDD.n5811 DVDD.n150 0.0443934
R27233 DVDD.n5167 DVDD.n466 0.0443934
R27234 DVDD.n4974 DVDD.n4944 0.0443934
R27235 DVDD.n791 DVDD.n790 0.0443934
R27236 DVDD.n4530 DVDD.n4503 0.0443934
R27237 DVDD.n3246 DVDD.n3088 0.0442838
R27238 DVDD.n3176 DVDD.n3125 0.0442838
R27239 DVDD.n3178 DVDD.n3174 0.0442838
R27240 DVDD.n3178 DVDD.n3177 0.0442838
R27241 DVDD.n3202 DVDD.n3124 0.0442838
R27242 DVDD.n3238 DVDD.n3236 0.0442838
R27243 DVDD.n3238 DVDD.n3237 0.0442838
R27244 DVDD.n3248 DVDD.n3247 0.0442838
R27245 DVDD.n5764 DVDD.n176 0.0440246
R27246 DVDD.n5222 DVDD.n562 0.0440246
R27247 DVDD.n646 DVDD.n612 0.0440246
R27248 DVDD.n846 DVDD.n722 0.0440246
R27249 DVDD.n4595 DVDD.n1053 0.0440246
R27250 DVDD.n5795 DVDD.n156 0.0436557
R27251 DVDD.n5151 DVDD.n464 0.0436557
R27252 DVDD.n4990 DVDD.n4942 0.0436557
R27253 DVDD.n772 DVDD.n755 0.0436557
R27254 DVDD.n4546 DVDD.n4501 0.0436557
R27255 DVDD.n3175 DVDD.n3124 0.043473
R27256 DVDD.n3247 DVDD.n3087 0.043473
R27257 DVDD.n5779 DVDD.n178 0.0432869
R27258 DVDD.n5206 DVDD.n493 0.0432869
R27259 DVDD.n662 DVDD.n614 0.0432869
R27260 DVDD.n830 DVDD.n712 0.0432869
R27261 DVDD.n4579 DVDD.n1017 0.0432869
R27262 DVDD.n5929 DVDD.n5928 0.0428146
R27263 DVDD.n5432 DVDD.n296 0.0428146
R27264 DVDD.n5784 DVDD.n190 0.0425492
R27265 DVDD.n5212 DVDD.n559 0.0425492
R27266 DVDD.n656 DVDD.n625 0.0425492
R27267 DVDD.n836 DVDD.n719 0.0425492
R27268 DVDD.n4585 DVDD.n1050 0.0425492
R27269 DVDD.n5801 DVDD.n153 0.0421803
R27270 DVDD.n5157 DVDD.n452 0.0421803
R27271 DVDD.n4984 DVDD.n675 0.0421803
R27272 DVDD.n778 DVDD.n777 0.0421803
R27273 DVDD.n4540 DVDD.n1076 0.0421803
R27274 DVDD.n5758 DVDD.n172 0.0418115
R27275 DVDD.n5228 DVDD.n489 0.0418115
R27276 DVDD.n640 DVDD.n608 0.0418115
R27277 DVDD.n852 DVDD.n708 0.0418115
R27278 DVDD.n4601 DVDD.n1013 0.0418115
R27279 DVDD.n5817 DVDD.n160 0.0414426
R27280 DVDD.n5173 DVDD.n471 0.0414426
R27281 DVDD.n4968 DVDD.n4949 0.0414426
R27282 DVDD.n796 DVDD.n747 0.0414426
R27283 DVDD.n4524 DVDD.n4507 0.0414426
R27284 DVDD.n2625 DVDD.n2624 0.0410978
R27285 DVDD.n5742 DVDD.n187 0.0410738
R27286 DVDD.n5243 DVDD.n566 0.0410738
R27287 DVDD.n5016 DVDD.n5015 0.0410738
R27288 DVDD.n4878 DVDD.n726 0.0410738
R27289 DVDD.n4616 DVDD.n1057 0.0410738
R27290 DVDD.n5834 DVDD.n146 0.0407049
R27291 DVDD.n5189 DVDD.n455 0.0407049
R27292 DVDD.n4952 DVDD.n678 0.0407049
R27293 DVDD.n813 DVDD.n812 0.0407049
R27294 DVDD.n1079 DVDD.n1074 0.0407049
R27295 DVDD.n5928 DVDD.n5927 0.0393914
R27296 DVDD.n5432 DVDD.n5431 0.0393914
R27297 DVDD.n5825 DVDD.n147 0.0384918
R27298 DVDD.n5181 DVDD.n457 0.0384918
R27299 DVDD.n4960 DVDD.n679 0.0384918
R27300 DVDD.n806 DVDD.n805 0.0384918
R27301 DVDD.n4516 DVDD.n1080 0.0384918
R27302 DVDD.n5750 DVDD.n186 0.038123
R27303 DVDD.n5236 DVDD.n565 0.038123
R27304 DVDD.n632 DVDD.n622 0.038123
R27305 DVDD.n860 DVDD.n725 0.038123
R27306 DVDD.n4609 DVDD.n1056 0.038123
R27307 DVDD.n2623 DVDD.n2499 0.03785
R27308 DVDD.n3240 DVDD.n3239 0.0377973
R27309 DVDD.n3179 DVDD.n3142 0.0377973
R27310 DVDD.n5809 DVDD.n159 0.0377541
R27311 DVDD.n5165 DVDD.n459 0.0377541
R27312 DVDD.n4976 DVDD.n681 0.0377541
R27313 DVDD.n787 DVDD.n749 0.0377541
R27314 DVDD.n4532 DVDD.n1082 0.0377541
R27315 DVDD.n5658 DVDD.n5657 0.0376798
R27316 DVDD.n5484 DVDD.n5483 0.0376798
R27317 DVDD.n5766 DVDD.n184 0.0373852
R27318 DVDD.n5220 DVDD.n490 0.0373852
R27319 DVDD.n648 DVDD.n620 0.0373852
R27320 DVDD.n844 DVDD.n709 0.0373852
R27321 DVDD.n4593 DVDD.n1014 0.0373852
R27322 DVDD.n1386 DVDD.n1307 0.0372431
R27323 DVDD.n1387 DVDD.n1311 0.0372431
R27324 DVDD.n1320 DVDD.n1219 0.0372431
R27325 DVDD.n1324 DVDD.n1221 0.0372431
R27326 DVDD.n154 DVDD.n142 0.0370164
R27327 DVDD.n473 DVDD.n461 0.0370164
R27328 DVDD.n4951 DVDD.n683 0.0370164
R27329 DVDD.n771 DVDD.n770 0.0370164
R27330 DVDD.n4509 DVDD.n1084 0.0370164
R27331 DVDD.n3245 DVDD.n3084 0.0369865
R27332 DVDD.n3201 DVDD.n3199 0.0369865
R27333 DVDD.n5777 DVDD.n182 0.0366475
R27334 DVDD.n5787 DVDD.n166 0.0366475
R27335 DVDD.n5847 DVDD.n135 0.0366475
R27336 DVDD.n5204 DVDD.n558 0.0366475
R27337 DVDD.n5198 DVDD.n556 0.0366475
R27338 DVDD.n5140 DVDD.n5139 0.0366475
R27339 DVDD.n664 DVDD.n618 0.0366475
R27340 DVDD.n5013 DVDD.n626 0.0366475
R27341 DVDD.n4994 DVDD.n424 0.0366475
R27342 DVDD.n828 DVDD.n718 0.0366475
R27343 DVDD.n822 DVDD.n716 0.0366475
R27344 DVDD.n758 DVDD.n400 0.0366475
R27345 DVDD.n4577 DVDD.n1049 0.0366475
R27346 DVDD.n4571 DVDD.n1047 0.0366475
R27347 DVDD.n4550 DVDD.n377 0.0366475
R27348 DVDD.n5772 DVDD.n171 0.0359098
R27349 DVDD.n5214 DVDD.n492 0.0359098
R27350 DVDD.n654 DVDD.n607 0.0359098
R27351 DVDD.n838 DVDD.n711 0.0359098
R27352 DVDD.n4587 DVDD.n1016 0.0359098
R27353 DVDD.n5803 DVDD.n157 0.035541
R27354 DVDD.n5159 DVDD.n472 0.035541
R27355 DVDD.n4982 DVDD.n4950 0.035541
R27356 DVDD.n780 DVDD.n779 0.035541
R27357 DVDD.n4538 DVDD.n4508 0.035541
R27358 DVDD.n3252 DVDD.n3086 0.0353649
R27359 DVDD.n3207 DVDD.n3122 0.0353649
R27360 DVDD.n5756 DVDD.n188 0.0351721
R27361 DVDD.n5230 DVDD.n563 0.0351721
R27362 DVDD.n638 DVDD.n623 0.0351721
R27363 DVDD.n854 DVDD.n723 0.0351721
R27364 DVDD.n4603 DVDD.n1054 0.0351721
R27365 DVDD.n5731 DVDD.n198 0.0348033
R27366 DVDD.n5819 DVDD.n149 0.0348033
R27367 DVDD.n5095 DVDD.n5094 0.0348033
R27368 DVDD.n5175 DVDD.n454 0.0348033
R27369 DVDD.n597 DVDD.n593 0.0348033
R27370 DVDD.n4966 DVDD.n677 0.0348033
R27371 DVDD.n876 DVDD.n735 0.0348033
R27372 DVDD.n798 DVDD.n797 0.0348033
R27373 DVDD.n1059 DVDD.n892 0.0348033
R27374 DVDD.n4522 DVDD.n1078 0.0348033
R27375 DVDD.n3235 DVDD.n3234 0.0345541
R27376 DVDD.n3164 DVDD.n3139 0.0345541
R27377 DVDD.n3232 DVDD.n3231 0.0344013
R27378 DVDD.n3227 DVDD.n3098 0.0344013
R27379 DVDD.n3170 DVDD.n3166 0.0344013
R27380 DVDD.n3167 DVDD.n3135 0.0344013
R27381 DVDD.n5835 DVDD.n164 0.0340656
R27382 DVDD.n5191 DVDD.n469 0.0340656
R27383 DVDD.n4947 DVDD.n673 0.0340656
R27384 DVDD.n815 DVDD.n814 0.0340656
R27385 DVDD.n4564 DVDD.n4563 0.0340656
R27386 DVDD.n1392 DVDD.n1309 0.0330202
R27387 DVDD.n1222 DVDD.n1214 0.0330202
R27388 DVDD.n5513 DVDD.n5512 0.0325451
R27389 DVDD.n4706 DVDD.n949 0.0325451
R27390 DVDD.n5733 DVDD.n198 0.0324979
R27391 DVDD.n5095 DVDD.n5089 0.0324979
R27392 DVDD.n596 DVDD.n593 0.0324979
R27393 DVDD.n878 DVDD.n735 0.0324979
R27394 DVDD.n896 DVDD.n892 0.0324979
R27395 DVDD.n1925 DVDD.n1923 0.03245
R27396 DVDD.n1926 DVDD.n1925 0.03245
R27397 DVDD.n3189 DVDD.n3133 0.03245
R27398 DVDD.n3193 DVDD.n3133 0.03245
R27399 DVDD.n3194 DVDD.n3193 0.03245
R27400 DVDD.n1924 DVDD.n1916 0.03245
R27401 DVDD.n1924 DVDD.n1921 0.03245
R27402 DVDD.n3676 DVDD.n1979 0.03245
R27403 DVDD.n3683 DVDD.n1979 0.03245
R27404 DVDD.n3685 DVDD.n3683 0.03245
R27405 DVDD.n3685 DVDD.n3684 0.03245
R27406 DVDD.n3684 DVDD.n1894 0.03245
R27407 DVDD.n3712 DVDD.n1894 0.03245
R27408 DVDD.n3713 DVDD.n3712 0.03245
R27409 DVDD.n3713 DVDD.n1888 0.03245
R27410 DVDD.n3721 DVDD.n1888 0.03245
R27411 DVDD.n3775 DVDD.n3755 0.03245
R27412 DVDD.n3763 DVDD.n3755 0.03245
R27413 DVDD.n3768 DVDD.n3763 0.03245
R27414 DVDD.n3768 DVDD.n3767 0.03245
R27415 DVDD.n3767 DVDD.n1664 0.03245
R27416 DVDD.n4292 DVDD.n1664 0.03245
R27417 DVDD.n4293 DVDD.n4292 0.03245
R27418 DVDD.n4293 DVDD.n1658 0.03245
R27419 DVDD.n4301 DVDD.n1658 0.03245
R27420 DVDD.n5737 DVDD.n193 0.0318525
R27421 DVDD.n5823 DVDD.n162 0.0318525
R27422 DVDD.n5097 DVDD.n569 0.0318525
R27423 DVDD.n5179 DVDD.n467 0.0318525
R27424 DVDD.n5021 DVDD.n594 0.0318525
R27425 DVDD.n4962 DVDD.n4945 0.0318525
R27426 DVDD.n872 DVDD.n737 0.0318525
R27427 DVDD.n804 DVDD.n803 0.0318525
R27428 DVDD.n1063 DVDD.n894 0.0318525
R27429 DVDD.n4518 DVDD.n4504 0.0318525
R27430 DVDD.n5849 DVDD.n135 0.0315574
R27431 DVDD.n5139 DVDD.n5138 0.0315574
R27432 DVDD.n428 DVDD.n424 0.0315574
R27433 DVDD.n404 DVDD.n400 0.0315574
R27434 DVDD.n381 DVDD.n377 0.0315574
R27435 DVDD.n3188 DVDD.n3134 0.03155
R27436 DVDD.n3187 DVDD.n3184 0.03155
R27437 DVDD.n3183 DVDD.n3132 0.03155
R27438 DVDD.n3196 DVDD.n3195 0.03155
R27439 DVDD.n5752 DVDD.n175 0.0314836
R27440 DVDD.n5234 DVDD.n487 0.0314836
R27441 DVDD.n634 DVDD.n611 0.0314836
R27442 DVDD.n858 DVDD.n706 0.0314836
R27443 DVDD.n4607 DVDD.n1011 0.0314836
R27444 DVDD.n5807 DVDD.n151 0.0311148
R27445 DVDD.n5163 DVDD.n465 0.0311148
R27446 DVDD.n4978 DVDD.n4943 0.0311148
R27447 DVDD.n786 DVDD.n785 0.0311148
R27448 DVDD.n4534 DVDD.n4502 0.0311148
R27449 DVDD.n2612 DVDD.n2505 0.0308261
R27450 DVDD.n2613 DVDD.n2612 0.0308261
R27451 DVDD.n2614 DVDD.n2613 0.0308261
R27452 DVDD.n2614 DVDD.n2503 0.0308261
R27453 DVDD.n2618 DVDD.n2503 0.0308261
R27454 DVDD.n2619 DVDD.n2618 0.0308261
R27455 DVDD.n2620 DVDD.n2619 0.0308261
R27456 DVDD.n2620 DVDD.n2501 0.0308261
R27457 DVDD.n2624 DVDD.n2501 0.0308261
R27458 DVDD.n2605 DVDD.n2507 0.0308261
R27459 DVDD.n5768 DVDD.n177 0.0307459
R27460 DVDD.n5218 DVDD.n561 0.0307459
R27461 DVDD.n650 DVDD.n613 0.0307459
R27462 DVDD.n842 DVDD.n721 0.0307459
R27463 DVDD.n4591 DVDD.n1052 0.0307459
R27464 DVDD.n5496 DVDD.n256 0.0305
R27465 DVDD.n5500 DVDD.n5499 0.0305
R27466 DVDD.n5495 DVDD.n5494 0.0305
R27467 DVDD.n5492 DVDD.n5491 0.0305
R27468 DVDD.n5838 DVDD.n5837 0.030377
R27469 DVDD.n5319 DVDD.n474 0.030377
R27470 DVDD.n5005 DVDD.n5004 0.030377
R27471 DVDD.n769 DVDD.n768 0.030377
R27472 DVDD.n4561 DVDD.n4560 0.030377
R27473 DVDD.n5775 DVDD.n179 0.0300082
R27474 DVDD.n5786 DVDD.n168 0.0300082
R27475 DVDD.n5845 DVDD.n138 0.0300082
R27476 DVDD.n5202 DVDD.n494 0.0300082
R27477 DVDD.n5200 DVDD.n495 0.0300082
R27478 DVDD.n5142 DVDD.n5141 0.0300082
R27479 DVDD.n666 DVDD.n615 0.0300082
R27480 DVDD.n668 DVDD.n606 0.0300082
R27481 DVDD.n4996 DVDD.n427 0.0300082
R27482 DVDD.n826 DVDD.n713 0.0300082
R27483 DVDD.n824 DVDD.n714 0.0300082
R27484 DVDD.n760 DVDD.n403 0.0300082
R27485 DVDD.n4575 DVDD.n1018 0.0300082
R27486 DVDD.n4573 DVDD.n1019 0.0300082
R27487 DVDD.n4552 DVDD.n380 0.0300082
R27488 DVDD.n1381 DVDD.n1312 0.0298119
R27489 DVDD.n1381 DVDD.n1308 0.0298119
R27490 DVDD.n1317 DVDD.n1217 0.0298119
R27491 DVDD.n1317 DVDD.n1215 0.0298119
R27492 DVDD.n5770 DVDD.n189 0.0292705
R27493 DVDD.n5216 DVDD.n560 0.0292705
R27494 DVDD.n652 DVDD.n624 0.0292705
R27495 DVDD.n840 DVDD.n720 0.0292705
R27496 DVDD.n4589 DVDD.n1051 0.0292705
R27497 DVDD.n937 DVDD.n936 0.0292629
R27498 DVDD.n956 DVDD.n955 0.0292629
R27499 DVDD.n5674 DVDD.n242 0.0292629
R27500 DVDD.n250 DVDD.n249 0.0292629
R27501 DVDD.n3232 DVDD.n3091 0.0291547
R27502 DVDD.n3242 DVDD.n3091 0.0291547
R27503 DVDD.n3243 DVDD.n3242 0.0291547
R27504 DVDD.n3243 DVDD.n3083 0.0291547
R27505 DVDD.n3186 DVDD.n3098 0.0291547
R27506 DVDD.n3186 DVDD.n3093 0.0291547
R27507 DVDD.n3093 DVDD.n3090 0.0291547
R27508 DVDD.n3090 DVDD.n3082 0.0291547
R27509 DVDD.n3166 DVDD.n3138 0.0291547
R27510 DVDD.n3140 DVDD.n3138 0.0291547
R27511 DVDD.n3140 DVDD.n3129 0.0291547
R27512 DVDD.n3129 DVDD.n3128 0.0291547
R27513 DVDD.n3182 DVDD.n3135 0.0291547
R27514 DVDD.n3182 DVDD.n3130 0.0291547
R27515 DVDD.n3197 DVDD.n3130 0.0291547
R27516 DVDD.n3197 DVDD.n3131 0.0291547
R27517 DVDD.n111 DVDD.n99 0.0290309
R27518 DVDD.n102 DVDD.n95 0.0290309
R27519 DVDD.n5409 DVDD.n338 0.0290309
R27520 DVDD.n349 DVDD.n342 0.0290309
R27521 DVDD.n940 DVDD.n916 0.0290309
R27522 DVDD.n958 DVDD.n923 0.0290309
R27523 DVDD.n5705 DVDD.n240 0.0290309
R27524 DVDD.n246 DVDD.n229 0.0290309
R27525 DVDD.n5805 DVDD.n152 0.0289016
R27526 DVDD.n5161 DVDD.n453 0.0289016
R27527 DVDD.n4980 DVDD.n676 0.0289016
R27528 DVDD.n783 DVDD.n751 0.0289016
R27529 DVDD.n4536 DVDD.n1077 0.0289016
R27530 DVDD.n5754 DVDD.n173 0.0285328
R27531 DVDD.n5232 DVDD.n488 0.0285328
R27532 DVDD.n636 DVDD.n609 0.0285328
R27533 DVDD.n856 DVDD.n707 0.0285328
R27534 DVDD.n4605 DVDD.n1012 0.0285328
R27535 DVDD.n2610 DVDD.n2609 0.0284
R27536 DVDD.n2611 DVDD.n2610 0.0284
R27537 DVDD.n2611 DVDD.n2504 0.0284
R27538 DVDD.n2615 DVDD.n2504 0.0284
R27539 DVDD.n2616 DVDD.n2615 0.0284
R27540 DVDD.n2617 DVDD.n2616 0.0284
R27541 DVDD.n2617 DVDD.n2502 0.0284
R27542 DVDD.n2621 DVDD.n2502 0.0284
R27543 DVDD.n2622 DVDD.n2621 0.0284
R27544 DVDD.n2623 DVDD.n2622 0.0284
R27545 DVDD.n5730 DVDD.n195 0.0281639
R27546 DVDD.n5821 DVDD.n161 0.0281639
R27547 DVDD.n5091 DVDD.n573 0.0281639
R27548 DVDD.n5177 DVDD.n470 0.0281639
R27549 DVDD.n599 DVDD.n590 0.0281639
R27550 DVDD.n4964 DVDD.n4948 0.0281639
R27551 DVDD.n874 DVDD.n738 0.0281639
R27552 DVDD.n800 DVDD.n799 0.0281639
R27553 DVDD.n1061 DVDD.n895 0.0281639
R27554 DVDD.n4520 DVDD.n4506 0.0281639
R27555 DVDD.n5498 DVDD.n5497 0.0277727
R27556 DVDD.n5493 DVDD.n262 0.0277727
R27557 DVDD.n5792 DVDD.n145 0.0274262
R27558 DVDD.n5194 DVDD.n456 0.0274262
R27559 DVDD.n5008 DVDD.n5007 0.0274262
R27560 DVDD.n818 DVDD.n740 0.0274262
R27561 DVDD.n4567 DVDD.n1071 0.0274262
R27562 DVDD.n1927 DVDD.n1926 0.027126
R27563 DVDD.n2709 DVDD.n2702 0.0271068
R27564 DVDD.n1393 DVDD.n1392 0.0270348
R27565 DVDD.n1555 DVDD.n1222 0.0270348
R27566 DVDD.n3279 DVDD.n3277 0.026913
R27567 DVDD.n3279 DVDD.n3278 0.026913
R27568 DVDD.n3278 DVDD.n2925 0.026913
R27569 DVDD.n3298 DVDD.n2925 0.026913
R27570 DVDD.n3299 DVDD.n3298 0.026913
R27571 DVDD.n3300 DVDD.n3299 0.026913
R27572 DVDD.n3300 DVDD.n2916 0.026913
R27573 DVDD.n3327 DVDD.n2916 0.026913
R27574 DVDD.n3328 DVDD.n3327 0.026913
R27575 DVDD.n3328 DVDD.n2914 0.026913
R27576 DVDD.n3332 DVDD.n2914 0.026913
R27577 DVDD.n3280 DVDD.n2926 0.026913
R27578 DVDD.n3301 DVDD.n2924 0.026913
R27579 DVDD.n3301 DVDD.n2917 0.026913
R27580 DVDD.n3330 DVDD.n3329 0.026913
R27581 DVDD.n3331 DVDD.n3330 0.026913
R27582 DVDD.n2943 DVDD.n2763 0.026913
R27583 DVDD.n2805 DVDD.n2767 0.026913
R27584 DVDD.n2806 DVDD.n2805 0.026913
R27585 DVDD.n2814 DVDD.n2813 0.026913
R27586 DVDD.n2815 DVDD.n2814 0.026913
R27587 DVDD.n2950 DVDD.n2937 0.026913
R27588 DVDD.n3276 DVDD.n2953 0.026913
R27589 DVDD.n2942 DVDD.n2941 0.026913
R27590 DVDD.n2942 DVDD.n2765 0.026913
R27591 DVDD.n3369 DVDD.n2765 0.026913
R27592 DVDD.n3369 DVDD.n3368 0.026913
R27593 DVDD.n3368 DVDD.n2766 0.026913
R27594 DVDD.n2804 DVDD.n2766 0.026913
R27595 DVDD.n2804 DVDD.n2803 0.026913
R27596 DVDD.n2811 DVDD.n2803 0.026913
R27597 DVDD.n2812 DVDD.n2811 0.026913
R27598 DVDD.n2812 DVDD.n2800 0.026913
R27599 DVDD.n2816 DVDD.n2800 0.026913
R27600 DVDD.n2819 DVDD.n2790 0.026913
R27601 DVDD.n2823 DVDD.n2822 0.026913
R27602 DVDD.n2831 DVDD.n2830 0.026913
R27603 DVDD.n2839 DVDD.n2838 0.026913
R27604 DVDD.n2847 DVDD.n2846 0.026913
R27605 DVDD.n2855 DVDD.n2798 0.026913
R27606 DVDD.n2820 DVDD.n2818 0.026913
R27607 DVDD.n2824 DVDD.n2821 0.026913
R27608 DVDD.n2826 DVDD.n2824 0.026913
R27609 DVDD.n2828 DVDD.n2826 0.026913
R27610 DVDD.n2829 DVDD.n2828 0.026913
R27611 DVDD.n2832 DVDD.n2829 0.026913
R27612 DVDD.n2834 DVDD.n2832 0.026913
R27613 DVDD.n2836 DVDD.n2834 0.026913
R27614 DVDD.n2837 DVDD.n2836 0.026913
R27615 DVDD.n2840 DVDD.n2837 0.026913
R27616 DVDD.n2842 DVDD.n2840 0.026913
R27617 DVDD.n2844 DVDD.n2842 0.026913
R27618 DVDD.n2845 DVDD.n2844 0.026913
R27619 DVDD.n2848 DVDD.n2845 0.026913
R27620 DVDD.n2850 DVDD.n2848 0.026913
R27621 DVDD.n2852 DVDD.n2850 0.026913
R27622 DVDD.n2854 DVDD.n2852 0.026913
R27623 DVDD.n2856 DVDD.n2854 0.026913
R27624 DVDD.n2857 DVDD.n2856 0.026913
R27625 DVDD.n3344 DVDD.n2857 0.026913
R27626 DVDD.n3343 DVDD.n2858 0.026913
R27627 DVDD.n2882 DVDD.n2858 0.026913
R27628 DVDD.n2884 DVDD.n2882 0.026913
R27629 DVDD.n2886 DVDD.n2884 0.026913
R27630 DVDD.n2888 DVDD.n2886 0.026913
R27631 DVDD.n2889 DVDD.n2888 0.026913
R27632 DVDD.n2892 DVDD.n2889 0.026913
R27633 DVDD.n2894 DVDD.n2892 0.026913
R27634 DVDD.n2896 DVDD.n2894 0.026913
R27635 DVDD.n2897 DVDD.n2896 0.026913
R27636 DVDD.n2900 DVDD.n2897 0.026913
R27637 DVDD.n2902 DVDD.n2900 0.026913
R27638 DVDD.n2904 DVDD.n2902 0.026913
R27639 DVDD.n2905 DVDD.n2904 0.026913
R27640 DVDD.n2908 DVDD.n2905 0.026913
R27641 DVDD.n2910 DVDD.n2908 0.026913
R27642 DVDD.n2912 DVDD.n2910 0.026913
R27643 DVDD.n2913 DVDD.n2912 0.026913
R27644 DVDD.n3336 DVDD.n3334 0.026913
R27645 DVDD.n2881 DVDD.n2860 0.026913
R27646 DVDD.n2891 DVDD.n2890 0.026913
R27647 DVDD.n2899 DVDD.n2898 0.026913
R27648 DVDD.n2907 DVDD.n2906 0.026913
R27649 DVDD.n3338 DVDD.n2880 0.026913
R27650 DVDD.n3335 DVDD.n2873 0.026913
R27651 DVDD.n2668 DVDD.n2625 0.026913
R27652 DVDD.n2668 DVDD.n2667 0.026913
R27653 DVDD.n2667 DVDD.n2664 0.026913
R27654 DVDD.n2664 DVDD.n2663 0.026913
R27655 DVDD.n2663 DVDD.n2661 0.026913
R27656 DVDD.n2661 DVDD.n2659 0.026913
R27657 DVDD.n2659 DVDD.n2657 0.026913
R27658 DVDD.n2657 DVDD.n2654 0.026913
R27659 DVDD.n2654 DVDD.n2653 0.026913
R27660 DVDD.n2628 DVDD.n2453 0.026913
R27661 DVDD.n2630 DVDD.n2628 0.026913
R27662 DVDD.n2631 DVDD.n2630 0.026913
R27663 DVDD.n2634 DVDD.n2631 0.026913
R27664 DVDD.n2636 DVDD.n2634 0.026913
R27665 DVDD.n2638 DVDD.n2636 0.026913
R27666 DVDD.n2639 DVDD.n2638 0.026913
R27667 DVDD.n2642 DVDD.n2639 0.026913
R27668 DVDD.n2644 DVDD.n2642 0.026913
R27669 DVDD.n2608 DVDD.n2508 0.026913
R27670 DVDD.n2633 DVDD.n2632 0.026913
R27671 DVDD.n2641 DVDD.n2640 0.026913
R27672 DVDD.n1385 DVDD.n1384 0.0264516
R27673 DVDD.n1322 DVDD.n1319 0.0264516
R27674 DVDD.n1321 DVDD.n1319 0.0264516
R27675 DVDD.n1384 DVDD.n1383 0.0264516
R27676 DVDD.n3174 DVDD.n3173 0.0264459
R27677 DVDD.n3236 DVDD.n3095 0.0264459
R27678 DVDD DVDD.n2913 0.0264239
R27679 DVDD.n2626 DVDD.n2443 0.0264239
R27680 DVDD.n2849 DVDD.n2796 0.0261793
R27681 DVDD.n2853 DVDD.n2781 0.0261793
R27682 DVDD.n2883 DVDD.n2869 0.0261793
R27683 DVDD.n2887 DVDD.n2875 0.0261793
R27684 DVDD.n2643 DVDD.n2451 0.0259348
R27685 DVDD.n3203 DVDD.n3202 0.0256351
R27686 DVDD.n3249 DVDD.n3248 0.0256351
R27687 DVDD.n2708 DVDD.n2702 0.0255998
R27688 DVDD.n2750 DVDD.n2734 0.0255952
R27689 DVDD.n3292 DVDD.n3291 0.0254457
R27690 DVDD.n3371 DVDD.n3370 0.0254457
R27691 DVDD.n5912 DVDD.n91 0.0253196
R27692 DVDD.n114 DVDD.n93 0.0253196
R27693 DVDD.n5415 DVDD.n345 0.0253196
R27694 DVDD.n5412 DVDD.n347 0.0253196
R27695 DVDD.n933 DVDD.n926 0.0253196
R27696 DVDD.n952 DVDD.n919 0.0253196
R27697 DVDD.n5670 DVDD.n232 0.0253196
R27698 DVDD.n252 DVDD.n238 0.0253196
R27699 DVDD.n5736 DVDD.n195 0.0252131
R27700 DVDD.n5821 DVDD.n148 0.0252131
R27701 DVDD.n5091 DVDD.n5088 0.0252131
R27702 DVDD.n5177 DVDD.n458 0.0252131
R27703 DVDD.n599 DVDD.n592 0.0252131
R27704 DVDD.n4964 DVDD.n680 0.0252131
R27705 DVDD.n874 DVDD.n736 0.0252131
R27706 DVDD.n800 DVDD.n745 0.0252131
R27707 DVDD.n1061 DVDD.n893 0.0252131
R27708 DVDD.n4520 DVDD.n1081 0.0252131
R27709 DVDD.n3118 DVDD.n3083 0.024917
R27710 DVDD.n3212 DVDD.n3082 0.024917
R27711 DVDD.n3128 DVDD.n3121 0.024917
R27712 DVDD.n3131 DVDD.n3120 0.024917
R27713 DVDD.n5913 DVDD.n89 0.0248557
R27714 DVDD.n109 DVDD.n94 0.0248557
R27715 DVDD.n5416 DVDD.n343 0.0248557
R27716 DVDD.n5419 DVDD.n352 0.0248557
R27717 DVDD.n941 DVDD.n927 0.0248557
R27718 DVDD.n942 DVDD.n920 0.0248557
R27719 DVDD.n257 DVDD.n233 0.0248557
R27720 DVDD.n244 DVDD.n239 0.0248557
R27721 DVDD.n5754 DVDD.n185 0.0248443
R27722 DVDD.n5232 DVDD.n564 0.0248443
R27723 DVDD.n636 DVDD.n621 0.0248443
R27724 DVDD.n856 DVDD.n724 0.0248443
R27725 DVDD.n4605 DVDD.n1055 0.0248443
R27726 DVDD.n2666 DVDD.n2665 0.0248
R27727 DVDD.n2656 DVDD.n2655 0.0248
R27728 DVDD.n2750 DVDD.n2735 0.0247609
R27729 DVDD.n2512 DVDD 0.0247148
R27730 DVDD.n2841 DVDD.n2784 0.024712
R27731 DVDD.n2895 DVDD.n2866 0.024712
R27732 DVDD.n5805 DVDD.n158 0.0244754
R27733 DVDD.n5161 DVDD.n460 0.0244754
R27734 DVDD.n4980 DVDD.n682 0.0244754
R27735 DVDD.n784 DVDD.n783 0.0244754
R27736 DVDD.n4536 DVDD.n1083 0.0244754
R27737 DVDD.n2635 DVDD.n2446 0.0244674
R27738 DVDD.n2662 DVDD.n2496 0.02435
R27739 DVDD.n5770 DVDD.n183 0.0241066
R27740 DVDD.n5216 DVDD.n491 0.0241066
R27741 DVDD.n652 DVDD.n619 0.0241066
R27742 DVDD.n840 DVDD.n710 0.0241066
R27743 DVDD.n4589 DVDD.n1015 0.0241066
R27744 DVDD.n3235 DVDD.n3094 0.0240135
R27745 DVDD.n3180 DVDD.n3139 0.0240135
R27746 DVDD.n1370 DVDD.n1329 0.024
R27747 DVDD.n3274 DVDD.n3272 0.0239783
R27748 DVDD.n2949 DVDD.n2939 0.0239783
R27749 DVDD.n2658 DVDD.n2492 0.0239
R27750 DVDD.n2016 DVDD 0.0238333
R27751 DVDD.n2015 DVDD 0.0238333
R27752 DVDD.n2020 DVDD 0.0238333
R27753 DVDD.n2019 DVDD 0.0238333
R27754 DVDD.n2024 DVDD 0.0238333
R27755 DVDD.n2023 DVDD 0.0238333
R27756 DVDD.n2028 DVDD 0.0238333
R27757 DVDD.n2027 DVDD 0.0238333
R27758 DVDD.n2032 DVDD 0.0238333
R27759 DVDD.n2031 DVDD 0.0238333
R27760 DVDD.n2036 DVDD 0.0238333
R27761 DVDD.n2035 DVDD 0.0238333
R27762 DVDD DVDD.n2038 0.0238333
R27763 DVDD.n5841 DVDD.n140 0.0237377
R27764 DVDD.n5147 DVDD.n463 0.0237377
R27765 DVDD.n5001 DVDD.n4941 0.0237377
R27766 DVDD.n765 DVDD.n756 0.0237377
R27767 DVDD.n4557 DVDD.n4500 0.0237377
R27768 DVDD.n5775 DVDD.n181 0.0233689
R27769 DVDD.n181 DVDD.n168 0.0233689
R27770 DVDD.n5843 DVDD.n136 0.0233689
R27771 DVDD.n5845 DVDD.n136 0.0233689
R27772 DVDD.n5202 DVDD.n557 0.0233689
R27773 DVDD.n5200 DVDD.n557 0.0233689
R27774 DVDD.n5145 DVDD.n5104 0.0233689
R27775 DVDD.n5142 DVDD.n5104 0.0233689
R27776 DVDD.n666 DVDD.n617 0.0233689
R27777 DVDD.n668 DVDD.n617 0.0233689
R27778 DVDD.n4999 DVDD.n425 0.0233689
R27779 DVDD.n4996 DVDD.n425 0.0233689
R27780 DVDD.n826 DVDD.n717 0.0233689
R27781 DVDD.n824 DVDD.n717 0.0233689
R27782 DVDD.n763 DVDD.n401 0.0233689
R27783 DVDD.n760 DVDD.n401 0.0233689
R27784 DVDD.n4575 DVDD.n1048 0.0233689
R27785 DVDD.n4573 DVDD.n1048 0.0233689
R27786 DVDD.n4555 DVDD.n378 0.0233689
R27787 DVDD.n4552 DVDD.n378 0.0233689
R27788 DVDD.n2833 DVDD.n2793 0.0232446
R27789 DVDD.n2903 DVDD.n2878 0.0232446
R27790 DVDD.n3253 DVDD.n3252 0.0232027
R27791 DVDD.n3200 DVDD.n3122 0.0232027
R27792 DVDD.n5838 DVDD.n140 0.023
R27793 DVDD.n474 DVDD.n463 0.023
R27794 DVDD.n5004 DVDD.n4941 0.023
R27795 DVDD.n768 DVDD.n756 0.023
R27796 DVDD.n4560 DVDD.n4500 0.023
R27797 DVDD.n3602 DVDD.n2454 0.023
R27798 DVDD.n2715 DVDD.n2702 0.0229382
R27799 DVDD.n1741 DVDD.n1739 0.0229381
R27800 DVDD.n2750 DVDD.n2742 0.0227712
R27801 DVDD.n1898 DVDD.n1896 0.0227688
R27802 DVDD.n5768 DVDD.n183 0.0226311
R27803 DVDD.n5218 DVDD.n491 0.0226311
R27804 DVDD.n650 DVDD.n619 0.0226311
R27805 DVDD.n842 DVDD.n710 0.0226311
R27806 DVDD.n4591 DVDD.n1015 0.0226311
R27807 DVDD.n2817 DVDD.n2789 0.0225217
R27808 DVDD.n3333 DVDD.n2870 0.0225217
R27809 DVDD.n5850 DVDD.n5849 0.0224209
R27810 DVDD.n5138 DVDD.n5137 0.0224209
R27811 DVDD.n5341 DVDD.n428 0.0224209
R27812 DVDD.n5362 DVDD.n404 0.0224209
R27813 DVDD.n5382 DVDD.n381 0.0224209
R27814 DVDD.n3203 DVDD.n3123 0.0223919
R27815 DVDD.n3205 DVDD.n3203 0.0223919
R27816 DVDD.n3249 DVDD.n3085 0.0223919
R27817 DVDD.n3251 DVDD.n3249 0.0223919
R27818 DVDD.n1742 DVDD 0.0223846
R27819 DVDD.n1386 DVDD.n1312 0.0223807
R27820 DVDD.n1387 DVDD.n1308 0.0223807
R27821 DVDD.n1320 DVDD.n1217 0.0223807
R27822 DVDD.n1324 DVDD.n1215 0.0223807
R27823 DVDD.n2827 DVDD.n2786 0.0222663
R27824 DVDD.n2909 DVDD.n2864 0.0222663
R27825 DVDD.n5807 DVDD.n158 0.0222623
R27826 DVDD.n5163 DVDD.n460 0.0222623
R27827 DVDD.n4978 DVDD.n682 0.0222623
R27828 DVDD.n785 DVDD.n784 0.0222623
R27829 DVDD.n4534 DVDD.n1083 0.0222623
R27830 DVDD.n5752 DVDD.n185 0.0218934
R27831 DVDD.n5234 DVDD.n564 0.0218934
R27832 DVDD.n634 DVDD.n621 0.0218934
R27833 DVDD.n858 DVDD.n724 0.0218934
R27834 DVDD.n4607 DVDD.n1055 0.0218934
R27835 DVDD.n1922 DVDD.n1901 0.0218
R27836 DVDD.n3192 DVDD.n3191 0.0218
R27837 DVDD.n3192 DVDD.n2738 0.0218
R27838 DVDD.n2825 DVDD.n2787 0.0217772
R27839 DVDD.n2911 DVDD.n2863 0.0217772
R27840 DVDD.n3253 DVDD.n3084 0.0215811
R27841 DVDD.n3201 DVDD.n3200 0.0215811
R27842 DVDD.n5737 DVDD.n5736 0.0215246
R27843 DVDD.n5823 DVDD.n148 0.0215246
R27844 DVDD.n5088 DVDD.n569 0.0215246
R27845 DVDD.n5179 DVDD.n458 0.0215246
R27846 DVDD.n594 DVDD.n592 0.0215246
R27847 DVDD.n4962 DVDD.n680 0.0215246
R27848 DVDD.n872 DVDD.n736 0.0215246
R27849 DVDD.n803 DVDD.n745 0.0215246
R27850 DVDD.n1063 DVDD.n893 0.0215246
R27851 DVDD.n4518 DVDD.n1081 0.0215246
R27852 DVDD.n5734 DVDD.n5733 0.0215141
R27853 DVDD.n5089 DVDD.n572 0.0215141
R27854 DVDD.n596 DVDD.n589 0.0215141
R27855 DVDD.n4774 DVDD.n878 0.0215141
R27856 DVDD.n4745 DVDD.n896 0.0215141
R27857 DVDD.n112 DVDD.n97 0.0211443
R27858 DVDD.n5910 DVDD.n96 0.0211443
R27859 DVDD.n5410 DVDD.n336 0.0211443
R27860 DVDD.n5413 DVDD.n335 0.0211443
R27861 DVDD.n931 DVDD.n917 0.0211443
R27862 DVDD.n950 DVDD.n924 0.0211443
R27863 DVDD.n5668 DVDD.n236 0.0211443
R27864 DVDD.n254 DVDD.n230 0.0211443
R27865 DVDD.n2629 DVDD.n2449 0.0210435
R27866 DVDD.n2716 DVDD 0.0209763
R27867 DVDD.n5955 DVDD.n28 0.0209627
R27868 DVDD.n4702 DVDD.n4701 0.0209627
R27869 DVDD.n2835 DVDD.n2794 0.0207989
R27870 DVDD.n2901 DVDD.n2877 0.0207989
R27871 DVDD.n3239 DVDD.n3094 0.0207703
R27872 DVDD.n3180 DVDD.n3179 0.0207703
R27873 DVDD.n110 DVDD.n100 0.0206804
R27874 DVDD.n5916 DVDD.n5915 0.0206804
R27875 DVDD.n5408 DVDD.n339 0.0206804
R27876 DVDD.n5418 DVDD.n341 0.0206804
R27877 DVDD.n1886 DVDD.n1861 0.020525
R27878 DVDD.n1954 DVDD 0.0204408
R27879 DVDD.n2963 DVDD 0.0202739
R27880 DVDD.n3061 DVDD.n3000 0.0201875
R27881 DVDD.n3009 DVDD.n3000 0.0201875
R27882 DVDD.n3054 DVDD.n3009 0.0201875
R27883 DVDD.n3054 DVDD.n3053 0.0201875
R27884 DVDD.n3053 DVDD.n3010 0.0201875
R27885 DVDD.n3046 DVDD.n3010 0.0201875
R27886 DVDD.n3046 DVDD.n3045 0.0201875
R27887 DVDD.n3281 DVDD.n2932 0.0200652
R27888 DVDD.n2944 DVDD.n2940 0.0200652
R27889 DVDD.n5617 DVDD.n5616 0.0197083
R27890 DVDD.n5517 DVDD.n30 0.0197083
R27891 DVDD.n5533 DVDD.n5532 0.0197083
R27892 DVDD.n5550 DVDD.n5549 0.0197083
R27893 DVDD.n4656 DVDD.n973 0.0197083
R27894 DVDD.n4685 DVDD.n4684 0.0197083
R27895 DVDD.n4668 DVDD.n4667 0.0197083
R27896 DVDD.n5442 DVDD.n5441 0.0197083
R27897 DVDD.n2637 DVDD.n2445 0.0195761
R27898 DVDD.n5650 DVDD.n5611 0.0193985
R27899 DVDD.n317 DVDD.n293 0.0193985
R27900 DVDD.n2843 DVDD.n2783 0.0193315
R27901 DVDD.n2893 DVDD.n2867 0.0193315
R27902 DVDD.n164 DVDD.n145 0.0193115
R27903 DVDD.n5191 DVDD.n456 0.0193115
R27904 DVDD.n5007 DVDD.n673 0.0193115
R27905 DVDD.n815 DVDD.n740 0.0193115
R27906 DVDD.n4564 DVDD.n1071 0.0193115
R27907 DVDD.n5646 DVDD.n50 0.0192435
R27908 DVDD.n5473 DVDD.n5472 0.0192435
R27909 DVDD.n5519 DVDD.n27 0.0190886
R27910 DVDD.n4699 DVDD.n4698 0.0190886
R27911 DVDD.n5629 DVDD.n63 0.0189337
R27912 DVDD.n5454 DVDD.n302 0.0189337
R27913 DVDD.n5535 DVDD.n12 0.0187788
R27914 DVDD.n4681 DVDD.n979 0.0187788
R27915 DVDD.n1339 DVDD.n1338 0.0186803
R27916 DVDD.n1341 DVDD.n1335 0.0186803
R27917 DVDD.n1335 DVDD.n1334 0.0186803
R27918 DVDD.n1332 DVDD.n1330 0.0186803
R27919 DVDD.n1365 DVDD.n1333 0.0186803
R27920 DVDD.n1367 DVDD.n1366 0.0186803
R27921 DVDD.n1334 DVDD.n1329 0.0186803
R27922 DVDD.n1366 DVDD.n1365 0.0186803
R27923 DVDD.n1369 DVDD.n1330 0.0186803
R27924 DVDD.n1341 DVDD.n1339 0.0186803
R27925 DVDD.n1338 DVDD.n1336 0.0186803
R27926 DVDD.n1333 DVDD.n1332 0.0186803
R27927 DVDD.n5613 DVDD.n57 0.0186239
R27928 DVDD.n5438 DVDD.n309 0.0186239
R27929 DVDD.n3297 DVDD.n3296 0.0185978
R27930 DVDD.n3326 DVDD.n3325 0.0185978
R27931 DVDD.n3367 DVDD.n3366 0.0185978
R27932 DVDD.n2810 DVDD.n2809 0.0185978
R27933 DVDD.n5731 DVDD.n5730 0.0185738
R27934 DVDD.n5819 DVDD.n161 0.0185738
R27935 DVDD.n5094 DVDD.n573 0.0185738
R27936 DVDD.n5175 DVDD.n470 0.0185738
R27937 DVDD.n597 DVDD.n590 0.0185738
R27938 DVDD.n4966 DVDD.n4948 0.0185738
R27939 DVDD.n876 DVDD.n738 0.0185738
R27940 DVDD.n799 DVDD.n798 0.0185738
R27941 DVDD.n1059 DVDD.n895 0.0185738
R27942 DVDD.n4522 DVDD.n4506 0.0185738
R27943 DVDD.n5921 DVDD.n83 0.018469
R27944 DVDD.n5552 DVDD.n20 0.018469
R27945 DVDD.n4664 DVDD.n4649 0.018469
R27946 DVDD.n5427 DVDD.n327 0.018469
R27947 DVDD.n3345 DVDD.n2791 0.0182974
R27948 DVDD.n3339 DVDD.n2871 0.0182974
R27949 DVDD.n3340 DVDD.n3339 0.0182974
R27950 DVDD.n3345 DVDD.n2788 0.0182974
R27951 DVDD.n5756 DVDD.n173 0.0182049
R27952 DVDD.n5230 DVDD.n488 0.0182049
R27953 DVDD.n638 DVDD.n609 0.0182049
R27954 DVDD.n854 DVDD.n707 0.0182049
R27955 DVDD.n4603 DVDD.n1012 0.0182049
R27956 DVDD.n5546 DVDD.n15 0.0181592
R27957 DVDD.n4670 DVDD.n982 0.0181592
R27958 DVDD.n2649 DVDD.n2452 0.0181087
R27959 DVDD.n2652 DVDD.n2498 0.01805
R27960 DVDD.n2851 DVDD.n2782 0.0178641
R27961 DVDD.n2851 DVDD.n2797 0.0178641
R27962 DVDD.n2885 DVDD.n2874 0.0178641
R27963 DVDD.n2885 DVDD.n2868 0.0178641
R27964 DVDD.n5634 DVDD.n5633 0.0178494
R27965 DVDD.n5529 DVDD.n24 0.0178494
R27966 DVDD.n4687 DVDD.n4653 0.0178494
R27967 DVDD.n5459 DVDD.n5458 0.0178494
R27968 DVDD.n5803 DVDD.n152 0.0178361
R27969 DVDD.n5159 DVDD.n453 0.0178361
R27970 DVDD.n4982 DVDD.n676 0.0178361
R27971 DVDD.n780 DVDD.n751 0.0178361
R27972 DVDD.n4538 DVDD.n1077 0.0178361
R27973 DVDD.n5708 DVDD.n225 0.0176945
R27974 DVDD.n962 DVDD.n944 0.0176945
R27975 DVDD.n1379 DVDD.n1378 0.0176362
R27976 DVDD.n2649 DVDD.n2444 0.0176196
R27977 DVDD.n2669 DVDD.n2494 0.0176
R27978 DVDD.n5772 DVDD.n189 0.0174672
R27979 DVDD.n5214 DVDD.n560 0.0174672
R27980 DVDD.n654 DVDD.n624 0.0174672
R27981 DVDD.n838 DVDD.n720 0.0174672
R27982 DVDD.n4587 DVDD.n1051 0.0174672
R27983 DVDD.n3194 DVDD.n2750 0.017375
R27984 DVDD.n5619 DVDD.n5575 0.0172298
R27985 DVDD.n5444 DVDD.n282 0.0172298
R27986 DVDD.n3297 DVDD.n3295 0.0171304
R27987 DVDD.n3326 DVDD.n2915 0.0171304
R27988 DVDD.n3367 DVDD.n2764 0.0171304
R27989 DVDD.n2810 DVDD.n2802 0.0171304
R27990 DVDD.n5661 DVDD.n5660 0.0170354
R27991 DVDD.n5487 DVDD.n5486 0.0170354
R27992 DVDD.n5911 DVDD.n92 0.0169691
R27993 DVDD.n113 DVDD.n92 0.0169691
R27994 DVDD.n5414 DVDD.n346 0.0169691
R27995 DVDD.n5411 DVDD.n346 0.0169691
R27996 DVDD.n929 DVDD.n925 0.0169691
R27997 DVDD.n929 DVDD.n918 0.0169691
R27998 DVDD.n5666 DVDD.n231 0.0169691
R27999 DVDD.n5666 DVDD.n237 0.0169691
R28000 DVDD.n5636 DVDD.n5608 0.01692
R28001 DVDD.n5461 DVDD.n290 0.01692
R28002 DVDD.n2403 DVDD.n2402 0.0169185
R28003 DVDD.n2012 DVDD.n2011 0.0169185
R28004 DVDD.n2040 DVDD.n2012 0.0169185
R28005 DVDD.n2010 DVDD.n2009 0.0169185
R28006 DVDD.n2041 DVDD.n2010 0.0169185
R28007 DVDD.n2008 DVDD.n2007 0.0169185
R28008 DVDD.n2042 DVDD.n2008 0.0169185
R28009 DVDD.n2006 DVDD.n2005 0.0169185
R28010 DVDD.n2006 DVDD.n1998 0.0169185
R28011 DVDD.n3672 DVDD.n1984 0.0169185
R28012 DVDD.n1996 DVDD.n1995 0.0169185
R28013 DVDD.n3668 DVDD.n1985 0.0169185
R28014 DVDD.n1994 DVDD.n1993 0.0169185
R28015 DVDD.n3669 DVDD.n1986 0.0169185
R28016 DVDD.n1992 DVDD.n1991 0.0169185
R28017 DVDD.n3670 DVDD.n1987 0.0169185
R28018 DVDD.n1990 DVDD.n1989 0.0169185
R28019 DVDD.n3675 DVDD.n1981 0.0169185
R28020 DVDD.n3732 DVDD.n3722 0.0169185
R28021 DVDD.n3732 DVDD.n1857 0.0169185
R28022 DVDD.n3753 DVDD.n3731 0.0169185
R28023 DVDD.n3731 DVDD.n1858 0.0169185
R28024 DVDD.n3752 DVDD.n3730 0.0169185
R28025 DVDD.n3730 DVDD.n1859 0.0169185
R28026 DVDD.n3751 DVDD.n3729 0.0169185
R28027 DVDD.n3729 DVDD.n1860 0.0169185
R28028 DVDD.n3750 DVDD.n1861 0.0169185
R28029 DVDD.n3749 DVDD.n3728 0.0169185
R28030 DVDD.n3728 DVDD.n1862 0.0169185
R28031 DVDD.n3748 DVDD.n3727 0.0169185
R28032 DVDD.n3727 DVDD.n1863 0.0169185
R28033 DVDD.n3747 DVDD.n3726 0.0169185
R28034 DVDD.n3726 DVDD.n1864 0.0169185
R28035 DVDD.n3746 DVDD.n3725 0.0169185
R28036 DVDD.n3725 DVDD.n1865 0.0169185
R28037 DVDD.n3745 DVDD.n3724 0.0169185
R28038 DVDD.n3724 DVDD.n1866 0.0169185
R28039 DVDD.n4343 DVDD.n1629 0.0169185
R28040 DVDD.n4341 DVDD.n1657 0.0169185
R28041 DVDD.n1656 DVDD.n1630 0.0169185
R28042 DVDD.n4340 DVDD.n1655 0.0169185
R28043 DVDD.n1654 DVDD.n1631 0.0169185
R28044 DVDD.n4339 DVDD.n1653 0.0169185
R28045 DVDD.n1652 DVDD.n1632 0.0169185
R28046 DVDD.n4338 DVDD.n1651 0.0169185
R28047 DVDD.n1650 DVDD.n1633 0.0169185
R28048 DVDD.n4337 DVDD.n1649 0.0169185
R28049 DVDD.n1648 DVDD.n1634 0.0169185
R28050 DVDD.n4336 DVDD.n1647 0.0169185
R28051 DVDD.n1646 DVDD.n1635 0.0169185
R28052 DVDD.n4335 DVDD.n1645 0.0169185
R28053 DVDD.n1644 DVDD.n1636 0.0169185
R28054 DVDD.n4334 DVDD.n1643 0.0169185
R28055 DVDD.n1642 DVDD.n1637 0.0169185
R28056 DVDD.n4333 DVDD.n1641 0.0169185
R28057 DVDD.n1640 DVDD.n1638 0.0169185
R28058 DVDD.n4346 DVDD.n1626 0.0169185
R28059 DVDD.n4386 DVDD.n1597 0.0169185
R28060 DVDD.n4384 DVDD.n1625 0.0169185
R28061 DVDD.n1624 DVDD.n1598 0.0169185
R28062 DVDD.n4383 DVDD.n1623 0.0169185
R28063 DVDD.n1622 DVDD.n1599 0.0169185
R28064 DVDD.n4382 DVDD.n1621 0.0169185
R28065 DVDD.n1620 DVDD.n1600 0.0169185
R28066 DVDD.n4381 DVDD.n1619 0.0169185
R28067 DVDD.n1618 DVDD.n1601 0.0169185
R28068 DVDD.n4380 DVDD.n1617 0.0169185
R28069 DVDD.n1616 DVDD.n1602 0.0169185
R28070 DVDD.n4379 DVDD.n1615 0.0169185
R28071 DVDD.n1614 DVDD.n1603 0.0169185
R28072 DVDD.n4378 DVDD.n1613 0.0169185
R28073 DVDD.n1612 DVDD.n1604 0.0169185
R28074 DVDD.n4377 DVDD.n1611 0.0169185
R28075 DVDD.n1610 DVDD.n1605 0.0169185
R28076 DVDD.n4376 DVDD.n1609 0.0169185
R28077 DVDD.n1608 DVDD.n1606 0.0169185
R28078 DVDD.n4389 DVDD.n1594 0.0169185
R28079 DVDD.n4414 DVDD.n1109 0.0169185
R28080 DVDD.n4399 DVDD.n1593 0.0169185
R28081 DVDD.n4402 DVDD.n1110 0.0169185
R28082 DVDD.n4398 DVDD.n1592 0.0169185
R28083 DVDD.n4403 DVDD.n1111 0.0169185
R28084 DVDD.n4397 DVDD.n1591 0.0169185
R28085 DVDD.n4404 DVDD.n1112 0.0169185
R28086 DVDD.n4396 DVDD.n1590 0.0169185
R28087 DVDD.n4405 DVDD.n1113 0.0169185
R28088 DVDD.n4395 DVDD.n1589 0.0169185
R28089 DVDD.n4406 DVDD.n1114 0.0169185
R28090 DVDD.n4394 DVDD.n1588 0.0169185
R28091 DVDD.n4407 DVDD.n1115 0.0169185
R28092 DVDD.n4393 DVDD.n1587 0.0169185
R28093 DVDD.n4408 DVDD.n1116 0.0169185
R28094 DVDD.n4392 DVDD.n1586 0.0169185
R28095 DVDD.n4409 DVDD.n1117 0.0169185
R28096 DVDD.n4391 DVDD.n1585 0.0169185
R28097 DVDD.n4410 DVDD.n1118 0.0169185
R28098 DVDD.n4390 DVDD.n1584 0.0169185
R28099 DVDD.n3776 DVDD.n1866 0.0169185
R28100 DVDD.n3744 DVDD.n1865 0.0169185
R28101 DVDD.n3743 DVDD.n1864 0.0169185
R28102 DVDD.n3742 DVDD.n1863 0.0169185
R28103 DVDD.n3741 DVDD.n1862 0.0169185
R28104 DVDD.n3740 DVDD.n1860 0.0169185
R28105 DVDD.n3739 DVDD.n1859 0.0169185
R28106 DVDD.n3738 DVDD.n1858 0.0169185
R28107 DVDD.n3737 DVDD.n1857 0.0169185
R28108 DVDD.n1990 DVDD.n1981 0.0169185
R28109 DVDD.n1989 DVDD.n1987 0.0169185
R28110 DVDD.n3670 DVDD.n1992 0.0169185
R28111 DVDD.n1991 DVDD.n1986 0.0169185
R28112 DVDD.n3669 DVDD.n1994 0.0169185
R28113 DVDD.n1993 DVDD.n1985 0.0169185
R28114 DVDD.n3668 DVDD.n1996 0.0169185
R28115 DVDD.n1995 DVDD.n1984 0.0169185
R28116 DVDD.n3673 DVDD.n3672 0.0169185
R28117 DVDD.n2405 DVDD.n1998 0.0169185
R28118 DVDD.n2042 DVDD.n2003 0.0169185
R28119 DVDD.n2005 DVDD.n2003 0.0169185
R28120 DVDD.n2041 DVDD.n2002 0.0169185
R28121 DVDD.n2007 DVDD.n2002 0.0169185
R28122 DVDD.n2040 DVDD.n2001 0.0169185
R28123 DVDD.n2009 DVDD.n2001 0.0169185
R28124 DVDD.n2402 DVDD.n2000 0.0169185
R28125 DVDD.n2011 DVDD.n2000 0.0169185
R28126 DVDD.n3778 DVDD.n3722 0.0169185
R28127 DVDD.n3753 DVDD.n3737 0.0169185
R28128 DVDD.n3752 DVDD.n3738 0.0169185
R28129 DVDD.n3751 DVDD.n3739 0.0169185
R28130 DVDD.n3750 DVDD.n3740 0.0169185
R28131 DVDD.n3749 DVDD.n1887 0.0169185
R28132 DVDD.n3748 DVDD.n3741 0.0169185
R28133 DVDD.n3747 DVDD.n3742 0.0169185
R28134 DVDD.n3746 DVDD.n3743 0.0169185
R28135 DVDD.n3745 DVDD.n3744 0.0169185
R28136 DVDD.n4390 DVDD.n1118 0.0169185
R28137 DVDD.n4410 DVDD.n1585 0.0169185
R28138 DVDD.n4391 DVDD.n1117 0.0169185
R28139 DVDD.n4409 DVDD.n1586 0.0169185
R28140 DVDD.n4392 DVDD.n1116 0.0169185
R28141 DVDD.n4408 DVDD.n1587 0.0169185
R28142 DVDD.n4393 DVDD.n1115 0.0169185
R28143 DVDD.n4407 DVDD.n1588 0.0169185
R28144 DVDD.n4394 DVDD.n1114 0.0169185
R28145 DVDD.n4406 DVDD.n1589 0.0169185
R28146 DVDD.n4395 DVDD.n1113 0.0169185
R28147 DVDD.n4405 DVDD.n1590 0.0169185
R28148 DVDD.n4396 DVDD.n1112 0.0169185
R28149 DVDD.n4404 DVDD.n1591 0.0169185
R28150 DVDD.n4397 DVDD.n1111 0.0169185
R28151 DVDD.n4403 DVDD.n1592 0.0169185
R28152 DVDD.n4398 DVDD.n1110 0.0169185
R28153 DVDD.n4402 DVDD.n1593 0.0169185
R28154 DVDD.n4399 DVDD.n1109 0.0169185
R28155 DVDD.n4415 DVDD.n4414 0.0169185
R28156 DVDD.n1606 DVDD.n1594 0.0169185
R28157 DVDD.n1609 DVDD.n1608 0.0169185
R28158 DVDD.n4376 DVDD.n1605 0.0169185
R28159 DVDD.n1611 DVDD.n1610 0.0169185
R28160 DVDD.n4377 DVDD.n1604 0.0169185
R28161 DVDD.n1613 DVDD.n1612 0.0169185
R28162 DVDD.n4378 DVDD.n1603 0.0169185
R28163 DVDD.n1615 DVDD.n1614 0.0169185
R28164 DVDD.n4379 DVDD.n1602 0.0169185
R28165 DVDD.n1617 DVDD.n1616 0.0169185
R28166 DVDD.n4380 DVDD.n1601 0.0169185
R28167 DVDD.n1619 DVDD.n1618 0.0169185
R28168 DVDD.n4381 DVDD.n1600 0.0169185
R28169 DVDD.n1621 DVDD.n1620 0.0169185
R28170 DVDD.n4382 DVDD.n1599 0.0169185
R28171 DVDD.n1623 DVDD.n1622 0.0169185
R28172 DVDD.n4383 DVDD.n1598 0.0169185
R28173 DVDD.n1625 DVDD.n1624 0.0169185
R28174 DVDD.n4384 DVDD.n1597 0.0169185
R28175 DVDD.n4387 DVDD.n4386 0.0169185
R28176 DVDD.n1638 DVDD.n1626 0.0169185
R28177 DVDD.n1641 DVDD.n1640 0.0169185
R28178 DVDD.n4333 DVDD.n1637 0.0169185
R28179 DVDD.n1643 DVDD.n1642 0.0169185
R28180 DVDD.n4334 DVDD.n1636 0.0169185
R28181 DVDD.n1645 DVDD.n1644 0.0169185
R28182 DVDD.n4335 DVDD.n1635 0.0169185
R28183 DVDD.n1647 DVDD.n1646 0.0169185
R28184 DVDD.n4336 DVDD.n1634 0.0169185
R28185 DVDD.n1649 DVDD.n1648 0.0169185
R28186 DVDD.n4337 DVDD.n1633 0.0169185
R28187 DVDD.n1651 DVDD.n1650 0.0169185
R28188 DVDD.n4338 DVDD.n1632 0.0169185
R28189 DVDD.n1653 DVDD.n1652 0.0169185
R28190 DVDD.n4339 DVDD.n1631 0.0169185
R28191 DVDD.n1655 DVDD.n1654 0.0169185
R28192 DVDD.n4340 DVDD.n1630 0.0169185
R28193 DVDD.n1657 DVDD.n1656 0.0169185
R28194 DVDD.n4341 DVDD.n1629 0.0169185
R28195 DVDD.n4344 DVDD.n4343 0.0169185
R28196 DVDD.n5777 DVDD.n179 0.0167295
R28197 DVDD.n5787 DVDD.n5786 0.0167295
R28198 DVDD.n5847 DVDD.n138 0.0167295
R28199 DVDD.n5204 DVDD.n494 0.0167295
R28200 DVDD.n5198 DVDD.n495 0.0167295
R28201 DVDD.n5141 DVDD.n5140 0.0167295
R28202 DVDD.n664 DVDD.n615 0.0167295
R28203 DVDD.n626 DVDD.n606 0.0167295
R28204 DVDD.n4994 DVDD.n427 0.0167295
R28205 DVDD.n828 DVDD.n713 0.0167295
R28206 DVDD.n822 DVDD.n714 0.0167295
R28207 DVDD.n758 DVDD.n403 0.0167295
R28208 DVDD.n4577 DVDD.n1018 0.0167295
R28209 DVDD.n4571 DVDD.n1019 0.0167295
R28210 DVDD.n4550 DVDD.n380 0.0167295
R28211 DVDD.n2660 DVDD.n2493 0.0167
R28212 DVDD.n3190 DVDD.n3189 0.0166964
R28213 DVDD.n5568 DVDD.n5567 0.0166102
R28214 DVDD.n275 DVDD.n274 0.0166102
R28215 DVDD.n3255 DVDD.n2986 0.016475
R28216 DVDD.n5644 DVDD.n66 0.0164553
R28217 DVDD.n5469 DVDD.n299 0.0164553
R28218 DVDD.n2843 DVDD.n2795 0.0163967
R28219 DVDD.n2893 DVDD.n2876 0.0163967
R28220 DVDD.n5837 DVDD.n142 0.0163607
R28221 DVDD.n5319 DVDD.n473 0.0163607
R28222 DVDD.n5005 DVDD.n4951 0.0163607
R28223 DVDD.n770 DVDD.n769 0.0163607
R28224 DVDD.n4561 DVDD.n4509 0.0163607
R28225 DVDD.n5521 DVDD.n9 0.0163003
R28226 DVDD.n4695 DVDD.n976 0.0163003
R28227 DVDD.n2660 DVDD.n2497 0.01625
R28228 DVDD.n2637 DVDD.n2450 0.0161522
R28229 DVDD.n5627 DVDD.n54 0.0161454
R28230 DVDD.n5452 DVDD.n312 0.0161454
R28231 DVDD.n5766 DVDD.n177 0.0159918
R28232 DVDD.n5220 DVDD.n561 0.0159918
R28233 DVDD.n648 DVDD.n613 0.0159918
R28234 DVDD.n844 DVDD.n721 0.0159918
R28235 DVDD.n4593 DVDD.n1052 0.0159918
R28236 DVDD.n5537 DVDD.n23 0.0159905
R28237 DVDD.n4679 DVDD.n4652 0.0159905
R28238 DVDD.n71 DVDD.n59 0.0158356
R28239 DVDD.n5436 DVDD.n306 0.0158356
R28240 DVDD.n5554 DVDD.n16 0.0156807
R28241 DVDD.n5560 DVDD.n8 0.0156807
R28242 DVDD.n4662 DVDD.n983 0.0156807
R28243 DVDD.n4646 DVDD.n267 0.0156807
R28244 DVDD.n3273 DVDD.n2932 0.015663
R28245 DVDD.n2948 DVDD.n2940 0.015663
R28246 DVDD.n2653 DVDD.n2651 0.0156593
R28247 DVDD.n5809 DVDD.n151 0.015623
R28248 DVDD.n5165 DVDD.n465 0.015623
R28249 DVDD.n4976 DVDD.n4943 0.015623
R28250 DVDD.n787 DVDD.n786 0.015623
R28251 DVDD.n4532 DVDD.n4502 0.015623
R28252 DVDD.n939 DVDD.n928 0.0155811
R28253 DVDD.n939 DVDD.n938 0.0155811
R28254 DVDD.n938 DVDD.n935 0.0155811
R28255 DVDD.n935 DVDD.n934 0.0155811
R28256 DVDD.n934 DVDD.n932 0.0155811
R28257 DVDD.n932 DVDD.n930 0.0155811
R28258 DVDD.n953 DVDD.n951 0.0155811
R28259 DVDD.n954 DVDD.n953 0.0155811
R28260 DVDD.n957 DVDD.n954 0.0155811
R28261 DVDD.n959 DVDD.n957 0.0155811
R28262 DVDD.n960 DVDD.n959 0.0155811
R28263 DVDD.n1923 DVDD.n1896 0.015575
R28264 DVDD.n3079 DVDD.n2750 0.015575
R28265 DVDD.n3691 DVDD.n1916 0.015575
R28266 DVDD.n3255 DVDD.n3080 0.015575
R28267 DVDD.n258 DVDD.n243 0.0154398
R28268 DVDD.n5673 DVDD.n243 0.0154398
R28269 DVDD.n5673 DVDD.n5672 0.0154398
R28270 DVDD.n5672 DVDD.n5671 0.0154398
R28271 DVDD.n5671 DVDD.n5669 0.0154398
R28272 DVDD.n5669 DVDD.n5667 0.0154398
R28273 DVDD.n255 DVDD.n253 0.0154398
R28274 DVDD.n253 DVDD.n251 0.0154398
R28275 DVDD.n251 DVDD.n248 0.0154398
R28276 DVDD.n248 DVDD.n247 0.0154398
R28277 DVDD.n247 DVDD.n245 0.0154398
R28278 DVDD.n5544 DVDD.n21 0.0153709
R28279 DVDD.n4672 DVDD.n4650 0.0153709
R28280 DVDD.n3527 DVDD.n2669 0.01535
R28281 DVDD.n104 DVDD.n98 0.0153356
R28282 DVDD.n5918 DVDD.n101 0.0153356
R28283 DVDD.n5421 DVDD.n337 0.0153356
R28284 DVDD.n5423 DVDD.n348 0.0153356
R28285 DVDD.n5421 DVDD.n344 0.0153356
R28286 DVDD.n104 DVDD.n90 0.0153356
R28287 DVDD.n101 DVDD.n88 0.0153356
R28288 DVDD.n348 DVDD.n334 0.0153356
R28289 DVDD.n3680 DVDD.n1976 0.0153088
R28290 DVDD.n3688 DVDD.n1976 0.0153088
R28291 DVDD.n3689 DVDD.n3688 0.0153088
R28292 DVDD.n3709 DVDD.n1892 0.0153088
R28293 DVDD.n3717 DVDD.n1892 0.0153088
R28294 DVDD.n3717 DVDD.n1890 0.0153088
R28295 DVDD.n3771 DVDD.n3757 0.0153088
R28296 DVDD.n3771 DVDD.n3759 0.0153088
R28297 DVDD.n3764 DVDD.n3759 0.0153088
R28298 DVDD.n4289 DVDD.n1662 0.0153088
R28299 DVDD.n4297 DVDD.n1662 0.0153088
R28300 DVDD.n4297 DVDD.n1660 0.0153088
R28301 DVDD.n5750 DVDD.n175 0.0152541
R28302 DVDD.n5236 DVDD.n487 0.0152541
R28303 DVDD.n632 DVDD.n611 0.0152541
R28304 DVDD.n860 DVDD.n706 0.0152541
R28305 DVDD.n4609 DVDD.n1011 0.0152541
R28306 DVDD.n5527 DVDD.n11 0.0150611
R28307 DVDD.n4689 DVDD.n978 0.0150611
R28308 DVDD.n1122 DVDD.n1119 0.015031
R28309 DVDD.n1581 DVDD.n1149 0.015031
R28310 DVDD.n1580 DVDD.n1123 0.015031
R28311 DVDD.n1148 DVDD.n1147 0.015031
R28312 DVDD.n1182 DVDD.n1124 0.015031
R28313 DVDD.n1146 DVDD.n1145 0.015031
R28314 DVDD.n1183 DVDD.n1125 0.015031
R28315 DVDD.n1144 DVDD.n1143 0.015031
R28316 DVDD.n1184 DVDD.n1126 0.015031
R28317 DVDD.n1142 DVDD.n1141 0.015031
R28318 DVDD.n1185 DVDD.n1127 0.015031
R28319 DVDD.n1140 DVDD.n1139 0.015031
R28320 DVDD.n1186 DVDD.n1128 0.015031
R28321 DVDD.n1138 DVDD.n1137 0.015031
R28322 DVDD.n1187 DVDD.n1129 0.015031
R28323 DVDD.n1136 DVDD.n1135 0.015031
R28324 DVDD.n1188 DVDD.n1130 0.015031
R28325 DVDD.n1134 DVDD.n1133 0.015031
R28326 DVDD.n1190 DVDD.n1189 0.015031
R28327 DVDD.n1578 DVDD.n1132 0.015031
R28328 DVDD.n1189 DVDD.n1132 0.015031
R28329 DVDD.n1190 DVDD.n1134 0.015031
R28330 DVDD.n1133 DVDD.n1130 0.015031
R28331 DVDD.n1188 DVDD.n1136 0.015031
R28332 DVDD.n1135 DVDD.n1129 0.015031
R28333 DVDD.n1187 DVDD.n1138 0.015031
R28334 DVDD.n1137 DVDD.n1128 0.015031
R28335 DVDD.n1186 DVDD.n1140 0.015031
R28336 DVDD.n1139 DVDD.n1127 0.015031
R28337 DVDD.n1185 DVDD.n1142 0.015031
R28338 DVDD.n1141 DVDD.n1126 0.015031
R28339 DVDD.n1184 DVDD.n1144 0.015031
R28340 DVDD.n1143 DVDD.n1125 0.015031
R28341 DVDD.n1183 DVDD.n1146 0.015031
R28342 DVDD.n1145 DVDD.n1124 0.015031
R28343 DVDD.n1182 DVDD.n1148 0.015031
R28344 DVDD.n1147 DVDD.n1123 0.015031
R28345 DVDD.n1581 DVDD.n1580 0.015031
R28346 DVDD.n1149 DVDD.n1122 0.015031
R28347 DVDD.n1583 DVDD.n1119 0.015031
R28348 DVDD.n1382 DVDD.n1307 0.0149495
R28349 DVDD.n1390 DVDD.n1311 0.0149495
R28350 DVDD.n1318 DVDD.n1219 0.0149495
R28351 DVDD.n1314 DVDD.n1221 0.0149495
R28352 DVDD.n2835 DVDD.n2785 0.0149293
R28353 DVDD.n2901 DVDD.n2865 0.0149293
R28354 DVDD.n2606 DVDD.n2509 0.0149069
R28355 DVDD.n2609 DVDD.n2506 0.0149069
R28356 DVDD.n2509 DVDD.n2506 0.0149069
R28357 DVDD.n2607 DVDD.n2606 0.0149069
R28358 DVDD.n5504 DVDD.n221 0.0149062
R28359 DVDD.n964 DVDD.n947 0.0149062
R28360 DVDD.n2652 DVDD.n2491 0.0149
R28361 DVDD.n5740 DVDD.n193 0.0148852
R28362 DVDD.n5825 DVDD.n162 0.0148852
R28363 DVDD.n5098 DVDD.n5097 0.0148852
R28364 DVDD.n5181 DVDD.n467 0.0148852
R28365 DVDD.n5021 DVDD.n5020 0.0148852
R28366 DVDD.n4960 DVDD.n4945 0.0148852
R28367 DVDD.n870 DVDD.n737 0.0148852
R28368 DVDD.n805 DVDD.n804 0.0148852
R28369 DVDD.n1066 DVDD.n894 0.0148852
R28370 DVDD.n4516 DVDD.n4504 0.0148852
R28371 DVDD.n2629 DVDD.n2447 0.0146848
R28372 DVDD.n5621 DVDD.n5605 0.0144415
R28373 DVDD.n5446 DVDD.n287 0.0144415
R28374 DVDD.n2198 DVDD.n2197 0.0142814
R28375 DVDD.n3471 DVDD.n3470 0.0142814
R28376 DVDD.n1363 DVDD.n1362 0.0141845
R28377 DVDD.n2956 DVDD.n2954 0.0141679
R28378 DVDD.n2936 DVDD.n2934 0.0141679
R28379 DVDD.n2952 DVDD.n2933 0.0141679
R28380 DVDD.n3275 DVDD.n2955 0.0141679
R28381 DVDD.n2937 DVDD.n2933 0.0141679
R28382 DVDD.n2951 DVDD.n2936 0.0141679
R28383 DVDD.n3276 DVDD.n3275 0.0141679
R28384 DVDD.n2957 DVDD.n2954 0.0141679
R28385 DVDD.n2648 DVDD.n2645 0.0141679
R28386 DVDD.n2645 DVDD.n2627 0.0141679
R28387 DVDD.n2650 DVDD.n2627 0.0141679
R28388 DVDD.n2648 DVDD.n2647 0.0141679
R28389 DVDD.n5638 DVDD.n5571 0.0141317
R28390 DVDD.n5463 DVDD.n278 0.0141317
R28391 DVDD.n1374 DVDD.n1328 0.0140776
R28392 DVDD.n1328 DVDD.n1327 0.0140776
R28393 DVDD.n2817 DVDD.n2790 0.013978
R28394 DVDD.n3333 DVDD.n2873 0.013978
R28395 DVDD.n2825 DVDD.n2792 0.0139511
R28396 DVDD.n2911 DVDD.n2879 0.0139511
R28397 DVDD.n5653 DVDD.n5652 0.0138219
R28398 DVDD.n5479 DVDD.n5478 0.0138219
R28399 DVDD.n2508 DVDD.n2505 0.0137065
R28400 DVDD.n5642 DVDD.n51 0.013667
R28401 DVDD.n5509 DVDD.n218 0.013667
R28402 DVDD.n4707 DVDD.n948 0.013667
R28403 DVDD.n5467 DVDD.n315 0.013667
R28404 DVDD DVDD.n2540 0.0135263
R28405 DVDD.n5523 DVDD.n26 0.013512
R28406 DVDD.n4693 DVDD.n4655 0.013512
R28407 DVDD.n3065 DVDD.n3061 0.0135078
R28408 DVDD.n2827 DVDD.n2792 0.013462
R28409 DVDD.n2909 DVDD.n2879 0.013462
R28410 DVDD.n3173 DVDD.n3154 0.0134255
R28411 DVDD.n3173 DVDD.n3155 0.0134255
R28412 DVDD.n3229 DVDD.n3095 0.0134255
R28413 DVDD.n3114 DVDD.n3095 0.0134255
R28414 DVDD.n963 DVDD.n961 0.0134017
R28415 DVDD.n965 DVDD.n963 0.0134017
R28416 DVDD.n969 DVDD.n968 0.0134017
R28417 DVDD.n4705 DVDD.n969 0.0134017
R28418 DVDD.n4705 DVDD.n4704 0.0134017
R28419 DVDD.n4704 DVDD.n4703 0.0134017
R28420 DVDD.n4703 DVDD.n970 0.0134017
R28421 DVDD.n4657 DVDD.n970 0.0134017
R28422 DVDD.n4697 DVDD.n4657 0.0134017
R28423 DVDD.n4697 DVDD.n4696 0.0134017
R28424 DVDD.n4696 DVDD.n4694 0.0134017
R28425 DVDD.n4694 DVDD.n4692 0.0134017
R28426 DVDD.n4692 DVDD.n4690 0.0134017
R28427 DVDD.n4690 DVDD.n4688 0.0134017
R28428 DVDD.n4688 DVDD.n4686 0.0134017
R28429 DVDD.n4686 DVDD.n4683 0.0134017
R28430 DVDD.n4683 DVDD.n4682 0.0134017
R28431 DVDD.n4682 DVDD.n4680 0.0134017
R28432 DVDD.n4677 DVDD.n4675 0.0134017
R28433 DVDD.n4675 DVDD.n4673 0.0134017
R28434 DVDD.n4673 DVDD.n4671 0.0134017
R28435 DVDD.n4671 DVDD.n4669 0.0134017
R28436 DVDD.n4669 DVDD.n4666 0.0134017
R28437 DVDD.n4666 DVDD.n4665 0.0134017
R28438 DVDD.n4665 DVDD.n4663 0.0134017
R28439 DVDD.n4663 DVDD.n4661 0.0134017
R28440 DVDD.n4661 DVDD.n4659 0.0134017
R28441 DVDD.n4659 DVDD.n265 0.0134017
R28442 DVDD.n5481 DVDD.n266 0.0134017
R28443 DVDD.n5481 DVDD.n5480 0.0134017
R28444 DVDD.n5480 DVDD.n269 0.0134017
R28445 DVDD.n318 DVDD.n269 0.0134017
R28446 DVDD.n319 DVDD.n318 0.0134017
R28447 DVDD.n5471 DVDD.n319 0.0134017
R28448 DVDD.n5471 DVDD.n5470 0.0134017
R28449 DVDD.n5470 DVDD.n5468 0.0134017
R28450 DVDD.n5468 DVDD.n5466 0.0134017
R28451 DVDD.n5466 DVDD.n5464 0.0134017
R28452 DVDD.n5464 DVDD.n5462 0.0134017
R28453 DVDD.n5462 DVDD.n5460 0.0134017
R28454 DVDD.n5456 DVDD.n5455 0.0134017
R28455 DVDD.n5455 DVDD.n5453 0.0134017
R28456 DVDD.n5453 DVDD.n5451 0.0134017
R28457 DVDD.n5451 DVDD.n5449 0.0134017
R28458 DVDD.n5449 DVDD.n5447 0.0134017
R28459 DVDD.n5447 DVDD.n5445 0.0134017
R28460 DVDD.n5445 DVDD.n5443 0.0134017
R28461 DVDD.n5443 DVDD.n5440 0.0134017
R28462 DVDD.n5440 DVDD.n5439 0.0134017
R28463 DVDD.n5439 DVDD.n5437 0.0134017
R28464 DVDD.n5437 DVDD.n5435 0.0134017
R28465 DVDD.n5435 DVDD.n5434 0.0134017
R28466 DVDD.n5434 DVDD.n5433 0.0134017
R28467 DVDD.n5433 DVDD.n320 0.0134017
R28468 DVDD.n330 DVDD.n320 0.0134017
R28469 DVDD.n332 DVDD.n330 0.0134017
R28470 DVDD.n5426 DVDD.n5425 0.0134017
R28471 DVDD.n5485 DVDD.n266 0.0134017
R28472 DVDD.n5659 DVDD.n5562 0.013372
R28473 DVDD.n5503 DVDD.n223 0.013372
R28474 DVDD.n5505 DVDD.n5503 0.013372
R28475 DVDD.n5510 DVDD.n5508 0.013372
R28476 DVDD.n5511 DVDD.n5510 0.013372
R28477 DVDD.n5514 DVDD.n5511 0.013372
R28478 DVDD.n5515 DVDD.n5514 0.013372
R28479 DVDD.n5516 DVDD.n5515 0.013372
R28480 DVDD.n5518 DVDD.n5516 0.013372
R28481 DVDD.n5520 DVDD.n5518 0.013372
R28482 DVDD.n5522 DVDD.n5520 0.013372
R28483 DVDD.n5524 DVDD.n5522 0.013372
R28484 DVDD.n5526 DVDD.n5524 0.013372
R28485 DVDD.n5528 DVDD.n5526 0.013372
R28486 DVDD.n5530 DVDD.n5528 0.013372
R28487 DVDD.n5531 DVDD.n5530 0.013372
R28488 DVDD.n5534 DVDD.n5531 0.013372
R28489 DVDD.n5536 DVDD.n5534 0.013372
R28490 DVDD.n5538 DVDD.n5536 0.013372
R28491 DVDD.n5543 DVDD.n5541 0.013372
R28492 DVDD.n5545 DVDD.n5543 0.013372
R28493 DVDD.n5547 DVDD.n5545 0.013372
R28494 DVDD.n5548 DVDD.n5547 0.013372
R28495 DVDD.n5551 DVDD.n5548 0.013372
R28496 DVDD.n5553 DVDD.n5551 0.013372
R28497 DVDD.n5555 DVDD.n5553 0.013372
R28498 DVDD.n5557 DVDD.n5555 0.013372
R28499 DVDD.n5559 DVDD.n5557 0.013372
R28500 DVDD.n5561 DVDD.n5559 0.013372
R28501 DVDD.n5655 DVDD.n5562 0.013372
R28502 DVDD.n5655 DVDD.n5654 0.013372
R28503 DVDD.n5654 DVDD.n5564 0.013372
R28504 DVDD.n5612 DVDD.n5564 0.013372
R28505 DVDD.n5648 DVDD.n5612 0.013372
R28506 DVDD.n5648 DVDD.n5647 0.013372
R28507 DVDD.n5647 DVDD.n5645 0.013372
R28508 DVDD.n5645 DVDD.n5643 0.013372
R28509 DVDD.n5643 DVDD.n5641 0.013372
R28510 DVDD.n5641 DVDD.n5639 0.013372
R28511 DVDD.n5639 DVDD.n5637 0.013372
R28512 DVDD.n5637 DVDD.n5635 0.013372
R28513 DVDD.n5631 DVDD.n5630 0.013372
R28514 DVDD.n5630 DVDD.n5628 0.013372
R28515 DVDD.n5628 DVDD.n5626 0.013372
R28516 DVDD.n5626 DVDD.n5624 0.013372
R28517 DVDD.n5624 DVDD.n5622 0.013372
R28518 DVDD.n5622 DVDD.n5620 0.013372
R28519 DVDD.n5620 DVDD.n5618 0.013372
R28520 DVDD.n5618 DVDD.n5615 0.013372
R28521 DVDD.n5615 DVDD.n5614 0.013372
R28522 DVDD.n5614 DVDD.n72 0.013372
R28523 DVDD.n5931 DVDD.n72 0.013372
R28524 DVDD.n5931 DVDD.n5930 0.013372
R28525 DVDD.n5930 DVDD.n73 0.013372
R28526 DVDD.n5926 DVDD.n73 0.013372
R28527 DVDD.n5926 DVDD.n5925 0.013372
R28528 DVDD.n5925 DVDD.n75 0.013372
R28529 DVDD.n5920 DVDD.n86 0.013372
R28530 DVDD.n5625 DVDD.n62 0.0133571
R28531 DVDD.n5450 DVDD.n303 0.0133571
R28532 DVDD.n3677 DVDD.n1980 0.0133273
R28533 DVDD.n3682 DVDD.n3681 0.0133273
R28534 DVDD.n3686 DVDD.n1978 0.0133273
R28535 DVDD.n3687 DVDD.n1975 0.0133273
R28536 DVDD.n3711 DVDD.n3710 0.0133273
R28537 DVDD.n3714 DVDD.n1893 0.0133273
R28538 DVDD.n3716 DVDD.n3715 0.0133273
R28539 DVDD.n3720 DVDD.n1889 0.0133273
R28540 DVDD.n1371 DVDD.n1200 0.0132218
R28541 DVDD.n5540 DVDD.n13 0.0132022
R28542 DVDD.n4676 DVDD.n980 0.0132022
R28543 DVDD.n5933 DVDD.n5932 0.0130473
R28544 DVDD.n308 DVDD.n294 0.0130473
R28545 DVDD.n5924 DVDD.n5923 0.0128924
R28546 DVDD.n5556 DVDD.n19 0.0128924
R28547 DVDD.n5558 DVDD.n18 0.0128924
R28548 DVDD.n4660 DVDD.n4648 0.0128924
R28549 DVDD.n4658 DVDD.n4647 0.0128924
R28550 DVDD.n326 DVDD.n323 0.0128924
R28551 DVDD.n5911 DVDD.n97 0.0127938
R28552 DVDD.n113 DVDD.n96 0.0127938
R28553 DVDD.n5414 DVDD.n336 0.0127938
R28554 DVDD.n5411 DVDD.n335 0.0127938
R28555 DVDD.n931 DVDD.n925 0.0127938
R28556 DVDD.n950 DVDD.n918 0.0127938
R28557 DVDD.n5668 DVDD.n231 0.0127938
R28558 DVDD.n254 DVDD.n237 0.0127938
R28559 DVDD.n2454 DVDD.n2447 0.0127283
R28560 DVDD.n5835 DVDD.n5834 0.0126721
R28561 DVDD.n5189 DVDD.n469 0.0126721
R28562 DVDD.n4952 DVDD.n4947 0.0126721
R28563 DVDD.n814 DVDD.n813 0.0126721
R28564 DVDD.n4563 DVDD.n1074 0.0126721
R28565 DVDD.n3045 DVDD.n3044 0.0126289
R28566 DVDD.n5542 DVDD.n14 0.0125826
R28567 DVDD.n4674 DVDD.n981 0.0125826
R28568 DVDD.n1370 DVDD.n1369 0.0125
R28569 DVDD.n2833 DVDD.n2785 0.0124837
R28570 DVDD.n2903 DVDD.n2865 0.0124837
R28571 DVDD.n1887 DVDD.n1886 0.012425
R28572 DVDD.n5525 DVDD.n25 0.0122728
R28573 DVDD.n4691 DVDD.n4654 0.0122728
R28574 DVDD.n5460 DVDD.n5457 0.0121532
R28575 DVDD.n5635 DVDD.n5632 0.0121263
R28576 DVDD.n5507 DVDD.n219 0.0121179
R28577 DVDD.n967 DVDD.n945 0.0121179
R28578 DVDD.n5817 DVDD.n149 0.0119344
R28579 DVDD.n5173 DVDD.n454 0.0119344
R28580 DVDD.n4968 DVDD.n677 0.0119344
R28581 DVDD.n797 DVDD.n796 0.0119344
R28582 DVDD.n4524 DVDD.n1078 0.0119344
R28583 DVDD.n3774 DVDD.n3756 0.011763
R28584 DVDD.n3761 DVDD.n3760 0.011763
R28585 DVDD.n3770 DVDD.n3769 0.011763
R28586 DVDD.n3766 DVDD.n3762 0.011763
R28587 DVDD.n4291 DVDD.n4290 0.011763
R28588 DVDD.n4294 DVDD.n1663 0.011763
R28589 DVDD.n4296 DVDD.n4295 0.011763
R28590 DVDD.n4300 DVDD.n1659 0.011763
R28591 DVDD.n1205 DVDD.n1193 0.0117585
R28592 DVDD.n3274 DVDD.n3273 0.01175
R28593 DVDD.n2949 DVDD.n2948 0.01175
R28594 DVDD.n3389 DVDD.n2738 0.01175
R28595 DVDD.n5623 DVDD.n5574 0.0116532
R28596 DVDD.n5448 DVDD.n281 0.0116532
R28597 DVDD.n5486 DVDD.n265 0.0116329
R28598 DVDD.n5660 DVDD.n5561 0.0116073
R28599 DVDD.n5758 DVDD.n188 0.0115656
R28600 DVDD.n5228 DVDD.n563 0.0115656
R28601 DVDD.n640 DVDD.n623 0.0115656
R28602 DVDD.n852 DVDD.n723 0.0115656
R28603 DVDD.n4601 DVDD.n1054 0.0115656
R28604 DVDD.n5640 DVDD.n5609 0.0113434
R28605 DVDD.n5465 DVDD.n291 0.0113434
R28606 DVDD.n2635 DVDD.n2450 0.0112609
R28607 DVDD.n5801 DVDD.n157 0.0111967
R28608 DVDD.n5157 DVDD.n472 0.0111967
R28609 DVDD.n4984 DVDD.n4950 0.0111967
R28610 DVDD.n779 DVDD.n778 0.0111967
R28611 DVDD.n4540 DVDD.n4508 0.0111967
R28612 DVDD.n5656 DVDD.n5563 0.0110336
R28613 DVDD.n5482 DVDD.n268 0.0110336
R28614 DVDD.n2841 DVDD.n2795 0.0110163
R28615 DVDD.n2895 DVDD.n2876 0.0110163
R28616 DVDD.n5640 DVDD.n65 0.0108787
R28617 DVDD.n5507 DVDD.n222 0.0108787
R28618 DVDD.n967 DVDD.n946 0.0108787
R28619 DVDD.n5465 DVDD.n300 0.0108787
R28620 DVDD.n190 DVDD.n171 0.0108279
R28621 DVDD.n5212 DVDD.n492 0.0108279
R28622 DVDD.n656 DVDD.n607 0.0108279
R28623 DVDD.n836 DVDD.n711 0.0108279
R28624 DVDD.n4585 DVDD.n1016 0.0108279
R28625 DVDD.n5525 DVDD.n10 0.0107238
R28626 DVDD.n4691 DVDD.n977 0.0107238
R28627 DVDD.n1577 DVDD.n1191 0.0105885
R28628 DVDD.n1203 DVDD.n1196 0.0105885
R28629 DVDD.n1204 DVDD.n1195 0.0105885
R28630 DVDD.n1575 DVDD.n1574 0.0105885
R28631 DVDD.n1574 DVDD.n1194 0.0105885
R28632 DVDD.n1204 DVDD.n1202 0.0105885
R28633 DVDD.n1203 DVDD.n1200 0.0105885
R28634 DVDD.n1199 DVDD.n1191 0.0105885
R28635 DVDD.n1198 DVDD.n1196 0.0105885
R28636 DVDD.n1201 DVDD.n1194 0.0105885
R28637 DVDD.n1202 DVDD.n1201 0.0105885
R28638 DVDD.n1199 DVDD.n1198 0.0105885
R28639 DVDD.n5623 DVDD.n55 0.0105688
R28640 DVDD.n5448 DVDD.n311 0.0105688
R28641 DVDD.n3707 DVDD.n1901 0.01055
R28642 DVDD.n5542 DVDD.n22 0.0104139
R28643 DVDD.n4674 DVDD.n4651 0.0104139
R28644 DVDD.n3404 DVDD.n2726 0.0104
R28645 DVDD.n3268 DVDD.n2959 0.0104
R28646 DVDD.n3381 DVDD.n3380 0.0104
R28647 DVDD.n3070 DVDD.n3069 0.0104
R28648 DVDD.n3678 DVDD.n1977 0.0103725
R28649 DVDD.n1977 DVDD.n1910 0.0103725
R28650 DVDD.n3708 DVDD.n1891 0.0103725
R28651 DVDD.n3718 DVDD.n1891 0.0103725
R28652 DVDD.n3772 DVDD.n3758 0.0103725
R28653 DVDD.n3758 DVDD.n1667 0.0103725
R28654 DVDD.n4288 DVDD.n1661 0.0103725
R28655 DVDD.n4298 DVDD.n1661 0.0103725
R28656 DVDD.n3295 DVDD.n3292 0.0102826
R28657 DVDD.n3329 DVDD.n2915 0.0102826
R28658 DVDD.n3370 DVDD.n2764 0.0102826
R28659 DVDD.n2813 DVDD.n2802 0.0102826
R28660 DVDD.n5929 DVDD.n48 0.010259
R28661 DVDD.n5475 DVDD.n296 0.010259
R28662 DVDD.n3234 DVDD.n3096 0.0102297
R28663 DVDD.n3164 DVDD.n3163 0.0102297
R28664 DVDD.n5927 DVDD.n74 0.0101041
R28665 DVDD.n5924 DVDD.n74 0.0101041
R28666 DVDD.n5556 DVDD.n17 0.0101041
R28667 DVDD.n5558 DVDD.n17 0.0101041
R28668 DVDD.n4660 DVDD.n984 0.0101041
R28669 DVDD.n4658 DVDD.n984 0.0101041
R28670 DVDD.n5431 DVDD.n5430 0.0101041
R28671 DVDD.n5430 DVDD.n323 0.0101041
R28672 DVDD.n5779 DVDD.n182 0.0100902
R28673 DVDD.n5790 DVDD.n166 0.0100902
R28674 DVDD.n5206 DVDD.n558 0.0100902
R28675 DVDD.n5196 DVDD.n556 0.0100902
R28676 DVDD.n662 DVDD.n618 0.0100902
R28677 DVDD.n5013 DVDD.n5012 0.0100902
R28678 DVDD.n830 DVDD.n718 0.0100902
R28679 DVDD.n820 DVDD.n716 0.0100902
R28680 DVDD.n4579 DVDD.n1049 0.0100902
R28681 DVDD.n4569 DVDD.n1047 0.0100902
R28682 DVDD.n3527 DVDD.n2499 0.00995
R28683 DVDD.n84 DVDD.n81 0.00994923
R28684 DVDD.n5428 DVDD.n329 0.00994923
R28685 DVDD.n3436 DVDD.n3435 0.00992
R28686 DVDD.n3437 DVDD.n2695 0.00992
R28687 DVDD.n3321 DVDD.n3319 0.00992
R28688 DVDD.n3358 DVDD.n3357 0.00992
R28689 DVDD.n3037 DVDD.n3036 0.00992
R28690 DVDD.n3035 DVDD.n3020 0.00992
R28691 DVDD.n5540 DVDD.n22 0.00979432
R28692 DVDD.n4676 DVDD.n4651 0.00979432
R28693 DVDD.n2643 DVDD.n2444 0.00979348
R28694 DVDD.n5795 DVDD.n154 0.00972131
R28695 DVDD.n5151 DVDD.n461 0.00972131
R28696 DVDD.n4990 DVDD.n683 0.00972131
R28697 DVDD.n772 DVDD.n771 0.00972131
R28698 DVDD.n4546 DVDD.n1084 0.00972131
R28699 DVDD.n3262 DVDD.n2958 0.00965
R28700 DVDD.n2935 DVDD.n2757 0.00965
R28701 DVDD.n2399 DVDD.n2398 0.00962857
R28702 DVDD.n2398 DVDD.n2043 0.00962857
R28703 DVDD.n2394 DVDD.n2043 0.00962857
R28704 DVDD.n2394 DVDD.n2045 0.00962857
R28705 DVDD.n2390 DVDD.n2045 0.00962857
R28706 DVDD.n2390 DVDD.n2047 0.00962857
R28707 DVDD.n2386 DVDD.n2047 0.00962857
R28708 DVDD.n2386 DVDD.n2049 0.00962857
R28709 DVDD.n2382 DVDD.n2049 0.00962857
R28710 DVDD.n2382 DVDD.n2051 0.00962857
R28711 DVDD.n2378 DVDD.n2051 0.00962857
R28712 DVDD.n2378 DVDD.n2053 0.00962857
R28713 DVDD.n2374 DVDD.n2053 0.00962857
R28714 DVDD.n2374 DVDD.n2055 0.00962857
R28715 DVDD.n2370 DVDD.n2055 0.00962857
R28716 DVDD.n2370 DVDD.n2057 0.00962857
R28717 DVDD.n2071 DVDD.n2057 0.00962857
R28718 DVDD.n2077 DVDD.n2071 0.00962857
R28719 DVDD.n2077 DVDD.n2069 0.00962857
R28720 DVDD.n2081 DVDD.n2069 0.00962857
R28721 DVDD.n2081 DVDD.n2067 0.00962857
R28722 DVDD.n2088 DVDD.n2067 0.00962857
R28723 DVDD.n2088 DVDD.n2064 0.00962857
R28724 DVDD.n2359 DVDD.n2064 0.00962857
R28725 DVDD.n2359 DVDD.n2065 0.00962857
R28726 DVDD.n2355 DVDD.n2065 0.00962857
R28727 DVDD.n2355 DVDD.n2092 0.00962857
R28728 DVDD.n2351 DVDD.n2092 0.00962857
R28729 DVDD.n2351 DVDD.n2095 0.00962857
R28730 DVDD.n2347 DVDD.n2095 0.00962857
R28731 DVDD.n2347 DVDD.n2097 0.00962857
R28732 DVDD.n2101 DVDD.n2097 0.00962857
R28733 DVDD.n2332 DVDD.n2101 0.00962857
R28734 DVDD.n2332 DVDD.n2102 0.00962857
R28735 DVDD.n2328 DVDD.n2102 0.00962857
R28736 DVDD.n2328 DVDD.n2105 0.00962857
R28737 DVDD.n2324 DVDD.n2105 0.00962857
R28738 DVDD.n2324 DVDD.n2107 0.00962857
R28739 DVDD.n2320 DVDD.n2107 0.00962857
R28740 DVDD.n2320 DVDD.n2109 0.00962857
R28741 DVDD.n2316 DVDD.n2109 0.00962857
R28742 DVDD.n2316 DVDD.n2111 0.00962857
R28743 DVDD.n2312 DVDD.n2111 0.00962857
R28744 DVDD.n2312 DVDD.n2113 0.00962857
R28745 DVDD.n2308 DVDD.n2113 0.00962857
R28746 DVDD.n2308 DVDD.n2115 0.00962857
R28747 DVDD.n2304 DVDD.n2115 0.00962857
R28748 DVDD.n2304 DVDD.n2117 0.00962857
R28749 DVDD.n2300 DVDD.n2117 0.00962857
R28750 DVDD.n2300 DVDD.n2119 0.00962857
R28751 DVDD.n2296 DVDD.n2119 0.00962857
R28752 DVDD.n2296 DVDD.n2121 0.00962857
R28753 DVDD.n2136 DVDD.n2121 0.00962857
R28754 DVDD.n2137 DVDD.n2136 0.00962857
R28755 DVDD.n2143 DVDD.n2137 0.00962857
R28756 DVDD.n2143 DVDD.n2133 0.00962857
R28757 DVDD.n2147 DVDD.n2133 0.00962857
R28758 DVDD.n2147 DVDD.n2131 0.00962857
R28759 DVDD.n2154 DVDD.n2131 0.00962857
R28760 DVDD.n2154 DVDD.n2128 0.00962857
R28761 DVDD.n2284 DVDD.n2128 0.00962857
R28762 DVDD.n2284 DVDD.n2129 0.00962857
R28763 DVDD.n2280 DVDD.n2129 0.00962857
R28764 DVDD.n2280 DVDD.n2158 0.00962857
R28765 DVDD.n2276 DVDD.n2158 0.00962857
R28766 DVDD.n2276 DVDD.n2161 0.00962857
R28767 DVDD.n2272 DVDD.n2161 0.00962857
R28768 DVDD.n2272 DVDD.n2163 0.00962857
R28769 DVDD.n2167 DVDD.n2163 0.00962857
R28770 DVDD.n2257 DVDD.n2167 0.00962857
R28771 DVDD.n2257 DVDD.n2168 0.00962857
R28772 DVDD.n2253 DVDD.n2168 0.00962857
R28773 DVDD.n2253 DVDD.n2171 0.00962857
R28774 DVDD.n2249 DVDD.n2171 0.00962857
R28775 DVDD.n2249 DVDD.n2173 0.00962857
R28776 DVDD.n2245 DVDD.n2173 0.00962857
R28777 DVDD.n2245 DVDD.n2175 0.00962857
R28778 DVDD.n2241 DVDD.n2175 0.00962857
R28779 DVDD.n2241 DVDD.n2177 0.00962857
R28780 DVDD.n2237 DVDD.n2177 0.00962857
R28781 DVDD.n2237 DVDD.n2179 0.00962857
R28782 DVDD.n2233 DVDD.n2179 0.00962857
R28783 DVDD.n2233 DVDD.n2181 0.00962857
R28784 DVDD.n2229 DVDD.n2181 0.00962857
R28785 DVDD.n2229 DVDD.n2183 0.00962857
R28786 DVDD.n2225 DVDD.n2183 0.00962857
R28787 DVDD.n2225 DVDD.n2185 0.00962857
R28788 DVDD.n2221 DVDD.n2185 0.00962857
R28789 DVDD.n2221 DVDD.n2187 0.00962857
R28790 DVDD.n2217 DVDD.n2187 0.00962857
R28791 DVDD.n2217 DVDD.n2189 0.00962857
R28792 DVDD.n2213 DVDD.n2189 0.00962857
R28793 DVDD.n2213 DVDD.n2191 0.00962857
R28794 DVDD.n2209 DVDD.n2191 0.00962857
R28795 DVDD.n2209 DVDD.n2193 0.00962857
R28796 DVDD.n2205 DVDD.n2193 0.00962857
R28797 DVDD.n2205 DVDD.n2195 0.00962857
R28798 DVDD.n2393 DVDD.n2004 0.00962857
R28799 DVDD.n2393 DVDD.n2392 0.00962857
R28800 DVDD.n2392 DVDD.n2391 0.00962857
R28801 DVDD.n2391 DVDD.n2046 0.00962857
R28802 DVDD.n2385 DVDD.n2046 0.00962857
R28803 DVDD.n2385 DVDD.n2384 0.00962857
R28804 DVDD.n2384 DVDD.n2383 0.00962857
R28805 DVDD.n2383 DVDD.n2050 0.00962857
R28806 DVDD.n2377 DVDD.n2050 0.00962857
R28807 DVDD.n2377 DVDD.n2376 0.00962857
R28808 DVDD.n2376 DVDD.n2375 0.00962857
R28809 DVDD.n2369 DVDD.n2058 0.00962857
R28810 DVDD.n2072 DVDD.n2059 0.00962857
R28811 DVDD.n2076 DVDD.n2072 0.00962857
R28812 DVDD.n2082 DVDD.n2068 0.00962857
R28813 DVDD.n2083 DVDD.n2082 0.00962857
R28814 DVDD.n2087 DVDD.n2083 0.00962857
R28815 DVDD.n2354 DVDD.n2093 0.00962857
R28816 DVDD.n2354 DVDD.n2353 0.00962857
R28817 DVDD.n2353 DVDD.n2352 0.00962857
R28818 DVDD.n2346 DVDD.n2098 0.00962857
R28819 DVDD.n2346 DVDD.n2345 0.00962857
R28820 DVDD.n2333 DVDD.n2100 0.00962857
R28821 DVDD.n2327 DVDD.n2100 0.00962857
R28822 DVDD.n2327 DVDD.n2326 0.00962857
R28823 DVDD.n2326 DVDD.n2325 0.00962857
R28824 DVDD.n2325 DVDD.n2106 0.00962857
R28825 DVDD.n2319 DVDD.n2106 0.00962857
R28826 DVDD.n2319 DVDD.n2318 0.00962857
R28827 DVDD.n2318 DVDD.n2317 0.00962857
R28828 DVDD.n2317 DVDD.n2110 0.00962857
R28829 DVDD.n2311 DVDD.n2110 0.00962857
R28830 DVDD.n2311 DVDD.n2310 0.00962857
R28831 DVDD.n2310 DVDD.n2309 0.00962857
R28832 DVDD.n2309 DVDD.n2114 0.00962857
R28833 DVDD.n2303 DVDD.n2114 0.00962857
R28834 DVDD.n2303 DVDD.n2302 0.00962857
R28835 DVDD.n2302 DVDD.n2301 0.00962857
R28836 DVDD.n2301 DVDD.n2118 0.00962857
R28837 DVDD.n2295 DVDD.n2294 0.00962857
R28838 DVDD.n2138 DVDD.n2123 0.00962857
R28839 DVDD.n2142 DVDD.n2138 0.00962857
R28840 DVDD.n2148 DVDD.n2132 0.00962857
R28841 DVDD.n2149 DVDD.n2148 0.00962857
R28842 DVDD.n2153 DVDD.n2149 0.00962857
R28843 DVDD.n2279 DVDD.n2159 0.00962857
R28844 DVDD.n2279 DVDD.n2278 0.00962857
R28845 DVDD.n2278 DVDD.n2277 0.00962857
R28846 DVDD.n2271 DVDD.n2164 0.00962857
R28847 DVDD.n2271 DVDD.n2270 0.00962857
R28848 DVDD.n2258 DVDD.n2166 0.00962857
R28849 DVDD.n2252 DVDD.n2166 0.00962857
R28850 DVDD.n2252 DVDD.n2251 0.00962857
R28851 DVDD.n2251 DVDD.n2250 0.00962857
R28852 DVDD.n2250 DVDD.n2172 0.00962857
R28853 DVDD.n2244 DVDD.n2172 0.00962857
R28854 DVDD.n2244 DVDD.n2243 0.00962857
R28855 DVDD.n2243 DVDD.n2242 0.00962857
R28856 DVDD.n2242 DVDD.n2176 0.00962857
R28857 DVDD.n2236 DVDD.n2176 0.00962857
R28858 DVDD.n2236 DVDD.n2235 0.00962857
R28859 DVDD.n2235 DVDD.n2234 0.00962857
R28860 DVDD.n2234 DVDD.n2180 0.00962857
R28861 DVDD.n2228 DVDD.n2180 0.00962857
R28862 DVDD.n2228 DVDD.n2227 0.00962857
R28863 DVDD.n2227 DVDD.n2226 0.00962857
R28864 DVDD.n2226 DVDD.n2184 0.00962857
R28865 DVDD.n2220 DVDD.n2184 0.00962857
R28866 DVDD.n2220 DVDD.n2219 0.00962857
R28867 DVDD.n2219 DVDD.n2218 0.00962857
R28868 DVDD.n2218 DVDD.n2188 0.00962857
R28869 DVDD.n2212 DVDD.n2188 0.00962857
R28870 DVDD.n2212 DVDD.n2211 0.00962857
R28871 DVDD.n2211 DVDD.n2210 0.00962857
R28872 DVDD.n2210 DVDD.n2192 0.00962857
R28873 DVDD.n2204 DVDD.n2192 0.00962857
R28874 DVDD.n3666 DVDD.n2406 0.00962857
R28875 DVDD.n3662 DVDD.n2406 0.00962857
R28876 DVDD.n3662 DVDD.n3661 0.00962857
R28877 DVDD.n3661 DVDD.n2408 0.00962857
R28878 DVDD.n3657 DVDD.n2408 0.00962857
R28879 DVDD.n3657 DVDD.n2410 0.00962857
R28880 DVDD.n3653 DVDD.n2410 0.00962857
R28881 DVDD.n3653 DVDD.n2413 0.00962857
R28882 DVDD.n3649 DVDD.n2413 0.00962857
R28883 DVDD.n3649 DVDD.n2415 0.00962857
R28884 DVDD.n3645 DVDD.n2415 0.00962857
R28885 DVDD.n3645 DVDD.n2417 0.00962857
R28886 DVDD.n3641 DVDD.n2417 0.00962857
R28887 DVDD.n3641 DVDD.n2419 0.00962857
R28888 DVDD.n3637 DVDD.n2419 0.00962857
R28889 DVDD.n3637 DVDD.n2421 0.00962857
R28890 DVDD.n3633 DVDD.n2421 0.00962857
R28891 DVDD.n3633 DVDD.n2423 0.00962857
R28892 DVDD.n3629 DVDD.n2423 0.00962857
R28893 DVDD.n3629 DVDD.n2425 0.00962857
R28894 DVDD.n3625 DVDD.n2425 0.00962857
R28895 DVDD.n3625 DVDD.n2427 0.00962857
R28896 DVDD.n3621 DVDD.n2427 0.00962857
R28897 DVDD.n3621 DVDD.n2429 0.00962857
R28898 DVDD.n3617 DVDD.n2429 0.00962857
R28899 DVDD.n3617 DVDD.n2434 0.00962857
R28900 DVDD.n3613 DVDD.n2434 0.00962857
R28901 DVDD.n3613 DVDD.n2436 0.00962857
R28902 DVDD.n3609 DVDD.n2436 0.00962857
R28903 DVDD.n3609 DVDD.n2439 0.00962857
R28904 DVDD.n3605 DVDD.n2439 0.00962857
R28905 DVDD.n3605 DVDD.n2441 0.00962857
R28906 DVDD.n3599 DVDD.n2441 0.00962857
R28907 DVDD.n3599 DVDD.n2456 0.00962857
R28908 DVDD.n3595 DVDD.n2456 0.00962857
R28909 DVDD.n3595 DVDD.n2458 0.00962857
R28910 DVDD.n3591 DVDD.n2458 0.00962857
R28911 DVDD.n3591 DVDD.n2460 0.00962857
R28912 DVDD.n3587 DVDD.n2460 0.00962857
R28913 DVDD.n3587 DVDD.n2462 0.00962857
R28914 DVDD.n3583 DVDD.n2462 0.00962857
R28915 DVDD.n3583 DVDD.n2464 0.00962857
R28916 DVDD.n3579 DVDD.n2464 0.00962857
R28917 DVDD.n3579 DVDD.n2466 0.00962857
R28918 DVDD.n3575 DVDD.n2466 0.00962857
R28919 DVDD.n3575 DVDD.n2468 0.00962857
R28920 DVDD.n3571 DVDD.n2468 0.00962857
R28921 DVDD.n3571 DVDD.n2470 0.00962857
R28922 DVDD.n3567 DVDD.n2470 0.00962857
R28923 DVDD.n3567 DVDD.n2472 0.00962857
R28924 DVDD.n3563 DVDD.n2472 0.00962857
R28925 DVDD.n3563 DVDD.n2474 0.00962857
R28926 DVDD.n3559 DVDD.n2474 0.00962857
R28927 DVDD.n3559 DVDD.n2476 0.00962857
R28928 DVDD.n3555 DVDD.n2476 0.00962857
R28929 DVDD.n3555 DVDD.n2478 0.00962857
R28930 DVDD.n3551 DVDD.n2478 0.00962857
R28931 DVDD.n3551 DVDD.n2480 0.00962857
R28932 DVDD.n3547 DVDD.n2480 0.00962857
R28933 DVDD.n3547 DVDD.n2482 0.00962857
R28934 DVDD.n3543 DVDD.n2482 0.00962857
R28935 DVDD.n3543 DVDD.n2484 0.00962857
R28936 DVDD.n3539 DVDD.n2484 0.00962857
R28937 DVDD.n3539 DVDD.n2486 0.00962857
R28938 DVDD.n3535 DVDD.n2486 0.00962857
R28939 DVDD.n3535 DVDD.n2488 0.00962857
R28940 DVDD.n3531 DVDD.n2488 0.00962857
R28941 DVDD.n3531 DVDD.n2490 0.00962857
R28942 DVDD.n2675 DVDD.n2490 0.00962857
R28943 DVDD.n2676 DVDD.n2675 0.00962857
R28944 DVDD.n2676 DVDD.n2671 0.00962857
R28945 DVDD.n3523 DVDD.n2671 0.00962857
R28946 DVDD.n3523 DVDD.n2673 0.00962857
R28947 DVDD.n3519 DVDD.n2673 0.00962857
R28948 DVDD.n3519 DVDD.n2680 0.00962857
R28949 DVDD.n3515 DVDD.n2680 0.00962857
R28950 DVDD.n3515 DVDD.n2682 0.00962857
R28951 DVDD.n3511 DVDD.n2682 0.00962857
R28952 DVDD.n3511 DVDD.n2684 0.00962857
R28953 DVDD.n3507 DVDD.n2684 0.00962857
R28954 DVDD.n3507 DVDD.n3453 0.00962857
R28955 DVDD.n3503 DVDD.n3453 0.00962857
R28956 DVDD.n3503 DVDD.n3455 0.00962857
R28957 DVDD.n3499 DVDD.n3455 0.00962857
R28958 DVDD.n3499 DVDD.n3457 0.00962857
R28959 DVDD.n3495 DVDD.n3457 0.00962857
R28960 DVDD.n3495 DVDD.n3459 0.00962857
R28961 DVDD.n3491 DVDD.n3459 0.00962857
R28962 DVDD.n3491 DVDD.n3461 0.00962857
R28963 DVDD.n3487 DVDD.n3461 0.00962857
R28964 DVDD.n3487 DVDD.n3463 0.00962857
R28965 DVDD.n3483 DVDD.n3463 0.00962857
R28966 DVDD.n3483 DVDD.n3465 0.00962857
R28967 DVDD.n3479 DVDD.n3465 0.00962857
R28968 DVDD.n3479 DVDD.n3467 0.00962857
R28969 DVDD.n3475 DVDD.n3467 0.00962857
R28970 DVDD.n3475 DVDD.n3469 0.00962857
R28971 DVDD.n3660 DVDD.n1988 0.00962857
R28972 DVDD.n3660 DVDD.n3659 0.00962857
R28973 DVDD.n3659 DVDD.n3658 0.00962857
R28974 DVDD.n3658 DVDD.n2409 0.00962857
R28975 DVDD.n3652 DVDD.n2409 0.00962857
R28976 DVDD.n3652 DVDD.n3651 0.00962857
R28977 DVDD.n3651 DVDD.n3650 0.00962857
R28978 DVDD.n3650 DVDD.n2414 0.00962857
R28979 DVDD.n3644 DVDD.n2414 0.00962857
R28980 DVDD.n3644 DVDD.n3643 0.00962857
R28981 DVDD.n3643 DVDD.n3642 0.00962857
R28982 DVDD.n3642 DVDD.n2418 0.00962857
R28983 DVDD.n3636 DVDD.n2418 0.00962857
R28984 DVDD.n3636 DVDD.n3635 0.00962857
R28985 DVDD.n3635 DVDD.n3634 0.00962857
R28986 DVDD.n3634 DVDD.n2422 0.00962857
R28987 DVDD.n3628 DVDD.n2422 0.00962857
R28988 DVDD.n3628 DVDD.n3627 0.00962857
R28989 DVDD.n3627 DVDD.n3626 0.00962857
R28990 DVDD.n3626 DVDD.n2426 0.00962857
R28991 DVDD.n3620 DVDD.n2426 0.00962857
R28992 DVDD.n3620 DVDD.n3619 0.00962857
R28993 DVDD.n3619 DVDD.n3618 0.00962857
R28994 DVDD.n3612 DVDD.n2437 0.00962857
R28995 DVDD.n3612 DVDD.n3611 0.00962857
R28996 DVDD.n3611 DVDD.n3610 0.00962857
R28997 DVDD.n3610 DVDD.n2438 0.00962857
R28998 DVDD.n3600 DVDD.n2455 0.00962857
R28999 DVDD.n3594 DVDD.n2455 0.00962857
R29000 DVDD.n3594 DVDD.n3593 0.00962857
R29001 DVDD.n3593 DVDD.n3592 0.00962857
R29002 DVDD.n3592 DVDD.n2459 0.00962857
R29003 DVDD.n3586 DVDD.n2459 0.00962857
R29004 DVDD.n3586 DVDD.n3585 0.00962857
R29005 DVDD.n3585 DVDD.n3584 0.00962857
R29006 DVDD.n3584 DVDD.n2463 0.00962857
R29007 DVDD.n3578 DVDD.n2463 0.00962857
R29008 DVDD.n3578 DVDD.n3577 0.00962857
R29009 DVDD.n3577 DVDD.n3576 0.00962857
R29010 DVDD.n3576 DVDD.n2467 0.00962857
R29011 DVDD.n3570 DVDD.n2467 0.00962857
R29012 DVDD.n3570 DVDD.n3569 0.00962857
R29013 DVDD.n3569 DVDD.n3568 0.00962857
R29014 DVDD.n3568 DVDD.n2471 0.00962857
R29015 DVDD.n3562 DVDD.n2471 0.00962857
R29016 DVDD.n3562 DVDD.n3561 0.00962857
R29017 DVDD.n3561 DVDD.n3560 0.00962857
R29018 DVDD.n3560 DVDD.n2475 0.00962857
R29019 DVDD.n3554 DVDD.n2475 0.00962857
R29020 DVDD.n3554 DVDD.n3553 0.00962857
R29021 DVDD.n3553 DVDD.n3552 0.00962857
R29022 DVDD.n3552 DVDD.n2479 0.00962857
R29023 DVDD.n3546 DVDD.n2479 0.00962857
R29024 DVDD.n3546 DVDD.n3545 0.00962857
R29025 DVDD.n3545 DVDD.n3544 0.00962857
R29026 DVDD.n3544 DVDD.n2483 0.00962857
R29027 DVDD.n3538 DVDD.n2483 0.00962857
R29028 DVDD.n3538 DVDD.n3537 0.00962857
R29029 DVDD.n3537 DVDD.n3536 0.00962857
R29030 DVDD.n3536 DVDD.n2487 0.00962857
R29031 DVDD.n3530 DVDD.n2487 0.00962857
R29032 DVDD.n3530 DVDD.n3529 0.00962857
R29033 DVDD.n3525 DVDD.n3524 0.00962857
R29034 DVDD.n3524 DVDD.n2672 0.00962857
R29035 DVDD.n3518 DVDD.n2672 0.00962857
R29036 DVDD.n3518 DVDD.n3517 0.00962857
R29037 DVDD.n3517 DVDD.n3516 0.00962857
R29038 DVDD.n3516 DVDD.n2681 0.00962857
R29039 DVDD.n3510 DVDD.n3509 0.00962857
R29040 DVDD.n3509 DVDD.n3508 0.00962857
R29041 DVDD.n3508 DVDD.n3452 0.00962857
R29042 DVDD.n3502 DVDD.n3452 0.00962857
R29043 DVDD.n3502 DVDD.n3501 0.00962857
R29044 DVDD.n3501 DVDD.n3500 0.00962857
R29045 DVDD.n3500 DVDD.n3456 0.00962857
R29046 DVDD.n3494 DVDD.n3456 0.00962857
R29047 DVDD.n3494 DVDD.n3493 0.00962857
R29048 DVDD.n3493 DVDD.n3492 0.00962857
R29049 DVDD.n3492 DVDD.n3460 0.00962857
R29050 DVDD.n3486 DVDD.n3460 0.00962857
R29051 DVDD.n3486 DVDD.n3485 0.00962857
R29052 DVDD.n3485 DVDD.n3484 0.00962857
R29053 DVDD.n3484 DVDD.n3464 0.00962857
R29054 DVDD.n3478 DVDD.n3464 0.00962857
R29055 DVDD.n3478 DVDD.n3477 0.00962857
R29056 DVDD.n3477 DVDD.n3476 0.00962857
R29057 DVDD.n3476 DVDD.n3468 0.00962857
R29058 DVDD.n1571 DVDD.n1205 0.00962857
R29059 DVDD.n1571 DVDD.n1206 0.00962857
R29060 DVDD.n1567 DVDD.n1206 0.00962857
R29061 DVDD.n1567 DVDD.n1208 0.00962857
R29062 DVDD.n1563 DVDD.n1208 0.00962857
R29063 DVDD.n1563 DVDD.n1211 0.00962857
R29064 DVDD.n1559 DVDD.n1211 0.00962857
R29065 DVDD.n1559 DVDD.n1213 0.00962857
R29066 DVDD.n1224 DVDD.n1213 0.00962857
R29067 DVDD.n1552 DVDD.n1224 0.00962857
R29068 DVDD.n1552 DVDD.n1225 0.00962857
R29069 DVDD.n1548 DVDD.n1225 0.00962857
R29070 DVDD.n1548 DVDD.n1228 0.00962857
R29071 DVDD.n1544 DVDD.n1228 0.00962857
R29072 DVDD.n1544 DVDD.n1230 0.00962857
R29073 DVDD.n1540 DVDD.n1230 0.00962857
R29074 DVDD.n1540 DVDD.n1232 0.00962857
R29075 DVDD.n1536 DVDD.n1232 0.00962857
R29076 DVDD.n1536 DVDD.n1234 0.00962857
R29077 DVDD.n1532 DVDD.n1234 0.00962857
R29078 DVDD.n1532 DVDD.n1236 0.00962857
R29079 DVDD.n1528 DVDD.n1236 0.00962857
R29080 DVDD.n1528 DVDD.n1238 0.00962857
R29081 DVDD.n1524 DVDD.n1238 0.00962857
R29082 DVDD.n1524 DVDD.n1240 0.00962857
R29083 DVDD.n1520 DVDD.n1240 0.00962857
R29084 DVDD.n1520 DVDD.n1242 0.00962857
R29085 DVDD.n1516 DVDD.n1242 0.00962857
R29086 DVDD.n1516 DVDD.n1244 0.00962857
R29087 DVDD.n1512 DVDD.n1244 0.00962857
R29088 DVDD.n1512 DVDD.n1246 0.00962857
R29089 DVDD.n1508 DVDD.n1246 0.00962857
R29090 DVDD.n1508 DVDD.n1248 0.00962857
R29091 DVDD.n1504 DVDD.n1248 0.00962857
R29092 DVDD.n1504 DVDD.n1250 0.00962857
R29093 DVDD.n1500 DVDD.n1250 0.00962857
R29094 DVDD.n1500 DVDD.n1252 0.00962857
R29095 DVDD.n1496 DVDD.n1252 0.00962857
R29096 DVDD.n1496 DVDD.n1254 0.00962857
R29097 DVDD.n1492 DVDD.n1254 0.00962857
R29098 DVDD.n1492 DVDD.n1256 0.00962857
R29099 DVDD.n1488 DVDD.n1256 0.00962857
R29100 DVDD.n1488 DVDD.n1258 0.00962857
R29101 DVDD.n1484 DVDD.n1258 0.00962857
R29102 DVDD.n1484 DVDD.n1260 0.00962857
R29103 DVDD.n1480 DVDD.n1260 0.00962857
R29104 DVDD.n1480 DVDD.n1262 0.00962857
R29105 DVDD.n1476 DVDD.n1262 0.00962857
R29106 DVDD.n1476 DVDD.n1264 0.00962857
R29107 DVDD.n1472 DVDD.n1264 0.00962857
R29108 DVDD.n1472 DVDD.n1266 0.00962857
R29109 DVDD.n1468 DVDD.n1266 0.00962857
R29110 DVDD.n1468 DVDD.n1268 0.00962857
R29111 DVDD.n1464 DVDD.n1268 0.00962857
R29112 DVDD.n1464 DVDD.n1270 0.00962857
R29113 DVDD.n1460 DVDD.n1270 0.00962857
R29114 DVDD.n1460 DVDD.n1272 0.00962857
R29115 DVDD.n1456 DVDD.n1272 0.00962857
R29116 DVDD.n1456 DVDD.n1274 0.00962857
R29117 DVDD.n1452 DVDD.n1274 0.00962857
R29118 DVDD.n1452 DVDD.n1276 0.00962857
R29119 DVDD.n1448 DVDD.n1276 0.00962857
R29120 DVDD.n1448 DVDD.n1278 0.00962857
R29121 DVDD.n1444 DVDD.n1278 0.00962857
R29122 DVDD.n1444 DVDD.n1280 0.00962857
R29123 DVDD.n1440 DVDD.n1280 0.00962857
R29124 DVDD.n1440 DVDD.n1282 0.00962857
R29125 DVDD.n1436 DVDD.n1282 0.00962857
R29126 DVDD.n1436 DVDD.n1284 0.00962857
R29127 DVDD.n1432 DVDD.n1284 0.00962857
R29128 DVDD.n1432 DVDD.n1286 0.00962857
R29129 DVDD.n1428 DVDD.n1286 0.00962857
R29130 DVDD.n1428 DVDD.n1288 0.00962857
R29131 DVDD.n1424 DVDD.n1288 0.00962857
R29132 DVDD.n1424 DVDD.n1290 0.00962857
R29133 DVDD.n1420 DVDD.n1290 0.00962857
R29134 DVDD.n1420 DVDD.n1292 0.00962857
R29135 DVDD.n1416 DVDD.n1292 0.00962857
R29136 DVDD.n1416 DVDD.n1294 0.00962857
R29137 DVDD.n1412 DVDD.n1294 0.00962857
R29138 DVDD.n1412 DVDD.n1296 0.00962857
R29139 DVDD.n1408 DVDD.n1296 0.00962857
R29140 DVDD.n1408 DVDD.n1298 0.00962857
R29141 DVDD.n1404 DVDD.n1298 0.00962857
R29142 DVDD.n1404 DVDD.n1300 0.00962857
R29143 DVDD.n1400 DVDD.n1300 0.00962857
R29144 DVDD.n1400 DVDD.n1302 0.00962857
R29145 DVDD.n1396 DVDD.n1302 0.00962857
R29146 DVDD.n1396 DVDD.n1304 0.00962857
R29147 DVDD.n1347 DVDD.n1304 0.00962857
R29148 DVDD.n1350 DVDD.n1347 0.00962857
R29149 DVDD.n1350 DVDD.n1345 0.00962857
R29150 DVDD.n1354 DVDD.n1345 0.00962857
R29151 DVDD.n1354 DVDD.n1343 0.00962857
R29152 DVDD.n1358 DVDD.n1343 0.00962857
R29153 DVDD.n1362 DVDD.n1361 0.00962857
R29154 DVDD.n1566 DVDD.n1209 0.00962857
R29155 DVDD.n1566 DVDD.n1565 0.00962857
R29156 DVDD.n1565 DVDD.n1564 0.00962857
R29157 DVDD.n1564 DVDD.n1210 0.00962857
R29158 DVDD.n1558 DVDD.n1210 0.00962857
R29159 DVDD.n1558 DVDD.n1557 0.00962857
R29160 DVDD.n1553 DVDD.n1223 0.00962857
R29161 DVDD.n1547 DVDD.n1223 0.00962857
R29162 DVDD.n1547 DVDD.n1546 0.00962857
R29163 DVDD.n1546 DVDD.n1545 0.00962857
R29164 DVDD.n1545 DVDD.n1229 0.00962857
R29165 DVDD.n1539 DVDD.n1229 0.00962857
R29166 DVDD.n1539 DVDD.n1538 0.00962857
R29167 DVDD.n1538 DVDD.n1537 0.00962857
R29168 DVDD.n1537 DVDD.n1233 0.00962857
R29169 DVDD.n1531 DVDD.n1233 0.00962857
R29170 DVDD.n1531 DVDD.n1530 0.00962857
R29171 DVDD.n1530 DVDD.n1529 0.00962857
R29172 DVDD.n1529 DVDD.n1237 0.00962857
R29173 DVDD.n1523 DVDD.n1237 0.00962857
R29174 DVDD.n1523 DVDD.n1522 0.00962857
R29175 DVDD.n1522 DVDD.n1521 0.00962857
R29176 DVDD.n1521 DVDD.n1241 0.00962857
R29177 DVDD.n1515 DVDD.n1241 0.00962857
R29178 DVDD.n1515 DVDD.n1514 0.00962857
R29179 DVDD.n1514 DVDD.n1513 0.00962857
R29180 DVDD.n1513 DVDD.n1245 0.00962857
R29181 DVDD.n1507 DVDD.n1245 0.00962857
R29182 DVDD.n1507 DVDD.n1506 0.00962857
R29183 DVDD.n1506 DVDD.n1505 0.00962857
R29184 DVDD.n1505 DVDD.n1249 0.00962857
R29185 DVDD.n1499 DVDD.n1249 0.00962857
R29186 DVDD.n1499 DVDD.n1498 0.00962857
R29187 DVDD.n1498 DVDD.n1497 0.00962857
R29188 DVDD.n1497 DVDD.n1253 0.00962857
R29189 DVDD.n1491 DVDD.n1253 0.00962857
R29190 DVDD.n1491 DVDD.n1490 0.00962857
R29191 DVDD.n1490 DVDD.n1489 0.00962857
R29192 DVDD.n1489 DVDD.n1257 0.00962857
R29193 DVDD.n1483 DVDD.n1257 0.00962857
R29194 DVDD.n1483 DVDD.n1482 0.00962857
R29195 DVDD.n1482 DVDD.n1481 0.00962857
R29196 DVDD.n1481 DVDD.n1261 0.00962857
R29197 DVDD.n1475 DVDD.n1261 0.00962857
R29198 DVDD.n1475 DVDD.n1474 0.00962857
R29199 DVDD.n1474 DVDD.n1473 0.00962857
R29200 DVDD.n1473 DVDD.n1265 0.00962857
R29201 DVDD.n1467 DVDD.n1265 0.00962857
R29202 DVDD.n1467 DVDD.n1466 0.00962857
R29203 DVDD.n1466 DVDD.n1465 0.00962857
R29204 DVDD.n1465 DVDD.n1269 0.00962857
R29205 DVDD.n1459 DVDD.n1269 0.00962857
R29206 DVDD.n1459 DVDD.n1458 0.00962857
R29207 DVDD.n1458 DVDD.n1457 0.00962857
R29208 DVDD.n1457 DVDD.n1273 0.00962857
R29209 DVDD.n1451 DVDD.n1273 0.00962857
R29210 DVDD.n1451 DVDD.n1450 0.00962857
R29211 DVDD.n1450 DVDD.n1449 0.00962857
R29212 DVDD.n1449 DVDD.n1277 0.00962857
R29213 DVDD.n1443 DVDD.n1277 0.00962857
R29214 DVDD.n1443 DVDD.n1442 0.00962857
R29215 DVDD.n1442 DVDD.n1441 0.00962857
R29216 DVDD.n1441 DVDD.n1281 0.00962857
R29217 DVDD.n1435 DVDD.n1281 0.00962857
R29218 DVDD.n1435 DVDD.n1434 0.00962857
R29219 DVDD.n1434 DVDD.n1433 0.00962857
R29220 DVDD.n1433 DVDD.n1285 0.00962857
R29221 DVDD.n1427 DVDD.n1285 0.00962857
R29222 DVDD.n1427 DVDD.n1426 0.00962857
R29223 DVDD.n1426 DVDD.n1425 0.00962857
R29224 DVDD.n1425 DVDD.n1289 0.00962857
R29225 DVDD.n1419 DVDD.n1289 0.00962857
R29226 DVDD.n1419 DVDD.n1418 0.00962857
R29227 DVDD.n1418 DVDD.n1417 0.00962857
R29228 DVDD.n1417 DVDD.n1293 0.00962857
R29229 DVDD.n1411 DVDD.n1293 0.00962857
R29230 DVDD.n1411 DVDD.n1410 0.00962857
R29231 DVDD.n1410 DVDD.n1409 0.00962857
R29232 DVDD.n1409 DVDD.n1297 0.00962857
R29233 DVDD.n1403 DVDD.n1297 0.00962857
R29234 DVDD.n1403 DVDD.n1402 0.00962857
R29235 DVDD.n1402 DVDD.n1401 0.00962857
R29236 DVDD.n1401 DVDD.n1301 0.00962857
R29237 DVDD.n1348 DVDD.n1310 0.00962857
R29238 DVDD.n1349 DVDD.n1348 0.00962857
R29239 DVDD.n1349 DVDD.n1344 0.00962857
R29240 DVDD.n1355 DVDD.n1344 0.00962857
R29241 DVDD.n1356 DVDD.n1355 0.00962857
R29242 DVDD.n1357 DVDD.n1356 0.00962857
R29243 DVDD.n2730 DVDD.n2725 0.00959
R29244 DVDD.n1337 DVDD.n1331 0.00956429
R29245 DVDD.n1364 DVDD.n1340 0.00956429
R29246 DVDD.n5426 DVDD.n333 0.00955202
R29247 DVDD.n2849 DVDD.n2782 0.00954891
R29248 DVDD.n2853 DVDD.n2797 0.00954891
R29249 DVDD.n2883 DVDD.n2874 0.00954891
R29250 DVDD.n2887 DVDD.n2868 0.00954891
R29251 DVDD.n86 DVDD.n85 0.00953114
R29252 DVDD.n5523 DVDD.n10 0.00948451
R29253 DVDD.n4693 DVDD.n977 0.00948451
R29254 DVDD.n3250 DVDD.n3086 0.00941892
R29255 DVDD.n3207 DVDD.n3206 0.00941892
R29256 DVDD.n5764 DVDD.n184 0.00935246
R29257 DVDD.n5222 DVDD.n490 0.00935246
R29258 DVDD.n646 DVDD.n620 0.00935246
R29259 DVDD.n846 DVDD.n709 0.00935246
R29260 DVDD.n4595 DVDD.n1014 0.00935246
R29261 DVDD.n3320 DVDD.n2861 0.00935
R29262 DVDD.n3346 DVDD.n2776 0.00935
R29263 DVDD.n3071 DVDD.n2991 0.00935
R29264 DVDD.n5509 DVDD.n222 0.0093296
R29265 DVDD.n948 DVDD.n946 0.0093296
R29266 DVDD.n2626 DVDD.n2452 0.00930435
R29267 DVDD.n2375 DVDD.n2054 0.00917857
R29268 DVDD.n5932 DVDD.n70 0.0091747
R29269 DVDD.n5476 DVDD.n294 0.0091747
R29270 DVDD.n110 DVDD.n89 0.00908247
R29271 DVDD.n5915 DVDD.n94 0.00908247
R29272 DVDD.n5408 DVDD.n343 0.00908247
R29273 DVDD.n5419 DVDD.n5418 0.00908247
R29274 DVDD.n927 DVDD.n915 0.00908247
R29275 DVDD.n4711 DVDD.n942 0.00908247
R29276 DVDD.n257 DVDD.n235 0.00908247
R29277 DVDD.n244 DVDD.n228 0.00908247
R29278 DVDD.n2658 DVDD.n2497 0.00905
R29279 DVDD.n4678 DVDD.n4677 0.00903179
R29280 DVDD.n5541 DVDD.n5539 0.00901211
R29281 DVDD.n5811 DVDD.n159 0.00898361
R29282 DVDD.n5167 DVDD.n459 0.00898361
R29283 DVDD.n4974 DVDD.n681 0.00898361
R29284 DVDD.n790 DVDD.n749 0.00898361
R29285 DVDD.n4530 DVDD.n1082 0.00898361
R29286 DVDD.n2152 DVDD.n2126 0.00892143
R29287 DVDD.n2164 DVDD.n2160 0.00892143
R29288 DVDD.n5625 DVDD.n5606 0.00886489
R29289 DVDD.n5450 DVDD.n288 0.00886489
R29290 DVDD.n3296 DVDD.n2924 0.00881522
R29291 DVDD.n3325 DVDD.n2917 0.00881522
R29292 DVDD.n3366 DVDD.n2767 0.00881522
R29293 DVDD.n2809 DVDD.n2806 0.00881522
R29294 DVDD.n2819 DVDD.n2788 0.00881522
R29295 DVDD.n3335 DVDD.n2871 0.00881522
R29296 DVDD.n2334 DVDD.n2099 0.00879286
R29297 DVDD.n3529 DVDD.n3528 0.00879286
R29298 DVDD.n2500 DVDD.n2495 0.00879286
R29299 DVDD.n3526 DVDD.n2670 0.00879286
R29300 DVDD.n1556 DVDD.n1218 0.00879286
R29301 DVDD.n1554 DVDD.n1553 0.00879286
R29302 DVDD.n2750 DVDD.n2736 0.00868173
R29303 DVDD.n112 DVDD.n91 0.00861856
R29304 DVDD.n5910 DVDD.n93 0.00861856
R29305 DVDD.n5410 DVDD.n345 0.00861856
R29306 DVDD.n5413 DVDD.n347 0.00861856
R29307 DVDD.n933 DVDD.n917 0.00861856
R29308 DVDD.n952 DVDD.n924 0.00861856
R29309 DVDD.n5670 DVDD.n236 0.00861856
R29310 DVDD.n252 DVDD.n230 0.00861856
R29311 DVDD.n5748 DVDD.n186 0.00861475
R29312 DVDD.n5238 DVDD.n565 0.00861475
R29313 DVDD.n630 DVDD.n622 0.00861475
R29314 DVDD.n862 DVDD.n725 0.00861475
R29315 DVDD.n4611 DVDD.n1056 0.00861475
R29316 DVDD.n2662 DVDD.n2493 0.0086
R29317 DVDD.n5642 DVDD.n5570 0.00855508
R29318 DVDD.n5467 DVDD.n277 0.00855508
R29319 DVDD.n2400 DVDD.n1997 0.00853571
R29320 DVDD.n2404 DVDD.n1999 0.00853571
R29321 DVDD.n2122 DVDD.n2118 0.00853571
R29322 DVDD.n3671 DVDD.n3667 0.00853571
R29323 DVDD.n3674 DVDD.n1983 0.00853571
R29324 DVDD.n3604 DVDD.n2442 0.00853571
R29325 DVDD.n3603 DVDD.n2448 0.00853571
R29326 DVDD.n3601 DVDD.n3600 0.00853571
R29327 DVDD.n3451 DVDD.n2681 0.00853571
R29328 DVDD.n4079 DVDD.n4078 0.0084875
R29329 DVDD.n4078 DVDD.n4048 0.0084875
R29330 DVDD.n4074 DVDD.n4048 0.0084875
R29331 DVDD.n4074 DVDD.n4050 0.0084875
R29332 DVDD.n4070 DVDD.n4050 0.0084875
R29333 DVDD.n4070 DVDD.n4053 0.0084875
R29334 DVDD.n4063 DVDD.n4053 0.0084875
R29335 DVDD.n4063 DVDD.n4060 0.0084875
R29336 DVDD.n4060 DVDD.n1723 0.0084875
R29337 DVDD.n4225 DVDD.n1723 0.0084875
R29338 DVDD.n1765 DVDD.n1727 0.0084875
R29339 DVDD.n1758 DVDD.n1727 0.0084875
R29340 DVDD.n1758 DVDD.n1731 0.0084875
R29341 DVDD.n1754 DVDD.n1731 0.0084875
R29342 DVDD.n1754 DVDD.n1733 0.0084875
R29343 DVDD.n1750 DVDD.n1733 0.0084875
R29344 DVDD.n1750 DVDD.n1736 0.0084875
R29345 DVDD.n1746 DVDD.n1736 0.0084875
R29346 DVDD.n1746 DVDD.n1738 0.0084875
R29347 DVDD.n4077 DVDD.n4044 0.0084875
R29348 DVDD.n4077 DVDD.n4076 0.0084875
R29349 DVDD.n4076 DVDD.n4075 0.0084875
R29350 DVDD.n4075 DVDD.n4049 0.0084875
R29351 DVDD.n1753 DVDD.n1734 0.0084875
R29352 DVDD.n1753 DVDD.n1752 0.0084875
R29353 DVDD.n1752 DVDD.n1751 0.0084875
R29354 DVDD.n1751 DVDD.n1735 0.0084875
R29355 DVDD.n1745 DVDD.n1735 0.0084875
R29356 DVDD.n1745 DVDD.n1744 0.0084875
R29357 DVDD.n3900 DVDD.n3899 0.0084875
R29358 DVDD.n3899 DVDD.n3898 0.0084875
R29359 DVDD.n3898 DVDD.n3873 0.0084875
R29360 DVDD.n3892 DVDD.n3873 0.0084875
R29361 DVDD.n3892 DVDD.n3891 0.0084875
R29362 DVDD.n3891 DVDD.n3890 0.0084875
R29363 DVDD.n3890 DVDD.n3878 0.0084875
R29364 DVDD.n3884 DVDD.n3878 0.0084875
R29365 DVDD.n3884 DVDD.n3883 0.0084875
R29366 DVDD.n3883 DVDD.n1794 0.0084875
R29367 DVDD.n4101 DVDD.n4100 0.0084875
R29368 DVDD.n4100 DVDD.n4099 0.0084875
R29369 DVDD.n4099 DVDD.n4036 0.0084875
R29370 DVDD.n4093 DVDD.n4036 0.0084875
R29371 DVDD.n4093 DVDD.n4092 0.0084875
R29372 DVDD.n4092 DVDD.n4091 0.0084875
R29373 DVDD.n4091 DVDD.n4040 0.0084875
R29374 DVDD.n4085 DVDD.n4040 0.0084875
R29375 DVDD.n4085 DVDD.n4084 0.0084875
R29376 DVDD.n3901 DVDD.n3872 0.0084875
R29377 DVDD.n3897 DVDD.n3872 0.0084875
R29378 DVDD.n3897 DVDD.n3874 0.0084875
R29379 DVDD.n3893 DVDD.n3874 0.0084875
R29380 DVDD.n3893 DVDD.n3877 0.0084875
R29381 DVDD.n3889 DVDD.n3877 0.0084875
R29382 DVDD.n3889 DVDD.n3879 0.0084875
R29383 DVDD.n3885 DVDD.n3879 0.0084875
R29384 DVDD.n3885 DVDD.n3882 0.0084875
R29385 DVDD.n3882 DVDD.n3881 0.0084875
R29386 DVDD.n4102 DVDD.n1793 0.0084875
R29387 DVDD.n4098 DVDD.n1793 0.0084875
R29388 DVDD.n4098 DVDD.n4037 0.0084875
R29389 DVDD.n4094 DVDD.n4037 0.0084875
R29390 DVDD.n4094 DVDD.n4039 0.0084875
R29391 DVDD.n4090 DVDD.n4039 0.0084875
R29392 DVDD.n4090 DVDD.n4041 0.0084875
R29393 DVDD.n4086 DVDD.n4041 0.0084875
R29394 DVDD.n4086 DVDD.n4043 0.0084875
R29395 DVDD.n3837 DVDD.n1828 0.0084875
R29396 DVDD.n3841 DVDD.n1828 0.0084875
R29397 DVDD.n3841 DVDD.n1826 0.0084875
R29398 DVDD.n3845 DVDD.n1826 0.0084875
R29399 DVDD.n3845 DVDD.n1824 0.0084875
R29400 DVDD.n3849 DVDD.n1824 0.0084875
R29401 DVDD.n3849 DVDD.n1822 0.0084875
R29402 DVDD.n3853 DVDD.n1822 0.0084875
R29403 DVDD.n3853 DVDD.n1820 0.0084875
R29404 DVDD.n3857 DVDD.n1820 0.0084875
R29405 DVDD.n3923 DVDD.n3860 0.0084875
R29406 DVDD.n3919 DVDD.n3860 0.0084875
R29407 DVDD.n3919 DVDD.n3862 0.0084875
R29408 DVDD.n3915 DVDD.n3862 0.0084875
R29409 DVDD.n3915 DVDD.n3864 0.0084875
R29410 DVDD.n3911 DVDD.n3864 0.0084875
R29411 DVDD.n3911 DVDD.n3866 0.0084875
R29412 DVDD.n3907 DVDD.n3866 0.0084875
R29413 DVDD.n3907 DVDD.n3868 0.0084875
R29414 DVDD.n4285 DVDD.n1669 0.0084875
R29415 DVDD.n4281 DVDD.n1669 0.0084875
R29416 DVDD.n4281 DVDD.n1672 0.0084875
R29417 DVDD.n4277 DVDD.n1672 0.0084875
R29418 DVDD.n4277 DVDD.n1674 0.0084875
R29419 DVDD.n4273 DVDD.n1674 0.0084875
R29420 DVDD.n4273 DVDD.n1676 0.0084875
R29421 DVDD.n4269 DVDD.n1676 0.0084875
R29422 DVDD.n4269 DVDD.n1678 0.0084875
R29423 DVDD.n4262 DVDD.n1678 0.0084875
R29424 DVDD.n3811 DVDD.n3809 0.0084875
R29425 DVDD.n3811 DVDD.n1839 0.0084875
R29426 DVDD.n3820 DVDD.n1839 0.0084875
R29427 DVDD.n3820 DVDD.n1837 0.0084875
R29428 DVDD.n3824 DVDD.n1837 0.0084875
R29429 DVDD.n3824 DVDD.n1835 0.0084875
R29430 DVDD.n3828 DVDD.n1835 0.0084875
R29431 DVDD.n3828 DVDD.n1833 0.0084875
R29432 DVDD.n3832 DVDD.n1833 0.0084875
R29433 DVDD.n3836 DVDD.n1827 0.0084875
R29434 DVDD.n3842 DVDD.n1827 0.0084875
R29435 DVDD.n3843 DVDD.n3842 0.0084875
R29436 DVDD.n3844 DVDD.n3843 0.0084875
R29437 DVDD.n3844 DVDD.n1823 0.0084875
R29438 DVDD.n3850 DVDD.n1823 0.0084875
R29439 DVDD.n3851 DVDD.n3850 0.0084875
R29440 DVDD.n3852 DVDD.n3851 0.0084875
R29441 DVDD.n3852 DVDD.n1819 0.0084875
R29442 DVDD.n3858 DVDD.n1819 0.0084875
R29443 DVDD.n3924 DVDD.n3859 0.0084875
R29444 DVDD.n3918 DVDD.n3859 0.0084875
R29445 DVDD.n3918 DVDD.n3917 0.0084875
R29446 DVDD.n3917 DVDD.n3916 0.0084875
R29447 DVDD.n3916 DVDD.n3863 0.0084875
R29448 DVDD.n3910 DVDD.n3863 0.0084875
R29449 DVDD.n3910 DVDD.n3909 0.0084875
R29450 DVDD.n3909 DVDD.n3908 0.0084875
R29451 DVDD.n3908 DVDD.n3867 0.0084875
R29452 DVDD.n4284 DVDD.n4283 0.0084875
R29453 DVDD.n4283 DVDD.n4282 0.0084875
R29454 DVDD.n4282 DVDD.n1671 0.0084875
R29455 DVDD.n4276 DVDD.n1671 0.0084875
R29456 DVDD.n4276 DVDD.n4275 0.0084875
R29457 DVDD.n4275 DVDD.n4274 0.0084875
R29458 DVDD.n3826 DVDD.n3825 0.0084875
R29459 DVDD.n3827 DVDD.n3826 0.0084875
R29460 DVDD.n3827 DVDD.n1832 0.0084875
R29461 DVDD.n3833 DVDD.n1832 0.0084875
R29462 DVDD.n5653 DVDD.n68 0.00840017
R29463 DVDD.n5479 DVDD.n270 0.00840017
R29464 DVDD.n3689 DVDD.n1896 0.00832155
R29465 DVDD.n3691 DVDD.n3690 0.00832155
R29466 DVDD.n4289 DVDD.n1666 0.00832155
R29467 DVDD.n3680 DVDD.n3679 0.00830425
R29468 DVDD.n3719 DVDD.n1890 0.00830425
R29469 DVDD.n3773 DVDD.n3757 0.00830425
R29470 DVDD.n4299 DVDD.n1660 0.00830425
R29471 DVDD.n968 DVDD.n966 0.00830347
R29472 DVDD.n5508 DVDD.n5506 0.00828547
R29473 DVDD.n2086 DVDD.n2062 0.00827857
R29474 DVDD.n2098 DVDD.n2094 0.00827857
R29475 DVDD.n5827 DVDD.n147 0.0082459
R29476 DVDD.n5183 DVDD.n457 0.0082459
R29477 DVDD.n4958 DVDD.n679 0.0082459
R29478 DVDD.n807 DVDD.n806 0.0082459
R29479 DVDD.n4514 DVDD.n1080 0.0082459
R29480 DVDD.n2259 DVDD.n2165 0.00815
R29481 DVDD.n5638 DVDD.n52 0.00809036
R29482 DVDD.n5504 DVDD.n219 0.00809036
R29483 DVDD.n964 DVDD.n945 0.00809036
R29484 DVDD.n5463 DVDD.n314 0.00809036
R29485 DVDD.n2846 DVDD.n2783 0.00808152
R29486 DVDD.n3347 DVDD.n2798 0.00808152
R29487 DVDD.n3342 DVDD.n2860 0.00808152
R29488 DVDD.n2891 DVDD.n2867 0.00808152
R29489 DVDD.n930 DVDD.n264 0.00804054
R29490 DVDD.n951 DVDD.n264 0.00804054
R29491 DVDD.n5667 DVDD.n5665 0.00796988
R29492 DVDD.n5665 DVDD.n255 0.00796988
R29493 DVDD.n3618 DVDD.n2433 0.00795714
R29494 DVDD.n5527 DVDD.n25 0.00793546
R29495 DVDD.n4689 DVDD.n4654 0.00793546
R29496 DVDD.n2640 DVDD.n2445 0.00783696
R29497 DVDD DVDD.n2195 0.00782857
R29498 DVDD.n2199 DVDD 0.00782857
R29499 DVDD DVDD.n3469 0.00782857
R29500 DVDD DVDD.n3468 0.00782857
R29501 DVDD.n1358 DVDD 0.00782857
R29502 DVDD.n1357 DVDD 0.00782857
R29503 DVDD.n3246 DVDD.n3245 0.0077973
R29504 DVDD.n3199 DVDD.n3125 0.0077973
R29505 DVDD.n5621 DVDD.n61 0.00778055
R29506 DVDD.n5446 DVDD.n304 0.00778055
R29507 DVDD.n2545 DVDD.n2544 0.00777531
R29508 DVDD.n2537 DVDD.n2530 0.00777531
R29509 DVDD.n2585 DVDD.n2527 0.00777531
R29510 DVDD.n2536 DVDD.n2526 0.00777531
R29511 DVDD.n2587 DVDD.n2533 0.00777531
R29512 DVDD.n2535 DVDD.n2525 0.00777531
R29513 DVDD.n2592 DVDD.n2534 0.00777531
R29514 DVDD.n2544 DVDD.n2528 0.00777531
R29515 DVDD.n2537 DVDD.n2528 0.00777531
R29516 DVDD.n2585 DVDD.n2530 0.00777531
R29517 DVDD.n2536 DVDD.n2532 0.00777531
R29518 DVDD.n2587 DVDD.n2526 0.00777531
R29519 DVDD.n2535 DVDD.n2533 0.00777531
R29520 DVDD.n2534 DVDD.n2525 0.00777531
R29521 DVDD.n2293 DVDD.n2123 0.00776429
R29522 DVDD.n1305 DVDD.n1301 0.00776429
R29523 DVDD.n1395 DVDD.n1394 0.00776429
R29524 DVDD.n5898 DVDD.n5897 0.00772462
R29525 DVDD.n5690 DVDD.n5689 0.00772462
R29526 DVDD.n5973 DVDD.n5972 0.00772462
R29527 DVDD.n5592 DVDD.n5591 0.00772462
R29528 DVDD.n2720 DVDD.n2719 0.00770384
R29529 DVDD.n2718 DVDD.n2702 0.00770384
R29530 DVDD.n2666 DVDD.n2494 0.0077
R29531 DVDD.n3832 DVDD.n1830 0.0077
R29532 DVDD.n3835 DVDD.n3833 0.0077
R29533 DVDD.n5544 DVDD.n14 0.00762565
R29534 DVDD.n4672 DVDD.n981 0.00762565
R29535 DVDD.n1937 DVDD.n1929 0.00760526
R29536 DVDD.n2532 DVDD.n2531 0.00754348
R29537 DVDD.n1385 DVDD.n1313 0.00751835
R29538 DVDD.n1322 DVDD.n1216 0.00751835
R29539 DVDD.n1323 DVDD.n1316 0.00751005
R29540 DVDD.n1325 DVDD.n1316 0.00751005
R29541 DVDD.n1389 DVDD.n1380 0.00751005
R29542 DVDD.n1389 DVDD.n1388 0.00751005
R29543 DVDD.n3709 DVDD.n1896 0.00748725
R29544 DVDD.n3764 DVDD.n1666 0.00748725
R29545 DVDD.n3765 DVDD.n1670 0.00748725
R29546 DVDD.n1928 DVDD.n1921 0.007475
R29547 DVDD.n3281 DVDD.n3280 0.00734783
R29548 DVDD.n2944 DVDD.n2943 0.00734783
R29549 DVDD.n2645 DVDD.n2644 0.00734783
R29550 DVDD.n5923 DVDD.n78 0.00731583
R29551 DVDD.n5554 DVDD.n19 0.00731583
R29552 DVDD.n5560 DVDD.n18 0.00731583
R29553 DVDD.n4662 DVDD.n4648 0.00731583
R29554 DVDD.n4647 DVDD.n4646 0.00731583
R29555 DVDD.n331 DVDD.n326 0.00731583
R29556 DVDD.n2655 DVDD.n2498 0.00725
R29557 DVDD.n3902 DVDD.n3868 0.00725
R29558 DVDD.n3871 DVDD.n3867 0.00725
R29559 DVDD.n1373 DVDD.n1372 0.00720213
R29560 DVDD.n1372 DVDD.n1326 0.00720213
R29561 DVDD.n1376 DVDD.n1375 0.00720213
R29562 DVDD.n1377 DVDD.n1376 0.00720213
R29563 DVDD.n3066 DVDD.n3065 0.00717969
R29564 DVDD.n1765 DVDD.n1724 0.0071375
R29565 DVDD.n2368 DVDD.n2059 0.00712143
R29566 DVDD.n1576 DVDD.n1197 0.00712143
R29567 DVDD.n1573 DVDD.n1572 0.00712143
R29568 DVDD.n1209 DVDD.n1192 0.00712143
R29569 DVDD.n2994 DVDD.n2993 0.0071
R29570 DVDD.n3382 DVDD.n2755 0.0071
R29571 DVDD.n3267 DVDD.n3266 0.0071
R29572 DVDD.n3403 DVDD.n3402 0.0071
R29573 DVDD.n2531 DVDD.n2527 0.00702174
R29574 DVDD.n5537 DVDD.n13 0.00700602
R29575 DVDD.n4679 DVDD.n980 0.00700602
R29576 DVDD.n1371 DVDD.n1195 0.00699624
R29577 DVDD.n2572 DVDD.n2551 0.00699429
R29578 DVDD.n2561 DVDD.n2553 0.00699429
R29579 DVDD.n2568 DVDD.n2550 0.00699429
R29580 DVDD.n2562 DVDD.n2532 0.00699429
R29581 DVDD.n2567 DVDD.n2549 0.00699429
R29582 DVDD.n2563 DVDD.n2554 0.00699429
R29583 DVDD.n2566 DVDD.n2548 0.00699429
R29584 DVDD.n2581 DVDD.n2555 0.00699429
R29585 DVDD.n2573 DVDD.n2572 0.00699429
R29586 DVDD.n2561 DVDD.n2551 0.00699429
R29587 DVDD.n2568 DVDD.n2553 0.00699429
R29588 DVDD.n2562 DVDD.n2550 0.00699429
R29589 DVDD.n2567 DVDD.n2532 0.00699429
R29590 DVDD.n2563 DVDD.n2549 0.00699429
R29591 DVDD.n2566 DVDD.n2554 0.00699429
R29592 DVDD.n2555 DVDD.n2548 0.00699429
R29593 DVDD.n2076 DVDD.n2075 0.00699286
R29594 DVDD.n2360 DVDD.n2063 0.00699286
R29595 DVDD.n3240 DVDD.n3088 0.00698649
R29596 DVDD.n3176 DVDD.n3142 0.00698649
R29597 DVDD.n4084 DVDD.n4083 0.0068
R29598 DVDD.n4046 DVDD.n4043 0.0068
R29599 DVDD.n3024 DVDD.n3023 0.00678
R29600 DVDD.n3356 DVDD.n2774 0.00678
R29601 DVDD.n3309 DVDD.n3308 0.00678
R29602 DVDD.n3438 DVDD.n2694 0.00678
R29603 DVDD.n5521 DVDD.n26 0.00669621
R29604 DVDD.n4695 DVDD.n4655 0.00669621
R29605 DVDD.n4101 DVDD.n4035 0.0066875
R29606 DVDD.n4102 DVDD.n1792 0.0066875
R29607 DVDD.n2203 DVDD.n2199 0.00667143
R29608 DVDD.n2838 DVDD.n2794 0.00661413
R29609 DVDD.n2899 DVDD.n2877 0.00661413
R29610 DVDD.n5502 DVDD.n103 0.00660465
R29611 DVDD.n5502 DVDD.n5501 0.00660465
R29612 DVDD.n2397 DVDD.n2396 0.00658571
R29613 DVDD.n2396 DVDD.n2395 0.00658571
R29614 DVDD.n2395 DVDD.n2044 0.00658571
R29615 DVDD.n2389 DVDD.n2044 0.00658571
R29616 DVDD.n2389 DVDD.n2388 0.00658571
R29617 DVDD.n2388 DVDD.n2387 0.00658571
R29618 DVDD.n2387 DVDD.n2048 0.00658571
R29619 DVDD.n2381 DVDD.n2048 0.00658571
R29620 DVDD.n2381 DVDD.n2380 0.00658571
R29621 DVDD.n2380 DVDD.n2379 0.00658571
R29622 DVDD.n2379 DVDD.n2052 0.00658571
R29623 DVDD.n2373 DVDD.n2052 0.00658571
R29624 DVDD.n2373 DVDD.n2372 0.00658571
R29625 DVDD.n2372 DVDD.n2371 0.00658571
R29626 DVDD.n2371 DVDD.n2056 0.00658571
R29627 DVDD.n2070 DVDD.n2056 0.00658571
R29628 DVDD.n2078 DVDD.n2070 0.00658571
R29629 DVDD.n2079 DVDD.n2078 0.00658571
R29630 DVDD.n2080 DVDD.n2079 0.00658571
R29631 DVDD.n2080 DVDD.n2066 0.00658571
R29632 DVDD.n2089 DVDD.n2066 0.00658571
R29633 DVDD.n2090 DVDD.n2089 0.00658571
R29634 DVDD.n2358 DVDD.n2090 0.00658571
R29635 DVDD.n2358 DVDD.n2357 0.00658571
R29636 DVDD.n2357 DVDD.n2356 0.00658571
R29637 DVDD.n2356 DVDD.n2091 0.00658571
R29638 DVDD.n2350 DVDD.n2091 0.00658571
R29639 DVDD.n2350 DVDD.n2349 0.00658571
R29640 DVDD.n2349 DVDD.n2348 0.00658571
R29641 DVDD.n2348 DVDD.n2096 0.00658571
R29642 DVDD.n2103 DVDD.n2096 0.00658571
R29643 DVDD.n2331 DVDD.n2103 0.00658571
R29644 DVDD.n2331 DVDD.n2330 0.00658571
R29645 DVDD.n2330 DVDD.n2329 0.00658571
R29646 DVDD.n2329 DVDD.n2104 0.00658571
R29647 DVDD.n2323 DVDD.n2104 0.00658571
R29648 DVDD.n2323 DVDD.n2322 0.00658571
R29649 DVDD.n2322 DVDD.n2321 0.00658571
R29650 DVDD.n2321 DVDD.n2108 0.00658571
R29651 DVDD.n2315 DVDD.n2108 0.00658571
R29652 DVDD.n2315 DVDD.n2314 0.00658571
R29653 DVDD.n2314 DVDD.n2313 0.00658571
R29654 DVDD.n2313 DVDD.n2112 0.00658571
R29655 DVDD.n2307 DVDD.n2112 0.00658571
R29656 DVDD.n2307 DVDD.n2306 0.00658571
R29657 DVDD.n2306 DVDD.n2305 0.00658571
R29658 DVDD.n2305 DVDD.n2116 0.00658571
R29659 DVDD.n2299 DVDD.n2116 0.00658571
R29660 DVDD.n2299 DVDD.n2298 0.00658571
R29661 DVDD.n2298 DVDD.n2297 0.00658571
R29662 DVDD.n2297 DVDD.n2120 0.00658571
R29663 DVDD.n2135 DVDD.n2120 0.00658571
R29664 DVDD.n2135 DVDD.n2134 0.00658571
R29665 DVDD.n2144 DVDD.n2134 0.00658571
R29666 DVDD.n2145 DVDD.n2144 0.00658571
R29667 DVDD.n2146 DVDD.n2145 0.00658571
R29668 DVDD.n2146 DVDD.n2130 0.00658571
R29669 DVDD.n2155 DVDD.n2130 0.00658571
R29670 DVDD.n2156 DVDD.n2155 0.00658571
R29671 DVDD.n2283 DVDD.n2156 0.00658571
R29672 DVDD.n2283 DVDD.n2282 0.00658571
R29673 DVDD.n2282 DVDD.n2281 0.00658571
R29674 DVDD.n2281 DVDD.n2157 0.00658571
R29675 DVDD.n2275 DVDD.n2157 0.00658571
R29676 DVDD.n2275 DVDD.n2274 0.00658571
R29677 DVDD.n2274 DVDD.n2273 0.00658571
R29678 DVDD.n2273 DVDD.n2162 0.00658571
R29679 DVDD.n2169 DVDD.n2162 0.00658571
R29680 DVDD.n2256 DVDD.n2169 0.00658571
R29681 DVDD.n2256 DVDD.n2255 0.00658571
R29682 DVDD.n2255 DVDD.n2254 0.00658571
R29683 DVDD.n2254 DVDD.n2170 0.00658571
R29684 DVDD.n2248 DVDD.n2170 0.00658571
R29685 DVDD.n2248 DVDD.n2247 0.00658571
R29686 DVDD.n2247 DVDD.n2246 0.00658571
R29687 DVDD.n2246 DVDD.n2174 0.00658571
R29688 DVDD.n2240 DVDD.n2174 0.00658571
R29689 DVDD.n2240 DVDD.n2239 0.00658571
R29690 DVDD.n2239 DVDD.n2238 0.00658571
R29691 DVDD.n2238 DVDD.n2178 0.00658571
R29692 DVDD.n2232 DVDD.n2178 0.00658571
R29693 DVDD.n2232 DVDD.n2231 0.00658571
R29694 DVDD.n2231 DVDD.n2230 0.00658571
R29695 DVDD.n2230 DVDD.n2182 0.00658571
R29696 DVDD.n2224 DVDD.n2182 0.00658571
R29697 DVDD.n2224 DVDD.n2223 0.00658571
R29698 DVDD.n2223 DVDD.n2222 0.00658571
R29699 DVDD.n2222 DVDD.n2186 0.00658571
R29700 DVDD.n2216 DVDD.n2186 0.00658571
R29701 DVDD.n2216 DVDD.n2215 0.00658571
R29702 DVDD.n2215 DVDD.n2214 0.00658571
R29703 DVDD.n2214 DVDD.n2190 0.00658571
R29704 DVDD.n2208 DVDD.n2190 0.00658571
R29705 DVDD.n2208 DVDD.n2207 0.00658571
R29706 DVDD.n2207 DVDD.n2206 0.00658571
R29707 DVDD.n2206 DVDD.n2194 0.00658571
R29708 DVDD.n2196 DVDD.n2194 0.00658571
R29709 DVDD.n3664 DVDD.n3663 0.00658571
R29710 DVDD.n3663 DVDD.n2407 0.00658571
R29711 DVDD.n2411 DVDD.n2407 0.00658571
R29712 DVDD.n3656 DVDD.n2411 0.00658571
R29713 DVDD.n3656 DVDD.n3655 0.00658571
R29714 DVDD.n3655 DVDD.n3654 0.00658571
R29715 DVDD.n3654 DVDD.n2412 0.00658571
R29716 DVDD.n3648 DVDD.n2412 0.00658571
R29717 DVDD.n3648 DVDD.n3647 0.00658571
R29718 DVDD.n3647 DVDD.n3646 0.00658571
R29719 DVDD.n3646 DVDD.n2416 0.00658571
R29720 DVDD.n3640 DVDD.n2416 0.00658571
R29721 DVDD.n3640 DVDD.n3639 0.00658571
R29722 DVDD.n3639 DVDD.n3638 0.00658571
R29723 DVDD.n3638 DVDD.n2420 0.00658571
R29724 DVDD.n3632 DVDD.n2420 0.00658571
R29725 DVDD.n3632 DVDD.n3631 0.00658571
R29726 DVDD.n3631 DVDD.n3630 0.00658571
R29727 DVDD.n3630 DVDD.n2424 0.00658571
R29728 DVDD.n3624 DVDD.n2424 0.00658571
R29729 DVDD.n3624 DVDD.n3623 0.00658571
R29730 DVDD.n3623 DVDD.n3622 0.00658571
R29731 DVDD.n3622 DVDD.n2428 0.00658571
R29732 DVDD.n3616 DVDD.n2428 0.00658571
R29733 DVDD.n3616 DVDD.n3615 0.00658571
R29734 DVDD.n3615 DVDD.n3614 0.00658571
R29735 DVDD.n3614 DVDD.n2435 0.00658571
R29736 DVDD.n3608 DVDD.n2435 0.00658571
R29737 DVDD.n3608 DVDD.n3607 0.00658571
R29738 DVDD.n3607 DVDD.n3606 0.00658571
R29739 DVDD.n3606 DVDD.n2440 0.00658571
R29740 DVDD.n3598 DVDD.n2440 0.00658571
R29741 DVDD.n3598 DVDD.n3597 0.00658571
R29742 DVDD.n3597 DVDD.n3596 0.00658571
R29743 DVDD.n3596 DVDD.n2457 0.00658571
R29744 DVDD.n3590 DVDD.n2457 0.00658571
R29745 DVDD.n3590 DVDD.n3589 0.00658571
R29746 DVDD.n3589 DVDD.n3588 0.00658571
R29747 DVDD.n3588 DVDD.n2461 0.00658571
R29748 DVDD.n3582 DVDD.n2461 0.00658571
R29749 DVDD.n3582 DVDD.n3581 0.00658571
R29750 DVDD.n3581 DVDD.n3580 0.00658571
R29751 DVDD.n3580 DVDD.n2465 0.00658571
R29752 DVDD.n3574 DVDD.n2465 0.00658571
R29753 DVDD.n3574 DVDD.n3573 0.00658571
R29754 DVDD.n3573 DVDD.n3572 0.00658571
R29755 DVDD.n3572 DVDD.n2469 0.00658571
R29756 DVDD.n3566 DVDD.n2469 0.00658571
R29757 DVDD.n3566 DVDD.n3565 0.00658571
R29758 DVDD.n3565 DVDD.n3564 0.00658571
R29759 DVDD.n3564 DVDD.n2473 0.00658571
R29760 DVDD.n3558 DVDD.n2473 0.00658571
R29761 DVDD.n3558 DVDD.n3557 0.00658571
R29762 DVDD.n3557 DVDD.n3556 0.00658571
R29763 DVDD.n3556 DVDD.n2477 0.00658571
R29764 DVDD.n3550 DVDD.n2477 0.00658571
R29765 DVDD.n3550 DVDD.n3549 0.00658571
R29766 DVDD.n3549 DVDD.n3548 0.00658571
R29767 DVDD.n3548 DVDD.n2481 0.00658571
R29768 DVDD.n3542 DVDD.n2481 0.00658571
R29769 DVDD.n3542 DVDD.n3541 0.00658571
R29770 DVDD.n3541 DVDD.n3540 0.00658571
R29771 DVDD.n3540 DVDD.n2485 0.00658571
R29772 DVDD.n3534 DVDD.n2485 0.00658571
R29773 DVDD.n3534 DVDD.n3533 0.00658571
R29774 DVDD.n3533 DVDD.n3532 0.00658571
R29775 DVDD.n3532 DVDD.n2489 0.00658571
R29776 DVDD.n2674 DVDD.n2489 0.00658571
R29777 DVDD.n2677 DVDD.n2674 0.00658571
R29778 DVDD.n2678 DVDD.n2677 0.00658571
R29779 DVDD.n3522 DVDD.n2678 0.00658571
R29780 DVDD.n3522 DVDD.n3521 0.00658571
R29781 DVDD.n3521 DVDD.n3520 0.00658571
R29782 DVDD.n3520 DVDD.n2679 0.00658571
R29783 DVDD.n3514 DVDD.n2679 0.00658571
R29784 DVDD.n3514 DVDD.n3513 0.00658571
R29785 DVDD.n3513 DVDD.n3512 0.00658571
R29786 DVDD.n3512 DVDD.n2683 0.00658571
R29787 DVDD.n3506 DVDD.n2683 0.00658571
R29788 DVDD.n3506 DVDD.n3505 0.00658571
R29789 DVDD.n3505 DVDD.n3504 0.00658571
R29790 DVDD.n3504 DVDD.n3454 0.00658571
R29791 DVDD.n3498 DVDD.n3454 0.00658571
R29792 DVDD.n3498 DVDD.n3497 0.00658571
R29793 DVDD.n3497 DVDD.n3496 0.00658571
R29794 DVDD.n3496 DVDD.n3458 0.00658571
R29795 DVDD.n3490 DVDD.n3458 0.00658571
R29796 DVDD.n3490 DVDD.n3489 0.00658571
R29797 DVDD.n3489 DVDD.n3488 0.00658571
R29798 DVDD.n3488 DVDD.n3462 0.00658571
R29799 DVDD.n3482 DVDD.n3462 0.00658571
R29800 DVDD.n3482 DVDD.n3481 0.00658571
R29801 DVDD.n3481 DVDD.n3480 0.00658571
R29802 DVDD.n3480 DVDD.n3466 0.00658571
R29803 DVDD.n3474 DVDD.n3466 0.00658571
R29804 DVDD.n3474 DVDD.n3473 0.00658571
R29805 DVDD.n3473 DVDD.n3472 0.00658571
R29806 DVDD.n1570 DVDD.n1569 0.00658571
R29807 DVDD.n1569 DVDD.n1568 0.00658571
R29808 DVDD.n1568 DVDD.n1207 0.00658571
R29809 DVDD.n1562 DVDD.n1207 0.00658571
R29810 DVDD.n1562 DVDD.n1561 0.00658571
R29811 DVDD.n1561 DVDD.n1560 0.00658571
R29812 DVDD.n1560 DVDD.n1212 0.00658571
R29813 DVDD.n1226 DVDD.n1212 0.00658571
R29814 DVDD.n1551 DVDD.n1226 0.00658571
R29815 DVDD.n1551 DVDD.n1550 0.00658571
R29816 DVDD.n1550 DVDD.n1549 0.00658571
R29817 DVDD.n1549 DVDD.n1227 0.00658571
R29818 DVDD.n1543 DVDD.n1227 0.00658571
R29819 DVDD.n1543 DVDD.n1542 0.00658571
R29820 DVDD.n1542 DVDD.n1541 0.00658571
R29821 DVDD.n1541 DVDD.n1231 0.00658571
R29822 DVDD.n1535 DVDD.n1231 0.00658571
R29823 DVDD.n1535 DVDD.n1534 0.00658571
R29824 DVDD.n1534 DVDD.n1533 0.00658571
R29825 DVDD.n1533 DVDD.n1235 0.00658571
R29826 DVDD.n1527 DVDD.n1235 0.00658571
R29827 DVDD.n1527 DVDD.n1526 0.00658571
R29828 DVDD.n1526 DVDD.n1525 0.00658571
R29829 DVDD.n1525 DVDD.n1239 0.00658571
R29830 DVDD.n1519 DVDD.n1239 0.00658571
R29831 DVDD.n1519 DVDD.n1518 0.00658571
R29832 DVDD.n1518 DVDD.n1517 0.00658571
R29833 DVDD.n1517 DVDD.n1243 0.00658571
R29834 DVDD.n1511 DVDD.n1243 0.00658571
R29835 DVDD.n1511 DVDD.n1510 0.00658571
R29836 DVDD.n1510 DVDD.n1509 0.00658571
R29837 DVDD.n1509 DVDD.n1247 0.00658571
R29838 DVDD.n1503 DVDD.n1247 0.00658571
R29839 DVDD.n1503 DVDD.n1502 0.00658571
R29840 DVDD.n1502 DVDD.n1501 0.00658571
R29841 DVDD.n1501 DVDD.n1251 0.00658571
R29842 DVDD.n1495 DVDD.n1251 0.00658571
R29843 DVDD.n1495 DVDD.n1494 0.00658571
R29844 DVDD.n1494 DVDD.n1493 0.00658571
R29845 DVDD.n1493 DVDD.n1255 0.00658571
R29846 DVDD.n1487 DVDD.n1255 0.00658571
R29847 DVDD.n1487 DVDD.n1486 0.00658571
R29848 DVDD.n1486 DVDD.n1485 0.00658571
R29849 DVDD.n1485 DVDD.n1259 0.00658571
R29850 DVDD.n1479 DVDD.n1259 0.00658571
R29851 DVDD.n1479 DVDD.n1478 0.00658571
R29852 DVDD.n1478 DVDD.n1477 0.00658571
R29853 DVDD.n1477 DVDD.n1263 0.00658571
R29854 DVDD.n1471 DVDD.n1263 0.00658571
R29855 DVDD.n1471 DVDD.n1470 0.00658571
R29856 DVDD.n1470 DVDD.n1469 0.00658571
R29857 DVDD.n1469 DVDD.n1267 0.00658571
R29858 DVDD.n1463 DVDD.n1267 0.00658571
R29859 DVDD.n1463 DVDD.n1462 0.00658571
R29860 DVDD.n1462 DVDD.n1461 0.00658571
R29861 DVDD.n1461 DVDD.n1271 0.00658571
R29862 DVDD.n1455 DVDD.n1271 0.00658571
R29863 DVDD.n1455 DVDD.n1454 0.00658571
R29864 DVDD.n1454 DVDD.n1453 0.00658571
R29865 DVDD.n1453 DVDD.n1275 0.00658571
R29866 DVDD.n1447 DVDD.n1275 0.00658571
R29867 DVDD.n1447 DVDD.n1446 0.00658571
R29868 DVDD.n1446 DVDD.n1445 0.00658571
R29869 DVDD.n1445 DVDD.n1279 0.00658571
R29870 DVDD.n1439 DVDD.n1279 0.00658571
R29871 DVDD.n1439 DVDD.n1438 0.00658571
R29872 DVDD.n1438 DVDD.n1437 0.00658571
R29873 DVDD.n1437 DVDD.n1283 0.00658571
R29874 DVDD.n1431 DVDD.n1283 0.00658571
R29875 DVDD.n1431 DVDD.n1430 0.00658571
R29876 DVDD.n1430 DVDD.n1429 0.00658571
R29877 DVDD.n1429 DVDD.n1287 0.00658571
R29878 DVDD.n1423 DVDD.n1287 0.00658571
R29879 DVDD.n1423 DVDD.n1422 0.00658571
R29880 DVDD.n1422 DVDD.n1421 0.00658571
R29881 DVDD.n1421 DVDD.n1291 0.00658571
R29882 DVDD.n1415 DVDD.n1291 0.00658571
R29883 DVDD.n1415 DVDD.n1414 0.00658571
R29884 DVDD.n1414 DVDD.n1413 0.00658571
R29885 DVDD.n1413 DVDD.n1295 0.00658571
R29886 DVDD.n1407 DVDD.n1295 0.00658571
R29887 DVDD.n1407 DVDD.n1406 0.00658571
R29888 DVDD.n1406 DVDD.n1405 0.00658571
R29889 DVDD.n1405 DVDD.n1299 0.00658571
R29890 DVDD.n1399 DVDD.n1299 0.00658571
R29891 DVDD.n1399 DVDD.n1398 0.00658571
R29892 DVDD.n1398 DVDD.n1397 0.00658571
R29893 DVDD.n1397 DVDD.n1303 0.00658571
R29894 DVDD.n1346 DVDD.n1303 0.00658571
R29895 DVDD.n1351 DVDD.n1346 0.00658571
R29896 DVDD.n1352 DVDD.n1351 0.00658571
R29897 DVDD.n1353 DVDD.n1352 0.00658571
R29898 DVDD.n1353 DVDD.n1342 0.00658571
R29899 DVDD.n1359 DVDD.n1342 0.00658571
R29900 DVDD.n1360 DVDD.n1359 0.00658571
R29901 DVDD.n5512 DVDD.n218 0.00654131
R29902 DVDD.n4707 DVDD.n4706 0.00654131
R29903 DVDD.n4880 DVDD.n703 0.0065
R29904 DVDD.n571 DVDD.n450 0.0065
R29905 DVDD.n909 DVDD.n359 0.0065
R29906 DVDD.n4881 DVDD.n4880 0.0065
R29907 DVDD.n990 DVDD.n358 0.0065
R29908 DVDD.n696 DVDD.n407 0.0065
R29909 DVDD.n4637 DVDD.n990 0.0065
R29910 DVDD.n4873 DVDD.n696 0.0065
R29911 DVDD.n5247 DVDD.n481 0.0065
R29912 DVDD.n4873 DVDD.n4804 0.0065
R29913 DVDD.n4637 DVDD.n908 0.0065
R29914 DVDD.n5712 DVDD.n38 0.0065
R29915 DVDD.n44 DVDD.n38 0.0065
R29916 DVDD.n5248 DVDD.n5247 0.0065
R29917 DVDD.n5248 DVDD.n448 0.0065
R29918 DVDD.n119 DVDD.n44 0.0065
R29919 DVDD.n5401 DVDD.n359 0.0065
R29920 DVDD.n4881 DVDD.n405 0.0065
R29921 DVDD.n5939 DVDD.n41 0.0065
R29922 DVDD.n5321 DVDD.n450 0.0065
R29923 DVDD.n5322 DVDD.n5321 0.0065
R29924 DVDD.n5940 DVDD.n40 0.0065
R29925 DVDD.n5940 DVDD.n5939 0.0065
R29926 DVDD.n4720 DVDD.n909 0.0065
R29927 DVDD.n4199 DVDD.n4198 0.00642084
R29928 DVDD.n71 DVDD.n69 0.0063864
R29929 DVDD.n5436 DVDD.n285 0.0063864
R29930 DVDD.n2632 DVDD.n2449 0.00636957
R29931 DVDD.n2142 DVDD.n2141 0.00635
R29932 DVDD.n2286 DVDD.n2285 0.00635
R29933 DVDD.n2285 DVDD.n2127 0.00635
R29934 DVDD.n1741 DVDD.n1738 0.00635
R29935 DVDD.n1744 DVDD.n1743 0.00635
R29936 DVDD.n1391 DVDD.n1389 0.00635
R29937 DVDD.n1316 DVDD.n1315 0.00635
R29938 DVDD.n3923 DVDD.n1818 0.0062375
R29939 DVDD.n3977 DVDD.n3924 0.0062375
R29940 DVDD.n84 DVDD.n78 0.0062315
R29941 DVDD.n331 DVDD.n329 0.0062315
R29942 DVDD.n5627 DVDD.n5573 0.00607659
R29943 DVDD.n5452 DVDD.n280 0.00607659
R29944 DVDD.n5831 DVDD.n146 0.00603279
R29945 DVDD.n5187 DVDD.n455 0.00603279
R29946 DVDD.n4955 DVDD.n678 0.00603279
R29947 DVDD.n812 DVDD.n811 0.00603279
R29948 DVDD.n4511 DVDD.n1079 0.00603279
R29949 DVDD.n4069 DVDD.n4054 0.0060125
R29950 DVDD.n4068 DVDD.n4055 0.0060125
R29951 DVDD.n4065 DVDD.n4064 0.0060125
R29952 DVDD.n4059 DVDD.n4057 0.0060125
R29953 DVDD.n4058 DVDD.n1721 0.0060125
R29954 DVDD.n4227 DVDD.n4226 0.0060125
R29955 DVDD.n1764 DVDD.n1728 0.0060125
R29956 DVDD.n1763 DVDD.n1729 0.0060125
R29957 DVDD.n1760 DVDD.n1759 0.0060125
R29958 DVDD.n1734 DVDD.n1730 0.0060125
R29959 DVDD.n3277 DVDD.n3276 0.00588043
R29960 DVDD.n3334 DVDD.n3332 0.00588043
R29961 DVDD.n3331 DVDD.n2873 0.00588043
R29962 DVDD.n2815 DVDD.n2790 0.00588043
R29963 DVDD.n2941 DVDD.n2937 0.00588043
R29964 DVDD.n2818 DVDD.n2816 0.00588043
R29965 DVDD.n2719 DVDD 0.00587887
R29966 DVDD.n2718 DVDD 0.00587887
R29967 DVDD.n1679 DVDD.n1675 0.00584375
R29968 DVDD.n4268 DVDD.n1680 0.00584375
R29969 DVDD.n4267 DVDD.n1681 0.00584375
R29970 DVDD.n4264 DVDD.n4263 0.00584375
R29971 DVDD.n3812 DVDD.n1843 0.00584375
R29972 DVDD.n3814 DVDD.n3813 0.00584375
R29973 DVDD.n3819 DVDD.n1840 0.00584375
R29974 DVDD.n3818 DVDD.n1841 0.00584375
R29975 DVDD.n3825 DVDD.n1836 0.00584375
R29976 DVDD.n2345 DVDD.n2344 0.00583571
R29977 DVDD.n4080 DVDD.n4047 0.005825
R29978 DVDD.n4051 DVDD.n4047 0.005825
R29979 DVDD.n4073 DVDD.n4051 0.005825
R29980 DVDD.n4073 DVDD.n4072 0.005825
R29981 DVDD.n4072 DVDD.n4071 0.005825
R29982 DVDD.n4071 DVDD.n4052 0.005825
R29983 DVDD.n4062 DVDD.n4052 0.005825
R29984 DVDD.n4062 DVDD.n4061 0.005825
R29985 DVDD.n4061 DVDD.n1725 0.005825
R29986 DVDD.n4224 DVDD.n1725 0.005825
R29987 DVDD.n1766 DVDD.n1726 0.005825
R29988 DVDD.n1757 DVDD.n1726 0.005825
R29989 DVDD.n1757 DVDD.n1756 0.005825
R29990 DVDD.n1756 DVDD.n1755 0.005825
R29991 DVDD.n1755 DVDD.n1732 0.005825
R29992 DVDD.n1749 DVDD.n1732 0.005825
R29993 DVDD.n1749 DVDD.n1748 0.005825
R29994 DVDD.n1748 DVDD.n1747 0.005825
R29995 DVDD.n1747 DVDD.n1737 0.005825
R29996 DVDD.n4286 DVDD.n1668 0.005825
R29997 DVDD.n4280 DVDD.n1668 0.005825
R29998 DVDD.n4280 DVDD.n4279 0.005825
R29999 DVDD.n4279 DVDD.n4278 0.005825
R30000 DVDD.n4278 DVDD.n1673 0.005825
R30001 DVDD.n4272 DVDD.n1673 0.005825
R30002 DVDD.n4272 DVDD.n4271 0.005825
R30003 DVDD.n4271 DVDD.n4270 0.005825
R30004 DVDD.n4270 DVDD.n1677 0.005825
R30005 DVDD.n4261 DVDD.n1677 0.005825
R30006 DVDD.n3810 DVDD.n1686 0.005825
R30007 DVDD.n3810 DVDD.n1838 0.005825
R30008 DVDD.n3821 DVDD.n1838 0.005825
R30009 DVDD.n3822 DVDD.n3821 0.005825
R30010 DVDD.n3823 DVDD.n3822 0.005825
R30011 DVDD.n3823 DVDD.n1834 0.005825
R30012 DVDD.n3829 DVDD.n1834 0.005825
R30013 DVDD.n3830 DVDD.n3829 0.005825
R30014 DVDD.n3831 DVDD.n3830 0.005825
R30015 DVDD.n3875 DVDD.n3869 0.005825
R30016 DVDD.n3896 DVDD.n3875 0.005825
R30017 DVDD.n3896 DVDD.n3895 0.005825
R30018 DVDD.n3895 DVDD.n3894 0.005825
R30019 DVDD.n3894 DVDD.n3876 0.005825
R30020 DVDD.n3888 DVDD.n3876 0.005825
R30021 DVDD.n3888 DVDD.n3887 0.005825
R30022 DVDD.n3887 DVDD.n3886 0.005825
R30023 DVDD.n3886 DVDD.n3880 0.005825
R30024 DVDD.n3880 DVDD.n1790 0.005825
R30025 DVDD.n4103 DVDD.n1791 0.005825
R30026 DVDD.n4097 DVDD.n1791 0.005825
R30027 DVDD.n4097 DVDD.n4096 0.005825
R30028 DVDD.n4096 DVDD.n4095 0.005825
R30029 DVDD.n4095 DVDD.n4038 0.005825
R30030 DVDD.n4089 DVDD.n4038 0.005825
R30031 DVDD.n4089 DVDD.n4088 0.005825
R30032 DVDD.n4088 DVDD.n4087 0.005825
R30033 DVDD.n4087 DVDD.n4042 0.005825
R30034 DVDD.n3839 DVDD.n3838 0.005825
R30035 DVDD.n3840 DVDD.n3839 0.005825
R30036 DVDD.n3840 DVDD.n1825 0.005825
R30037 DVDD.n3846 DVDD.n1825 0.005825
R30038 DVDD.n3847 DVDD.n3846 0.005825
R30039 DVDD.n3848 DVDD.n3847 0.005825
R30040 DVDD.n3848 DVDD.n1821 0.005825
R30041 DVDD.n3854 DVDD.n1821 0.005825
R30042 DVDD.n3855 DVDD.n3854 0.005825
R30043 DVDD.n3856 DVDD.n3855 0.005825
R30044 DVDD.n3922 DVDD.n3921 0.005825
R30045 DVDD.n3921 DVDD.n3920 0.005825
R30046 DVDD.n3920 DVDD.n3861 0.005825
R30047 DVDD.n3914 DVDD.n3861 0.005825
R30048 DVDD.n3914 DVDD.n3913 0.005825
R30049 DVDD.n3913 DVDD.n3912 0.005825
R30050 DVDD.n3912 DVDD.n3865 0.005825
R30051 DVDD.n3906 DVDD.n3865 0.005825
R30052 DVDD.n3906 DVDD.n3905 0.005825
R30053 DVDD.n3809 DVDD.n1685 0.0057875
R30054 DVDD.n3808 DVDD.n3807 0.0057875
R30055 DVDD.n5644 DVDD.n5610 0.00576678
R30056 DVDD.n5469 DVDD.n292 0.00576678
R30057 DVDD.n3707 DVDD.n1910 0.00571437
R30058 DVDD.n4288 DVDD.n4287 0.00571437
R30059 DVDD.n2361 DVDD.n2360 0.00570714
R30060 DVDD.n5745 DVDD.n187 0.00566393
R30061 DVDD.n5243 DVDD.n5242 0.00566393
R30062 DVDD.n5015 DVDD.n604 0.00566393
R30063 DVDD.n4878 DVDD.n727 0.00566393
R30064 DVDD.n4616 DVDD.n4615 0.00566393
R30065 DVDD.n2823 DVDD.n2787 0.00563587
R30066 DVDD.n2880 DVDD.n2863 0.00563587
R30067 DVDD.n5567 DVDD.n49 0.00561188
R30068 DVDD.n274 DVDD.n272 0.00561188
R30069 DVDD.n966 DVDD.n965 0.00559827
R30070 DVDD.n5506 DVDD.n5505 0.00558651
R30071 DVDD.n3691 DVDD.n1895 0.00550579
R30072 DVDD.n2399 DVDD.n2039 0.00548841
R30073 DVDD.n3666 DVDD.n3665 0.00548841
R30074 DVDD.n2717 DVDD.n2701 0.00530256
R30075 DVDD.n5636 DVDD.n64 0.00530207
R30076 DVDD.n225 DVDD.n221 0.00530207
R30077 DVDD.n962 DVDD.n947 0.00530207
R30078 DVDD.n5461 DVDD.n301 0.00530207
R30079 DVDD.n3831 DVDD.n1829 0.0053
R30080 DVDD.n5815 DVDD.n160 0.00529508
R30081 DVDD.n5171 DVDD.n471 0.00529508
R30082 DVDD.n4971 DVDD.n4949 0.00529508
R30083 DVDD.n793 DVDD.n747 0.00529508
R30084 DVDD.n4527 DVDD.n4507 0.00529508
R30085 DVDD.n2270 DVDD.n2269 0.00519286
R30086 DVDD.n3708 DVDD.n3707 0.00515817
R30087 DVDD.n4287 DVDD.n1667 0.00515817
R30088 DVDD.n5529 DVDD.n11 0.00514716
R30089 DVDD.n4687 DVDD.n978 0.00514716
R30090 DVDD.n2830 DVDD.n2786 0.00514674
R30091 DVDD.n2907 DVDD.n2864 0.00514674
R30092 DVDD.n3905 DVDD.n3904 0.005
R30093 DVDD.n5619 DVDD.n56 0.00499225
R30094 DVDD.n5444 DVDD.n310 0.00499225
R30095 DVDD.n2269 DVDD.n2165 0.00493571
R30096 DVDD.n5761 DVDD.n172 0.00492623
R30097 DVDD.n5226 DVDD.n489 0.00492623
R30098 DVDD.n643 DVDD.n608 0.00492623
R30099 DVDD.n850 DVDD.n708 0.00492623
R30100 DVDD.n4599 DVDD.n1013 0.00492623
R30101 DVDD.n4223 DVDD.n1766 0.004925
R30102 DVDD.n5913 DVDD.n99 0.00490722
R30103 DVDD.n109 DVDD.n95 0.00490722
R30104 DVDD.n5416 DVDD.n338 0.00490722
R30105 DVDD.n352 DVDD.n342 0.00490722
R30106 DVDD.n941 DVDD.n940 0.00490722
R30107 DVDD.n958 DVDD.n920 0.00490722
R30108 DVDD.n240 DVDD.n233 0.00490722
R30109 DVDD.n246 DVDD.n239 0.00490722
R30110 DVDD.n1944 DVDD.n1943 0.00489803
R30111 DVDD.n1968 DVDD.n1956 0.00489803
R30112 DVDD.n1950 DVDD.n1920 0.00488868
R30113 DVDD.n3701 DVDD.n3700 0.00488868
R30114 DVDD.n4680 DVDD.n4678 0.00486994
R30115 DVDD.n5539 DVDD.n5538 0.00485986
R30116 DVDD.n5546 DVDD.n21 0.00483735
R30117 DVDD.n4670 DVDD.n4650 0.00483735
R30118 DVDD.n1670 DVDD.n1665 0.00477578
R30119 DVDD.n4331 DVDD.n4330 0.00476
R30120 DVDD.n4330 DVDD.n4329 0.00476
R30121 DVDD.n4329 DVDD.n4328 0.00476
R30122 DVDD.n4328 DVDD.n4306 0.00476
R30123 DVDD.n4324 DVDD.n4306 0.00476
R30124 DVDD.n4324 DVDD.n4323 0.00476
R30125 DVDD.n4323 DVDD.n4322 0.00476
R30126 DVDD.n4322 DVDD.n4312 0.00476
R30127 DVDD.n4318 DVDD.n4312 0.00476
R30128 DVDD.n4318 DVDD.n4317 0.00476
R30129 DVDD.n4317 DVDD.n913 0.00476
R30130 DVDD.n4714 DVDD.n913 0.00476
R30131 DVDD.n4714 DVDD.n911 0.00476
R30132 DVDD.n4718 DVDD.n911 0.00476
R30133 DVDD.n4722 DVDD.n906 0.00476
R30134 DVDD.n4726 DVDD.n906 0.00476
R30135 DVDD.n4726 DVDD.n904 0.00476
R30136 DVDD.n4730 DVDD.n904 0.00476
R30137 DVDD.n4730 DVDD.n902 0.00476
R30138 DVDD.n4734 DVDD.n902 0.00476
R30139 DVDD.n4734 DVDD.n900 0.00476
R30140 DVDD.n4738 DVDD.n900 0.00476
R30141 DVDD.n4738 DVDD.n898 0.00476
R30142 DVDD.n4742 DVDD.n898 0.00476
R30143 DVDD.n4742 DVDD.n890 0.00476
R30144 DVDD.n4748 DVDD.n890 0.00476
R30145 DVDD.n4748 DVDD.n888 0.00476
R30146 DVDD.n4752 DVDD.n888 0.00476
R30147 DVDD.n4752 DVDD.n886 0.00476
R30148 DVDD.n4756 DVDD.n886 0.00476
R30149 DVDD.n4756 DVDD.n884 0.00476
R30150 DVDD.n4760 DVDD.n884 0.00476
R30151 DVDD.n4760 DVDD.n882 0.00476
R30152 DVDD.n4764 DVDD.n882 0.00476
R30153 DVDD.n4764 DVDD.n880 0.00476
R30154 DVDD.n4770 DVDD.n880 0.00476
R30155 DVDD.n4770 DVDD.n732 0.00476
R30156 DVDD.n4803 DVDD.n734 0.00476
R30157 DVDD.n4799 DVDD.n734 0.00476
R30158 DVDD.n4799 DVDD.n4798 0.00476
R30159 DVDD.n4798 DVDD.n4797 0.00476
R30160 DVDD.n4797 DVDD.n4781 0.00476
R30161 DVDD.n4793 DVDD.n4781 0.00476
R30162 DVDD.n4793 DVDD.n4792 0.00476
R30163 DVDD.n4792 DVDD.n4791 0.00476
R30164 DVDD.n4791 DVDD.n4788 0.00476
R30165 DVDD.n4788 DVDD.n587 0.00476
R30166 DVDD.n5024 DVDD.n587 0.00476
R30167 DVDD.n5024 DVDD.n585 0.00476
R30168 DVDD.n5028 DVDD.n585 0.00476
R30169 DVDD.n5028 DVDD.n583 0.00476
R30170 DVDD.n5032 DVDD.n583 0.00476
R30171 DVDD.n5032 DVDD.n581 0.00476
R30172 DVDD.n5036 DVDD.n581 0.00476
R30173 DVDD.n5036 DVDD.n579 0.00476
R30174 DVDD.n5040 DVDD.n579 0.00476
R30175 DVDD.n5040 DVDD.n577 0.00476
R30176 DVDD.n5044 DVDD.n577 0.00476
R30177 DVDD.n5044 DVDD.n575 0.00476
R30178 DVDD.n5048 DVDD.n575 0.00476
R30179 DVDD.n5086 DVDD.n5085 0.00476
R30180 DVDD.n5085 DVDD.n5053 0.00476
R30181 DVDD.n5081 DVDD.n5053 0.00476
R30182 DVDD.n5081 DVDD.n5080 0.00476
R30183 DVDD.n5080 DVDD.n5079 0.00476
R30184 DVDD.n5079 DVDD.n5059 0.00476
R30185 DVDD.n5075 DVDD.n5059 0.00476
R30186 DVDD.n5075 DVDD.n5074 0.00476
R30187 DVDD.n5074 DVDD.n5073 0.00476
R30188 DVDD.n5073 DVDD.n5065 0.00476
R30189 DVDD.n5069 DVDD.n5065 0.00476
R30190 DVDD.n5069 DVDD.n200 0.00476
R30191 DVDD.n5728 DVDD.n200 0.00476
R30192 DVDD.n5728 DVDD.n5727 0.00476
R30193 DVDD.n5727 DVDD.n5726 0.00476
R30194 DVDD.n5726 DVDD.n204 0.00476
R30195 DVDD.n5722 DVDD.n204 0.00476
R30196 DVDD.n5722 DVDD.n5721 0.00476
R30197 DVDD.n5721 DVDD.n5720 0.00476
R30198 DVDD.n5720 DVDD.n210 0.00476
R30199 DVDD.n5716 DVDD.n210 0.00476
R30200 DVDD.n5716 DVDD.n5715 0.00476
R30201 DVDD.n5715 DVDD.n5714 0.00476
R30202 DVDD.n5711 DVDD.n217 0.00476
R30203 DVDD.n5702 DVDD.n217 0.00476
R30204 DVDD.n5702 DVDD.n5701 0.00476
R30205 DVDD.n5701 DVDD.n5700 0.00476
R30206 DVDD.n5700 DVDD.n5699 0.00476
R30207 DVDD.n5699 DVDD.n5680 0.00476
R30208 DVDD.n5695 DVDD.n5680 0.00476
R30209 DVDD.n5695 DVDD.n5694 0.00476
R30210 DVDD.n5694 DVDD.n5693 0.00476
R30211 DVDD.n5693 DVDD.n5686 0.00476
R30212 DVDD.n4374 DVDD.n4373 0.00476
R30213 DVDD.n4373 DVDD.n4372 0.00476
R30214 DVDD.n4372 DVDD.n4371 0.00476
R30215 DVDD.n4371 DVDD.n4351 0.00476
R30216 DVDD.n4367 DVDD.n4351 0.00476
R30217 DVDD.n4367 DVDD.n4366 0.00476
R30218 DVDD.n4366 DVDD.n4365 0.00476
R30219 DVDD.n4365 DVDD.n4357 0.00476
R30220 DVDD.n4361 DVDD.n4357 0.00476
R30221 DVDD.n4361 DVDD.n985 0.00476
R30222 DVDD.n4644 DVDD.n985 0.00476
R30223 DVDD.n4644 DVDD.n4643 0.00476
R30224 DVDD.n4643 DVDD.n4641 0.00476
R30225 DVDD.n4641 DVDD.n4639 0.00476
R30226 DVDD.n4636 DVDD.n992 0.00476
R30227 DVDD.n4632 DVDD.n992 0.00476
R30228 DVDD.n4632 DVDD.n4631 0.00476
R30229 DVDD.n4631 DVDD.n4630 0.00476
R30230 DVDD.n4630 DVDD.n998 0.00476
R30231 DVDD.n4626 DVDD.n998 0.00476
R30232 DVDD.n4626 DVDD.n4625 0.00476
R30233 DVDD.n4625 DVDD.n4624 0.00476
R30234 DVDD.n4624 DVDD.n1004 0.00476
R30235 DVDD.n4620 DVDD.n1004 0.00476
R30236 DVDD.n4620 DVDD.n4619 0.00476
R30237 DVDD.n4619 DVDD.n1009 0.00476
R30238 DVDD.n1044 DVDD.n1009 0.00476
R30239 DVDD.n1044 DVDD.n1043 0.00476
R30240 DVDD.n1043 DVDD.n1042 0.00476
R30241 DVDD.n1042 DVDD.n1025 0.00476
R30242 DVDD.n1038 DVDD.n1025 0.00476
R30243 DVDD.n1038 DVDD.n1037 0.00476
R30244 DVDD.n1037 DVDD.n1036 0.00476
R30245 DVDD.n1036 DVDD.n1033 0.00476
R30246 DVDD.n1033 DVDD.n729 0.00476
R30247 DVDD.n4875 DVDD.n729 0.00476
R30248 DVDD.n4875 DVDD.n4874 0.00476
R30249 DVDD.n4872 DVDD.n4871 0.00476
R30250 DVDD.n4871 DVDD.n4807 0.00476
R30251 DVDD.n4867 DVDD.n4807 0.00476
R30252 DVDD.n4867 DVDD.n4866 0.00476
R30253 DVDD.n4866 DVDD.n4865 0.00476
R30254 DVDD.n4865 DVDD.n4813 0.00476
R30255 DVDD.n4861 DVDD.n4813 0.00476
R30256 DVDD.n4861 DVDD.n4860 0.00476
R30257 DVDD.n4860 DVDD.n4859 0.00476
R30258 DVDD.n4859 DVDD.n4856 0.00476
R30259 DVDD.n4856 DVDD.n4855 0.00476
R30260 DVDD.n4855 DVDD.n4854 0.00476
R30261 DVDD.n4854 DVDD.n4853 0.00476
R30262 DVDD.n4853 DVDD.n4823 0.00476
R30263 DVDD.n4849 DVDD.n4823 0.00476
R30264 DVDD.n4849 DVDD.n4848 0.00476
R30265 DVDD.n4848 DVDD.n4847 0.00476
R30266 DVDD.n4847 DVDD.n4829 0.00476
R30267 DVDD.n4843 DVDD.n4829 0.00476
R30268 DVDD.n4843 DVDD.n4842 0.00476
R30269 DVDD.n4842 DVDD.n4841 0.00476
R30270 DVDD.n4841 DVDD.n4837 0.00476
R30271 DVDD.n4837 DVDD.n482 0.00476
R30272 DVDD.n5246 DVDD.n484 0.00476
R30273 DVDD.n553 DVDD.n484 0.00476
R30274 DVDD.n553 DVDD.n552 0.00476
R30275 DVDD.n552 DVDD.n551 0.00476
R30276 DVDD.n551 DVDD.n501 0.00476
R30277 DVDD.n547 DVDD.n501 0.00476
R30278 DVDD.n547 DVDD.n546 0.00476
R30279 DVDD.n546 DVDD.n545 0.00476
R30280 DVDD.n545 DVDD.n507 0.00476
R30281 DVDD.n541 DVDD.n507 0.00476
R30282 DVDD.n541 DVDD.n540 0.00476
R30283 DVDD.n540 DVDD.n539 0.00476
R30284 DVDD.n539 DVDD.n538 0.00476
R30285 DVDD.n538 DVDD.n513 0.00476
R30286 DVDD.n534 DVDD.n513 0.00476
R30287 DVDD.n534 DVDD.n533 0.00476
R30288 DVDD.n533 DVDD.n532 0.00476
R30289 DVDD.n532 DVDD.n519 0.00476
R30290 DVDD.n528 DVDD.n519 0.00476
R30291 DVDD.n528 DVDD.n527 0.00476
R30292 DVDD.n527 DVDD.n526 0.00476
R30293 DVDD.n526 DVDD.n37 0.00476
R30294 DVDD.n5942 DVDD.n37 0.00476
R30295 DVDD.n5952 DVDD.n33 0.00476
R30296 DVDD.n5952 DVDD.n5951 0.00476
R30297 DVDD.n5951 DVDD.n5949 0.00476
R30298 DVDD.n5949 DVDD.n6 0.00476
R30299 DVDD.n5959 DVDD.n6 0.00476
R30300 DVDD.n5959 DVDD.n4 0.00476
R30301 DVDD.n5964 DVDD.n4 0.00476
R30302 DVDD.n5964 DVDD.n2 0.00476
R30303 DVDD.n5968 DVDD.n2 0.00476
R30304 DVDD.n5969 DVDD.n5968 0.00476
R30305 DVDD.n4411 DVDD.n1107 0.00476
R30306 DVDD.n4418 DVDD.n1107 0.00476
R30307 DVDD.n4418 DVDD.n1105 0.00476
R30308 DVDD.n4422 DVDD.n1105 0.00476
R30309 DVDD.n4422 DVDD.n1103 0.00476
R30310 DVDD.n4426 DVDD.n1103 0.00476
R30311 DVDD.n4426 DVDD.n1101 0.00476
R30312 DVDD.n4430 DVDD.n1101 0.00476
R30313 DVDD.n4430 DVDD.n1099 0.00476
R30314 DVDD.n4434 DVDD.n1099 0.00476
R30315 DVDD.n4434 DVDD.n1097 0.00476
R30316 DVDD.n4438 DVDD.n1097 0.00476
R30317 DVDD.n4439 DVDD.n4438 0.00476
R30318 DVDD.n4440 DVDD.n4439 0.00476
R30319 DVDD.n4447 DVDD.n4444 0.00476
R30320 DVDD.n4447 DVDD.n1093 0.00476
R30321 DVDD.n4451 DVDD.n1093 0.00476
R30322 DVDD.n4451 DVDD.n1091 0.00476
R30323 DVDD.n4455 DVDD.n1091 0.00476
R30324 DVDD.n4455 DVDD.n1089 0.00476
R30325 DVDD.n4459 DVDD.n1089 0.00476
R30326 DVDD.n4459 DVDD.n1087 0.00476
R30327 DVDD.n4463 DVDD.n1087 0.00476
R30328 DVDD.n4463 DVDD.n1085 0.00476
R30329 DVDD.n4498 DVDD.n1085 0.00476
R30330 DVDD.n4498 DVDD.n4497 0.00476
R30331 DVDD.n4497 DVDD.n4468 0.00476
R30332 DVDD.n4493 DVDD.n4468 0.00476
R30333 DVDD.n4493 DVDD.n4492 0.00476
R30334 DVDD.n4492 DVDD.n4491 0.00476
R30335 DVDD.n4491 DVDD.n4474 0.00476
R30336 DVDD.n4487 DVDD.n4474 0.00476
R30337 DVDD.n4487 DVDD.n4486 0.00476
R30338 DVDD.n4486 DVDD.n4485 0.00476
R30339 DVDD.n4485 DVDD.n4481 0.00476
R30340 DVDD.n4481 DVDD.n701 0.00476
R30341 DVDD.n4883 DVDD.n701 0.00476
R30342 DVDD.n4887 DVDD.n694 0.00476
R30343 DVDD.n4891 DVDD.n694 0.00476
R30344 DVDD.n4891 DVDD.n692 0.00476
R30345 DVDD.n4895 DVDD.n692 0.00476
R30346 DVDD.n4895 DVDD.n690 0.00476
R30347 DVDD.n4899 DVDD.n690 0.00476
R30348 DVDD.n4899 DVDD.n688 0.00476
R30349 DVDD.n4903 DVDD.n688 0.00476
R30350 DVDD.n4903 DVDD.n686 0.00476
R30351 DVDD.n4907 DVDD.n686 0.00476
R30352 DVDD.n4907 DVDD.n684 0.00476
R30353 DVDD.n4939 DVDD.n684 0.00476
R30354 DVDD.n4939 DVDD.n4938 0.00476
R30355 DVDD.n4938 DVDD.n4912 0.00476
R30356 DVDD.n4934 DVDD.n4912 0.00476
R30357 DVDD.n4934 DVDD.n4933 0.00476
R30358 DVDD.n4933 DVDD.n4932 0.00476
R30359 DVDD.n4932 DVDD.n4918 0.00476
R30360 DVDD.n4928 DVDD.n4918 0.00476
R30361 DVDD.n4928 DVDD.n4927 0.00476
R30362 DVDD.n4927 DVDD.n4926 0.00476
R30363 DVDD.n4926 DVDD.n480 0.00476
R30364 DVDD.n5249 DVDD.n480 0.00476
R30365 DVDD.n5316 DVDD.n476 0.00476
R30366 DVDD.n5316 DVDD.n5315 0.00476
R30367 DVDD.n5315 DVDD.n5314 0.00476
R30368 DVDD.n5314 DVDD.n5256 0.00476
R30369 DVDD.n5310 DVDD.n5256 0.00476
R30370 DVDD.n5310 DVDD.n5309 0.00476
R30371 DVDD.n5309 DVDD.n5308 0.00476
R30372 DVDD.n5308 DVDD.n5262 0.00476
R30373 DVDD.n5304 DVDD.n5262 0.00476
R30374 DVDD.n5304 DVDD.n5303 0.00476
R30375 DVDD.n5303 DVDD.n5302 0.00476
R30376 DVDD.n5302 DVDD.n5300 0.00476
R30377 DVDD.n5300 DVDD.n5299 0.00476
R30378 DVDD.n5299 DVDD.n5298 0.00476
R30379 DVDD.n5298 DVDD.n5271 0.00476
R30380 DVDD.n5294 DVDD.n5271 0.00476
R30381 DVDD.n5294 DVDD.n5293 0.00476
R30382 DVDD.n5293 DVDD.n5292 0.00476
R30383 DVDD.n5292 DVDD.n5277 0.00476
R30384 DVDD.n5288 DVDD.n5277 0.00476
R30385 DVDD.n5288 DVDD.n5287 0.00476
R30386 DVDD.n5287 DVDD.n5286 0.00476
R30387 DVDD.n5286 DVDD.n5284 0.00476
R30388 DVDD.n5937 DVDD.n5936 0.00476
R30389 DVDD.n5936 DVDD.n47 0.00476
R30390 DVDD.n5578 DVDD.n47 0.00476
R30391 DVDD.n5602 DVDD.n5578 0.00476
R30392 DVDD.n5602 DVDD.n5601 0.00476
R30393 DVDD.n5601 DVDD.n5600 0.00476
R30394 DVDD.n5600 DVDD.n5584 0.00476
R30395 DVDD.n5596 DVDD.n5584 0.00476
R30396 DVDD.n5596 DVDD.n5595 0.00476
R30397 DVDD.n5595 DVDD.n5594 0.00476
R30398 DVDD.n1180 DVDD.n1179 0.00476
R30399 DVDD.n1179 DVDD.n1178 0.00476
R30400 DVDD.n1178 DVDD.n1177 0.00476
R30401 DVDD.n1177 DVDD.n1154 0.00476
R30402 DVDD.n1173 DVDD.n1154 0.00476
R30403 DVDD.n1173 DVDD.n1172 0.00476
R30404 DVDD.n1172 DVDD.n1171 0.00476
R30405 DVDD.n1171 DVDD.n1160 0.00476
R30406 DVDD.n1167 DVDD.n1160 0.00476
R30407 DVDD.n1167 DVDD.n1166 0.00476
R30408 DVDD.n1166 DVDD.n354 0.00476
R30409 DVDD.n5406 DVDD.n354 0.00476
R30410 DVDD.n5406 DVDD.n5405 0.00476
R30411 DVDD.n5405 DVDD.n5403 0.00476
R30412 DVDD.n5399 DVDD.n5398 0.00476
R30413 DVDD.n5398 DVDD.n5397 0.00476
R30414 DVDD.n5397 DVDD.n364 0.00476
R30415 DVDD.n5393 DVDD.n364 0.00476
R30416 DVDD.n5393 DVDD.n5392 0.00476
R30417 DVDD.n5392 DVDD.n5391 0.00476
R30418 DVDD.n5391 DVDD.n370 0.00476
R30419 DVDD.n5387 DVDD.n370 0.00476
R30420 DVDD.n5387 DVDD.n5386 0.00476
R30421 DVDD.n5386 DVDD.n5385 0.00476
R30422 DVDD.n5385 DVDD.n376 0.00476
R30423 DVDD.n5379 DVDD.n376 0.00476
R30424 DVDD.n5379 DVDD.n5378 0.00476
R30425 DVDD.n5378 DVDD.n5377 0.00476
R30426 DVDD.n5377 DVDD.n387 0.00476
R30427 DVDD.n5373 DVDD.n387 0.00476
R30428 DVDD.n5373 DVDD.n5372 0.00476
R30429 DVDD.n5372 DVDD.n5371 0.00476
R30430 DVDD.n5371 DVDD.n393 0.00476
R30431 DVDD.n5367 DVDD.n393 0.00476
R30432 DVDD.n5367 DVDD.n5366 0.00476
R30433 DVDD.n5366 DVDD.n5365 0.00476
R30434 DVDD.n5365 DVDD.n399 0.00476
R30435 DVDD.n5359 DVDD.n5358 0.00476
R30436 DVDD.n5358 DVDD.n5357 0.00476
R30437 DVDD.n5357 DVDD.n411 0.00476
R30438 DVDD.n5353 DVDD.n411 0.00476
R30439 DVDD.n5353 DVDD.n5352 0.00476
R30440 DVDD.n5352 DVDD.n5351 0.00476
R30441 DVDD.n5351 DVDD.n417 0.00476
R30442 DVDD.n5347 DVDD.n417 0.00476
R30443 DVDD.n5347 DVDD.n5346 0.00476
R30444 DVDD.n5346 DVDD.n5345 0.00476
R30445 DVDD.n5345 DVDD.n423 0.00476
R30446 DVDD.n430 DVDD.n423 0.00476
R30447 DVDD.n5338 DVDD.n430 0.00476
R30448 DVDD.n5338 DVDD.n5337 0.00476
R30449 DVDD.n5337 DVDD.n5336 0.00476
R30450 DVDD.n5336 DVDD.n436 0.00476
R30451 DVDD.n5332 DVDD.n436 0.00476
R30452 DVDD.n5332 DVDD.n5331 0.00476
R30453 DVDD.n5331 DVDD.n5330 0.00476
R30454 DVDD.n5330 DVDD.n442 0.00476
R30455 DVDD.n5326 DVDD.n442 0.00476
R30456 DVDD.n5326 DVDD.n5325 0.00476
R30457 DVDD.n5325 DVDD.n5324 0.00476
R30458 DVDD.n5134 DVDD.n5108 0.00476
R30459 DVDD.n5134 DVDD.n5133 0.00476
R30460 DVDD.n5133 DVDD.n5132 0.00476
R30461 DVDD.n5132 DVDD.n5113 0.00476
R30462 DVDD.n5128 DVDD.n5113 0.00476
R30463 DVDD.n5128 DVDD.n5127 0.00476
R30464 DVDD.n5127 DVDD.n5126 0.00476
R30465 DVDD.n5126 DVDD.n5119 0.00476
R30466 DVDD.n5122 DVDD.n5119 0.00476
R30467 DVDD.n5122 DVDD.n133 0.00476
R30468 DVDD.n5853 DVDD.n133 0.00476
R30469 DVDD.n5853 DVDD.n131 0.00476
R30470 DVDD.n5857 DVDD.n131 0.00476
R30471 DVDD.n5857 DVDD.n129 0.00476
R30472 DVDD.n5861 DVDD.n129 0.00476
R30473 DVDD.n5861 DVDD.n127 0.00476
R30474 DVDD.n5865 DVDD.n127 0.00476
R30475 DVDD.n5865 DVDD.n125 0.00476
R30476 DVDD.n5869 DVDD.n125 0.00476
R30477 DVDD.n5869 DVDD.n123 0.00476
R30478 DVDD.n5873 DVDD.n123 0.00476
R30479 DVDD.n5873 DVDD.n121 0.00476
R30480 DVDD.n5877 DVDD.n121 0.00476
R30481 DVDD.n5882 DVDD.n5881 0.00476
R30482 DVDD.n5884 DVDD.n5882 0.00476
R30483 DVDD.n5884 DVDD.n117 0.00476
R30484 DVDD.n5908 DVDD.n117 0.00476
R30485 DVDD.n5908 DVDD.n5907 0.00476
R30486 DVDD.n5907 DVDD.n5906 0.00476
R30487 DVDD.n5906 DVDD.n5890 0.00476
R30488 DVDD.n5902 DVDD.n5890 0.00476
R30489 DVDD.n5902 DVDD.n5901 0.00476
R30490 DVDD.n5901 DVDD.n5900 0.00476
R30491 DVDD.n3436 DVDD.n2689 0.00476
R30492 DVDD.n3443 DVDD.n2690 0.00476
R30493 DVDD.n2690 DVDD.n1915 0.00476
R30494 DVDD.n1941 DVDD.n1914 0.00476
R30495 DVDD.n1941 DVDD.n1938 0.00476
R30496 DVDD.n2975 DVDD.n2968 0.00476
R30497 DVDD.n2979 DVDD.n2968 0.00476
R30498 DVDD.n2979 DVDD.n2969 0.00476
R30499 DVDD.n3392 DVDD.n2733 0.00476
R30500 DVDD.n3392 DVDD.n2728 0.00476
R30501 DVDD.n3400 DVDD.n2728 0.00476
R30502 DVDD.n3400 DVDD.n2726 0.00476
R30503 DVDD.n3404 DVDD.n2723 0.00476
R30504 DVDD.n3412 DVDD.n2723 0.00476
R30505 DVDD.n3412 DVDD.n2721 0.00476
R30506 DVDD.n3416 DVDD.n2721 0.00476
R30507 DVDD.n3425 DVDD.n2699 0.00476
R30508 DVDD.n3430 DVDD.n2699 0.00476
R30509 DVDD.n3430 DVDD.n2700 0.00476
R30510 DVDD.n2700 DVDD.n2695 0.00476
R30511 DVDD.n3437 DVDD.n2691 0.00476
R30512 DVDD.n3442 DVDD.n2691 0.00476
R30513 DVDD.n3442 DVDD.n2693 0.00476
R30514 DVDD.n2693 DVDD.n2692 0.00476
R30515 DVDD.n1942 DVDD.n1940 0.00476
R30516 DVDD.n1943 DVDD.n1942 0.00476
R30517 DVDD.n3104 DVDD.n3103 0.00476
R30518 DVDD.n3103 DVDD.n3102 0.00476
R30519 DVDD.n3102 DVDD.n3101 0.00476
R30520 DVDD.n3259 DVDD.n3257 0.00476
R30521 DVDD.n3259 DVDD.n2961 0.00476
R30522 DVDD.n3264 DVDD.n2961 0.00476
R30523 DVDD.n3264 DVDD.n2959 0.00476
R30524 DVDD.n3268 DVDD.n2930 0.00476
R30525 DVDD.n3284 DVDD.n2930 0.00476
R30526 DVDD.n3284 DVDD.n2928 0.00476
R30527 DVDD.n3288 DVDD.n2928 0.00476
R30528 DVDD.n3304 DVDD.n2922 0.00476
R30529 DVDD.n3304 DVDD.n2920 0.00476
R30530 DVDD.n3322 DVDD.n2920 0.00476
R30531 DVDD.n3322 DVDD.n3321 0.00476
R30532 DVDD.n3319 DVDD.n3318 0.00476
R30533 DVDD.n3318 DVDD.n3317 0.00476
R30534 DVDD.n3317 DVDD.n3314 0.00476
R30535 DVDD.n3314 DVDD.n3313 0.00476
R30536 DVDD.n1952 DVDD.n1951 0.00476
R30537 DVDD.n1951 DVDD.n1950 0.00476
R30538 DVDD.n3261 DVDD.n3260 0.00476
R30539 DVDD.n3263 DVDD.n3261 0.00476
R30540 DVDD.n3263 DVDD.n3262 0.00476
R30541 DVDD.n3316 DVDD.n3315 0.00476
R30542 DVDD.n3315 DVDD.n1917 0.00476
R30543 DVDD.n1953 DVDD.n1918 0.00476
R30544 DVDD.n1949 DVDD.n1918 0.00476
R30545 DVDD.n2753 DVDD.n2752 0.00476
R30546 DVDD.n2756 DVDD.n2753 0.00476
R30547 DVDD.n2757 DVDD.n2756 0.00476
R30548 DVDD.n3350 DVDD.n3349 0.00476
R30549 DVDD.n3350 DVDD.n1973 0.00476
R30550 DVDD.n1972 DVDD.n1955 0.00476
R30551 DVDD.n1957 DVDD.n1955 0.00476
R30552 DVDD.n3160 DVDD.n3156 0.00476
R30553 DVDD.n3160 DVDD.n3159 0.00476
R30554 DVDD.n3159 DVDD.n3158 0.00476
R30555 DVDD.n3387 DVDD.n3386 0.00476
R30556 DVDD.n3386 DVDD.n3385 0.00476
R30557 DVDD.n3385 DVDD.n2754 0.00476
R30558 DVDD.n3381 DVDD.n2754 0.00476
R30559 DVDD.n3380 DVDD.n3379 0.00476
R30560 DVDD.n3379 DVDD.n2760 0.00476
R30561 DVDD.n3375 DVDD.n2760 0.00476
R30562 DVDD.n3375 DVDD.n3374 0.00476
R30563 DVDD.n3363 DVDD.n2771 0.00476
R30564 DVDD.n3363 DVDD.n2772 0.00476
R30565 DVDD.n3359 DVDD.n2772 0.00476
R30566 DVDD.n3359 DVDD.n3358 0.00476
R30567 DVDD.n3357 DVDD.n2778 0.00476
R30568 DVDD.n3353 DVDD.n2778 0.00476
R30569 DVDD.n3353 DVDD.n3352 0.00476
R30570 DVDD.n3352 DVDD.n3351 0.00476
R30571 DVDD.n1971 DVDD.n1970 0.00476
R30572 DVDD.n1970 DVDD.n1956 0.00476
R30573 DVDD.n3076 DVDD.n3075 0.00476
R30574 DVDD.n3075 DVDD.n3074 0.00476
R30575 DVDD.n3074 DVDD.n2990 0.00476
R30576 DVDD.n3070 DVDD.n2990 0.00476
R30577 DVDD.n3069 DVDD.n2995 0.00476
R30578 DVDD.n3058 DVDD.n2995 0.00476
R30579 DVDD.n3058 DVDD.n3057 0.00476
R30580 DVDD.n3057 DVDD.n3006 0.00476
R30581 DVDD.n3050 DVDD.n3049 0.00476
R30582 DVDD.n3049 DVDD.n3014 0.00476
R30583 DVDD.n3038 DVDD.n3014 0.00476
R30584 DVDD.n3038 DVDD.n3037 0.00476
R30585 DVDD.n3036 DVDD.n3025 0.00476
R30586 DVDD.n3032 DVDD.n3025 0.00476
R30587 DVDD.n3032 DVDD.n3031 0.00476
R30588 DVDD.n3031 DVDD.n3030 0.00476
R30589 DVDD.n3705 DVDD.n1913 0.00476
R30590 DVDD.n3701 DVDD.n1913 0.00476
R30591 DVDD.n3077 DVDD.n2987 0.00476
R30592 DVDD.n3073 DVDD.n2987 0.00476
R30593 DVDD.n3073 DVDD.n3072 0.00476
R30594 DVDD.n3072 DVDD.n3071 0.00476
R30595 DVDD.n3039 DVDD.n3020 0.00476
R30596 DVDD.n3035 DVDD.n3034 0.00476
R30597 DVDD.n3034 DVDD.n3033 0.00476
R30598 DVDD.n3033 DVDD.n3026 0.00476
R30599 DVDD.n3026 DVDD.n1974 0.00476
R30600 DVDD.n3704 DVDD.n3703 0.00476
R30601 DVDD.n3703 DVDD.n3702 0.00476
R30602 DVDD.n3735 DVDD.n3734 0.00476
R30603 DVDD.n3734 DVDD.n1855 0.00476
R30604 DVDD.n3783 DVDD.n1855 0.00476
R30605 DVDD.n3783 DVDD.n1853 0.00476
R30606 DVDD.n3787 DVDD.n1853 0.00476
R30607 DVDD.n3787 DVDD.n1851 0.00476
R30608 DVDD.n3791 DVDD.n1851 0.00476
R30609 DVDD.n3791 DVDD.n1849 0.00476
R30610 DVDD.n3795 DVDD.n1849 0.00476
R30611 DVDD.n3795 DVDD.n1847 0.00476
R30612 DVDD.n3800 DVDD.n1847 0.00476
R30613 DVDD.n3800 DVDD.n1845 0.00476
R30614 DVDD.n3804 DVDD.n1845 0.00476
R30615 DVDD.n3805 DVDD.n3804 0.00476
R30616 DVDD.n4258 DVDD.n1689 0.00476
R30617 DVDD.n4254 DVDD.n1689 0.00476
R30618 DVDD.n4254 DVDD.n4253 0.00476
R30619 DVDD.n4253 DVDD.n1694 0.00476
R30620 DVDD.n4249 DVDD.n1694 0.00476
R30621 DVDD.n4249 DVDD.n4248 0.00476
R30622 DVDD.n4248 DVDD.n1699 0.00476
R30623 DVDD.n4244 DVDD.n1699 0.00476
R30624 DVDD.n4244 DVDD.n4243 0.00476
R30625 DVDD.n4243 DVDD.n4242 0.00476
R30626 DVDD.n4242 DVDD.n1705 0.00476
R30627 DVDD.n3937 DVDD.n1705 0.00476
R30628 DVDD.n3958 DVDD.n3937 0.00476
R30629 DVDD.n3958 DVDD.n3957 0.00476
R30630 DVDD.n3957 DVDD.n3956 0.00476
R30631 DVDD.n3956 DVDD.n3943 0.00476
R30632 DVDD.n3951 DVDD.n3943 0.00476
R30633 DVDD.n3951 DVDD.n3950 0.00476
R30634 DVDD.n3950 DVDD.n3949 0.00476
R30635 DVDD.n3949 DVDD.n3928 0.00476
R30636 DVDD.n3971 DVDD.n3928 0.00476
R30637 DVDD.n3971 DVDD.n3926 0.00476
R30638 DVDD.n3975 DVDD.n3926 0.00476
R30639 DVDD.n3979 DVDD.n1816 0.00476
R30640 DVDD.n3983 DVDD.n1816 0.00476
R30641 DVDD.n3983 DVDD.n1814 0.00476
R30642 DVDD.n3987 DVDD.n1814 0.00476
R30643 DVDD.n3987 DVDD.n1812 0.00476
R30644 DVDD.n3991 DVDD.n1812 0.00476
R30645 DVDD.n3991 DVDD.n1810 0.00476
R30646 DVDD.n3999 DVDD.n1810 0.00476
R30647 DVDD.n3999 DVDD.n1808 0.00476
R30648 DVDD.n4003 DVDD.n1808 0.00476
R30649 DVDD.n4003 DVDD.n1806 0.00476
R30650 DVDD.n4007 DVDD.n1806 0.00476
R30651 DVDD.n4007 DVDD.n1804 0.00476
R30652 DVDD.n4011 DVDD.n1804 0.00476
R30653 DVDD.n4011 DVDD.n1802 0.00476
R30654 DVDD.n4019 DVDD.n1802 0.00476
R30655 DVDD.n4019 DVDD.n1800 0.00476
R30656 DVDD.n4023 DVDD.n1800 0.00476
R30657 DVDD.n4023 DVDD.n1798 0.00476
R30658 DVDD.n4028 DVDD.n1798 0.00476
R30659 DVDD.n4028 DVDD.n1796 0.00476
R30660 DVDD.n4032 DVDD.n1796 0.00476
R30661 DVDD.n4033 DVDD.n4032 0.00476
R30662 DVDD.n4119 DVDD.n1788 0.00476
R30663 DVDD.n4119 DVDD.n4118 0.00476
R30664 DVDD.n4118 DVDD.n4117 0.00476
R30665 DVDD.n4117 DVDD.n4109 0.00476
R30666 DVDD.n4112 DVDD.n4109 0.00476
R30667 DVDD.n4112 DVDD.n1783 0.00476
R30668 DVDD.n4131 DVDD.n1783 0.00476
R30669 DVDD.n4131 DVDD.n1781 0.00476
R30670 DVDD.n4135 DVDD.n1781 0.00476
R30671 DVDD.n4135 DVDD.n1779 0.00476
R30672 DVDD.n4143 DVDD.n1779 0.00476
R30673 DVDD.n4143 DVDD.n1777 0.00476
R30674 DVDD.n4147 DVDD.n1777 0.00476
R30675 DVDD.n4147 DVDD.n1776 0.00476
R30676 DVDD.n4153 DVDD.n1776 0.00476
R30677 DVDD.n4153 DVDD.n1774 0.00476
R30678 DVDD.n4157 DVDD.n1774 0.00476
R30679 DVDD.n4157 DVDD.n1772 0.00476
R30680 DVDD.n4163 DVDD.n1772 0.00476
R30681 DVDD.n4163 DVDD.n1770 0.00476
R30682 DVDD.n4167 DVDD.n1770 0.00476
R30683 DVDD.n4167 DVDD.n1768 0.00476
R30684 DVDD.n4171 DVDD.n1768 0.00476
R30685 DVDD.n4221 DVDD.n4174 0.00476
R30686 DVDD.n4217 DVDD.n4174 0.00476
R30687 DVDD.n4217 DVDD.n4216 0.00476
R30688 DVDD.n4216 DVDD.n4215 0.00476
R30689 DVDD.n4215 DVDD.n4182 0.00476
R30690 DVDD.n4211 DVDD.n4182 0.00476
R30691 DVDD.n4211 DVDD.n4210 0.00476
R30692 DVDD.n4210 DVDD.n4209 0.00476
R30693 DVDD.n4209 DVDD.n4188 0.00476
R30694 DVDD.n4193 DVDD.n4188 0.00476
R30695 DVDD.n4198 DVDD.n4197 0.00476
R30696 DVDD.n3782 DVDD.n3780 0.00476
R30697 DVDD.n3782 DVDD.n3781 0.00476
R30698 DVDD.n3789 DVDD.n3788 0.00476
R30699 DVDD.n3790 DVDD.n3789 0.00476
R30700 DVDD.n3790 DVDD.n1848 0.00476
R30701 DVDD.n3796 DVDD.n1848 0.00476
R30702 DVDD.n3797 DVDD.n3796 0.00476
R30703 DVDD.n3799 DVDD.n3797 0.00476
R30704 DVDD.n3799 DVDD.n3798 0.00476
R30705 DVDD.n3798 DVDD.n1844 0.00476
R30706 DVDD.n3806 DVDD.n1844 0.00476
R30707 DVDD.n4257 DVDD.n4256 0.00476
R30708 DVDD.n4256 DVDD.n4255 0.00476
R30709 DVDD.n4252 DVDD.n4251 0.00476
R30710 DVDD.n4251 DVDD.n4250 0.00476
R30711 DVDD.n4247 DVDD.n4246 0.00476
R30712 DVDD.n4246 DVDD.n4245 0.00476
R30713 DVDD.n4245 DVDD.n1700 0.00476
R30714 DVDD.n3935 DVDD.n1707 0.00476
R30715 DVDD.n3959 DVDD.n3936 0.00476
R30716 DVDD.n3955 DVDD.n3936 0.00476
R30717 DVDD.n3953 DVDD.n3952 0.00476
R30718 DVDD.n3952 DVDD.n3944 0.00476
R30719 DVDD.n3944 DVDD.n3929 0.00476
R30720 DVDD.n3970 DVDD.n3968 0.00476
R30721 DVDD.n3970 DVDD.n3969 0.00476
R30722 DVDD.n3978 DVDD.n1815 0.00476
R30723 DVDD.n3984 DVDD.n1815 0.00476
R30724 DVDD.n3985 DVDD.n3984 0.00476
R30725 DVDD.n3986 DVDD.n3985 0.00476
R30726 DVDD.n3986 DVDD.n1811 0.00476
R30727 DVDD.n3992 DVDD.n1811 0.00476
R30728 DVDD.n3993 DVDD.n3992 0.00476
R30729 DVDD.n3998 DVDD.n3993 0.00476
R30730 DVDD.n4004 DVDD.n1807 0.00476
R30731 DVDD.n4005 DVDD.n4004 0.00476
R30732 DVDD.n4006 DVDD.n4005 0.00476
R30733 DVDD.n4006 DVDD.n1803 0.00476
R30734 DVDD.n4012 DVDD.n1803 0.00476
R30735 DVDD.n4018 DVDD.n4017 0.00476
R30736 DVDD.n4018 DVDD.n1799 0.00476
R30737 DVDD.n4024 DVDD.n1799 0.00476
R30738 DVDD.n4025 DVDD.n4024 0.00476
R30739 DVDD.n4027 DVDD.n4025 0.00476
R30740 DVDD.n4027 DVDD.n4026 0.00476
R30741 DVDD.n4026 DVDD.n1795 0.00476
R30742 DVDD.n4034 DVDD.n1795 0.00476
R30743 DVDD.n4120 DVDD.n1787 0.00476
R30744 DVDD.n4116 DVDD.n1787 0.00476
R30745 DVDD.n4114 DVDD.n4113 0.00476
R30746 DVDD.n4113 DVDD.n1784 0.00476
R30747 DVDD.n4130 DVDD.n1784 0.00476
R30748 DVDD.n4136 DVDD.n1780 0.00476
R30749 DVDD.n4137 DVDD.n4136 0.00476
R30750 DVDD.n4142 DVDD.n4141 0.00476
R30751 DVDD.n4152 DVDD.n4151 0.00476
R30752 DVDD.n4152 DVDD.n1773 0.00476
R30753 DVDD.n4158 DVDD.n1773 0.00476
R30754 DVDD.n4162 DVDD.n4160 0.00476
R30755 DVDD.n4162 DVDD.n4161 0.00476
R30756 DVDD.n4169 DVDD.n4168 0.00476
R30757 DVDD.n4170 DVDD.n4169 0.00476
R30758 DVDD.n4220 DVDD.n4219 0.00476
R30759 DVDD.n4219 DVDD.n4218 0.00476
R30760 DVDD.n4218 DVDD.n4178 0.00476
R30761 DVDD.n4214 DVDD.n4178 0.00476
R30762 DVDD.n4214 DVDD.n4213 0.00476
R30763 DVDD.n4213 DVDD.n4212 0.00476
R30764 DVDD.n4212 DVDD.n4183 0.00476
R30765 DVDD.n4208 DVDD.n4183 0.00476
R30766 DVDD.n4208 DVDD.n4207 0.00476
R30767 DVDD.n4196 DVDD.n4191 0.00476
R30768 DVDD.n1176 DVDD.n1131 0.00476
R30769 DVDD.n1176 DVDD.n1175 0.00476
R30770 DVDD.n1175 DVDD.n1174 0.00476
R30771 DVDD.n1174 DVDD.n1155 0.00476
R30772 DVDD.n1170 DVDD.n1155 0.00476
R30773 DVDD.n1170 DVDD.n1169 0.00476
R30774 DVDD.n1169 DVDD.n1168 0.00476
R30775 DVDD.n1168 DVDD.n1161 0.00476
R30776 DVDD.n5400 DVDD.n360 0.00476
R30777 DVDD.n5396 DVDD.n360 0.00476
R30778 DVDD.n5396 DVDD.n5395 0.00476
R30779 DVDD.n5395 DVDD.n5394 0.00476
R30780 DVDD.n5394 DVDD.n365 0.00476
R30781 DVDD.n5390 DVDD.n365 0.00476
R30782 DVDD.n5390 DVDD.n5389 0.00476
R30783 DVDD.n5389 DVDD.n5388 0.00476
R30784 DVDD.n5388 DVDD.n371 0.00476
R30785 DVDD.n5384 DVDD.n371 0.00476
R30786 DVDD.n5380 DVDD.n382 0.00476
R30787 DVDD.n5376 DVDD.n382 0.00476
R30788 DVDD.n5376 DVDD.n5375 0.00476
R30789 DVDD.n5375 DVDD.n5374 0.00476
R30790 DVDD.n5374 DVDD.n388 0.00476
R30791 DVDD.n5370 DVDD.n388 0.00476
R30792 DVDD.n5370 DVDD.n5369 0.00476
R30793 DVDD.n5369 DVDD.n5368 0.00476
R30794 DVDD.n5368 DVDD.n394 0.00476
R30795 DVDD.n5364 DVDD.n394 0.00476
R30796 DVDD.n5360 DVDD.n406 0.00476
R30797 DVDD.n5356 DVDD.n406 0.00476
R30798 DVDD.n5356 DVDD.n5355 0.00476
R30799 DVDD.n5355 DVDD.n5354 0.00476
R30800 DVDD.n5354 DVDD.n412 0.00476
R30801 DVDD.n5350 DVDD.n412 0.00476
R30802 DVDD.n5350 DVDD.n5349 0.00476
R30803 DVDD.n5349 DVDD.n5348 0.00476
R30804 DVDD.n5348 DVDD.n418 0.00476
R30805 DVDD.n5344 DVDD.n418 0.00476
R30806 DVDD.n5344 DVDD.n5343 0.00476
R30807 DVDD.n5339 DVDD.n429 0.00476
R30808 DVDD.n5335 DVDD.n429 0.00476
R30809 DVDD.n5335 DVDD.n5334 0.00476
R30810 DVDD.n5334 DVDD.n5333 0.00476
R30811 DVDD.n5333 DVDD.n437 0.00476
R30812 DVDD.n5329 DVDD.n437 0.00476
R30813 DVDD.n5329 DVDD.n5328 0.00476
R30814 DVDD.n5328 DVDD.n5327 0.00476
R30815 DVDD.n5327 DVDD.n443 0.00476
R30816 DVDD.n5323 DVDD.n443 0.00476
R30817 DVDD.n5135 DVDD.n5107 0.00476
R30818 DVDD.n5131 DVDD.n5107 0.00476
R30819 DVDD.n5131 DVDD.n5130 0.00476
R30820 DVDD.n5130 DVDD.n5129 0.00476
R30821 DVDD.n5129 DVDD.n5114 0.00476
R30822 DVDD.n5125 DVDD.n5114 0.00476
R30823 DVDD.n5125 DVDD.n5124 0.00476
R30824 DVDD.n5124 DVDD.n5123 0.00476
R30825 DVDD.n5123 DVDD.n134 0.00476
R30826 DVDD.n5852 DVDD.n134 0.00476
R30827 DVDD.n5859 DVDD.n5858 0.00476
R30828 DVDD.n5860 DVDD.n5859 0.00476
R30829 DVDD.n5860 DVDD.n126 0.00476
R30830 DVDD.n5866 DVDD.n126 0.00476
R30831 DVDD.n5867 DVDD.n5866 0.00476
R30832 DVDD.n5868 DVDD.n5867 0.00476
R30833 DVDD.n5868 DVDD.n122 0.00476
R30834 DVDD.n5874 DVDD.n122 0.00476
R30835 DVDD.n5875 DVDD.n5874 0.00476
R30836 DVDD.n5876 DVDD.n5875 0.00476
R30837 DVDD.n5909 DVDD.n115 0.00476
R30838 DVDD.n5905 DVDD.n115 0.00476
R30839 DVDD.n5905 DVDD.n5904 0.00476
R30840 DVDD.n5904 DVDD.n5903 0.00476
R30841 DVDD.n5903 DVDD.n5891 0.00476
R30842 DVDD.n5899 DVDD.n5891 0.00476
R30843 DVDD.n4417 DVDD.n1104 0.00476
R30844 DVDD.n4423 DVDD.n1104 0.00476
R30845 DVDD.n4424 DVDD.n4423 0.00476
R30846 DVDD.n4425 DVDD.n4424 0.00476
R30847 DVDD.n4425 DVDD.n1100 0.00476
R30848 DVDD.n4431 DVDD.n1100 0.00476
R30849 DVDD.n4432 DVDD.n4431 0.00476
R30850 DVDD.n4433 DVDD.n4432 0.00476
R30851 DVDD.n4446 DVDD.n4445 0.00476
R30852 DVDD.n4446 DVDD.n1092 0.00476
R30853 DVDD.n4452 DVDD.n1092 0.00476
R30854 DVDD.n4453 DVDD.n4452 0.00476
R30855 DVDD.n4454 DVDD.n4453 0.00476
R30856 DVDD.n4454 DVDD.n1088 0.00476
R30857 DVDD.n4460 DVDD.n1088 0.00476
R30858 DVDD.n4461 DVDD.n4460 0.00476
R30859 DVDD.n4462 DVDD.n4461 0.00476
R30860 DVDD.n4462 DVDD.n1075 0.00476
R30861 DVDD.n4496 DVDD.n4495 0.00476
R30862 DVDD.n4495 DVDD.n4494 0.00476
R30863 DVDD.n4494 DVDD.n4469 0.00476
R30864 DVDD.n4490 DVDD.n4469 0.00476
R30865 DVDD.n4490 DVDD.n4489 0.00476
R30866 DVDD.n4489 DVDD.n4488 0.00476
R30867 DVDD.n4488 DVDD.n4475 0.00476
R30868 DVDD.n4484 DVDD.n4475 0.00476
R30869 DVDD.n4484 DVDD.n4483 0.00476
R30870 DVDD.n4483 DVDD.n4482 0.00476
R30871 DVDD.n4889 DVDD.n4888 0.00476
R30872 DVDD.n4890 DVDD.n4889 0.00476
R30873 DVDD.n4890 DVDD.n691 0.00476
R30874 DVDD.n4896 DVDD.n691 0.00476
R30875 DVDD.n4897 DVDD.n4896 0.00476
R30876 DVDD.n4898 DVDD.n4897 0.00476
R30877 DVDD.n4898 DVDD.n687 0.00476
R30878 DVDD.n4904 DVDD.n687 0.00476
R30879 DVDD.n4905 DVDD.n4904 0.00476
R30880 DVDD.n4906 DVDD.n4905 0.00476
R30881 DVDD.n4906 DVDD.n674 0.00476
R30882 DVDD.n4937 DVDD.n4936 0.00476
R30883 DVDD.n4936 DVDD.n4935 0.00476
R30884 DVDD.n4935 DVDD.n4913 0.00476
R30885 DVDD.n4931 DVDD.n4913 0.00476
R30886 DVDD.n4931 DVDD.n4930 0.00476
R30887 DVDD.n4930 DVDD.n4929 0.00476
R30888 DVDD.n4929 DVDD.n4919 0.00476
R30889 DVDD.n4925 DVDD.n4919 0.00476
R30890 DVDD.n4925 DVDD.n4924 0.00476
R30891 DVDD.n4924 DVDD.n451 0.00476
R30892 DVDD.n5317 DVDD.n475 0.00476
R30893 DVDD.n5313 DVDD.n475 0.00476
R30894 DVDD.n5313 DVDD.n5312 0.00476
R30895 DVDD.n5312 DVDD.n5311 0.00476
R30896 DVDD.n5311 DVDD.n5257 0.00476
R30897 DVDD.n5307 DVDD.n5257 0.00476
R30898 DVDD.n5307 DVDD.n5306 0.00476
R30899 DVDD.n5306 DVDD.n5305 0.00476
R30900 DVDD.n5305 DVDD.n5263 0.00476
R30901 DVDD.n5301 DVDD.n5263 0.00476
R30902 DVDD.n5297 DVDD.n155 0.00476
R30903 DVDD.n5297 DVDD.n5296 0.00476
R30904 DVDD.n5296 DVDD.n5295 0.00476
R30905 DVDD.n5295 DVDD.n5272 0.00476
R30906 DVDD.n5291 DVDD.n5272 0.00476
R30907 DVDD.n5291 DVDD.n5290 0.00476
R30908 DVDD.n5290 DVDD.n5289 0.00476
R30909 DVDD.n5289 DVDD.n5278 0.00476
R30910 DVDD.n5285 DVDD.n5278 0.00476
R30911 DVDD.n5285 DVDD.n42 0.00476
R30912 DVDD.n5603 DVDD.n5577 0.00476
R30913 DVDD.n5599 DVDD.n5577 0.00476
R30914 DVDD.n5599 DVDD.n5598 0.00476
R30915 DVDD.n5598 DVDD.n5597 0.00476
R30916 DVDD.n5597 DVDD.n5585 0.00476
R30917 DVDD.n5593 DVDD.n5585 0.00476
R30918 DVDD.n4370 DVDD.n1607 0.00476
R30919 DVDD.n4370 DVDD.n4369 0.00476
R30920 DVDD.n4369 DVDD.n4368 0.00476
R30921 DVDD.n4368 DVDD.n4352 0.00476
R30922 DVDD.n4364 DVDD.n4352 0.00476
R30923 DVDD.n4364 DVDD.n4363 0.00476
R30924 DVDD.n4363 DVDD.n4362 0.00476
R30925 DVDD.n4362 DVDD.n975 0.00476
R30926 DVDD.n4635 DVDD.n4634 0.00476
R30927 DVDD.n4634 DVDD.n4633 0.00476
R30928 DVDD.n4633 DVDD.n993 0.00476
R30929 DVDD.n4629 DVDD.n993 0.00476
R30930 DVDD.n4629 DVDD.n4628 0.00476
R30931 DVDD.n4628 DVDD.n4627 0.00476
R30932 DVDD.n4627 DVDD.n999 0.00476
R30933 DVDD.n4623 DVDD.n999 0.00476
R30934 DVDD.n4623 DVDD.n4622 0.00476
R30935 DVDD.n4622 DVDD.n4621 0.00476
R30936 DVDD.n1046 DVDD.n1045 0.00476
R30937 DVDD.n1045 DVDD.n1020 0.00476
R30938 DVDD.n1041 DVDD.n1020 0.00476
R30939 DVDD.n1041 DVDD.n1040 0.00476
R30940 DVDD.n1040 DVDD.n1039 0.00476
R30941 DVDD.n1039 DVDD.n1026 0.00476
R30942 DVDD.n1035 DVDD.n1026 0.00476
R30943 DVDD.n1035 DVDD.n1034 0.00476
R30944 DVDD.n1034 DVDD.n728 0.00476
R30945 DVDD.n4876 DVDD.n728 0.00476
R30946 DVDD.n4870 DVDD.n715 0.00476
R30947 DVDD.n4870 DVDD.n4869 0.00476
R30948 DVDD.n4869 DVDD.n4868 0.00476
R30949 DVDD.n4868 DVDD.n4808 0.00476
R30950 DVDD.n4864 DVDD.n4808 0.00476
R30951 DVDD.n4864 DVDD.n4863 0.00476
R30952 DVDD.n4863 DVDD.n4862 0.00476
R30953 DVDD.n4862 DVDD.n4814 0.00476
R30954 DVDD.n4858 DVDD.n4814 0.00476
R30955 DVDD.n4858 DVDD.n4857 0.00476
R30956 DVDD.n4857 DVDD.n605 0.00476
R30957 DVDD.n4852 DVDD.n4851 0.00476
R30958 DVDD.n4851 DVDD.n4850 0.00476
R30959 DVDD.n4850 DVDD.n4824 0.00476
R30960 DVDD.n4846 DVDD.n4824 0.00476
R30961 DVDD.n4846 DVDD.n4845 0.00476
R30962 DVDD.n4845 DVDD.n4844 0.00476
R30963 DVDD.n4844 DVDD.n4830 0.00476
R30964 DVDD.n4840 DVDD.n4830 0.00476
R30965 DVDD.n4840 DVDD.n4839 0.00476
R30966 DVDD.n4839 DVDD.n4838 0.00476
R30967 DVDD.n555 DVDD.n554 0.00476
R30968 DVDD.n554 DVDD.n496 0.00476
R30969 DVDD.n550 DVDD.n496 0.00476
R30970 DVDD.n550 DVDD.n549 0.00476
R30971 DVDD.n549 DVDD.n548 0.00476
R30972 DVDD.n548 DVDD.n502 0.00476
R30973 DVDD.n544 DVDD.n502 0.00476
R30974 DVDD.n544 DVDD.n543 0.00476
R30975 DVDD.n543 DVDD.n542 0.00476
R30976 DVDD.n542 DVDD.n170 0.00476
R30977 DVDD.n537 DVDD.n536 0.00476
R30978 DVDD.n536 DVDD.n535 0.00476
R30979 DVDD.n535 DVDD.n514 0.00476
R30980 DVDD.n531 DVDD.n514 0.00476
R30981 DVDD.n531 DVDD.n530 0.00476
R30982 DVDD.n530 DVDD.n529 0.00476
R30983 DVDD.n529 DVDD.n520 0.00476
R30984 DVDD.n525 DVDD.n520 0.00476
R30985 DVDD.n525 DVDD.n39 0.00476
R30986 DVDD.n5941 DVDD.n39 0.00476
R30987 DVDD.n5958 DVDD.n5957 0.00476
R30988 DVDD.n5958 DVDD.n3 0.00476
R30989 DVDD.n5965 DVDD.n3 0.00476
R30990 DVDD.n5966 DVDD.n5965 0.00476
R30991 DVDD.n5967 DVDD.n5966 0.00476
R30992 DVDD.n5967 DVDD.n0 0.00476
R30993 DVDD.n4327 DVDD.n1639 0.00476
R30994 DVDD.n4327 DVDD.n4326 0.00476
R30995 DVDD.n4326 DVDD.n4325 0.00476
R30996 DVDD.n4325 DVDD.n4307 0.00476
R30997 DVDD.n4321 DVDD.n4307 0.00476
R30998 DVDD.n4321 DVDD.n4320 0.00476
R30999 DVDD.n4320 DVDD.n4319 0.00476
R31000 DVDD.n4319 DVDD.n4313 0.00476
R31001 DVDD.n4721 DVDD.n905 0.00476
R31002 DVDD.n4727 DVDD.n905 0.00476
R31003 DVDD.n4728 DVDD.n4727 0.00476
R31004 DVDD.n4729 DVDD.n4728 0.00476
R31005 DVDD.n4729 DVDD.n901 0.00476
R31006 DVDD.n4735 DVDD.n901 0.00476
R31007 DVDD.n4736 DVDD.n4735 0.00476
R31008 DVDD.n4737 DVDD.n4736 0.00476
R31009 DVDD.n4737 DVDD.n897 0.00476
R31010 DVDD.n4743 DVDD.n897 0.00476
R31011 DVDD.n4747 DVDD.n887 0.00476
R31012 DVDD.n4753 DVDD.n887 0.00476
R31013 DVDD.n4754 DVDD.n4753 0.00476
R31014 DVDD.n4755 DVDD.n4754 0.00476
R31015 DVDD.n4755 DVDD.n883 0.00476
R31016 DVDD.n4761 DVDD.n883 0.00476
R31017 DVDD.n4762 DVDD.n4761 0.00476
R31018 DVDD.n4763 DVDD.n4762 0.00476
R31019 DVDD.n4763 DVDD.n879 0.00476
R31020 DVDD.n4771 DVDD.n879 0.00476
R31021 DVDD.n4802 DVDD.n4801 0.00476
R31022 DVDD.n4801 DVDD.n4800 0.00476
R31023 DVDD.n4800 DVDD.n4776 0.00476
R31024 DVDD.n4796 DVDD.n4776 0.00476
R31025 DVDD.n4796 DVDD.n4795 0.00476
R31026 DVDD.n4795 DVDD.n4794 0.00476
R31027 DVDD.n4794 DVDD.n4782 0.00476
R31028 DVDD.n4790 DVDD.n4782 0.00476
R31029 DVDD.n4790 DVDD.n4789 0.00476
R31030 DVDD.n4789 DVDD.n588 0.00476
R31031 DVDD.n5023 DVDD.n588 0.00476
R31032 DVDD.n5030 DVDD.n5029 0.00476
R31033 DVDD.n5031 DVDD.n5030 0.00476
R31034 DVDD.n5031 DVDD.n580 0.00476
R31035 DVDD.n5037 DVDD.n580 0.00476
R31036 DVDD.n5038 DVDD.n5037 0.00476
R31037 DVDD.n5039 DVDD.n5038 0.00476
R31038 DVDD.n5039 DVDD.n576 0.00476
R31039 DVDD.n5045 DVDD.n576 0.00476
R31040 DVDD.n5046 DVDD.n5045 0.00476
R31041 DVDD.n5047 DVDD.n5046 0.00476
R31042 DVDD.n5084 DVDD.n5083 0.00476
R31043 DVDD.n5083 DVDD.n5082 0.00476
R31044 DVDD.n5082 DVDD.n5054 0.00476
R31045 DVDD.n5078 DVDD.n5054 0.00476
R31046 DVDD.n5078 DVDD.n5077 0.00476
R31047 DVDD.n5077 DVDD.n5076 0.00476
R31048 DVDD.n5076 DVDD.n5060 0.00476
R31049 DVDD.n5072 DVDD.n5060 0.00476
R31050 DVDD.n5072 DVDD.n5071 0.00476
R31051 DVDD.n5071 DVDD.n5070 0.00476
R31052 DVDD.n5729 DVDD.n199 0.00476
R31053 DVDD.n5725 DVDD.n199 0.00476
R31054 DVDD.n5725 DVDD.n5724 0.00476
R31055 DVDD.n5724 DVDD.n5723 0.00476
R31056 DVDD.n5723 DVDD.n205 0.00476
R31057 DVDD.n5719 DVDD.n205 0.00476
R31058 DVDD.n5719 DVDD.n5718 0.00476
R31059 DVDD.n5718 DVDD.n5717 0.00476
R31060 DVDD.n5717 DVDD.n211 0.00476
R31061 DVDD.n5713 DVDD.n211 0.00476
R31062 DVDD.n5698 DVDD.n234 0.00476
R31063 DVDD.n5698 DVDD.n5697 0.00476
R31064 DVDD.n5697 DVDD.n5696 0.00476
R31065 DVDD.n5696 DVDD.n5681 0.00476
R31066 DVDD.n5692 DVDD.n5681 0.00476
R31067 DVDD.n5692 DVDD.n5691 0.00476
R31068 DVDD.n3212 DVDD.n3211 0.00473767
R31069 DVDD.n3209 DVDD.n3120 0.00473767
R31070 DVDD.n5342 DVDD.n426 0.00473
R31071 DVDD.n5340 DVDD.n5339 0.00473
R31072 DVDD.n5006 DVDD.n4940 0.00473
R31073 DVDD.n4937 DVDD.n672 0.00473
R31074 DVDD.n5014 DVDD.n616 0.00473
R31075 DVDD.n4852 DVDD.n603 0.00473
R31076 DVDD.n5022 DVDD.n591 0.00473
R31077 DVDD.n5029 DVDD.n584 0.00473
R31078 DVDD.n4081 DVDD.n4042 0.0047
R31079 DVDD.n3233 DVDD.n3105 0.00464
R31080 DVDD.n3185 DVDD.n3092 0.00464
R31081 DVDD.n3241 DVDD.n3089 0.00464
R31082 DVDD.n3244 DVDD.n3081 0.00464
R31083 DVDD.n3260 DVDD.n2962 0.00464
R31084 DVDD.n3165 DVDD.n3136 0.00464
R31085 DVDD.n3181 DVDD.n3137 0.00464
R31086 DVDD.n3141 DVDD.n3126 0.00464
R31087 DVDD.n3198 DVDD.n3127 0.00464
R31088 DVDD.n3208 DVDD.n2752 0.00464
R31089 DVDD.n4104 DVDD.n4103 0.004625
R31090 DVDD.n5420 DVDD.n260 0.0045724
R31091 DVDD.n261 DVDD.n260 0.0045724
R31092 DVDD.n5799 DVDD.n153 0.00455738
R31093 DVDD.n5155 DVDD.n452 0.00455738
R31094 DVDD.n4987 DVDD.n675 0.00455738
R31095 DVDD.n777 DVDD.n776 0.00455738
R31096 DVDD.n4543 DVDD.n1076 0.00455738
R31097 DVDD.n3955 DVDD.n3954 0.00455
R31098 DVDD.n83 DVDD.n81 0.00452754
R31099 DVDD.n5552 DVDD.n16 0.00452754
R31100 DVDD.n5658 DVDD.n8 0.00452754
R31101 DVDD.n4664 DVDD.n983 0.00452754
R31102 DVDD.n5484 DVDD.n267 0.00452754
R31103 DVDD.n5428 DVDD.n5427 0.00452754
R31104 DVDD.n4767 DVDD.n697 0.0045
R31105 DVDD.n5050 DVDD.n477 0.0045
R31106 DVDD.n4442 DVDD.n1094 0.0045
R31107 DVDD.n4885 DVDD.n697 0.0045
R31108 DVDD.n4442 DVDD.n1095 0.0045
R31109 DVDD.n4885 DVDD.n699 0.0045
R31110 DVDD.n5879 DVDD.n35 0.0045
R31111 DVDD.n5251 DVDD.n477 0.0045
R31112 DVDD.n5251 DVDD.n478 0.0045
R31113 DVDD.n5944 DVDD.n34 0.0045
R31114 DVDD.n5944 DVDD.n35 0.0045
R31115 DVDD.n1094 DVDD.n907 0.0045
R31116 DVDD.n5912 DVDD.n98 0.0044433
R31117 DVDD.n114 DVDD.n88 0.0044433
R31118 DVDD.n5415 DVDD.n337 0.0044433
R31119 DVDD.n5412 DVDD.n334 0.0044433
R31120 DVDD.n936 DVDD.n926 0.0044433
R31121 DVDD.n955 DVDD.n919 0.0044433
R31122 DVDD.n242 DVDD.n232 0.0044433
R31123 DVDD.n250 DVDD.n238 0.0044433
R31124 DVDD.n4129 DVDD.n1780 0.00443
R31125 DVDD.n2361 DVDD.n2062 0.00442143
R31126 DVDD.n2605 DVDD.n2508 0.00441304
R31127 DVDD.n1740 DVDD.n1737 0.0044
R31128 DVDD.n4016 DVDD.n4012 0.00437
R31129 DVDD.n5852 DVDD.n5851 0.00437
R31130 DVDD.n137 DVDD.n130 0.00437
R31131 DVDD.n5301 DVDD.n143 0.00437
R31132 DVDD.n5836 DVDD.n144 0.00437
R31133 DVDD.n5785 DVDD.n170 0.00437
R31134 DVDD.n180 DVDD.n169 0.00437
R31135 DVDD.n5070 DVDD.n196 0.00437
R31136 DVDD.n5735 DVDD.n197 0.00437
R31137 DVDD.n333 DVDD.n332 0.00434971
R31138 DVDD.n85 DVDD.n75 0.00434083
R31139 DVDD.n3922 DVDD.n1817 0.004325
R31140 DVDD.n3444 DVDD.n2689 0.00431
R31141 DVDD.n5383 DVDD.n379 0.00431
R31142 DVDD.n5381 DVDD.n5380 0.00431
R31143 DVDD.n4562 DVDD.n4499 0.00431
R31144 DVDD.n4496 DVDD.n1073 0.00431
R31145 DVDD.n4618 DVDD.n1005 0.00431
R31146 DVDD.n4617 DVDD.n1046 0.00431
R31147 DVDD.n4744 DVDD.n891 0.00431
R31148 DVDD.n4747 DVDD.n4746 0.00431
R31149 DVDD.n2344 DVDD.n2099 0.00429286
R31150 DVDD.n3754 DVDD.n3736 0.00425
R31151 DVDD.n3779 DVDD.n1856 0.00425
R31152 DVDD.n3997 DVDD.n1807 0.00425
R31153 DVDD.n1579 DVDD.n1181 0.00425
R31154 DVDD.n1582 DVDD.n1121 0.00425
R31155 DVDD.n4412 DVDD.n4400 0.00425
R31156 DVDD.n4416 DVDD.n1108 0.00425
R31157 DVDD.n4385 DVDD.n4375 0.00425
R31158 DVDD.n4388 DVDD.n1596 0.00425
R31159 DVDD.n4342 DVDD.n4332 0.00425
R31160 DVDD.n4345 DVDD.n1628 0.00425
R31161 DVDD.n5535 DVDD.n23 0.00421773
R31162 DVDD.n4681 DVDD.n4652 0.00421773
R31163 DVDD.n2974 DVDD.n2973 0.00419
R31164 DVDD.n2971 DVDD.n2967 0.00419
R31165 DVDD.n2981 DVDD.n2980 0.00419
R31166 DVDD.n2965 DVDD.n2732 0.00419
R31167 DVDD.n3395 DVDD.n3393 0.00419
R31168 DVDD.n3394 DVDD.n2729 0.00419
R31169 DVDD.n3399 DVDD.n3398 0.00419
R31170 DVDD.n3341 DVDD.n2862 0.00419
R31171 DVDD.n2872 DVDD.n2859 0.00419
R31172 DVDD.n2799 DVDD.n2777 0.00419
R31173 DVDD.n3348 DVDD.n2780 0.00419
R31174 DVDD.n4150 DVDD.n4148 0.00419
R31175 DVDD.n4200 DVDD.n4191 0.00419
R31176 DVDD.n5784 DVDD.n5783 0.00418852
R31177 DVDD.n5210 DVDD.n559 0.00418852
R31178 DVDD.n659 DVDD.n625 0.00418852
R31179 DVDD.n834 DVDD.n719 0.00418852
R31180 DVDD.n4583 DVDD.n1050 0.00418852
R31181 DVDD.n2831 DVDD.n2793 0.00416848
R31182 DVDD.n2906 DVDD.n2878 0.00416848
R31183 DVDD.n2717 DVDD 0.00408591
R31184 DVDD.n4241 DVDD.n1706 0.00407
R31185 DVDD.n4241 DVDD.n4240 0.00407
R31186 DVDD.n3760 DVDD.n3756 0.00404577
R31187 DVDD.n3770 DVDD.n3761 0.00404577
R31188 DVDD.n3769 DVDD.n3762 0.00404577
R31189 DVDD.n3766 DVDD.n3765 0.00404577
R31190 DVDD.n4290 DVDD.n1665 0.00404577
R31191 DVDD.n4291 DVDD.n1663 0.00404577
R31192 DVDD.n4296 DVDD.n4294 0.00404577
R31193 DVDD.n4295 DVDD.n1659 0.00404577
R31194 DVDD.n5712 DVDD.n5711 0.00404
R31195 DVDD.n38 DVDD.n33 0.00404
R31196 DVDD.n5937 DVDD.n44 0.00404
R31197 DVDD.n5881 DVDD.n119 0.00404
R31198 DVDD.n4221 DVDD.n1724 0.00404
R31199 DVDD.n80 DVDD.n41 0.00404
R31200 DVDD.n5939 DVDD.n5938 0.00404
R31201 DVDD.n5940 DVDD.n32 0.00404
R31202 DVDD.n5710 DVDD.n40 0.00404
R31203 DVDD.n4260 DVDD.n1686 0.004025
R31204 DVDD.n3271 DVDD.n3269 0.00401
R31205 DVDD.n3270 DVDD.n2931 0.00401
R31206 DVDD.n3283 DVDD.n3282 0.00401
R31207 DVDD.n3290 DVDD.n2927 0.00401
R31208 DVDD.n3293 DVDD.n2923 0.00401
R31209 DVDD.n3303 DVDD.n3302 0.00401
R31210 DVDD.n3324 DVDD.n2918 0.00401
R31211 DVDD.n3323 DVDD.n2919 0.00401
R31212 DVDD.n2938 DVDD.n2758 0.00401
R31213 DVDD.n2947 DVDD.n2759 0.00401
R31214 DVDD.n2946 DVDD.n2945 0.00401
R31215 DVDD.n3372 DVDD.n2762 0.00401
R31216 DVDD.n3365 DVDD.n2769 0.00401
R31217 DVDD.n3364 DVDD.n2770 0.00401
R31218 DVDD.n2808 DVDD.n2807 0.00401
R31219 DVDD.n2801 DVDD.n2775 0.00401
R31220 DVDD.n3406 DVDD.n3405 0.00395
R31221 DVDD.n3409 DVDD.n2724 0.00395
R31222 DVDD.n3411 DVDD.n3410 0.00395
R31223 DVDD.n3418 DVDD.n2706 0.00395
R31224 DVDD.n3424 DVDD.n3423 0.00395
R31225 DVDD.n2704 DVDD.n2698 0.00395
R31226 DVDD.n3432 DVDD.n3431 0.00395
R31227 DVDD.n3434 DVDD.n2696 0.00395
R31228 DVDD.n4148 DVDD.n1712 0.00395
R31229 DVDD DVDD.n5686 0.00392
R31230 DVDD.n5969 DVDD 0.00392
R31231 DVDD.n5594 DVDD 0.00392
R31232 DVDD.n5900 DVDD 0.00392
R31233 DVDD.n4193 DVDD 0.00392
R31234 DVDD DVDD.n4189 0.00392
R31235 DVDD.n5899 DVDD 0.00392
R31236 DVDD.n5593 DVDD 0.00392
R31237 DVDD DVDD.n0 0.00392
R31238 DVDD.n5691 DVDD 0.00392
R31239 DVDD.n5519 DVDD.n9 0.00390792
R31240 DVDD.n4698 DVDD.n976 0.00390792
R31241 DVDD.n3007 DVDD.n3001 0.00386
R31242 DVDD.n3047 DVDD.n3015 0.00386
R31243 DVDD.n5086 DVDD.n481 0.0038
R31244 DVDD.n5247 DVDD.n5246 0.0038
R31245 DVDD.n5248 DVDD.n476 0.0038
R31246 DVDD.n5108 DVDD.n448 0.0038
R31247 DVDD.n1792 DVDD.n1788 0.0038
R31248 DVDD.n4035 DVDD.n1786 0.0038
R31249 DVDD.n2141 DVDD.n2132 0.00377857
R31250 DVDD.n2286 DVDD.n2126 0.00377857
R31251 DVDD.n2159 DVDD.n2127 0.00377857
R31252 DVDD.n3255 DVDD 0.00376574
R31253 DVDD DVDD.n2750 0.00376574
R31254 DVDD DVDD.n1896 0.00376574
R31255 DVDD.n3691 DVDD 0.00376574
R31256 DVDD.n2822 DVDD.n2791 0.00367935
R31257 DVDD.n3340 DVDD.n3338 0.00367935
R31258 DVDD.n4079 DVDD.n4046 0.00365
R31259 DVDD.n4083 DVDD.n4044 0.00365
R31260 DVDD.n4161 DVDD.n1769 0.00365
R31261 DVDD.n5613 DVDD.n5576 0.00359811
R31262 DVDD.n5438 DVDD.n283 0.00359811
R31263 DVDD.n3048 DVDD.n3011 0.00359
R31264 DVDD.n4250 DVDD.n1695 0.00359
R31265 DVDD.n350 DVDD.n340 0.00357827
R31266 DVDD.n5422 DVDD.n351 0.00357827
R31267 DVDD.n106 DVDD.n105 0.00357827
R31268 DVDD.n5919 DVDD.n87 0.00357827
R31269 DVDD.n351 DVDD.n350 0.00357827
R31270 DVDD.n105 DVDD.n87 0.00357827
R31271 DVDD.n5424 DVDD.n340 0.00357827
R31272 DVDD.n5917 DVDD.n106 0.00357827
R31273 DVDD.n4804 DVDD.n4803 0.00356
R31274 DVDD.n4873 DVDD.n4872 0.00356
R31275 DVDD.n4887 DVDD.n696 0.00356
R31276 DVDD.n5359 DVDD.n407 0.00356
R31277 DVDD.n3979 DVDD.n1818 0.00356
R31278 DVDD.n3978 DVDD.n3977 0.00356
R31279 DVDD.n4252 DVDD.n1691 0.00353
R31280 DVDD.n4121 DVDD.n1786 0.00353
R31281 DVDD.n3056 DVDD.n3055 0.00347
R31282 DVDD.n4160 DVDD.n4159 0.00347
R31283 DVDD.n2204 DVDD.n2203 0.00345714
R31284 DVDD.n191 DVDD.n178 0.00345082
R31285 DVDD.n5209 DVDD.n493 0.00345082
R31286 DVDD.n660 DVDD.n614 0.00345082
R31287 DVDD.n833 DVDD.n712 0.00345082
R31288 DVDD.n4582 DVDD.n1017 0.00345082
R31289 DVDD.n3272 DVDD.n2956 0.00343478
R31290 DVDD.n2939 DVDD.n2934 0.00343478
R31291 DVDD.n3976 DVDD.n3925 0.00341
R31292 DVDD.n2974 DVDD.n2970 0.00338032
R31293 DVDD.n3060 DVDD.n3059 0.00335
R31294 DVDD.n1152 DVDD.n1151 0.00334
R31295 DVDD.n1153 DVDD.n1152 0.00334
R31296 DVDD.n1156 DVDD.n1153 0.00334
R31297 DVDD.n1157 DVDD.n1156 0.00334
R31298 DVDD.n1158 DVDD.n1157 0.00334
R31299 DVDD.n1159 DVDD.n1158 0.00334
R31300 DVDD.n1162 DVDD.n1159 0.00334
R31301 DVDD.n1163 DVDD.n1162 0.00334
R31302 DVDD.n1165 DVDD.n1163 0.00334
R31303 DVDD.n1165 DVDD.n1164 0.00334
R31304 DVDD.n1164 DVDD.n355 0.00334
R31305 DVDD.n356 DVDD.n355 0.00334
R31306 DVDD.n357 DVDD.n356 0.00334
R31307 DVDD.n362 DVDD.n361 0.00334
R31308 DVDD.n363 DVDD.n362 0.00334
R31309 DVDD.n366 DVDD.n363 0.00334
R31310 DVDD.n367 DVDD.n366 0.00334
R31311 DVDD.n368 DVDD.n367 0.00334
R31312 DVDD.n369 DVDD.n368 0.00334
R31313 DVDD.n372 DVDD.n369 0.00334
R31314 DVDD.n373 DVDD.n372 0.00334
R31315 DVDD.n374 DVDD.n373 0.00334
R31316 DVDD.n375 DVDD.n374 0.00334
R31317 DVDD.n383 DVDD.n375 0.00334
R31318 DVDD.n384 DVDD.n383 0.00334
R31319 DVDD.n385 DVDD.n384 0.00334
R31320 DVDD.n386 DVDD.n385 0.00334
R31321 DVDD.n389 DVDD.n386 0.00334
R31322 DVDD.n390 DVDD.n389 0.00334
R31323 DVDD.n391 DVDD.n390 0.00334
R31324 DVDD.n392 DVDD.n391 0.00334
R31325 DVDD.n395 DVDD.n392 0.00334
R31326 DVDD.n396 DVDD.n395 0.00334
R31327 DVDD.n397 DVDD.n396 0.00334
R31328 DVDD.n398 DVDD.n397 0.00334
R31329 DVDD.n698 DVDD.n398 0.00334
R31330 DVDD.n409 DVDD.n408 0.00334
R31331 DVDD.n410 DVDD.n409 0.00334
R31332 DVDD.n413 DVDD.n410 0.00334
R31333 DVDD.n414 DVDD.n413 0.00334
R31334 DVDD.n415 DVDD.n414 0.00334
R31335 DVDD.n416 DVDD.n415 0.00334
R31336 DVDD.n419 DVDD.n416 0.00334
R31337 DVDD.n420 DVDD.n419 0.00334
R31338 DVDD.n421 DVDD.n420 0.00334
R31339 DVDD.n422 DVDD.n421 0.00334
R31340 DVDD.n431 DVDD.n422 0.00334
R31341 DVDD.n432 DVDD.n431 0.00334
R31342 DVDD.n433 DVDD.n432 0.00334
R31343 DVDD.n434 DVDD.n433 0.00334
R31344 DVDD.n435 DVDD.n434 0.00334
R31345 DVDD.n438 DVDD.n435 0.00334
R31346 DVDD.n439 DVDD.n438 0.00334
R31347 DVDD.n440 DVDD.n439 0.00334
R31348 DVDD.n441 DVDD.n440 0.00334
R31349 DVDD.n444 DVDD.n441 0.00334
R31350 DVDD.n445 DVDD.n444 0.00334
R31351 DVDD.n446 DVDD.n445 0.00334
R31352 DVDD.n447 DVDD.n446 0.00334
R31353 DVDD.n5110 DVDD.n5109 0.00334
R31354 DVDD.n5111 DVDD.n5110 0.00334
R31355 DVDD.n5112 DVDD.n5111 0.00334
R31356 DVDD.n5115 DVDD.n5112 0.00334
R31357 DVDD.n5116 DVDD.n5115 0.00334
R31358 DVDD.n5117 DVDD.n5116 0.00334
R31359 DVDD.n5118 DVDD.n5117 0.00334
R31360 DVDD.n5120 DVDD.n5118 0.00334
R31361 DVDD.n5121 DVDD.n5120 0.00334
R31362 DVDD.n5121 DVDD.n132 0.00334
R31363 DVDD.n5854 DVDD.n132 0.00334
R31364 DVDD.n5855 DVDD.n5854 0.00334
R31365 DVDD.n5856 DVDD.n5855 0.00334
R31366 DVDD.n5856 DVDD.n128 0.00334
R31367 DVDD.n5862 DVDD.n128 0.00334
R31368 DVDD.n5863 DVDD.n5862 0.00334
R31369 DVDD.n5864 DVDD.n5863 0.00334
R31370 DVDD.n5864 DVDD.n124 0.00334
R31371 DVDD.n5870 DVDD.n124 0.00334
R31372 DVDD.n5871 DVDD.n5870 0.00334
R31373 DVDD.n5872 DVDD.n5871 0.00334
R31374 DVDD.n5872 DVDD.n120 0.00334
R31375 DVDD.n5878 DVDD.n120 0.00334
R31376 DVDD.n5880 DVDD.n118 0.00334
R31377 DVDD.n5885 DVDD.n118 0.00334
R31378 DVDD.n5886 DVDD.n5885 0.00334
R31379 DVDD.n5887 DVDD.n5886 0.00334
R31380 DVDD.n5888 DVDD.n5887 0.00334
R31381 DVDD.n5889 DVDD.n5888 0.00334
R31382 DVDD.n5892 DVDD.n5889 0.00334
R31383 DVDD.n5893 DVDD.n5892 0.00334
R31384 DVDD.n5894 DVDD.n5893 0.00334
R31385 DVDD.n5895 DVDD.n5894 0.00334
R31386 DVDD.n4419 DVDD.n1106 0.00334
R31387 DVDD.n4420 DVDD.n4419 0.00334
R31388 DVDD.n4421 DVDD.n4420 0.00334
R31389 DVDD.n4421 DVDD.n1102 0.00334
R31390 DVDD.n4427 DVDD.n1102 0.00334
R31391 DVDD.n4428 DVDD.n4427 0.00334
R31392 DVDD.n4429 DVDD.n4428 0.00334
R31393 DVDD.n4429 DVDD.n1098 0.00334
R31394 DVDD.n4435 DVDD.n1098 0.00334
R31395 DVDD.n4436 DVDD.n4435 0.00334
R31396 DVDD.n4437 DVDD.n4436 0.00334
R31397 DVDD.n4437 DVDD.n1096 0.00334
R31398 DVDD.n4441 DVDD.n1096 0.00334
R31399 DVDD.n4448 DVDD.n4443 0.00334
R31400 DVDD.n4449 DVDD.n4448 0.00334
R31401 DVDD.n4450 DVDD.n4449 0.00334
R31402 DVDD.n4450 DVDD.n1090 0.00334
R31403 DVDD.n4456 DVDD.n1090 0.00334
R31404 DVDD.n4457 DVDD.n4456 0.00334
R31405 DVDD.n4458 DVDD.n4457 0.00334
R31406 DVDD.n4458 DVDD.n1086 0.00334
R31407 DVDD.n4464 DVDD.n1086 0.00334
R31408 DVDD.n4465 DVDD.n4464 0.00334
R31409 DVDD.n4466 DVDD.n4465 0.00334
R31410 DVDD.n4467 DVDD.n4466 0.00334
R31411 DVDD.n4470 DVDD.n4467 0.00334
R31412 DVDD.n4471 DVDD.n4470 0.00334
R31413 DVDD.n4472 DVDD.n4471 0.00334
R31414 DVDD.n4473 DVDD.n4472 0.00334
R31415 DVDD.n4476 DVDD.n4473 0.00334
R31416 DVDD.n4477 DVDD.n4476 0.00334
R31417 DVDD.n4478 DVDD.n4477 0.00334
R31418 DVDD.n4479 DVDD.n4478 0.00334
R31419 DVDD.n4480 DVDD.n4479 0.00334
R31420 DVDD.n4480 DVDD.n700 0.00334
R31421 DVDD.n4884 DVDD.n700 0.00334
R31422 DVDD.n4886 DVDD.n693 0.00334
R31423 DVDD.n4892 DVDD.n693 0.00334
R31424 DVDD.n4893 DVDD.n4892 0.00334
R31425 DVDD.n4894 DVDD.n4893 0.00334
R31426 DVDD.n4894 DVDD.n689 0.00334
R31427 DVDD.n4900 DVDD.n689 0.00334
R31428 DVDD.n4901 DVDD.n4900 0.00334
R31429 DVDD.n4902 DVDD.n4901 0.00334
R31430 DVDD.n4902 DVDD.n685 0.00334
R31431 DVDD.n4908 DVDD.n685 0.00334
R31432 DVDD.n4909 DVDD.n4908 0.00334
R31433 DVDD.n4910 DVDD.n4909 0.00334
R31434 DVDD.n4911 DVDD.n4910 0.00334
R31435 DVDD.n4914 DVDD.n4911 0.00334
R31436 DVDD.n4915 DVDD.n4914 0.00334
R31437 DVDD.n4916 DVDD.n4915 0.00334
R31438 DVDD.n4917 DVDD.n4916 0.00334
R31439 DVDD.n4920 DVDD.n4917 0.00334
R31440 DVDD.n4921 DVDD.n4920 0.00334
R31441 DVDD.n4922 DVDD.n4921 0.00334
R31442 DVDD.n4923 DVDD.n4922 0.00334
R31443 DVDD.n4923 DVDD.n479 0.00334
R31444 DVDD.n5250 DVDD.n479 0.00334
R31445 DVDD.n5253 DVDD.n5252 0.00334
R31446 DVDD.n5254 DVDD.n5253 0.00334
R31447 DVDD.n5255 DVDD.n5254 0.00334
R31448 DVDD.n5258 DVDD.n5255 0.00334
R31449 DVDD.n5259 DVDD.n5258 0.00334
R31450 DVDD.n5260 DVDD.n5259 0.00334
R31451 DVDD.n5261 DVDD.n5260 0.00334
R31452 DVDD.n5264 DVDD.n5261 0.00334
R31453 DVDD.n5265 DVDD.n5264 0.00334
R31454 DVDD.n5266 DVDD.n5265 0.00334
R31455 DVDD.n5267 DVDD.n5266 0.00334
R31456 DVDD.n5268 DVDD.n5267 0.00334
R31457 DVDD.n5269 DVDD.n5268 0.00334
R31458 DVDD.n5270 DVDD.n5269 0.00334
R31459 DVDD.n5273 DVDD.n5270 0.00334
R31460 DVDD.n5274 DVDD.n5273 0.00334
R31461 DVDD.n5275 DVDD.n5274 0.00334
R31462 DVDD.n5276 DVDD.n5275 0.00334
R31463 DVDD.n5279 DVDD.n5276 0.00334
R31464 DVDD.n5280 DVDD.n5279 0.00334
R31465 DVDD.n5281 DVDD.n5280 0.00334
R31466 DVDD.n5282 DVDD.n5281 0.00334
R31467 DVDD.n5283 DVDD.n5282 0.00334
R31468 DVDD.n46 DVDD.n45 0.00334
R31469 DVDD.n5579 DVDD.n46 0.00334
R31470 DVDD.n5580 DVDD.n5579 0.00334
R31471 DVDD.n5581 DVDD.n5580 0.00334
R31472 DVDD.n5582 DVDD.n5581 0.00334
R31473 DVDD.n5583 DVDD.n5582 0.00334
R31474 DVDD.n5586 DVDD.n5583 0.00334
R31475 DVDD.n5587 DVDD.n5586 0.00334
R31476 DVDD.n5588 DVDD.n5587 0.00334
R31477 DVDD.n5589 DVDD.n5588 0.00334
R31478 DVDD.n4349 DVDD.n4348 0.00334
R31479 DVDD.n4350 DVDD.n4349 0.00334
R31480 DVDD.n4353 DVDD.n4350 0.00334
R31481 DVDD.n4354 DVDD.n4353 0.00334
R31482 DVDD.n4355 DVDD.n4354 0.00334
R31483 DVDD.n4356 DVDD.n4355 0.00334
R31484 DVDD.n4358 DVDD.n4356 0.00334
R31485 DVDD.n4360 DVDD.n4358 0.00334
R31486 DVDD.n4360 DVDD.n4359 0.00334
R31487 DVDD.n4359 DVDD.n986 0.00334
R31488 DVDD.n987 DVDD.n986 0.00334
R31489 DVDD.n988 DVDD.n987 0.00334
R31490 DVDD.n989 DVDD.n988 0.00334
R31491 DVDD.n994 DVDD.n991 0.00334
R31492 DVDD.n995 DVDD.n994 0.00334
R31493 DVDD.n996 DVDD.n995 0.00334
R31494 DVDD.n997 DVDD.n996 0.00334
R31495 DVDD.n1000 DVDD.n997 0.00334
R31496 DVDD.n1001 DVDD.n1000 0.00334
R31497 DVDD.n1002 DVDD.n1001 0.00334
R31498 DVDD.n1003 DVDD.n1002 0.00334
R31499 DVDD.n1006 DVDD.n1003 0.00334
R31500 DVDD.n1007 DVDD.n1006 0.00334
R31501 DVDD.n1008 DVDD.n1007 0.00334
R31502 DVDD.n1021 DVDD.n1008 0.00334
R31503 DVDD.n1022 DVDD.n1021 0.00334
R31504 DVDD.n1023 DVDD.n1022 0.00334
R31505 DVDD.n1024 DVDD.n1023 0.00334
R31506 DVDD.n1027 DVDD.n1024 0.00334
R31507 DVDD.n1028 DVDD.n1027 0.00334
R31508 DVDD.n1029 DVDD.n1028 0.00334
R31509 DVDD.n1030 DVDD.n1029 0.00334
R31510 DVDD.n1032 DVDD.n1030 0.00334
R31511 DVDD.n1032 DVDD.n1031 0.00334
R31512 DVDD.n1031 DVDD.n730 0.00334
R31513 DVDD.n731 DVDD.n730 0.00334
R31514 DVDD.n4806 DVDD.n4805 0.00334
R31515 DVDD.n4809 DVDD.n4806 0.00334
R31516 DVDD.n4810 DVDD.n4809 0.00334
R31517 DVDD.n4811 DVDD.n4810 0.00334
R31518 DVDD.n4812 DVDD.n4811 0.00334
R31519 DVDD.n4815 DVDD.n4812 0.00334
R31520 DVDD.n4816 DVDD.n4815 0.00334
R31521 DVDD.n4817 DVDD.n4816 0.00334
R31522 DVDD.n4818 DVDD.n4817 0.00334
R31523 DVDD.n4819 DVDD.n4818 0.00334
R31524 DVDD.n4820 DVDD.n4819 0.00334
R31525 DVDD.n4821 DVDD.n4820 0.00334
R31526 DVDD.n4822 DVDD.n4821 0.00334
R31527 DVDD.n4825 DVDD.n4822 0.00334
R31528 DVDD.n4826 DVDD.n4825 0.00334
R31529 DVDD.n4827 DVDD.n4826 0.00334
R31530 DVDD.n4828 DVDD.n4827 0.00334
R31531 DVDD.n4831 DVDD.n4828 0.00334
R31532 DVDD.n4832 DVDD.n4831 0.00334
R31533 DVDD.n4833 DVDD.n4832 0.00334
R31534 DVDD.n4834 DVDD.n4833 0.00334
R31535 DVDD.n4836 DVDD.n4834 0.00334
R31536 DVDD.n4836 DVDD.n4835 0.00334
R31537 DVDD.n497 DVDD.n483 0.00334
R31538 DVDD.n498 DVDD.n497 0.00334
R31539 DVDD.n499 DVDD.n498 0.00334
R31540 DVDD.n500 DVDD.n499 0.00334
R31541 DVDD.n503 DVDD.n500 0.00334
R31542 DVDD.n504 DVDD.n503 0.00334
R31543 DVDD.n505 DVDD.n504 0.00334
R31544 DVDD.n506 DVDD.n505 0.00334
R31545 DVDD.n508 DVDD.n506 0.00334
R31546 DVDD.n509 DVDD.n508 0.00334
R31547 DVDD.n510 DVDD.n509 0.00334
R31548 DVDD.n511 DVDD.n510 0.00334
R31549 DVDD.n512 DVDD.n511 0.00334
R31550 DVDD.n515 DVDD.n512 0.00334
R31551 DVDD.n516 DVDD.n515 0.00334
R31552 DVDD.n517 DVDD.n516 0.00334
R31553 DVDD.n518 DVDD.n517 0.00334
R31554 DVDD.n521 DVDD.n518 0.00334
R31555 DVDD.n522 DVDD.n521 0.00334
R31556 DVDD.n523 DVDD.n522 0.00334
R31557 DVDD.n524 DVDD.n523 0.00334
R31558 DVDD.n524 DVDD.n36 0.00334
R31559 DVDD.n5943 DVDD.n36 0.00334
R31560 DVDD.n5946 DVDD.n5945 0.00334
R31561 DVDD.n5947 DVDD.n5946 0.00334
R31562 DVDD.n5948 DVDD.n5947 0.00334
R31563 DVDD.n5948 DVDD.n5 0.00334
R31564 DVDD.n5960 DVDD.n5 0.00334
R31565 DVDD.n5961 DVDD.n5960 0.00334
R31566 DVDD.n5963 DVDD.n5961 0.00334
R31567 DVDD.n5963 DVDD.n5962 0.00334
R31568 DVDD.n5962 DVDD.n1 0.00334
R31569 DVDD.n5970 DVDD.n1 0.00334
R31570 DVDD.n4304 DVDD.n4303 0.00334
R31571 DVDD.n4305 DVDD.n4304 0.00334
R31572 DVDD.n4308 DVDD.n4305 0.00334
R31573 DVDD.n4309 DVDD.n4308 0.00334
R31574 DVDD.n4310 DVDD.n4309 0.00334
R31575 DVDD.n4311 DVDD.n4310 0.00334
R31576 DVDD.n4314 DVDD.n4311 0.00334
R31577 DVDD.n4315 DVDD.n4314 0.00334
R31578 DVDD.n4316 DVDD.n4315 0.00334
R31579 DVDD.n4316 DVDD.n912 0.00334
R31580 DVDD.n4715 DVDD.n912 0.00334
R31581 DVDD.n4716 DVDD.n4715 0.00334
R31582 DVDD.n4717 DVDD.n4716 0.00334
R31583 DVDD.n4724 DVDD.n4723 0.00334
R31584 DVDD.n4725 DVDD.n4724 0.00334
R31585 DVDD.n4725 DVDD.n903 0.00334
R31586 DVDD.n4731 DVDD.n903 0.00334
R31587 DVDD.n4732 DVDD.n4731 0.00334
R31588 DVDD.n4733 DVDD.n4732 0.00334
R31589 DVDD.n4733 DVDD.n899 0.00334
R31590 DVDD.n4739 DVDD.n899 0.00334
R31591 DVDD.n4740 DVDD.n4739 0.00334
R31592 DVDD.n4741 DVDD.n4740 0.00334
R31593 DVDD.n4741 DVDD.n889 0.00334
R31594 DVDD.n4749 DVDD.n889 0.00334
R31595 DVDD.n4750 DVDD.n4749 0.00334
R31596 DVDD.n4751 DVDD.n4750 0.00334
R31597 DVDD.n4751 DVDD.n885 0.00334
R31598 DVDD.n4757 DVDD.n885 0.00334
R31599 DVDD.n4758 DVDD.n4757 0.00334
R31600 DVDD.n4759 DVDD.n4758 0.00334
R31601 DVDD.n4759 DVDD.n881 0.00334
R31602 DVDD.n4765 DVDD.n881 0.00334
R31603 DVDD.n4766 DVDD.n4765 0.00334
R31604 DVDD.n4769 DVDD.n4766 0.00334
R31605 DVDD.n4769 DVDD.n4768 0.00334
R31606 DVDD.n4777 DVDD.n733 0.00334
R31607 DVDD.n4778 DVDD.n4777 0.00334
R31608 DVDD.n4779 DVDD.n4778 0.00334
R31609 DVDD.n4780 DVDD.n4779 0.00334
R31610 DVDD.n4783 DVDD.n4780 0.00334
R31611 DVDD.n4784 DVDD.n4783 0.00334
R31612 DVDD.n4785 DVDD.n4784 0.00334
R31613 DVDD.n4786 DVDD.n4785 0.00334
R31614 DVDD.n4787 DVDD.n4786 0.00334
R31615 DVDD.n4787 DVDD.n586 0.00334
R31616 DVDD.n5025 DVDD.n586 0.00334
R31617 DVDD.n5026 DVDD.n5025 0.00334
R31618 DVDD.n5027 DVDD.n5026 0.00334
R31619 DVDD.n5027 DVDD.n582 0.00334
R31620 DVDD.n5033 DVDD.n582 0.00334
R31621 DVDD.n5034 DVDD.n5033 0.00334
R31622 DVDD.n5035 DVDD.n5034 0.00334
R31623 DVDD.n5035 DVDD.n578 0.00334
R31624 DVDD.n5041 DVDD.n578 0.00334
R31625 DVDD.n5042 DVDD.n5041 0.00334
R31626 DVDD.n5043 DVDD.n5042 0.00334
R31627 DVDD.n5043 DVDD.n574 0.00334
R31628 DVDD.n5049 DVDD.n574 0.00334
R31629 DVDD.n5052 DVDD.n5051 0.00334
R31630 DVDD.n5055 DVDD.n5052 0.00334
R31631 DVDD.n5056 DVDD.n5055 0.00334
R31632 DVDD.n5057 DVDD.n5056 0.00334
R31633 DVDD.n5058 DVDD.n5057 0.00334
R31634 DVDD.n5061 DVDD.n5058 0.00334
R31635 DVDD.n5062 DVDD.n5061 0.00334
R31636 DVDD.n5063 DVDD.n5062 0.00334
R31637 DVDD.n5064 DVDD.n5063 0.00334
R31638 DVDD.n5066 DVDD.n5064 0.00334
R31639 DVDD.n5068 DVDD.n5066 0.00334
R31640 DVDD.n5068 DVDD.n5067 0.00334
R31641 DVDD.n5067 DVDD.n201 0.00334
R31642 DVDD.n202 DVDD.n201 0.00334
R31643 DVDD.n203 DVDD.n202 0.00334
R31644 DVDD.n206 DVDD.n203 0.00334
R31645 DVDD.n207 DVDD.n206 0.00334
R31646 DVDD.n208 DVDD.n207 0.00334
R31647 DVDD.n209 DVDD.n208 0.00334
R31648 DVDD.n212 DVDD.n209 0.00334
R31649 DVDD.n213 DVDD.n212 0.00334
R31650 DVDD.n214 DVDD.n213 0.00334
R31651 DVDD.n215 DVDD.n214 0.00334
R31652 DVDD.n5675 DVDD.n216 0.00334
R31653 DVDD.n5676 DVDD.n5675 0.00334
R31654 DVDD.n5677 DVDD.n5676 0.00334
R31655 DVDD.n5678 DVDD.n5677 0.00334
R31656 DVDD.n5679 DVDD.n5678 0.00334
R31657 DVDD.n5682 DVDD.n5679 0.00334
R31658 DVDD.n5683 DVDD.n5682 0.00334
R31659 DVDD.n5684 DVDD.n5683 0.00334
R31660 DVDD.n5685 DVDD.n5684 0.00334
R31661 DVDD.n5687 DVDD.n5685 0.00334
R31662 DVDD.n5688 DVDD.n5687 0.00334
R31663 DVDD.n2988 DVDD.n2737 0.00334
R31664 DVDD.n2989 DVDD.n2988 0.00334
R31665 DVDD.n2992 DVDD.n2989 0.00334
R31666 DVDD.n2993 DVDD.n2992 0.00334
R31667 DVDD.n3002 DVDD.n2994 0.00334
R31668 DVDD.n3003 DVDD.n3002 0.00334
R31669 DVDD.n3004 DVDD.n3003 0.00334
R31670 DVDD.n3005 DVDD.n3004 0.00334
R31671 DVDD.n3013 DVDD.n3012 0.00334
R31672 DVDD.n3021 DVDD.n3013 0.00334
R31673 DVDD.n3022 DVDD.n3021 0.00334
R31674 DVDD.n3023 DVDD.n3022 0.00334
R31675 DVDD.n3027 DVDD.n3024 0.00334
R31676 DVDD.n3028 DVDD.n3027 0.00334
R31677 DVDD.n3029 DVDD.n3028 0.00334
R31678 DVDD.n3029 DVDD.n1911 0.00334
R31679 DVDD.n3706 DVDD.n1912 0.00334
R31680 DVDD.n3161 DVDD.n3157 0.00334
R31681 DVDD.n3157 DVDD.n2748 0.00334
R31682 DVDD.n3388 DVDD.n2749 0.00334
R31683 DVDD.n3384 DVDD.n2749 0.00334
R31684 DVDD.n3384 DVDD.n3383 0.00334
R31685 DVDD.n3383 DVDD.n3382 0.00334
R31686 DVDD.n3378 DVDD.n2755 0.00334
R31687 DVDD.n3378 DVDD.n3377 0.00334
R31688 DVDD.n3377 DVDD.n3376 0.00334
R31689 DVDD.n3376 DVDD.n2761 0.00334
R31690 DVDD.n3362 DVDD.n2773 0.00334
R31691 DVDD.n3362 DVDD.n3361 0.00334
R31692 DVDD.n3361 DVDD.n3360 0.00334
R31693 DVDD.n3360 DVDD.n2774 0.00334
R31694 DVDD.n3356 DVDD.n3355 0.00334
R31695 DVDD.n3355 DVDD.n3354 0.00334
R31696 DVDD.n3354 DVDD.n2779 0.00334
R31697 DVDD.n2779 DVDD.n1908 0.00334
R31698 DVDD.n1969 DVDD.n1907 0.00334
R31699 DVDD.n3100 DVDD.n3099 0.00334
R31700 DVDD.n3100 DVDD.n2744 0.00334
R31701 DVDD.n3258 DVDD.n2743 0.00334
R31702 DVDD.n3258 DVDD.n2960 0.00334
R31703 DVDD.n3265 DVDD.n2960 0.00334
R31704 DVDD.n3266 DVDD.n3265 0.00334
R31705 DVDD.n3267 DVDD.n2929 0.00334
R31706 DVDD.n3285 DVDD.n2929 0.00334
R31707 DVDD.n3286 DVDD.n3285 0.00334
R31708 DVDD.n3287 DVDD.n3286 0.00334
R31709 DVDD.n3305 DVDD.n2921 0.00334
R31710 DVDD.n3306 DVDD.n3305 0.00334
R31711 DVDD.n3307 DVDD.n3306 0.00334
R31712 DVDD.n3308 DVDD.n3307 0.00334
R31713 DVDD.n3310 DVDD.n3309 0.00334
R31714 DVDD.n3311 DVDD.n3310 0.00334
R31715 DVDD.n3312 DVDD.n3311 0.00334
R31716 DVDD.n3312 DVDD.n1904 0.00334
R31717 DVDD.n1919 DVDD.n1903 0.00334
R31718 DVDD.n2978 DVDD.n2977 0.00334
R31719 DVDD.n2978 DVDD.n2739 0.00334
R31720 DVDD.n3391 DVDD.n3390 0.00334
R31721 DVDD.n3391 DVDD.n2727 0.00334
R31722 DVDD.n3401 DVDD.n2727 0.00334
R31723 DVDD.n3402 DVDD.n3401 0.00334
R31724 DVDD.n3403 DVDD.n2722 0.00334
R31725 DVDD.n3413 DVDD.n2722 0.00334
R31726 DVDD.n3414 DVDD.n3413 0.00334
R31727 DVDD.n3415 DVDD.n3414 0.00334
R31728 DVDD.n3427 DVDD.n3426 0.00334
R31729 DVDD.n3429 DVDD.n3427 0.00334
R31730 DVDD.n3429 DVDD.n3428 0.00334
R31731 DVDD.n3428 DVDD.n2694 0.00334
R31732 DVDD.n3439 DVDD.n3438 0.00334
R31733 DVDD.n3441 DVDD.n3439 0.00334
R31734 DVDD.n3441 DVDD.n3440 0.00334
R31735 DVDD.n3440 DVDD.n1900 0.00334
R31736 DVDD.n1939 DVDD.n1899 0.00334
R31737 DVDD.n3733 DVDD.n1854 0.00334
R31738 DVDD.n3784 DVDD.n1854 0.00334
R31739 DVDD.n3785 DVDD.n3784 0.00334
R31740 DVDD.n3786 DVDD.n3785 0.00334
R31741 DVDD.n3786 DVDD.n1850 0.00334
R31742 DVDD.n3792 DVDD.n1850 0.00334
R31743 DVDD.n3793 DVDD.n3792 0.00334
R31744 DVDD.n3794 DVDD.n3793 0.00334
R31745 DVDD.n3794 DVDD.n1846 0.00334
R31746 DVDD.n3801 DVDD.n1846 0.00334
R31747 DVDD.n3802 DVDD.n3801 0.00334
R31748 DVDD.n3803 DVDD.n3802 0.00334
R31749 DVDD.n3803 DVDD.n1687 0.00334
R31750 DVDD.n4259 DVDD.n1688 0.00334
R31751 DVDD.n1692 DVDD.n1688 0.00334
R31752 DVDD.n1693 DVDD.n1692 0.00334
R31753 DVDD.n1696 DVDD.n1693 0.00334
R31754 DVDD.n1697 DVDD.n1696 0.00334
R31755 DVDD.n1698 DVDD.n1697 0.00334
R31756 DVDD.n1701 DVDD.n1698 0.00334
R31757 DVDD.n1702 DVDD.n1701 0.00334
R31758 DVDD.n1703 DVDD.n1702 0.00334
R31759 DVDD.n1704 DVDD.n1703 0.00334
R31760 DVDD.n3938 DVDD.n1704 0.00334
R31761 DVDD.n3939 DVDD.n3938 0.00334
R31762 DVDD.n3940 DVDD.n3939 0.00334
R31763 DVDD.n3941 DVDD.n3940 0.00334
R31764 DVDD.n3942 DVDD.n3941 0.00334
R31765 DVDD.n3945 DVDD.n3942 0.00334
R31766 DVDD.n3946 DVDD.n3945 0.00334
R31767 DVDD.n3947 DVDD.n3946 0.00334
R31768 DVDD.n3948 DVDD.n3947 0.00334
R31769 DVDD.n3948 DVDD.n3927 0.00334
R31770 DVDD.n3972 DVDD.n3927 0.00334
R31771 DVDD.n3973 DVDD.n3972 0.00334
R31772 DVDD.n3974 DVDD.n3973 0.00334
R31773 DVDD.n3981 DVDD.n3980 0.00334
R31774 DVDD.n3982 DVDD.n3981 0.00334
R31775 DVDD.n3982 DVDD.n1813 0.00334
R31776 DVDD.n3988 DVDD.n1813 0.00334
R31777 DVDD.n3989 DVDD.n3988 0.00334
R31778 DVDD.n3990 DVDD.n3989 0.00334
R31779 DVDD.n3990 DVDD.n1809 0.00334
R31780 DVDD.n4000 DVDD.n1809 0.00334
R31781 DVDD.n4001 DVDD.n4000 0.00334
R31782 DVDD.n4002 DVDD.n4001 0.00334
R31783 DVDD.n4002 DVDD.n1805 0.00334
R31784 DVDD.n4008 DVDD.n1805 0.00334
R31785 DVDD.n4009 DVDD.n4008 0.00334
R31786 DVDD.n4010 DVDD.n4009 0.00334
R31787 DVDD.n4010 DVDD.n1801 0.00334
R31788 DVDD.n4020 DVDD.n1801 0.00334
R31789 DVDD.n4021 DVDD.n4020 0.00334
R31790 DVDD.n4022 DVDD.n4021 0.00334
R31791 DVDD.n4022 DVDD.n1797 0.00334
R31792 DVDD.n4029 DVDD.n1797 0.00334
R31793 DVDD.n4030 DVDD.n4029 0.00334
R31794 DVDD.n4031 DVDD.n4030 0.00334
R31795 DVDD.n4031 DVDD.n1789 0.00334
R31796 DVDD.n4106 DVDD.n4105 0.00334
R31797 DVDD.n4107 DVDD.n4106 0.00334
R31798 DVDD.n4108 DVDD.n4107 0.00334
R31799 DVDD.n4110 DVDD.n4108 0.00334
R31800 DVDD.n4111 DVDD.n4110 0.00334
R31801 DVDD.n4111 DVDD.n1782 0.00334
R31802 DVDD.n4132 DVDD.n1782 0.00334
R31803 DVDD.n4133 DVDD.n4132 0.00334
R31804 DVDD.n4134 DVDD.n4133 0.00334
R31805 DVDD.n4134 DVDD.n1778 0.00334
R31806 DVDD.n4144 DVDD.n1778 0.00334
R31807 DVDD.n4145 DVDD.n4144 0.00334
R31808 DVDD.n4146 DVDD.n4145 0.00334
R31809 DVDD.n4146 DVDD.n1775 0.00334
R31810 DVDD.n4154 DVDD.n1775 0.00334
R31811 DVDD.n4155 DVDD.n4154 0.00334
R31812 DVDD.n4156 DVDD.n4155 0.00334
R31813 DVDD.n4156 DVDD.n1771 0.00334
R31814 DVDD.n4164 DVDD.n1771 0.00334
R31815 DVDD.n4165 DVDD.n4164 0.00334
R31816 DVDD.n4166 DVDD.n4165 0.00334
R31817 DVDD.n4166 DVDD.n1767 0.00334
R31818 DVDD.n4172 DVDD.n1767 0.00334
R31819 DVDD.n4222 DVDD.n4173 0.00334
R31820 DVDD.n4179 DVDD.n4173 0.00334
R31821 DVDD.n4180 DVDD.n4179 0.00334
R31822 DVDD.n4181 DVDD.n4180 0.00334
R31823 DVDD.n4184 DVDD.n4181 0.00334
R31824 DVDD.n4185 DVDD.n4184 0.00334
R31825 DVDD.n4186 DVDD.n4185 0.00334
R31826 DVDD.n4187 DVDD.n4186 0.00334
R31827 DVDD.n4192 DVDD.n4187 0.00334
R31828 DVDD.n4194 DVDD.n4192 0.00334
R31829 DVDD.n4195 DVDD.n4194 0.00334
R31830 DVDD.n4722 DVDD.n908 0.00332
R31831 DVDD.n4637 DVDD.n4636 0.00332
R31832 DVDD.n4444 DVDD.n990 0.00332
R31833 DVDD.n5399 DVDD.n358 0.00332
R31834 DVDD.n4258 DVDD.n1685 0.00332
R31835 DVDD.n5401 DVDD.n5400 0.00332
R31836 DVDD.n4445 DVDD.n359 0.00332
R31837 DVDD.n4635 DVDD.n909 0.00332
R31838 DVDD.n4721 DVDD.n4720 0.00332
R31839 DVDD.n5404 DVDD.n322 0.00329
R31840 DVDD.n295 DVDD.n284 0.00329
R31841 DVDD.n5474 DVDD.n297 0.00329
R31842 DVDD.n4642 DVDD.n974 0.00329
R31843 DVDD.n4640 DVDD.n972 0.00329
R31844 DVDD.n921 DVDD.n910 0.00329
R31845 DVDD.n5629 DVDD.n5607 0.0032883
R31846 DVDD.n5454 DVDD.n289 0.0032883
R31847 DVDD.n3040 DVDD.n3019 0.00323
R31848 DVDD.n4257 DVDD.n1690 0.00323
R31849 DVDD.n4116 DVDD.n4115 0.00323
R31850 DVDD.n5922 DVDD.n82 0.00323
R31851 DVDD.n5935 DVDD.n43 0.00323
R31852 DVDD.n5934 DVDD.n58 0.00323
R31853 DVDD.n5954 DVDD.n5953 0.00323
R31854 DVDD.n5950 DVDD.n29 0.00323
R31855 DVDD.n5709 DVDD.n220 0.00323
R31856 DVDD.n3900 DVDD.n3871 0.0032
R31857 DVDD.n3902 DVDD.n3901 0.0032
R31858 DVDD.n4262 DVDD.n1685 0.0032
R31859 DVDD.n3697 DVDD.n3693 0.00314706
R31860 DVDD.n4274 DVDD.n1675 0.00314375
R31861 DVDD.n1680 DVDD.n1679 0.00314375
R31862 DVDD.n4268 DVDD.n4267 0.00314375
R31863 DVDD.n4264 DVDD.n1681 0.00314375
R31864 DVDD.n4263 DVDD.n1684 0.00314375
R31865 DVDD.n3808 DVDD.n1843 0.00314375
R31866 DVDD.n3814 DVDD.n3812 0.00314375
R31867 DVDD.n3813 DVDD.n1840 0.00314375
R31868 DVDD.n3819 DVDD.n3818 0.00314375
R31869 DVDD.n1841 DVDD.n1836 0.00314375
R31870 DVDD.n2075 DVDD.n2068 0.00313571
R31871 DVDD.n2093 DVDD.n2063 0.00313571
R31872 DVDD.n3968 DVDD.n3967 0.00311
R31873 DVDD.n4331 DVDD.n4302 0.00309529
R31874 DVDD.n4374 DVDD.n4347 0.00309529
R31875 DVDD.n4411 DVDD.n4401 0.00309529
R31876 DVDD.n1180 DVDD.n1150 0.00309529
R31877 DVDD.n2976 DVDD.n2975 0.00309529
R31878 DVDD.n3104 DVDD.n3097 0.00309529
R31879 DVDD.n3162 DVDD.n3156 0.00309529
R31880 DVDD.n3735 DVDD.n3723 0.00309529
R31881 DVDD.n5798 DVDD.n156 0.00308197
R31882 DVDD.n5154 DVDD.n464 0.00308197
R31883 DVDD.n4988 DVDD.n4942 0.00308197
R31884 DVDD.n755 DVDD.n753 0.00308197
R31885 DVDD.n4544 DVDD.n4501 0.00308197
R31886 DVDD.n5883 DVDD.n77 0.00302
R31887 DVDD.n116 DVDD.n79 0.00302
R31888 DVDD.n5565 DVDD.n58 0.00302
R31889 DVDD.n5651 DVDD.n5566 0.00302
R31890 DVDD.n5950 DVDD.n31 0.00302
R31891 DVDD.n5956 DVDD.n7 0.00302
R31892 DVDD.n5703 DVDD.n224 0.00302
R31893 DVDD.n5707 DVDD.n227 0.00302
R31894 DVDD.n2369 DVDD.n2368 0.00300714
R31895 DVDD.n1573 DVDD.n1197 0.00300714
R31896 DVDD.n1572 DVDD.n1192 0.00300714
R31897 DVDD.n5646 DVDD.n5569 0.00297849
R31898 DVDD.n5472 DVDD.n276 0.00297849
R31899 DVDD.n4054 DVDD.n4049 0.002975
R31900 DVDD.n4069 DVDD.n4068 0.002975
R31901 DVDD.n4065 DVDD.n4055 0.002975
R31902 DVDD.n4064 DVDD.n4057 0.002975
R31903 DVDD.n4059 DVDD.n4058 0.002975
R31904 DVDD.n4227 DVDD.n1721 0.002975
R31905 DVDD.n1764 DVDD.n1763 0.002975
R31906 DVDD.n1760 DVDD.n1729 0.002975
R31907 DVDD.n1759 DVDD.n1730 0.002975
R31908 DVDD.n5429 DVDD.n328 0.00296
R31909 DVDD.n5407 DVDD.n321 0.00296
R31910 DVDD.n273 DVDD.n271 0.00296
R31911 DVDD.n5477 DVDD.n284 0.00296
R31912 DVDD.n4700 DVDD.n4645 0.00296
R31913 DVDD.n4642 DVDD.n971 0.00296
R31914 DVDD.n4709 DVDD.n4708 0.00296
R31915 DVDD.n4713 DVDD.n914 0.00296
R31916 DVDD.n2633 DVDD.n2446 0.00294565
R31917 DVDD.n3781 DVDD.n1852 0.00287
R31918 DVDD.n5364 DVDD.n5363 0.00287
R31919 DVDD.n4482 DVDD.n702 0.00287
R31920 DVDD.n4877 DVDD.n4876 0.00287
R31921 DVDD.n4773 DVDD.n4771 0.00287
R31922 DVDD.n5880 DVDD.n5879 0.00286
R31923 DVDD.n45 DVDD.n35 0.00286
R31924 DVDD.n5945 DVDD.n5944 0.00286
R31925 DVDD.n216 DVDD.n34 0.00286
R31926 DVDD.n4223 DVDD.n4222 0.00286
R31927 DVDD.n5611 DVDD.n67 0.00282358
R31928 DVDD.n317 DVDD.n298 0.00282358
R31929 DVDD.n3068 DVDD.n3067 0.00281
R31930 DVDD.n5106 DVDD.n449 0.00281
R31931 DVDD.n5136 DVDD.n5135 0.00281
R31932 DVDD.n5320 DVDD.n462 0.00281
R31933 DVDD.n5318 DVDD.n5317 0.00281
R31934 DVDD.n5245 DVDD.n485 0.00281
R31935 DVDD.n5244 DVDD.n555 0.00281
R31936 DVDD.n5096 DVDD.n5087 0.00281
R31937 DVDD.n5084 DVDD.n570 0.00281
R31938 DVDD DVDD.n5895 0.00278
R31939 DVDD DVDD.n5589 0.00278
R31940 DVDD DVDD.n5970 0.00278
R31941 DVDD.n3255 DVDD.n2964 0.00275
R31942 DVDD.n3691 DVDD.n1915 0.00275
R31943 DVDD.n2969 DVDD.n2750 0.00275
R31944 DVDD.n3425 DVDD.n2702 0.00275
R31945 DVDD.n2692 DVDD.n1896 0.00275
R31946 DVDD.n3101 DVDD.n2750 0.00275
R31947 DVDD.n2922 DVDD.n2702 0.00275
R31948 DVDD.n3313 DVDD.n1896 0.00275
R31949 DVDD.n3691 DVDD.n1917 0.00275
R31950 DVDD.n3691 DVDD.n1973 0.00275
R31951 DVDD.n3158 DVDD.n2750 0.00275
R31952 DVDD.n2771 DVDD.n2702 0.00275
R31953 DVDD.n3351 DVDD.n1896 0.00275
R31954 DVDD.n3050 DVDD.n2702 0.00275
R31955 DVDD.n3030 DVDD.n1896 0.00275
R31956 DVDD.n3691 DVDD.n1974 0.00275
R31957 DVDD.n3837 DVDD.n1830 0.00275
R31958 DVDD.n3857 DVDD.n1818 0.00275
R31959 DVDD.n3836 DVDD.n3835 0.00275
R31960 DVDD.n3977 DVDD.n3858 0.00275
R31961 DVDD.n4206 DVDD.n4189 0.00275
R31962 DVDD.n5762 DVDD.n176 0.00271311
R31963 DVDD.n5225 DVDD.n562 0.00271311
R31964 DVDD.n644 DVDD.n612 0.00271311
R31965 DVDD.n849 DVDD.n722 0.00271311
R31966 DVDD.n4598 DVDD.n1053 0.00271311
R31967 DVDD.n2839 DVDD.n2784 0.00270109
R31968 DVDD.n2898 DVDD.n2866 0.00270109
R31969 DVDD.n5109 DVDD.n478 0.0027
R31970 DVDD.n5252 DVDD.n5251 0.0027
R31971 DVDD.n483 DVDD.n477 0.0027
R31972 DVDD.n5051 DVDD.n5050 0.0027
R31973 DVDD.n4105 DVDD.n4104 0.0027
R31974 DVDD.n3052 DVDD.n3051 0.00269
R31975 DVDD.n3960 DVDD.n3935 0.00269
R31976 DVDD.n4140 DVDD.n4137 0.00269
R31977 DVDD.n3389 DVDD 0.00267716
R31978 DVDD.n3707 DVDD 0.00267716
R31979 DVDD.n5955 DVDD.n30 0.00266867
R31980 DVDD.n4701 DVDD.n973 0.00266867
R31981 DVDD.n3255 DVDD.n3254 0.00263
R31982 DVDD.n3255 DVDD.n3078 0.00263
R31983 DVDD.n4177 DVDD.n1722 0.00263
R31984 DVDD.n4081 DVDD.n4080 0.0026
R31985 DVDD.n3960 DVDD.n3959 0.00257
R31986 DVDD.n4142 DVDD.n4140 0.00257
R31987 DVDD.n699 DVDD.n408 0.00254
R31988 DVDD.n4886 DVDD.n4885 0.00254
R31989 DVDD.n4805 DVDD.n697 0.00254
R31990 DVDD.n4767 DVDD.n733 0.00254
R31991 DVDD.n3980 DVDD.n1817 0.00254
R31992 DVDD.n5634 DVDD.n53 0.00251377
R31993 DVDD.n5459 DVDD.n313 0.00251377
R31994 DVDD.n3417 DVDD.n2720 0.00251
R31995 DVDD.n3691 DVDD.n1914 0.00251
R31996 DVDD.n2750 DVDD.n2733 0.00251
R31997 DVDD.n3416 DVDD.n2702 0.00251
R31998 DVDD.n1940 DVDD.n1896 0.00251
R31999 DVDD.n3257 DVDD.n2750 0.00251
R32000 DVDD.n3288 DVDD.n2702 0.00251
R32001 DVDD.n1952 DVDD.n1896 0.00251
R32002 DVDD.n3256 DVDD.n3255 0.00251
R32003 DVDD.n3289 DVDD.n2720 0.00251
R32004 DVDD.n3691 DVDD.n1953 0.00251
R32005 DVDD.n3255 DVDD.n2751 0.00251
R32006 DVDD.n3373 DVDD.n2720 0.00251
R32007 DVDD.n3691 DVDD.n1972 0.00251
R32008 DVDD.n3387 DVDD.n2750 0.00251
R32009 DVDD.n3374 DVDD.n2702 0.00251
R32010 DVDD.n1971 DVDD.n1896 0.00251
R32011 DVDD.n3076 DVDD.n2750 0.00251
R32012 DVDD.n3006 DVDD.n2702 0.00251
R32013 DVDD.n3705 DVDD.n1896 0.00251
R32014 DVDD.n3255 DVDD.n3077 0.00251
R32015 DVDD.n3008 DVDD.n2720 0.00251
R32016 DVDD.n3704 DVDD.n3691 0.00251
R32017 DVDD.n4207 DVDD.n4206 0.00251
R32018 DVDD.n3681 DVDD.n1980 0.00248146
R32019 DVDD.n3682 DVDD.n1978 0.00248146
R32020 DVDD.n3687 DVDD.n3686 0.00248146
R32021 DVDD.n3690 DVDD.n1975 0.00248146
R32022 DVDD.n3710 DVDD.n1895 0.00248146
R32023 DVDD.n3711 DVDD.n1893 0.00248146
R32024 DVDD.n3716 DVDD.n3714 0.00248146
R32025 DVDD.n3715 DVDD.n1889 0.00248146
R32026 DVDD.n3067 DVDD.n2996 0.00245
R32027 DVDD.n5136 DVDD.n5106 0.00245
R32028 DVDD.n5318 DVDD.n462 0.00245
R32029 DVDD.n5245 DVDD.n5244 0.00245
R32030 DVDD.n5087 DVDD.n570 0.00245
R32031 DVDD.n3788 DVDD.n1852 0.00239
R32032 DVDD.n5363 DVDD.n402 0.00239
R32033 DVDD.n5361 DVDD.n5360 0.00239
R32034 DVDD.n4882 DVDD.n702 0.00239
R32035 DVDD.n4888 DVDD.n695 0.00239
R32036 DVDD.n4877 DVDD.n704 0.00239
R32037 DVDD.n4879 DVDD.n715 0.00239
R32038 DVDD.n4773 DVDD.n4772 0.00239
R32039 DVDD.n4802 DVDD.n4775 0.00239
R32040 DVDD.n1095 DVDD.n361 0.00238
R32041 DVDD.n4443 DVDD.n4442 0.00238
R32042 DVDD.n1094 DVDD.n991 0.00238
R32043 DVDD.n4723 DVDD.n907 0.00238
R32044 DVDD.n4260 DVDD.n4259 0.00238
R32045 DVDD.n2294 DVDD.n2293 0.00236429
R32046 DVDD.n1395 DVDD.n1305 0.00236429
R32047 DVDD.n1394 DVDD.n1310 0.00236429
R32048 DVDD.n5633 DVDD.n5572 0.00235886
R32049 DVDD.n5532 DVDD.n24 0.00235886
R32050 DVDD.n4685 DVDD.n4653 0.00235886
R32051 DVDD.n5458 DVDD.n279 0.00235886
R32052 DVDD.n5814 DVDD.n150 0.00234426
R32053 DVDD.n5170 DVDD.n466 0.00234426
R32054 DVDD.n4972 DVDD.n4944 0.00234426
R32055 DVDD.n792 DVDD.n791 0.00234426
R32056 DVDD.n4528 DVDD.n4503 0.00234426
R32057 DVDD.n2197 DVDD 0.0023
R32058 DVDD.n3471 DVDD 0.0023
R32059 DVDD.n4035 DVDD.n1794 0.0023
R32060 DVDD.n4261 DVDD.n4260 0.0023
R32061 DVDD.n3904 DVDD.n3869 0.0023
R32062 DVDD.n3881 DVDD.n1792 0.0023
R32063 DVDD.n4285 DVDD.n1666 0.0023
R32064 DVDD.n4284 DVDD.n1670 0.0023
R32065 DVDD.n1361 DVDD 0.0023
R32066 DVDD.n4433 DVDD.n271 0.0023
R32067 DVDD.n5477 DVDD.n273 0.0023
R32068 DVDD.n4700 DVDD.n975 0.0023
R32069 DVDD.n4645 DVDD.n971 0.0023
R32070 DVDD.n5486 DVDD.n5485 0.00226879
R32071 DVDD.n5660 DVDD.n5659 0.00226471
R32072 DVDD.n5566 DVDD.n5565 0.00224
R32073 DVDD.n5651 DVDD.n5603 0.00224
R32074 DVDD.n31 DVDD.n7 0.00224
R32075 DVDD.n5957 DVDD.n5956 0.00224
R32076 DVDD.n1368 DVDD 0.00223571
R32077 DVDD.n5617 DVDD.n60 0.00220396
R32078 DVDD.n5442 DVDD.n305 0.00220396
R32079 DVDD.n2437 DVDD.n2433 0.00217143
R32080 DVDD.n3967 DVDD.n3929 0.00215
R32081 DVDD.n108 DVDD.n76 0.00206
R32082 DVDD.n5704 DVDD.n226 0.00206
R32083 DVDD.n5549 DVDD.n15 0.00204905
R32084 DVDD.n4668 DVDD.n982 0.00204905
R32085 DVDD.n3040 DVDD.n3039 0.00203
R32086 DVDD.n4115 DVDD.n4114 0.00203
R32087 DVDD.n5922 DVDD.n80 0.00203
R32088 DVDD.n82 DVDD.n76 0.00203
R32089 DVDD.n5938 DVDD.n43 0.00203
R32090 DVDD.n5935 DVDD.n5934 0.00203
R32091 DVDD.n5954 DVDD.n32 0.00203
R32092 DVDD.n5953 DVDD.n29 0.00203
R32093 DVDD.n5710 DVDD.n5709 0.00203
R32094 DVDD.n226 DVDD.n220 0.00203
R32095 DVDD.n3012 DVDD.n2701 0.002
R32096 DVDD.n3707 DVDD.n1911 0.002
R32097 DVDD.n3389 DVDD.n2748 0.002
R32098 DVDD.n2773 DVDD.n2701 0.002
R32099 DVDD.n3707 DVDD.n1908 0.002
R32100 DVDD.n3389 DVDD.n2744 0.002
R32101 DVDD.n2921 DVDD.n2701 0.002
R32102 DVDD.n3707 DVDD.n1904 0.002
R32103 DVDD.n3389 DVDD.n2739 0.002
R32104 DVDD.n3426 DVDD.n2701 0.002
R32105 DVDD.n3707 DVDD.n1900 0.002
R32106 DVDD.n3294 DVDD.n2720 0.002
R32107 DVDD.n2768 DVDD.n2720 0.002
R32108 DVDD.n3838 DVDD.n1829 0.002
R32109 DVDD.n3856 DVDD.n1817 0.002
R32110 DVDD.n1161 DVDD.n325 0.002
R32111 DVDD.n353 DVDD.n328 0.002
R32112 DVDD.n5417 DVDD.n5407 0.002
R32113 DVDD.n4313 DVDD.n943 0.002
R32114 DVDD.n4710 DVDD.n4709 0.002
R32115 DVDD.n4713 DVDD.n4712 0.002
R32116 DVDD.n2259 DVDD.n2258 0.00197857
R32117 DVDD.n5746 DVDD.n174 0.00197541
R32118 DVDD.n567 DVDD.n486 0.00197541
R32119 DVDD.n628 DVDD.n610 0.00197541
R32120 DVDD.n864 DVDD.n705 0.00197541
R32121 DVDD.n1058 DVDD.n1010 0.00197541
R32122 DVDD.n5404 DVDD.n324 0.00197
R32123 DVDD.n5402 DVDD.n322 0.00197
R32124 DVDD.n297 DVDD.n295 0.00197
R32125 DVDD.n5474 DVDD.n307 0.00197
R32126 DVDD.n4640 DVDD.n974 0.00197
R32127 DVDD.n4638 DVDD.n972 0.00197
R32128 DVDD.n922 DVDD.n921 0.00197
R32129 DVDD.n4719 DVDD.n910 0.00197
R32130 DVDD.n3291 DVDD.n2926 0.00196739
R32131 DVDD.n3371 DVDD.n2763 0.00196739
R32132 DVDD.n4718 DVDD.n908 0.00194
R32133 DVDD.n4639 DVDD.n4637 0.00194
R32134 DVDD.n4440 DVDD.n990 0.00194
R32135 DVDD.n5403 DVDD.n358 0.00194
R32136 DVDD.n3255 DVDD.n2985 0.00194
R32137 DVDD.n2720 DVDD.n2703 0.00194
R32138 DVDD.n3805 DVDD.n1685 0.00194
R32139 DVDD.n3807 DVDD.n3806 0.00194
R32140 DVDD.n5402 DVDD.n5401 0.00194
R32141 DVDD.n359 DVDD.n307 0.00194
R32142 DVDD.n4638 DVDD.n909 0.00194
R32143 DVDD.n4720 DVDD.n4719 0.00194
R32144 DVDD.n3060 DVDD.n2996 0.00191
R32145 DVDD.n4220 DVDD.n4177 0.00191
R32146 DVDD.n2087 DVDD.n2086 0.00185
R32147 DVDD.n2352 DVDD.n2094 0.00185
R32148 DVDD.n4225 DVDD.n1724 0.00185
R32149 DVDD.n4226 DVDD.n1722 0.00185
R32150 DVDD.n3969 DVDD.n3925 0.00185
R32151 DVDD.n3389 DVDD.n2737 0.00184
R32152 DVDD.n3005 DVDD.n2701 0.00184
R32153 DVDD.n3707 DVDD.n3706 0.00184
R32154 DVDD.n3389 DVDD.n3388 0.00184
R32155 DVDD.n2761 DVDD.n2701 0.00184
R32156 DVDD.n3707 DVDD.n1907 0.00184
R32157 DVDD.n3389 DVDD.n2743 0.00184
R32158 DVDD.n3287 DVDD.n2701 0.00184
R32159 DVDD.n3707 DVDD.n1903 0.00184
R32160 DVDD.n3390 DVDD.n3389 0.00184
R32161 DVDD.n3415 DVDD.n2701 0.00184
R32162 DVDD.n3707 DVDD.n1899 0.00184
R32163 DVDD.n3055 DVDD.n3008 0.00179
R32164 DVDD.n4159 DVDD.n4158 0.00179
R32165 DVDD.n5417 DVDD.n324 0.00179
R32166 DVDD.n4712 DVDD.n922 0.00179
R32167 DVDD.n5457 DVDD.n5456 0.00174855
R32168 DVDD.n5632 DVDD.n5631 0.00174567
R32169 DVDD.n5550 DVDD.n20 0.00173924
R32170 DVDD.n4667 DVDD.n4649 0.00173924
R32171 DVDD.n4255 DVDD.n1691 0.00173
R32172 DVDD.n4121 DVDD.n4120 0.00173
R32173 DVDD.n4804 DVDD.n732 0.0017
R32174 DVDD.n4874 DVDD.n4873 0.0017
R32175 DVDD.n4883 DVDD.n696 0.0017
R32176 DVDD.n407 DVDD.n399 0.0017
R32177 DVDD.n4287 DVDD.n4286 0.0017
R32178 DVDD.n4104 DVDD.n1790 0.0017
R32179 DVDD.n3975 DVDD.n1818 0.0017
R32180 DVDD.n3977 DVDD.n3976 0.0017
R32181 DVDD.n405 DVDD.n402 0.0017
R32182 DVDD.n4882 DVDD.n4881 0.0017
R32183 DVDD.n4880 DVDD.n704 0.0017
R32184 DVDD.n4772 DVDD.n703 0.0017
R32185 DVDD.n3051 DVDD.n3011 0.00167
R32186 DVDD.n4247 DVDD.n1695 0.00167
R32187 DVDD.n5361 DVDD.n405 0.00167
R32188 DVDD.n5883 DVDD.n108 0.00167
R32189 DVDD.n116 DVDD.n107 0.00167
R32190 DVDD.n5914 DVDD.n5909 0.00167
R32191 DVDD.n4881 DVDD.n695 0.00167
R32192 DVDD.n4880 DVDD.n4879 0.00167
R32193 DVDD.n4775 DVDD.n703 0.00167
R32194 DVDD.n5704 DVDD.n5703 0.00167
R32195 DVDD.n241 DVDD.n227 0.00167
R32196 DVDD.n5706 DVDD.n234 0.00167
R32197 DVDD DVDD.n1741 0.00165261
R32198 DVDD.n1743 DVDD 0.00165261
R32199 DVDD.n1728 DVDD.n1722 0.001625
R32200 DVDD.n4168 DVDD.n1769 0.00161
R32201 DVDD.n5830 DVDD.n163 0.00160656
R32202 DVDD.n5186 DVDD.n468 0.00160656
R32203 DVDD.n4956 DVDD.n4946 0.00160656
R32204 DVDD.n744 DVDD.n742 0.00160656
R32205 DVDD.n4512 DVDD.n4505 0.00160656
R32206 DVDD.n2401 DVDD.n2400 0.00159286
R32207 DVDD.n1999 DVDD.n1997 0.00159286
R32208 DVDD.n2404 DVDD.n2004 0.00159286
R32209 DVDD.n2295 DVDD.n2122 0.00159286
R32210 DVDD.n3667 DVDD.n1982 0.00159286
R32211 DVDD.n3671 DVDD.n1983 0.00159286
R32212 DVDD.n3674 DVDD.n1988 0.00159286
R32213 DVDD.n2442 DVDD.n2438 0.00159286
R32214 DVDD.n3604 DVDD.n3603 0.00159286
R32215 DVDD.n3601 DVDD.n2448 0.00159286
R32216 DVDD.n3510 DVDD.n3451 0.00159286
R32217 DVDD.n3068 DVDD.n2991 0.00155
R32218 DVDD.n5322 DVDD.n449 0.00149
R32219 DVDD.n5321 DVDD.n5320 0.00149
R32220 DVDD.n485 DVDD.n450 0.00149
R32221 DVDD.n5096 DVDD.n571 0.00149
R32222 DVDD.n2641 DVDD.n2451 0.00147826
R32223 DVDD.n1095 DVDD.n357 0.00146
R32224 DVDD.n4442 DVDD.n4441 0.00146
R32225 DVDD.n1094 DVDD.n989 0.00146
R32226 DVDD.n4717 DVDD.n907 0.00146
R32227 DVDD.n5048 DVDD.n481 0.00146
R32228 DVDD.n5247 DVDD.n482 0.00146
R32229 DVDD.n5249 DVDD.n5248 0.00146
R32230 DVDD.n5324 DVDD.n448 0.00146
R32231 DVDD.n4260 DVDD.n1687 0.00146
R32232 DVDD.n4033 DVDD.n1792 0.00146
R32233 DVDD.n4035 DVDD.n4034 0.00146
R32234 DVDD.n5323 DVDD.n5322 0.00146
R32235 DVDD.n5321 DVDD.n451 0.00146
R32236 DVDD.n4838 DVDD.n450 0.00146
R32237 DVDD.n5047 DVDD.n571 0.00146
R32238 DVDD.n1945 DVDD.n1938 0.00143
R32239 DVDD.n1949 DVDD.n1948 0.00143
R32240 DVDD.n1967 DVDD.n1957 0.00143
R32241 DVDD.n3702 DVDD.n3699 0.00143
R32242 DVDD.n5533 DVDD.n12 0.00142943
R32243 DVDD.n4684 DVDD.n979 0.00142943
R32244 DVDD.n2656 DVDD.n2492 0.0014
R32245 DVDD.n3188 DVDD.n3187 0.0014
R32246 DVDD.n3184 DVDD.n3183 0.0014
R32247 DVDD.n3196 DVDD.n3132 0.0014
R32248 DVDD.n3195 DVDD.n2986 0.0014
R32249 DVDD.n3210 DVDD.n3080 0.0014
R32250 DVDD.n4224 DVDD.n4223 0.0014
R32251 DVDD.n5689 DVDD 0.00134
R32252 DVDD.n5972 DVDD 0.00134
R32253 DVDD.n5591 DVDD 0.00134
R32254 DVDD.n5897 DVDD 0.00134
R32255 DVDD.n4197 DVDD 0.00134
R32256 DVDD.n4196 DVDD 0.00134
R32257 DVDD.n2334 DVDD.n2333 0.00133571
R32258 DVDD.n3528 DVDD.n2495 0.00133571
R32259 DVDD.n2670 DVDD.n2500 0.00133571
R32260 DVDD.n3526 DVDD.n3525 0.00133571
R32261 DVDD.n1557 DVDD.n1556 0.00133571
R32262 DVDD.n1554 DVDD.n1218 0.00133571
R32263 DVDD.n3177 DVDD.n3175 0.00131081
R32264 DVDD.n3237 DVDD.n3087 0.00131081
R32265 DVDD.n3405 DVDD.n2725 0.00131
R32266 DVDD.n3406 DVDD.n2724 0.00131
R32267 DVDD.n3411 DVDD.n3409 0.00131
R32268 DVDD.n3410 DVDD.n2706 0.00131
R32269 DVDD.n3418 DVDD.n3417 0.00131
R32270 DVDD.n3424 DVDD.n2703 0.00131
R32271 DVDD.n3423 DVDD.n2704 0.00131
R32272 DVDD.n3431 DVDD.n2698 0.00131
R32273 DVDD.n3432 DVDD.n2696 0.00131
R32274 DVDD.n3435 DVDD.n3434 0.00131
R32275 DVDD.n4141 DVDD.n1712 0.00131
R32276 DVDD.n699 DVDD.n698 0.0013
R32277 DVDD.n4885 DVDD.n4884 0.0013
R32278 DVDD.n731 DVDD.n697 0.0013
R32279 DVDD.n4768 DVDD.n4767 0.0013
R32280 DVDD.n3974 DVDD.n1817 0.0013
R32281 DVDD.n5563 DVDD.n68 0.00127453
R32282 DVDD.n5652 DVDD.n49 0.00127453
R32283 DVDD.n5568 DVDD.n67 0.00127453
R32284 DVDD.n5569 DVDD.n66 0.00127453
R32285 DVDD.n5610 DVDD.n51 0.00127453
R32286 DVDD.n5570 DVDD.n65 0.00127453
R32287 DVDD.n5609 DVDD.n52 0.00127453
R32288 DVDD.n5571 DVDD.n64 0.00127453
R32289 DVDD.n5608 DVDD.n53 0.00127453
R32290 DVDD.n5572 DVDD.n63 0.00127453
R32291 DVDD.n5607 DVDD.n54 0.00127453
R32292 DVDD.n5573 DVDD.n62 0.00127453
R32293 DVDD.n5606 DVDD.n55 0.00127453
R32294 DVDD.n5574 DVDD.n61 0.00127453
R32295 DVDD.n5605 DVDD.n56 0.00127453
R32296 DVDD.n5575 DVDD.n60 0.00127453
R32297 DVDD.n5604 DVDD.n57 0.00127453
R32298 DVDD.n5576 DVDD.n59 0.00127453
R32299 DVDD.n5933 DVDD.n69 0.00127453
R32300 DVDD.n70 DVDD.n48 0.00127453
R32301 DVDD.n270 DVDD.n268 0.00127453
R32302 DVDD.n5478 DVDD.n272 0.00127453
R32303 DVDD.n298 DVDD.n275 0.00127453
R32304 DVDD.n299 DVDD.n276 0.00127453
R32305 DVDD.n315 DVDD.n292 0.00127453
R32306 DVDD.n300 DVDD.n277 0.00127453
R32307 DVDD.n314 DVDD.n291 0.00127453
R32308 DVDD.n301 DVDD.n278 0.00127453
R32309 DVDD.n313 DVDD.n290 0.00127453
R32310 DVDD.n302 DVDD.n279 0.00127453
R32311 DVDD.n312 DVDD.n289 0.00127453
R32312 DVDD.n303 DVDD.n280 0.00127453
R32313 DVDD.n311 DVDD.n288 0.00127453
R32314 DVDD.n304 DVDD.n281 0.00127453
R32315 DVDD.n310 DVDD.n287 0.00127453
R32316 DVDD.n305 DVDD.n282 0.00127453
R32317 DVDD.n309 DVDD.n286 0.00127453
R32318 DVDD.n306 DVDD.n283 0.00127453
R32319 DVDD.n308 DVDD.n285 0.00127453
R32320 DVDD.n5476 DVDD.n5475 0.00127453
R32321 DVDD DVDD.n1740 0.00126841
R32322 DVDD.n3269 DVDD.n2958 0.00125
R32323 DVDD.n3271 DVDD.n3270 0.00125
R32324 DVDD.n3283 DVDD.n2931 0.00125
R32325 DVDD.n3282 DVDD.n2927 0.00125
R32326 DVDD.n3290 DVDD.n3289 0.00125
R32327 DVDD.n3294 DVDD.n3293 0.00125
R32328 DVDD.n3303 DVDD.n2923 0.00125
R32329 DVDD.n3302 DVDD.n2918 0.00125
R32330 DVDD.n3324 DVDD.n3323 0.00125
R32331 DVDD.n3320 DVDD.n2919 0.00125
R32332 DVDD.n2935 DVDD.n2758 0.00125
R32333 DVDD.n2938 DVDD.n2759 0.00125
R32334 DVDD.n2947 DVDD.n2946 0.00125
R32335 DVDD.n2945 DVDD.n2762 0.00125
R32336 DVDD.n3373 DVDD.n3372 0.00125
R32337 DVDD.n2769 DVDD.n2768 0.00125
R32338 DVDD.n3365 DVDD.n3364 0.00125
R32339 DVDD.n2807 DVDD.n2770 0.00125
R32340 DVDD.n2808 DVDD.n2775 0.00125
R32341 DVDD.n2801 DVDD.n2776 0.00125
R32342 DVDD.n5420 DVDD.n103 0.00124896
R32343 DVDD.n2847 DVDD.n2796 0.0012337
R32344 DVDD.n2855 DVDD.n2781 0.0012337
R32345 DVDD.n2881 DVDD.n2869 0.0012337
R32346 DVDD.n2890 DVDD.n2875 0.0012337
R32347 DVDD.n5714 DVDD.n5712 0.00122
R32348 DVDD.n5942 DVDD.n38 0.00122
R32349 DVDD.n5284 DVDD.n44 0.00122
R32350 DVDD.n5877 DVDD.n119 0.00122
R32351 DVDD.n4171 DVDD.n1724 0.00122
R32352 DVDD.n4170 DVDD.n1722 0.00122
R32353 DVDD.n5876 DVDD.n41 0.00122
R32354 DVDD.n5939 DVDD.n42 0.00122
R32355 DVDD.n5941 DVDD.n5940 0.00122
R32356 DVDD.n5713 DVDD.n40 0.00122
R32357 DVDD.n2153 DVDD.n2152 0.00120714
R32358 DVDD.n2277 DVDD.n2160 0.00120714
R32359 DVDD.n3064 DVDD 0.00119767
R32360 DVDD.n3043 DVDD 0.00119767
R32361 DVDD.n2999 DVDD 0.00119767
R32362 DVDD.n3018 DVDD 0.00119767
R32363 DVDD.n1706 DVDD.n1700 0.00119
R32364 DVDD.n4240 DVDD.n1707 0.00119
R32365 DVDD.n478 DVDD.n447 0.00114
R32366 DVDD.n5251 DVDD.n5250 0.00114
R32367 DVDD.n4835 DVDD.n477 0.00114
R32368 DVDD.n5050 DVDD.n5049 0.00114
R32369 DVDD.n4104 DVDD.n1789 0.00114
R32370 DVDD.n3019 DVDD.n3015 0.00113
R32371 DVDD.n5517 DVDD.n27 0.00111962
R32372 DVDD.n4699 DVDD.n4656 0.00111962
R32373 DVDD.n2973 DVDD.n2971 0.00107
R32374 DVDD.n2980 DVDD.n2967 0.00107
R32375 DVDD.n2981 DVDD.n2964 0.00107
R32376 DVDD.n2985 DVDD.n2965 0.00107
R32377 DVDD.n3393 DVDD.n2732 0.00107
R32378 DVDD.n3395 DVDD.n3394 0.00107
R32379 DVDD.n3399 DVDD.n2729 0.00107
R32380 DVDD.n3398 DVDD.n2730 0.00107
R32381 DVDD.n2862 DVDD.n2861 0.00107
R32382 DVDD.n3341 DVDD.n2872 0.00107
R32383 DVDD.n3316 DVDD.n2859 0.00107
R32384 DVDD.n3346 DVDD.n2777 0.00107
R32385 DVDD.n2799 DVDD.n2780 0.00107
R32386 DVDD.n3349 DVDD.n3348 0.00107
R32387 DVDD.n4151 DVDD.n4150 0.00107
R32388 DVDD.n107 DVDD.n77 0.00107
R32389 DVDD.n5914 DVDD.n79 0.00107
R32390 DVDD.n241 DVDD.n224 0.00107
R32391 DVDD.n5707 DVDD.n5706 0.00107
R32392 DVDD.n5896 DVDD 0.00106
R32393 DVDD.n5590 DVDD 0.00106
R32394 DVDD.n5971 DVDD 0.00106
R32395 DVDD.n3059 DVDD.n3001 0.00101
R32396 DVDD.n3777 DVDD.n3736 0.00101
R32397 DVDD.n3754 DVDD.n1856 0.00101
R32398 DVDD.n3780 DVDD.n3779 0.00101
R32399 DVDD.n3998 DVDD.n3997 0.00101
R32400 DVDD.n1181 DVDD.n1120 0.00101
R32401 DVDD.n1579 DVDD.n1121 0.00101
R32402 DVDD.n1582 DVDD.n1131 0.00101
R32403 DVDD.n4413 DVDD.n4412 0.00101
R32404 DVDD.n4400 DVDD.n1108 0.00101
R32405 DVDD.n4417 DVDD.n4416 0.00101
R32406 DVDD.n4375 DVDD.n1595 0.00101
R32407 DVDD.n4385 DVDD.n1596 0.00101
R32408 DVDD.n4388 DVDD.n1607 0.00101
R32409 DVDD.n4332 DVDD.n1627 0.00101
R32410 DVDD.n4342 DVDD.n1628 0.00101
R32411 DVDD.n4345 DVDD.n1639 0.00101
R32412 DVDD.n3337 DVDD 0.00098913
R32413 DVDD.n2646 DVDD.n2443 0.00098913
R32414 DVDD.n5879 DVDD.n5878 0.00098
R32415 DVDD.n5283 DVDD.n35 0.00098
R32416 DVDD.n5944 DVDD.n5943 0.00098
R32417 DVDD.n215 DVDD.n34 0.00098
R32418 DVDD.n4223 DVDD.n4172 0.00098
R32419 DVDD.n5649 DVDD.n50 0.000964716
R32420 DVDD.n5473 DVDD.n316 0.000964716
R32421 DVDD.n2058 DVDD.n2054 0.00095
R32422 DVDD.n2665 DVDD.n2496 0.00095
R32423 DVDD.n3444 DVDD.n3443 0.00095
R32424 DVDD.n5384 DVDD.n5383 0.00095
R32425 DVDD.n5381 DVDD.n379 0.00095
R32426 DVDD.n4562 DVDD.n1075 0.00095
R32427 DVDD.n4499 DVDD.n1073 0.00095
R32428 DVDD.n4621 DVDD.n1005 0.00095
R32429 DVDD.n4618 DVDD.n4617 0.00095
R32430 DVDD.n4744 DVDD.n4743 0.00095
R32431 DVDD.n4746 DVDD.n891 0.00095
R32432 DVDD.n1383 DVDD.n1306 0.000912844
R32433 DVDD.n1321 DVDD.n1220 0.000912844
R32434 DVDD.n3056 DVDD.n3007 0.00089
R32435 DVDD.n4017 DVDD.n4016 0.00089
R32436 DVDD.n5851 DVDD.n137 0.00089
R32437 DVDD.n5858 DVDD.n130 0.00089
R32438 DVDD.n144 DVDD.n143 0.00089
R32439 DVDD.n5836 DVDD.n155 0.00089
R32440 DVDD.n5785 DVDD.n180 0.00089
R32441 DVDD.n537 DVDD.n169 0.00089
R32442 DVDD.n197 DVDD.n196 0.00089
R32443 DVDD.n5735 DVDD.n5729 0.00089
R32444 DVDD.n4130 DVDD.n4129 0.00083
R32445 DVDD.n5650 DVDD.n5649 0.000809811
R32446 DVDD.n5616 DVDD.n5604 0.000809811
R32447 DVDD.n316 DVDD.n293 0.000809811
R32448 DVDD.n5441 DVDD.n286 0.000809811
R32449 DVDD.n5429 DVDD.n325 0.0008
R32450 DVDD.n353 DVDD.n321 0.0008
R32451 DVDD.n4708 DVDD.n943 0.0008
R32452 DVDD.n4710 DVDD.n914 0.0008
R32453 DVDD.n3048 DVDD.n3047 0.00077
R32454 DVDD.n111 DVDD.n90 0.000731959
R32455 DVDD.n5918 DVDD.n102 0.000731959
R32456 DVDD.n5409 DVDD.n344 0.000731959
R32457 DVDD.n5423 DVDD.n349 0.000731959
R32458 DVDD.n937 DVDD.n916 0.000731959
R32459 DVDD.n956 DVDD.n923 0.000731959
R32460 DVDD.n5705 DVDD.n5674 0.000731959
R32461 DVDD.n249 DVDD.n229 0.000731959
R32462 DVDD.n3954 DVDD.n3953 0.00071
R32463 DVDD.n2196 DVDD 0.000671429
R32464 DVDD.n3472 DVDD 0.000671429
R32465 DVDD.n1360 DVDD 0.000671429
R32466 DVDD.n3185 DVDD.n3105 0.00062
R32467 DVDD.n3241 DVDD.n3092 0.00062
R32468 DVDD.n3244 DVDD.n3089 0.00062
R32469 DVDD.n3254 DVDD.n3081 0.00062
R32470 DVDD.n3256 DVDD.n2962 0.00062
R32471 DVDD.n3181 DVDD.n3136 0.00062
R32472 DVDD.n3141 DVDD.n3137 0.00062
R32473 DVDD.n3198 DVDD.n3126 0.00062
R32474 DVDD.n3127 DVDD.n3078 0.00062
R32475 DVDD.n3208 DVDD.n2751 0.00062
R32476 DVDD.n3807 DVDD.n1690 0.00059
R32477 DVDD.n5896 DVDD 0.00058
R32478 DVDD.n5590 DVDD 0.00058
R32479 DVDD.n5971 DVDD 0.00058
R32480 DVDD.n5688 DVDD 0.00058
R32481 DVDD.n4195 DVDD 0.00058
R32482 DVDD.n1368 DVDD.n1337 0.000564286
R32483 DVDD.n1340 DVDD.n1331 0.000564286
R32484 DVDD.n3052 DVDD.n2720 0.00056
R32485 DVDD.n3807 DVDD.n1684 0.00055625
R32486 DVDD.n5343 DVDD.n5342 0.00053
R32487 DVDD.n5340 DVDD.n426 0.00053
R32488 DVDD.n5006 DVDD.n674 0.00053
R32489 DVDD.n4940 DVDD.n672 0.00053
R32490 DVDD.n5014 DVDD.n605 0.00053
R32491 DVDD.n616 DVDD.n603 0.00053
R32492 DVDD.n5023 DVDD.n5022 0.00053
R32493 DVDD.n591 DVDD.n584 0.00053
R32494 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t4 14.2306
R32495 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t3 13.9076
R32496 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t1 11.6919
R32497 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t0 4.40522
R32498 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t2 4.13853
R32499 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.n0 4.13772
R32500 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t4 35.5619
R32501 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t2 35.5619
R32502 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t5 34.9362
R32503 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t3 34.9362
R32504 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.B 6.58393
R32505 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.B GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.n1 4.4005
R32506 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.B GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.n0 4.00161
R32507 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t0 3.08699
R32508 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z 2.76118
R32509 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t3 35.9269
R32510 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t2 30.9212
R32511 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A 23.5268
R32512 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.n0 4.0005
R32513 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t1 3.23447
R32514 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_1.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D.n0 1.15854
R32515 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D.t1 0.5465
R32516 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D.t0 0.5465
R32517 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS 11.0117
R32518 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS.t1 11.0117
R32519 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS.t0 11.0117
R32520 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS.t1 11.0117
R32521 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n6 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t9 79.2576
R32522 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t13 79.2576
R32523 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t3 79.2576
R32524 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t5 79.2576
R32525 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n6 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t6 77.8672
R32526 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t7 77.8672
R32527 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t2 77.8672
R32528 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t12 77.8672
R32529 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t10 37.5434
R32530 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t4 37.5434
R32531 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t8 25.3941
R32532 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t11 25.3941
R32533 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 12.2973
R32534 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n8 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n7 8.47471
R32535 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n0 8.44221
R32536 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n7 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 6.07313
R32537 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 6.07313
R32538 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n8 5.15345
R32539 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n2 5.13701
R32540 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n3 5.13701
R32541 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n4 5.13701
R32542 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n6 5.13701
R32543 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n1 4.34849
R32544 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n8 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 3.78055
R32545 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t0 2.33587
R32546 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 2.08654
R32547 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n7 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n5 2.07524
R32548 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.ndrive_x_<0>.t3 89.2634
R32549 GF_NI_BI_T_BASE_0.ndrive_x_<0>.t0 GF_NI_BI_T_BASE_0.ndrive_x_<0>.n0 7.28458
R32550 GF_NI_BI_T_BASE_0.ndrive_x_<0>.n0 GF_NI_BI_T_BASE_0.ndrive_x_<0>.t2 6.03391
R32551 GF_NI_BI_T_BASE_0.ndrive_x_<0>.n0 GF_NI_BI_T_BASE_0.ndrive_x_<0> 1.45646
R32552 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.ndrive_x_<0>.t0 0.951421
R32553 GF_NI_BI_T_BASE_0.ndrive_x_<0>.t1 GF_NI_BI_T_BASE_0.ndrive_x_<0> 0.773893
R32554 GF_NI_BI_T_BASE_0.ndrive_y_<0> GF_NI_BI_T_BASE_0.ndrive_y_<0>.t5 90.6729
R32555 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n0 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t4 5.90425
R32556 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n1 GF_NI_BI_T_BASE_0.ndrive_y_<0> 3.52102
R32557 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n3 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t3 2.41832
R32558 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n0 GF_NI_BI_T_BASE_0.ndrive_y_<0> 1.5749
R32559 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n4 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n3 1.48076
R32560 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n2 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n1 1.48076
R32561 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n2 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n0 1.09118
R32562 GF_NI_BI_T_BASE_0.ndrive_y_<0> GF_NI_BI_T_BASE_0.ndrive_y_<0>.n4 0.9455
R32563 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n3 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n2 0.578395
R32564 GF_NI_BI_T_BASE_0.ndrive_y_<0> GF_NI_BI_T_BASE_0.ndrive_y_<0>.t2 0.500893
R32565 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n4 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t0 0.360167
R32566 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n1 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t1 0.360167
R32567 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t1 37.5434
R32568 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t2 37.5434
R32569 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t4 29.034
R32570 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t7 28.9248
R32571 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t6 28.9248
R32572 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t12 28.9248
R32573 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t11 28.9248
R32574 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t8 25.3941
R32575 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t9 25.3941
R32576 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t10 24.9104
R32577 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t3 24.8782
R32578 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t5 24.5969
R32579 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 10.2118
R32580 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n2 8.44221
R32581 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n1 5.94601
R32582 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n3 4.40816
R32583 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t0 2.75597
R32584 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314531_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB.t0 2.36868
R32585 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314531_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB.t1 2.08654
R32586 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t10 30.5934
R32587 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t9 30.5934
R32588 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t4 30.5934
R32589 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t2 30.5934
R32590 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t5 29.0913
R32591 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t1 28.7684
R32592 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t12 28.7684
R32593 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t3 28.7684
R32594 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t6 15.5342
R32595 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t11 15.2112
R32596 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t8 14.2306
R32597 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t7 13.9076
R32598 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 13.3452
R32599 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t0 11.0117
R32600 PAD.n6374 PAD.n6373 4.5005
R32601 PAD.n6374 PAD.n5982 4.5005
R32602 PAD.n6374 PAD.n5981 4.5005
R32603 PAD.n6374 PAD.n5980 4.5005
R32604 PAD.n11507 PAD.n11156 4.5005
R32605 PAD.n11302 PAD.n11156 4.5005
R32606 PAD.n11509 PAD.n11156 4.5005
R32607 PAD.n11156 PAD.n11100 4.5005
R32608 PAD.n6373 PAD.n6032 4.5005
R32609 PAD.n6032 PAD.n5981 4.5005
R32610 PAD.n6032 PAD.n5979 4.5005
R32611 PAD.n11507 PAD.n11154 4.5005
R32612 PAD.n11302 PAD.n11154 4.5005
R32613 PAD.n11509 PAD.n11154 4.5005
R32614 PAD.n11507 PAD.n11158 4.5005
R32615 PAD.n11509 PAD.n11158 4.5005
R32616 PAD.n11158 PAD.n11105 4.5005
R32617 PAD.n11507 PAD.n11153 4.5005
R32618 PAD.n11509 PAD.n11153 4.5005
R32619 PAD.n11153 PAD.n11105 4.5005
R32620 PAD.n11507 PAD.n11160 4.5005
R32621 PAD.n11509 PAD.n11160 4.5005
R32622 PAD.n11160 PAD.n11105 4.5005
R32623 PAD.n11507 PAD.n11152 4.5005
R32624 PAD.n11509 PAD.n11152 4.5005
R32625 PAD.n11152 PAD.n11105 4.5005
R32626 PAD.n11507 PAD.n11162 4.5005
R32627 PAD.n11509 PAD.n11162 4.5005
R32628 PAD.n11162 PAD.n11105 4.5005
R32629 PAD.n11507 PAD.n11151 4.5005
R32630 PAD.n11509 PAD.n11151 4.5005
R32631 PAD.n11151 PAD.n11105 4.5005
R32632 PAD.n11507 PAD.n11164 4.5005
R32633 PAD.n11509 PAD.n11164 4.5005
R32634 PAD.n11164 PAD.n11105 4.5005
R32635 PAD.n11507 PAD.n11150 4.5005
R32636 PAD.n11509 PAD.n11150 4.5005
R32637 PAD.n11150 PAD.n11105 4.5005
R32638 PAD.n11507 PAD.n11166 4.5005
R32639 PAD.n11509 PAD.n11166 4.5005
R32640 PAD.n11166 PAD.n11105 4.5005
R32641 PAD.n11507 PAD.n11149 4.5005
R32642 PAD.n11509 PAD.n11149 4.5005
R32643 PAD.n11149 PAD.n11105 4.5005
R32644 PAD.n11507 PAD.n11168 4.5005
R32645 PAD.n11509 PAD.n11168 4.5005
R32646 PAD.n11168 PAD.n11105 4.5005
R32647 PAD.n11507 PAD.n11148 4.5005
R32648 PAD.n11509 PAD.n11148 4.5005
R32649 PAD.n11148 PAD.n11105 4.5005
R32650 PAD.n11507 PAD.n11170 4.5005
R32651 PAD.n11509 PAD.n11170 4.5005
R32652 PAD.n11170 PAD.n11105 4.5005
R32653 PAD.n11507 PAD.n11147 4.5005
R32654 PAD.n11509 PAD.n11147 4.5005
R32655 PAD.n11147 PAD.n11105 4.5005
R32656 PAD.n11507 PAD.n11172 4.5005
R32657 PAD.n11509 PAD.n11172 4.5005
R32658 PAD.n11172 PAD.n11105 4.5005
R32659 PAD.n11507 PAD.n11146 4.5005
R32660 PAD.n11509 PAD.n11146 4.5005
R32661 PAD.n11146 PAD.n11105 4.5005
R32662 PAD.n11507 PAD.n11174 4.5005
R32663 PAD.n11509 PAD.n11174 4.5005
R32664 PAD.n11174 PAD.n11105 4.5005
R32665 PAD.n11507 PAD.n11145 4.5005
R32666 PAD.n11509 PAD.n11145 4.5005
R32667 PAD.n11145 PAD.n11105 4.5005
R32668 PAD.n11507 PAD.n11176 4.5005
R32669 PAD.n11509 PAD.n11176 4.5005
R32670 PAD.n11176 PAD.n11105 4.5005
R32671 PAD.n11507 PAD.n11144 4.5005
R32672 PAD.n11509 PAD.n11144 4.5005
R32673 PAD.n11144 PAD.n11105 4.5005
R32674 PAD.n11507 PAD.n11178 4.5005
R32675 PAD.n11509 PAD.n11178 4.5005
R32676 PAD.n11178 PAD.n11105 4.5005
R32677 PAD.n11507 PAD.n11143 4.5005
R32678 PAD.n11509 PAD.n11143 4.5005
R32679 PAD.n11143 PAD.n11105 4.5005
R32680 PAD.n11507 PAD.n11180 4.5005
R32681 PAD.n11509 PAD.n11180 4.5005
R32682 PAD.n11180 PAD.n11105 4.5005
R32683 PAD.n11507 PAD.n11142 4.5005
R32684 PAD.n11509 PAD.n11142 4.5005
R32685 PAD.n11142 PAD.n11105 4.5005
R32686 PAD.n11507 PAD.n11182 4.5005
R32687 PAD.n11509 PAD.n11182 4.5005
R32688 PAD.n11182 PAD.n11105 4.5005
R32689 PAD.n11507 PAD.n11141 4.5005
R32690 PAD.n11509 PAD.n11141 4.5005
R32691 PAD.n11141 PAD.n11105 4.5005
R32692 PAD.n11507 PAD.n11184 4.5005
R32693 PAD.n11509 PAD.n11184 4.5005
R32694 PAD.n11184 PAD.n11105 4.5005
R32695 PAD.n11507 PAD.n11140 4.5005
R32696 PAD.n11509 PAD.n11140 4.5005
R32697 PAD.n11140 PAD.n11105 4.5005
R32698 PAD.n11507 PAD.n11186 4.5005
R32699 PAD.n11509 PAD.n11186 4.5005
R32700 PAD.n11186 PAD.n11105 4.5005
R32701 PAD.n11507 PAD.n11139 4.5005
R32702 PAD.n11509 PAD.n11139 4.5005
R32703 PAD.n11139 PAD.n11105 4.5005
R32704 PAD.n11507 PAD.n11188 4.5005
R32705 PAD.n11509 PAD.n11188 4.5005
R32706 PAD.n11188 PAD.n11105 4.5005
R32707 PAD.n11507 PAD.n11138 4.5005
R32708 PAD.n11509 PAD.n11138 4.5005
R32709 PAD.n11138 PAD.n11105 4.5005
R32710 PAD.n11507 PAD.n11190 4.5005
R32711 PAD.n11509 PAD.n11190 4.5005
R32712 PAD.n11190 PAD.n11105 4.5005
R32713 PAD.n11507 PAD.n11137 4.5005
R32714 PAD.n11509 PAD.n11137 4.5005
R32715 PAD.n11137 PAD.n11105 4.5005
R32716 PAD.n11507 PAD.n11192 4.5005
R32717 PAD.n11509 PAD.n11192 4.5005
R32718 PAD.n11192 PAD.n11105 4.5005
R32719 PAD.n11507 PAD.n11136 4.5005
R32720 PAD.n11509 PAD.n11136 4.5005
R32721 PAD.n11136 PAD.n11105 4.5005
R32722 PAD.n11507 PAD.n11194 4.5005
R32723 PAD.n11509 PAD.n11194 4.5005
R32724 PAD.n11194 PAD.n11105 4.5005
R32725 PAD.n11507 PAD.n11135 4.5005
R32726 PAD.n11509 PAD.n11135 4.5005
R32727 PAD.n11135 PAD.n11105 4.5005
R32728 PAD.n11507 PAD.n11196 4.5005
R32729 PAD.n11509 PAD.n11196 4.5005
R32730 PAD.n11196 PAD.n11105 4.5005
R32731 PAD.n11507 PAD.n11134 4.5005
R32732 PAD.n11509 PAD.n11134 4.5005
R32733 PAD.n11134 PAD.n11105 4.5005
R32734 PAD.n11507 PAD.n11198 4.5005
R32735 PAD.n11509 PAD.n11198 4.5005
R32736 PAD.n11198 PAD.n11105 4.5005
R32737 PAD.n11507 PAD.n11133 4.5005
R32738 PAD.n11509 PAD.n11133 4.5005
R32739 PAD.n11133 PAD.n11105 4.5005
R32740 PAD.n11507 PAD.n11200 4.5005
R32741 PAD.n11509 PAD.n11200 4.5005
R32742 PAD.n11200 PAD.n11105 4.5005
R32743 PAD.n11507 PAD.n11132 4.5005
R32744 PAD.n11509 PAD.n11132 4.5005
R32745 PAD.n11132 PAD.n11105 4.5005
R32746 PAD.n11507 PAD.n11202 4.5005
R32747 PAD.n11509 PAD.n11202 4.5005
R32748 PAD.n11202 PAD.n11105 4.5005
R32749 PAD.n11507 PAD.n11131 4.5005
R32750 PAD.n11509 PAD.n11131 4.5005
R32751 PAD.n11131 PAD.n11105 4.5005
R32752 PAD.n11507 PAD.n11204 4.5005
R32753 PAD.n11509 PAD.n11204 4.5005
R32754 PAD.n11204 PAD.n11105 4.5005
R32755 PAD.n11507 PAD.n11130 4.5005
R32756 PAD.n11509 PAD.n11130 4.5005
R32757 PAD.n11130 PAD.n11105 4.5005
R32758 PAD.n11507 PAD.n11206 4.5005
R32759 PAD.n11509 PAD.n11206 4.5005
R32760 PAD.n11206 PAD.n11105 4.5005
R32761 PAD.n11507 PAD.n11129 4.5005
R32762 PAD.n11509 PAD.n11129 4.5005
R32763 PAD.n11129 PAD.n11105 4.5005
R32764 PAD.n11507 PAD.n11208 4.5005
R32765 PAD.n11509 PAD.n11208 4.5005
R32766 PAD.n11208 PAD.n11105 4.5005
R32767 PAD.n11507 PAD.n11128 4.5005
R32768 PAD.n11509 PAD.n11128 4.5005
R32769 PAD.n11128 PAD.n11105 4.5005
R32770 PAD.n11507 PAD.n11210 4.5005
R32771 PAD.n11509 PAD.n11210 4.5005
R32772 PAD.n11210 PAD.n11105 4.5005
R32773 PAD.n11507 PAD.n11127 4.5005
R32774 PAD.n11509 PAD.n11127 4.5005
R32775 PAD.n11127 PAD.n11105 4.5005
R32776 PAD.n11507 PAD.n11212 4.5005
R32777 PAD.n11509 PAD.n11212 4.5005
R32778 PAD.n11212 PAD.n11105 4.5005
R32779 PAD.n11507 PAD.n11126 4.5005
R32780 PAD.n11509 PAD.n11126 4.5005
R32781 PAD.n11126 PAD.n11105 4.5005
R32782 PAD.n11507 PAD.n11214 4.5005
R32783 PAD.n11509 PAD.n11214 4.5005
R32784 PAD.n11214 PAD.n11105 4.5005
R32785 PAD.n11507 PAD.n11125 4.5005
R32786 PAD.n11509 PAD.n11125 4.5005
R32787 PAD.n11125 PAD.n11105 4.5005
R32788 PAD.n11507 PAD.n11216 4.5005
R32789 PAD.n11509 PAD.n11216 4.5005
R32790 PAD.n11216 PAD.n11105 4.5005
R32791 PAD.n11507 PAD.n11124 4.5005
R32792 PAD.n11509 PAD.n11124 4.5005
R32793 PAD.n11124 PAD.n11105 4.5005
R32794 PAD.n11507 PAD.n11218 4.5005
R32795 PAD.n11509 PAD.n11218 4.5005
R32796 PAD.n11218 PAD.n11105 4.5005
R32797 PAD.n11507 PAD.n11123 4.5005
R32798 PAD.n11509 PAD.n11123 4.5005
R32799 PAD.n11123 PAD.n11105 4.5005
R32800 PAD.n11507 PAD.n11220 4.5005
R32801 PAD.n11509 PAD.n11220 4.5005
R32802 PAD.n11220 PAD.n11105 4.5005
R32803 PAD.n11507 PAD.n11122 4.5005
R32804 PAD.n11509 PAD.n11122 4.5005
R32805 PAD.n11122 PAD.n11105 4.5005
R32806 PAD.n11507 PAD.n11222 4.5005
R32807 PAD.n11509 PAD.n11222 4.5005
R32808 PAD.n11222 PAD.n11105 4.5005
R32809 PAD.n11507 PAD.n11121 4.5005
R32810 PAD.n11509 PAD.n11121 4.5005
R32811 PAD.n11121 PAD.n11105 4.5005
R32812 PAD.n11507 PAD.n11224 4.5005
R32813 PAD.n11509 PAD.n11224 4.5005
R32814 PAD.n11224 PAD.n11105 4.5005
R32815 PAD.n11507 PAD.n11120 4.5005
R32816 PAD.n11509 PAD.n11120 4.5005
R32817 PAD.n11120 PAD.n11105 4.5005
R32818 PAD.n11507 PAD.n11226 4.5005
R32819 PAD.n11509 PAD.n11226 4.5005
R32820 PAD.n11226 PAD.n11105 4.5005
R32821 PAD.n11507 PAD.n11119 4.5005
R32822 PAD.n11509 PAD.n11119 4.5005
R32823 PAD.n11119 PAD.n11105 4.5005
R32824 PAD.n11507 PAD.n11228 4.5005
R32825 PAD.n11509 PAD.n11228 4.5005
R32826 PAD.n11228 PAD.n11105 4.5005
R32827 PAD.n11507 PAD.n11118 4.5005
R32828 PAD.n11509 PAD.n11118 4.5005
R32829 PAD.n11118 PAD.n11105 4.5005
R32830 PAD.n11507 PAD.n11230 4.5005
R32831 PAD.n11509 PAD.n11230 4.5005
R32832 PAD.n11230 PAD.n11105 4.5005
R32833 PAD.n11507 PAD.n11117 4.5005
R32834 PAD.n11509 PAD.n11117 4.5005
R32835 PAD.n11117 PAD.n11105 4.5005
R32836 PAD.n11507 PAD.n11232 4.5005
R32837 PAD.n11509 PAD.n11232 4.5005
R32838 PAD.n11232 PAD.n11105 4.5005
R32839 PAD.n11507 PAD.n11116 4.5005
R32840 PAD.n11509 PAD.n11116 4.5005
R32841 PAD.n11116 PAD.n11105 4.5005
R32842 PAD.n11507 PAD.n11234 4.5005
R32843 PAD.n11509 PAD.n11234 4.5005
R32844 PAD.n11234 PAD.n11105 4.5005
R32845 PAD.n11507 PAD.n11115 4.5005
R32846 PAD.n11509 PAD.n11115 4.5005
R32847 PAD.n11115 PAD.n11105 4.5005
R32848 PAD.n11507 PAD.n11236 4.5005
R32849 PAD.n11509 PAD.n11236 4.5005
R32850 PAD.n11236 PAD.n11105 4.5005
R32851 PAD.n11507 PAD.n11114 4.5005
R32852 PAD.n11509 PAD.n11114 4.5005
R32853 PAD.n11114 PAD.n11105 4.5005
R32854 PAD.n11507 PAD.n11238 4.5005
R32855 PAD.n11509 PAD.n11238 4.5005
R32856 PAD.n11238 PAD.n11105 4.5005
R32857 PAD.n11507 PAD.n11113 4.5005
R32858 PAD.n11509 PAD.n11113 4.5005
R32859 PAD.n11113 PAD.n11105 4.5005
R32860 PAD.n11507 PAD.n11240 4.5005
R32861 PAD.n11509 PAD.n11240 4.5005
R32862 PAD.n11240 PAD.n11105 4.5005
R32863 PAD.n11507 PAD.n11112 4.5005
R32864 PAD.n11509 PAD.n11112 4.5005
R32865 PAD.n11112 PAD.n11105 4.5005
R32866 PAD.n11507 PAD.n11242 4.5005
R32867 PAD.n11509 PAD.n11242 4.5005
R32868 PAD.n11242 PAD.n11105 4.5005
R32869 PAD.n11507 PAD.n11111 4.5005
R32870 PAD.n11509 PAD.n11111 4.5005
R32871 PAD.n11111 PAD.n11105 4.5005
R32872 PAD.n11507 PAD.n11244 4.5005
R32873 PAD.n11509 PAD.n11244 4.5005
R32874 PAD.n11244 PAD.n11105 4.5005
R32875 PAD.n11507 PAD.n11110 4.5005
R32876 PAD.n11509 PAD.n11110 4.5005
R32877 PAD.n11110 PAD.n11105 4.5005
R32878 PAD.n11507 PAD.n11246 4.5005
R32879 PAD.n11509 PAD.n11246 4.5005
R32880 PAD.n11246 PAD.n11105 4.5005
R32881 PAD.n11507 PAD.n11109 4.5005
R32882 PAD.n11509 PAD.n11109 4.5005
R32883 PAD.n11109 PAD.n11105 4.5005
R32884 PAD.n11507 PAD.n11248 4.5005
R32885 PAD.n11509 PAD.n11248 4.5005
R32886 PAD.n11248 PAD.n11105 4.5005
R32887 PAD.n11507 PAD.n11108 4.5005
R32888 PAD.n11509 PAD.n11108 4.5005
R32889 PAD.n11108 PAD.n11105 4.5005
R32890 PAD.n11507 PAD.n11250 4.5005
R32891 PAD.n11509 PAD.n11250 4.5005
R32892 PAD.n11250 PAD.n11105 4.5005
R32893 PAD.n11507 PAD.n11107 4.5005
R32894 PAD.n11509 PAD.n11107 4.5005
R32895 PAD.n11107 PAD.n11105 4.5005
R32896 PAD.n11507 PAD.n11252 4.5005
R32897 PAD.n11509 PAD.n11252 4.5005
R32898 PAD.n11252 PAD.n11105 4.5005
R32899 PAD.n11507 PAD.n11106 4.5005
R32900 PAD.n11509 PAD.n11106 4.5005
R32901 PAD.n11106 PAD.n11100 4.5005
R32902 PAD.n11106 PAD.n11105 4.5005
R32903 PAD.n5969 PAD.n5963 4.5005
R32904 PAD.n5969 PAD.n5964 4.5005
R32905 PAD.n5969 PAD.n5962 4.5005
R32906 PAD.n5969 PAD.n5965 4.5005
R32907 PAD.n6386 PAD.n5969 4.5005
R32908 PAD.n11104 PAD.n11096 4.5005
R32909 PAD.n11104 PAD.n11099 4.5005
R32910 PAD.n11513 PAD.n11104 4.5005
R32911 PAD.n6387 PAD.n5963 4.5005
R32912 PAD.n6387 PAD.n5964 4.5005
R32913 PAD.n6387 PAD.n5962 4.5005
R32914 PAD.n6387 PAD.n5965 4.5005
R32915 PAD.n6387 PAD.n6386 4.5005
R32916 PAD.n11514 PAD.n11097 4.5005
R32917 PAD.n11514 PAD.n11098 4.5005
R32918 PAD.n11514 PAD.n11096 4.5005
R32919 PAD.n11514 PAD.n11099 4.5005
R32920 PAD.n11514 PAD.n11513 4.5005
R32921 PAD.n5968 PAD.n5963 4.5005
R32922 PAD.n5968 PAD.n5964 4.5005
R32923 PAD.n5968 PAD.n5962 4.5005
R32924 PAD.n5968 PAD.n5965 4.5005
R32925 PAD.n6386 PAD.n5968 4.5005
R32926 PAD.n11102 PAD.n11097 4.5005
R32927 PAD.n11102 PAD.n11098 4.5005
R32928 PAD.n11102 PAD.n11096 4.5005
R32929 PAD.n11102 PAD.n11099 4.5005
R32930 PAD.n11513 PAD.n11102 4.5005
R32931 PAD.n6385 PAD.n5963 4.5005
R32932 PAD.n6385 PAD.n5964 4.5005
R32933 PAD.n6385 PAD.n5962 4.5005
R32934 PAD.n6385 PAD.n5965 4.5005
R32935 PAD.n6386 PAD.n6385 4.5005
R32936 PAD.n11512 PAD.n11097 4.5005
R32937 PAD.n11512 PAD.n11098 4.5005
R32938 PAD.n11512 PAD.n11096 4.5005
R32939 PAD.n11512 PAD.n11099 4.5005
R32940 PAD.n11513 PAD.n11512 4.5005
R32941 PAD.n11085 PAD.n21 4.5005
R32942 PAD.n10837 PAD.n21 4.5005
R32943 PAD.n367 PAD.n74 4.5005
R32944 PAD.n367 PAD.n366 4.5005
R32945 PAD.n10716 PAD.n415 4.5005
R32946 PAD.n10716 PAD.n10715 4.5005
R32947 PAD.n523 PAD.n435 4.5005
R32948 PAD.n770 PAD.n435 4.5005
R32949 PAD.n10388 PAD.n824 4.5005
R32950 PAD.n10388 PAD.n10387 4.5005
R32951 PAD.n10106 PAD.n1132 4.5005
R32952 PAD.n10353 PAD.n1132 4.5005
R32953 PAD.n1481 PAD.n1140 4.5005
R32954 PAD.n1294 PAD.n1140 4.5005
R32955 PAD.n9998 PAD.n1531 4.5005
R32956 PAD.n9998 PAD.n9997 4.5005
R32957 PAD.n1599 PAD.n1594 4.5005
R32958 PAD.n1685 PAD.n1594 4.5005
R32959 PAD.n9712 PAD.n1984 4.5005
R32960 PAD.n9712 PAD.n9711 4.5005
R32961 PAD.n9445 PAD.n2088 4.5005
R32962 PAD.n9445 PAD.n9444 4.5005
R32963 PAD.n2151 PAD.n2139 4.5005
R32964 PAD.n2236 PAD.n2139 4.5005
R32965 PAD.n2498 PAD.n2487 4.5005
R32966 PAD.n2583 PAD.n2487 4.5005
R32967 PAD.n9140 PAD.n2876 4.5005
R32968 PAD.n9140 PAD.n9139 4.5005
R32969 PAD.n8819 PAD.n2891 4.5005
R32970 PAD.n8570 PAD.n2891 4.5005
R32971 PAD.n8517 PAD.n2994 4.5005
R32972 PAD.n8517 PAD.n8516 4.5005
R32973 PAD.n8492 PAD.n3338 4.5005
R32974 PAD.n8492 PAD.n8491 4.5005
R32975 PAD.n8468 PAD.n3683 4.5005
R32976 PAD.n8468 PAD.n8467 4.5005
R32977 PAD.n8444 PAD.n4025 4.5005
R32978 PAD.n8444 PAD.n8443 4.5005
R32979 PAD.n4420 PAD.n4333 4.5005
R32980 PAD.n4667 PAD.n4333 4.5005
R32981 PAD.n8395 PAD.n4673 4.5005
R32982 PAD.n4832 PAD.n4673 4.5005
R32983 PAD.n4847 PAD.n4843 4.5005
R32984 PAD.n4932 PAD.n4843 4.5005
R32985 PAD.n8161 PAD.n5183 4.5005
R32986 PAD.n7971 PAD.n5183 4.5005
R32987 PAD.n5211 PAD.n5197 4.5005
R32988 PAD.n5296 PAD.n5197 4.5005
R32989 PAD.n7518 PAD.n7207 4.5005
R32990 PAD.n7269 PAD.n7207 4.5005
R32991 PAD.n7780 PAD.n7105 4.5005
R32992 PAD.n7531 PAD.n7105 4.5005
R32993 PAD.n6719 PAD.n6713 4.5005
R32994 PAD.n6804 PAD.n6713 4.5005
R32995 PAD.n5892 PAD.n5551 4.5005
R32996 PAD.n5702 PAD.n5551 4.5005
R32997 PAD.n6690 PAD.n6689 4.5005
R32998 PAD.n6689 PAD.n6688 4.5005
R32999 PAD.n6034 PAD.n5979 4.5005
R33000 PAD.n6034 PAD.n5980 4.5005
R33001 PAD.n6034 PAD.n5981 4.5005
R33002 PAD.n6373 PAD.n6034 4.5005
R33003 PAD.n6030 PAD.n5979 4.5005
R33004 PAD.n6030 PAD.n5981 4.5005
R33005 PAD.n6373 PAD.n6030 4.5005
R33006 PAD.n6037 PAD.n5979 4.5005
R33007 PAD.n6037 PAD.n5981 4.5005
R33008 PAD.n6373 PAD.n6037 4.5005
R33009 PAD.n6029 PAD.n5979 4.5005
R33010 PAD.n6029 PAD.n5981 4.5005
R33011 PAD.n6373 PAD.n6029 4.5005
R33012 PAD.n6040 PAD.n5979 4.5005
R33013 PAD.n6040 PAD.n5981 4.5005
R33014 PAD.n6373 PAD.n6040 4.5005
R33015 PAD.n6028 PAD.n5979 4.5005
R33016 PAD.n6028 PAD.n5981 4.5005
R33017 PAD.n6373 PAD.n6028 4.5005
R33018 PAD.n6043 PAD.n5979 4.5005
R33019 PAD.n6043 PAD.n5981 4.5005
R33020 PAD.n6373 PAD.n6043 4.5005
R33021 PAD.n6027 PAD.n5979 4.5005
R33022 PAD.n6027 PAD.n5981 4.5005
R33023 PAD.n6373 PAD.n6027 4.5005
R33024 PAD.n6046 PAD.n5979 4.5005
R33025 PAD.n6046 PAD.n5981 4.5005
R33026 PAD.n6373 PAD.n6046 4.5005
R33027 PAD.n6026 PAD.n5979 4.5005
R33028 PAD.n6026 PAD.n5981 4.5005
R33029 PAD.n6373 PAD.n6026 4.5005
R33030 PAD.n6049 PAD.n5979 4.5005
R33031 PAD.n6049 PAD.n5981 4.5005
R33032 PAD.n6373 PAD.n6049 4.5005
R33033 PAD.n6025 PAD.n5979 4.5005
R33034 PAD.n6025 PAD.n5981 4.5005
R33035 PAD.n6373 PAD.n6025 4.5005
R33036 PAD.n6052 PAD.n5979 4.5005
R33037 PAD.n6052 PAD.n5981 4.5005
R33038 PAD.n6373 PAD.n6052 4.5005
R33039 PAD.n6024 PAD.n5979 4.5005
R33040 PAD.n6024 PAD.n5981 4.5005
R33041 PAD.n6373 PAD.n6024 4.5005
R33042 PAD.n6055 PAD.n5979 4.5005
R33043 PAD.n6055 PAD.n5981 4.5005
R33044 PAD.n6373 PAD.n6055 4.5005
R33045 PAD.n6023 PAD.n5979 4.5005
R33046 PAD.n6023 PAD.n5981 4.5005
R33047 PAD.n6373 PAD.n6023 4.5005
R33048 PAD.n6058 PAD.n5979 4.5005
R33049 PAD.n6058 PAD.n5981 4.5005
R33050 PAD.n6373 PAD.n6058 4.5005
R33051 PAD.n6022 PAD.n5979 4.5005
R33052 PAD.n6022 PAD.n5981 4.5005
R33053 PAD.n6373 PAD.n6022 4.5005
R33054 PAD.n6061 PAD.n5979 4.5005
R33055 PAD.n6061 PAD.n5981 4.5005
R33056 PAD.n6373 PAD.n6061 4.5005
R33057 PAD.n6021 PAD.n5979 4.5005
R33058 PAD.n6021 PAD.n5981 4.5005
R33059 PAD.n6373 PAD.n6021 4.5005
R33060 PAD.n6064 PAD.n5979 4.5005
R33061 PAD.n6064 PAD.n5981 4.5005
R33062 PAD.n6373 PAD.n6064 4.5005
R33063 PAD.n6020 PAD.n5979 4.5005
R33064 PAD.n6020 PAD.n5981 4.5005
R33065 PAD.n6373 PAD.n6020 4.5005
R33066 PAD.n6067 PAD.n5979 4.5005
R33067 PAD.n6067 PAD.n5981 4.5005
R33068 PAD.n6373 PAD.n6067 4.5005
R33069 PAD.n6019 PAD.n5979 4.5005
R33070 PAD.n6019 PAD.n5981 4.5005
R33071 PAD.n6373 PAD.n6019 4.5005
R33072 PAD.n6070 PAD.n5979 4.5005
R33073 PAD.n6070 PAD.n5981 4.5005
R33074 PAD.n6373 PAD.n6070 4.5005
R33075 PAD.n6018 PAD.n5979 4.5005
R33076 PAD.n6018 PAD.n5981 4.5005
R33077 PAD.n6373 PAD.n6018 4.5005
R33078 PAD.n6073 PAD.n5979 4.5005
R33079 PAD.n6073 PAD.n5981 4.5005
R33080 PAD.n6373 PAD.n6073 4.5005
R33081 PAD.n6017 PAD.n5979 4.5005
R33082 PAD.n6017 PAD.n5981 4.5005
R33083 PAD.n6373 PAD.n6017 4.5005
R33084 PAD.n6076 PAD.n5979 4.5005
R33085 PAD.n6076 PAD.n5981 4.5005
R33086 PAD.n6373 PAD.n6076 4.5005
R33087 PAD.n6016 PAD.n5979 4.5005
R33088 PAD.n6016 PAD.n5981 4.5005
R33089 PAD.n6373 PAD.n6016 4.5005
R33090 PAD.n6079 PAD.n5979 4.5005
R33091 PAD.n6079 PAD.n5981 4.5005
R33092 PAD.n6373 PAD.n6079 4.5005
R33093 PAD.n6015 PAD.n5979 4.5005
R33094 PAD.n6015 PAD.n5981 4.5005
R33095 PAD.n6373 PAD.n6015 4.5005
R33096 PAD.n6082 PAD.n5979 4.5005
R33097 PAD.n6082 PAD.n5981 4.5005
R33098 PAD.n6373 PAD.n6082 4.5005
R33099 PAD.n6014 PAD.n5979 4.5005
R33100 PAD.n6014 PAD.n5981 4.5005
R33101 PAD.n6373 PAD.n6014 4.5005
R33102 PAD.n6085 PAD.n5979 4.5005
R33103 PAD.n6085 PAD.n5981 4.5005
R33104 PAD.n6373 PAD.n6085 4.5005
R33105 PAD.n6013 PAD.n5979 4.5005
R33106 PAD.n6013 PAD.n5981 4.5005
R33107 PAD.n6373 PAD.n6013 4.5005
R33108 PAD.n6088 PAD.n5979 4.5005
R33109 PAD.n6088 PAD.n5981 4.5005
R33110 PAD.n6373 PAD.n6088 4.5005
R33111 PAD.n6012 PAD.n5979 4.5005
R33112 PAD.n6012 PAD.n5981 4.5005
R33113 PAD.n6373 PAD.n6012 4.5005
R33114 PAD.n6091 PAD.n5979 4.5005
R33115 PAD.n6091 PAD.n5981 4.5005
R33116 PAD.n6373 PAD.n6091 4.5005
R33117 PAD.n6011 PAD.n5979 4.5005
R33118 PAD.n6011 PAD.n5981 4.5005
R33119 PAD.n6373 PAD.n6011 4.5005
R33120 PAD.n6094 PAD.n5979 4.5005
R33121 PAD.n6094 PAD.n5981 4.5005
R33122 PAD.n6373 PAD.n6094 4.5005
R33123 PAD.n6010 PAD.n5979 4.5005
R33124 PAD.n6010 PAD.n5981 4.5005
R33125 PAD.n6373 PAD.n6010 4.5005
R33126 PAD.n6097 PAD.n5979 4.5005
R33127 PAD.n6097 PAD.n5981 4.5005
R33128 PAD.n6373 PAD.n6097 4.5005
R33129 PAD.n6009 PAD.n5979 4.5005
R33130 PAD.n6009 PAD.n5981 4.5005
R33131 PAD.n6373 PAD.n6009 4.5005
R33132 PAD.n6100 PAD.n5979 4.5005
R33133 PAD.n6100 PAD.n5981 4.5005
R33134 PAD.n6373 PAD.n6100 4.5005
R33135 PAD.n6008 PAD.n5979 4.5005
R33136 PAD.n6008 PAD.n5981 4.5005
R33137 PAD.n6373 PAD.n6008 4.5005
R33138 PAD.n6103 PAD.n5979 4.5005
R33139 PAD.n6103 PAD.n5981 4.5005
R33140 PAD.n6373 PAD.n6103 4.5005
R33141 PAD.n6007 PAD.n5979 4.5005
R33142 PAD.n6007 PAD.n5981 4.5005
R33143 PAD.n6373 PAD.n6007 4.5005
R33144 PAD.n6106 PAD.n5979 4.5005
R33145 PAD.n6106 PAD.n5981 4.5005
R33146 PAD.n6373 PAD.n6106 4.5005
R33147 PAD.n6006 PAD.n5979 4.5005
R33148 PAD.n6006 PAD.n5981 4.5005
R33149 PAD.n6373 PAD.n6006 4.5005
R33150 PAD.n6109 PAD.n5979 4.5005
R33151 PAD.n6109 PAD.n5981 4.5005
R33152 PAD.n6373 PAD.n6109 4.5005
R33153 PAD.n6005 PAD.n5979 4.5005
R33154 PAD.n6005 PAD.n5981 4.5005
R33155 PAD.n6373 PAD.n6005 4.5005
R33156 PAD.n6112 PAD.n5979 4.5005
R33157 PAD.n6112 PAD.n5981 4.5005
R33158 PAD.n6373 PAD.n6112 4.5005
R33159 PAD.n6004 PAD.n5979 4.5005
R33160 PAD.n6004 PAD.n5981 4.5005
R33161 PAD.n6373 PAD.n6004 4.5005
R33162 PAD.n6115 PAD.n5979 4.5005
R33163 PAD.n6115 PAD.n5981 4.5005
R33164 PAD.n6373 PAD.n6115 4.5005
R33165 PAD.n6003 PAD.n5979 4.5005
R33166 PAD.n6003 PAD.n5981 4.5005
R33167 PAD.n6373 PAD.n6003 4.5005
R33168 PAD.n6118 PAD.n5979 4.5005
R33169 PAD.n6118 PAD.n5981 4.5005
R33170 PAD.n6373 PAD.n6118 4.5005
R33171 PAD.n6002 PAD.n5979 4.5005
R33172 PAD.n6002 PAD.n5981 4.5005
R33173 PAD.n6373 PAD.n6002 4.5005
R33174 PAD.n6121 PAD.n5979 4.5005
R33175 PAD.n6121 PAD.n5981 4.5005
R33176 PAD.n6373 PAD.n6121 4.5005
R33177 PAD.n6001 PAD.n5979 4.5005
R33178 PAD.n6001 PAD.n5981 4.5005
R33179 PAD.n6373 PAD.n6001 4.5005
R33180 PAD.n6124 PAD.n5979 4.5005
R33181 PAD.n6124 PAD.n5981 4.5005
R33182 PAD.n6373 PAD.n6124 4.5005
R33183 PAD.n6000 PAD.n5979 4.5005
R33184 PAD.n6000 PAD.n5981 4.5005
R33185 PAD.n6373 PAD.n6000 4.5005
R33186 PAD.n6127 PAD.n5979 4.5005
R33187 PAD.n6127 PAD.n5981 4.5005
R33188 PAD.n6373 PAD.n6127 4.5005
R33189 PAD.n5999 PAD.n5979 4.5005
R33190 PAD.n5999 PAD.n5981 4.5005
R33191 PAD.n6373 PAD.n5999 4.5005
R33192 PAD.n6130 PAD.n5979 4.5005
R33193 PAD.n6130 PAD.n5981 4.5005
R33194 PAD.n6373 PAD.n6130 4.5005
R33195 PAD.n5998 PAD.n5979 4.5005
R33196 PAD.n5998 PAD.n5981 4.5005
R33197 PAD.n6373 PAD.n5998 4.5005
R33198 PAD.n6133 PAD.n5979 4.5005
R33199 PAD.n6133 PAD.n5981 4.5005
R33200 PAD.n6373 PAD.n6133 4.5005
R33201 PAD.n5997 PAD.n5979 4.5005
R33202 PAD.n5997 PAD.n5981 4.5005
R33203 PAD.n6373 PAD.n5997 4.5005
R33204 PAD.n6136 PAD.n5979 4.5005
R33205 PAD.n6136 PAD.n5981 4.5005
R33206 PAD.n6373 PAD.n6136 4.5005
R33207 PAD.n5996 PAD.n5979 4.5005
R33208 PAD.n5996 PAD.n5981 4.5005
R33209 PAD.n6373 PAD.n5996 4.5005
R33210 PAD.n6139 PAD.n5979 4.5005
R33211 PAD.n6139 PAD.n5981 4.5005
R33212 PAD.n6373 PAD.n6139 4.5005
R33213 PAD.n5995 PAD.n5979 4.5005
R33214 PAD.n5995 PAD.n5981 4.5005
R33215 PAD.n6373 PAD.n5995 4.5005
R33216 PAD.n6142 PAD.n5979 4.5005
R33217 PAD.n6142 PAD.n5981 4.5005
R33218 PAD.n6373 PAD.n6142 4.5005
R33219 PAD.n5994 PAD.n5979 4.5005
R33220 PAD.n5994 PAD.n5981 4.5005
R33221 PAD.n6373 PAD.n5994 4.5005
R33222 PAD.n6145 PAD.n5979 4.5005
R33223 PAD.n6145 PAD.n5981 4.5005
R33224 PAD.n6373 PAD.n6145 4.5005
R33225 PAD.n5993 PAD.n5979 4.5005
R33226 PAD.n5993 PAD.n5981 4.5005
R33227 PAD.n6373 PAD.n5993 4.5005
R33228 PAD.n6148 PAD.n5979 4.5005
R33229 PAD.n6148 PAD.n5981 4.5005
R33230 PAD.n6373 PAD.n6148 4.5005
R33231 PAD.n5992 PAD.n5979 4.5005
R33232 PAD.n5992 PAD.n5981 4.5005
R33233 PAD.n6373 PAD.n5992 4.5005
R33234 PAD.n6151 PAD.n5979 4.5005
R33235 PAD.n6151 PAD.n5981 4.5005
R33236 PAD.n6373 PAD.n6151 4.5005
R33237 PAD.n5991 PAD.n5979 4.5005
R33238 PAD.n5991 PAD.n5981 4.5005
R33239 PAD.n6373 PAD.n5991 4.5005
R33240 PAD.n6154 PAD.n5979 4.5005
R33241 PAD.n6154 PAD.n5981 4.5005
R33242 PAD.n6373 PAD.n6154 4.5005
R33243 PAD.n5990 PAD.n5979 4.5005
R33244 PAD.n5990 PAD.n5981 4.5005
R33245 PAD.n6373 PAD.n5990 4.5005
R33246 PAD.n6157 PAD.n5979 4.5005
R33247 PAD.n6157 PAD.n5981 4.5005
R33248 PAD.n6373 PAD.n6157 4.5005
R33249 PAD.n5989 PAD.n5979 4.5005
R33250 PAD.n5989 PAD.n5981 4.5005
R33251 PAD.n6373 PAD.n5989 4.5005
R33252 PAD.n6160 PAD.n5979 4.5005
R33253 PAD.n6160 PAD.n5981 4.5005
R33254 PAD.n6373 PAD.n6160 4.5005
R33255 PAD.n5988 PAD.n5979 4.5005
R33256 PAD.n5988 PAD.n5981 4.5005
R33257 PAD.n6373 PAD.n5988 4.5005
R33258 PAD.n6163 PAD.n5979 4.5005
R33259 PAD.n6163 PAD.n5981 4.5005
R33260 PAD.n6373 PAD.n6163 4.5005
R33261 PAD.n5987 PAD.n5979 4.5005
R33262 PAD.n5987 PAD.n5981 4.5005
R33263 PAD.n6373 PAD.n5987 4.5005
R33264 PAD.n6166 PAD.n5979 4.5005
R33265 PAD.n6166 PAD.n5981 4.5005
R33266 PAD.n6373 PAD.n6166 4.5005
R33267 PAD.n5986 PAD.n5979 4.5005
R33268 PAD.n5986 PAD.n5981 4.5005
R33269 PAD.n6373 PAD.n5986 4.5005
R33270 PAD.n6169 PAD.n5979 4.5005
R33271 PAD.n6169 PAD.n5981 4.5005
R33272 PAD.n6373 PAD.n6169 4.5005
R33273 PAD.n5985 PAD.n5979 4.5005
R33274 PAD.n5985 PAD.n5981 4.5005
R33275 PAD.n6373 PAD.n5985 4.5005
R33276 PAD.n6172 PAD.n5979 4.5005
R33277 PAD.n6172 PAD.n5981 4.5005
R33278 PAD.n6373 PAD.n6172 4.5005
R33279 PAD.n5984 PAD.n5979 4.5005
R33280 PAD.n5984 PAD.n5981 4.5005
R33281 PAD.n6373 PAD.n5984 4.5005
R33282 PAD.n6175 PAD.n5979 4.5005
R33283 PAD.n6175 PAD.n5981 4.5005
R33284 PAD.n6373 PAD.n6175 4.5005
R33285 PAD.n5983 PAD.n5979 4.5005
R33286 PAD.n5983 PAD.n5981 4.5005
R33287 PAD.n6373 PAD.n5983 4.5005
R33288 PAD.n6372 PAD.n5979 4.5005
R33289 PAD.n6372 PAD.n5980 4.5005
R33290 PAD.n6372 PAD.n5981 4.5005
R33291 PAD.n6373 PAD.n6372 4.5005
R33292 PAD.n11508 PAD.n11105 4.5005
R33293 PAD.n11508 PAD.n11100 4.5005
R33294 PAD.n11509 PAD.n11508 4.5005
R33295 PAD.n11508 PAD.n11302 4.5005
R33296 PAD.n11508 PAD.n11507 4.5005
R33297 PAD.n6374 PAD.n5979 4.5005
R33298 PAD.n4 PAD 4.06833
R33299 PAD.n2 PAD.n1 3.98767
R33300 PAD.n8 PAD.n7 3.98767
R33301 PAD.n7808 PAD.n7807 2.65427
R33302 PAD.n3 PAD.n2 2.64417
R33303 PAD.n7 PAD.n6 2.64417
R33304 PAD.n5 PAD.n4 2.64417
R33305 PAD.n0 PAD.t4 2.55406
R33306 PAD.n11539 PAD.n11538 2.53369
R33307 PAD.n11104 PAD.n11103 2.25086
R33308 PAD.n7518 PAD.n7517 2.2505
R33309 PAD.n7209 PAD.n7201 2.2505
R33310 PAD.n7513 PAD.n7512 2.2505
R33311 PAD.n7510 PAD.n7509 2.2505
R33312 PAD.n7507 PAD.n7506 2.2505
R33313 PAD.n7499 PAD.n7229 2.2505
R33314 PAD.n7502 PAD.n7501 2.2505
R33315 PAD.n7498 PAD.n7497 2.2505
R33316 PAD.n7495 PAD.n7494 2.2505
R33317 PAD.n7487 PAD.n7231 2.2505
R33318 PAD.n7490 PAD.n7489 2.2505
R33319 PAD.n7486 PAD.n7485 2.2505
R33320 PAD.n7483 PAD.n7482 2.2505
R33321 PAD.n7475 PAD.n7233 2.2505
R33322 PAD.n7478 PAD.n7477 2.2505
R33323 PAD.n7474 PAD.n7473 2.2505
R33324 PAD.n7471 PAD.n7470 2.2505
R33325 PAD.n7463 PAD.n7235 2.2505
R33326 PAD.n7466 PAD.n7465 2.2505
R33327 PAD.n7462 PAD.n7461 2.2505
R33328 PAD.n7459 PAD.n7458 2.2505
R33329 PAD.n7451 PAD.n7237 2.2505
R33330 PAD.n7454 PAD.n7453 2.2505
R33331 PAD.n7450 PAD.n7449 2.2505
R33332 PAD.n7447 PAD.n7446 2.2505
R33333 PAD.n7439 PAD.n7239 2.2505
R33334 PAD.n7442 PAD.n7441 2.2505
R33335 PAD.n7438 PAD.n7437 2.2505
R33336 PAD.n7435 PAD.n7434 2.2505
R33337 PAD.n7427 PAD.n7241 2.2505
R33338 PAD.n7430 PAD.n7429 2.2505
R33339 PAD.n7426 PAD.n7425 2.2505
R33340 PAD.n7423 PAD.n7422 2.2505
R33341 PAD.n7415 PAD.n7243 2.2505
R33342 PAD.n7418 PAD.n7417 2.2505
R33343 PAD.n7414 PAD.n7413 2.2505
R33344 PAD.n7411 PAD.n7410 2.2505
R33345 PAD.n7403 PAD.n7245 2.2505
R33346 PAD.n7406 PAD.n7405 2.2505
R33347 PAD.n7402 PAD.n7401 2.2505
R33348 PAD.n7399 PAD.n7398 2.2505
R33349 PAD.n7391 PAD.n7247 2.2505
R33350 PAD.n7394 PAD.n7393 2.2505
R33351 PAD.n7390 PAD.n7389 2.2505
R33352 PAD.n7387 PAD.n7386 2.2505
R33353 PAD.n7379 PAD.n7249 2.2505
R33354 PAD.n7382 PAD.n7381 2.2505
R33355 PAD.n7378 PAD.n7377 2.2505
R33356 PAD.n7375 PAD.n7374 2.2505
R33357 PAD.n7367 PAD.n7251 2.2505
R33358 PAD.n7370 PAD.n7369 2.2505
R33359 PAD.n7366 PAD.n7365 2.2505
R33360 PAD.n7363 PAD.n7362 2.2505
R33361 PAD.n7355 PAD.n7253 2.2505
R33362 PAD.n7358 PAD.n7357 2.2505
R33363 PAD.n7354 PAD.n7353 2.2505
R33364 PAD.n7351 PAD.n7350 2.2505
R33365 PAD.n7343 PAD.n7255 2.2505
R33366 PAD.n7346 PAD.n7345 2.2505
R33367 PAD.n7342 PAD.n7341 2.2505
R33368 PAD.n7339 PAD.n7338 2.2505
R33369 PAD.n7331 PAD.n7257 2.2505
R33370 PAD.n7334 PAD.n7333 2.2505
R33371 PAD.n7330 PAD.n7329 2.2505
R33372 PAD.n7327 PAD.n7326 2.2505
R33373 PAD.n7319 PAD.n7259 2.2505
R33374 PAD.n7322 PAD.n7321 2.2505
R33375 PAD.n7318 PAD.n7317 2.2505
R33376 PAD.n7315 PAD.n7314 2.2505
R33377 PAD.n7307 PAD.n7261 2.2505
R33378 PAD.n7310 PAD.n7309 2.2505
R33379 PAD.n7306 PAD.n7305 2.2505
R33380 PAD.n7303 PAD.n7302 2.2505
R33381 PAD.n7295 PAD.n7263 2.2505
R33382 PAD.n7298 PAD.n7297 2.2505
R33383 PAD.n7294 PAD.n7293 2.2505
R33384 PAD.n7291 PAD.n7290 2.2505
R33385 PAD.n7283 PAD.n7265 2.2505
R33386 PAD.n7286 PAD.n7285 2.2505
R33387 PAD.n7282 PAD.n7281 2.2505
R33388 PAD.n7279 PAD.n7278 2.2505
R33389 PAD.n7271 PAD.n7267 2.2505
R33390 PAD.n7274 PAD.n7273 2.2505
R33391 PAD.n7270 PAD.n7269 2.2505
R33392 PAD.n7270 PAD.n7268 2.2505
R33393 PAD.n7275 PAD.n7274 2.2505
R33394 PAD.n7276 PAD.n7267 2.2505
R33395 PAD.n7278 PAD.n7277 2.2505
R33396 PAD.n7282 PAD.n7266 2.2505
R33397 PAD.n7287 PAD.n7286 2.2505
R33398 PAD.n7288 PAD.n7265 2.2505
R33399 PAD.n7290 PAD.n7289 2.2505
R33400 PAD.n7294 PAD.n7264 2.2505
R33401 PAD.n7299 PAD.n7298 2.2505
R33402 PAD.n7300 PAD.n7263 2.2505
R33403 PAD.n7302 PAD.n7301 2.2505
R33404 PAD.n7306 PAD.n7262 2.2505
R33405 PAD.n7311 PAD.n7310 2.2505
R33406 PAD.n7312 PAD.n7261 2.2505
R33407 PAD.n7314 PAD.n7313 2.2505
R33408 PAD.n7318 PAD.n7260 2.2505
R33409 PAD.n7323 PAD.n7322 2.2505
R33410 PAD.n7324 PAD.n7259 2.2505
R33411 PAD.n7326 PAD.n7325 2.2505
R33412 PAD.n7330 PAD.n7258 2.2505
R33413 PAD.n7335 PAD.n7334 2.2505
R33414 PAD.n7336 PAD.n7257 2.2505
R33415 PAD.n7338 PAD.n7337 2.2505
R33416 PAD.n7342 PAD.n7256 2.2505
R33417 PAD.n7347 PAD.n7346 2.2505
R33418 PAD.n7348 PAD.n7255 2.2505
R33419 PAD.n7350 PAD.n7349 2.2505
R33420 PAD.n7354 PAD.n7254 2.2505
R33421 PAD.n7359 PAD.n7358 2.2505
R33422 PAD.n7360 PAD.n7253 2.2505
R33423 PAD.n7362 PAD.n7361 2.2505
R33424 PAD.n7366 PAD.n7252 2.2505
R33425 PAD.n7371 PAD.n7370 2.2505
R33426 PAD.n7372 PAD.n7251 2.2505
R33427 PAD.n7374 PAD.n7373 2.2505
R33428 PAD.n7378 PAD.n7250 2.2505
R33429 PAD.n7383 PAD.n7382 2.2505
R33430 PAD.n7384 PAD.n7249 2.2505
R33431 PAD.n7386 PAD.n7385 2.2505
R33432 PAD.n7390 PAD.n7248 2.2505
R33433 PAD.n7395 PAD.n7394 2.2505
R33434 PAD.n7396 PAD.n7247 2.2505
R33435 PAD.n7398 PAD.n7397 2.2505
R33436 PAD.n7402 PAD.n7246 2.2505
R33437 PAD.n7407 PAD.n7406 2.2505
R33438 PAD.n7408 PAD.n7245 2.2505
R33439 PAD.n7410 PAD.n7409 2.2505
R33440 PAD.n7414 PAD.n7244 2.2505
R33441 PAD.n7419 PAD.n7418 2.2505
R33442 PAD.n7420 PAD.n7243 2.2505
R33443 PAD.n7422 PAD.n7421 2.2505
R33444 PAD.n7426 PAD.n7242 2.2505
R33445 PAD.n7431 PAD.n7430 2.2505
R33446 PAD.n7432 PAD.n7241 2.2505
R33447 PAD.n7434 PAD.n7433 2.2505
R33448 PAD.n7438 PAD.n7240 2.2505
R33449 PAD.n7443 PAD.n7442 2.2505
R33450 PAD.n7444 PAD.n7239 2.2505
R33451 PAD.n7446 PAD.n7445 2.2505
R33452 PAD.n7450 PAD.n7238 2.2505
R33453 PAD.n7455 PAD.n7454 2.2505
R33454 PAD.n7456 PAD.n7237 2.2505
R33455 PAD.n7458 PAD.n7457 2.2505
R33456 PAD.n7462 PAD.n7236 2.2505
R33457 PAD.n7467 PAD.n7466 2.2505
R33458 PAD.n7468 PAD.n7235 2.2505
R33459 PAD.n7470 PAD.n7469 2.2505
R33460 PAD.n7474 PAD.n7234 2.2505
R33461 PAD.n7479 PAD.n7478 2.2505
R33462 PAD.n7480 PAD.n7233 2.2505
R33463 PAD.n7482 PAD.n7481 2.2505
R33464 PAD.n7486 PAD.n7232 2.2505
R33465 PAD.n7491 PAD.n7490 2.2505
R33466 PAD.n7492 PAD.n7231 2.2505
R33467 PAD.n7494 PAD.n7493 2.2505
R33468 PAD.n7498 PAD.n7230 2.2505
R33469 PAD.n7503 PAD.n7502 2.2505
R33470 PAD.n7504 PAD.n7229 2.2505
R33471 PAD.n7506 PAD.n7505 2.2505
R33472 PAD.n7510 PAD.n7228 2.2505
R33473 PAD.n7514 PAD.n7513 2.2505
R33474 PAD.n7515 PAD.n7209 2.2505
R33475 PAD.n7517 PAD.n7516 2.2505
R33476 PAD.n10695 PAD.n415 2.2505
R33477 PAD.n10694 PAD.n10693 2.2505
R33478 PAD.n10691 PAD.n10417 2.2505
R33479 PAD.n10415 PAD.n10414 2.2505
R33480 PAD.n10687 PAD.n10686 2.2505
R33481 PAD.n10684 PAD.n10683 2.2505
R33482 PAD.n10682 PAD.n10422 2.2505
R33483 PAD.n10420 PAD.n10419 2.2505
R33484 PAD.n10678 PAD.n10677 2.2505
R33485 PAD.n10675 PAD.n10674 2.2505
R33486 PAD.n10673 PAD.n10427 2.2505
R33487 PAD.n10425 PAD.n10424 2.2505
R33488 PAD.n10669 PAD.n10668 2.2505
R33489 PAD.n10666 PAD.n10665 2.2505
R33490 PAD.n10664 PAD.n10432 2.2505
R33491 PAD.n10430 PAD.n10429 2.2505
R33492 PAD.n10660 PAD.n10659 2.2505
R33493 PAD.n10657 PAD.n10656 2.2505
R33494 PAD.n10655 PAD.n10437 2.2505
R33495 PAD.n10435 PAD.n10434 2.2505
R33496 PAD.n10651 PAD.n10650 2.2505
R33497 PAD.n10648 PAD.n10647 2.2505
R33498 PAD.n10646 PAD.n10442 2.2505
R33499 PAD.n10440 PAD.n10439 2.2505
R33500 PAD.n10642 PAD.n10641 2.2505
R33501 PAD.n10639 PAD.n10638 2.2505
R33502 PAD.n10637 PAD.n10447 2.2505
R33503 PAD.n10445 PAD.n10444 2.2505
R33504 PAD.n10633 PAD.n10632 2.2505
R33505 PAD.n10630 PAD.n10629 2.2505
R33506 PAD.n10628 PAD.n10452 2.2505
R33507 PAD.n10450 PAD.n10449 2.2505
R33508 PAD.n10624 PAD.n10623 2.2505
R33509 PAD.n10621 PAD.n10620 2.2505
R33510 PAD.n10619 PAD.n10457 2.2505
R33511 PAD.n10455 PAD.n10454 2.2505
R33512 PAD.n10615 PAD.n10614 2.2505
R33513 PAD.n10612 PAD.n10611 2.2505
R33514 PAD.n10610 PAD.n10462 2.2505
R33515 PAD.n10460 PAD.n10459 2.2505
R33516 PAD.n10606 PAD.n10605 2.2505
R33517 PAD.n10603 PAD.n10602 2.2505
R33518 PAD.n10601 PAD.n10467 2.2505
R33519 PAD.n10465 PAD.n10464 2.2505
R33520 PAD.n10597 PAD.n10596 2.2505
R33521 PAD.n10594 PAD.n10593 2.2505
R33522 PAD.n10592 PAD.n10472 2.2505
R33523 PAD.n10470 PAD.n10469 2.2505
R33524 PAD.n10588 PAD.n10587 2.2505
R33525 PAD.n10585 PAD.n10584 2.2505
R33526 PAD.n10583 PAD.n10477 2.2505
R33527 PAD.n10475 PAD.n10474 2.2505
R33528 PAD.n10579 PAD.n10578 2.2505
R33529 PAD.n10576 PAD.n10575 2.2505
R33530 PAD.n10574 PAD.n10482 2.2505
R33531 PAD.n10480 PAD.n10479 2.2505
R33532 PAD.n10570 PAD.n10569 2.2505
R33533 PAD.n10567 PAD.n10566 2.2505
R33534 PAD.n10565 PAD.n10487 2.2505
R33535 PAD.n10485 PAD.n10484 2.2505
R33536 PAD.n10561 PAD.n10560 2.2505
R33537 PAD.n10558 PAD.n10557 2.2505
R33538 PAD.n10556 PAD.n10492 2.2505
R33539 PAD.n10490 PAD.n10489 2.2505
R33540 PAD.n10552 PAD.n10551 2.2505
R33541 PAD.n10549 PAD.n10548 2.2505
R33542 PAD.n10547 PAD.n10497 2.2505
R33543 PAD.n10495 PAD.n10494 2.2505
R33544 PAD.n10543 PAD.n10542 2.2505
R33545 PAD.n10540 PAD.n10539 2.2505
R33546 PAD.n10538 PAD.n10502 2.2505
R33547 PAD.n10500 PAD.n10499 2.2505
R33548 PAD.n10534 PAD.n10533 2.2505
R33549 PAD.n10531 PAD.n10530 2.2505
R33550 PAD.n10529 PAD.n10507 2.2505
R33551 PAD.n10505 PAD.n10504 2.2505
R33552 PAD.n10525 PAD.n10524 2.2505
R33553 PAD.n10522 PAD.n10521 2.2505
R33554 PAD.n10520 PAD.n10512 2.2505
R33555 PAD.n10510 PAD.n10509 2.2505
R33556 PAD.n10516 PAD.n10515 2.2505
R33557 PAD.n10513 PAD.n420 2.2505
R33558 PAD.n10713 PAD.n10712 2.2505
R33559 PAD.n10715 PAD.n416 2.2505
R33560 PAD.n10710 PAD.n416 2.2505
R33561 PAD.n10712 PAD.n10711 2.2505
R33562 PAD.n421 PAD.n420 2.2505
R33563 PAD.n10517 PAD.n10516 2.2505
R33564 PAD.n10518 PAD.n10509 2.2505
R33565 PAD.n10520 PAD.n10519 2.2505
R33566 PAD.n10521 PAD.n10508 2.2505
R33567 PAD.n10526 PAD.n10525 2.2505
R33568 PAD.n10527 PAD.n10504 2.2505
R33569 PAD.n10529 PAD.n10528 2.2505
R33570 PAD.n10530 PAD.n10503 2.2505
R33571 PAD.n10535 PAD.n10534 2.2505
R33572 PAD.n10536 PAD.n10499 2.2505
R33573 PAD.n10538 PAD.n10537 2.2505
R33574 PAD.n10539 PAD.n10498 2.2505
R33575 PAD.n10544 PAD.n10543 2.2505
R33576 PAD.n10545 PAD.n10494 2.2505
R33577 PAD.n10547 PAD.n10546 2.2505
R33578 PAD.n10548 PAD.n10493 2.2505
R33579 PAD.n10553 PAD.n10552 2.2505
R33580 PAD.n10554 PAD.n10489 2.2505
R33581 PAD.n10556 PAD.n10555 2.2505
R33582 PAD.n10557 PAD.n10488 2.2505
R33583 PAD.n10562 PAD.n10561 2.2505
R33584 PAD.n10563 PAD.n10484 2.2505
R33585 PAD.n10565 PAD.n10564 2.2505
R33586 PAD.n10566 PAD.n10483 2.2505
R33587 PAD.n10571 PAD.n10570 2.2505
R33588 PAD.n10572 PAD.n10479 2.2505
R33589 PAD.n10574 PAD.n10573 2.2505
R33590 PAD.n10575 PAD.n10478 2.2505
R33591 PAD.n10580 PAD.n10579 2.2505
R33592 PAD.n10581 PAD.n10474 2.2505
R33593 PAD.n10583 PAD.n10582 2.2505
R33594 PAD.n10584 PAD.n10473 2.2505
R33595 PAD.n10589 PAD.n10588 2.2505
R33596 PAD.n10590 PAD.n10469 2.2505
R33597 PAD.n10592 PAD.n10591 2.2505
R33598 PAD.n10593 PAD.n10468 2.2505
R33599 PAD.n10598 PAD.n10597 2.2505
R33600 PAD.n10599 PAD.n10464 2.2505
R33601 PAD.n10601 PAD.n10600 2.2505
R33602 PAD.n10602 PAD.n10463 2.2505
R33603 PAD.n10607 PAD.n10606 2.2505
R33604 PAD.n10608 PAD.n10459 2.2505
R33605 PAD.n10610 PAD.n10609 2.2505
R33606 PAD.n10611 PAD.n10458 2.2505
R33607 PAD.n10616 PAD.n10615 2.2505
R33608 PAD.n10617 PAD.n10454 2.2505
R33609 PAD.n10619 PAD.n10618 2.2505
R33610 PAD.n10620 PAD.n10453 2.2505
R33611 PAD.n10625 PAD.n10624 2.2505
R33612 PAD.n10626 PAD.n10449 2.2505
R33613 PAD.n10628 PAD.n10627 2.2505
R33614 PAD.n10629 PAD.n10448 2.2505
R33615 PAD.n10634 PAD.n10633 2.2505
R33616 PAD.n10635 PAD.n10444 2.2505
R33617 PAD.n10637 PAD.n10636 2.2505
R33618 PAD.n10638 PAD.n10443 2.2505
R33619 PAD.n10643 PAD.n10642 2.2505
R33620 PAD.n10644 PAD.n10439 2.2505
R33621 PAD.n10646 PAD.n10645 2.2505
R33622 PAD.n10647 PAD.n10438 2.2505
R33623 PAD.n10652 PAD.n10651 2.2505
R33624 PAD.n10653 PAD.n10434 2.2505
R33625 PAD.n10655 PAD.n10654 2.2505
R33626 PAD.n10656 PAD.n10433 2.2505
R33627 PAD.n10661 PAD.n10660 2.2505
R33628 PAD.n10662 PAD.n10429 2.2505
R33629 PAD.n10664 PAD.n10663 2.2505
R33630 PAD.n10665 PAD.n10428 2.2505
R33631 PAD.n10670 PAD.n10669 2.2505
R33632 PAD.n10671 PAD.n10424 2.2505
R33633 PAD.n10673 PAD.n10672 2.2505
R33634 PAD.n10674 PAD.n10423 2.2505
R33635 PAD.n10679 PAD.n10678 2.2505
R33636 PAD.n10680 PAD.n10419 2.2505
R33637 PAD.n10682 PAD.n10681 2.2505
R33638 PAD.n10683 PAD.n10418 2.2505
R33639 PAD.n10688 PAD.n10687 2.2505
R33640 PAD.n10689 PAD.n10414 2.2505
R33641 PAD.n10691 PAD.n10690 2.2505
R33642 PAD.n10694 PAD.n10413 2.2505
R33643 PAD.n10696 PAD.n10695 2.2505
R33644 PAD.n523 PAD.n522 2.2505
R33645 PAD.n525 PAD.n520 2.2505
R33646 PAD.n530 PAD.n529 2.2505
R33647 PAD.n527 PAD.n518 2.2505
R33648 PAD.n535 PAD.n534 2.2505
R33649 PAD.n537 PAD.n516 2.2505
R33650 PAD.n542 PAD.n541 2.2505
R33651 PAD.n539 PAD.n514 2.2505
R33652 PAD.n547 PAD.n546 2.2505
R33653 PAD.n549 PAD.n512 2.2505
R33654 PAD.n554 PAD.n553 2.2505
R33655 PAD.n551 PAD.n510 2.2505
R33656 PAD.n559 PAD.n558 2.2505
R33657 PAD.n561 PAD.n508 2.2505
R33658 PAD.n566 PAD.n565 2.2505
R33659 PAD.n563 PAD.n506 2.2505
R33660 PAD.n571 PAD.n570 2.2505
R33661 PAD.n573 PAD.n504 2.2505
R33662 PAD.n578 PAD.n577 2.2505
R33663 PAD.n575 PAD.n502 2.2505
R33664 PAD.n583 PAD.n582 2.2505
R33665 PAD.n585 PAD.n500 2.2505
R33666 PAD.n590 PAD.n589 2.2505
R33667 PAD.n587 PAD.n498 2.2505
R33668 PAD.n595 PAD.n594 2.2505
R33669 PAD.n597 PAD.n496 2.2505
R33670 PAD.n602 PAD.n601 2.2505
R33671 PAD.n599 PAD.n494 2.2505
R33672 PAD.n607 PAD.n606 2.2505
R33673 PAD.n609 PAD.n492 2.2505
R33674 PAD.n614 PAD.n613 2.2505
R33675 PAD.n611 PAD.n490 2.2505
R33676 PAD.n619 PAD.n618 2.2505
R33677 PAD.n621 PAD.n488 2.2505
R33678 PAD.n626 PAD.n625 2.2505
R33679 PAD.n623 PAD.n486 2.2505
R33680 PAD.n631 PAD.n630 2.2505
R33681 PAD.n633 PAD.n484 2.2505
R33682 PAD.n638 PAD.n637 2.2505
R33683 PAD.n635 PAD.n482 2.2505
R33684 PAD.n643 PAD.n642 2.2505
R33685 PAD.n645 PAD.n480 2.2505
R33686 PAD.n650 PAD.n649 2.2505
R33687 PAD.n647 PAD.n478 2.2505
R33688 PAD.n655 PAD.n654 2.2505
R33689 PAD.n657 PAD.n476 2.2505
R33690 PAD.n662 PAD.n661 2.2505
R33691 PAD.n659 PAD.n474 2.2505
R33692 PAD.n667 PAD.n666 2.2505
R33693 PAD.n669 PAD.n472 2.2505
R33694 PAD.n674 PAD.n673 2.2505
R33695 PAD.n671 PAD.n470 2.2505
R33696 PAD.n679 PAD.n678 2.2505
R33697 PAD.n681 PAD.n468 2.2505
R33698 PAD.n686 PAD.n685 2.2505
R33699 PAD.n683 PAD.n466 2.2505
R33700 PAD.n691 PAD.n690 2.2505
R33701 PAD.n693 PAD.n464 2.2505
R33702 PAD.n698 PAD.n697 2.2505
R33703 PAD.n695 PAD.n462 2.2505
R33704 PAD.n703 PAD.n702 2.2505
R33705 PAD.n705 PAD.n460 2.2505
R33706 PAD.n710 PAD.n709 2.2505
R33707 PAD.n707 PAD.n458 2.2505
R33708 PAD.n715 PAD.n714 2.2505
R33709 PAD.n717 PAD.n456 2.2505
R33710 PAD.n722 PAD.n721 2.2505
R33711 PAD.n719 PAD.n454 2.2505
R33712 PAD.n727 PAD.n726 2.2505
R33713 PAD.n729 PAD.n452 2.2505
R33714 PAD.n734 PAD.n733 2.2505
R33715 PAD.n731 PAD.n450 2.2505
R33716 PAD.n739 PAD.n738 2.2505
R33717 PAD.n741 PAD.n448 2.2505
R33718 PAD.n746 PAD.n745 2.2505
R33719 PAD.n743 PAD.n446 2.2505
R33720 PAD.n751 PAD.n750 2.2505
R33721 PAD.n753 PAD.n444 2.2505
R33722 PAD.n758 PAD.n757 2.2505
R33723 PAD.n755 PAD.n442 2.2505
R33724 PAD.n764 PAD.n763 2.2505
R33725 PAD.n766 PAD.n440 2.2505
R33726 PAD.n768 PAD.n439 2.2505
R33727 PAD.n771 PAD.n770 2.2505
R33728 PAD.n772 PAD.n771 2.2505
R33729 PAD.n439 PAD.n438 2.2505
R33730 PAD.n761 PAD.n440 2.2505
R33731 PAD.n763 PAD.n762 2.2505
R33732 PAD.n760 PAD.n442 2.2505
R33733 PAD.n759 PAD.n758 2.2505
R33734 PAD.n444 PAD.n443 2.2505
R33735 PAD.n750 PAD.n749 2.2505
R33736 PAD.n748 PAD.n446 2.2505
R33737 PAD.n747 PAD.n746 2.2505
R33738 PAD.n448 PAD.n447 2.2505
R33739 PAD.n738 PAD.n737 2.2505
R33740 PAD.n736 PAD.n450 2.2505
R33741 PAD.n735 PAD.n734 2.2505
R33742 PAD.n452 PAD.n451 2.2505
R33743 PAD.n726 PAD.n725 2.2505
R33744 PAD.n724 PAD.n454 2.2505
R33745 PAD.n723 PAD.n722 2.2505
R33746 PAD.n456 PAD.n455 2.2505
R33747 PAD.n714 PAD.n713 2.2505
R33748 PAD.n712 PAD.n458 2.2505
R33749 PAD.n711 PAD.n710 2.2505
R33750 PAD.n460 PAD.n459 2.2505
R33751 PAD.n702 PAD.n701 2.2505
R33752 PAD.n700 PAD.n462 2.2505
R33753 PAD.n699 PAD.n698 2.2505
R33754 PAD.n464 PAD.n463 2.2505
R33755 PAD.n690 PAD.n689 2.2505
R33756 PAD.n688 PAD.n466 2.2505
R33757 PAD.n687 PAD.n686 2.2505
R33758 PAD.n468 PAD.n467 2.2505
R33759 PAD.n678 PAD.n677 2.2505
R33760 PAD.n676 PAD.n470 2.2505
R33761 PAD.n675 PAD.n674 2.2505
R33762 PAD.n472 PAD.n471 2.2505
R33763 PAD.n666 PAD.n665 2.2505
R33764 PAD.n664 PAD.n474 2.2505
R33765 PAD.n663 PAD.n662 2.2505
R33766 PAD.n476 PAD.n475 2.2505
R33767 PAD.n654 PAD.n653 2.2505
R33768 PAD.n652 PAD.n478 2.2505
R33769 PAD.n651 PAD.n650 2.2505
R33770 PAD.n480 PAD.n479 2.2505
R33771 PAD.n642 PAD.n641 2.2505
R33772 PAD.n640 PAD.n482 2.2505
R33773 PAD.n639 PAD.n638 2.2505
R33774 PAD.n484 PAD.n483 2.2505
R33775 PAD.n630 PAD.n629 2.2505
R33776 PAD.n628 PAD.n486 2.2505
R33777 PAD.n627 PAD.n626 2.2505
R33778 PAD.n488 PAD.n487 2.2505
R33779 PAD.n618 PAD.n617 2.2505
R33780 PAD.n616 PAD.n490 2.2505
R33781 PAD.n615 PAD.n614 2.2505
R33782 PAD.n492 PAD.n491 2.2505
R33783 PAD.n606 PAD.n605 2.2505
R33784 PAD.n604 PAD.n494 2.2505
R33785 PAD.n603 PAD.n602 2.2505
R33786 PAD.n496 PAD.n495 2.2505
R33787 PAD.n594 PAD.n593 2.2505
R33788 PAD.n592 PAD.n498 2.2505
R33789 PAD.n591 PAD.n590 2.2505
R33790 PAD.n500 PAD.n499 2.2505
R33791 PAD.n582 PAD.n581 2.2505
R33792 PAD.n580 PAD.n502 2.2505
R33793 PAD.n579 PAD.n578 2.2505
R33794 PAD.n504 PAD.n503 2.2505
R33795 PAD.n570 PAD.n569 2.2505
R33796 PAD.n568 PAD.n506 2.2505
R33797 PAD.n567 PAD.n566 2.2505
R33798 PAD.n508 PAD.n507 2.2505
R33799 PAD.n558 PAD.n557 2.2505
R33800 PAD.n556 PAD.n510 2.2505
R33801 PAD.n555 PAD.n554 2.2505
R33802 PAD.n512 PAD.n511 2.2505
R33803 PAD.n546 PAD.n545 2.2505
R33804 PAD.n544 PAD.n514 2.2505
R33805 PAD.n543 PAD.n542 2.2505
R33806 PAD.n516 PAD.n515 2.2505
R33807 PAD.n534 PAD.n533 2.2505
R33808 PAD.n532 PAD.n518 2.2505
R33809 PAD.n531 PAD.n530 2.2505
R33810 PAD.n520 PAD.n519 2.2505
R33811 PAD.n522 PAD.n521 2.2505
R33812 PAD.n872 PAD.n824 2.2505
R33813 PAD.n871 PAD.n870 2.2505
R33814 PAD.n877 PAD.n876 2.2505
R33815 PAD.n880 PAD.n879 2.2505
R33816 PAD.n884 PAD.n883 2.2505
R33817 PAD.n881 PAD.n867 2.2505
R33818 PAD.n889 PAD.n888 2.2505
R33819 PAD.n892 PAD.n891 2.2505
R33820 PAD.n896 PAD.n895 2.2505
R33821 PAD.n893 PAD.n865 2.2505
R33822 PAD.n901 PAD.n900 2.2505
R33823 PAD.n904 PAD.n903 2.2505
R33824 PAD.n908 PAD.n907 2.2505
R33825 PAD.n905 PAD.n863 2.2505
R33826 PAD.n913 PAD.n912 2.2505
R33827 PAD.n916 PAD.n915 2.2505
R33828 PAD.n920 PAD.n919 2.2505
R33829 PAD.n917 PAD.n861 2.2505
R33830 PAD.n925 PAD.n924 2.2505
R33831 PAD.n928 PAD.n927 2.2505
R33832 PAD.n932 PAD.n931 2.2505
R33833 PAD.n929 PAD.n859 2.2505
R33834 PAD.n937 PAD.n936 2.2505
R33835 PAD.n940 PAD.n939 2.2505
R33836 PAD.n944 PAD.n943 2.2505
R33837 PAD.n941 PAD.n857 2.2505
R33838 PAD.n949 PAD.n948 2.2505
R33839 PAD.n952 PAD.n951 2.2505
R33840 PAD.n956 PAD.n955 2.2505
R33841 PAD.n953 PAD.n855 2.2505
R33842 PAD.n961 PAD.n960 2.2505
R33843 PAD.n964 PAD.n963 2.2505
R33844 PAD.n968 PAD.n967 2.2505
R33845 PAD.n965 PAD.n853 2.2505
R33846 PAD.n973 PAD.n972 2.2505
R33847 PAD.n976 PAD.n975 2.2505
R33848 PAD.n980 PAD.n979 2.2505
R33849 PAD.n977 PAD.n851 2.2505
R33850 PAD.n985 PAD.n984 2.2505
R33851 PAD.n988 PAD.n987 2.2505
R33852 PAD.n992 PAD.n991 2.2505
R33853 PAD.n989 PAD.n849 2.2505
R33854 PAD.n997 PAD.n996 2.2505
R33855 PAD.n1000 PAD.n999 2.2505
R33856 PAD.n1004 PAD.n1003 2.2505
R33857 PAD.n1001 PAD.n847 2.2505
R33858 PAD.n1009 PAD.n1008 2.2505
R33859 PAD.n1012 PAD.n1011 2.2505
R33860 PAD.n1016 PAD.n1015 2.2505
R33861 PAD.n1013 PAD.n845 2.2505
R33862 PAD.n1021 PAD.n1020 2.2505
R33863 PAD.n1024 PAD.n1023 2.2505
R33864 PAD.n1028 PAD.n1027 2.2505
R33865 PAD.n1025 PAD.n843 2.2505
R33866 PAD.n1033 PAD.n1032 2.2505
R33867 PAD.n1036 PAD.n1035 2.2505
R33868 PAD.n1040 PAD.n1039 2.2505
R33869 PAD.n1037 PAD.n841 2.2505
R33870 PAD.n1045 PAD.n1044 2.2505
R33871 PAD.n1048 PAD.n1047 2.2505
R33872 PAD.n1052 PAD.n1051 2.2505
R33873 PAD.n1049 PAD.n839 2.2505
R33874 PAD.n1057 PAD.n1056 2.2505
R33875 PAD.n1060 PAD.n1059 2.2505
R33876 PAD.n1064 PAD.n1063 2.2505
R33877 PAD.n1061 PAD.n837 2.2505
R33878 PAD.n1069 PAD.n1068 2.2505
R33879 PAD.n1072 PAD.n1071 2.2505
R33880 PAD.n1076 PAD.n1075 2.2505
R33881 PAD.n1073 PAD.n835 2.2505
R33882 PAD.n1081 PAD.n1080 2.2505
R33883 PAD.n1084 PAD.n1083 2.2505
R33884 PAD.n1088 PAD.n1087 2.2505
R33885 PAD.n1085 PAD.n833 2.2505
R33886 PAD.n1093 PAD.n1092 2.2505
R33887 PAD.n1096 PAD.n1095 2.2505
R33888 PAD.n1100 PAD.n1099 2.2505
R33889 PAD.n1097 PAD.n831 2.2505
R33890 PAD.n1105 PAD.n1104 2.2505
R33891 PAD.n1108 PAD.n1107 2.2505
R33892 PAD.n1112 PAD.n1111 2.2505
R33893 PAD.n1109 PAD.n829 2.2505
R33894 PAD.n10385 PAD.n10384 2.2505
R33895 PAD.n10387 PAD.n826 2.2505
R33896 PAD.n10382 PAD.n826 2.2505
R33897 PAD.n10384 PAD.n10383 2.2505
R33898 PAD.n1114 PAD.n829 2.2505
R33899 PAD.n1113 PAD.n1112 2.2505
R33900 PAD.n1108 PAD.n830 2.2505
R33901 PAD.n1104 PAD.n1103 2.2505
R33902 PAD.n1102 PAD.n831 2.2505
R33903 PAD.n1101 PAD.n1100 2.2505
R33904 PAD.n1096 PAD.n832 2.2505
R33905 PAD.n1092 PAD.n1091 2.2505
R33906 PAD.n1090 PAD.n833 2.2505
R33907 PAD.n1089 PAD.n1088 2.2505
R33908 PAD.n1084 PAD.n834 2.2505
R33909 PAD.n1080 PAD.n1079 2.2505
R33910 PAD.n1078 PAD.n835 2.2505
R33911 PAD.n1077 PAD.n1076 2.2505
R33912 PAD.n1072 PAD.n836 2.2505
R33913 PAD.n1068 PAD.n1067 2.2505
R33914 PAD.n1066 PAD.n837 2.2505
R33915 PAD.n1065 PAD.n1064 2.2505
R33916 PAD.n1060 PAD.n838 2.2505
R33917 PAD.n1056 PAD.n1055 2.2505
R33918 PAD.n1054 PAD.n839 2.2505
R33919 PAD.n1053 PAD.n1052 2.2505
R33920 PAD.n1048 PAD.n840 2.2505
R33921 PAD.n1044 PAD.n1043 2.2505
R33922 PAD.n1042 PAD.n841 2.2505
R33923 PAD.n1041 PAD.n1040 2.2505
R33924 PAD.n1036 PAD.n842 2.2505
R33925 PAD.n1032 PAD.n1031 2.2505
R33926 PAD.n1030 PAD.n843 2.2505
R33927 PAD.n1029 PAD.n1028 2.2505
R33928 PAD.n1024 PAD.n844 2.2505
R33929 PAD.n1020 PAD.n1019 2.2505
R33930 PAD.n1018 PAD.n845 2.2505
R33931 PAD.n1017 PAD.n1016 2.2505
R33932 PAD.n1012 PAD.n846 2.2505
R33933 PAD.n1008 PAD.n1007 2.2505
R33934 PAD.n1006 PAD.n847 2.2505
R33935 PAD.n1005 PAD.n1004 2.2505
R33936 PAD.n1000 PAD.n848 2.2505
R33937 PAD.n996 PAD.n995 2.2505
R33938 PAD.n994 PAD.n849 2.2505
R33939 PAD.n993 PAD.n992 2.2505
R33940 PAD.n988 PAD.n850 2.2505
R33941 PAD.n984 PAD.n983 2.2505
R33942 PAD.n982 PAD.n851 2.2505
R33943 PAD.n981 PAD.n980 2.2505
R33944 PAD.n976 PAD.n852 2.2505
R33945 PAD.n972 PAD.n971 2.2505
R33946 PAD.n970 PAD.n853 2.2505
R33947 PAD.n969 PAD.n968 2.2505
R33948 PAD.n964 PAD.n854 2.2505
R33949 PAD.n960 PAD.n959 2.2505
R33950 PAD.n958 PAD.n855 2.2505
R33951 PAD.n957 PAD.n956 2.2505
R33952 PAD.n952 PAD.n856 2.2505
R33953 PAD.n948 PAD.n947 2.2505
R33954 PAD.n946 PAD.n857 2.2505
R33955 PAD.n945 PAD.n944 2.2505
R33956 PAD.n940 PAD.n858 2.2505
R33957 PAD.n936 PAD.n935 2.2505
R33958 PAD.n934 PAD.n859 2.2505
R33959 PAD.n933 PAD.n932 2.2505
R33960 PAD.n928 PAD.n860 2.2505
R33961 PAD.n924 PAD.n923 2.2505
R33962 PAD.n922 PAD.n861 2.2505
R33963 PAD.n921 PAD.n920 2.2505
R33964 PAD.n916 PAD.n862 2.2505
R33965 PAD.n912 PAD.n911 2.2505
R33966 PAD.n910 PAD.n863 2.2505
R33967 PAD.n909 PAD.n908 2.2505
R33968 PAD.n904 PAD.n864 2.2505
R33969 PAD.n900 PAD.n899 2.2505
R33970 PAD.n898 PAD.n865 2.2505
R33971 PAD.n897 PAD.n896 2.2505
R33972 PAD.n892 PAD.n866 2.2505
R33973 PAD.n888 PAD.n887 2.2505
R33974 PAD.n886 PAD.n867 2.2505
R33975 PAD.n885 PAD.n884 2.2505
R33976 PAD.n880 PAD.n868 2.2505
R33977 PAD.n876 PAD.n875 2.2505
R33978 PAD.n874 PAD.n871 2.2505
R33979 PAD.n873 PAD.n872 2.2505
R33980 PAD.n10106 PAD.n10105 2.2505
R33981 PAD.n10108 PAD.n10104 2.2505
R33982 PAD.n10113 PAD.n10112 2.2505
R33983 PAD.n10110 PAD.n10102 2.2505
R33984 PAD.n10118 PAD.n10117 2.2505
R33985 PAD.n10120 PAD.n10100 2.2505
R33986 PAD.n10125 PAD.n10124 2.2505
R33987 PAD.n10122 PAD.n10098 2.2505
R33988 PAD.n10130 PAD.n10129 2.2505
R33989 PAD.n10132 PAD.n10096 2.2505
R33990 PAD.n10137 PAD.n10136 2.2505
R33991 PAD.n10134 PAD.n10094 2.2505
R33992 PAD.n10142 PAD.n10141 2.2505
R33993 PAD.n10144 PAD.n10092 2.2505
R33994 PAD.n10149 PAD.n10148 2.2505
R33995 PAD.n10146 PAD.n10090 2.2505
R33996 PAD.n10154 PAD.n10153 2.2505
R33997 PAD.n10156 PAD.n10088 2.2505
R33998 PAD.n10161 PAD.n10160 2.2505
R33999 PAD.n10158 PAD.n10086 2.2505
R34000 PAD.n10166 PAD.n10165 2.2505
R34001 PAD.n10168 PAD.n10084 2.2505
R34002 PAD.n10173 PAD.n10172 2.2505
R34003 PAD.n10170 PAD.n10082 2.2505
R34004 PAD.n10178 PAD.n10177 2.2505
R34005 PAD.n10180 PAD.n10080 2.2505
R34006 PAD.n10185 PAD.n10184 2.2505
R34007 PAD.n10182 PAD.n10078 2.2505
R34008 PAD.n10190 PAD.n10189 2.2505
R34009 PAD.n10192 PAD.n10076 2.2505
R34010 PAD.n10197 PAD.n10196 2.2505
R34011 PAD.n10194 PAD.n10074 2.2505
R34012 PAD.n10202 PAD.n10201 2.2505
R34013 PAD.n10204 PAD.n10072 2.2505
R34014 PAD.n10209 PAD.n10208 2.2505
R34015 PAD.n10206 PAD.n10070 2.2505
R34016 PAD.n10214 PAD.n10213 2.2505
R34017 PAD.n10216 PAD.n10068 2.2505
R34018 PAD.n10221 PAD.n10220 2.2505
R34019 PAD.n10218 PAD.n10066 2.2505
R34020 PAD.n10226 PAD.n10225 2.2505
R34021 PAD.n10228 PAD.n10064 2.2505
R34022 PAD.n10233 PAD.n10232 2.2505
R34023 PAD.n10230 PAD.n10062 2.2505
R34024 PAD.n10238 PAD.n10237 2.2505
R34025 PAD.n10240 PAD.n10060 2.2505
R34026 PAD.n10245 PAD.n10244 2.2505
R34027 PAD.n10242 PAD.n10058 2.2505
R34028 PAD.n10250 PAD.n10249 2.2505
R34029 PAD.n10252 PAD.n10056 2.2505
R34030 PAD.n10257 PAD.n10256 2.2505
R34031 PAD.n10254 PAD.n10054 2.2505
R34032 PAD.n10262 PAD.n10261 2.2505
R34033 PAD.n10264 PAD.n10052 2.2505
R34034 PAD.n10269 PAD.n10268 2.2505
R34035 PAD.n10266 PAD.n10050 2.2505
R34036 PAD.n10274 PAD.n10273 2.2505
R34037 PAD.n10276 PAD.n10048 2.2505
R34038 PAD.n10281 PAD.n10280 2.2505
R34039 PAD.n10278 PAD.n10046 2.2505
R34040 PAD.n10286 PAD.n10285 2.2505
R34041 PAD.n10288 PAD.n10044 2.2505
R34042 PAD.n10293 PAD.n10292 2.2505
R34043 PAD.n10290 PAD.n10042 2.2505
R34044 PAD.n10298 PAD.n10297 2.2505
R34045 PAD.n10300 PAD.n10040 2.2505
R34046 PAD.n10305 PAD.n10304 2.2505
R34047 PAD.n10302 PAD.n10038 2.2505
R34048 PAD.n10310 PAD.n10309 2.2505
R34049 PAD.n10312 PAD.n10036 2.2505
R34050 PAD.n10317 PAD.n10316 2.2505
R34051 PAD.n10314 PAD.n10034 2.2505
R34052 PAD.n10322 PAD.n10321 2.2505
R34053 PAD.n10324 PAD.n10032 2.2505
R34054 PAD.n10329 PAD.n10328 2.2505
R34055 PAD.n10326 PAD.n10030 2.2505
R34056 PAD.n10334 PAD.n10333 2.2505
R34057 PAD.n10336 PAD.n10028 2.2505
R34058 PAD.n10341 PAD.n10340 2.2505
R34059 PAD.n10338 PAD.n10026 2.2505
R34060 PAD.n10347 PAD.n10346 2.2505
R34061 PAD.n10349 PAD.n10024 2.2505
R34062 PAD.n10351 PAD.n10023 2.2505
R34063 PAD.n10354 PAD.n10353 2.2505
R34064 PAD.n10355 PAD.n10354 2.2505
R34065 PAD.n10023 PAD.n10022 2.2505
R34066 PAD.n10344 PAD.n10024 2.2505
R34067 PAD.n10346 PAD.n10345 2.2505
R34068 PAD.n10343 PAD.n10026 2.2505
R34069 PAD.n10342 PAD.n10341 2.2505
R34070 PAD.n10028 PAD.n10027 2.2505
R34071 PAD.n10333 PAD.n10332 2.2505
R34072 PAD.n10331 PAD.n10030 2.2505
R34073 PAD.n10330 PAD.n10329 2.2505
R34074 PAD.n10032 PAD.n10031 2.2505
R34075 PAD.n10321 PAD.n10320 2.2505
R34076 PAD.n10319 PAD.n10034 2.2505
R34077 PAD.n10318 PAD.n10317 2.2505
R34078 PAD.n10036 PAD.n10035 2.2505
R34079 PAD.n10309 PAD.n10308 2.2505
R34080 PAD.n10307 PAD.n10038 2.2505
R34081 PAD.n10306 PAD.n10305 2.2505
R34082 PAD.n10040 PAD.n10039 2.2505
R34083 PAD.n10297 PAD.n10296 2.2505
R34084 PAD.n10295 PAD.n10042 2.2505
R34085 PAD.n10294 PAD.n10293 2.2505
R34086 PAD.n10044 PAD.n10043 2.2505
R34087 PAD.n10285 PAD.n10284 2.2505
R34088 PAD.n10283 PAD.n10046 2.2505
R34089 PAD.n10282 PAD.n10281 2.2505
R34090 PAD.n10048 PAD.n10047 2.2505
R34091 PAD.n10273 PAD.n10272 2.2505
R34092 PAD.n10271 PAD.n10050 2.2505
R34093 PAD.n10270 PAD.n10269 2.2505
R34094 PAD.n10052 PAD.n10051 2.2505
R34095 PAD.n10261 PAD.n10260 2.2505
R34096 PAD.n10259 PAD.n10054 2.2505
R34097 PAD.n10258 PAD.n10257 2.2505
R34098 PAD.n10056 PAD.n10055 2.2505
R34099 PAD.n10249 PAD.n10248 2.2505
R34100 PAD.n10247 PAD.n10058 2.2505
R34101 PAD.n10246 PAD.n10245 2.2505
R34102 PAD.n10060 PAD.n10059 2.2505
R34103 PAD.n10237 PAD.n10236 2.2505
R34104 PAD.n10235 PAD.n10062 2.2505
R34105 PAD.n10234 PAD.n10233 2.2505
R34106 PAD.n10064 PAD.n10063 2.2505
R34107 PAD.n10225 PAD.n10224 2.2505
R34108 PAD.n10223 PAD.n10066 2.2505
R34109 PAD.n10222 PAD.n10221 2.2505
R34110 PAD.n10068 PAD.n10067 2.2505
R34111 PAD.n10213 PAD.n10212 2.2505
R34112 PAD.n10211 PAD.n10070 2.2505
R34113 PAD.n10210 PAD.n10209 2.2505
R34114 PAD.n10072 PAD.n10071 2.2505
R34115 PAD.n10201 PAD.n10200 2.2505
R34116 PAD.n10199 PAD.n10074 2.2505
R34117 PAD.n10198 PAD.n10197 2.2505
R34118 PAD.n10076 PAD.n10075 2.2505
R34119 PAD.n10189 PAD.n10188 2.2505
R34120 PAD.n10187 PAD.n10078 2.2505
R34121 PAD.n10186 PAD.n10185 2.2505
R34122 PAD.n10080 PAD.n10079 2.2505
R34123 PAD.n10177 PAD.n10176 2.2505
R34124 PAD.n10175 PAD.n10082 2.2505
R34125 PAD.n10174 PAD.n10173 2.2505
R34126 PAD.n10084 PAD.n10083 2.2505
R34127 PAD.n10165 PAD.n10164 2.2505
R34128 PAD.n10163 PAD.n10086 2.2505
R34129 PAD.n10162 PAD.n10161 2.2505
R34130 PAD.n10088 PAD.n10087 2.2505
R34131 PAD.n10153 PAD.n10152 2.2505
R34132 PAD.n10151 PAD.n10090 2.2505
R34133 PAD.n10150 PAD.n10149 2.2505
R34134 PAD.n10092 PAD.n10091 2.2505
R34135 PAD.n10141 PAD.n10140 2.2505
R34136 PAD.n10139 PAD.n10094 2.2505
R34137 PAD.n10138 PAD.n10137 2.2505
R34138 PAD.n10096 PAD.n10095 2.2505
R34139 PAD.n10129 PAD.n10128 2.2505
R34140 PAD.n10127 PAD.n10098 2.2505
R34141 PAD.n10126 PAD.n10125 2.2505
R34142 PAD.n10100 PAD.n10099 2.2505
R34143 PAD.n10117 PAD.n10116 2.2505
R34144 PAD.n10115 PAD.n10102 2.2505
R34145 PAD.n10114 PAD.n10113 2.2505
R34146 PAD.n10104 PAD.n10103 2.2505
R34147 PAD.n10105 PAD.n1124 2.2505
R34148 PAD.n1481 PAD.n1480 2.2505
R34149 PAD.n1479 PAD.n1190 2.2505
R34150 PAD.n1193 PAD.n1192 2.2505
R34151 PAD.n1475 PAD.n1474 2.2505
R34152 PAD.n1472 PAD.n1471 2.2505
R34153 PAD.n1470 PAD.n1198 2.2505
R34154 PAD.n1196 PAD.n1195 2.2505
R34155 PAD.n1466 PAD.n1465 2.2505
R34156 PAD.n1463 PAD.n1462 2.2505
R34157 PAD.n1461 PAD.n1203 2.2505
R34158 PAD.n1201 PAD.n1200 2.2505
R34159 PAD.n1457 PAD.n1456 2.2505
R34160 PAD.n1454 PAD.n1453 2.2505
R34161 PAD.n1452 PAD.n1208 2.2505
R34162 PAD.n1206 PAD.n1205 2.2505
R34163 PAD.n1448 PAD.n1447 2.2505
R34164 PAD.n1445 PAD.n1444 2.2505
R34165 PAD.n1443 PAD.n1213 2.2505
R34166 PAD.n1211 PAD.n1210 2.2505
R34167 PAD.n1439 PAD.n1438 2.2505
R34168 PAD.n1436 PAD.n1435 2.2505
R34169 PAD.n1434 PAD.n1218 2.2505
R34170 PAD.n1216 PAD.n1215 2.2505
R34171 PAD.n1430 PAD.n1429 2.2505
R34172 PAD.n1427 PAD.n1426 2.2505
R34173 PAD.n1425 PAD.n1223 2.2505
R34174 PAD.n1221 PAD.n1220 2.2505
R34175 PAD.n1421 PAD.n1420 2.2505
R34176 PAD.n1418 PAD.n1417 2.2505
R34177 PAD.n1416 PAD.n1228 2.2505
R34178 PAD.n1226 PAD.n1225 2.2505
R34179 PAD.n1412 PAD.n1411 2.2505
R34180 PAD.n1409 PAD.n1408 2.2505
R34181 PAD.n1407 PAD.n1233 2.2505
R34182 PAD.n1231 PAD.n1230 2.2505
R34183 PAD.n1403 PAD.n1402 2.2505
R34184 PAD.n1400 PAD.n1399 2.2505
R34185 PAD.n1398 PAD.n1238 2.2505
R34186 PAD.n1236 PAD.n1235 2.2505
R34187 PAD.n1394 PAD.n1393 2.2505
R34188 PAD.n1391 PAD.n1390 2.2505
R34189 PAD.n1389 PAD.n1243 2.2505
R34190 PAD.n1241 PAD.n1240 2.2505
R34191 PAD.n1385 PAD.n1384 2.2505
R34192 PAD.n1382 PAD.n1381 2.2505
R34193 PAD.n1380 PAD.n1248 2.2505
R34194 PAD.n1246 PAD.n1245 2.2505
R34195 PAD.n1376 PAD.n1375 2.2505
R34196 PAD.n1373 PAD.n1372 2.2505
R34197 PAD.n1371 PAD.n1253 2.2505
R34198 PAD.n1251 PAD.n1250 2.2505
R34199 PAD.n1367 PAD.n1366 2.2505
R34200 PAD.n1364 PAD.n1363 2.2505
R34201 PAD.n1362 PAD.n1258 2.2505
R34202 PAD.n1256 PAD.n1255 2.2505
R34203 PAD.n1358 PAD.n1357 2.2505
R34204 PAD.n1355 PAD.n1354 2.2505
R34205 PAD.n1353 PAD.n1263 2.2505
R34206 PAD.n1261 PAD.n1260 2.2505
R34207 PAD.n1349 PAD.n1348 2.2505
R34208 PAD.n1346 PAD.n1345 2.2505
R34209 PAD.n1344 PAD.n1268 2.2505
R34210 PAD.n1266 PAD.n1265 2.2505
R34211 PAD.n1340 PAD.n1339 2.2505
R34212 PAD.n1337 PAD.n1336 2.2505
R34213 PAD.n1335 PAD.n1273 2.2505
R34214 PAD.n1271 PAD.n1270 2.2505
R34215 PAD.n1331 PAD.n1330 2.2505
R34216 PAD.n1328 PAD.n1327 2.2505
R34217 PAD.n1326 PAD.n1278 2.2505
R34218 PAD.n1276 PAD.n1275 2.2505
R34219 PAD.n1322 PAD.n1321 2.2505
R34220 PAD.n1319 PAD.n1318 2.2505
R34221 PAD.n1317 PAD.n1283 2.2505
R34222 PAD.n1281 PAD.n1280 2.2505
R34223 PAD.n1313 PAD.n1312 2.2505
R34224 PAD.n1310 PAD.n1309 2.2505
R34225 PAD.n1308 PAD.n1288 2.2505
R34226 PAD.n1286 PAD.n1285 2.2505
R34227 PAD.n1304 PAD.n1303 2.2505
R34228 PAD.n1301 PAD.n1300 2.2505
R34229 PAD.n1299 PAD.n1293 2.2505
R34230 PAD.n1291 PAD.n1290 2.2505
R34231 PAD.n1295 PAD.n1294 2.2505
R34232 PAD.n1296 PAD.n1295 2.2505
R34233 PAD.n1297 PAD.n1290 2.2505
R34234 PAD.n1299 PAD.n1298 2.2505
R34235 PAD.n1300 PAD.n1289 2.2505
R34236 PAD.n1305 PAD.n1304 2.2505
R34237 PAD.n1306 PAD.n1285 2.2505
R34238 PAD.n1308 PAD.n1307 2.2505
R34239 PAD.n1309 PAD.n1284 2.2505
R34240 PAD.n1314 PAD.n1313 2.2505
R34241 PAD.n1315 PAD.n1280 2.2505
R34242 PAD.n1317 PAD.n1316 2.2505
R34243 PAD.n1318 PAD.n1279 2.2505
R34244 PAD.n1323 PAD.n1322 2.2505
R34245 PAD.n1324 PAD.n1275 2.2505
R34246 PAD.n1326 PAD.n1325 2.2505
R34247 PAD.n1327 PAD.n1274 2.2505
R34248 PAD.n1332 PAD.n1331 2.2505
R34249 PAD.n1333 PAD.n1270 2.2505
R34250 PAD.n1335 PAD.n1334 2.2505
R34251 PAD.n1336 PAD.n1269 2.2505
R34252 PAD.n1341 PAD.n1340 2.2505
R34253 PAD.n1342 PAD.n1265 2.2505
R34254 PAD.n1344 PAD.n1343 2.2505
R34255 PAD.n1345 PAD.n1264 2.2505
R34256 PAD.n1350 PAD.n1349 2.2505
R34257 PAD.n1351 PAD.n1260 2.2505
R34258 PAD.n1353 PAD.n1352 2.2505
R34259 PAD.n1354 PAD.n1259 2.2505
R34260 PAD.n1359 PAD.n1358 2.2505
R34261 PAD.n1360 PAD.n1255 2.2505
R34262 PAD.n1362 PAD.n1361 2.2505
R34263 PAD.n1363 PAD.n1254 2.2505
R34264 PAD.n1368 PAD.n1367 2.2505
R34265 PAD.n1369 PAD.n1250 2.2505
R34266 PAD.n1371 PAD.n1370 2.2505
R34267 PAD.n1372 PAD.n1249 2.2505
R34268 PAD.n1377 PAD.n1376 2.2505
R34269 PAD.n1378 PAD.n1245 2.2505
R34270 PAD.n1380 PAD.n1379 2.2505
R34271 PAD.n1381 PAD.n1244 2.2505
R34272 PAD.n1386 PAD.n1385 2.2505
R34273 PAD.n1387 PAD.n1240 2.2505
R34274 PAD.n1389 PAD.n1388 2.2505
R34275 PAD.n1390 PAD.n1239 2.2505
R34276 PAD.n1395 PAD.n1394 2.2505
R34277 PAD.n1396 PAD.n1235 2.2505
R34278 PAD.n1398 PAD.n1397 2.2505
R34279 PAD.n1399 PAD.n1234 2.2505
R34280 PAD.n1404 PAD.n1403 2.2505
R34281 PAD.n1405 PAD.n1230 2.2505
R34282 PAD.n1407 PAD.n1406 2.2505
R34283 PAD.n1408 PAD.n1229 2.2505
R34284 PAD.n1413 PAD.n1412 2.2505
R34285 PAD.n1414 PAD.n1225 2.2505
R34286 PAD.n1416 PAD.n1415 2.2505
R34287 PAD.n1417 PAD.n1224 2.2505
R34288 PAD.n1422 PAD.n1421 2.2505
R34289 PAD.n1423 PAD.n1220 2.2505
R34290 PAD.n1425 PAD.n1424 2.2505
R34291 PAD.n1426 PAD.n1219 2.2505
R34292 PAD.n1431 PAD.n1430 2.2505
R34293 PAD.n1432 PAD.n1215 2.2505
R34294 PAD.n1434 PAD.n1433 2.2505
R34295 PAD.n1435 PAD.n1214 2.2505
R34296 PAD.n1440 PAD.n1439 2.2505
R34297 PAD.n1441 PAD.n1210 2.2505
R34298 PAD.n1443 PAD.n1442 2.2505
R34299 PAD.n1444 PAD.n1209 2.2505
R34300 PAD.n1449 PAD.n1448 2.2505
R34301 PAD.n1450 PAD.n1205 2.2505
R34302 PAD.n1452 PAD.n1451 2.2505
R34303 PAD.n1453 PAD.n1204 2.2505
R34304 PAD.n1458 PAD.n1457 2.2505
R34305 PAD.n1459 PAD.n1200 2.2505
R34306 PAD.n1461 PAD.n1460 2.2505
R34307 PAD.n1462 PAD.n1199 2.2505
R34308 PAD.n1467 PAD.n1466 2.2505
R34309 PAD.n1468 PAD.n1195 2.2505
R34310 PAD.n1470 PAD.n1469 2.2505
R34311 PAD.n1471 PAD.n1194 2.2505
R34312 PAD.n1476 PAD.n1475 2.2505
R34313 PAD.n1477 PAD.n1193 2.2505
R34314 PAD.n1479 PAD.n1478 2.2505
R34315 PAD.n1480 PAD.n1145 2.2505
R34316 PAD.n9749 PAD.n1531 2.2505
R34317 PAD.n1579 PAD.n1578 2.2505
R34318 PAD.n9754 PAD.n9753 2.2505
R34319 PAD.n9757 PAD.n9756 2.2505
R34320 PAD.n9761 PAD.n9760 2.2505
R34321 PAD.n9758 PAD.n1575 2.2505
R34322 PAD.n9766 PAD.n9765 2.2505
R34323 PAD.n9769 PAD.n9768 2.2505
R34324 PAD.n9773 PAD.n9772 2.2505
R34325 PAD.n9770 PAD.n1573 2.2505
R34326 PAD.n9778 PAD.n9777 2.2505
R34327 PAD.n9781 PAD.n9780 2.2505
R34328 PAD.n9785 PAD.n9784 2.2505
R34329 PAD.n9782 PAD.n1571 2.2505
R34330 PAD.n9790 PAD.n9789 2.2505
R34331 PAD.n9793 PAD.n9792 2.2505
R34332 PAD.n9797 PAD.n9796 2.2505
R34333 PAD.n9794 PAD.n1569 2.2505
R34334 PAD.n9802 PAD.n9801 2.2505
R34335 PAD.n9805 PAD.n9804 2.2505
R34336 PAD.n9809 PAD.n9808 2.2505
R34337 PAD.n9806 PAD.n1567 2.2505
R34338 PAD.n9814 PAD.n9813 2.2505
R34339 PAD.n9817 PAD.n9816 2.2505
R34340 PAD.n9821 PAD.n9820 2.2505
R34341 PAD.n9818 PAD.n1565 2.2505
R34342 PAD.n9826 PAD.n9825 2.2505
R34343 PAD.n9829 PAD.n9828 2.2505
R34344 PAD.n9833 PAD.n9832 2.2505
R34345 PAD.n9830 PAD.n1563 2.2505
R34346 PAD.n9838 PAD.n9837 2.2505
R34347 PAD.n9841 PAD.n9840 2.2505
R34348 PAD.n9845 PAD.n9844 2.2505
R34349 PAD.n9842 PAD.n1561 2.2505
R34350 PAD.n9850 PAD.n9849 2.2505
R34351 PAD.n9853 PAD.n9852 2.2505
R34352 PAD.n9857 PAD.n9856 2.2505
R34353 PAD.n9854 PAD.n1559 2.2505
R34354 PAD.n9862 PAD.n9861 2.2505
R34355 PAD.n9865 PAD.n9864 2.2505
R34356 PAD.n9869 PAD.n9868 2.2505
R34357 PAD.n9866 PAD.n1557 2.2505
R34358 PAD.n9874 PAD.n9873 2.2505
R34359 PAD.n9877 PAD.n9876 2.2505
R34360 PAD.n9881 PAD.n9880 2.2505
R34361 PAD.n9878 PAD.n1555 2.2505
R34362 PAD.n9886 PAD.n9885 2.2505
R34363 PAD.n9889 PAD.n9888 2.2505
R34364 PAD.n9893 PAD.n9892 2.2505
R34365 PAD.n9890 PAD.n1553 2.2505
R34366 PAD.n9898 PAD.n9897 2.2505
R34367 PAD.n9901 PAD.n9900 2.2505
R34368 PAD.n9905 PAD.n9904 2.2505
R34369 PAD.n9902 PAD.n1551 2.2505
R34370 PAD.n9910 PAD.n9909 2.2505
R34371 PAD.n9913 PAD.n9912 2.2505
R34372 PAD.n9917 PAD.n9916 2.2505
R34373 PAD.n9914 PAD.n1549 2.2505
R34374 PAD.n9922 PAD.n9921 2.2505
R34375 PAD.n9925 PAD.n9924 2.2505
R34376 PAD.n9929 PAD.n9928 2.2505
R34377 PAD.n9926 PAD.n1547 2.2505
R34378 PAD.n9934 PAD.n9933 2.2505
R34379 PAD.n9937 PAD.n9936 2.2505
R34380 PAD.n9941 PAD.n9940 2.2505
R34381 PAD.n9938 PAD.n1545 2.2505
R34382 PAD.n9946 PAD.n9945 2.2505
R34383 PAD.n9949 PAD.n9948 2.2505
R34384 PAD.n9953 PAD.n9952 2.2505
R34385 PAD.n9950 PAD.n1543 2.2505
R34386 PAD.n9958 PAD.n9957 2.2505
R34387 PAD.n9961 PAD.n9960 2.2505
R34388 PAD.n9965 PAD.n9964 2.2505
R34389 PAD.n9962 PAD.n1541 2.2505
R34390 PAD.n9970 PAD.n9969 2.2505
R34391 PAD.n9973 PAD.n9972 2.2505
R34392 PAD.n9977 PAD.n9976 2.2505
R34393 PAD.n9974 PAD.n1539 2.2505
R34394 PAD.n9982 PAD.n9981 2.2505
R34395 PAD.n9985 PAD.n9984 2.2505
R34396 PAD.n9989 PAD.n9988 2.2505
R34397 PAD.n9986 PAD.n1537 2.2505
R34398 PAD.n9995 PAD.n9994 2.2505
R34399 PAD.n9997 PAD.n1535 2.2505
R34400 PAD.n9992 PAD.n1535 2.2505
R34401 PAD.n9994 PAD.n9993 2.2505
R34402 PAD.n9991 PAD.n1537 2.2505
R34403 PAD.n9990 PAD.n9989 2.2505
R34404 PAD.n9985 PAD.n1538 2.2505
R34405 PAD.n9981 PAD.n9980 2.2505
R34406 PAD.n9979 PAD.n1539 2.2505
R34407 PAD.n9978 PAD.n9977 2.2505
R34408 PAD.n9973 PAD.n1540 2.2505
R34409 PAD.n9969 PAD.n9968 2.2505
R34410 PAD.n9967 PAD.n1541 2.2505
R34411 PAD.n9966 PAD.n9965 2.2505
R34412 PAD.n9961 PAD.n1542 2.2505
R34413 PAD.n9957 PAD.n9956 2.2505
R34414 PAD.n9955 PAD.n1543 2.2505
R34415 PAD.n9954 PAD.n9953 2.2505
R34416 PAD.n9949 PAD.n1544 2.2505
R34417 PAD.n9945 PAD.n9944 2.2505
R34418 PAD.n9943 PAD.n1545 2.2505
R34419 PAD.n9942 PAD.n9941 2.2505
R34420 PAD.n9937 PAD.n1546 2.2505
R34421 PAD.n9933 PAD.n9932 2.2505
R34422 PAD.n9931 PAD.n1547 2.2505
R34423 PAD.n9930 PAD.n9929 2.2505
R34424 PAD.n9925 PAD.n1548 2.2505
R34425 PAD.n9921 PAD.n9920 2.2505
R34426 PAD.n9919 PAD.n1549 2.2505
R34427 PAD.n9918 PAD.n9917 2.2505
R34428 PAD.n9913 PAD.n1550 2.2505
R34429 PAD.n9909 PAD.n9908 2.2505
R34430 PAD.n9907 PAD.n1551 2.2505
R34431 PAD.n9906 PAD.n9905 2.2505
R34432 PAD.n9901 PAD.n1552 2.2505
R34433 PAD.n9897 PAD.n9896 2.2505
R34434 PAD.n9895 PAD.n1553 2.2505
R34435 PAD.n9894 PAD.n9893 2.2505
R34436 PAD.n9889 PAD.n1554 2.2505
R34437 PAD.n9885 PAD.n9884 2.2505
R34438 PAD.n9883 PAD.n1555 2.2505
R34439 PAD.n9882 PAD.n9881 2.2505
R34440 PAD.n9877 PAD.n1556 2.2505
R34441 PAD.n9873 PAD.n9872 2.2505
R34442 PAD.n9871 PAD.n1557 2.2505
R34443 PAD.n9870 PAD.n9869 2.2505
R34444 PAD.n9865 PAD.n1558 2.2505
R34445 PAD.n9861 PAD.n9860 2.2505
R34446 PAD.n9859 PAD.n1559 2.2505
R34447 PAD.n9858 PAD.n9857 2.2505
R34448 PAD.n9853 PAD.n1560 2.2505
R34449 PAD.n9849 PAD.n9848 2.2505
R34450 PAD.n9847 PAD.n1561 2.2505
R34451 PAD.n9846 PAD.n9845 2.2505
R34452 PAD.n9841 PAD.n1562 2.2505
R34453 PAD.n9837 PAD.n9836 2.2505
R34454 PAD.n9835 PAD.n1563 2.2505
R34455 PAD.n9834 PAD.n9833 2.2505
R34456 PAD.n9829 PAD.n1564 2.2505
R34457 PAD.n9825 PAD.n9824 2.2505
R34458 PAD.n9823 PAD.n1565 2.2505
R34459 PAD.n9822 PAD.n9821 2.2505
R34460 PAD.n9817 PAD.n1566 2.2505
R34461 PAD.n9813 PAD.n9812 2.2505
R34462 PAD.n9811 PAD.n1567 2.2505
R34463 PAD.n9810 PAD.n9809 2.2505
R34464 PAD.n9805 PAD.n1568 2.2505
R34465 PAD.n9801 PAD.n9800 2.2505
R34466 PAD.n9799 PAD.n1569 2.2505
R34467 PAD.n9798 PAD.n9797 2.2505
R34468 PAD.n9793 PAD.n1570 2.2505
R34469 PAD.n9789 PAD.n9788 2.2505
R34470 PAD.n9787 PAD.n1571 2.2505
R34471 PAD.n9786 PAD.n9785 2.2505
R34472 PAD.n9781 PAD.n1572 2.2505
R34473 PAD.n9777 PAD.n9776 2.2505
R34474 PAD.n9775 PAD.n1573 2.2505
R34475 PAD.n9774 PAD.n9773 2.2505
R34476 PAD.n9769 PAD.n1574 2.2505
R34477 PAD.n9765 PAD.n9764 2.2505
R34478 PAD.n9763 PAD.n1575 2.2505
R34479 PAD.n9762 PAD.n9761 2.2505
R34480 PAD.n9757 PAD.n1576 2.2505
R34481 PAD.n9753 PAD.n9752 2.2505
R34482 PAD.n9751 PAD.n1579 2.2505
R34483 PAD.n9750 PAD.n9749 2.2505
R34484 PAD.n1931 PAD.n1599 2.2505
R34485 PAD.n1930 PAD.n1929 2.2505
R34486 PAD.n1927 PAD.n1600 2.2505
R34487 PAD.n1925 PAD.n1924 2.2505
R34488 PAD.n1917 PAD.n1603 2.2505
R34489 PAD.n1920 PAD.n1919 2.2505
R34490 PAD.n1915 PAD.n1606 2.2505
R34491 PAD.n1913 PAD.n1912 2.2505
R34492 PAD.n1905 PAD.n1608 2.2505
R34493 PAD.n1908 PAD.n1907 2.2505
R34494 PAD.n1903 PAD.n1610 2.2505
R34495 PAD.n1901 PAD.n1900 2.2505
R34496 PAD.n1893 PAD.n1612 2.2505
R34497 PAD.n1896 PAD.n1895 2.2505
R34498 PAD.n1891 PAD.n1614 2.2505
R34499 PAD.n1889 PAD.n1888 2.2505
R34500 PAD.n1881 PAD.n1616 2.2505
R34501 PAD.n1884 PAD.n1883 2.2505
R34502 PAD.n1879 PAD.n1618 2.2505
R34503 PAD.n1877 PAD.n1876 2.2505
R34504 PAD.n1869 PAD.n1620 2.2505
R34505 PAD.n1872 PAD.n1871 2.2505
R34506 PAD.n1867 PAD.n1622 2.2505
R34507 PAD.n1865 PAD.n1864 2.2505
R34508 PAD.n1857 PAD.n1624 2.2505
R34509 PAD.n1860 PAD.n1859 2.2505
R34510 PAD.n1855 PAD.n1626 2.2505
R34511 PAD.n1853 PAD.n1852 2.2505
R34512 PAD.n1845 PAD.n1628 2.2505
R34513 PAD.n1848 PAD.n1847 2.2505
R34514 PAD.n1843 PAD.n1630 2.2505
R34515 PAD.n1841 PAD.n1840 2.2505
R34516 PAD.n1833 PAD.n1632 2.2505
R34517 PAD.n1836 PAD.n1835 2.2505
R34518 PAD.n1831 PAD.n1634 2.2505
R34519 PAD.n1829 PAD.n1828 2.2505
R34520 PAD.n1821 PAD.n1636 2.2505
R34521 PAD.n1824 PAD.n1823 2.2505
R34522 PAD.n1819 PAD.n1638 2.2505
R34523 PAD.n1817 PAD.n1816 2.2505
R34524 PAD.n1809 PAD.n1640 2.2505
R34525 PAD.n1812 PAD.n1811 2.2505
R34526 PAD.n1807 PAD.n1642 2.2505
R34527 PAD.n1805 PAD.n1804 2.2505
R34528 PAD.n1797 PAD.n1644 2.2505
R34529 PAD.n1800 PAD.n1799 2.2505
R34530 PAD.n1795 PAD.n1646 2.2505
R34531 PAD.n1793 PAD.n1792 2.2505
R34532 PAD.n1785 PAD.n1648 2.2505
R34533 PAD.n1788 PAD.n1787 2.2505
R34534 PAD.n1783 PAD.n1650 2.2505
R34535 PAD.n1781 PAD.n1780 2.2505
R34536 PAD.n1773 PAD.n1652 2.2505
R34537 PAD.n1776 PAD.n1775 2.2505
R34538 PAD.n1771 PAD.n1654 2.2505
R34539 PAD.n1769 PAD.n1768 2.2505
R34540 PAD.n1761 PAD.n1656 2.2505
R34541 PAD.n1764 PAD.n1763 2.2505
R34542 PAD.n1759 PAD.n1658 2.2505
R34543 PAD.n1757 PAD.n1756 2.2505
R34544 PAD.n1749 PAD.n1660 2.2505
R34545 PAD.n1752 PAD.n1751 2.2505
R34546 PAD.n1747 PAD.n1662 2.2505
R34547 PAD.n1745 PAD.n1744 2.2505
R34548 PAD.n1737 PAD.n1664 2.2505
R34549 PAD.n1740 PAD.n1739 2.2505
R34550 PAD.n1735 PAD.n1666 2.2505
R34551 PAD.n1733 PAD.n1732 2.2505
R34552 PAD.n1725 PAD.n1668 2.2505
R34553 PAD.n1728 PAD.n1727 2.2505
R34554 PAD.n1723 PAD.n1670 2.2505
R34555 PAD.n1721 PAD.n1720 2.2505
R34556 PAD.n1713 PAD.n1672 2.2505
R34557 PAD.n1716 PAD.n1715 2.2505
R34558 PAD.n1711 PAD.n1674 2.2505
R34559 PAD.n1709 PAD.n1708 2.2505
R34560 PAD.n1701 PAD.n1676 2.2505
R34561 PAD.n1704 PAD.n1703 2.2505
R34562 PAD.n1699 PAD.n1678 2.2505
R34563 PAD.n1697 PAD.n1696 2.2505
R34564 PAD.n1689 PAD.n1680 2.2505
R34565 PAD.n1692 PAD.n1691 2.2505
R34566 PAD.n1687 PAD.n1682 2.2505
R34567 PAD.n1685 PAD.n1684 2.2505
R34568 PAD.n1684 PAD.n1683 2.2505
R34569 PAD.n1682 PAD.n1681 2.2505
R34570 PAD.n1693 PAD.n1692 2.2505
R34571 PAD.n1694 PAD.n1680 2.2505
R34572 PAD.n1696 PAD.n1695 2.2505
R34573 PAD.n1678 PAD.n1677 2.2505
R34574 PAD.n1705 PAD.n1704 2.2505
R34575 PAD.n1706 PAD.n1676 2.2505
R34576 PAD.n1708 PAD.n1707 2.2505
R34577 PAD.n1674 PAD.n1673 2.2505
R34578 PAD.n1717 PAD.n1716 2.2505
R34579 PAD.n1718 PAD.n1672 2.2505
R34580 PAD.n1720 PAD.n1719 2.2505
R34581 PAD.n1670 PAD.n1669 2.2505
R34582 PAD.n1729 PAD.n1728 2.2505
R34583 PAD.n1730 PAD.n1668 2.2505
R34584 PAD.n1732 PAD.n1731 2.2505
R34585 PAD.n1666 PAD.n1665 2.2505
R34586 PAD.n1741 PAD.n1740 2.2505
R34587 PAD.n1742 PAD.n1664 2.2505
R34588 PAD.n1744 PAD.n1743 2.2505
R34589 PAD.n1662 PAD.n1661 2.2505
R34590 PAD.n1753 PAD.n1752 2.2505
R34591 PAD.n1754 PAD.n1660 2.2505
R34592 PAD.n1756 PAD.n1755 2.2505
R34593 PAD.n1658 PAD.n1657 2.2505
R34594 PAD.n1765 PAD.n1764 2.2505
R34595 PAD.n1766 PAD.n1656 2.2505
R34596 PAD.n1768 PAD.n1767 2.2505
R34597 PAD.n1654 PAD.n1653 2.2505
R34598 PAD.n1777 PAD.n1776 2.2505
R34599 PAD.n1778 PAD.n1652 2.2505
R34600 PAD.n1780 PAD.n1779 2.2505
R34601 PAD.n1650 PAD.n1649 2.2505
R34602 PAD.n1789 PAD.n1788 2.2505
R34603 PAD.n1790 PAD.n1648 2.2505
R34604 PAD.n1792 PAD.n1791 2.2505
R34605 PAD.n1646 PAD.n1645 2.2505
R34606 PAD.n1801 PAD.n1800 2.2505
R34607 PAD.n1802 PAD.n1644 2.2505
R34608 PAD.n1804 PAD.n1803 2.2505
R34609 PAD.n1642 PAD.n1641 2.2505
R34610 PAD.n1813 PAD.n1812 2.2505
R34611 PAD.n1814 PAD.n1640 2.2505
R34612 PAD.n1816 PAD.n1815 2.2505
R34613 PAD.n1638 PAD.n1637 2.2505
R34614 PAD.n1825 PAD.n1824 2.2505
R34615 PAD.n1826 PAD.n1636 2.2505
R34616 PAD.n1828 PAD.n1827 2.2505
R34617 PAD.n1634 PAD.n1633 2.2505
R34618 PAD.n1837 PAD.n1836 2.2505
R34619 PAD.n1838 PAD.n1632 2.2505
R34620 PAD.n1840 PAD.n1839 2.2505
R34621 PAD.n1630 PAD.n1629 2.2505
R34622 PAD.n1849 PAD.n1848 2.2505
R34623 PAD.n1850 PAD.n1628 2.2505
R34624 PAD.n1852 PAD.n1851 2.2505
R34625 PAD.n1626 PAD.n1625 2.2505
R34626 PAD.n1861 PAD.n1860 2.2505
R34627 PAD.n1862 PAD.n1624 2.2505
R34628 PAD.n1864 PAD.n1863 2.2505
R34629 PAD.n1622 PAD.n1621 2.2505
R34630 PAD.n1873 PAD.n1872 2.2505
R34631 PAD.n1874 PAD.n1620 2.2505
R34632 PAD.n1876 PAD.n1875 2.2505
R34633 PAD.n1618 PAD.n1617 2.2505
R34634 PAD.n1885 PAD.n1884 2.2505
R34635 PAD.n1886 PAD.n1616 2.2505
R34636 PAD.n1888 PAD.n1887 2.2505
R34637 PAD.n1614 PAD.n1613 2.2505
R34638 PAD.n1897 PAD.n1896 2.2505
R34639 PAD.n1898 PAD.n1612 2.2505
R34640 PAD.n1900 PAD.n1899 2.2505
R34641 PAD.n1610 PAD.n1609 2.2505
R34642 PAD.n1909 PAD.n1908 2.2505
R34643 PAD.n1910 PAD.n1608 2.2505
R34644 PAD.n1912 PAD.n1911 2.2505
R34645 PAD.n1606 PAD.n1605 2.2505
R34646 PAD.n1921 PAD.n1920 2.2505
R34647 PAD.n1922 PAD.n1603 2.2505
R34648 PAD.n1924 PAD.n1923 2.2505
R34649 PAD.n1604 PAD.n1600 2.2505
R34650 PAD.n1930 PAD.n1598 2.2505
R34651 PAD.n1932 PAD.n1931 2.2505
R34652 PAD.n9463 PAD.n1984 2.2505
R34653 PAD.n2031 PAD.n2030 2.2505
R34654 PAD.n9468 PAD.n9467 2.2505
R34655 PAD.n9471 PAD.n9470 2.2505
R34656 PAD.n9475 PAD.n9474 2.2505
R34657 PAD.n9472 PAD.n2027 2.2505
R34658 PAD.n9480 PAD.n9479 2.2505
R34659 PAD.n9483 PAD.n9482 2.2505
R34660 PAD.n9487 PAD.n9486 2.2505
R34661 PAD.n9484 PAD.n2025 2.2505
R34662 PAD.n9492 PAD.n9491 2.2505
R34663 PAD.n9495 PAD.n9494 2.2505
R34664 PAD.n9499 PAD.n9498 2.2505
R34665 PAD.n9496 PAD.n2023 2.2505
R34666 PAD.n9504 PAD.n9503 2.2505
R34667 PAD.n9507 PAD.n9506 2.2505
R34668 PAD.n9511 PAD.n9510 2.2505
R34669 PAD.n9508 PAD.n2021 2.2505
R34670 PAD.n9516 PAD.n9515 2.2505
R34671 PAD.n9519 PAD.n9518 2.2505
R34672 PAD.n9523 PAD.n9522 2.2505
R34673 PAD.n9520 PAD.n2019 2.2505
R34674 PAD.n9528 PAD.n9527 2.2505
R34675 PAD.n9531 PAD.n9530 2.2505
R34676 PAD.n9535 PAD.n9534 2.2505
R34677 PAD.n9532 PAD.n2017 2.2505
R34678 PAD.n9540 PAD.n9539 2.2505
R34679 PAD.n9543 PAD.n9542 2.2505
R34680 PAD.n9547 PAD.n9546 2.2505
R34681 PAD.n9544 PAD.n2015 2.2505
R34682 PAD.n9552 PAD.n9551 2.2505
R34683 PAD.n9555 PAD.n9554 2.2505
R34684 PAD.n9559 PAD.n9558 2.2505
R34685 PAD.n9556 PAD.n2013 2.2505
R34686 PAD.n9564 PAD.n9563 2.2505
R34687 PAD.n9567 PAD.n9566 2.2505
R34688 PAD.n9571 PAD.n9570 2.2505
R34689 PAD.n9568 PAD.n2011 2.2505
R34690 PAD.n9576 PAD.n9575 2.2505
R34691 PAD.n9579 PAD.n9578 2.2505
R34692 PAD.n9583 PAD.n9582 2.2505
R34693 PAD.n9580 PAD.n2009 2.2505
R34694 PAD.n9588 PAD.n9587 2.2505
R34695 PAD.n9591 PAD.n9590 2.2505
R34696 PAD.n9595 PAD.n9594 2.2505
R34697 PAD.n9592 PAD.n2007 2.2505
R34698 PAD.n9600 PAD.n9599 2.2505
R34699 PAD.n9603 PAD.n9602 2.2505
R34700 PAD.n9607 PAD.n9606 2.2505
R34701 PAD.n9604 PAD.n2005 2.2505
R34702 PAD.n9612 PAD.n9611 2.2505
R34703 PAD.n9615 PAD.n9614 2.2505
R34704 PAD.n9619 PAD.n9618 2.2505
R34705 PAD.n9616 PAD.n2003 2.2505
R34706 PAD.n9624 PAD.n9623 2.2505
R34707 PAD.n9627 PAD.n9626 2.2505
R34708 PAD.n9631 PAD.n9630 2.2505
R34709 PAD.n9628 PAD.n2001 2.2505
R34710 PAD.n9636 PAD.n9635 2.2505
R34711 PAD.n9639 PAD.n9638 2.2505
R34712 PAD.n9643 PAD.n9642 2.2505
R34713 PAD.n9640 PAD.n1999 2.2505
R34714 PAD.n9648 PAD.n9647 2.2505
R34715 PAD.n9651 PAD.n9650 2.2505
R34716 PAD.n9655 PAD.n9654 2.2505
R34717 PAD.n9652 PAD.n1997 2.2505
R34718 PAD.n9660 PAD.n9659 2.2505
R34719 PAD.n9663 PAD.n9662 2.2505
R34720 PAD.n9667 PAD.n9666 2.2505
R34721 PAD.n9664 PAD.n1995 2.2505
R34722 PAD.n9672 PAD.n9671 2.2505
R34723 PAD.n9675 PAD.n9674 2.2505
R34724 PAD.n9679 PAD.n9678 2.2505
R34725 PAD.n9676 PAD.n1993 2.2505
R34726 PAD.n9684 PAD.n9683 2.2505
R34727 PAD.n9687 PAD.n9686 2.2505
R34728 PAD.n9691 PAD.n9690 2.2505
R34729 PAD.n9688 PAD.n1991 2.2505
R34730 PAD.n9696 PAD.n9695 2.2505
R34731 PAD.n9699 PAD.n9698 2.2505
R34732 PAD.n9703 PAD.n9702 2.2505
R34733 PAD.n9700 PAD.n1989 2.2505
R34734 PAD.n9709 PAD.n9708 2.2505
R34735 PAD.n9711 PAD.n1987 2.2505
R34736 PAD.n9706 PAD.n1987 2.2505
R34737 PAD.n9708 PAD.n9707 2.2505
R34738 PAD.n9705 PAD.n1989 2.2505
R34739 PAD.n9704 PAD.n9703 2.2505
R34740 PAD.n9699 PAD.n1990 2.2505
R34741 PAD.n9695 PAD.n9694 2.2505
R34742 PAD.n9693 PAD.n1991 2.2505
R34743 PAD.n9692 PAD.n9691 2.2505
R34744 PAD.n9687 PAD.n1992 2.2505
R34745 PAD.n9683 PAD.n9682 2.2505
R34746 PAD.n9681 PAD.n1993 2.2505
R34747 PAD.n9680 PAD.n9679 2.2505
R34748 PAD.n9675 PAD.n1994 2.2505
R34749 PAD.n9671 PAD.n9670 2.2505
R34750 PAD.n9669 PAD.n1995 2.2505
R34751 PAD.n9668 PAD.n9667 2.2505
R34752 PAD.n9663 PAD.n1996 2.2505
R34753 PAD.n9659 PAD.n9658 2.2505
R34754 PAD.n9657 PAD.n1997 2.2505
R34755 PAD.n9656 PAD.n9655 2.2505
R34756 PAD.n9651 PAD.n1998 2.2505
R34757 PAD.n9647 PAD.n9646 2.2505
R34758 PAD.n9645 PAD.n1999 2.2505
R34759 PAD.n9644 PAD.n9643 2.2505
R34760 PAD.n9639 PAD.n2000 2.2505
R34761 PAD.n9635 PAD.n9634 2.2505
R34762 PAD.n9633 PAD.n2001 2.2505
R34763 PAD.n9632 PAD.n9631 2.2505
R34764 PAD.n9627 PAD.n2002 2.2505
R34765 PAD.n9623 PAD.n9622 2.2505
R34766 PAD.n9621 PAD.n2003 2.2505
R34767 PAD.n9620 PAD.n9619 2.2505
R34768 PAD.n9615 PAD.n2004 2.2505
R34769 PAD.n9611 PAD.n9610 2.2505
R34770 PAD.n9609 PAD.n2005 2.2505
R34771 PAD.n9608 PAD.n9607 2.2505
R34772 PAD.n9603 PAD.n2006 2.2505
R34773 PAD.n9599 PAD.n9598 2.2505
R34774 PAD.n9597 PAD.n2007 2.2505
R34775 PAD.n9596 PAD.n9595 2.2505
R34776 PAD.n9591 PAD.n2008 2.2505
R34777 PAD.n9587 PAD.n9586 2.2505
R34778 PAD.n9585 PAD.n2009 2.2505
R34779 PAD.n9584 PAD.n9583 2.2505
R34780 PAD.n9579 PAD.n2010 2.2505
R34781 PAD.n9575 PAD.n9574 2.2505
R34782 PAD.n9573 PAD.n2011 2.2505
R34783 PAD.n9572 PAD.n9571 2.2505
R34784 PAD.n9567 PAD.n2012 2.2505
R34785 PAD.n9563 PAD.n9562 2.2505
R34786 PAD.n9561 PAD.n2013 2.2505
R34787 PAD.n9560 PAD.n9559 2.2505
R34788 PAD.n9555 PAD.n2014 2.2505
R34789 PAD.n9551 PAD.n9550 2.2505
R34790 PAD.n9549 PAD.n2015 2.2505
R34791 PAD.n9548 PAD.n9547 2.2505
R34792 PAD.n9543 PAD.n2016 2.2505
R34793 PAD.n9539 PAD.n9538 2.2505
R34794 PAD.n9537 PAD.n2017 2.2505
R34795 PAD.n9536 PAD.n9535 2.2505
R34796 PAD.n9531 PAD.n2018 2.2505
R34797 PAD.n9527 PAD.n9526 2.2505
R34798 PAD.n9525 PAD.n2019 2.2505
R34799 PAD.n9524 PAD.n9523 2.2505
R34800 PAD.n9519 PAD.n2020 2.2505
R34801 PAD.n9515 PAD.n9514 2.2505
R34802 PAD.n9513 PAD.n2021 2.2505
R34803 PAD.n9512 PAD.n9511 2.2505
R34804 PAD.n9507 PAD.n2022 2.2505
R34805 PAD.n9503 PAD.n9502 2.2505
R34806 PAD.n9501 PAD.n2023 2.2505
R34807 PAD.n9500 PAD.n9499 2.2505
R34808 PAD.n9495 PAD.n2024 2.2505
R34809 PAD.n9491 PAD.n9490 2.2505
R34810 PAD.n9489 PAD.n2025 2.2505
R34811 PAD.n9488 PAD.n9487 2.2505
R34812 PAD.n9483 PAD.n2026 2.2505
R34813 PAD.n9479 PAD.n9478 2.2505
R34814 PAD.n9477 PAD.n2027 2.2505
R34815 PAD.n9476 PAD.n9475 2.2505
R34816 PAD.n9471 PAD.n2028 2.2505
R34817 PAD.n9467 PAD.n9466 2.2505
R34818 PAD.n9465 PAD.n2031 2.2505
R34819 PAD.n9464 PAD.n9463 2.2505
R34820 PAD.n9197 PAD.n2088 2.2505
R34821 PAD.n2134 PAD.n2133 2.2505
R34822 PAD.n9202 PAD.n9201 2.2505
R34823 PAD.n9205 PAD.n9204 2.2505
R34824 PAD.n9209 PAD.n9208 2.2505
R34825 PAD.n9206 PAD.n2130 2.2505
R34826 PAD.n9214 PAD.n9213 2.2505
R34827 PAD.n9217 PAD.n9216 2.2505
R34828 PAD.n9221 PAD.n9220 2.2505
R34829 PAD.n9218 PAD.n2128 2.2505
R34830 PAD.n9226 PAD.n9225 2.2505
R34831 PAD.n9229 PAD.n9228 2.2505
R34832 PAD.n9233 PAD.n9232 2.2505
R34833 PAD.n9230 PAD.n2126 2.2505
R34834 PAD.n9238 PAD.n9237 2.2505
R34835 PAD.n9241 PAD.n9240 2.2505
R34836 PAD.n9245 PAD.n9244 2.2505
R34837 PAD.n9242 PAD.n2124 2.2505
R34838 PAD.n9250 PAD.n9249 2.2505
R34839 PAD.n9253 PAD.n9252 2.2505
R34840 PAD.n9257 PAD.n9256 2.2505
R34841 PAD.n9254 PAD.n2122 2.2505
R34842 PAD.n9262 PAD.n9261 2.2505
R34843 PAD.n9265 PAD.n9264 2.2505
R34844 PAD.n9269 PAD.n9268 2.2505
R34845 PAD.n9266 PAD.n2120 2.2505
R34846 PAD.n9274 PAD.n9273 2.2505
R34847 PAD.n9277 PAD.n9276 2.2505
R34848 PAD.n9281 PAD.n9280 2.2505
R34849 PAD.n9278 PAD.n2118 2.2505
R34850 PAD.n9286 PAD.n9285 2.2505
R34851 PAD.n9289 PAD.n9288 2.2505
R34852 PAD.n9293 PAD.n9292 2.2505
R34853 PAD.n9290 PAD.n2116 2.2505
R34854 PAD.n9298 PAD.n9297 2.2505
R34855 PAD.n9301 PAD.n9300 2.2505
R34856 PAD.n9305 PAD.n9304 2.2505
R34857 PAD.n9302 PAD.n2114 2.2505
R34858 PAD.n9310 PAD.n9309 2.2505
R34859 PAD.n9313 PAD.n9312 2.2505
R34860 PAD.n9317 PAD.n9316 2.2505
R34861 PAD.n9314 PAD.n2112 2.2505
R34862 PAD.n9322 PAD.n9321 2.2505
R34863 PAD.n9325 PAD.n9324 2.2505
R34864 PAD.n9329 PAD.n9328 2.2505
R34865 PAD.n9326 PAD.n2110 2.2505
R34866 PAD.n9334 PAD.n9333 2.2505
R34867 PAD.n9337 PAD.n9336 2.2505
R34868 PAD.n9341 PAD.n9340 2.2505
R34869 PAD.n9338 PAD.n2108 2.2505
R34870 PAD.n9346 PAD.n9345 2.2505
R34871 PAD.n9349 PAD.n9348 2.2505
R34872 PAD.n9353 PAD.n9352 2.2505
R34873 PAD.n9350 PAD.n2106 2.2505
R34874 PAD.n9358 PAD.n9357 2.2505
R34875 PAD.n9361 PAD.n9360 2.2505
R34876 PAD.n9365 PAD.n9364 2.2505
R34877 PAD.n9362 PAD.n2104 2.2505
R34878 PAD.n9370 PAD.n9369 2.2505
R34879 PAD.n9373 PAD.n9372 2.2505
R34880 PAD.n9377 PAD.n9376 2.2505
R34881 PAD.n9374 PAD.n2102 2.2505
R34882 PAD.n9382 PAD.n9381 2.2505
R34883 PAD.n9385 PAD.n9384 2.2505
R34884 PAD.n9389 PAD.n9388 2.2505
R34885 PAD.n9386 PAD.n2100 2.2505
R34886 PAD.n9394 PAD.n9393 2.2505
R34887 PAD.n9397 PAD.n9396 2.2505
R34888 PAD.n9401 PAD.n9400 2.2505
R34889 PAD.n9398 PAD.n2098 2.2505
R34890 PAD.n9406 PAD.n9405 2.2505
R34891 PAD.n9409 PAD.n9408 2.2505
R34892 PAD.n9413 PAD.n9412 2.2505
R34893 PAD.n9410 PAD.n2096 2.2505
R34894 PAD.n9418 PAD.n9417 2.2505
R34895 PAD.n9421 PAD.n9420 2.2505
R34896 PAD.n9425 PAD.n9424 2.2505
R34897 PAD.n9422 PAD.n2094 2.2505
R34898 PAD.n9430 PAD.n9429 2.2505
R34899 PAD.n9433 PAD.n9432 2.2505
R34900 PAD.n9437 PAD.n9436 2.2505
R34901 PAD.n9434 PAD.n2092 2.2505
R34902 PAD.n9442 PAD.n9441 2.2505
R34903 PAD.n9444 PAD.n2090 2.2505
R34904 PAD.n2090 PAD.n2040 2.2505
R34905 PAD.n9441 PAD.n9440 2.2505
R34906 PAD.n9439 PAD.n2092 2.2505
R34907 PAD.n9438 PAD.n9437 2.2505
R34908 PAD.n9433 PAD.n2093 2.2505
R34909 PAD.n9429 PAD.n9428 2.2505
R34910 PAD.n9427 PAD.n2094 2.2505
R34911 PAD.n9426 PAD.n9425 2.2505
R34912 PAD.n9421 PAD.n2095 2.2505
R34913 PAD.n9417 PAD.n9416 2.2505
R34914 PAD.n9415 PAD.n2096 2.2505
R34915 PAD.n9414 PAD.n9413 2.2505
R34916 PAD.n9409 PAD.n2097 2.2505
R34917 PAD.n9405 PAD.n9404 2.2505
R34918 PAD.n9403 PAD.n2098 2.2505
R34919 PAD.n9402 PAD.n9401 2.2505
R34920 PAD.n9397 PAD.n2099 2.2505
R34921 PAD.n9393 PAD.n9392 2.2505
R34922 PAD.n9391 PAD.n2100 2.2505
R34923 PAD.n9390 PAD.n9389 2.2505
R34924 PAD.n9385 PAD.n2101 2.2505
R34925 PAD.n9381 PAD.n9380 2.2505
R34926 PAD.n9379 PAD.n2102 2.2505
R34927 PAD.n9378 PAD.n9377 2.2505
R34928 PAD.n9373 PAD.n2103 2.2505
R34929 PAD.n9369 PAD.n9368 2.2505
R34930 PAD.n9367 PAD.n2104 2.2505
R34931 PAD.n9366 PAD.n9365 2.2505
R34932 PAD.n9361 PAD.n2105 2.2505
R34933 PAD.n9357 PAD.n9356 2.2505
R34934 PAD.n9355 PAD.n2106 2.2505
R34935 PAD.n9354 PAD.n9353 2.2505
R34936 PAD.n9349 PAD.n2107 2.2505
R34937 PAD.n9345 PAD.n9344 2.2505
R34938 PAD.n9343 PAD.n2108 2.2505
R34939 PAD.n9342 PAD.n9341 2.2505
R34940 PAD.n9337 PAD.n2109 2.2505
R34941 PAD.n9333 PAD.n9332 2.2505
R34942 PAD.n9331 PAD.n2110 2.2505
R34943 PAD.n9330 PAD.n9329 2.2505
R34944 PAD.n9325 PAD.n2111 2.2505
R34945 PAD.n9321 PAD.n9320 2.2505
R34946 PAD.n9319 PAD.n2112 2.2505
R34947 PAD.n9318 PAD.n9317 2.2505
R34948 PAD.n9313 PAD.n2113 2.2505
R34949 PAD.n9309 PAD.n9308 2.2505
R34950 PAD.n9307 PAD.n2114 2.2505
R34951 PAD.n9306 PAD.n9305 2.2505
R34952 PAD.n9301 PAD.n2115 2.2505
R34953 PAD.n9297 PAD.n9296 2.2505
R34954 PAD.n9295 PAD.n2116 2.2505
R34955 PAD.n9294 PAD.n9293 2.2505
R34956 PAD.n9289 PAD.n2117 2.2505
R34957 PAD.n9285 PAD.n9284 2.2505
R34958 PAD.n9283 PAD.n2118 2.2505
R34959 PAD.n9282 PAD.n9281 2.2505
R34960 PAD.n9277 PAD.n2119 2.2505
R34961 PAD.n9273 PAD.n9272 2.2505
R34962 PAD.n9271 PAD.n2120 2.2505
R34963 PAD.n9270 PAD.n9269 2.2505
R34964 PAD.n9265 PAD.n2121 2.2505
R34965 PAD.n9261 PAD.n9260 2.2505
R34966 PAD.n9259 PAD.n2122 2.2505
R34967 PAD.n9258 PAD.n9257 2.2505
R34968 PAD.n9253 PAD.n2123 2.2505
R34969 PAD.n9249 PAD.n9248 2.2505
R34970 PAD.n9247 PAD.n2124 2.2505
R34971 PAD.n9246 PAD.n9245 2.2505
R34972 PAD.n9241 PAD.n2125 2.2505
R34973 PAD.n9237 PAD.n9236 2.2505
R34974 PAD.n9235 PAD.n2126 2.2505
R34975 PAD.n9234 PAD.n9233 2.2505
R34976 PAD.n9229 PAD.n2127 2.2505
R34977 PAD.n9225 PAD.n9224 2.2505
R34978 PAD.n9223 PAD.n2128 2.2505
R34979 PAD.n9222 PAD.n9221 2.2505
R34980 PAD.n9217 PAD.n2129 2.2505
R34981 PAD.n9213 PAD.n9212 2.2505
R34982 PAD.n9211 PAD.n2130 2.2505
R34983 PAD.n9210 PAD.n9209 2.2505
R34984 PAD.n9205 PAD.n2131 2.2505
R34985 PAD.n9201 PAD.n9200 2.2505
R34986 PAD.n9199 PAD.n2134 2.2505
R34987 PAD.n9198 PAD.n9197 2.2505
R34988 PAD.n2482 PAD.n2151 2.2505
R34989 PAD.n2481 PAD.n2480 2.2505
R34990 PAD.n2478 PAD.n2152 2.2505
R34991 PAD.n2476 PAD.n2475 2.2505
R34992 PAD.n2468 PAD.n2155 2.2505
R34993 PAD.n2471 PAD.n2470 2.2505
R34994 PAD.n2466 PAD.n2158 2.2505
R34995 PAD.n2464 PAD.n2463 2.2505
R34996 PAD.n2456 PAD.n2160 2.2505
R34997 PAD.n2459 PAD.n2458 2.2505
R34998 PAD.n2454 PAD.n2162 2.2505
R34999 PAD.n2452 PAD.n2451 2.2505
R35000 PAD.n2444 PAD.n2164 2.2505
R35001 PAD.n2447 PAD.n2446 2.2505
R35002 PAD.n2442 PAD.n2166 2.2505
R35003 PAD.n2440 PAD.n2439 2.2505
R35004 PAD.n2432 PAD.n2168 2.2505
R35005 PAD.n2435 PAD.n2434 2.2505
R35006 PAD.n2430 PAD.n2170 2.2505
R35007 PAD.n2428 PAD.n2427 2.2505
R35008 PAD.n2420 PAD.n2172 2.2505
R35009 PAD.n2423 PAD.n2422 2.2505
R35010 PAD.n2418 PAD.n2174 2.2505
R35011 PAD.n2416 PAD.n2415 2.2505
R35012 PAD.n2408 PAD.n2176 2.2505
R35013 PAD.n2411 PAD.n2410 2.2505
R35014 PAD.n2406 PAD.n2178 2.2505
R35015 PAD.n2404 PAD.n2403 2.2505
R35016 PAD.n2396 PAD.n2180 2.2505
R35017 PAD.n2399 PAD.n2398 2.2505
R35018 PAD.n2394 PAD.n2182 2.2505
R35019 PAD.n2392 PAD.n2391 2.2505
R35020 PAD.n2384 PAD.n2184 2.2505
R35021 PAD.n2387 PAD.n2386 2.2505
R35022 PAD.n2382 PAD.n2186 2.2505
R35023 PAD.n2380 PAD.n2379 2.2505
R35024 PAD.n2372 PAD.n2188 2.2505
R35025 PAD.n2375 PAD.n2374 2.2505
R35026 PAD.n2370 PAD.n2190 2.2505
R35027 PAD.n2368 PAD.n2367 2.2505
R35028 PAD.n2360 PAD.n2192 2.2505
R35029 PAD.n2363 PAD.n2362 2.2505
R35030 PAD.n2358 PAD.n2194 2.2505
R35031 PAD.n2356 PAD.n2355 2.2505
R35032 PAD.n2348 PAD.n2196 2.2505
R35033 PAD.n2351 PAD.n2350 2.2505
R35034 PAD.n2346 PAD.n2198 2.2505
R35035 PAD.n2344 PAD.n2343 2.2505
R35036 PAD.n2336 PAD.n2200 2.2505
R35037 PAD.n2339 PAD.n2338 2.2505
R35038 PAD.n2334 PAD.n2202 2.2505
R35039 PAD.n2332 PAD.n2331 2.2505
R35040 PAD.n2324 PAD.n2204 2.2505
R35041 PAD.n2327 PAD.n2326 2.2505
R35042 PAD.n2322 PAD.n2206 2.2505
R35043 PAD.n2320 PAD.n2319 2.2505
R35044 PAD.n2312 PAD.n2208 2.2505
R35045 PAD.n2315 PAD.n2314 2.2505
R35046 PAD.n2310 PAD.n2210 2.2505
R35047 PAD.n2308 PAD.n2307 2.2505
R35048 PAD.n2300 PAD.n2212 2.2505
R35049 PAD.n2303 PAD.n2302 2.2505
R35050 PAD.n2298 PAD.n2214 2.2505
R35051 PAD.n2296 PAD.n2295 2.2505
R35052 PAD.n2288 PAD.n2216 2.2505
R35053 PAD.n2291 PAD.n2290 2.2505
R35054 PAD.n2286 PAD.n2218 2.2505
R35055 PAD.n2284 PAD.n2283 2.2505
R35056 PAD.n2276 PAD.n2220 2.2505
R35057 PAD.n2279 PAD.n2278 2.2505
R35058 PAD.n2274 PAD.n2222 2.2505
R35059 PAD.n2272 PAD.n2271 2.2505
R35060 PAD.n2264 PAD.n2224 2.2505
R35061 PAD.n2267 PAD.n2266 2.2505
R35062 PAD.n2262 PAD.n2226 2.2505
R35063 PAD.n2260 PAD.n2259 2.2505
R35064 PAD.n2252 PAD.n2228 2.2505
R35065 PAD.n2255 PAD.n2254 2.2505
R35066 PAD.n2250 PAD.n2230 2.2505
R35067 PAD.n2248 PAD.n2247 2.2505
R35068 PAD.n2240 PAD.n2232 2.2505
R35069 PAD.n2243 PAD.n2242 2.2505
R35070 PAD.n2238 PAD.n2234 2.2505
R35071 PAD.n2236 PAD.n2235 2.2505
R35072 PAD.n2235 PAD.n2142 2.2505
R35073 PAD.n2234 PAD.n2233 2.2505
R35074 PAD.n2244 PAD.n2243 2.2505
R35075 PAD.n2245 PAD.n2232 2.2505
R35076 PAD.n2247 PAD.n2246 2.2505
R35077 PAD.n2230 PAD.n2229 2.2505
R35078 PAD.n2256 PAD.n2255 2.2505
R35079 PAD.n2257 PAD.n2228 2.2505
R35080 PAD.n2259 PAD.n2258 2.2505
R35081 PAD.n2226 PAD.n2225 2.2505
R35082 PAD.n2268 PAD.n2267 2.2505
R35083 PAD.n2269 PAD.n2224 2.2505
R35084 PAD.n2271 PAD.n2270 2.2505
R35085 PAD.n2222 PAD.n2221 2.2505
R35086 PAD.n2280 PAD.n2279 2.2505
R35087 PAD.n2281 PAD.n2220 2.2505
R35088 PAD.n2283 PAD.n2282 2.2505
R35089 PAD.n2218 PAD.n2217 2.2505
R35090 PAD.n2292 PAD.n2291 2.2505
R35091 PAD.n2293 PAD.n2216 2.2505
R35092 PAD.n2295 PAD.n2294 2.2505
R35093 PAD.n2214 PAD.n2213 2.2505
R35094 PAD.n2304 PAD.n2303 2.2505
R35095 PAD.n2305 PAD.n2212 2.2505
R35096 PAD.n2307 PAD.n2306 2.2505
R35097 PAD.n2210 PAD.n2209 2.2505
R35098 PAD.n2316 PAD.n2315 2.2505
R35099 PAD.n2317 PAD.n2208 2.2505
R35100 PAD.n2319 PAD.n2318 2.2505
R35101 PAD.n2206 PAD.n2205 2.2505
R35102 PAD.n2328 PAD.n2327 2.2505
R35103 PAD.n2329 PAD.n2204 2.2505
R35104 PAD.n2331 PAD.n2330 2.2505
R35105 PAD.n2202 PAD.n2201 2.2505
R35106 PAD.n2340 PAD.n2339 2.2505
R35107 PAD.n2341 PAD.n2200 2.2505
R35108 PAD.n2343 PAD.n2342 2.2505
R35109 PAD.n2198 PAD.n2197 2.2505
R35110 PAD.n2352 PAD.n2351 2.2505
R35111 PAD.n2353 PAD.n2196 2.2505
R35112 PAD.n2355 PAD.n2354 2.2505
R35113 PAD.n2194 PAD.n2193 2.2505
R35114 PAD.n2364 PAD.n2363 2.2505
R35115 PAD.n2365 PAD.n2192 2.2505
R35116 PAD.n2367 PAD.n2366 2.2505
R35117 PAD.n2190 PAD.n2189 2.2505
R35118 PAD.n2376 PAD.n2375 2.2505
R35119 PAD.n2377 PAD.n2188 2.2505
R35120 PAD.n2379 PAD.n2378 2.2505
R35121 PAD.n2186 PAD.n2185 2.2505
R35122 PAD.n2388 PAD.n2387 2.2505
R35123 PAD.n2389 PAD.n2184 2.2505
R35124 PAD.n2391 PAD.n2390 2.2505
R35125 PAD.n2182 PAD.n2181 2.2505
R35126 PAD.n2400 PAD.n2399 2.2505
R35127 PAD.n2401 PAD.n2180 2.2505
R35128 PAD.n2403 PAD.n2402 2.2505
R35129 PAD.n2178 PAD.n2177 2.2505
R35130 PAD.n2412 PAD.n2411 2.2505
R35131 PAD.n2413 PAD.n2176 2.2505
R35132 PAD.n2415 PAD.n2414 2.2505
R35133 PAD.n2174 PAD.n2173 2.2505
R35134 PAD.n2424 PAD.n2423 2.2505
R35135 PAD.n2425 PAD.n2172 2.2505
R35136 PAD.n2427 PAD.n2426 2.2505
R35137 PAD.n2170 PAD.n2169 2.2505
R35138 PAD.n2436 PAD.n2435 2.2505
R35139 PAD.n2437 PAD.n2168 2.2505
R35140 PAD.n2439 PAD.n2438 2.2505
R35141 PAD.n2166 PAD.n2165 2.2505
R35142 PAD.n2448 PAD.n2447 2.2505
R35143 PAD.n2449 PAD.n2164 2.2505
R35144 PAD.n2451 PAD.n2450 2.2505
R35145 PAD.n2162 PAD.n2161 2.2505
R35146 PAD.n2460 PAD.n2459 2.2505
R35147 PAD.n2461 PAD.n2160 2.2505
R35148 PAD.n2463 PAD.n2462 2.2505
R35149 PAD.n2158 PAD.n2157 2.2505
R35150 PAD.n2472 PAD.n2471 2.2505
R35151 PAD.n2473 PAD.n2155 2.2505
R35152 PAD.n2475 PAD.n2474 2.2505
R35153 PAD.n2156 PAD.n2152 2.2505
R35154 PAD.n2481 PAD.n2150 2.2505
R35155 PAD.n2483 PAD.n2482 2.2505
R35156 PAD.n2829 PAD.n2498 2.2505
R35157 PAD.n2828 PAD.n2827 2.2505
R35158 PAD.n2825 PAD.n2499 2.2505
R35159 PAD.n2823 PAD.n2822 2.2505
R35160 PAD.n2815 PAD.n2502 2.2505
R35161 PAD.n2818 PAD.n2817 2.2505
R35162 PAD.n2813 PAD.n2505 2.2505
R35163 PAD.n2811 PAD.n2810 2.2505
R35164 PAD.n2803 PAD.n2507 2.2505
R35165 PAD.n2806 PAD.n2805 2.2505
R35166 PAD.n2801 PAD.n2509 2.2505
R35167 PAD.n2799 PAD.n2798 2.2505
R35168 PAD.n2791 PAD.n2511 2.2505
R35169 PAD.n2794 PAD.n2793 2.2505
R35170 PAD.n2789 PAD.n2513 2.2505
R35171 PAD.n2787 PAD.n2786 2.2505
R35172 PAD.n2779 PAD.n2515 2.2505
R35173 PAD.n2782 PAD.n2781 2.2505
R35174 PAD.n2777 PAD.n2517 2.2505
R35175 PAD.n2775 PAD.n2774 2.2505
R35176 PAD.n2767 PAD.n2519 2.2505
R35177 PAD.n2770 PAD.n2769 2.2505
R35178 PAD.n2765 PAD.n2521 2.2505
R35179 PAD.n2763 PAD.n2762 2.2505
R35180 PAD.n2755 PAD.n2523 2.2505
R35181 PAD.n2758 PAD.n2757 2.2505
R35182 PAD.n2753 PAD.n2525 2.2505
R35183 PAD.n2751 PAD.n2750 2.2505
R35184 PAD.n2743 PAD.n2527 2.2505
R35185 PAD.n2746 PAD.n2745 2.2505
R35186 PAD.n2741 PAD.n2529 2.2505
R35187 PAD.n2739 PAD.n2738 2.2505
R35188 PAD.n2731 PAD.n2531 2.2505
R35189 PAD.n2734 PAD.n2733 2.2505
R35190 PAD.n2729 PAD.n2533 2.2505
R35191 PAD.n2727 PAD.n2726 2.2505
R35192 PAD.n2719 PAD.n2535 2.2505
R35193 PAD.n2722 PAD.n2721 2.2505
R35194 PAD.n2717 PAD.n2537 2.2505
R35195 PAD.n2715 PAD.n2714 2.2505
R35196 PAD.n2707 PAD.n2539 2.2505
R35197 PAD.n2710 PAD.n2709 2.2505
R35198 PAD.n2705 PAD.n2541 2.2505
R35199 PAD.n2703 PAD.n2702 2.2505
R35200 PAD.n2695 PAD.n2543 2.2505
R35201 PAD.n2698 PAD.n2697 2.2505
R35202 PAD.n2693 PAD.n2545 2.2505
R35203 PAD.n2691 PAD.n2690 2.2505
R35204 PAD.n2683 PAD.n2547 2.2505
R35205 PAD.n2686 PAD.n2685 2.2505
R35206 PAD.n2681 PAD.n2549 2.2505
R35207 PAD.n2679 PAD.n2678 2.2505
R35208 PAD.n2671 PAD.n2551 2.2505
R35209 PAD.n2674 PAD.n2673 2.2505
R35210 PAD.n2669 PAD.n2553 2.2505
R35211 PAD.n2667 PAD.n2666 2.2505
R35212 PAD.n2659 PAD.n2555 2.2505
R35213 PAD.n2662 PAD.n2661 2.2505
R35214 PAD.n2657 PAD.n2557 2.2505
R35215 PAD.n2655 PAD.n2654 2.2505
R35216 PAD.n2647 PAD.n2559 2.2505
R35217 PAD.n2650 PAD.n2649 2.2505
R35218 PAD.n2645 PAD.n2561 2.2505
R35219 PAD.n2643 PAD.n2642 2.2505
R35220 PAD.n2635 PAD.n2563 2.2505
R35221 PAD.n2638 PAD.n2637 2.2505
R35222 PAD.n2633 PAD.n2565 2.2505
R35223 PAD.n2631 PAD.n2630 2.2505
R35224 PAD.n2623 PAD.n2567 2.2505
R35225 PAD.n2626 PAD.n2625 2.2505
R35226 PAD.n2621 PAD.n2569 2.2505
R35227 PAD.n2619 PAD.n2618 2.2505
R35228 PAD.n2611 PAD.n2571 2.2505
R35229 PAD.n2614 PAD.n2613 2.2505
R35230 PAD.n2609 PAD.n2573 2.2505
R35231 PAD.n2607 PAD.n2606 2.2505
R35232 PAD.n2599 PAD.n2575 2.2505
R35233 PAD.n2602 PAD.n2601 2.2505
R35234 PAD.n2597 PAD.n2577 2.2505
R35235 PAD.n2595 PAD.n2594 2.2505
R35236 PAD.n2587 PAD.n2579 2.2505
R35237 PAD.n2590 PAD.n2589 2.2505
R35238 PAD.n2585 PAD.n2581 2.2505
R35239 PAD.n2583 PAD.n2582 2.2505
R35240 PAD.n2582 PAD.n2490 2.2505
R35241 PAD.n2581 PAD.n2580 2.2505
R35242 PAD.n2591 PAD.n2590 2.2505
R35243 PAD.n2592 PAD.n2579 2.2505
R35244 PAD.n2594 PAD.n2593 2.2505
R35245 PAD.n2577 PAD.n2576 2.2505
R35246 PAD.n2603 PAD.n2602 2.2505
R35247 PAD.n2604 PAD.n2575 2.2505
R35248 PAD.n2606 PAD.n2605 2.2505
R35249 PAD.n2573 PAD.n2572 2.2505
R35250 PAD.n2615 PAD.n2614 2.2505
R35251 PAD.n2616 PAD.n2571 2.2505
R35252 PAD.n2618 PAD.n2617 2.2505
R35253 PAD.n2569 PAD.n2568 2.2505
R35254 PAD.n2627 PAD.n2626 2.2505
R35255 PAD.n2628 PAD.n2567 2.2505
R35256 PAD.n2630 PAD.n2629 2.2505
R35257 PAD.n2565 PAD.n2564 2.2505
R35258 PAD.n2639 PAD.n2638 2.2505
R35259 PAD.n2640 PAD.n2563 2.2505
R35260 PAD.n2642 PAD.n2641 2.2505
R35261 PAD.n2561 PAD.n2560 2.2505
R35262 PAD.n2651 PAD.n2650 2.2505
R35263 PAD.n2652 PAD.n2559 2.2505
R35264 PAD.n2654 PAD.n2653 2.2505
R35265 PAD.n2557 PAD.n2556 2.2505
R35266 PAD.n2663 PAD.n2662 2.2505
R35267 PAD.n2664 PAD.n2555 2.2505
R35268 PAD.n2666 PAD.n2665 2.2505
R35269 PAD.n2553 PAD.n2552 2.2505
R35270 PAD.n2675 PAD.n2674 2.2505
R35271 PAD.n2676 PAD.n2551 2.2505
R35272 PAD.n2678 PAD.n2677 2.2505
R35273 PAD.n2549 PAD.n2548 2.2505
R35274 PAD.n2687 PAD.n2686 2.2505
R35275 PAD.n2688 PAD.n2547 2.2505
R35276 PAD.n2690 PAD.n2689 2.2505
R35277 PAD.n2545 PAD.n2544 2.2505
R35278 PAD.n2699 PAD.n2698 2.2505
R35279 PAD.n2700 PAD.n2543 2.2505
R35280 PAD.n2702 PAD.n2701 2.2505
R35281 PAD.n2541 PAD.n2540 2.2505
R35282 PAD.n2711 PAD.n2710 2.2505
R35283 PAD.n2712 PAD.n2539 2.2505
R35284 PAD.n2714 PAD.n2713 2.2505
R35285 PAD.n2537 PAD.n2536 2.2505
R35286 PAD.n2723 PAD.n2722 2.2505
R35287 PAD.n2724 PAD.n2535 2.2505
R35288 PAD.n2726 PAD.n2725 2.2505
R35289 PAD.n2533 PAD.n2532 2.2505
R35290 PAD.n2735 PAD.n2734 2.2505
R35291 PAD.n2736 PAD.n2531 2.2505
R35292 PAD.n2738 PAD.n2737 2.2505
R35293 PAD.n2529 PAD.n2528 2.2505
R35294 PAD.n2747 PAD.n2746 2.2505
R35295 PAD.n2748 PAD.n2527 2.2505
R35296 PAD.n2750 PAD.n2749 2.2505
R35297 PAD.n2525 PAD.n2524 2.2505
R35298 PAD.n2759 PAD.n2758 2.2505
R35299 PAD.n2760 PAD.n2523 2.2505
R35300 PAD.n2762 PAD.n2761 2.2505
R35301 PAD.n2521 PAD.n2520 2.2505
R35302 PAD.n2771 PAD.n2770 2.2505
R35303 PAD.n2772 PAD.n2519 2.2505
R35304 PAD.n2774 PAD.n2773 2.2505
R35305 PAD.n2517 PAD.n2516 2.2505
R35306 PAD.n2783 PAD.n2782 2.2505
R35307 PAD.n2784 PAD.n2515 2.2505
R35308 PAD.n2786 PAD.n2785 2.2505
R35309 PAD.n2513 PAD.n2512 2.2505
R35310 PAD.n2795 PAD.n2794 2.2505
R35311 PAD.n2796 PAD.n2511 2.2505
R35312 PAD.n2798 PAD.n2797 2.2505
R35313 PAD.n2509 PAD.n2508 2.2505
R35314 PAD.n2807 PAD.n2806 2.2505
R35315 PAD.n2808 PAD.n2507 2.2505
R35316 PAD.n2810 PAD.n2809 2.2505
R35317 PAD.n2505 PAD.n2504 2.2505
R35318 PAD.n2819 PAD.n2818 2.2505
R35319 PAD.n2820 PAD.n2502 2.2505
R35320 PAD.n2822 PAD.n2821 2.2505
R35321 PAD.n2503 PAD.n2499 2.2505
R35322 PAD.n2828 PAD.n2497 2.2505
R35323 PAD.n2830 PAD.n2829 2.2505
R35324 PAD.n9119 PAD.n2876 2.2505
R35325 PAD.n9118 PAD.n9117 2.2505
R35326 PAD.n9115 PAD.n8841 2.2505
R35327 PAD.n8839 PAD.n8838 2.2505
R35328 PAD.n9111 PAD.n9110 2.2505
R35329 PAD.n9108 PAD.n9107 2.2505
R35330 PAD.n9106 PAD.n8846 2.2505
R35331 PAD.n8844 PAD.n8843 2.2505
R35332 PAD.n9102 PAD.n9101 2.2505
R35333 PAD.n9099 PAD.n9098 2.2505
R35334 PAD.n9097 PAD.n8851 2.2505
R35335 PAD.n8849 PAD.n8848 2.2505
R35336 PAD.n9093 PAD.n9092 2.2505
R35337 PAD.n9090 PAD.n9089 2.2505
R35338 PAD.n9088 PAD.n8856 2.2505
R35339 PAD.n8854 PAD.n8853 2.2505
R35340 PAD.n9084 PAD.n9083 2.2505
R35341 PAD.n9081 PAD.n9080 2.2505
R35342 PAD.n9079 PAD.n8861 2.2505
R35343 PAD.n8859 PAD.n8858 2.2505
R35344 PAD.n9075 PAD.n9074 2.2505
R35345 PAD.n9072 PAD.n9071 2.2505
R35346 PAD.n9070 PAD.n8866 2.2505
R35347 PAD.n8864 PAD.n8863 2.2505
R35348 PAD.n9066 PAD.n9065 2.2505
R35349 PAD.n9063 PAD.n9062 2.2505
R35350 PAD.n9061 PAD.n8871 2.2505
R35351 PAD.n8869 PAD.n8868 2.2505
R35352 PAD.n9057 PAD.n9056 2.2505
R35353 PAD.n9054 PAD.n9053 2.2505
R35354 PAD.n9052 PAD.n8876 2.2505
R35355 PAD.n8874 PAD.n8873 2.2505
R35356 PAD.n9048 PAD.n9047 2.2505
R35357 PAD.n9045 PAD.n9044 2.2505
R35358 PAD.n9043 PAD.n8881 2.2505
R35359 PAD.n8879 PAD.n8878 2.2505
R35360 PAD.n9039 PAD.n9038 2.2505
R35361 PAD.n9036 PAD.n9035 2.2505
R35362 PAD.n9034 PAD.n8886 2.2505
R35363 PAD.n8884 PAD.n8883 2.2505
R35364 PAD.n9030 PAD.n9029 2.2505
R35365 PAD.n9027 PAD.n9026 2.2505
R35366 PAD.n9025 PAD.n8891 2.2505
R35367 PAD.n8889 PAD.n8888 2.2505
R35368 PAD.n9021 PAD.n9020 2.2505
R35369 PAD.n9018 PAD.n9017 2.2505
R35370 PAD.n9016 PAD.n8896 2.2505
R35371 PAD.n8894 PAD.n8893 2.2505
R35372 PAD.n9012 PAD.n9011 2.2505
R35373 PAD.n9009 PAD.n9008 2.2505
R35374 PAD.n9007 PAD.n8901 2.2505
R35375 PAD.n8899 PAD.n8898 2.2505
R35376 PAD.n9003 PAD.n9002 2.2505
R35377 PAD.n9000 PAD.n8999 2.2505
R35378 PAD.n8998 PAD.n8906 2.2505
R35379 PAD.n8904 PAD.n8903 2.2505
R35380 PAD.n8994 PAD.n8993 2.2505
R35381 PAD.n8991 PAD.n8990 2.2505
R35382 PAD.n8989 PAD.n8911 2.2505
R35383 PAD.n8909 PAD.n8908 2.2505
R35384 PAD.n8985 PAD.n8984 2.2505
R35385 PAD.n8982 PAD.n8981 2.2505
R35386 PAD.n8980 PAD.n8916 2.2505
R35387 PAD.n8914 PAD.n8913 2.2505
R35388 PAD.n8976 PAD.n8975 2.2505
R35389 PAD.n8973 PAD.n8972 2.2505
R35390 PAD.n8971 PAD.n8921 2.2505
R35391 PAD.n8919 PAD.n8918 2.2505
R35392 PAD.n8967 PAD.n8966 2.2505
R35393 PAD.n8964 PAD.n8963 2.2505
R35394 PAD.n8962 PAD.n8926 2.2505
R35395 PAD.n8924 PAD.n8923 2.2505
R35396 PAD.n8958 PAD.n8957 2.2505
R35397 PAD.n8955 PAD.n8954 2.2505
R35398 PAD.n8953 PAD.n8931 2.2505
R35399 PAD.n8929 PAD.n8928 2.2505
R35400 PAD.n8949 PAD.n8948 2.2505
R35401 PAD.n8946 PAD.n8945 2.2505
R35402 PAD.n8944 PAD.n8936 2.2505
R35403 PAD.n8934 PAD.n8933 2.2505
R35404 PAD.n8940 PAD.n8939 2.2505
R35405 PAD.n8937 PAD.n2880 2.2505
R35406 PAD.n9137 PAD.n9136 2.2505
R35407 PAD.n9139 PAD.n2877 2.2505
R35408 PAD.n9134 PAD.n2877 2.2505
R35409 PAD.n9136 PAD.n9135 2.2505
R35410 PAD.n2881 PAD.n2880 2.2505
R35411 PAD.n8941 PAD.n8940 2.2505
R35412 PAD.n8942 PAD.n8933 2.2505
R35413 PAD.n8944 PAD.n8943 2.2505
R35414 PAD.n8945 PAD.n8932 2.2505
R35415 PAD.n8950 PAD.n8949 2.2505
R35416 PAD.n8951 PAD.n8928 2.2505
R35417 PAD.n8953 PAD.n8952 2.2505
R35418 PAD.n8954 PAD.n8927 2.2505
R35419 PAD.n8959 PAD.n8958 2.2505
R35420 PAD.n8960 PAD.n8923 2.2505
R35421 PAD.n8962 PAD.n8961 2.2505
R35422 PAD.n8963 PAD.n8922 2.2505
R35423 PAD.n8968 PAD.n8967 2.2505
R35424 PAD.n8969 PAD.n8918 2.2505
R35425 PAD.n8971 PAD.n8970 2.2505
R35426 PAD.n8972 PAD.n8917 2.2505
R35427 PAD.n8977 PAD.n8976 2.2505
R35428 PAD.n8978 PAD.n8913 2.2505
R35429 PAD.n8980 PAD.n8979 2.2505
R35430 PAD.n8981 PAD.n8912 2.2505
R35431 PAD.n8986 PAD.n8985 2.2505
R35432 PAD.n8987 PAD.n8908 2.2505
R35433 PAD.n8989 PAD.n8988 2.2505
R35434 PAD.n8990 PAD.n8907 2.2505
R35435 PAD.n8995 PAD.n8994 2.2505
R35436 PAD.n8996 PAD.n8903 2.2505
R35437 PAD.n8998 PAD.n8997 2.2505
R35438 PAD.n8999 PAD.n8902 2.2505
R35439 PAD.n9004 PAD.n9003 2.2505
R35440 PAD.n9005 PAD.n8898 2.2505
R35441 PAD.n9007 PAD.n9006 2.2505
R35442 PAD.n9008 PAD.n8897 2.2505
R35443 PAD.n9013 PAD.n9012 2.2505
R35444 PAD.n9014 PAD.n8893 2.2505
R35445 PAD.n9016 PAD.n9015 2.2505
R35446 PAD.n9017 PAD.n8892 2.2505
R35447 PAD.n9022 PAD.n9021 2.2505
R35448 PAD.n9023 PAD.n8888 2.2505
R35449 PAD.n9025 PAD.n9024 2.2505
R35450 PAD.n9026 PAD.n8887 2.2505
R35451 PAD.n9031 PAD.n9030 2.2505
R35452 PAD.n9032 PAD.n8883 2.2505
R35453 PAD.n9034 PAD.n9033 2.2505
R35454 PAD.n9035 PAD.n8882 2.2505
R35455 PAD.n9040 PAD.n9039 2.2505
R35456 PAD.n9041 PAD.n8878 2.2505
R35457 PAD.n9043 PAD.n9042 2.2505
R35458 PAD.n9044 PAD.n8877 2.2505
R35459 PAD.n9049 PAD.n9048 2.2505
R35460 PAD.n9050 PAD.n8873 2.2505
R35461 PAD.n9052 PAD.n9051 2.2505
R35462 PAD.n9053 PAD.n8872 2.2505
R35463 PAD.n9058 PAD.n9057 2.2505
R35464 PAD.n9059 PAD.n8868 2.2505
R35465 PAD.n9061 PAD.n9060 2.2505
R35466 PAD.n9062 PAD.n8867 2.2505
R35467 PAD.n9067 PAD.n9066 2.2505
R35468 PAD.n9068 PAD.n8863 2.2505
R35469 PAD.n9070 PAD.n9069 2.2505
R35470 PAD.n9071 PAD.n8862 2.2505
R35471 PAD.n9076 PAD.n9075 2.2505
R35472 PAD.n9077 PAD.n8858 2.2505
R35473 PAD.n9079 PAD.n9078 2.2505
R35474 PAD.n9080 PAD.n8857 2.2505
R35475 PAD.n9085 PAD.n9084 2.2505
R35476 PAD.n9086 PAD.n8853 2.2505
R35477 PAD.n9088 PAD.n9087 2.2505
R35478 PAD.n9089 PAD.n8852 2.2505
R35479 PAD.n9094 PAD.n9093 2.2505
R35480 PAD.n9095 PAD.n8848 2.2505
R35481 PAD.n9097 PAD.n9096 2.2505
R35482 PAD.n9098 PAD.n8847 2.2505
R35483 PAD.n9103 PAD.n9102 2.2505
R35484 PAD.n9104 PAD.n8843 2.2505
R35485 PAD.n9106 PAD.n9105 2.2505
R35486 PAD.n9107 PAD.n8842 2.2505
R35487 PAD.n9112 PAD.n9111 2.2505
R35488 PAD.n9113 PAD.n8838 2.2505
R35489 PAD.n9115 PAD.n9114 2.2505
R35490 PAD.n9118 PAD.n8837 2.2505
R35491 PAD.n9120 PAD.n9119 2.2505
R35492 PAD.n8819 PAD.n8818 2.2505
R35493 PAD.n8529 PAD.n8528 2.2505
R35494 PAD.n8814 PAD.n8813 2.2505
R35495 PAD.n8811 PAD.n8810 2.2505
R35496 PAD.n8808 PAD.n8807 2.2505
R35497 PAD.n8800 PAD.n8531 2.2505
R35498 PAD.n8803 PAD.n8802 2.2505
R35499 PAD.n8799 PAD.n8798 2.2505
R35500 PAD.n8796 PAD.n8795 2.2505
R35501 PAD.n8788 PAD.n8533 2.2505
R35502 PAD.n8791 PAD.n8790 2.2505
R35503 PAD.n8787 PAD.n8786 2.2505
R35504 PAD.n8784 PAD.n8783 2.2505
R35505 PAD.n8776 PAD.n8535 2.2505
R35506 PAD.n8779 PAD.n8778 2.2505
R35507 PAD.n8775 PAD.n8774 2.2505
R35508 PAD.n8772 PAD.n8771 2.2505
R35509 PAD.n8764 PAD.n8537 2.2505
R35510 PAD.n8767 PAD.n8766 2.2505
R35511 PAD.n8763 PAD.n8762 2.2505
R35512 PAD.n8760 PAD.n8759 2.2505
R35513 PAD.n8752 PAD.n8539 2.2505
R35514 PAD.n8755 PAD.n8754 2.2505
R35515 PAD.n8751 PAD.n8750 2.2505
R35516 PAD.n8748 PAD.n8747 2.2505
R35517 PAD.n8740 PAD.n8541 2.2505
R35518 PAD.n8743 PAD.n8742 2.2505
R35519 PAD.n8739 PAD.n8738 2.2505
R35520 PAD.n8736 PAD.n8735 2.2505
R35521 PAD.n8728 PAD.n8543 2.2505
R35522 PAD.n8731 PAD.n8730 2.2505
R35523 PAD.n8727 PAD.n8726 2.2505
R35524 PAD.n8724 PAD.n8723 2.2505
R35525 PAD.n8716 PAD.n8545 2.2505
R35526 PAD.n8719 PAD.n8718 2.2505
R35527 PAD.n8715 PAD.n8714 2.2505
R35528 PAD.n8712 PAD.n8711 2.2505
R35529 PAD.n8704 PAD.n8547 2.2505
R35530 PAD.n8707 PAD.n8706 2.2505
R35531 PAD.n8703 PAD.n8702 2.2505
R35532 PAD.n8700 PAD.n8699 2.2505
R35533 PAD.n8692 PAD.n8549 2.2505
R35534 PAD.n8695 PAD.n8694 2.2505
R35535 PAD.n8691 PAD.n8690 2.2505
R35536 PAD.n8688 PAD.n8687 2.2505
R35537 PAD.n8680 PAD.n8551 2.2505
R35538 PAD.n8683 PAD.n8682 2.2505
R35539 PAD.n8679 PAD.n8678 2.2505
R35540 PAD.n8676 PAD.n8675 2.2505
R35541 PAD.n8668 PAD.n8553 2.2505
R35542 PAD.n8671 PAD.n8670 2.2505
R35543 PAD.n8667 PAD.n8666 2.2505
R35544 PAD.n8664 PAD.n8663 2.2505
R35545 PAD.n8656 PAD.n8555 2.2505
R35546 PAD.n8659 PAD.n8658 2.2505
R35547 PAD.n8655 PAD.n8654 2.2505
R35548 PAD.n8652 PAD.n8651 2.2505
R35549 PAD.n8644 PAD.n8557 2.2505
R35550 PAD.n8647 PAD.n8646 2.2505
R35551 PAD.n8643 PAD.n8642 2.2505
R35552 PAD.n8640 PAD.n8639 2.2505
R35553 PAD.n8632 PAD.n8559 2.2505
R35554 PAD.n8635 PAD.n8634 2.2505
R35555 PAD.n8631 PAD.n8630 2.2505
R35556 PAD.n8628 PAD.n8627 2.2505
R35557 PAD.n8620 PAD.n8561 2.2505
R35558 PAD.n8623 PAD.n8622 2.2505
R35559 PAD.n8619 PAD.n8618 2.2505
R35560 PAD.n8616 PAD.n8615 2.2505
R35561 PAD.n8608 PAD.n8563 2.2505
R35562 PAD.n8611 PAD.n8610 2.2505
R35563 PAD.n8607 PAD.n8606 2.2505
R35564 PAD.n8604 PAD.n8603 2.2505
R35565 PAD.n8596 PAD.n8565 2.2505
R35566 PAD.n8599 PAD.n8598 2.2505
R35567 PAD.n8595 PAD.n8594 2.2505
R35568 PAD.n8592 PAD.n8591 2.2505
R35569 PAD.n8584 PAD.n8567 2.2505
R35570 PAD.n8587 PAD.n8586 2.2505
R35571 PAD.n8583 PAD.n8582 2.2505
R35572 PAD.n8580 PAD.n8579 2.2505
R35573 PAD.n8572 PAD.n8569 2.2505
R35574 PAD.n8575 PAD.n8574 2.2505
R35575 PAD.n8571 PAD.n8570 2.2505
R35576 PAD.n8571 PAD.n2898 2.2505
R35577 PAD.n8576 PAD.n8575 2.2505
R35578 PAD.n8577 PAD.n8569 2.2505
R35579 PAD.n8579 PAD.n8578 2.2505
R35580 PAD.n8583 PAD.n8568 2.2505
R35581 PAD.n8588 PAD.n8587 2.2505
R35582 PAD.n8589 PAD.n8567 2.2505
R35583 PAD.n8591 PAD.n8590 2.2505
R35584 PAD.n8595 PAD.n8566 2.2505
R35585 PAD.n8600 PAD.n8599 2.2505
R35586 PAD.n8601 PAD.n8565 2.2505
R35587 PAD.n8603 PAD.n8602 2.2505
R35588 PAD.n8607 PAD.n8564 2.2505
R35589 PAD.n8612 PAD.n8611 2.2505
R35590 PAD.n8613 PAD.n8563 2.2505
R35591 PAD.n8615 PAD.n8614 2.2505
R35592 PAD.n8619 PAD.n8562 2.2505
R35593 PAD.n8624 PAD.n8623 2.2505
R35594 PAD.n8625 PAD.n8561 2.2505
R35595 PAD.n8627 PAD.n8626 2.2505
R35596 PAD.n8631 PAD.n8560 2.2505
R35597 PAD.n8636 PAD.n8635 2.2505
R35598 PAD.n8637 PAD.n8559 2.2505
R35599 PAD.n8639 PAD.n8638 2.2505
R35600 PAD.n8643 PAD.n8558 2.2505
R35601 PAD.n8648 PAD.n8647 2.2505
R35602 PAD.n8649 PAD.n8557 2.2505
R35603 PAD.n8651 PAD.n8650 2.2505
R35604 PAD.n8655 PAD.n8556 2.2505
R35605 PAD.n8660 PAD.n8659 2.2505
R35606 PAD.n8661 PAD.n8555 2.2505
R35607 PAD.n8663 PAD.n8662 2.2505
R35608 PAD.n8667 PAD.n8554 2.2505
R35609 PAD.n8672 PAD.n8671 2.2505
R35610 PAD.n8673 PAD.n8553 2.2505
R35611 PAD.n8675 PAD.n8674 2.2505
R35612 PAD.n8679 PAD.n8552 2.2505
R35613 PAD.n8684 PAD.n8683 2.2505
R35614 PAD.n8685 PAD.n8551 2.2505
R35615 PAD.n8687 PAD.n8686 2.2505
R35616 PAD.n8691 PAD.n8550 2.2505
R35617 PAD.n8696 PAD.n8695 2.2505
R35618 PAD.n8697 PAD.n8549 2.2505
R35619 PAD.n8699 PAD.n8698 2.2505
R35620 PAD.n8703 PAD.n8548 2.2505
R35621 PAD.n8708 PAD.n8707 2.2505
R35622 PAD.n8709 PAD.n8547 2.2505
R35623 PAD.n8711 PAD.n8710 2.2505
R35624 PAD.n8715 PAD.n8546 2.2505
R35625 PAD.n8720 PAD.n8719 2.2505
R35626 PAD.n8721 PAD.n8545 2.2505
R35627 PAD.n8723 PAD.n8722 2.2505
R35628 PAD.n8727 PAD.n8544 2.2505
R35629 PAD.n8732 PAD.n8731 2.2505
R35630 PAD.n8733 PAD.n8543 2.2505
R35631 PAD.n8735 PAD.n8734 2.2505
R35632 PAD.n8739 PAD.n8542 2.2505
R35633 PAD.n8744 PAD.n8743 2.2505
R35634 PAD.n8745 PAD.n8541 2.2505
R35635 PAD.n8747 PAD.n8746 2.2505
R35636 PAD.n8751 PAD.n8540 2.2505
R35637 PAD.n8756 PAD.n8755 2.2505
R35638 PAD.n8757 PAD.n8539 2.2505
R35639 PAD.n8759 PAD.n8758 2.2505
R35640 PAD.n8763 PAD.n8538 2.2505
R35641 PAD.n8768 PAD.n8767 2.2505
R35642 PAD.n8769 PAD.n8537 2.2505
R35643 PAD.n8771 PAD.n8770 2.2505
R35644 PAD.n8775 PAD.n8536 2.2505
R35645 PAD.n8780 PAD.n8779 2.2505
R35646 PAD.n8781 PAD.n8535 2.2505
R35647 PAD.n8783 PAD.n8782 2.2505
R35648 PAD.n8787 PAD.n8534 2.2505
R35649 PAD.n8792 PAD.n8791 2.2505
R35650 PAD.n8793 PAD.n8533 2.2505
R35651 PAD.n8795 PAD.n8794 2.2505
R35652 PAD.n8799 PAD.n8532 2.2505
R35653 PAD.n8804 PAD.n8803 2.2505
R35654 PAD.n8805 PAD.n8531 2.2505
R35655 PAD.n8807 PAD.n8806 2.2505
R35656 PAD.n8811 PAD.n8530 2.2505
R35657 PAD.n8815 PAD.n8814 2.2505
R35658 PAD.n8816 PAD.n8529 2.2505
R35659 PAD.n8818 PAD.n8817 2.2505
R35660 PAD.n3041 PAD.n2994 2.2505
R35661 PAD.n3040 PAD.n3039 2.2505
R35662 PAD.n3046 PAD.n3045 2.2505
R35663 PAD.n3049 PAD.n3048 2.2505
R35664 PAD.n3053 PAD.n3052 2.2505
R35665 PAD.n3050 PAD.n3036 2.2505
R35666 PAD.n3058 PAD.n3057 2.2505
R35667 PAD.n3061 PAD.n3060 2.2505
R35668 PAD.n3065 PAD.n3064 2.2505
R35669 PAD.n3062 PAD.n3034 2.2505
R35670 PAD.n3070 PAD.n3069 2.2505
R35671 PAD.n3073 PAD.n3072 2.2505
R35672 PAD.n3077 PAD.n3076 2.2505
R35673 PAD.n3074 PAD.n3032 2.2505
R35674 PAD.n3082 PAD.n3081 2.2505
R35675 PAD.n3085 PAD.n3084 2.2505
R35676 PAD.n3089 PAD.n3088 2.2505
R35677 PAD.n3086 PAD.n3030 2.2505
R35678 PAD.n3094 PAD.n3093 2.2505
R35679 PAD.n3097 PAD.n3096 2.2505
R35680 PAD.n3101 PAD.n3100 2.2505
R35681 PAD.n3098 PAD.n3028 2.2505
R35682 PAD.n3106 PAD.n3105 2.2505
R35683 PAD.n3109 PAD.n3108 2.2505
R35684 PAD.n3113 PAD.n3112 2.2505
R35685 PAD.n3110 PAD.n3026 2.2505
R35686 PAD.n3118 PAD.n3117 2.2505
R35687 PAD.n3121 PAD.n3120 2.2505
R35688 PAD.n3125 PAD.n3124 2.2505
R35689 PAD.n3122 PAD.n3024 2.2505
R35690 PAD.n3130 PAD.n3129 2.2505
R35691 PAD.n3133 PAD.n3132 2.2505
R35692 PAD.n3137 PAD.n3136 2.2505
R35693 PAD.n3134 PAD.n3022 2.2505
R35694 PAD.n3142 PAD.n3141 2.2505
R35695 PAD.n3145 PAD.n3144 2.2505
R35696 PAD.n3149 PAD.n3148 2.2505
R35697 PAD.n3146 PAD.n3020 2.2505
R35698 PAD.n3154 PAD.n3153 2.2505
R35699 PAD.n3157 PAD.n3156 2.2505
R35700 PAD.n3161 PAD.n3160 2.2505
R35701 PAD.n3158 PAD.n3018 2.2505
R35702 PAD.n3166 PAD.n3165 2.2505
R35703 PAD.n3169 PAD.n3168 2.2505
R35704 PAD.n3173 PAD.n3172 2.2505
R35705 PAD.n3170 PAD.n3016 2.2505
R35706 PAD.n3178 PAD.n3177 2.2505
R35707 PAD.n3181 PAD.n3180 2.2505
R35708 PAD.n3185 PAD.n3184 2.2505
R35709 PAD.n3182 PAD.n3014 2.2505
R35710 PAD.n3190 PAD.n3189 2.2505
R35711 PAD.n3193 PAD.n3192 2.2505
R35712 PAD.n3197 PAD.n3196 2.2505
R35713 PAD.n3194 PAD.n3012 2.2505
R35714 PAD.n3202 PAD.n3201 2.2505
R35715 PAD.n3205 PAD.n3204 2.2505
R35716 PAD.n3209 PAD.n3208 2.2505
R35717 PAD.n3206 PAD.n3010 2.2505
R35718 PAD.n3214 PAD.n3213 2.2505
R35719 PAD.n3217 PAD.n3216 2.2505
R35720 PAD.n3221 PAD.n3220 2.2505
R35721 PAD.n3218 PAD.n3008 2.2505
R35722 PAD.n3226 PAD.n3225 2.2505
R35723 PAD.n3229 PAD.n3228 2.2505
R35724 PAD.n3233 PAD.n3232 2.2505
R35725 PAD.n3230 PAD.n3006 2.2505
R35726 PAD.n3238 PAD.n3237 2.2505
R35727 PAD.n3241 PAD.n3240 2.2505
R35728 PAD.n3245 PAD.n3244 2.2505
R35729 PAD.n3242 PAD.n3004 2.2505
R35730 PAD.n3250 PAD.n3249 2.2505
R35731 PAD.n3253 PAD.n3252 2.2505
R35732 PAD.n3257 PAD.n3256 2.2505
R35733 PAD.n3254 PAD.n3002 2.2505
R35734 PAD.n3262 PAD.n3261 2.2505
R35735 PAD.n3265 PAD.n3264 2.2505
R35736 PAD.n3269 PAD.n3268 2.2505
R35737 PAD.n3266 PAD.n3000 2.2505
R35738 PAD.n3274 PAD.n3273 2.2505
R35739 PAD.n3277 PAD.n3276 2.2505
R35740 PAD.n3281 PAD.n3280 2.2505
R35741 PAD.n3278 PAD.n2998 2.2505
R35742 PAD.n8514 PAD.n8513 2.2505
R35743 PAD.n8516 PAD.n2995 2.2505
R35744 PAD.n8511 PAD.n2995 2.2505
R35745 PAD.n8513 PAD.n8512 2.2505
R35746 PAD.n3283 PAD.n2998 2.2505
R35747 PAD.n3282 PAD.n3281 2.2505
R35748 PAD.n3277 PAD.n2999 2.2505
R35749 PAD.n3273 PAD.n3272 2.2505
R35750 PAD.n3271 PAD.n3000 2.2505
R35751 PAD.n3270 PAD.n3269 2.2505
R35752 PAD.n3265 PAD.n3001 2.2505
R35753 PAD.n3261 PAD.n3260 2.2505
R35754 PAD.n3259 PAD.n3002 2.2505
R35755 PAD.n3258 PAD.n3257 2.2505
R35756 PAD.n3253 PAD.n3003 2.2505
R35757 PAD.n3249 PAD.n3248 2.2505
R35758 PAD.n3247 PAD.n3004 2.2505
R35759 PAD.n3246 PAD.n3245 2.2505
R35760 PAD.n3241 PAD.n3005 2.2505
R35761 PAD.n3237 PAD.n3236 2.2505
R35762 PAD.n3235 PAD.n3006 2.2505
R35763 PAD.n3234 PAD.n3233 2.2505
R35764 PAD.n3229 PAD.n3007 2.2505
R35765 PAD.n3225 PAD.n3224 2.2505
R35766 PAD.n3223 PAD.n3008 2.2505
R35767 PAD.n3222 PAD.n3221 2.2505
R35768 PAD.n3217 PAD.n3009 2.2505
R35769 PAD.n3213 PAD.n3212 2.2505
R35770 PAD.n3211 PAD.n3010 2.2505
R35771 PAD.n3210 PAD.n3209 2.2505
R35772 PAD.n3205 PAD.n3011 2.2505
R35773 PAD.n3201 PAD.n3200 2.2505
R35774 PAD.n3199 PAD.n3012 2.2505
R35775 PAD.n3198 PAD.n3197 2.2505
R35776 PAD.n3193 PAD.n3013 2.2505
R35777 PAD.n3189 PAD.n3188 2.2505
R35778 PAD.n3187 PAD.n3014 2.2505
R35779 PAD.n3186 PAD.n3185 2.2505
R35780 PAD.n3181 PAD.n3015 2.2505
R35781 PAD.n3177 PAD.n3176 2.2505
R35782 PAD.n3175 PAD.n3016 2.2505
R35783 PAD.n3174 PAD.n3173 2.2505
R35784 PAD.n3169 PAD.n3017 2.2505
R35785 PAD.n3165 PAD.n3164 2.2505
R35786 PAD.n3163 PAD.n3018 2.2505
R35787 PAD.n3162 PAD.n3161 2.2505
R35788 PAD.n3157 PAD.n3019 2.2505
R35789 PAD.n3153 PAD.n3152 2.2505
R35790 PAD.n3151 PAD.n3020 2.2505
R35791 PAD.n3150 PAD.n3149 2.2505
R35792 PAD.n3145 PAD.n3021 2.2505
R35793 PAD.n3141 PAD.n3140 2.2505
R35794 PAD.n3139 PAD.n3022 2.2505
R35795 PAD.n3138 PAD.n3137 2.2505
R35796 PAD.n3133 PAD.n3023 2.2505
R35797 PAD.n3129 PAD.n3128 2.2505
R35798 PAD.n3127 PAD.n3024 2.2505
R35799 PAD.n3126 PAD.n3125 2.2505
R35800 PAD.n3121 PAD.n3025 2.2505
R35801 PAD.n3117 PAD.n3116 2.2505
R35802 PAD.n3115 PAD.n3026 2.2505
R35803 PAD.n3114 PAD.n3113 2.2505
R35804 PAD.n3109 PAD.n3027 2.2505
R35805 PAD.n3105 PAD.n3104 2.2505
R35806 PAD.n3103 PAD.n3028 2.2505
R35807 PAD.n3102 PAD.n3101 2.2505
R35808 PAD.n3097 PAD.n3029 2.2505
R35809 PAD.n3093 PAD.n3092 2.2505
R35810 PAD.n3091 PAD.n3030 2.2505
R35811 PAD.n3090 PAD.n3089 2.2505
R35812 PAD.n3085 PAD.n3031 2.2505
R35813 PAD.n3081 PAD.n3080 2.2505
R35814 PAD.n3079 PAD.n3032 2.2505
R35815 PAD.n3078 PAD.n3077 2.2505
R35816 PAD.n3073 PAD.n3033 2.2505
R35817 PAD.n3069 PAD.n3068 2.2505
R35818 PAD.n3067 PAD.n3034 2.2505
R35819 PAD.n3066 PAD.n3065 2.2505
R35820 PAD.n3061 PAD.n3035 2.2505
R35821 PAD.n3057 PAD.n3056 2.2505
R35822 PAD.n3055 PAD.n3036 2.2505
R35823 PAD.n3054 PAD.n3053 2.2505
R35824 PAD.n3049 PAD.n3037 2.2505
R35825 PAD.n3045 PAD.n3044 2.2505
R35826 PAD.n3043 PAD.n3040 2.2505
R35827 PAD.n3042 PAD.n3041 2.2505
R35828 PAD.n3386 PAD.n3338 2.2505
R35829 PAD.n3385 PAD.n3384 2.2505
R35830 PAD.n3391 PAD.n3390 2.2505
R35831 PAD.n3394 PAD.n3393 2.2505
R35832 PAD.n3398 PAD.n3397 2.2505
R35833 PAD.n3395 PAD.n3381 2.2505
R35834 PAD.n3403 PAD.n3402 2.2505
R35835 PAD.n3406 PAD.n3405 2.2505
R35836 PAD.n3410 PAD.n3409 2.2505
R35837 PAD.n3407 PAD.n3379 2.2505
R35838 PAD.n3415 PAD.n3414 2.2505
R35839 PAD.n3418 PAD.n3417 2.2505
R35840 PAD.n3422 PAD.n3421 2.2505
R35841 PAD.n3419 PAD.n3377 2.2505
R35842 PAD.n3427 PAD.n3426 2.2505
R35843 PAD.n3430 PAD.n3429 2.2505
R35844 PAD.n3434 PAD.n3433 2.2505
R35845 PAD.n3431 PAD.n3375 2.2505
R35846 PAD.n3439 PAD.n3438 2.2505
R35847 PAD.n3442 PAD.n3441 2.2505
R35848 PAD.n3446 PAD.n3445 2.2505
R35849 PAD.n3443 PAD.n3373 2.2505
R35850 PAD.n3451 PAD.n3450 2.2505
R35851 PAD.n3454 PAD.n3453 2.2505
R35852 PAD.n3458 PAD.n3457 2.2505
R35853 PAD.n3455 PAD.n3371 2.2505
R35854 PAD.n3463 PAD.n3462 2.2505
R35855 PAD.n3466 PAD.n3465 2.2505
R35856 PAD.n3470 PAD.n3469 2.2505
R35857 PAD.n3467 PAD.n3369 2.2505
R35858 PAD.n3475 PAD.n3474 2.2505
R35859 PAD.n3478 PAD.n3477 2.2505
R35860 PAD.n3482 PAD.n3481 2.2505
R35861 PAD.n3479 PAD.n3367 2.2505
R35862 PAD.n3487 PAD.n3486 2.2505
R35863 PAD.n3490 PAD.n3489 2.2505
R35864 PAD.n3494 PAD.n3493 2.2505
R35865 PAD.n3491 PAD.n3365 2.2505
R35866 PAD.n3499 PAD.n3498 2.2505
R35867 PAD.n3502 PAD.n3501 2.2505
R35868 PAD.n3506 PAD.n3505 2.2505
R35869 PAD.n3503 PAD.n3363 2.2505
R35870 PAD.n3511 PAD.n3510 2.2505
R35871 PAD.n3514 PAD.n3513 2.2505
R35872 PAD.n3518 PAD.n3517 2.2505
R35873 PAD.n3515 PAD.n3361 2.2505
R35874 PAD.n3523 PAD.n3522 2.2505
R35875 PAD.n3526 PAD.n3525 2.2505
R35876 PAD.n3530 PAD.n3529 2.2505
R35877 PAD.n3527 PAD.n3359 2.2505
R35878 PAD.n3535 PAD.n3534 2.2505
R35879 PAD.n3538 PAD.n3537 2.2505
R35880 PAD.n3542 PAD.n3541 2.2505
R35881 PAD.n3539 PAD.n3357 2.2505
R35882 PAD.n3547 PAD.n3546 2.2505
R35883 PAD.n3550 PAD.n3549 2.2505
R35884 PAD.n3554 PAD.n3553 2.2505
R35885 PAD.n3551 PAD.n3355 2.2505
R35886 PAD.n3559 PAD.n3558 2.2505
R35887 PAD.n3562 PAD.n3561 2.2505
R35888 PAD.n3566 PAD.n3565 2.2505
R35889 PAD.n3563 PAD.n3353 2.2505
R35890 PAD.n3571 PAD.n3570 2.2505
R35891 PAD.n3574 PAD.n3573 2.2505
R35892 PAD.n3578 PAD.n3577 2.2505
R35893 PAD.n3575 PAD.n3351 2.2505
R35894 PAD.n3583 PAD.n3582 2.2505
R35895 PAD.n3586 PAD.n3585 2.2505
R35896 PAD.n3590 PAD.n3589 2.2505
R35897 PAD.n3587 PAD.n3349 2.2505
R35898 PAD.n3595 PAD.n3594 2.2505
R35899 PAD.n3598 PAD.n3597 2.2505
R35900 PAD.n3602 PAD.n3601 2.2505
R35901 PAD.n3599 PAD.n3347 2.2505
R35902 PAD.n3607 PAD.n3606 2.2505
R35903 PAD.n3610 PAD.n3609 2.2505
R35904 PAD.n3614 PAD.n3613 2.2505
R35905 PAD.n3611 PAD.n3345 2.2505
R35906 PAD.n3619 PAD.n3618 2.2505
R35907 PAD.n3622 PAD.n3621 2.2505
R35908 PAD.n3626 PAD.n3625 2.2505
R35909 PAD.n3623 PAD.n3343 2.2505
R35910 PAD.n8489 PAD.n8488 2.2505
R35911 PAD.n8491 PAD.n3340 2.2505
R35912 PAD.n8486 PAD.n3340 2.2505
R35913 PAD.n8488 PAD.n8487 2.2505
R35914 PAD.n3628 PAD.n3343 2.2505
R35915 PAD.n3627 PAD.n3626 2.2505
R35916 PAD.n3622 PAD.n3344 2.2505
R35917 PAD.n3618 PAD.n3617 2.2505
R35918 PAD.n3616 PAD.n3345 2.2505
R35919 PAD.n3615 PAD.n3614 2.2505
R35920 PAD.n3610 PAD.n3346 2.2505
R35921 PAD.n3606 PAD.n3605 2.2505
R35922 PAD.n3604 PAD.n3347 2.2505
R35923 PAD.n3603 PAD.n3602 2.2505
R35924 PAD.n3598 PAD.n3348 2.2505
R35925 PAD.n3594 PAD.n3593 2.2505
R35926 PAD.n3592 PAD.n3349 2.2505
R35927 PAD.n3591 PAD.n3590 2.2505
R35928 PAD.n3586 PAD.n3350 2.2505
R35929 PAD.n3582 PAD.n3581 2.2505
R35930 PAD.n3580 PAD.n3351 2.2505
R35931 PAD.n3579 PAD.n3578 2.2505
R35932 PAD.n3574 PAD.n3352 2.2505
R35933 PAD.n3570 PAD.n3569 2.2505
R35934 PAD.n3568 PAD.n3353 2.2505
R35935 PAD.n3567 PAD.n3566 2.2505
R35936 PAD.n3562 PAD.n3354 2.2505
R35937 PAD.n3558 PAD.n3557 2.2505
R35938 PAD.n3556 PAD.n3355 2.2505
R35939 PAD.n3555 PAD.n3554 2.2505
R35940 PAD.n3550 PAD.n3356 2.2505
R35941 PAD.n3546 PAD.n3545 2.2505
R35942 PAD.n3544 PAD.n3357 2.2505
R35943 PAD.n3543 PAD.n3542 2.2505
R35944 PAD.n3538 PAD.n3358 2.2505
R35945 PAD.n3534 PAD.n3533 2.2505
R35946 PAD.n3532 PAD.n3359 2.2505
R35947 PAD.n3531 PAD.n3530 2.2505
R35948 PAD.n3526 PAD.n3360 2.2505
R35949 PAD.n3522 PAD.n3521 2.2505
R35950 PAD.n3520 PAD.n3361 2.2505
R35951 PAD.n3519 PAD.n3518 2.2505
R35952 PAD.n3514 PAD.n3362 2.2505
R35953 PAD.n3510 PAD.n3509 2.2505
R35954 PAD.n3508 PAD.n3363 2.2505
R35955 PAD.n3507 PAD.n3506 2.2505
R35956 PAD.n3502 PAD.n3364 2.2505
R35957 PAD.n3498 PAD.n3497 2.2505
R35958 PAD.n3496 PAD.n3365 2.2505
R35959 PAD.n3495 PAD.n3494 2.2505
R35960 PAD.n3490 PAD.n3366 2.2505
R35961 PAD.n3486 PAD.n3485 2.2505
R35962 PAD.n3484 PAD.n3367 2.2505
R35963 PAD.n3483 PAD.n3482 2.2505
R35964 PAD.n3478 PAD.n3368 2.2505
R35965 PAD.n3474 PAD.n3473 2.2505
R35966 PAD.n3472 PAD.n3369 2.2505
R35967 PAD.n3471 PAD.n3470 2.2505
R35968 PAD.n3466 PAD.n3370 2.2505
R35969 PAD.n3462 PAD.n3461 2.2505
R35970 PAD.n3460 PAD.n3371 2.2505
R35971 PAD.n3459 PAD.n3458 2.2505
R35972 PAD.n3454 PAD.n3372 2.2505
R35973 PAD.n3450 PAD.n3449 2.2505
R35974 PAD.n3448 PAD.n3373 2.2505
R35975 PAD.n3447 PAD.n3446 2.2505
R35976 PAD.n3442 PAD.n3374 2.2505
R35977 PAD.n3438 PAD.n3437 2.2505
R35978 PAD.n3436 PAD.n3375 2.2505
R35979 PAD.n3435 PAD.n3434 2.2505
R35980 PAD.n3430 PAD.n3376 2.2505
R35981 PAD.n3426 PAD.n3425 2.2505
R35982 PAD.n3424 PAD.n3377 2.2505
R35983 PAD.n3423 PAD.n3422 2.2505
R35984 PAD.n3418 PAD.n3378 2.2505
R35985 PAD.n3414 PAD.n3413 2.2505
R35986 PAD.n3412 PAD.n3379 2.2505
R35987 PAD.n3411 PAD.n3410 2.2505
R35988 PAD.n3406 PAD.n3380 2.2505
R35989 PAD.n3402 PAD.n3401 2.2505
R35990 PAD.n3400 PAD.n3381 2.2505
R35991 PAD.n3399 PAD.n3398 2.2505
R35992 PAD.n3394 PAD.n3382 2.2505
R35993 PAD.n3390 PAD.n3389 2.2505
R35994 PAD.n3388 PAD.n3385 2.2505
R35995 PAD.n3387 PAD.n3386 2.2505
R35996 PAD.n3731 PAD.n3683 2.2505
R35997 PAD.n3730 PAD.n3729 2.2505
R35998 PAD.n3736 PAD.n3735 2.2505
R35999 PAD.n3739 PAD.n3738 2.2505
R36000 PAD.n3743 PAD.n3742 2.2505
R36001 PAD.n3740 PAD.n3726 2.2505
R36002 PAD.n3748 PAD.n3747 2.2505
R36003 PAD.n3751 PAD.n3750 2.2505
R36004 PAD.n3755 PAD.n3754 2.2505
R36005 PAD.n3752 PAD.n3724 2.2505
R36006 PAD.n3760 PAD.n3759 2.2505
R36007 PAD.n3763 PAD.n3762 2.2505
R36008 PAD.n3767 PAD.n3766 2.2505
R36009 PAD.n3764 PAD.n3722 2.2505
R36010 PAD.n3772 PAD.n3771 2.2505
R36011 PAD.n3775 PAD.n3774 2.2505
R36012 PAD.n3779 PAD.n3778 2.2505
R36013 PAD.n3776 PAD.n3720 2.2505
R36014 PAD.n3784 PAD.n3783 2.2505
R36015 PAD.n3787 PAD.n3786 2.2505
R36016 PAD.n3791 PAD.n3790 2.2505
R36017 PAD.n3788 PAD.n3718 2.2505
R36018 PAD.n3796 PAD.n3795 2.2505
R36019 PAD.n3799 PAD.n3798 2.2505
R36020 PAD.n3803 PAD.n3802 2.2505
R36021 PAD.n3800 PAD.n3716 2.2505
R36022 PAD.n3808 PAD.n3807 2.2505
R36023 PAD.n3811 PAD.n3810 2.2505
R36024 PAD.n3815 PAD.n3814 2.2505
R36025 PAD.n3812 PAD.n3714 2.2505
R36026 PAD.n3820 PAD.n3819 2.2505
R36027 PAD.n3823 PAD.n3822 2.2505
R36028 PAD.n3827 PAD.n3826 2.2505
R36029 PAD.n3824 PAD.n3712 2.2505
R36030 PAD.n3832 PAD.n3831 2.2505
R36031 PAD.n3835 PAD.n3834 2.2505
R36032 PAD.n3839 PAD.n3838 2.2505
R36033 PAD.n3836 PAD.n3710 2.2505
R36034 PAD.n3844 PAD.n3843 2.2505
R36035 PAD.n3847 PAD.n3846 2.2505
R36036 PAD.n3851 PAD.n3850 2.2505
R36037 PAD.n3848 PAD.n3708 2.2505
R36038 PAD.n3856 PAD.n3855 2.2505
R36039 PAD.n3859 PAD.n3858 2.2505
R36040 PAD.n3863 PAD.n3862 2.2505
R36041 PAD.n3860 PAD.n3706 2.2505
R36042 PAD.n3868 PAD.n3867 2.2505
R36043 PAD.n3871 PAD.n3870 2.2505
R36044 PAD.n3875 PAD.n3874 2.2505
R36045 PAD.n3872 PAD.n3704 2.2505
R36046 PAD.n3880 PAD.n3879 2.2505
R36047 PAD.n3883 PAD.n3882 2.2505
R36048 PAD.n3887 PAD.n3886 2.2505
R36049 PAD.n3884 PAD.n3702 2.2505
R36050 PAD.n3892 PAD.n3891 2.2505
R36051 PAD.n3895 PAD.n3894 2.2505
R36052 PAD.n3899 PAD.n3898 2.2505
R36053 PAD.n3896 PAD.n3700 2.2505
R36054 PAD.n3904 PAD.n3903 2.2505
R36055 PAD.n3907 PAD.n3906 2.2505
R36056 PAD.n3911 PAD.n3910 2.2505
R36057 PAD.n3908 PAD.n3698 2.2505
R36058 PAD.n3916 PAD.n3915 2.2505
R36059 PAD.n3919 PAD.n3918 2.2505
R36060 PAD.n3923 PAD.n3922 2.2505
R36061 PAD.n3920 PAD.n3696 2.2505
R36062 PAD.n3928 PAD.n3927 2.2505
R36063 PAD.n3931 PAD.n3930 2.2505
R36064 PAD.n3935 PAD.n3934 2.2505
R36065 PAD.n3932 PAD.n3694 2.2505
R36066 PAD.n3940 PAD.n3939 2.2505
R36067 PAD.n3943 PAD.n3942 2.2505
R36068 PAD.n3947 PAD.n3946 2.2505
R36069 PAD.n3944 PAD.n3692 2.2505
R36070 PAD.n3952 PAD.n3951 2.2505
R36071 PAD.n3955 PAD.n3954 2.2505
R36072 PAD.n3959 PAD.n3958 2.2505
R36073 PAD.n3956 PAD.n3690 2.2505
R36074 PAD.n3964 PAD.n3963 2.2505
R36075 PAD.n3967 PAD.n3966 2.2505
R36076 PAD.n3971 PAD.n3970 2.2505
R36077 PAD.n3968 PAD.n3688 2.2505
R36078 PAD.n8465 PAD.n8464 2.2505
R36079 PAD.n8467 PAD.n3685 2.2505
R36080 PAD.n8462 PAD.n3685 2.2505
R36081 PAD.n8464 PAD.n8463 2.2505
R36082 PAD.n3973 PAD.n3688 2.2505
R36083 PAD.n3972 PAD.n3971 2.2505
R36084 PAD.n3967 PAD.n3689 2.2505
R36085 PAD.n3963 PAD.n3962 2.2505
R36086 PAD.n3961 PAD.n3690 2.2505
R36087 PAD.n3960 PAD.n3959 2.2505
R36088 PAD.n3955 PAD.n3691 2.2505
R36089 PAD.n3951 PAD.n3950 2.2505
R36090 PAD.n3949 PAD.n3692 2.2505
R36091 PAD.n3948 PAD.n3947 2.2505
R36092 PAD.n3943 PAD.n3693 2.2505
R36093 PAD.n3939 PAD.n3938 2.2505
R36094 PAD.n3937 PAD.n3694 2.2505
R36095 PAD.n3936 PAD.n3935 2.2505
R36096 PAD.n3931 PAD.n3695 2.2505
R36097 PAD.n3927 PAD.n3926 2.2505
R36098 PAD.n3925 PAD.n3696 2.2505
R36099 PAD.n3924 PAD.n3923 2.2505
R36100 PAD.n3919 PAD.n3697 2.2505
R36101 PAD.n3915 PAD.n3914 2.2505
R36102 PAD.n3913 PAD.n3698 2.2505
R36103 PAD.n3912 PAD.n3911 2.2505
R36104 PAD.n3907 PAD.n3699 2.2505
R36105 PAD.n3903 PAD.n3902 2.2505
R36106 PAD.n3901 PAD.n3700 2.2505
R36107 PAD.n3900 PAD.n3899 2.2505
R36108 PAD.n3895 PAD.n3701 2.2505
R36109 PAD.n3891 PAD.n3890 2.2505
R36110 PAD.n3889 PAD.n3702 2.2505
R36111 PAD.n3888 PAD.n3887 2.2505
R36112 PAD.n3883 PAD.n3703 2.2505
R36113 PAD.n3879 PAD.n3878 2.2505
R36114 PAD.n3877 PAD.n3704 2.2505
R36115 PAD.n3876 PAD.n3875 2.2505
R36116 PAD.n3871 PAD.n3705 2.2505
R36117 PAD.n3867 PAD.n3866 2.2505
R36118 PAD.n3865 PAD.n3706 2.2505
R36119 PAD.n3864 PAD.n3863 2.2505
R36120 PAD.n3859 PAD.n3707 2.2505
R36121 PAD.n3855 PAD.n3854 2.2505
R36122 PAD.n3853 PAD.n3708 2.2505
R36123 PAD.n3852 PAD.n3851 2.2505
R36124 PAD.n3847 PAD.n3709 2.2505
R36125 PAD.n3843 PAD.n3842 2.2505
R36126 PAD.n3841 PAD.n3710 2.2505
R36127 PAD.n3840 PAD.n3839 2.2505
R36128 PAD.n3835 PAD.n3711 2.2505
R36129 PAD.n3831 PAD.n3830 2.2505
R36130 PAD.n3829 PAD.n3712 2.2505
R36131 PAD.n3828 PAD.n3827 2.2505
R36132 PAD.n3823 PAD.n3713 2.2505
R36133 PAD.n3819 PAD.n3818 2.2505
R36134 PAD.n3817 PAD.n3714 2.2505
R36135 PAD.n3816 PAD.n3815 2.2505
R36136 PAD.n3811 PAD.n3715 2.2505
R36137 PAD.n3807 PAD.n3806 2.2505
R36138 PAD.n3805 PAD.n3716 2.2505
R36139 PAD.n3804 PAD.n3803 2.2505
R36140 PAD.n3799 PAD.n3717 2.2505
R36141 PAD.n3795 PAD.n3794 2.2505
R36142 PAD.n3793 PAD.n3718 2.2505
R36143 PAD.n3792 PAD.n3791 2.2505
R36144 PAD.n3787 PAD.n3719 2.2505
R36145 PAD.n3783 PAD.n3782 2.2505
R36146 PAD.n3781 PAD.n3720 2.2505
R36147 PAD.n3780 PAD.n3779 2.2505
R36148 PAD.n3775 PAD.n3721 2.2505
R36149 PAD.n3771 PAD.n3770 2.2505
R36150 PAD.n3769 PAD.n3722 2.2505
R36151 PAD.n3768 PAD.n3767 2.2505
R36152 PAD.n3763 PAD.n3723 2.2505
R36153 PAD.n3759 PAD.n3758 2.2505
R36154 PAD.n3757 PAD.n3724 2.2505
R36155 PAD.n3756 PAD.n3755 2.2505
R36156 PAD.n3751 PAD.n3725 2.2505
R36157 PAD.n3747 PAD.n3746 2.2505
R36158 PAD.n3745 PAD.n3726 2.2505
R36159 PAD.n3744 PAD.n3743 2.2505
R36160 PAD.n3739 PAD.n3727 2.2505
R36161 PAD.n3735 PAD.n3734 2.2505
R36162 PAD.n3733 PAD.n3730 2.2505
R36163 PAD.n3732 PAD.n3731 2.2505
R36164 PAD.n4072 PAD.n4025 2.2505
R36165 PAD.n4071 PAD.n4070 2.2505
R36166 PAD.n4077 PAD.n4076 2.2505
R36167 PAD.n4080 PAD.n4079 2.2505
R36168 PAD.n4084 PAD.n4083 2.2505
R36169 PAD.n4081 PAD.n4067 2.2505
R36170 PAD.n4089 PAD.n4088 2.2505
R36171 PAD.n4092 PAD.n4091 2.2505
R36172 PAD.n4096 PAD.n4095 2.2505
R36173 PAD.n4093 PAD.n4065 2.2505
R36174 PAD.n4101 PAD.n4100 2.2505
R36175 PAD.n4104 PAD.n4103 2.2505
R36176 PAD.n4108 PAD.n4107 2.2505
R36177 PAD.n4105 PAD.n4063 2.2505
R36178 PAD.n4113 PAD.n4112 2.2505
R36179 PAD.n4116 PAD.n4115 2.2505
R36180 PAD.n4120 PAD.n4119 2.2505
R36181 PAD.n4117 PAD.n4061 2.2505
R36182 PAD.n4125 PAD.n4124 2.2505
R36183 PAD.n4128 PAD.n4127 2.2505
R36184 PAD.n4132 PAD.n4131 2.2505
R36185 PAD.n4129 PAD.n4059 2.2505
R36186 PAD.n4137 PAD.n4136 2.2505
R36187 PAD.n4140 PAD.n4139 2.2505
R36188 PAD.n4144 PAD.n4143 2.2505
R36189 PAD.n4141 PAD.n4057 2.2505
R36190 PAD.n4149 PAD.n4148 2.2505
R36191 PAD.n4152 PAD.n4151 2.2505
R36192 PAD.n4156 PAD.n4155 2.2505
R36193 PAD.n4153 PAD.n4055 2.2505
R36194 PAD.n4161 PAD.n4160 2.2505
R36195 PAD.n4164 PAD.n4163 2.2505
R36196 PAD.n4168 PAD.n4167 2.2505
R36197 PAD.n4165 PAD.n4053 2.2505
R36198 PAD.n4173 PAD.n4172 2.2505
R36199 PAD.n4176 PAD.n4175 2.2505
R36200 PAD.n4180 PAD.n4179 2.2505
R36201 PAD.n4177 PAD.n4051 2.2505
R36202 PAD.n4185 PAD.n4184 2.2505
R36203 PAD.n4188 PAD.n4187 2.2505
R36204 PAD.n4192 PAD.n4191 2.2505
R36205 PAD.n4189 PAD.n4049 2.2505
R36206 PAD.n4197 PAD.n4196 2.2505
R36207 PAD.n4200 PAD.n4199 2.2505
R36208 PAD.n4204 PAD.n4203 2.2505
R36209 PAD.n4201 PAD.n4047 2.2505
R36210 PAD.n4209 PAD.n4208 2.2505
R36211 PAD.n4212 PAD.n4211 2.2505
R36212 PAD.n4216 PAD.n4215 2.2505
R36213 PAD.n4213 PAD.n4045 2.2505
R36214 PAD.n4221 PAD.n4220 2.2505
R36215 PAD.n4224 PAD.n4223 2.2505
R36216 PAD.n4228 PAD.n4227 2.2505
R36217 PAD.n4225 PAD.n4043 2.2505
R36218 PAD.n4233 PAD.n4232 2.2505
R36219 PAD.n4236 PAD.n4235 2.2505
R36220 PAD.n4240 PAD.n4239 2.2505
R36221 PAD.n4237 PAD.n4041 2.2505
R36222 PAD.n4245 PAD.n4244 2.2505
R36223 PAD.n4248 PAD.n4247 2.2505
R36224 PAD.n4252 PAD.n4251 2.2505
R36225 PAD.n4249 PAD.n4039 2.2505
R36226 PAD.n4257 PAD.n4256 2.2505
R36227 PAD.n4260 PAD.n4259 2.2505
R36228 PAD.n4264 PAD.n4263 2.2505
R36229 PAD.n4261 PAD.n4037 2.2505
R36230 PAD.n4269 PAD.n4268 2.2505
R36231 PAD.n4272 PAD.n4271 2.2505
R36232 PAD.n4276 PAD.n4275 2.2505
R36233 PAD.n4273 PAD.n4035 2.2505
R36234 PAD.n4281 PAD.n4280 2.2505
R36235 PAD.n4284 PAD.n4283 2.2505
R36236 PAD.n4288 PAD.n4287 2.2505
R36237 PAD.n4285 PAD.n4033 2.2505
R36238 PAD.n4293 PAD.n4292 2.2505
R36239 PAD.n4296 PAD.n4295 2.2505
R36240 PAD.n4300 PAD.n4299 2.2505
R36241 PAD.n4297 PAD.n4031 2.2505
R36242 PAD.n4305 PAD.n4304 2.2505
R36243 PAD.n4308 PAD.n4307 2.2505
R36244 PAD.n4312 PAD.n4311 2.2505
R36245 PAD.n4309 PAD.n4029 2.2505
R36246 PAD.n8441 PAD.n8440 2.2505
R36247 PAD.n8443 PAD.n4026 2.2505
R36248 PAD.n8438 PAD.n4026 2.2505
R36249 PAD.n8440 PAD.n8439 2.2505
R36250 PAD.n4314 PAD.n4029 2.2505
R36251 PAD.n4313 PAD.n4312 2.2505
R36252 PAD.n4308 PAD.n4030 2.2505
R36253 PAD.n4304 PAD.n4303 2.2505
R36254 PAD.n4302 PAD.n4031 2.2505
R36255 PAD.n4301 PAD.n4300 2.2505
R36256 PAD.n4296 PAD.n4032 2.2505
R36257 PAD.n4292 PAD.n4291 2.2505
R36258 PAD.n4290 PAD.n4033 2.2505
R36259 PAD.n4289 PAD.n4288 2.2505
R36260 PAD.n4284 PAD.n4034 2.2505
R36261 PAD.n4280 PAD.n4279 2.2505
R36262 PAD.n4278 PAD.n4035 2.2505
R36263 PAD.n4277 PAD.n4276 2.2505
R36264 PAD.n4272 PAD.n4036 2.2505
R36265 PAD.n4268 PAD.n4267 2.2505
R36266 PAD.n4266 PAD.n4037 2.2505
R36267 PAD.n4265 PAD.n4264 2.2505
R36268 PAD.n4260 PAD.n4038 2.2505
R36269 PAD.n4256 PAD.n4255 2.2505
R36270 PAD.n4254 PAD.n4039 2.2505
R36271 PAD.n4253 PAD.n4252 2.2505
R36272 PAD.n4248 PAD.n4040 2.2505
R36273 PAD.n4244 PAD.n4243 2.2505
R36274 PAD.n4242 PAD.n4041 2.2505
R36275 PAD.n4241 PAD.n4240 2.2505
R36276 PAD.n4236 PAD.n4042 2.2505
R36277 PAD.n4232 PAD.n4231 2.2505
R36278 PAD.n4230 PAD.n4043 2.2505
R36279 PAD.n4229 PAD.n4228 2.2505
R36280 PAD.n4224 PAD.n4044 2.2505
R36281 PAD.n4220 PAD.n4219 2.2505
R36282 PAD.n4218 PAD.n4045 2.2505
R36283 PAD.n4217 PAD.n4216 2.2505
R36284 PAD.n4212 PAD.n4046 2.2505
R36285 PAD.n4208 PAD.n4207 2.2505
R36286 PAD.n4206 PAD.n4047 2.2505
R36287 PAD.n4205 PAD.n4204 2.2505
R36288 PAD.n4200 PAD.n4048 2.2505
R36289 PAD.n4196 PAD.n4195 2.2505
R36290 PAD.n4194 PAD.n4049 2.2505
R36291 PAD.n4193 PAD.n4192 2.2505
R36292 PAD.n4188 PAD.n4050 2.2505
R36293 PAD.n4184 PAD.n4183 2.2505
R36294 PAD.n4182 PAD.n4051 2.2505
R36295 PAD.n4181 PAD.n4180 2.2505
R36296 PAD.n4176 PAD.n4052 2.2505
R36297 PAD.n4172 PAD.n4171 2.2505
R36298 PAD.n4170 PAD.n4053 2.2505
R36299 PAD.n4169 PAD.n4168 2.2505
R36300 PAD.n4164 PAD.n4054 2.2505
R36301 PAD.n4160 PAD.n4159 2.2505
R36302 PAD.n4158 PAD.n4055 2.2505
R36303 PAD.n4157 PAD.n4156 2.2505
R36304 PAD.n4152 PAD.n4056 2.2505
R36305 PAD.n4148 PAD.n4147 2.2505
R36306 PAD.n4146 PAD.n4057 2.2505
R36307 PAD.n4145 PAD.n4144 2.2505
R36308 PAD.n4140 PAD.n4058 2.2505
R36309 PAD.n4136 PAD.n4135 2.2505
R36310 PAD.n4134 PAD.n4059 2.2505
R36311 PAD.n4133 PAD.n4132 2.2505
R36312 PAD.n4128 PAD.n4060 2.2505
R36313 PAD.n4124 PAD.n4123 2.2505
R36314 PAD.n4122 PAD.n4061 2.2505
R36315 PAD.n4121 PAD.n4120 2.2505
R36316 PAD.n4116 PAD.n4062 2.2505
R36317 PAD.n4112 PAD.n4111 2.2505
R36318 PAD.n4110 PAD.n4063 2.2505
R36319 PAD.n4109 PAD.n4108 2.2505
R36320 PAD.n4104 PAD.n4064 2.2505
R36321 PAD.n4100 PAD.n4099 2.2505
R36322 PAD.n4098 PAD.n4065 2.2505
R36323 PAD.n4097 PAD.n4096 2.2505
R36324 PAD.n4092 PAD.n4066 2.2505
R36325 PAD.n4088 PAD.n4087 2.2505
R36326 PAD.n4086 PAD.n4067 2.2505
R36327 PAD.n4085 PAD.n4084 2.2505
R36328 PAD.n4080 PAD.n4068 2.2505
R36329 PAD.n4076 PAD.n4075 2.2505
R36330 PAD.n4074 PAD.n4071 2.2505
R36331 PAD.n4073 PAD.n4072 2.2505
R36332 PAD.n4420 PAD.n4419 2.2505
R36333 PAD.n4422 PAD.n4418 2.2505
R36334 PAD.n4427 PAD.n4426 2.2505
R36335 PAD.n4424 PAD.n4416 2.2505
R36336 PAD.n4432 PAD.n4431 2.2505
R36337 PAD.n4434 PAD.n4414 2.2505
R36338 PAD.n4439 PAD.n4438 2.2505
R36339 PAD.n4436 PAD.n4412 2.2505
R36340 PAD.n4444 PAD.n4443 2.2505
R36341 PAD.n4446 PAD.n4410 2.2505
R36342 PAD.n4451 PAD.n4450 2.2505
R36343 PAD.n4448 PAD.n4408 2.2505
R36344 PAD.n4456 PAD.n4455 2.2505
R36345 PAD.n4458 PAD.n4406 2.2505
R36346 PAD.n4463 PAD.n4462 2.2505
R36347 PAD.n4460 PAD.n4404 2.2505
R36348 PAD.n4468 PAD.n4467 2.2505
R36349 PAD.n4470 PAD.n4402 2.2505
R36350 PAD.n4475 PAD.n4474 2.2505
R36351 PAD.n4472 PAD.n4400 2.2505
R36352 PAD.n4480 PAD.n4479 2.2505
R36353 PAD.n4482 PAD.n4398 2.2505
R36354 PAD.n4487 PAD.n4486 2.2505
R36355 PAD.n4484 PAD.n4396 2.2505
R36356 PAD.n4492 PAD.n4491 2.2505
R36357 PAD.n4494 PAD.n4394 2.2505
R36358 PAD.n4499 PAD.n4498 2.2505
R36359 PAD.n4496 PAD.n4392 2.2505
R36360 PAD.n4504 PAD.n4503 2.2505
R36361 PAD.n4506 PAD.n4390 2.2505
R36362 PAD.n4511 PAD.n4510 2.2505
R36363 PAD.n4508 PAD.n4388 2.2505
R36364 PAD.n4516 PAD.n4515 2.2505
R36365 PAD.n4518 PAD.n4386 2.2505
R36366 PAD.n4523 PAD.n4522 2.2505
R36367 PAD.n4520 PAD.n4384 2.2505
R36368 PAD.n4528 PAD.n4527 2.2505
R36369 PAD.n4530 PAD.n4382 2.2505
R36370 PAD.n4535 PAD.n4534 2.2505
R36371 PAD.n4532 PAD.n4380 2.2505
R36372 PAD.n4540 PAD.n4539 2.2505
R36373 PAD.n4542 PAD.n4378 2.2505
R36374 PAD.n4547 PAD.n4546 2.2505
R36375 PAD.n4544 PAD.n4376 2.2505
R36376 PAD.n4552 PAD.n4551 2.2505
R36377 PAD.n4554 PAD.n4374 2.2505
R36378 PAD.n4559 PAD.n4558 2.2505
R36379 PAD.n4556 PAD.n4372 2.2505
R36380 PAD.n4564 PAD.n4563 2.2505
R36381 PAD.n4566 PAD.n4370 2.2505
R36382 PAD.n4571 PAD.n4570 2.2505
R36383 PAD.n4568 PAD.n4368 2.2505
R36384 PAD.n4576 PAD.n4575 2.2505
R36385 PAD.n4578 PAD.n4366 2.2505
R36386 PAD.n4583 PAD.n4582 2.2505
R36387 PAD.n4580 PAD.n4364 2.2505
R36388 PAD.n4588 PAD.n4587 2.2505
R36389 PAD.n4590 PAD.n4362 2.2505
R36390 PAD.n4595 PAD.n4594 2.2505
R36391 PAD.n4592 PAD.n4360 2.2505
R36392 PAD.n4600 PAD.n4599 2.2505
R36393 PAD.n4602 PAD.n4358 2.2505
R36394 PAD.n4607 PAD.n4606 2.2505
R36395 PAD.n4604 PAD.n4356 2.2505
R36396 PAD.n4612 PAD.n4611 2.2505
R36397 PAD.n4614 PAD.n4354 2.2505
R36398 PAD.n4619 PAD.n4618 2.2505
R36399 PAD.n4616 PAD.n4352 2.2505
R36400 PAD.n4624 PAD.n4623 2.2505
R36401 PAD.n4626 PAD.n4350 2.2505
R36402 PAD.n4631 PAD.n4630 2.2505
R36403 PAD.n4628 PAD.n4348 2.2505
R36404 PAD.n4636 PAD.n4635 2.2505
R36405 PAD.n4638 PAD.n4346 2.2505
R36406 PAD.n4643 PAD.n4642 2.2505
R36407 PAD.n4640 PAD.n4344 2.2505
R36408 PAD.n4648 PAD.n4647 2.2505
R36409 PAD.n4650 PAD.n4342 2.2505
R36410 PAD.n4655 PAD.n4654 2.2505
R36411 PAD.n4652 PAD.n4340 2.2505
R36412 PAD.n4661 PAD.n4660 2.2505
R36413 PAD.n4663 PAD.n4338 2.2505
R36414 PAD.n4665 PAD.n4337 2.2505
R36415 PAD.n4668 PAD.n4667 2.2505
R36416 PAD.n4669 PAD.n4668 2.2505
R36417 PAD.n4337 PAD.n4336 2.2505
R36418 PAD.n4658 PAD.n4338 2.2505
R36419 PAD.n4660 PAD.n4659 2.2505
R36420 PAD.n4657 PAD.n4340 2.2505
R36421 PAD.n4656 PAD.n4655 2.2505
R36422 PAD.n4342 PAD.n4341 2.2505
R36423 PAD.n4647 PAD.n4646 2.2505
R36424 PAD.n4645 PAD.n4344 2.2505
R36425 PAD.n4644 PAD.n4643 2.2505
R36426 PAD.n4346 PAD.n4345 2.2505
R36427 PAD.n4635 PAD.n4634 2.2505
R36428 PAD.n4633 PAD.n4348 2.2505
R36429 PAD.n4632 PAD.n4631 2.2505
R36430 PAD.n4350 PAD.n4349 2.2505
R36431 PAD.n4623 PAD.n4622 2.2505
R36432 PAD.n4621 PAD.n4352 2.2505
R36433 PAD.n4620 PAD.n4619 2.2505
R36434 PAD.n4354 PAD.n4353 2.2505
R36435 PAD.n4611 PAD.n4610 2.2505
R36436 PAD.n4609 PAD.n4356 2.2505
R36437 PAD.n4608 PAD.n4607 2.2505
R36438 PAD.n4358 PAD.n4357 2.2505
R36439 PAD.n4599 PAD.n4598 2.2505
R36440 PAD.n4597 PAD.n4360 2.2505
R36441 PAD.n4596 PAD.n4595 2.2505
R36442 PAD.n4362 PAD.n4361 2.2505
R36443 PAD.n4587 PAD.n4586 2.2505
R36444 PAD.n4585 PAD.n4364 2.2505
R36445 PAD.n4584 PAD.n4583 2.2505
R36446 PAD.n4366 PAD.n4365 2.2505
R36447 PAD.n4575 PAD.n4574 2.2505
R36448 PAD.n4573 PAD.n4368 2.2505
R36449 PAD.n4572 PAD.n4571 2.2505
R36450 PAD.n4370 PAD.n4369 2.2505
R36451 PAD.n4563 PAD.n4562 2.2505
R36452 PAD.n4561 PAD.n4372 2.2505
R36453 PAD.n4560 PAD.n4559 2.2505
R36454 PAD.n4374 PAD.n4373 2.2505
R36455 PAD.n4551 PAD.n4550 2.2505
R36456 PAD.n4549 PAD.n4376 2.2505
R36457 PAD.n4548 PAD.n4547 2.2505
R36458 PAD.n4378 PAD.n4377 2.2505
R36459 PAD.n4539 PAD.n4538 2.2505
R36460 PAD.n4537 PAD.n4380 2.2505
R36461 PAD.n4536 PAD.n4535 2.2505
R36462 PAD.n4382 PAD.n4381 2.2505
R36463 PAD.n4527 PAD.n4526 2.2505
R36464 PAD.n4525 PAD.n4384 2.2505
R36465 PAD.n4524 PAD.n4523 2.2505
R36466 PAD.n4386 PAD.n4385 2.2505
R36467 PAD.n4515 PAD.n4514 2.2505
R36468 PAD.n4513 PAD.n4388 2.2505
R36469 PAD.n4512 PAD.n4511 2.2505
R36470 PAD.n4390 PAD.n4389 2.2505
R36471 PAD.n4503 PAD.n4502 2.2505
R36472 PAD.n4501 PAD.n4392 2.2505
R36473 PAD.n4500 PAD.n4499 2.2505
R36474 PAD.n4394 PAD.n4393 2.2505
R36475 PAD.n4491 PAD.n4490 2.2505
R36476 PAD.n4489 PAD.n4396 2.2505
R36477 PAD.n4488 PAD.n4487 2.2505
R36478 PAD.n4398 PAD.n4397 2.2505
R36479 PAD.n4479 PAD.n4478 2.2505
R36480 PAD.n4477 PAD.n4400 2.2505
R36481 PAD.n4476 PAD.n4475 2.2505
R36482 PAD.n4402 PAD.n4401 2.2505
R36483 PAD.n4467 PAD.n4466 2.2505
R36484 PAD.n4465 PAD.n4404 2.2505
R36485 PAD.n4464 PAD.n4463 2.2505
R36486 PAD.n4406 PAD.n4405 2.2505
R36487 PAD.n4455 PAD.n4454 2.2505
R36488 PAD.n4453 PAD.n4408 2.2505
R36489 PAD.n4452 PAD.n4451 2.2505
R36490 PAD.n4410 PAD.n4409 2.2505
R36491 PAD.n4443 PAD.n4442 2.2505
R36492 PAD.n4441 PAD.n4412 2.2505
R36493 PAD.n4440 PAD.n4439 2.2505
R36494 PAD.n4414 PAD.n4413 2.2505
R36495 PAD.n4431 PAD.n4430 2.2505
R36496 PAD.n4429 PAD.n4416 2.2505
R36497 PAD.n4428 PAD.n4427 2.2505
R36498 PAD.n4418 PAD.n4417 2.2505
R36499 PAD.n4419 PAD.n4325 2.2505
R36500 PAD.n8395 PAD.n8394 2.2505
R36501 PAD.n8393 PAD.n4725 2.2505
R36502 PAD.n4728 PAD.n4727 2.2505
R36503 PAD.n8389 PAD.n8388 2.2505
R36504 PAD.n8386 PAD.n8385 2.2505
R36505 PAD.n8384 PAD.n4733 2.2505
R36506 PAD.n4731 PAD.n4730 2.2505
R36507 PAD.n8380 PAD.n8379 2.2505
R36508 PAD.n8377 PAD.n8376 2.2505
R36509 PAD.n8375 PAD.n4738 2.2505
R36510 PAD.n4736 PAD.n4735 2.2505
R36511 PAD.n8371 PAD.n8370 2.2505
R36512 PAD.n8368 PAD.n8367 2.2505
R36513 PAD.n8366 PAD.n4743 2.2505
R36514 PAD.n4741 PAD.n4740 2.2505
R36515 PAD.n8362 PAD.n8361 2.2505
R36516 PAD.n8359 PAD.n8358 2.2505
R36517 PAD.n8357 PAD.n4748 2.2505
R36518 PAD.n4746 PAD.n4745 2.2505
R36519 PAD.n8353 PAD.n8352 2.2505
R36520 PAD.n8350 PAD.n8349 2.2505
R36521 PAD.n8348 PAD.n4753 2.2505
R36522 PAD.n4751 PAD.n4750 2.2505
R36523 PAD.n8344 PAD.n8343 2.2505
R36524 PAD.n8341 PAD.n8340 2.2505
R36525 PAD.n8339 PAD.n4758 2.2505
R36526 PAD.n4756 PAD.n4755 2.2505
R36527 PAD.n8335 PAD.n8334 2.2505
R36528 PAD.n8332 PAD.n8331 2.2505
R36529 PAD.n8330 PAD.n4763 2.2505
R36530 PAD.n4761 PAD.n4760 2.2505
R36531 PAD.n8326 PAD.n8325 2.2505
R36532 PAD.n8323 PAD.n8322 2.2505
R36533 PAD.n8321 PAD.n4768 2.2505
R36534 PAD.n4766 PAD.n4765 2.2505
R36535 PAD.n8317 PAD.n8316 2.2505
R36536 PAD.n8314 PAD.n8313 2.2505
R36537 PAD.n8312 PAD.n4773 2.2505
R36538 PAD.n4771 PAD.n4770 2.2505
R36539 PAD.n8308 PAD.n8307 2.2505
R36540 PAD.n8305 PAD.n8304 2.2505
R36541 PAD.n8303 PAD.n4778 2.2505
R36542 PAD.n4776 PAD.n4775 2.2505
R36543 PAD.n8299 PAD.n8298 2.2505
R36544 PAD.n8296 PAD.n8295 2.2505
R36545 PAD.n8294 PAD.n4783 2.2505
R36546 PAD.n4781 PAD.n4780 2.2505
R36547 PAD.n8290 PAD.n8289 2.2505
R36548 PAD.n8287 PAD.n8286 2.2505
R36549 PAD.n8285 PAD.n4788 2.2505
R36550 PAD.n4786 PAD.n4785 2.2505
R36551 PAD.n8281 PAD.n8280 2.2505
R36552 PAD.n8278 PAD.n8277 2.2505
R36553 PAD.n8276 PAD.n4793 2.2505
R36554 PAD.n4791 PAD.n4790 2.2505
R36555 PAD.n8272 PAD.n8271 2.2505
R36556 PAD.n8269 PAD.n8268 2.2505
R36557 PAD.n8267 PAD.n4798 2.2505
R36558 PAD.n4796 PAD.n4795 2.2505
R36559 PAD.n8263 PAD.n8262 2.2505
R36560 PAD.n8260 PAD.n8259 2.2505
R36561 PAD.n8258 PAD.n4803 2.2505
R36562 PAD.n4801 PAD.n4800 2.2505
R36563 PAD.n8254 PAD.n8253 2.2505
R36564 PAD.n8251 PAD.n8250 2.2505
R36565 PAD.n8249 PAD.n4808 2.2505
R36566 PAD.n4806 PAD.n4805 2.2505
R36567 PAD.n8245 PAD.n8244 2.2505
R36568 PAD.n8242 PAD.n8241 2.2505
R36569 PAD.n8240 PAD.n4813 2.2505
R36570 PAD.n4811 PAD.n4810 2.2505
R36571 PAD.n8236 PAD.n8235 2.2505
R36572 PAD.n8233 PAD.n8232 2.2505
R36573 PAD.n8231 PAD.n4818 2.2505
R36574 PAD.n4816 PAD.n4815 2.2505
R36575 PAD.n8227 PAD.n8226 2.2505
R36576 PAD.n8224 PAD.n8223 2.2505
R36577 PAD.n8222 PAD.n4823 2.2505
R36578 PAD.n4821 PAD.n4820 2.2505
R36579 PAD.n8218 PAD.n8217 2.2505
R36580 PAD.n8215 PAD.n8214 2.2505
R36581 PAD.n8213 PAD.n4828 2.2505
R36582 PAD.n4826 PAD.n4825 2.2505
R36583 PAD.n4832 PAD.n4829 2.2505
R36584 PAD.n8210 PAD.n4829 2.2505
R36585 PAD.n8211 PAD.n4825 2.2505
R36586 PAD.n8213 PAD.n8212 2.2505
R36587 PAD.n8214 PAD.n4824 2.2505
R36588 PAD.n8219 PAD.n8218 2.2505
R36589 PAD.n8220 PAD.n4820 2.2505
R36590 PAD.n8222 PAD.n8221 2.2505
R36591 PAD.n8223 PAD.n4819 2.2505
R36592 PAD.n8228 PAD.n8227 2.2505
R36593 PAD.n8229 PAD.n4815 2.2505
R36594 PAD.n8231 PAD.n8230 2.2505
R36595 PAD.n8232 PAD.n4814 2.2505
R36596 PAD.n8237 PAD.n8236 2.2505
R36597 PAD.n8238 PAD.n4810 2.2505
R36598 PAD.n8240 PAD.n8239 2.2505
R36599 PAD.n8241 PAD.n4809 2.2505
R36600 PAD.n8246 PAD.n8245 2.2505
R36601 PAD.n8247 PAD.n4805 2.2505
R36602 PAD.n8249 PAD.n8248 2.2505
R36603 PAD.n8250 PAD.n4804 2.2505
R36604 PAD.n8255 PAD.n8254 2.2505
R36605 PAD.n8256 PAD.n4800 2.2505
R36606 PAD.n8258 PAD.n8257 2.2505
R36607 PAD.n8259 PAD.n4799 2.2505
R36608 PAD.n8264 PAD.n8263 2.2505
R36609 PAD.n8265 PAD.n4795 2.2505
R36610 PAD.n8267 PAD.n8266 2.2505
R36611 PAD.n8268 PAD.n4794 2.2505
R36612 PAD.n8273 PAD.n8272 2.2505
R36613 PAD.n8274 PAD.n4790 2.2505
R36614 PAD.n8276 PAD.n8275 2.2505
R36615 PAD.n8277 PAD.n4789 2.2505
R36616 PAD.n8282 PAD.n8281 2.2505
R36617 PAD.n8283 PAD.n4785 2.2505
R36618 PAD.n8285 PAD.n8284 2.2505
R36619 PAD.n8286 PAD.n4784 2.2505
R36620 PAD.n8291 PAD.n8290 2.2505
R36621 PAD.n8292 PAD.n4780 2.2505
R36622 PAD.n8294 PAD.n8293 2.2505
R36623 PAD.n8295 PAD.n4779 2.2505
R36624 PAD.n8300 PAD.n8299 2.2505
R36625 PAD.n8301 PAD.n4775 2.2505
R36626 PAD.n8303 PAD.n8302 2.2505
R36627 PAD.n8304 PAD.n4774 2.2505
R36628 PAD.n8309 PAD.n8308 2.2505
R36629 PAD.n8310 PAD.n4770 2.2505
R36630 PAD.n8312 PAD.n8311 2.2505
R36631 PAD.n8313 PAD.n4769 2.2505
R36632 PAD.n8318 PAD.n8317 2.2505
R36633 PAD.n8319 PAD.n4765 2.2505
R36634 PAD.n8321 PAD.n8320 2.2505
R36635 PAD.n8322 PAD.n4764 2.2505
R36636 PAD.n8327 PAD.n8326 2.2505
R36637 PAD.n8328 PAD.n4760 2.2505
R36638 PAD.n8330 PAD.n8329 2.2505
R36639 PAD.n8331 PAD.n4759 2.2505
R36640 PAD.n8336 PAD.n8335 2.2505
R36641 PAD.n8337 PAD.n4755 2.2505
R36642 PAD.n8339 PAD.n8338 2.2505
R36643 PAD.n8340 PAD.n4754 2.2505
R36644 PAD.n8345 PAD.n8344 2.2505
R36645 PAD.n8346 PAD.n4750 2.2505
R36646 PAD.n8348 PAD.n8347 2.2505
R36647 PAD.n8349 PAD.n4749 2.2505
R36648 PAD.n8354 PAD.n8353 2.2505
R36649 PAD.n8355 PAD.n4745 2.2505
R36650 PAD.n8357 PAD.n8356 2.2505
R36651 PAD.n8358 PAD.n4744 2.2505
R36652 PAD.n8363 PAD.n8362 2.2505
R36653 PAD.n8364 PAD.n4740 2.2505
R36654 PAD.n8366 PAD.n8365 2.2505
R36655 PAD.n8367 PAD.n4739 2.2505
R36656 PAD.n8372 PAD.n8371 2.2505
R36657 PAD.n8373 PAD.n4735 2.2505
R36658 PAD.n8375 PAD.n8374 2.2505
R36659 PAD.n8376 PAD.n4734 2.2505
R36660 PAD.n8381 PAD.n8380 2.2505
R36661 PAD.n8382 PAD.n4730 2.2505
R36662 PAD.n8384 PAD.n8383 2.2505
R36663 PAD.n8385 PAD.n4729 2.2505
R36664 PAD.n8390 PAD.n8389 2.2505
R36665 PAD.n8391 PAD.n4728 2.2505
R36666 PAD.n8393 PAD.n8392 2.2505
R36667 PAD.n8394 PAD.n4676 2.2505
R36668 PAD.n5178 PAD.n4847 2.2505
R36669 PAD.n5177 PAD.n5176 2.2505
R36670 PAD.n5174 PAD.n4848 2.2505
R36671 PAD.n5172 PAD.n5171 2.2505
R36672 PAD.n5164 PAD.n4851 2.2505
R36673 PAD.n5167 PAD.n5166 2.2505
R36674 PAD.n5162 PAD.n4854 2.2505
R36675 PAD.n5160 PAD.n5159 2.2505
R36676 PAD.n5152 PAD.n4856 2.2505
R36677 PAD.n5155 PAD.n5154 2.2505
R36678 PAD.n5150 PAD.n4858 2.2505
R36679 PAD.n5148 PAD.n5147 2.2505
R36680 PAD.n5140 PAD.n4860 2.2505
R36681 PAD.n5143 PAD.n5142 2.2505
R36682 PAD.n5138 PAD.n4862 2.2505
R36683 PAD.n5136 PAD.n5135 2.2505
R36684 PAD.n5128 PAD.n4864 2.2505
R36685 PAD.n5131 PAD.n5130 2.2505
R36686 PAD.n5126 PAD.n4866 2.2505
R36687 PAD.n5124 PAD.n5123 2.2505
R36688 PAD.n5116 PAD.n4868 2.2505
R36689 PAD.n5119 PAD.n5118 2.2505
R36690 PAD.n5114 PAD.n4870 2.2505
R36691 PAD.n5112 PAD.n5111 2.2505
R36692 PAD.n5104 PAD.n4872 2.2505
R36693 PAD.n5107 PAD.n5106 2.2505
R36694 PAD.n5102 PAD.n4874 2.2505
R36695 PAD.n5100 PAD.n5099 2.2505
R36696 PAD.n5092 PAD.n4876 2.2505
R36697 PAD.n5095 PAD.n5094 2.2505
R36698 PAD.n5090 PAD.n4878 2.2505
R36699 PAD.n5088 PAD.n5087 2.2505
R36700 PAD.n5080 PAD.n4880 2.2505
R36701 PAD.n5083 PAD.n5082 2.2505
R36702 PAD.n5078 PAD.n4882 2.2505
R36703 PAD.n5076 PAD.n5075 2.2505
R36704 PAD.n5068 PAD.n4884 2.2505
R36705 PAD.n5071 PAD.n5070 2.2505
R36706 PAD.n5066 PAD.n4886 2.2505
R36707 PAD.n5064 PAD.n5063 2.2505
R36708 PAD.n5056 PAD.n4888 2.2505
R36709 PAD.n5059 PAD.n5058 2.2505
R36710 PAD.n5054 PAD.n4890 2.2505
R36711 PAD.n5052 PAD.n5051 2.2505
R36712 PAD.n5044 PAD.n4892 2.2505
R36713 PAD.n5047 PAD.n5046 2.2505
R36714 PAD.n5042 PAD.n4894 2.2505
R36715 PAD.n5040 PAD.n5039 2.2505
R36716 PAD.n5032 PAD.n4896 2.2505
R36717 PAD.n5035 PAD.n5034 2.2505
R36718 PAD.n5030 PAD.n4898 2.2505
R36719 PAD.n5028 PAD.n5027 2.2505
R36720 PAD.n5020 PAD.n4900 2.2505
R36721 PAD.n5023 PAD.n5022 2.2505
R36722 PAD.n5018 PAD.n4902 2.2505
R36723 PAD.n5016 PAD.n5015 2.2505
R36724 PAD.n5008 PAD.n4904 2.2505
R36725 PAD.n5011 PAD.n5010 2.2505
R36726 PAD.n5006 PAD.n4906 2.2505
R36727 PAD.n5004 PAD.n5003 2.2505
R36728 PAD.n4996 PAD.n4908 2.2505
R36729 PAD.n4999 PAD.n4998 2.2505
R36730 PAD.n4994 PAD.n4910 2.2505
R36731 PAD.n4992 PAD.n4991 2.2505
R36732 PAD.n4984 PAD.n4912 2.2505
R36733 PAD.n4987 PAD.n4986 2.2505
R36734 PAD.n4982 PAD.n4914 2.2505
R36735 PAD.n4980 PAD.n4979 2.2505
R36736 PAD.n4972 PAD.n4916 2.2505
R36737 PAD.n4975 PAD.n4974 2.2505
R36738 PAD.n4970 PAD.n4918 2.2505
R36739 PAD.n4968 PAD.n4967 2.2505
R36740 PAD.n4960 PAD.n4920 2.2505
R36741 PAD.n4963 PAD.n4962 2.2505
R36742 PAD.n4958 PAD.n4922 2.2505
R36743 PAD.n4956 PAD.n4955 2.2505
R36744 PAD.n4948 PAD.n4924 2.2505
R36745 PAD.n4951 PAD.n4950 2.2505
R36746 PAD.n4946 PAD.n4926 2.2505
R36747 PAD.n4944 PAD.n4943 2.2505
R36748 PAD.n4936 PAD.n4928 2.2505
R36749 PAD.n4939 PAD.n4938 2.2505
R36750 PAD.n4934 PAD.n4930 2.2505
R36751 PAD.n4932 PAD.n4931 2.2505
R36752 PAD.n4931 PAD.n4835 2.2505
R36753 PAD.n4930 PAD.n4929 2.2505
R36754 PAD.n4940 PAD.n4939 2.2505
R36755 PAD.n4941 PAD.n4928 2.2505
R36756 PAD.n4943 PAD.n4942 2.2505
R36757 PAD.n4926 PAD.n4925 2.2505
R36758 PAD.n4952 PAD.n4951 2.2505
R36759 PAD.n4953 PAD.n4924 2.2505
R36760 PAD.n4955 PAD.n4954 2.2505
R36761 PAD.n4922 PAD.n4921 2.2505
R36762 PAD.n4964 PAD.n4963 2.2505
R36763 PAD.n4965 PAD.n4920 2.2505
R36764 PAD.n4967 PAD.n4966 2.2505
R36765 PAD.n4918 PAD.n4917 2.2505
R36766 PAD.n4976 PAD.n4975 2.2505
R36767 PAD.n4977 PAD.n4916 2.2505
R36768 PAD.n4979 PAD.n4978 2.2505
R36769 PAD.n4914 PAD.n4913 2.2505
R36770 PAD.n4988 PAD.n4987 2.2505
R36771 PAD.n4989 PAD.n4912 2.2505
R36772 PAD.n4991 PAD.n4990 2.2505
R36773 PAD.n4910 PAD.n4909 2.2505
R36774 PAD.n5000 PAD.n4999 2.2505
R36775 PAD.n5001 PAD.n4908 2.2505
R36776 PAD.n5003 PAD.n5002 2.2505
R36777 PAD.n4906 PAD.n4905 2.2505
R36778 PAD.n5012 PAD.n5011 2.2505
R36779 PAD.n5013 PAD.n4904 2.2505
R36780 PAD.n5015 PAD.n5014 2.2505
R36781 PAD.n4902 PAD.n4901 2.2505
R36782 PAD.n5024 PAD.n5023 2.2505
R36783 PAD.n5025 PAD.n4900 2.2505
R36784 PAD.n5027 PAD.n5026 2.2505
R36785 PAD.n4898 PAD.n4897 2.2505
R36786 PAD.n5036 PAD.n5035 2.2505
R36787 PAD.n5037 PAD.n4896 2.2505
R36788 PAD.n5039 PAD.n5038 2.2505
R36789 PAD.n4894 PAD.n4893 2.2505
R36790 PAD.n5048 PAD.n5047 2.2505
R36791 PAD.n5049 PAD.n4892 2.2505
R36792 PAD.n5051 PAD.n5050 2.2505
R36793 PAD.n4890 PAD.n4889 2.2505
R36794 PAD.n5060 PAD.n5059 2.2505
R36795 PAD.n5061 PAD.n4888 2.2505
R36796 PAD.n5063 PAD.n5062 2.2505
R36797 PAD.n4886 PAD.n4885 2.2505
R36798 PAD.n5072 PAD.n5071 2.2505
R36799 PAD.n5073 PAD.n4884 2.2505
R36800 PAD.n5075 PAD.n5074 2.2505
R36801 PAD.n4882 PAD.n4881 2.2505
R36802 PAD.n5084 PAD.n5083 2.2505
R36803 PAD.n5085 PAD.n4880 2.2505
R36804 PAD.n5087 PAD.n5086 2.2505
R36805 PAD.n4878 PAD.n4877 2.2505
R36806 PAD.n5096 PAD.n5095 2.2505
R36807 PAD.n5097 PAD.n4876 2.2505
R36808 PAD.n5099 PAD.n5098 2.2505
R36809 PAD.n4874 PAD.n4873 2.2505
R36810 PAD.n5108 PAD.n5107 2.2505
R36811 PAD.n5109 PAD.n4872 2.2505
R36812 PAD.n5111 PAD.n5110 2.2505
R36813 PAD.n4870 PAD.n4869 2.2505
R36814 PAD.n5120 PAD.n5119 2.2505
R36815 PAD.n5121 PAD.n4868 2.2505
R36816 PAD.n5123 PAD.n5122 2.2505
R36817 PAD.n4866 PAD.n4865 2.2505
R36818 PAD.n5132 PAD.n5131 2.2505
R36819 PAD.n5133 PAD.n4864 2.2505
R36820 PAD.n5135 PAD.n5134 2.2505
R36821 PAD.n4862 PAD.n4861 2.2505
R36822 PAD.n5144 PAD.n5143 2.2505
R36823 PAD.n5145 PAD.n4860 2.2505
R36824 PAD.n5147 PAD.n5146 2.2505
R36825 PAD.n4858 PAD.n4857 2.2505
R36826 PAD.n5156 PAD.n5155 2.2505
R36827 PAD.n5157 PAD.n4856 2.2505
R36828 PAD.n5159 PAD.n5158 2.2505
R36829 PAD.n4854 PAD.n4853 2.2505
R36830 PAD.n5168 PAD.n5167 2.2505
R36831 PAD.n5169 PAD.n4851 2.2505
R36832 PAD.n5171 PAD.n5170 2.2505
R36833 PAD.n4852 PAD.n4848 2.2505
R36834 PAD.n5177 PAD.n4846 2.2505
R36835 PAD.n5179 PAD.n5178 2.2505
R36836 PAD.n8161 PAD.n8160 2.2505
R36837 PAD.n8159 PAD.n7871 2.2505
R36838 PAD.n7874 PAD.n7873 2.2505
R36839 PAD.n8155 PAD.n8154 2.2505
R36840 PAD.n8152 PAD.n8151 2.2505
R36841 PAD.n8150 PAD.n7879 2.2505
R36842 PAD.n7877 PAD.n7876 2.2505
R36843 PAD.n8146 PAD.n8145 2.2505
R36844 PAD.n8143 PAD.n8142 2.2505
R36845 PAD.n8141 PAD.n7884 2.2505
R36846 PAD.n7882 PAD.n7881 2.2505
R36847 PAD.n8137 PAD.n8136 2.2505
R36848 PAD.n8134 PAD.n8133 2.2505
R36849 PAD.n8132 PAD.n7889 2.2505
R36850 PAD.n7887 PAD.n7886 2.2505
R36851 PAD.n8128 PAD.n8127 2.2505
R36852 PAD.n8125 PAD.n8124 2.2505
R36853 PAD.n8123 PAD.n7894 2.2505
R36854 PAD.n7892 PAD.n7891 2.2505
R36855 PAD.n8119 PAD.n8118 2.2505
R36856 PAD.n8116 PAD.n8115 2.2505
R36857 PAD.n8114 PAD.n7899 2.2505
R36858 PAD.n7897 PAD.n7896 2.2505
R36859 PAD.n8110 PAD.n8109 2.2505
R36860 PAD.n8107 PAD.n8106 2.2505
R36861 PAD.n8105 PAD.n7904 2.2505
R36862 PAD.n7902 PAD.n7901 2.2505
R36863 PAD.n8101 PAD.n8100 2.2505
R36864 PAD.n8098 PAD.n8097 2.2505
R36865 PAD.n8096 PAD.n7909 2.2505
R36866 PAD.n7907 PAD.n7906 2.2505
R36867 PAD.n8092 PAD.n8091 2.2505
R36868 PAD.n8089 PAD.n8088 2.2505
R36869 PAD.n8087 PAD.n7914 2.2505
R36870 PAD.n7912 PAD.n7911 2.2505
R36871 PAD.n8083 PAD.n8082 2.2505
R36872 PAD.n8080 PAD.n8079 2.2505
R36873 PAD.n8078 PAD.n7919 2.2505
R36874 PAD.n7917 PAD.n7916 2.2505
R36875 PAD.n8074 PAD.n8073 2.2505
R36876 PAD.n8071 PAD.n8070 2.2505
R36877 PAD.n8069 PAD.n7924 2.2505
R36878 PAD.n7922 PAD.n7921 2.2505
R36879 PAD.n8065 PAD.n8064 2.2505
R36880 PAD.n8062 PAD.n8061 2.2505
R36881 PAD.n8060 PAD.n7929 2.2505
R36882 PAD.n7927 PAD.n7926 2.2505
R36883 PAD.n8056 PAD.n8055 2.2505
R36884 PAD.n8053 PAD.n8052 2.2505
R36885 PAD.n8051 PAD.n7934 2.2505
R36886 PAD.n7932 PAD.n7931 2.2505
R36887 PAD.n8047 PAD.n8046 2.2505
R36888 PAD.n8044 PAD.n8043 2.2505
R36889 PAD.n8042 PAD.n7939 2.2505
R36890 PAD.n7937 PAD.n7936 2.2505
R36891 PAD.n8038 PAD.n8037 2.2505
R36892 PAD.n8035 PAD.n8034 2.2505
R36893 PAD.n8033 PAD.n7944 2.2505
R36894 PAD.n7942 PAD.n7941 2.2505
R36895 PAD.n8029 PAD.n8028 2.2505
R36896 PAD.n8026 PAD.n8025 2.2505
R36897 PAD.n8024 PAD.n7949 2.2505
R36898 PAD.n7947 PAD.n7946 2.2505
R36899 PAD.n8020 PAD.n8019 2.2505
R36900 PAD.n8017 PAD.n8016 2.2505
R36901 PAD.n8015 PAD.n7954 2.2505
R36902 PAD.n7952 PAD.n7951 2.2505
R36903 PAD.n8011 PAD.n8010 2.2505
R36904 PAD.n8008 PAD.n8007 2.2505
R36905 PAD.n8006 PAD.n7959 2.2505
R36906 PAD.n7957 PAD.n7956 2.2505
R36907 PAD.n8002 PAD.n8001 2.2505
R36908 PAD.n7999 PAD.n7998 2.2505
R36909 PAD.n7997 PAD.n7964 2.2505
R36910 PAD.n7962 PAD.n7961 2.2505
R36911 PAD.n7993 PAD.n7992 2.2505
R36912 PAD.n7990 PAD.n7989 2.2505
R36913 PAD.n7988 PAD.n7969 2.2505
R36914 PAD.n7967 PAD.n7966 2.2505
R36915 PAD.n7984 PAD.n7983 2.2505
R36916 PAD.n7981 PAD.n7980 2.2505
R36917 PAD.n7979 PAD.n7976 2.2505
R36918 PAD.n7974 PAD.n7973 2.2505
R36919 PAD.n7972 PAD.n7971 2.2505
R36920 PAD.n7972 PAD.n5186 2.2505
R36921 PAD.n7977 PAD.n7973 2.2505
R36922 PAD.n7979 PAD.n7978 2.2505
R36923 PAD.n7980 PAD.n7970 2.2505
R36924 PAD.n7985 PAD.n7984 2.2505
R36925 PAD.n7986 PAD.n7966 2.2505
R36926 PAD.n7988 PAD.n7987 2.2505
R36927 PAD.n7989 PAD.n7965 2.2505
R36928 PAD.n7994 PAD.n7993 2.2505
R36929 PAD.n7995 PAD.n7961 2.2505
R36930 PAD.n7997 PAD.n7996 2.2505
R36931 PAD.n7998 PAD.n7960 2.2505
R36932 PAD.n8003 PAD.n8002 2.2505
R36933 PAD.n8004 PAD.n7956 2.2505
R36934 PAD.n8006 PAD.n8005 2.2505
R36935 PAD.n8007 PAD.n7955 2.2505
R36936 PAD.n8012 PAD.n8011 2.2505
R36937 PAD.n8013 PAD.n7951 2.2505
R36938 PAD.n8015 PAD.n8014 2.2505
R36939 PAD.n8016 PAD.n7950 2.2505
R36940 PAD.n8021 PAD.n8020 2.2505
R36941 PAD.n8022 PAD.n7946 2.2505
R36942 PAD.n8024 PAD.n8023 2.2505
R36943 PAD.n8025 PAD.n7945 2.2505
R36944 PAD.n8030 PAD.n8029 2.2505
R36945 PAD.n8031 PAD.n7941 2.2505
R36946 PAD.n8033 PAD.n8032 2.2505
R36947 PAD.n8034 PAD.n7940 2.2505
R36948 PAD.n8039 PAD.n8038 2.2505
R36949 PAD.n8040 PAD.n7936 2.2505
R36950 PAD.n8042 PAD.n8041 2.2505
R36951 PAD.n8043 PAD.n7935 2.2505
R36952 PAD.n8048 PAD.n8047 2.2505
R36953 PAD.n8049 PAD.n7931 2.2505
R36954 PAD.n8051 PAD.n8050 2.2505
R36955 PAD.n8052 PAD.n7930 2.2505
R36956 PAD.n8057 PAD.n8056 2.2505
R36957 PAD.n8058 PAD.n7926 2.2505
R36958 PAD.n8060 PAD.n8059 2.2505
R36959 PAD.n8061 PAD.n7925 2.2505
R36960 PAD.n8066 PAD.n8065 2.2505
R36961 PAD.n8067 PAD.n7921 2.2505
R36962 PAD.n8069 PAD.n8068 2.2505
R36963 PAD.n8070 PAD.n7920 2.2505
R36964 PAD.n8075 PAD.n8074 2.2505
R36965 PAD.n8076 PAD.n7916 2.2505
R36966 PAD.n8078 PAD.n8077 2.2505
R36967 PAD.n8079 PAD.n7915 2.2505
R36968 PAD.n8084 PAD.n8083 2.2505
R36969 PAD.n8085 PAD.n7911 2.2505
R36970 PAD.n8087 PAD.n8086 2.2505
R36971 PAD.n8088 PAD.n7910 2.2505
R36972 PAD.n8093 PAD.n8092 2.2505
R36973 PAD.n8094 PAD.n7906 2.2505
R36974 PAD.n8096 PAD.n8095 2.2505
R36975 PAD.n8097 PAD.n7905 2.2505
R36976 PAD.n8102 PAD.n8101 2.2505
R36977 PAD.n8103 PAD.n7901 2.2505
R36978 PAD.n8105 PAD.n8104 2.2505
R36979 PAD.n8106 PAD.n7900 2.2505
R36980 PAD.n8111 PAD.n8110 2.2505
R36981 PAD.n8112 PAD.n7896 2.2505
R36982 PAD.n8114 PAD.n8113 2.2505
R36983 PAD.n8115 PAD.n7895 2.2505
R36984 PAD.n8120 PAD.n8119 2.2505
R36985 PAD.n8121 PAD.n7891 2.2505
R36986 PAD.n8123 PAD.n8122 2.2505
R36987 PAD.n8124 PAD.n7890 2.2505
R36988 PAD.n8129 PAD.n8128 2.2505
R36989 PAD.n8130 PAD.n7886 2.2505
R36990 PAD.n8132 PAD.n8131 2.2505
R36991 PAD.n8133 PAD.n7885 2.2505
R36992 PAD.n8138 PAD.n8137 2.2505
R36993 PAD.n8139 PAD.n7881 2.2505
R36994 PAD.n8141 PAD.n8140 2.2505
R36995 PAD.n8142 PAD.n7880 2.2505
R36996 PAD.n8147 PAD.n8146 2.2505
R36997 PAD.n8148 PAD.n7876 2.2505
R36998 PAD.n8150 PAD.n8149 2.2505
R36999 PAD.n8151 PAD.n7875 2.2505
R37000 PAD.n8156 PAD.n8155 2.2505
R37001 PAD.n8157 PAD.n7874 2.2505
R37002 PAD.n8159 PAD.n8158 2.2505
R37003 PAD.n8160 PAD.n5193 2.2505
R37004 PAD.n5542 PAD.n5211 2.2505
R37005 PAD.n5541 PAD.n5540 2.2505
R37006 PAD.n5538 PAD.n5212 2.2505
R37007 PAD.n5536 PAD.n5535 2.2505
R37008 PAD.n5528 PAD.n5215 2.2505
R37009 PAD.n5531 PAD.n5530 2.2505
R37010 PAD.n5526 PAD.n5218 2.2505
R37011 PAD.n5524 PAD.n5523 2.2505
R37012 PAD.n5516 PAD.n5220 2.2505
R37013 PAD.n5519 PAD.n5518 2.2505
R37014 PAD.n5514 PAD.n5222 2.2505
R37015 PAD.n5512 PAD.n5511 2.2505
R37016 PAD.n5504 PAD.n5224 2.2505
R37017 PAD.n5507 PAD.n5506 2.2505
R37018 PAD.n5502 PAD.n5226 2.2505
R37019 PAD.n5500 PAD.n5499 2.2505
R37020 PAD.n5492 PAD.n5228 2.2505
R37021 PAD.n5495 PAD.n5494 2.2505
R37022 PAD.n5490 PAD.n5230 2.2505
R37023 PAD.n5488 PAD.n5487 2.2505
R37024 PAD.n5480 PAD.n5232 2.2505
R37025 PAD.n5483 PAD.n5482 2.2505
R37026 PAD.n5478 PAD.n5234 2.2505
R37027 PAD.n5476 PAD.n5475 2.2505
R37028 PAD.n5468 PAD.n5236 2.2505
R37029 PAD.n5471 PAD.n5470 2.2505
R37030 PAD.n5466 PAD.n5238 2.2505
R37031 PAD.n5464 PAD.n5463 2.2505
R37032 PAD.n5456 PAD.n5240 2.2505
R37033 PAD.n5459 PAD.n5458 2.2505
R37034 PAD.n5454 PAD.n5242 2.2505
R37035 PAD.n5452 PAD.n5451 2.2505
R37036 PAD.n5444 PAD.n5244 2.2505
R37037 PAD.n5447 PAD.n5446 2.2505
R37038 PAD.n5442 PAD.n5246 2.2505
R37039 PAD.n5440 PAD.n5439 2.2505
R37040 PAD.n5432 PAD.n5248 2.2505
R37041 PAD.n5435 PAD.n5434 2.2505
R37042 PAD.n5430 PAD.n5250 2.2505
R37043 PAD.n5428 PAD.n5427 2.2505
R37044 PAD.n5420 PAD.n5252 2.2505
R37045 PAD.n5423 PAD.n5422 2.2505
R37046 PAD.n5418 PAD.n5254 2.2505
R37047 PAD.n5416 PAD.n5415 2.2505
R37048 PAD.n5408 PAD.n5256 2.2505
R37049 PAD.n5411 PAD.n5410 2.2505
R37050 PAD.n5406 PAD.n5258 2.2505
R37051 PAD.n5404 PAD.n5403 2.2505
R37052 PAD.n5396 PAD.n5260 2.2505
R37053 PAD.n5399 PAD.n5398 2.2505
R37054 PAD.n5394 PAD.n5262 2.2505
R37055 PAD.n5392 PAD.n5391 2.2505
R37056 PAD.n5384 PAD.n5264 2.2505
R37057 PAD.n5387 PAD.n5386 2.2505
R37058 PAD.n5382 PAD.n5266 2.2505
R37059 PAD.n5380 PAD.n5379 2.2505
R37060 PAD.n5372 PAD.n5268 2.2505
R37061 PAD.n5375 PAD.n5374 2.2505
R37062 PAD.n5370 PAD.n5270 2.2505
R37063 PAD.n5368 PAD.n5367 2.2505
R37064 PAD.n5360 PAD.n5272 2.2505
R37065 PAD.n5363 PAD.n5362 2.2505
R37066 PAD.n5358 PAD.n5274 2.2505
R37067 PAD.n5356 PAD.n5355 2.2505
R37068 PAD.n5348 PAD.n5276 2.2505
R37069 PAD.n5351 PAD.n5350 2.2505
R37070 PAD.n5346 PAD.n5278 2.2505
R37071 PAD.n5344 PAD.n5343 2.2505
R37072 PAD.n5336 PAD.n5280 2.2505
R37073 PAD.n5339 PAD.n5338 2.2505
R37074 PAD.n5334 PAD.n5282 2.2505
R37075 PAD.n5332 PAD.n5331 2.2505
R37076 PAD.n5324 PAD.n5284 2.2505
R37077 PAD.n5327 PAD.n5326 2.2505
R37078 PAD.n5322 PAD.n5286 2.2505
R37079 PAD.n5320 PAD.n5319 2.2505
R37080 PAD.n5312 PAD.n5288 2.2505
R37081 PAD.n5315 PAD.n5314 2.2505
R37082 PAD.n5310 PAD.n5290 2.2505
R37083 PAD.n5308 PAD.n5307 2.2505
R37084 PAD.n5300 PAD.n5292 2.2505
R37085 PAD.n5303 PAD.n5302 2.2505
R37086 PAD.n5298 PAD.n5294 2.2505
R37087 PAD.n5296 PAD.n5295 2.2505
R37088 PAD.n5295 PAD.n5200 2.2505
R37089 PAD.n5294 PAD.n5293 2.2505
R37090 PAD.n5304 PAD.n5303 2.2505
R37091 PAD.n5305 PAD.n5292 2.2505
R37092 PAD.n5307 PAD.n5306 2.2505
R37093 PAD.n5290 PAD.n5289 2.2505
R37094 PAD.n5316 PAD.n5315 2.2505
R37095 PAD.n5317 PAD.n5288 2.2505
R37096 PAD.n5319 PAD.n5318 2.2505
R37097 PAD.n5286 PAD.n5285 2.2505
R37098 PAD.n5328 PAD.n5327 2.2505
R37099 PAD.n5329 PAD.n5284 2.2505
R37100 PAD.n5331 PAD.n5330 2.2505
R37101 PAD.n5282 PAD.n5281 2.2505
R37102 PAD.n5340 PAD.n5339 2.2505
R37103 PAD.n5341 PAD.n5280 2.2505
R37104 PAD.n5343 PAD.n5342 2.2505
R37105 PAD.n5278 PAD.n5277 2.2505
R37106 PAD.n5352 PAD.n5351 2.2505
R37107 PAD.n5353 PAD.n5276 2.2505
R37108 PAD.n5355 PAD.n5354 2.2505
R37109 PAD.n5274 PAD.n5273 2.2505
R37110 PAD.n5364 PAD.n5363 2.2505
R37111 PAD.n5365 PAD.n5272 2.2505
R37112 PAD.n5367 PAD.n5366 2.2505
R37113 PAD.n5270 PAD.n5269 2.2505
R37114 PAD.n5376 PAD.n5375 2.2505
R37115 PAD.n5377 PAD.n5268 2.2505
R37116 PAD.n5379 PAD.n5378 2.2505
R37117 PAD.n5266 PAD.n5265 2.2505
R37118 PAD.n5388 PAD.n5387 2.2505
R37119 PAD.n5389 PAD.n5264 2.2505
R37120 PAD.n5391 PAD.n5390 2.2505
R37121 PAD.n5262 PAD.n5261 2.2505
R37122 PAD.n5400 PAD.n5399 2.2505
R37123 PAD.n5401 PAD.n5260 2.2505
R37124 PAD.n5403 PAD.n5402 2.2505
R37125 PAD.n5258 PAD.n5257 2.2505
R37126 PAD.n5412 PAD.n5411 2.2505
R37127 PAD.n5413 PAD.n5256 2.2505
R37128 PAD.n5415 PAD.n5414 2.2505
R37129 PAD.n5254 PAD.n5253 2.2505
R37130 PAD.n5424 PAD.n5423 2.2505
R37131 PAD.n5425 PAD.n5252 2.2505
R37132 PAD.n5427 PAD.n5426 2.2505
R37133 PAD.n5250 PAD.n5249 2.2505
R37134 PAD.n5436 PAD.n5435 2.2505
R37135 PAD.n5437 PAD.n5248 2.2505
R37136 PAD.n5439 PAD.n5438 2.2505
R37137 PAD.n5246 PAD.n5245 2.2505
R37138 PAD.n5448 PAD.n5447 2.2505
R37139 PAD.n5449 PAD.n5244 2.2505
R37140 PAD.n5451 PAD.n5450 2.2505
R37141 PAD.n5242 PAD.n5241 2.2505
R37142 PAD.n5460 PAD.n5459 2.2505
R37143 PAD.n5461 PAD.n5240 2.2505
R37144 PAD.n5463 PAD.n5462 2.2505
R37145 PAD.n5238 PAD.n5237 2.2505
R37146 PAD.n5472 PAD.n5471 2.2505
R37147 PAD.n5473 PAD.n5236 2.2505
R37148 PAD.n5475 PAD.n5474 2.2505
R37149 PAD.n5234 PAD.n5233 2.2505
R37150 PAD.n5484 PAD.n5483 2.2505
R37151 PAD.n5485 PAD.n5232 2.2505
R37152 PAD.n5487 PAD.n5486 2.2505
R37153 PAD.n5230 PAD.n5229 2.2505
R37154 PAD.n5496 PAD.n5495 2.2505
R37155 PAD.n5497 PAD.n5228 2.2505
R37156 PAD.n5499 PAD.n5498 2.2505
R37157 PAD.n5226 PAD.n5225 2.2505
R37158 PAD.n5508 PAD.n5507 2.2505
R37159 PAD.n5509 PAD.n5224 2.2505
R37160 PAD.n5511 PAD.n5510 2.2505
R37161 PAD.n5222 PAD.n5221 2.2505
R37162 PAD.n5520 PAD.n5519 2.2505
R37163 PAD.n5521 PAD.n5220 2.2505
R37164 PAD.n5523 PAD.n5522 2.2505
R37165 PAD.n5218 PAD.n5217 2.2505
R37166 PAD.n5532 PAD.n5531 2.2505
R37167 PAD.n5533 PAD.n5215 2.2505
R37168 PAD.n5535 PAD.n5534 2.2505
R37169 PAD.n5216 PAD.n5212 2.2505
R37170 PAD.n5541 PAD.n5210 2.2505
R37171 PAD.n5543 PAD.n5542 2.2505
R37172 PAD.n7780 PAD.n7779 2.2505
R37173 PAD.n7106 PAD.n7104 2.2505
R37174 PAD.n7775 PAD.n7774 2.2505
R37175 PAD.n7772 PAD.n7771 2.2505
R37176 PAD.n7769 PAD.n7768 2.2505
R37177 PAD.n7761 PAD.n7108 2.2505
R37178 PAD.n7764 PAD.n7763 2.2505
R37179 PAD.n7760 PAD.n7759 2.2505
R37180 PAD.n7757 PAD.n7756 2.2505
R37181 PAD.n7749 PAD.n7110 2.2505
R37182 PAD.n7752 PAD.n7751 2.2505
R37183 PAD.n7748 PAD.n7747 2.2505
R37184 PAD.n7745 PAD.n7744 2.2505
R37185 PAD.n7737 PAD.n7112 2.2505
R37186 PAD.n7740 PAD.n7739 2.2505
R37187 PAD.n7736 PAD.n7735 2.2505
R37188 PAD.n7733 PAD.n7732 2.2505
R37189 PAD.n7725 PAD.n7114 2.2505
R37190 PAD.n7728 PAD.n7727 2.2505
R37191 PAD.n7724 PAD.n7723 2.2505
R37192 PAD.n7721 PAD.n7720 2.2505
R37193 PAD.n7713 PAD.n7116 2.2505
R37194 PAD.n7716 PAD.n7715 2.2505
R37195 PAD.n7712 PAD.n7711 2.2505
R37196 PAD.n7709 PAD.n7708 2.2505
R37197 PAD.n7701 PAD.n7118 2.2505
R37198 PAD.n7704 PAD.n7703 2.2505
R37199 PAD.n7700 PAD.n7699 2.2505
R37200 PAD.n7697 PAD.n7696 2.2505
R37201 PAD.n7689 PAD.n7120 2.2505
R37202 PAD.n7692 PAD.n7691 2.2505
R37203 PAD.n7688 PAD.n7687 2.2505
R37204 PAD.n7685 PAD.n7684 2.2505
R37205 PAD.n7677 PAD.n7122 2.2505
R37206 PAD.n7680 PAD.n7679 2.2505
R37207 PAD.n7676 PAD.n7675 2.2505
R37208 PAD.n7673 PAD.n7672 2.2505
R37209 PAD.n7665 PAD.n7124 2.2505
R37210 PAD.n7668 PAD.n7667 2.2505
R37211 PAD.n7664 PAD.n7663 2.2505
R37212 PAD.n7661 PAD.n7660 2.2505
R37213 PAD.n7653 PAD.n7126 2.2505
R37214 PAD.n7656 PAD.n7655 2.2505
R37215 PAD.n7652 PAD.n7651 2.2505
R37216 PAD.n7649 PAD.n7648 2.2505
R37217 PAD.n7641 PAD.n7128 2.2505
R37218 PAD.n7644 PAD.n7643 2.2505
R37219 PAD.n7640 PAD.n7639 2.2505
R37220 PAD.n7637 PAD.n7636 2.2505
R37221 PAD.n7629 PAD.n7130 2.2505
R37222 PAD.n7632 PAD.n7631 2.2505
R37223 PAD.n7628 PAD.n7627 2.2505
R37224 PAD.n7625 PAD.n7624 2.2505
R37225 PAD.n7617 PAD.n7132 2.2505
R37226 PAD.n7620 PAD.n7619 2.2505
R37227 PAD.n7616 PAD.n7615 2.2505
R37228 PAD.n7613 PAD.n7612 2.2505
R37229 PAD.n7605 PAD.n7134 2.2505
R37230 PAD.n7608 PAD.n7607 2.2505
R37231 PAD.n7604 PAD.n7603 2.2505
R37232 PAD.n7601 PAD.n7600 2.2505
R37233 PAD.n7593 PAD.n7136 2.2505
R37234 PAD.n7596 PAD.n7595 2.2505
R37235 PAD.n7592 PAD.n7591 2.2505
R37236 PAD.n7589 PAD.n7588 2.2505
R37237 PAD.n7581 PAD.n7138 2.2505
R37238 PAD.n7584 PAD.n7583 2.2505
R37239 PAD.n7580 PAD.n7579 2.2505
R37240 PAD.n7577 PAD.n7576 2.2505
R37241 PAD.n7569 PAD.n7140 2.2505
R37242 PAD.n7572 PAD.n7571 2.2505
R37243 PAD.n7568 PAD.n7567 2.2505
R37244 PAD.n7565 PAD.n7564 2.2505
R37245 PAD.n7557 PAD.n7142 2.2505
R37246 PAD.n7560 PAD.n7559 2.2505
R37247 PAD.n7556 PAD.n7555 2.2505
R37248 PAD.n7553 PAD.n7552 2.2505
R37249 PAD.n7545 PAD.n7144 2.2505
R37250 PAD.n7548 PAD.n7547 2.2505
R37251 PAD.n7544 PAD.n7543 2.2505
R37252 PAD.n7541 PAD.n7540 2.2505
R37253 PAD.n7533 PAD.n7146 2.2505
R37254 PAD.n7536 PAD.n7535 2.2505
R37255 PAD.n7532 PAD.n7531 2.2505
R37256 PAD.n7532 PAD.n7147 2.2505
R37257 PAD.n7537 PAD.n7536 2.2505
R37258 PAD.n7538 PAD.n7146 2.2505
R37259 PAD.n7540 PAD.n7539 2.2505
R37260 PAD.n7544 PAD.n7145 2.2505
R37261 PAD.n7549 PAD.n7548 2.2505
R37262 PAD.n7550 PAD.n7144 2.2505
R37263 PAD.n7552 PAD.n7551 2.2505
R37264 PAD.n7556 PAD.n7143 2.2505
R37265 PAD.n7561 PAD.n7560 2.2505
R37266 PAD.n7562 PAD.n7142 2.2505
R37267 PAD.n7564 PAD.n7563 2.2505
R37268 PAD.n7568 PAD.n7141 2.2505
R37269 PAD.n7573 PAD.n7572 2.2505
R37270 PAD.n7574 PAD.n7140 2.2505
R37271 PAD.n7576 PAD.n7575 2.2505
R37272 PAD.n7580 PAD.n7139 2.2505
R37273 PAD.n7585 PAD.n7584 2.2505
R37274 PAD.n7586 PAD.n7138 2.2505
R37275 PAD.n7588 PAD.n7587 2.2505
R37276 PAD.n7592 PAD.n7137 2.2505
R37277 PAD.n7597 PAD.n7596 2.2505
R37278 PAD.n7598 PAD.n7136 2.2505
R37279 PAD.n7600 PAD.n7599 2.2505
R37280 PAD.n7604 PAD.n7135 2.2505
R37281 PAD.n7609 PAD.n7608 2.2505
R37282 PAD.n7610 PAD.n7134 2.2505
R37283 PAD.n7612 PAD.n7611 2.2505
R37284 PAD.n7616 PAD.n7133 2.2505
R37285 PAD.n7621 PAD.n7620 2.2505
R37286 PAD.n7622 PAD.n7132 2.2505
R37287 PAD.n7624 PAD.n7623 2.2505
R37288 PAD.n7628 PAD.n7131 2.2505
R37289 PAD.n7633 PAD.n7632 2.2505
R37290 PAD.n7634 PAD.n7130 2.2505
R37291 PAD.n7636 PAD.n7635 2.2505
R37292 PAD.n7640 PAD.n7129 2.2505
R37293 PAD.n7645 PAD.n7644 2.2505
R37294 PAD.n7646 PAD.n7128 2.2505
R37295 PAD.n7648 PAD.n7647 2.2505
R37296 PAD.n7652 PAD.n7127 2.2505
R37297 PAD.n7657 PAD.n7656 2.2505
R37298 PAD.n7658 PAD.n7126 2.2505
R37299 PAD.n7660 PAD.n7659 2.2505
R37300 PAD.n7664 PAD.n7125 2.2505
R37301 PAD.n7669 PAD.n7668 2.2505
R37302 PAD.n7670 PAD.n7124 2.2505
R37303 PAD.n7672 PAD.n7671 2.2505
R37304 PAD.n7676 PAD.n7123 2.2505
R37305 PAD.n7681 PAD.n7680 2.2505
R37306 PAD.n7682 PAD.n7122 2.2505
R37307 PAD.n7684 PAD.n7683 2.2505
R37308 PAD.n7688 PAD.n7121 2.2505
R37309 PAD.n7693 PAD.n7692 2.2505
R37310 PAD.n7694 PAD.n7120 2.2505
R37311 PAD.n7696 PAD.n7695 2.2505
R37312 PAD.n7700 PAD.n7119 2.2505
R37313 PAD.n7705 PAD.n7704 2.2505
R37314 PAD.n7706 PAD.n7118 2.2505
R37315 PAD.n7708 PAD.n7707 2.2505
R37316 PAD.n7712 PAD.n7117 2.2505
R37317 PAD.n7717 PAD.n7716 2.2505
R37318 PAD.n7718 PAD.n7116 2.2505
R37319 PAD.n7720 PAD.n7719 2.2505
R37320 PAD.n7724 PAD.n7115 2.2505
R37321 PAD.n7729 PAD.n7728 2.2505
R37322 PAD.n7730 PAD.n7114 2.2505
R37323 PAD.n7732 PAD.n7731 2.2505
R37324 PAD.n7736 PAD.n7113 2.2505
R37325 PAD.n7741 PAD.n7740 2.2505
R37326 PAD.n7742 PAD.n7112 2.2505
R37327 PAD.n7744 PAD.n7743 2.2505
R37328 PAD.n7748 PAD.n7111 2.2505
R37329 PAD.n7753 PAD.n7752 2.2505
R37330 PAD.n7754 PAD.n7110 2.2505
R37331 PAD.n7756 PAD.n7755 2.2505
R37332 PAD.n7760 PAD.n7109 2.2505
R37333 PAD.n7765 PAD.n7764 2.2505
R37334 PAD.n7766 PAD.n7108 2.2505
R37335 PAD.n7768 PAD.n7767 2.2505
R37336 PAD.n7772 PAD.n7107 2.2505
R37337 PAD.n7776 PAD.n7775 2.2505
R37338 PAD.n7777 PAD.n7106 2.2505
R37339 PAD.n7779 PAD.n7778 2.2505
R37340 PAD.n7050 PAD.n6719 2.2505
R37341 PAD.n7049 PAD.n7048 2.2505
R37342 PAD.n7046 PAD.n6720 2.2505
R37343 PAD.n7044 PAD.n7043 2.2505
R37344 PAD.n7036 PAD.n6723 2.2505
R37345 PAD.n7039 PAD.n7038 2.2505
R37346 PAD.n7034 PAD.n6726 2.2505
R37347 PAD.n7032 PAD.n7031 2.2505
R37348 PAD.n7024 PAD.n6728 2.2505
R37349 PAD.n7027 PAD.n7026 2.2505
R37350 PAD.n7022 PAD.n6730 2.2505
R37351 PAD.n7020 PAD.n7019 2.2505
R37352 PAD.n7012 PAD.n6732 2.2505
R37353 PAD.n7015 PAD.n7014 2.2505
R37354 PAD.n7010 PAD.n6734 2.2505
R37355 PAD.n7008 PAD.n7007 2.2505
R37356 PAD.n7000 PAD.n6736 2.2505
R37357 PAD.n7003 PAD.n7002 2.2505
R37358 PAD.n6998 PAD.n6738 2.2505
R37359 PAD.n6996 PAD.n6995 2.2505
R37360 PAD.n6988 PAD.n6740 2.2505
R37361 PAD.n6991 PAD.n6990 2.2505
R37362 PAD.n6986 PAD.n6742 2.2505
R37363 PAD.n6984 PAD.n6983 2.2505
R37364 PAD.n6976 PAD.n6744 2.2505
R37365 PAD.n6979 PAD.n6978 2.2505
R37366 PAD.n6974 PAD.n6746 2.2505
R37367 PAD.n6972 PAD.n6971 2.2505
R37368 PAD.n6964 PAD.n6748 2.2505
R37369 PAD.n6967 PAD.n6966 2.2505
R37370 PAD.n6962 PAD.n6750 2.2505
R37371 PAD.n6960 PAD.n6959 2.2505
R37372 PAD.n6952 PAD.n6752 2.2505
R37373 PAD.n6955 PAD.n6954 2.2505
R37374 PAD.n6950 PAD.n6754 2.2505
R37375 PAD.n6948 PAD.n6947 2.2505
R37376 PAD.n6940 PAD.n6756 2.2505
R37377 PAD.n6943 PAD.n6942 2.2505
R37378 PAD.n6938 PAD.n6758 2.2505
R37379 PAD.n6936 PAD.n6935 2.2505
R37380 PAD.n6928 PAD.n6760 2.2505
R37381 PAD.n6931 PAD.n6930 2.2505
R37382 PAD.n6926 PAD.n6762 2.2505
R37383 PAD.n6924 PAD.n6923 2.2505
R37384 PAD.n6916 PAD.n6764 2.2505
R37385 PAD.n6919 PAD.n6918 2.2505
R37386 PAD.n6914 PAD.n6766 2.2505
R37387 PAD.n6912 PAD.n6911 2.2505
R37388 PAD.n6904 PAD.n6768 2.2505
R37389 PAD.n6907 PAD.n6906 2.2505
R37390 PAD.n6902 PAD.n6770 2.2505
R37391 PAD.n6900 PAD.n6899 2.2505
R37392 PAD.n6892 PAD.n6772 2.2505
R37393 PAD.n6895 PAD.n6894 2.2505
R37394 PAD.n6890 PAD.n6774 2.2505
R37395 PAD.n6888 PAD.n6887 2.2505
R37396 PAD.n6880 PAD.n6776 2.2505
R37397 PAD.n6883 PAD.n6882 2.2505
R37398 PAD.n6878 PAD.n6778 2.2505
R37399 PAD.n6876 PAD.n6875 2.2505
R37400 PAD.n6868 PAD.n6780 2.2505
R37401 PAD.n6871 PAD.n6870 2.2505
R37402 PAD.n6866 PAD.n6782 2.2505
R37403 PAD.n6864 PAD.n6863 2.2505
R37404 PAD.n6856 PAD.n6784 2.2505
R37405 PAD.n6859 PAD.n6858 2.2505
R37406 PAD.n6854 PAD.n6786 2.2505
R37407 PAD.n6852 PAD.n6851 2.2505
R37408 PAD.n6844 PAD.n6788 2.2505
R37409 PAD.n6847 PAD.n6846 2.2505
R37410 PAD.n6842 PAD.n6790 2.2505
R37411 PAD.n6840 PAD.n6839 2.2505
R37412 PAD.n6832 PAD.n6792 2.2505
R37413 PAD.n6835 PAD.n6834 2.2505
R37414 PAD.n6830 PAD.n6794 2.2505
R37415 PAD.n6828 PAD.n6827 2.2505
R37416 PAD.n6820 PAD.n6796 2.2505
R37417 PAD.n6823 PAD.n6822 2.2505
R37418 PAD.n6818 PAD.n6798 2.2505
R37419 PAD.n6816 PAD.n6815 2.2505
R37420 PAD.n6808 PAD.n6800 2.2505
R37421 PAD.n6811 PAD.n6810 2.2505
R37422 PAD.n6806 PAD.n6802 2.2505
R37423 PAD.n6804 PAD.n6803 2.2505
R37424 PAD.n6803 PAD.n6705 2.2505
R37425 PAD.n6802 PAD.n6801 2.2505
R37426 PAD.n6812 PAD.n6811 2.2505
R37427 PAD.n6813 PAD.n6800 2.2505
R37428 PAD.n6815 PAD.n6814 2.2505
R37429 PAD.n6798 PAD.n6797 2.2505
R37430 PAD.n6824 PAD.n6823 2.2505
R37431 PAD.n6825 PAD.n6796 2.2505
R37432 PAD.n6827 PAD.n6826 2.2505
R37433 PAD.n6794 PAD.n6793 2.2505
R37434 PAD.n6836 PAD.n6835 2.2505
R37435 PAD.n6837 PAD.n6792 2.2505
R37436 PAD.n6839 PAD.n6838 2.2505
R37437 PAD.n6790 PAD.n6789 2.2505
R37438 PAD.n6848 PAD.n6847 2.2505
R37439 PAD.n6849 PAD.n6788 2.2505
R37440 PAD.n6851 PAD.n6850 2.2505
R37441 PAD.n6786 PAD.n6785 2.2505
R37442 PAD.n6860 PAD.n6859 2.2505
R37443 PAD.n6861 PAD.n6784 2.2505
R37444 PAD.n6863 PAD.n6862 2.2505
R37445 PAD.n6782 PAD.n6781 2.2505
R37446 PAD.n6872 PAD.n6871 2.2505
R37447 PAD.n6873 PAD.n6780 2.2505
R37448 PAD.n6875 PAD.n6874 2.2505
R37449 PAD.n6778 PAD.n6777 2.2505
R37450 PAD.n6884 PAD.n6883 2.2505
R37451 PAD.n6885 PAD.n6776 2.2505
R37452 PAD.n6887 PAD.n6886 2.2505
R37453 PAD.n6774 PAD.n6773 2.2505
R37454 PAD.n6896 PAD.n6895 2.2505
R37455 PAD.n6897 PAD.n6772 2.2505
R37456 PAD.n6899 PAD.n6898 2.2505
R37457 PAD.n6770 PAD.n6769 2.2505
R37458 PAD.n6908 PAD.n6907 2.2505
R37459 PAD.n6909 PAD.n6768 2.2505
R37460 PAD.n6911 PAD.n6910 2.2505
R37461 PAD.n6766 PAD.n6765 2.2505
R37462 PAD.n6920 PAD.n6919 2.2505
R37463 PAD.n6921 PAD.n6764 2.2505
R37464 PAD.n6923 PAD.n6922 2.2505
R37465 PAD.n6762 PAD.n6761 2.2505
R37466 PAD.n6932 PAD.n6931 2.2505
R37467 PAD.n6933 PAD.n6760 2.2505
R37468 PAD.n6935 PAD.n6934 2.2505
R37469 PAD.n6758 PAD.n6757 2.2505
R37470 PAD.n6944 PAD.n6943 2.2505
R37471 PAD.n6945 PAD.n6756 2.2505
R37472 PAD.n6947 PAD.n6946 2.2505
R37473 PAD.n6754 PAD.n6753 2.2505
R37474 PAD.n6956 PAD.n6955 2.2505
R37475 PAD.n6957 PAD.n6752 2.2505
R37476 PAD.n6959 PAD.n6958 2.2505
R37477 PAD.n6750 PAD.n6749 2.2505
R37478 PAD.n6968 PAD.n6967 2.2505
R37479 PAD.n6969 PAD.n6748 2.2505
R37480 PAD.n6971 PAD.n6970 2.2505
R37481 PAD.n6746 PAD.n6745 2.2505
R37482 PAD.n6980 PAD.n6979 2.2505
R37483 PAD.n6981 PAD.n6744 2.2505
R37484 PAD.n6983 PAD.n6982 2.2505
R37485 PAD.n6742 PAD.n6741 2.2505
R37486 PAD.n6992 PAD.n6991 2.2505
R37487 PAD.n6993 PAD.n6740 2.2505
R37488 PAD.n6995 PAD.n6994 2.2505
R37489 PAD.n6738 PAD.n6737 2.2505
R37490 PAD.n7004 PAD.n7003 2.2505
R37491 PAD.n7005 PAD.n6736 2.2505
R37492 PAD.n7007 PAD.n7006 2.2505
R37493 PAD.n6734 PAD.n6733 2.2505
R37494 PAD.n7016 PAD.n7015 2.2505
R37495 PAD.n7017 PAD.n6732 2.2505
R37496 PAD.n7019 PAD.n7018 2.2505
R37497 PAD.n6730 PAD.n6729 2.2505
R37498 PAD.n7028 PAD.n7027 2.2505
R37499 PAD.n7029 PAD.n6728 2.2505
R37500 PAD.n7031 PAD.n7030 2.2505
R37501 PAD.n6726 PAD.n6725 2.2505
R37502 PAD.n7040 PAD.n7039 2.2505
R37503 PAD.n7041 PAD.n6723 2.2505
R37504 PAD.n7043 PAD.n7042 2.2505
R37505 PAD.n6724 PAD.n6720 2.2505
R37506 PAD.n7049 PAD.n6718 2.2505
R37507 PAD.n7051 PAD.n7050 2.2505
R37508 PAD.n5892 PAD.n5891 2.2505
R37509 PAD.n5890 PAD.n5602 2.2505
R37510 PAD.n5605 PAD.n5604 2.2505
R37511 PAD.n5886 PAD.n5885 2.2505
R37512 PAD.n5883 PAD.n5882 2.2505
R37513 PAD.n5881 PAD.n5610 2.2505
R37514 PAD.n5608 PAD.n5607 2.2505
R37515 PAD.n5877 PAD.n5876 2.2505
R37516 PAD.n5874 PAD.n5873 2.2505
R37517 PAD.n5872 PAD.n5615 2.2505
R37518 PAD.n5613 PAD.n5612 2.2505
R37519 PAD.n5868 PAD.n5867 2.2505
R37520 PAD.n5865 PAD.n5864 2.2505
R37521 PAD.n5863 PAD.n5620 2.2505
R37522 PAD.n5618 PAD.n5617 2.2505
R37523 PAD.n5859 PAD.n5858 2.2505
R37524 PAD.n5856 PAD.n5855 2.2505
R37525 PAD.n5854 PAD.n5625 2.2505
R37526 PAD.n5623 PAD.n5622 2.2505
R37527 PAD.n5850 PAD.n5849 2.2505
R37528 PAD.n5847 PAD.n5846 2.2505
R37529 PAD.n5845 PAD.n5630 2.2505
R37530 PAD.n5628 PAD.n5627 2.2505
R37531 PAD.n5841 PAD.n5840 2.2505
R37532 PAD.n5838 PAD.n5837 2.2505
R37533 PAD.n5836 PAD.n5635 2.2505
R37534 PAD.n5633 PAD.n5632 2.2505
R37535 PAD.n5832 PAD.n5831 2.2505
R37536 PAD.n5829 PAD.n5828 2.2505
R37537 PAD.n5827 PAD.n5640 2.2505
R37538 PAD.n5638 PAD.n5637 2.2505
R37539 PAD.n5823 PAD.n5822 2.2505
R37540 PAD.n5820 PAD.n5819 2.2505
R37541 PAD.n5818 PAD.n5645 2.2505
R37542 PAD.n5643 PAD.n5642 2.2505
R37543 PAD.n5814 PAD.n5813 2.2505
R37544 PAD.n5811 PAD.n5810 2.2505
R37545 PAD.n5809 PAD.n5650 2.2505
R37546 PAD.n5648 PAD.n5647 2.2505
R37547 PAD.n5805 PAD.n5804 2.2505
R37548 PAD.n5802 PAD.n5801 2.2505
R37549 PAD.n5800 PAD.n5655 2.2505
R37550 PAD.n5653 PAD.n5652 2.2505
R37551 PAD.n5796 PAD.n5795 2.2505
R37552 PAD.n5793 PAD.n5792 2.2505
R37553 PAD.n5791 PAD.n5660 2.2505
R37554 PAD.n5658 PAD.n5657 2.2505
R37555 PAD.n5787 PAD.n5786 2.2505
R37556 PAD.n5784 PAD.n5783 2.2505
R37557 PAD.n5782 PAD.n5665 2.2505
R37558 PAD.n5663 PAD.n5662 2.2505
R37559 PAD.n5778 PAD.n5777 2.2505
R37560 PAD.n5775 PAD.n5774 2.2505
R37561 PAD.n5773 PAD.n5670 2.2505
R37562 PAD.n5668 PAD.n5667 2.2505
R37563 PAD.n5769 PAD.n5768 2.2505
R37564 PAD.n5766 PAD.n5765 2.2505
R37565 PAD.n5764 PAD.n5675 2.2505
R37566 PAD.n5673 PAD.n5672 2.2505
R37567 PAD.n5760 PAD.n5759 2.2505
R37568 PAD.n5757 PAD.n5756 2.2505
R37569 PAD.n5755 PAD.n5680 2.2505
R37570 PAD.n5678 PAD.n5677 2.2505
R37571 PAD.n5751 PAD.n5750 2.2505
R37572 PAD.n5748 PAD.n5747 2.2505
R37573 PAD.n5746 PAD.n5685 2.2505
R37574 PAD.n5683 PAD.n5682 2.2505
R37575 PAD.n5742 PAD.n5741 2.2505
R37576 PAD.n5739 PAD.n5738 2.2505
R37577 PAD.n5737 PAD.n5690 2.2505
R37578 PAD.n5688 PAD.n5687 2.2505
R37579 PAD.n5733 PAD.n5732 2.2505
R37580 PAD.n5730 PAD.n5729 2.2505
R37581 PAD.n5728 PAD.n5695 2.2505
R37582 PAD.n5693 PAD.n5692 2.2505
R37583 PAD.n5724 PAD.n5723 2.2505
R37584 PAD.n5721 PAD.n5720 2.2505
R37585 PAD.n5719 PAD.n5700 2.2505
R37586 PAD.n5698 PAD.n5697 2.2505
R37587 PAD.n5715 PAD.n5714 2.2505
R37588 PAD.n5712 PAD.n5711 2.2505
R37589 PAD.n5710 PAD.n5707 2.2505
R37590 PAD.n5705 PAD.n5704 2.2505
R37591 PAD.n5703 PAD.n5702 2.2505
R37592 PAD.n5703 PAD.n5557 2.2505
R37593 PAD.n5708 PAD.n5704 2.2505
R37594 PAD.n5710 PAD.n5709 2.2505
R37595 PAD.n5711 PAD.n5701 2.2505
R37596 PAD.n5716 PAD.n5715 2.2505
R37597 PAD.n5717 PAD.n5697 2.2505
R37598 PAD.n5719 PAD.n5718 2.2505
R37599 PAD.n5720 PAD.n5696 2.2505
R37600 PAD.n5725 PAD.n5724 2.2505
R37601 PAD.n5726 PAD.n5692 2.2505
R37602 PAD.n5728 PAD.n5727 2.2505
R37603 PAD.n5729 PAD.n5691 2.2505
R37604 PAD.n5734 PAD.n5733 2.2505
R37605 PAD.n5735 PAD.n5687 2.2505
R37606 PAD.n5737 PAD.n5736 2.2505
R37607 PAD.n5738 PAD.n5686 2.2505
R37608 PAD.n5743 PAD.n5742 2.2505
R37609 PAD.n5744 PAD.n5682 2.2505
R37610 PAD.n5746 PAD.n5745 2.2505
R37611 PAD.n5747 PAD.n5681 2.2505
R37612 PAD.n5752 PAD.n5751 2.2505
R37613 PAD.n5753 PAD.n5677 2.2505
R37614 PAD.n5755 PAD.n5754 2.2505
R37615 PAD.n5756 PAD.n5676 2.2505
R37616 PAD.n5761 PAD.n5760 2.2505
R37617 PAD.n5762 PAD.n5672 2.2505
R37618 PAD.n5764 PAD.n5763 2.2505
R37619 PAD.n5765 PAD.n5671 2.2505
R37620 PAD.n5770 PAD.n5769 2.2505
R37621 PAD.n5771 PAD.n5667 2.2505
R37622 PAD.n5773 PAD.n5772 2.2505
R37623 PAD.n5774 PAD.n5666 2.2505
R37624 PAD.n5779 PAD.n5778 2.2505
R37625 PAD.n5780 PAD.n5662 2.2505
R37626 PAD.n5782 PAD.n5781 2.2505
R37627 PAD.n5783 PAD.n5661 2.2505
R37628 PAD.n5788 PAD.n5787 2.2505
R37629 PAD.n5789 PAD.n5657 2.2505
R37630 PAD.n5791 PAD.n5790 2.2505
R37631 PAD.n5792 PAD.n5656 2.2505
R37632 PAD.n5797 PAD.n5796 2.2505
R37633 PAD.n5798 PAD.n5652 2.2505
R37634 PAD.n5800 PAD.n5799 2.2505
R37635 PAD.n5801 PAD.n5651 2.2505
R37636 PAD.n5806 PAD.n5805 2.2505
R37637 PAD.n5807 PAD.n5647 2.2505
R37638 PAD.n5809 PAD.n5808 2.2505
R37639 PAD.n5810 PAD.n5646 2.2505
R37640 PAD.n5815 PAD.n5814 2.2505
R37641 PAD.n5816 PAD.n5642 2.2505
R37642 PAD.n5818 PAD.n5817 2.2505
R37643 PAD.n5819 PAD.n5641 2.2505
R37644 PAD.n5824 PAD.n5823 2.2505
R37645 PAD.n5825 PAD.n5637 2.2505
R37646 PAD.n5827 PAD.n5826 2.2505
R37647 PAD.n5828 PAD.n5636 2.2505
R37648 PAD.n5833 PAD.n5832 2.2505
R37649 PAD.n5834 PAD.n5632 2.2505
R37650 PAD.n5836 PAD.n5835 2.2505
R37651 PAD.n5837 PAD.n5631 2.2505
R37652 PAD.n5842 PAD.n5841 2.2505
R37653 PAD.n5843 PAD.n5627 2.2505
R37654 PAD.n5845 PAD.n5844 2.2505
R37655 PAD.n5846 PAD.n5626 2.2505
R37656 PAD.n5851 PAD.n5850 2.2505
R37657 PAD.n5852 PAD.n5622 2.2505
R37658 PAD.n5854 PAD.n5853 2.2505
R37659 PAD.n5855 PAD.n5621 2.2505
R37660 PAD.n5860 PAD.n5859 2.2505
R37661 PAD.n5861 PAD.n5617 2.2505
R37662 PAD.n5863 PAD.n5862 2.2505
R37663 PAD.n5864 PAD.n5616 2.2505
R37664 PAD.n5869 PAD.n5868 2.2505
R37665 PAD.n5870 PAD.n5612 2.2505
R37666 PAD.n5872 PAD.n5871 2.2505
R37667 PAD.n5873 PAD.n5611 2.2505
R37668 PAD.n5878 PAD.n5877 2.2505
R37669 PAD.n5879 PAD.n5607 2.2505
R37670 PAD.n5881 PAD.n5880 2.2505
R37671 PAD.n5882 PAD.n5606 2.2505
R37672 PAD.n5887 PAD.n5886 2.2505
R37673 PAD.n5888 PAD.n5605 2.2505
R37674 PAD.n5890 PAD.n5889 2.2505
R37675 PAD.n5891 PAD.n5545 2.2505
R37676 PAD.n6687 PAD.n5951 2.2505
R37677 PAD.n6672 PAD.n5950 2.2505
R37678 PAD.n6673 PAD.n6439 2.2505
R37679 PAD.n6675 PAD.n6674 2.2505
R37680 PAD.n6671 PAD.n6438 2.2505
R37681 PAD.n6670 PAD.n6669 2.2505
R37682 PAD.n6667 PAD.n6440 2.2505
R37683 PAD.n6665 PAD.n6663 2.2505
R37684 PAD.n6662 PAD.n6442 2.2505
R37685 PAD.n6661 PAD.n6660 2.2505
R37686 PAD.n6658 PAD.n6443 2.2505
R37687 PAD.n6656 PAD.n6654 2.2505
R37688 PAD.n6653 PAD.n6445 2.2505
R37689 PAD.n6652 PAD.n6651 2.2505
R37690 PAD.n6649 PAD.n6446 2.2505
R37691 PAD.n6647 PAD.n6645 2.2505
R37692 PAD.n6644 PAD.n6448 2.2505
R37693 PAD.n6643 PAD.n6642 2.2505
R37694 PAD.n6640 PAD.n6449 2.2505
R37695 PAD.n6638 PAD.n6636 2.2505
R37696 PAD.n6635 PAD.n6451 2.2505
R37697 PAD.n6634 PAD.n6633 2.2505
R37698 PAD.n6631 PAD.n6452 2.2505
R37699 PAD.n6629 PAD.n6627 2.2505
R37700 PAD.n6626 PAD.n6454 2.2505
R37701 PAD.n6625 PAD.n6624 2.2505
R37702 PAD.n6622 PAD.n6455 2.2505
R37703 PAD.n6620 PAD.n6618 2.2505
R37704 PAD.n6617 PAD.n6457 2.2505
R37705 PAD.n6616 PAD.n6615 2.2505
R37706 PAD.n6613 PAD.n6458 2.2505
R37707 PAD.n6611 PAD.n6609 2.2505
R37708 PAD.n6608 PAD.n6460 2.2505
R37709 PAD.n6607 PAD.n6606 2.2505
R37710 PAD.n6604 PAD.n6461 2.2505
R37711 PAD.n6602 PAD.n6600 2.2505
R37712 PAD.n6599 PAD.n6463 2.2505
R37713 PAD.n6598 PAD.n6597 2.2505
R37714 PAD.n6595 PAD.n6464 2.2505
R37715 PAD.n6593 PAD.n6591 2.2505
R37716 PAD.n6590 PAD.n6466 2.2505
R37717 PAD.n6589 PAD.n6588 2.2505
R37718 PAD.n6586 PAD.n6467 2.2505
R37719 PAD.n6584 PAD.n6582 2.2505
R37720 PAD.n6581 PAD.n6469 2.2505
R37721 PAD.n6580 PAD.n6579 2.2505
R37722 PAD.n6577 PAD.n6470 2.2505
R37723 PAD.n6575 PAD.n6573 2.2505
R37724 PAD.n6572 PAD.n6472 2.2505
R37725 PAD.n6571 PAD.n6570 2.2505
R37726 PAD.n6568 PAD.n6473 2.2505
R37727 PAD.n6566 PAD.n6564 2.2505
R37728 PAD.n6563 PAD.n6475 2.2505
R37729 PAD.n6562 PAD.n6561 2.2505
R37730 PAD.n6559 PAD.n6476 2.2505
R37731 PAD.n6557 PAD.n6555 2.2505
R37732 PAD.n6554 PAD.n6478 2.2505
R37733 PAD.n6553 PAD.n6552 2.2505
R37734 PAD.n6550 PAD.n6479 2.2505
R37735 PAD.n6548 PAD.n6546 2.2505
R37736 PAD.n6545 PAD.n6481 2.2505
R37737 PAD.n6544 PAD.n6543 2.2505
R37738 PAD.n6541 PAD.n6482 2.2505
R37739 PAD.n6539 PAD.n6537 2.2505
R37740 PAD.n6536 PAD.n6484 2.2505
R37741 PAD.n6535 PAD.n6534 2.2505
R37742 PAD.n6532 PAD.n6485 2.2505
R37743 PAD.n6530 PAD.n6528 2.2505
R37744 PAD.n6527 PAD.n6487 2.2505
R37745 PAD.n6526 PAD.n6525 2.2505
R37746 PAD.n6523 PAD.n6488 2.2505
R37747 PAD.n6521 PAD.n6519 2.2505
R37748 PAD.n6518 PAD.n6490 2.2505
R37749 PAD.n6517 PAD.n6516 2.2505
R37750 PAD.n6514 PAD.n6491 2.2505
R37751 PAD.n6512 PAD.n6510 2.2505
R37752 PAD.n6509 PAD.n6493 2.2505
R37753 PAD.n6508 PAD.n6507 2.2505
R37754 PAD.n6505 PAD.n6494 2.2505
R37755 PAD.n6503 PAD.n6501 2.2505
R37756 PAD.n6500 PAD.n6496 2.2505
R37757 PAD.n6499 PAD.n6498 2.2505
R37758 PAD.n5900 PAD.n5898 2.2505
R37759 PAD.n6692 PAD.n6691 2.2505
R37760 PAD.n75 PAD.n26 2.2505
R37761 PAD.n363 PAD.n362 2.2505
R37762 PAD.n361 PAD.n76 2.2505
R37763 PAD.n360 PAD.n359 2.2505
R37764 PAD.n355 PAD.n77 2.2505
R37765 PAD.n351 PAD.n350 2.2505
R37766 PAD.n349 PAD.n78 2.2505
R37767 PAD.n348 PAD.n347 2.2505
R37768 PAD.n343 PAD.n79 2.2505
R37769 PAD.n339 PAD.n338 2.2505
R37770 PAD.n337 PAD.n80 2.2505
R37771 PAD.n336 PAD.n335 2.2505
R37772 PAD.n331 PAD.n81 2.2505
R37773 PAD.n327 PAD.n326 2.2505
R37774 PAD.n325 PAD.n82 2.2505
R37775 PAD.n324 PAD.n323 2.2505
R37776 PAD.n319 PAD.n83 2.2505
R37777 PAD.n315 PAD.n314 2.2505
R37778 PAD.n313 PAD.n84 2.2505
R37779 PAD.n312 PAD.n311 2.2505
R37780 PAD.n307 PAD.n85 2.2505
R37781 PAD.n303 PAD.n302 2.2505
R37782 PAD.n301 PAD.n86 2.2505
R37783 PAD.n300 PAD.n299 2.2505
R37784 PAD.n295 PAD.n87 2.2505
R37785 PAD.n291 PAD.n290 2.2505
R37786 PAD.n289 PAD.n88 2.2505
R37787 PAD.n288 PAD.n287 2.2505
R37788 PAD.n283 PAD.n89 2.2505
R37789 PAD.n279 PAD.n278 2.2505
R37790 PAD.n277 PAD.n90 2.2505
R37791 PAD.n276 PAD.n275 2.2505
R37792 PAD.n271 PAD.n91 2.2505
R37793 PAD.n267 PAD.n266 2.2505
R37794 PAD.n265 PAD.n92 2.2505
R37795 PAD.n264 PAD.n263 2.2505
R37796 PAD.n259 PAD.n93 2.2505
R37797 PAD.n255 PAD.n254 2.2505
R37798 PAD.n253 PAD.n94 2.2505
R37799 PAD.n252 PAD.n251 2.2505
R37800 PAD.n247 PAD.n95 2.2505
R37801 PAD.n243 PAD.n242 2.2505
R37802 PAD.n241 PAD.n96 2.2505
R37803 PAD.n240 PAD.n239 2.2505
R37804 PAD.n235 PAD.n97 2.2505
R37805 PAD.n231 PAD.n230 2.2505
R37806 PAD.n229 PAD.n98 2.2505
R37807 PAD.n228 PAD.n227 2.2505
R37808 PAD.n223 PAD.n99 2.2505
R37809 PAD.n219 PAD.n218 2.2505
R37810 PAD.n217 PAD.n100 2.2505
R37811 PAD.n216 PAD.n215 2.2505
R37812 PAD.n211 PAD.n101 2.2505
R37813 PAD.n207 PAD.n206 2.2505
R37814 PAD.n205 PAD.n102 2.2505
R37815 PAD.n204 PAD.n203 2.2505
R37816 PAD.n199 PAD.n103 2.2505
R37817 PAD.n195 PAD.n194 2.2505
R37818 PAD.n193 PAD.n104 2.2505
R37819 PAD.n192 PAD.n191 2.2505
R37820 PAD.n187 PAD.n105 2.2505
R37821 PAD.n183 PAD.n182 2.2505
R37822 PAD.n181 PAD.n106 2.2505
R37823 PAD.n180 PAD.n179 2.2505
R37824 PAD.n175 PAD.n107 2.2505
R37825 PAD.n171 PAD.n170 2.2505
R37826 PAD.n169 PAD.n108 2.2505
R37827 PAD.n168 PAD.n167 2.2505
R37828 PAD.n163 PAD.n109 2.2505
R37829 PAD.n159 PAD.n158 2.2505
R37830 PAD.n157 PAD.n110 2.2505
R37831 PAD.n156 PAD.n155 2.2505
R37832 PAD.n151 PAD.n111 2.2505
R37833 PAD.n147 PAD.n146 2.2505
R37834 PAD.n145 PAD.n112 2.2505
R37835 PAD.n144 PAD.n143 2.2505
R37836 PAD.n139 PAD.n113 2.2505
R37837 PAD.n135 PAD.n134 2.2505
R37838 PAD.n133 PAD.n114 2.2505
R37839 PAD.n132 PAD.n131 2.2505
R37840 PAD.n127 PAD.n115 2.2505
R37841 PAD.n123 PAD.n122 2.2505
R37842 PAD.n121 PAD.n118 2.2505
R37843 PAD.n120 PAD.n119 2.2505
R37844 PAD.n119 PAD.n74 2.2505
R37845 PAD.n118 PAD.n117 2.2505
R37846 PAD.n124 PAD.n123 2.2505
R37847 PAD.n127 PAD.n126 2.2505
R37848 PAD.n131 PAD.n130 2.2505
R37849 PAD.n128 PAD.n114 2.2505
R37850 PAD.n136 PAD.n135 2.2505
R37851 PAD.n139 PAD.n138 2.2505
R37852 PAD.n143 PAD.n142 2.2505
R37853 PAD.n140 PAD.n112 2.2505
R37854 PAD.n148 PAD.n147 2.2505
R37855 PAD.n151 PAD.n150 2.2505
R37856 PAD.n155 PAD.n154 2.2505
R37857 PAD.n152 PAD.n110 2.2505
R37858 PAD.n160 PAD.n159 2.2505
R37859 PAD.n163 PAD.n162 2.2505
R37860 PAD.n167 PAD.n166 2.2505
R37861 PAD.n164 PAD.n108 2.2505
R37862 PAD.n172 PAD.n171 2.2505
R37863 PAD.n175 PAD.n174 2.2505
R37864 PAD.n179 PAD.n178 2.2505
R37865 PAD.n176 PAD.n106 2.2505
R37866 PAD.n184 PAD.n183 2.2505
R37867 PAD.n187 PAD.n186 2.2505
R37868 PAD.n191 PAD.n190 2.2505
R37869 PAD.n188 PAD.n104 2.2505
R37870 PAD.n196 PAD.n195 2.2505
R37871 PAD.n199 PAD.n198 2.2505
R37872 PAD.n203 PAD.n202 2.2505
R37873 PAD.n200 PAD.n102 2.2505
R37874 PAD.n208 PAD.n207 2.2505
R37875 PAD.n211 PAD.n210 2.2505
R37876 PAD.n215 PAD.n214 2.2505
R37877 PAD.n212 PAD.n100 2.2505
R37878 PAD.n220 PAD.n219 2.2505
R37879 PAD.n223 PAD.n222 2.2505
R37880 PAD.n227 PAD.n226 2.2505
R37881 PAD.n224 PAD.n98 2.2505
R37882 PAD.n232 PAD.n231 2.2505
R37883 PAD.n235 PAD.n234 2.2505
R37884 PAD.n239 PAD.n238 2.2505
R37885 PAD.n236 PAD.n96 2.2505
R37886 PAD.n244 PAD.n243 2.2505
R37887 PAD.n247 PAD.n246 2.2505
R37888 PAD.n251 PAD.n250 2.2505
R37889 PAD.n248 PAD.n94 2.2505
R37890 PAD.n256 PAD.n255 2.2505
R37891 PAD.n259 PAD.n258 2.2505
R37892 PAD.n263 PAD.n262 2.2505
R37893 PAD.n260 PAD.n92 2.2505
R37894 PAD.n268 PAD.n267 2.2505
R37895 PAD.n271 PAD.n270 2.2505
R37896 PAD.n275 PAD.n274 2.2505
R37897 PAD.n272 PAD.n90 2.2505
R37898 PAD.n280 PAD.n279 2.2505
R37899 PAD.n283 PAD.n282 2.2505
R37900 PAD.n287 PAD.n286 2.2505
R37901 PAD.n284 PAD.n88 2.2505
R37902 PAD.n292 PAD.n291 2.2505
R37903 PAD.n295 PAD.n294 2.2505
R37904 PAD.n299 PAD.n298 2.2505
R37905 PAD.n296 PAD.n86 2.2505
R37906 PAD.n304 PAD.n303 2.2505
R37907 PAD.n307 PAD.n306 2.2505
R37908 PAD.n311 PAD.n310 2.2505
R37909 PAD.n308 PAD.n84 2.2505
R37910 PAD.n316 PAD.n315 2.2505
R37911 PAD.n319 PAD.n318 2.2505
R37912 PAD.n323 PAD.n322 2.2505
R37913 PAD.n320 PAD.n82 2.2505
R37914 PAD.n328 PAD.n327 2.2505
R37915 PAD.n331 PAD.n330 2.2505
R37916 PAD.n335 PAD.n334 2.2505
R37917 PAD.n332 PAD.n80 2.2505
R37918 PAD.n340 PAD.n339 2.2505
R37919 PAD.n343 PAD.n342 2.2505
R37920 PAD.n347 PAD.n346 2.2505
R37921 PAD.n344 PAD.n78 2.2505
R37922 PAD.n352 PAD.n351 2.2505
R37923 PAD.n355 PAD.n354 2.2505
R37924 PAD.n359 PAD.n358 2.2505
R37925 PAD.n356 PAD.n76 2.2505
R37926 PAD.n364 PAD.n363 2.2505
R37927 PAD.n366 PAD.n75 2.2505
R37928 PAD.n6381 PAD.n6380 2.2505
R37929 PAD.n6379 PAD.n5977 2.2505
R37930 PAD.n6378 PAD.n5952 2.2505
R37931 PAD.n6685 PAD.n5953 2.2505
R37932 PAD.n5559 PAD.n5558 2.2505
R37933 PAD.n6703 PAD.n6702 2.2505
R37934 PAD.n7799 PAD.n7798 2.2505
R37935 PAD.n7797 PAD.n5556 2.2505
R37936 PAD.n7795 PAD.n7794 2.2505
R37937 PAD.n6708 PAD.n6706 2.2505
R37938 PAD.n7153 PAD.n7152 2.2505
R37939 PAD.n7527 PAD.n7526 2.2505
R37940 PAD.n7525 PAD.n7151 2.2505
R37941 PAD.n7524 PAD.n7523 2.2505
R37942 PAD.n7204 PAD.n7203 2.2505
R37943 PAD.n5202 PAD.n5201 2.2505
R37944 PAD.n7823 PAD.n7822 2.2505
R37945 PAD.n7826 PAD.n7825 2.2505
R37946 PAD.n5188 PAD.n5187 2.2505
R37947 PAD.n8178 PAD.n8177 2.2505
R37948 PAD.n8181 PAD.n8180 2.2505
R37949 PAD.n4837 PAD.n4836 2.2505
R37950 PAD.n8198 PAD.n8197 2.2505
R37951 PAD.n8201 PAD.n8200 2.2505
R37952 PAD.n8202 PAD.n4830 2.2505
R37953 PAD.n8208 PAD.n8207 2.2505
R37954 PAD.n4671 PAD.n4670 2.2505
R37955 PAD.n8413 PAD.n8412 2.2505
R37956 PAD.n8417 PAD.n8416 2.2505
R37957 PAD.n8415 PAD.n4317 2.2505
R37958 PAD.n8433 PAD.n4315 2.2505
R37959 PAD.n8436 PAD.n8435 2.2505
R37960 PAD.n4316 PAD.n3975 2.2505
R37961 PAD.n8457 PAD.n3974 2.2505
R37962 PAD.n8460 PAD.n8459 2.2505
R37963 PAD.n3630 PAD.n3629 2.2505
R37964 PAD.n8483 PAD.n8482 2.2505
R37965 PAD.n8484 PAD.n3285 2.2505
R37966 PAD.n8505 PAD.n3284 2.2505
R37967 PAD.n8509 PAD.n8508 2.2505
R37968 PAD.n2900 PAD.n2899 2.2505
R37969 PAD.n8825 PAD.n8824 2.2505
R37970 PAD.n8827 PAD.n2896 2.2505
R37971 PAD.n8829 PAD.n8828 2.2505
R37972 PAD.n2897 PAD.n2882 2.2505
R37973 PAD.n9132 PAD.n9131 2.2505
R37974 PAD.n2492 PAD.n2491 2.2505
R37975 PAD.n9155 PAD.n9154 2.2505
R37976 PAD.n9158 PAD.n9157 2.2505
R37977 PAD.n2144 PAD.n2143 2.2505
R37978 PAD.n9179 PAD.n9178 2.2505
R37979 PAD.n9182 PAD.n9181 2.2505
R37980 PAD.n2042 PAD.n2041 2.2505
R37981 PAD.n9449 PAD.n9448 2.2505
R37982 PAD.n9451 PAD.n2039 2.2505
R37983 PAD.n9453 PAD.n9452 2.2505
R37984 PAD.n9716 PAD.n9715 2.2505
R37985 PAD.n9717 PAD.n1938 2.2505
R37986 PAD.n9719 PAD.n9718 2.2505
R37987 PAD.n9736 PAD.n9735 2.2505
R37988 PAD.n9737 PAD.n1588 2.2505
R37989 PAD.n9739 PAD.n9738 2.2505
R37990 PAD.n10002 PAD.n10001 2.2505
R37991 PAD.n10003 PAD.n1485 2.2505
R37992 PAD.n10005 PAD.n10004 2.2505
R37993 PAD.n10020 PAD.n10019 2.2505
R37994 PAD.n10021 PAD.n1135 2.2505
R37995 PAD.n10359 PAD.n10358 2.2505
R37996 PAD.n10356 PAD.n1116 2.2505
R37997 PAD.n10376 PAD.n1115 2.2505
R37998 PAD.n10380 PAD.n10379 2.2505
R37999 PAD.n774 PAD.n773 2.2505
R38000 PAD.n10401 PAD.n10400 2.2505
R38001 PAD.n10405 PAD.n10404 2.2505
R38002 PAD.n10403 PAD.n423 2.2505
R38003 PAD.n10704 PAD.n422 2.2505
R38004 PAD.n10708 PAD.n10707 2.2505
R38005 PAD.n28 PAD.n27 2.2505
R38006 PAD.n10731 PAD.n10730 2.2505
R38007 PAD.n10733 PAD.n24 2.2505
R38008 PAD.n11530 PAD.n11529 2.2505
R38009 PAD.n11528 PAD.n25 2.2505
R38010 PAD.n11526 PAD.n11525 2.2505
R38011 PAD.n10737 PAD.n10735 2.2505
R38012 PAD.n11504 PAD.n11503 2.2505
R38013 PAD.n10838 PAD.n10734 2.2505
R38014 PAD.n10840 PAD.n10839 2.2505
R38015 PAD.n10835 PAD.n10834 2.2505
R38016 PAD.n10849 PAD.n10848 2.2505
R38017 PAD.n10850 PAD.n10833 2.2505
R38018 PAD.n10852 PAD.n10851 2.2505
R38019 PAD.n10831 PAD.n10830 2.2505
R38020 PAD.n10861 PAD.n10860 2.2505
R38021 PAD.n10862 PAD.n10829 2.2505
R38022 PAD.n10864 PAD.n10863 2.2505
R38023 PAD.n10827 PAD.n10826 2.2505
R38024 PAD.n10873 PAD.n10872 2.2505
R38025 PAD.n10874 PAD.n10825 2.2505
R38026 PAD.n10876 PAD.n10875 2.2505
R38027 PAD.n10823 PAD.n10822 2.2505
R38028 PAD.n10885 PAD.n10884 2.2505
R38029 PAD.n10886 PAD.n10821 2.2505
R38030 PAD.n10888 PAD.n10887 2.2505
R38031 PAD.n10819 PAD.n10818 2.2505
R38032 PAD.n10897 PAD.n10896 2.2505
R38033 PAD.n10898 PAD.n10817 2.2505
R38034 PAD.n10900 PAD.n10899 2.2505
R38035 PAD.n10815 PAD.n10814 2.2505
R38036 PAD.n10909 PAD.n10908 2.2505
R38037 PAD.n10910 PAD.n10813 2.2505
R38038 PAD.n10912 PAD.n10911 2.2505
R38039 PAD.n10811 PAD.n10810 2.2505
R38040 PAD.n10921 PAD.n10920 2.2505
R38041 PAD.n10922 PAD.n10809 2.2505
R38042 PAD.n10924 PAD.n10923 2.2505
R38043 PAD.n10807 PAD.n10806 2.2505
R38044 PAD.n10933 PAD.n10932 2.2505
R38045 PAD.n10934 PAD.n10805 2.2505
R38046 PAD.n10936 PAD.n10935 2.2505
R38047 PAD.n10803 PAD.n10802 2.2505
R38048 PAD.n10945 PAD.n10944 2.2505
R38049 PAD.n10946 PAD.n10801 2.2505
R38050 PAD.n10948 PAD.n10947 2.2505
R38051 PAD.n10799 PAD.n10798 2.2505
R38052 PAD.n10957 PAD.n10956 2.2505
R38053 PAD.n10958 PAD.n10797 2.2505
R38054 PAD.n10960 PAD.n10959 2.2505
R38055 PAD.n10795 PAD.n10794 2.2505
R38056 PAD.n10969 PAD.n10968 2.2505
R38057 PAD.n10970 PAD.n10793 2.2505
R38058 PAD.n10972 PAD.n10971 2.2505
R38059 PAD.n10791 PAD.n10790 2.2505
R38060 PAD.n10981 PAD.n10980 2.2505
R38061 PAD.n10982 PAD.n10789 2.2505
R38062 PAD.n10984 PAD.n10983 2.2505
R38063 PAD.n10787 PAD.n10786 2.2505
R38064 PAD.n10993 PAD.n10992 2.2505
R38065 PAD.n10994 PAD.n10785 2.2505
R38066 PAD.n10996 PAD.n10995 2.2505
R38067 PAD.n10783 PAD.n10782 2.2505
R38068 PAD.n11005 PAD.n11004 2.2505
R38069 PAD.n11006 PAD.n10781 2.2505
R38070 PAD.n11008 PAD.n11007 2.2505
R38071 PAD.n10779 PAD.n10778 2.2505
R38072 PAD.n11017 PAD.n11016 2.2505
R38073 PAD.n11018 PAD.n10777 2.2505
R38074 PAD.n11020 PAD.n11019 2.2505
R38075 PAD.n10775 PAD.n10774 2.2505
R38076 PAD.n11029 PAD.n11028 2.2505
R38077 PAD.n11030 PAD.n10773 2.2505
R38078 PAD.n11032 PAD.n11031 2.2505
R38079 PAD.n10771 PAD.n10770 2.2505
R38080 PAD.n11041 PAD.n11040 2.2505
R38081 PAD.n11042 PAD.n10769 2.2505
R38082 PAD.n11044 PAD.n11043 2.2505
R38083 PAD.n10767 PAD.n10766 2.2505
R38084 PAD.n11053 PAD.n11052 2.2505
R38085 PAD.n11054 PAD.n10765 2.2505
R38086 PAD.n11056 PAD.n11055 2.2505
R38087 PAD.n10763 PAD.n10762 2.2505
R38088 PAD.n11065 PAD.n11064 2.2505
R38089 PAD.n11066 PAD.n10761 2.2505
R38090 PAD.n11068 PAD.n11067 2.2505
R38091 PAD.n10759 PAD.n10758 2.2505
R38092 PAD.n11077 PAD.n11076 2.2505
R38093 PAD.n11078 PAD.n10757 2.2505
R38094 PAD.n11080 PAD.n11079 2.2505
R38095 PAD.n10749 PAD.n10747 2.2505
R38096 PAD.n11087 PAD.n11086 2.2505
R38097 PAD.n11086 PAD.n11085 2.2505
R38098 PAD.n11083 PAD.n10749 2.2505
R38099 PAD.n11081 PAD.n11080 2.2505
R38100 PAD.n11073 PAD.n10757 2.2505
R38101 PAD.n11076 PAD.n11075 2.2505
R38102 PAD.n11071 PAD.n10759 2.2505
R38103 PAD.n11069 PAD.n11068 2.2505
R38104 PAD.n11061 PAD.n10761 2.2505
R38105 PAD.n11064 PAD.n11063 2.2505
R38106 PAD.n11059 PAD.n10763 2.2505
R38107 PAD.n11057 PAD.n11056 2.2505
R38108 PAD.n11049 PAD.n10765 2.2505
R38109 PAD.n11052 PAD.n11051 2.2505
R38110 PAD.n11047 PAD.n10767 2.2505
R38111 PAD.n11045 PAD.n11044 2.2505
R38112 PAD.n11037 PAD.n10769 2.2505
R38113 PAD.n11040 PAD.n11039 2.2505
R38114 PAD.n11035 PAD.n10771 2.2505
R38115 PAD.n11033 PAD.n11032 2.2505
R38116 PAD.n11025 PAD.n10773 2.2505
R38117 PAD.n11028 PAD.n11027 2.2505
R38118 PAD.n11023 PAD.n10775 2.2505
R38119 PAD.n11021 PAD.n11020 2.2505
R38120 PAD.n11013 PAD.n10777 2.2505
R38121 PAD.n11016 PAD.n11015 2.2505
R38122 PAD.n11011 PAD.n10779 2.2505
R38123 PAD.n11009 PAD.n11008 2.2505
R38124 PAD.n11001 PAD.n10781 2.2505
R38125 PAD.n11004 PAD.n11003 2.2505
R38126 PAD.n10999 PAD.n10783 2.2505
R38127 PAD.n10997 PAD.n10996 2.2505
R38128 PAD.n10989 PAD.n10785 2.2505
R38129 PAD.n10992 PAD.n10991 2.2505
R38130 PAD.n10987 PAD.n10787 2.2505
R38131 PAD.n10985 PAD.n10984 2.2505
R38132 PAD.n10977 PAD.n10789 2.2505
R38133 PAD.n10980 PAD.n10979 2.2505
R38134 PAD.n10975 PAD.n10791 2.2505
R38135 PAD.n10973 PAD.n10972 2.2505
R38136 PAD.n10965 PAD.n10793 2.2505
R38137 PAD.n10968 PAD.n10967 2.2505
R38138 PAD.n10963 PAD.n10795 2.2505
R38139 PAD.n10961 PAD.n10960 2.2505
R38140 PAD.n10953 PAD.n10797 2.2505
R38141 PAD.n10956 PAD.n10955 2.2505
R38142 PAD.n10951 PAD.n10799 2.2505
R38143 PAD.n10949 PAD.n10948 2.2505
R38144 PAD.n10941 PAD.n10801 2.2505
R38145 PAD.n10944 PAD.n10943 2.2505
R38146 PAD.n10939 PAD.n10803 2.2505
R38147 PAD.n10937 PAD.n10936 2.2505
R38148 PAD.n10929 PAD.n10805 2.2505
R38149 PAD.n10932 PAD.n10931 2.2505
R38150 PAD.n10927 PAD.n10807 2.2505
R38151 PAD.n10925 PAD.n10924 2.2505
R38152 PAD.n10917 PAD.n10809 2.2505
R38153 PAD.n10920 PAD.n10919 2.2505
R38154 PAD.n10915 PAD.n10811 2.2505
R38155 PAD.n10913 PAD.n10912 2.2505
R38156 PAD.n10905 PAD.n10813 2.2505
R38157 PAD.n10908 PAD.n10907 2.2505
R38158 PAD.n10903 PAD.n10815 2.2505
R38159 PAD.n10901 PAD.n10900 2.2505
R38160 PAD.n10893 PAD.n10817 2.2505
R38161 PAD.n10896 PAD.n10895 2.2505
R38162 PAD.n10891 PAD.n10819 2.2505
R38163 PAD.n10889 PAD.n10888 2.2505
R38164 PAD.n10881 PAD.n10821 2.2505
R38165 PAD.n10884 PAD.n10883 2.2505
R38166 PAD.n10879 PAD.n10823 2.2505
R38167 PAD.n10877 PAD.n10876 2.2505
R38168 PAD.n10869 PAD.n10825 2.2505
R38169 PAD.n10872 PAD.n10871 2.2505
R38170 PAD.n10867 PAD.n10827 2.2505
R38171 PAD.n10865 PAD.n10864 2.2505
R38172 PAD.n10857 PAD.n10829 2.2505
R38173 PAD.n10860 PAD.n10859 2.2505
R38174 PAD.n10855 PAD.n10831 2.2505
R38175 PAD.n10853 PAD.n10852 2.2505
R38176 PAD.n10845 PAD.n10833 2.2505
R38177 PAD.n10848 PAD.n10847 2.2505
R38178 PAD.n10843 PAD.n10835 2.2505
R38179 PAD.n10841 PAD.n10840 2.2505
R38180 PAD.n10838 PAD.n10837 2.2505
R38181 PAD.n6382 PAD.n6381 2.2505
R38182 PAD.n5977 PAD.n5975 2.2505
R38183 PAD.n5973 PAD.n5952 2.2505
R38184 PAD.n6685 PAD.n6684 2.2505
R38185 PAD.n5560 PAD.n5559 2.2505
R38186 PAD.n6702 PAD.n6701 2.2505
R38187 PAD.n7800 PAD.n7799 2.2505
R38188 PAD.n5556 PAD.n5554 2.2505
R38189 PAD.n7794 PAD.n7793 2.2505
R38190 PAD.n6710 PAD.n6708 2.2505
R38191 PAD.n7152 PAD.n7149 2.2505
R38192 PAD.n7529 PAD.n7527 2.2505
R38193 PAD.n7151 PAD.n7150 2.2505
R38194 PAD.n7523 PAD.n7522 2.2505
R38195 PAD.n7205 PAD.n7204 2.2505
R38196 PAD.n5203 PAD.n5202 2.2505
R38197 PAD.n7822 PAD.n7821 2.2505
R38198 PAD.n7827 PAD.n7826 2.2505
R38199 PAD.n5189 PAD.n5188 2.2505
R38200 PAD.n8177 PAD.n8176 2.2505
R38201 PAD.n8182 PAD.n8181 2.2505
R38202 PAD.n4838 PAD.n4837 2.2505
R38203 PAD.n8197 PAD.n8196 2.2505
R38204 PAD.n8201 PAD.n4833 2.2505
R38205 PAD.n8203 PAD.n8202 2.2505
R38206 PAD.n8207 PAD.n8206 2.2505
R38207 PAD.n4672 PAD.n4671 2.2505
R38208 PAD.n8412 PAD.n8411 2.2505
R38209 PAD.n8418 PAD.n8417 2.2505
R38210 PAD.n4318 PAD.n4317 2.2505
R38211 PAD.n8433 PAD.n8432 2.2505
R38212 PAD.n8435 PAD.n3976 2.2505
R38213 PAD.n8455 PAD.n3975 2.2505
R38214 PAD.n8457 PAD.n8456 2.2505
R38215 PAD.n8459 PAD.n3632 2.2505
R38216 PAD.n8480 PAD.n3630 2.2505
R38217 PAD.n8482 PAD.n8481 2.2505
R38218 PAD.n3286 PAD.n3285 2.2505
R38219 PAD.n8505 PAD.n8504 2.2505
R38220 PAD.n8508 PAD.n8507 2.2505
R38221 PAD.n2902 PAD.n2900 2.2505
R38222 PAD.n8824 PAD.n8823 2.2505
R38223 PAD.n2896 PAD.n2893 2.2505
R38224 PAD.n8830 PAD.n8829 2.2505
R38225 PAD.n2897 PAD.n2895 2.2505
R38226 PAD.n9131 PAD.n9130 2.2505
R38227 PAD.n2493 PAD.n2492 2.2505
R38228 PAD.n9154 PAD.n9153 2.2505
R38229 PAD.n9159 PAD.n9158 2.2505
R38230 PAD.n2145 PAD.n2144 2.2505
R38231 PAD.n9178 PAD.n9177 2.2505
R38232 PAD.n9183 PAD.n9182 2.2505
R38233 PAD.n2044 PAD.n2042 2.2505
R38234 PAD.n9448 PAD.n9447 2.2505
R38235 PAD.n2039 PAD.n2038 2.2505
R38236 PAD.n9454 PAD.n9453 2.2505
R38237 PAD.n9715 PAD.n9714 2.2505
R38238 PAD.n1938 PAD.n1937 2.2505
R38239 PAD.n9720 PAD.n9719 2.2505
R38240 PAD.n9735 PAD.n9734 2.2505
R38241 PAD.n1588 PAD.n1587 2.2505
R38242 PAD.n9740 PAD.n9739 2.2505
R38243 PAD.n10001 PAD.n10000 2.2505
R38244 PAD.n1485 PAD.n1484 2.2505
R38245 PAD.n10006 PAD.n10005 2.2505
R38246 PAD.n10019 PAD.n10018 2.2505
R38247 PAD.n1135 PAD.n1133 2.2505
R38248 PAD.n10360 PAD.n10359 2.2505
R38249 PAD.n1117 PAD.n1116 2.2505
R38250 PAD.n10376 PAD.n10375 2.2505
R38251 PAD.n10379 PAD.n10378 2.2505
R38252 PAD.n775 PAD.n774 2.2505
R38253 PAD.n10400 PAD.n10399 2.2505
R38254 PAD.n10406 PAD.n10405 2.2505
R38255 PAD.n424 PAD.n423 2.2505
R38256 PAD.n10704 PAD.n10703 2.2505
R38257 PAD.n10707 PAD.n10706 2.2505
R38258 PAD.n30 PAD.n28 2.2505
R38259 PAD.n10730 PAD.n10729 2.2505
R38260 PAD.n24 PAD.n22 2.2505
R38261 PAD.n11531 PAD.n11530 2.2505
R38262 PAD.n25 PAD.n23 2.2505
R38263 PAD.n11525 PAD.n11524 2.2505
R38264 PAD.n10739 PAD.n10737 2.2505
R38265 PAD.n11503 PAD.n11502 2.2505
R38266 PAD.n6691 PAD.n6690 2.2505
R38267 PAD.n5905 PAD.n5900 2.2505
R38268 PAD.n6498 PAD.n6497 2.2505
R38269 PAD.n6496 PAD.n6495 2.2505
R38270 PAD.n6503 PAD.n6502 2.2505
R38271 PAD.n6505 PAD.n6504 2.2505
R38272 PAD.n6507 PAD.n6506 2.2505
R38273 PAD.n6493 PAD.n6492 2.2505
R38274 PAD.n6512 PAD.n6511 2.2505
R38275 PAD.n6514 PAD.n6513 2.2505
R38276 PAD.n6516 PAD.n6515 2.2505
R38277 PAD.n6490 PAD.n6489 2.2505
R38278 PAD.n6521 PAD.n6520 2.2505
R38279 PAD.n6523 PAD.n6522 2.2505
R38280 PAD.n6525 PAD.n6524 2.2505
R38281 PAD.n6487 PAD.n6486 2.2505
R38282 PAD.n6530 PAD.n6529 2.2505
R38283 PAD.n6532 PAD.n6531 2.2505
R38284 PAD.n6534 PAD.n6533 2.2505
R38285 PAD.n6484 PAD.n6483 2.2505
R38286 PAD.n6539 PAD.n6538 2.2505
R38287 PAD.n6541 PAD.n6540 2.2505
R38288 PAD.n6543 PAD.n6542 2.2505
R38289 PAD.n6481 PAD.n6480 2.2505
R38290 PAD.n6548 PAD.n6547 2.2505
R38291 PAD.n6550 PAD.n6549 2.2505
R38292 PAD.n6552 PAD.n6551 2.2505
R38293 PAD.n6478 PAD.n6477 2.2505
R38294 PAD.n6557 PAD.n6556 2.2505
R38295 PAD.n6559 PAD.n6558 2.2505
R38296 PAD.n6561 PAD.n6560 2.2505
R38297 PAD.n6475 PAD.n6474 2.2505
R38298 PAD.n6566 PAD.n6565 2.2505
R38299 PAD.n6568 PAD.n6567 2.2505
R38300 PAD.n6570 PAD.n6569 2.2505
R38301 PAD.n6472 PAD.n6471 2.2505
R38302 PAD.n6575 PAD.n6574 2.2505
R38303 PAD.n6577 PAD.n6576 2.2505
R38304 PAD.n6579 PAD.n6578 2.2505
R38305 PAD.n6469 PAD.n6468 2.2505
R38306 PAD.n6584 PAD.n6583 2.2505
R38307 PAD.n6586 PAD.n6585 2.2505
R38308 PAD.n6588 PAD.n6587 2.2505
R38309 PAD.n6466 PAD.n6465 2.2505
R38310 PAD.n6593 PAD.n6592 2.2505
R38311 PAD.n6595 PAD.n6594 2.2505
R38312 PAD.n6597 PAD.n6596 2.2505
R38313 PAD.n6463 PAD.n6462 2.2505
R38314 PAD.n6602 PAD.n6601 2.2505
R38315 PAD.n6604 PAD.n6603 2.2505
R38316 PAD.n6606 PAD.n6605 2.2505
R38317 PAD.n6460 PAD.n6459 2.2505
R38318 PAD.n6611 PAD.n6610 2.2505
R38319 PAD.n6613 PAD.n6612 2.2505
R38320 PAD.n6615 PAD.n6614 2.2505
R38321 PAD.n6457 PAD.n6456 2.2505
R38322 PAD.n6620 PAD.n6619 2.2505
R38323 PAD.n6622 PAD.n6621 2.2505
R38324 PAD.n6624 PAD.n6623 2.2505
R38325 PAD.n6454 PAD.n6453 2.2505
R38326 PAD.n6629 PAD.n6628 2.2505
R38327 PAD.n6631 PAD.n6630 2.2505
R38328 PAD.n6633 PAD.n6632 2.2505
R38329 PAD.n6451 PAD.n6450 2.2505
R38330 PAD.n6638 PAD.n6637 2.2505
R38331 PAD.n6640 PAD.n6639 2.2505
R38332 PAD.n6642 PAD.n6641 2.2505
R38333 PAD.n6448 PAD.n6447 2.2505
R38334 PAD.n6647 PAD.n6646 2.2505
R38335 PAD.n6649 PAD.n6648 2.2505
R38336 PAD.n6651 PAD.n6650 2.2505
R38337 PAD.n6445 PAD.n6444 2.2505
R38338 PAD.n6656 PAD.n6655 2.2505
R38339 PAD.n6658 PAD.n6657 2.2505
R38340 PAD.n6660 PAD.n6659 2.2505
R38341 PAD.n6442 PAD.n6441 2.2505
R38342 PAD.n6665 PAD.n6664 2.2505
R38343 PAD.n6667 PAD.n6666 2.2505
R38344 PAD.n6669 PAD.n6668 2.2505
R38345 PAD.n6438 PAD.n6437 2.2505
R38346 PAD.n6676 PAD.n6675 2.2505
R38347 PAD.n6439 PAD.n6436 2.2505
R38348 PAD.n5950 PAD.n5949 2.2505
R38349 PAD.n6688 PAD.n6687 2.2505
R38350 PAD.n6383 PAD.n6382 2.2505
R38351 PAD.n5975 PAD.n5974 2.2505
R38352 PAD.n5973 PAD.n5904 2.2505
R38353 PAD.n6684 PAD.n6683 2.2505
R38354 PAD.n6680 PAD.n5560 2.2505
R38355 PAD.n6701 PAD.n6700 2.2505
R38356 PAD.n7801 PAD.n7800 2.2505
R38357 PAD.n6711 PAD.n5554 2.2505
R38358 PAD.n7793 PAD.n7792 2.2505
R38359 PAD.n7059 PAD.n6710 2.2505
R38360 PAD.n7149 PAD.n7061 2.2505
R38361 PAD.n7529 PAD.n7528 2.2505
R38362 PAD.n7215 PAD.n7150 2.2505
R38363 PAD.n7522 PAD.n7521 2.2505
R38364 PAD.n7206 PAD.n7205 2.2505
R38365 PAD.n7222 PAD.n5203 2.2505
R38366 PAD.n7821 PAD.n7820 2.2505
R38367 PAD.n7828 PAD.n7827 2.2505
R38368 PAD.n8164 PAD.n5189 2.2505
R38369 PAD.n8176 PAD.n8175 2.2505
R38370 PAD.n8183 PAD.n8182 2.2505
R38371 PAD.n8185 PAD.n4838 2.2505
R38372 PAD.n8196 PAD.n8195 2.2505
R38373 PAD.n4842 PAD.n4833 2.2505
R38374 PAD.n8203 PAD.n4682 2.2505
R38375 PAD.n8206 PAD.n8205 2.2505
R38376 PAD.n8408 PAD.n4672 2.2505
R38377 PAD.n8411 PAD.n8410 2.2505
R38378 PAD.n8419 PAD.n8418 2.2505
R38379 PAD.n4319 PAD.n4318 2.2505
R38380 PAD.n8432 PAD.n8431 2.2505
R38381 PAD.n3983 PAD.n3976 2.2505
R38382 PAD.n8455 PAD.n8454 2.2505
R38383 PAD.n8456 PAD.n3641 2.2505
R38384 PAD.n3684 PAD.n3632 2.2505
R38385 PAD.n8480 PAD.n8479 2.2505
R38386 PAD.n8481 PAD.n3296 2.2505
R38387 PAD.n3339 PAD.n3286 2.2505
R38388 PAD.n8504 PAD.n8503 2.2505
R38389 PAD.n8507 PAD.n2952 2.2505
R38390 PAD.n8518 PAD.n2902 2.2505
R38391 PAD.n8823 PAD.n8822 2.2505
R38392 PAD.n2946 PAD.n2893 2.2505
R38393 PAD.n8831 PAD.n8830 2.2505
R38394 PAD.n2895 PAD.n2894 2.2505
R38395 PAD.n9130 PAD.n9129 2.2505
R38396 PAD.n9142 PAD.n2493 2.2505
R38397 PAD.n9153 PAD.n9152 2.2505
R38398 PAD.n9160 PAD.n9159 2.2505
R38399 PAD.n9162 PAD.n2145 2.2505
R38400 PAD.n9177 PAD.n9176 2.2505
R38401 PAD.n9184 PAD.n9183 2.2505
R38402 PAD.n9186 PAD.n2044 2.2505
R38403 PAD.n9447 PAD.n9446 2.2505
R38404 PAD.n2038 PAD.n2037 2.2505
R38405 PAD.n9455 PAD.n9454 2.2505
R38406 PAD.n9714 PAD.n9713 2.2505
R38407 PAD.n1985 PAD.n1937 2.2505
R38408 PAD.n9721 PAD.n9720 2.2505
R38409 PAD.n9734 PAD.n9733 2.2505
R38410 PAD.n1587 PAD.n1586 2.2505
R38411 PAD.n9741 PAD.n9740 2.2505
R38412 PAD.n10000 PAD.n9999 2.2505
R38413 PAD.n1533 PAD.n1484 2.2505
R38414 PAD.n10007 PAD.n10006 2.2505
R38415 PAD.n10018 PAD.n10017 2.2505
R38416 PAD.n1142 PAD.n1133 2.2505
R38417 PAD.n10361 PAD.n10360 2.2505
R38418 PAD.n1118 PAD.n1117 2.2505
R38419 PAD.n10375 PAD.n10374 2.2505
R38420 PAD.n10378 PAD.n782 2.2505
R38421 PAD.n825 PAD.n775 2.2505
R38422 PAD.n10399 PAD.n10398 2.2505
R38423 PAD.n10407 PAD.n10406 2.2505
R38424 PAD.n425 PAD.n424 2.2505
R38425 PAD.n10703 PAD.n10702 2.2505
R38426 PAD.n10706 PAD.n373 2.2505
R38427 PAD.n10718 PAD.n30 2.2505
R38428 PAD.n10729 PAD.n10728 2.2505
R38429 PAD.n22 PAD.n20 2.2505
R38430 PAD.n11532 PAD.n11531 2.2505
R38431 PAD.n10754 PAD.n23 2.2505
R38432 PAD.n11524 PAD.n11523 2.2505
R38433 PAD.n10741 PAD.n10739 2.2505
R38434 PAD.n11502 PAD.n11501 2.2505
R38435 PAD.n11155 PAD.n11105 2.24752
R38436 PAD.n6031 PAD.n5980 2.24752
R38437 PAD.n11157 PAD.n11100 2.24752
R38438 PAD.n11302 PAD.n11254 2.24752
R38439 PAD.n11159 PAD.n11100 2.24752
R38440 PAD.n11302 PAD.n11255 2.24752
R38441 PAD.n11161 PAD.n11100 2.24752
R38442 PAD.n11302 PAD.n11256 2.24752
R38443 PAD.n11163 PAD.n11100 2.24752
R38444 PAD.n11302 PAD.n11257 2.24752
R38445 PAD.n11165 PAD.n11100 2.24752
R38446 PAD.n11302 PAD.n11258 2.24752
R38447 PAD.n11167 PAD.n11100 2.24752
R38448 PAD.n11302 PAD.n11259 2.24752
R38449 PAD.n11169 PAD.n11100 2.24752
R38450 PAD.n11302 PAD.n11260 2.24752
R38451 PAD.n11171 PAD.n11100 2.24752
R38452 PAD.n11302 PAD.n11261 2.24752
R38453 PAD.n11173 PAD.n11100 2.24752
R38454 PAD.n11302 PAD.n11262 2.24752
R38455 PAD.n11175 PAD.n11100 2.24752
R38456 PAD.n11302 PAD.n11263 2.24752
R38457 PAD.n11177 PAD.n11100 2.24752
R38458 PAD.n11302 PAD.n11264 2.24752
R38459 PAD.n11179 PAD.n11100 2.24752
R38460 PAD.n11302 PAD.n11265 2.24752
R38461 PAD.n11181 PAD.n11100 2.24752
R38462 PAD.n11302 PAD.n11266 2.24752
R38463 PAD.n11183 PAD.n11100 2.24752
R38464 PAD.n11302 PAD.n11267 2.24752
R38465 PAD.n11185 PAD.n11100 2.24752
R38466 PAD.n11302 PAD.n11268 2.24752
R38467 PAD.n11187 PAD.n11100 2.24752
R38468 PAD.n11302 PAD.n11269 2.24752
R38469 PAD.n11189 PAD.n11100 2.24752
R38470 PAD.n11302 PAD.n11270 2.24752
R38471 PAD.n11191 PAD.n11100 2.24752
R38472 PAD.n11302 PAD.n11271 2.24752
R38473 PAD.n11193 PAD.n11100 2.24752
R38474 PAD.n11302 PAD.n11272 2.24752
R38475 PAD.n11195 PAD.n11100 2.24752
R38476 PAD.n11302 PAD.n11273 2.24752
R38477 PAD.n11197 PAD.n11100 2.24752
R38478 PAD.n11302 PAD.n11274 2.24752
R38479 PAD.n11199 PAD.n11100 2.24752
R38480 PAD.n11302 PAD.n11275 2.24752
R38481 PAD.n11201 PAD.n11100 2.24752
R38482 PAD.n11302 PAD.n11276 2.24752
R38483 PAD.n11203 PAD.n11100 2.24752
R38484 PAD.n11302 PAD.n11277 2.24752
R38485 PAD.n11205 PAD.n11100 2.24752
R38486 PAD.n11302 PAD.n11278 2.24752
R38487 PAD.n11207 PAD.n11100 2.24752
R38488 PAD.n11302 PAD.n11279 2.24752
R38489 PAD.n11209 PAD.n11100 2.24752
R38490 PAD.n11302 PAD.n11280 2.24752
R38491 PAD.n11211 PAD.n11100 2.24752
R38492 PAD.n11302 PAD.n11281 2.24752
R38493 PAD.n11213 PAD.n11100 2.24752
R38494 PAD.n11302 PAD.n11282 2.24752
R38495 PAD.n11215 PAD.n11100 2.24752
R38496 PAD.n11302 PAD.n11283 2.24752
R38497 PAD.n11217 PAD.n11100 2.24752
R38498 PAD.n11302 PAD.n11284 2.24752
R38499 PAD.n11219 PAD.n11100 2.24752
R38500 PAD.n11302 PAD.n11285 2.24752
R38501 PAD.n11221 PAD.n11100 2.24752
R38502 PAD.n11302 PAD.n11286 2.24752
R38503 PAD.n11223 PAD.n11100 2.24752
R38504 PAD.n11302 PAD.n11287 2.24752
R38505 PAD.n11225 PAD.n11100 2.24752
R38506 PAD.n11302 PAD.n11288 2.24752
R38507 PAD.n11227 PAD.n11100 2.24752
R38508 PAD.n11302 PAD.n11289 2.24752
R38509 PAD.n11229 PAD.n11100 2.24752
R38510 PAD.n11302 PAD.n11290 2.24752
R38511 PAD.n11231 PAD.n11100 2.24752
R38512 PAD.n11302 PAD.n11291 2.24752
R38513 PAD.n11233 PAD.n11100 2.24752
R38514 PAD.n11302 PAD.n11292 2.24752
R38515 PAD.n11235 PAD.n11100 2.24752
R38516 PAD.n11302 PAD.n11293 2.24752
R38517 PAD.n11237 PAD.n11100 2.24752
R38518 PAD.n11302 PAD.n11294 2.24752
R38519 PAD.n11239 PAD.n11100 2.24752
R38520 PAD.n11302 PAD.n11295 2.24752
R38521 PAD.n11241 PAD.n11100 2.24752
R38522 PAD.n11302 PAD.n11296 2.24752
R38523 PAD.n11243 PAD.n11100 2.24752
R38524 PAD.n11302 PAD.n11297 2.24752
R38525 PAD.n11245 PAD.n11100 2.24752
R38526 PAD.n11302 PAD.n11298 2.24752
R38527 PAD.n11247 PAD.n11100 2.24752
R38528 PAD.n11302 PAD.n11299 2.24752
R38529 PAD.n11249 PAD.n11100 2.24752
R38530 PAD.n11302 PAD.n11300 2.24752
R38531 PAD.n11251 PAD.n11100 2.24752
R38532 PAD.n11302 PAD.n11301 2.24752
R38533 PAD.n5966 PAD.n5961 2.24752
R38534 PAD.n11510 PAD.n11095 2.24752
R38535 PAD.n6384 PAD.n5966 2.24752
R38536 PAD.n11511 PAD.n11510 2.24752
R38537 PAD.n6033 PAD.n5982 2.24752
R38538 PAD.n6035 PAD.n5980 2.24752
R38539 PAD.n6036 PAD.n5982 2.24752
R38540 PAD.n6038 PAD.n5980 2.24752
R38541 PAD.n6039 PAD.n5982 2.24752
R38542 PAD.n6041 PAD.n5980 2.24752
R38543 PAD.n6042 PAD.n5982 2.24752
R38544 PAD.n6044 PAD.n5980 2.24752
R38545 PAD.n6045 PAD.n5982 2.24752
R38546 PAD.n6047 PAD.n5980 2.24752
R38547 PAD.n6048 PAD.n5982 2.24752
R38548 PAD.n6050 PAD.n5980 2.24752
R38549 PAD.n6051 PAD.n5982 2.24752
R38550 PAD.n6053 PAD.n5980 2.24752
R38551 PAD.n6054 PAD.n5982 2.24752
R38552 PAD.n6056 PAD.n5980 2.24752
R38553 PAD.n6057 PAD.n5982 2.24752
R38554 PAD.n6059 PAD.n5980 2.24752
R38555 PAD.n6060 PAD.n5982 2.24752
R38556 PAD.n6062 PAD.n5980 2.24752
R38557 PAD.n6063 PAD.n5982 2.24752
R38558 PAD.n6065 PAD.n5980 2.24752
R38559 PAD.n6066 PAD.n5982 2.24752
R38560 PAD.n6068 PAD.n5980 2.24752
R38561 PAD.n6069 PAD.n5982 2.24752
R38562 PAD.n6071 PAD.n5980 2.24752
R38563 PAD.n6072 PAD.n5982 2.24752
R38564 PAD.n6074 PAD.n5980 2.24752
R38565 PAD.n6075 PAD.n5982 2.24752
R38566 PAD.n6077 PAD.n5980 2.24752
R38567 PAD.n6078 PAD.n5982 2.24752
R38568 PAD.n6080 PAD.n5980 2.24752
R38569 PAD.n6081 PAD.n5982 2.24752
R38570 PAD.n6083 PAD.n5980 2.24752
R38571 PAD.n6084 PAD.n5982 2.24752
R38572 PAD.n6086 PAD.n5980 2.24752
R38573 PAD.n6087 PAD.n5982 2.24752
R38574 PAD.n6089 PAD.n5980 2.24752
R38575 PAD.n6090 PAD.n5982 2.24752
R38576 PAD.n6092 PAD.n5980 2.24752
R38577 PAD.n6093 PAD.n5982 2.24752
R38578 PAD.n6095 PAD.n5980 2.24752
R38579 PAD.n6096 PAD.n5982 2.24752
R38580 PAD.n6098 PAD.n5980 2.24752
R38581 PAD.n6099 PAD.n5982 2.24752
R38582 PAD.n6101 PAD.n5980 2.24752
R38583 PAD.n6102 PAD.n5982 2.24752
R38584 PAD.n6104 PAD.n5980 2.24752
R38585 PAD.n6105 PAD.n5982 2.24752
R38586 PAD.n6107 PAD.n5980 2.24752
R38587 PAD.n6108 PAD.n5982 2.24752
R38588 PAD.n6110 PAD.n5980 2.24752
R38589 PAD.n6111 PAD.n5982 2.24752
R38590 PAD.n6113 PAD.n5980 2.24752
R38591 PAD.n6114 PAD.n5982 2.24752
R38592 PAD.n6116 PAD.n5980 2.24752
R38593 PAD.n6117 PAD.n5982 2.24752
R38594 PAD.n6119 PAD.n5980 2.24752
R38595 PAD.n6120 PAD.n5982 2.24752
R38596 PAD.n6122 PAD.n5980 2.24752
R38597 PAD.n6123 PAD.n5982 2.24752
R38598 PAD.n6125 PAD.n5980 2.24752
R38599 PAD.n6126 PAD.n5982 2.24752
R38600 PAD.n6128 PAD.n5980 2.24752
R38601 PAD.n6129 PAD.n5982 2.24752
R38602 PAD.n6131 PAD.n5980 2.24752
R38603 PAD.n6132 PAD.n5982 2.24752
R38604 PAD.n6134 PAD.n5980 2.24752
R38605 PAD.n6135 PAD.n5982 2.24752
R38606 PAD.n6137 PAD.n5980 2.24752
R38607 PAD.n6138 PAD.n5982 2.24752
R38608 PAD.n6140 PAD.n5980 2.24752
R38609 PAD.n6141 PAD.n5982 2.24752
R38610 PAD.n6143 PAD.n5980 2.24752
R38611 PAD.n6144 PAD.n5982 2.24752
R38612 PAD.n6146 PAD.n5980 2.24752
R38613 PAD.n6147 PAD.n5982 2.24752
R38614 PAD.n6149 PAD.n5980 2.24752
R38615 PAD.n6150 PAD.n5982 2.24752
R38616 PAD.n6152 PAD.n5980 2.24752
R38617 PAD.n6153 PAD.n5982 2.24752
R38618 PAD.n6155 PAD.n5980 2.24752
R38619 PAD.n6156 PAD.n5982 2.24752
R38620 PAD.n6158 PAD.n5980 2.24752
R38621 PAD.n6159 PAD.n5982 2.24752
R38622 PAD.n6161 PAD.n5980 2.24752
R38623 PAD.n6162 PAD.n5982 2.24752
R38624 PAD.n6164 PAD.n5980 2.24752
R38625 PAD.n6165 PAD.n5982 2.24752
R38626 PAD.n6167 PAD.n5980 2.24752
R38627 PAD.n6168 PAD.n5982 2.24752
R38628 PAD.n6170 PAD.n5980 2.24752
R38629 PAD.n6171 PAD.n5982 2.24752
R38630 PAD.n6173 PAD.n5980 2.24752
R38631 PAD.n6174 PAD.n5982 2.24752
R38632 PAD.n6176 PAD.n5982 2.24752
R38633 PAD.n11084 PAD.n10755 2.24164
R38634 PAD.n11082 PAD.n21 2.24164
R38635 PAD.n10756 PAD.n10755 2.24164
R38636 PAD.n11074 PAD.n21 2.24164
R38637 PAD.n11072 PAD.n10755 2.24164
R38638 PAD.n11070 PAD.n21 2.24164
R38639 PAD.n10760 PAD.n10755 2.24164
R38640 PAD.n11062 PAD.n21 2.24164
R38641 PAD.n11060 PAD.n10755 2.24164
R38642 PAD.n11058 PAD.n21 2.24164
R38643 PAD.n10764 PAD.n10755 2.24164
R38644 PAD.n11050 PAD.n21 2.24164
R38645 PAD.n11048 PAD.n10755 2.24164
R38646 PAD.n11046 PAD.n21 2.24164
R38647 PAD.n10768 PAD.n10755 2.24164
R38648 PAD.n11038 PAD.n21 2.24164
R38649 PAD.n11036 PAD.n10755 2.24164
R38650 PAD.n11034 PAD.n21 2.24164
R38651 PAD.n10772 PAD.n10755 2.24164
R38652 PAD.n11026 PAD.n21 2.24164
R38653 PAD.n11024 PAD.n10755 2.24164
R38654 PAD.n11022 PAD.n21 2.24164
R38655 PAD.n10776 PAD.n10755 2.24164
R38656 PAD.n11014 PAD.n21 2.24164
R38657 PAD.n11012 PAD.n10755 2.24164
R38658 PAD.n11010 PAD.n21 2.24164
R38659 PAD.n10780 PAD.n10755 2.24164
R38660 PAD.n11002 PAD.n21 2.24164
R38661 PAD.n11000 PAD.n10755 2.24164
R38662 PAD.n10998 PAD.n21 2.24164
R38663 PAD.n10784 PAD.n10755 2.24164
R38664 PAD.n10990 PAD.n21 2.24164
R38665 PAD.n10988 PAD.n10755 2.24164
R38666 PAD.n10986 PAD.n21 2.24164
R38667 PAD.n10788 PAD.n10755 2.24164
R38668 PAD.n10978 PAD.n21 2.24164
R38669 PAD.n10976 PAD.n10755 2.24164
R38670 PAD.n10974 PAD.n21 2.24164
R38671 PAD.n10792 PAD.n10755 2.24164
R38672 PAD.n10966 PAD.n21 2.24164
R38673 PAD.n10964 PAD.n10755 2.24164
R38674 PAD.n10962 PAD.n21 2.24164
R38675 PAD.n10796 PAD.n10755 2.24164
R38676 PAD.n10954 PAD.n21 2.24164
R38677 PAD.n10952 PAD.n10755 2.24164
R38678 PAD.n10950 PAD.n21 2.24164
R38679 PAD.n10800 PAD.n10755 2.24164
R38680 PAD.n10942 PAD.n21 2.24164
R38681 PAD.n10940 PAD.n10755 2.24164
R38682 PAD.n10938 PAD.n21 2.24164
R38683 PAD.n10804 PAD.n10755 2.24164
R38684 PAD.n10930 PAD.n21 2.24164
R38685 PAD.n10928 PAD.n10755 2.24164
R38686 PAD.n10926 PAD.n21 2.24164
R38687 PAD.n10808 PAD.n10755 2.24164
R38688 PAD.n10918 PAD.n21 2.24164
R38689 PAD.n10916 PAD.n10755 2.24164
R38690 PAD.n10914 PAD.n21 2.24164
R38691 PAD.n10812 PAD.n10755 2.24164
R38692 PAD.n10906 PAD.n21 2.24164
R38693 PAD.n10904 PAD.n10755 2.24164
R38694 PAD.n10902 PAD.n21 2.24164
R38695 PAD.n10816 PAD.n10755 2.24164
R38696 PAD.n10894 PAD.n21 2.24164
R38697 PAD.n10892 PAD.n10755 2.24164
R38698 PAD.n10890 PAD.n21 2.24164
R38699 PAD.n10820 PAD.n10755 2.24164
R38700 PAD.n10882 PAD.n21 2.24164
R38701 PAD.n10880 PAD.n10755 2.24164
R38702 PAD.n10878 PAD.n21 2.24164
R38703 PAD.n10824 PAD.n10755 2.24164
R38704 PAD.n10870 PAD.n21 2.24164
R38705 PAD.n10868 PAD.n10755 2.24164
R38706 PAD.n10866 PAD.n21 2.24164
R38707 PAD.n10828 PAD.n10755 2.24164
R38708 PAD.n10858 PAD.n21 2.24164
R38709 PAD.n10856 PAD.n10755 2.24164
R38710 PAD.n10854 PAD.n21 2.24164
R38711 PAD.n10832 PAD.n10755 2.24164
R38712 PAD.n10846 PAD.n21 2.24164
R38713 PAD.n10844 PAD.n10755 2.24164
R38714 PAD.n10842 PAD.n21 2.24164
R38715 PAD.n10836 PAD.n10755 2.24164
R38716 PAD.n116 PAD.n32 2.24164
R38717 PAD.n367 PAD.n73 2.24164
R38718 PAD.n125 PAD.n32 2.24164
R38719 PAD.n367 PAD.n72 2.24164
R38720 PAD.n129 PAD.n32 2.24164
R38721 PAD.n367 PAD.n71 2.24164
R38722 PAD.n137 PAD.n32 2.24164
R38723 PAD.n367 PAD.n70 2.24164
R38724 PAD.n141 PAD.n32 2.24164
R38725 PAD.n367 PAD.n69 2.24164
R38726 PAD.n149 PAD.n32 2.24164
R38727 PAD.n367 PAD.n68 2.24164
R38728 PAD.n153 PAD.n32 2.24164
R38729 PAD.n367 PAD.n67 2.24164
R38730 PAD.n161 PAD.n32 2.24164
R38731 PAD.n367 PAD.n66 2.24164
R38732 PAD.n165 PAD.n32 2.24164
R38733 PAD.n367 PAD.n65 2.24164
R38734 PAD.n173 PAD.n32 2.24164
R38735 PAD.n367 PAD.n64 2.24164
R38736 PAD.n177 PAD.n32 2.24164
R38737 PAD.n367 PAD.n63 2.24164
R38738 PAD.n185 PAD.n32 2.24164
R38739 PAD.n367 PAD.n62 2.24164
R38740 PAD.n189 PAD.n32 2.24164
R38741 PAD.n367 PAD.n61 2.24164
R38742 PAD.n197 PAD.n32 2.24164
R38743 PAD.n367 PAD.n60 2.24164
R38744 PAD.n201 PAD.n32 2.24164
R38745 PAD.n367 PAD.n59 2.24164
R38746 PAD.n209 PAD.n32 2.24164
R38747 PAD.n367 PAD.n58 2.24164
R38748 PAD.n213 PAD.n32 2.24164
R38749 PAD.n367 PAD.n57 2.24164
R38750 PAD.n221 PAD.n32 2.24164
R38751 PAD.n367 PAD.n56 2.24164
R38752 PAD.n225 PAD.n32 2.24164
R38753 PAD.n367 PAD.n55 2.24164
R38754 PAD.n233 PAD.n32 2.24164
R38755 PAD.n367 PAD.n54 2.24164
R38756 PAD.n237 PAD.n32 2.24164
R38757 PAD.n367 PAD.n53 2.24164
R38758 PAD.n245 PAD.n32 2.24164
R38759 PAD.n367 PAD.n52 2.24164
R38760 PAD.n249 PAD.n32 2.24164
R38761 PAD.n367 PAD.n51 2.24164
R38762 PAD.n257 PAD.n32 2.24164
R38763 PAD.n367 PAD.n50 2.24164
R38764 PAD.n261 PAD.n32 2.24164
R38765 PAD.n367 PAD.n49 2.24164
R38766 PAD.n269 PAD.n32 2.24164
R38767 PAD.n367 PAD.n48 2.24164
R38768 PAD.n273 PAD.n32 2.24164
R38769 PAD.n367 PAD.n47 2.24164
R38770 PAD.n281 PAD.n32 2.24164
R38771 PAD.n367 PAD.n46 2.24164
R38772 PAD.n285 PAD.n32 2.24164
R38773 PAD.n367 PAD.n45 2.24164
R38774 PAD.n293 PAD.n32 2.24164
R38775 PAD.n367 PAD.n44 2.24164
R38776 PAD.n297 PAD.n32 2.24164
R38777 PAD.n367 PAD.n43 2.24164
R38778 PAD.n305 PAD.n32 2.24164
R38779 PAD.n367 PAD.n42 2.24164
R38780 PAD.n309 PAD.n32 2.24164
R38781 PAD.n367 PAD.n41 2.24164
R38782 PAD.n317 PAD.n32 2.24164
R38783 PAD.n367 PAD.n40 2.24164
R38784 PAD.n321 PAD.n32 2.24164
R38785 PAD.n367 PAD.n39 2.24164
R38786 PAD.n329 PAD.n32 2.24164
R38787 PAD.n367 PAD.n38 2.24164
R38788 PAD.n333 PAD.n32 2.24164
R38789 PAD.n367 PAD.n37 2.24164
R38790 PAD.n341 PAD.n32 2.24164
R38791 PAD.n367 PAD.n36 2.24164
R38792 PAD.n345 PAD.n32 2.24164
R38793 PAD.n367 PAD.n35 2.24164
R38794 PAD.n353 PAD.n32 2.24164
R38795 PAD.n367 PAD.n34 2.24164
R38796 PAD.n357 PAD.n32 2.24164
R38797 PAD.n367 PAD.n33 2.24164
R38798 PAD.n365 PAD.n32 2.24164
R38799 PAD.n10692 PAD.n419 2.24164
R38800 PAD.n10716 PAD.n414 2.24164
R38801 PAD.n10416 PAD.n419 2.24164
R38802 PAD.n10716 PAD.n413 2.24164
R38803 PAD.n10685 PAD.n419 2.24164
R38804 PAD.n10716 PAD.n412 2.24164
R38805 PAD.n10421 PAD.n419 2.24164
R38806 PAD.n10716 PAD.n411 2.24164
R38807 PAD.n10676 PAD.n419 2.24164
R38808 PAD.n10716 PAD.n410 2.24164
R38809 PAD.n10426 PAD.n419 2.24164
R38810 PAD.n10716 PAD.n409 2.24164
R38811 PAD.n10667 PAD.n419 2.24164
R38812 PAD.n10716 PAD.n408 2.24164
R38813 PAD.n10431 PAD.n419 2.24164
R38814 PAD.n10716 PAD.n407 2.24164
R38815 PAD.n10658 PAD.n419 2.24164
R38816 PAD.n10716 PAD.n406 2.24164
R38817 PAD.n10436 PAD.n419 2.24164
R38818 PAD.n10716 PAD.n405 2.24164
R38819 PAD.n10649 PAD.n419 2.24164
R38820 PAD.n10716 PAD.n404 2.24164
R38821 PAD.n10441 PAD.n419 2.24164
R38822 PAD.n10716 PAD.n403 2.24164
R38823 PAD.n10640 PAD.n419 2.24164
R38824 PAD.n10716 PAD.n402 2.24164
R38825 PAD.n10446 PAD.n419 2.24164
R38826 PAD.n10716 PAD.n401 2.24164
R38827 PAD.n10631 PAD.n419 2.24164
R38828 PAD.n10716 PAD.n400 2.24164
R38829 PAD.n10451 PAD.n419 2.24164
R38830 PAD.n10716 PAD.n399 2.24164
R38831 PAD.n10622 PAD.n419 2.24164
R38832 PAD.n10716 PAD.n398 2.24164
R38833 PAD.n10456 PAD.n419 2.24164
R38834 PAD.n10716 PAD.n397 2.24164
R38835 PAD.n10613 PAD.n419 2.24164
R38836 PAD.n10716 PAD.n396 2.24164
R38837 PAD.n10461 PAD.n419 2.24164
R38838 PAD.n10716 PAD.n395 2.24164
R38839 PAD.n10604 PAD.n419 2.24164
R38840 PAD.n10716 PAD.n394 2.24164
R38841 PAD.n10466 PAD.n419 2.24164
R38842 PAD.n10716 PAD.n393 2.24164
R38843 PAD.n10595 PAD.n419 2.24164
R38844 PAD.n10716 PAD.n392 2.24164
R38845 PAD.n10471 PAD.n419 2.24164
R38846 PAD.n10716 PAD.n391 2.24164
R38847 PAD.n10586 PAD.n419 2.24164
R38848 PAD.n10716 PAD.n390 2.24164
R38849 PAD.n10476 PAD.n419 2.24164
R38850 PAD.n10716 PAD.n389 2.24164
R38851 PAD.n10577 PAD.n419 2.24164
R38852 PAD.n10716 PAD.n388 2.24164
R38853 PAD.n10481 PAD.n419 2.24164
R38854 PAD.n10716 PAD.n387 2.24164
R38855 PAD.n10568 PAD.n419 2.24164
R38856 PAD.n10716 PAD.n386 2.24164
R38857 PAD.n10486 PAD.n419 2.24164
R38858 PAD.n10716 PAD.n385 2.24164
R38859 PAD.n10559 PAD.n419 2.24164
R38860 PAD.n10716 PAD.n384 2.24164
R38861 PAD.n10491 PAD.n419 2.24164
R38862 PAD.n10716 PAD.n383 2.24164
R38863 PAD.n10550 PAD.n419 2.24164
R38864 PAD.n10716 PAD.n382 2.24164
R38865 PAD.n10496 PAD.n419 2.24164
R38866 PAD.n10716 PAD.n381 2.24164
R38867 PAD.n10541 PAD.n419 2.24164
R38868 PAD.n10716 PAD.n380 2.24164
R38869 PAD.n10501 PAD.n419 2.24164
R38870 PAD.n10716 PAD.n379 2.24164
R38871 PAD.n10532 PAD.n419 2.24164
R38872 PAD.n10716 PAD.n378 2.24164
R38873 PAD.n10506 PAD.n419 2.24164
R38874 PAD.n10716 PAD.n377 2.24164
R38875 PAD.n10523 PAD.n419 2.24164
R38876 PAD.n10716 PAD.n376 2.24164
R38877 PAD.n10511 PAD.n419 2.24164
R38878 PAD.n10716 PAD.n375 2.24164
R38879 PAD.n10514 PAD.n419 2.24164
R38880 PAD.n10716 PAD.n374 2.24164
R38881 PAD.n10714 PAD.n419 2.24164
R38882 PAD.n524 PAD.n433 2.24164
R38883 PAD.n526 PAD.n435 2.24164
R38884 PAD.n528 PAD.n433 2.24164
R38885 PAD.n517 PAD.n435 2.24164
R38886 PAD.n536 PAD.n433 2.24164
R38887 PAD.n538 PAD.n435 2.24164
R38888 PAD.n540 PAD.n433 2.24164
R38889 PAD.n513 PAD.n435 2.24164
R38890 PAD.n548 PAD.n433 2.24164
R38891 PAD.n550 PAD.n435 2.24164
R38892 PAD.n552 PAD.n433 2.24164
R38893 PAD.n509 PAD.n435 2.24164
R38894 PAD.n560 PAD.n433 2.24164
R38895 PAD.n562 PAD.n435 2.24164
R38896 PAD.n564 PAD.n433 2.24164
R38897 PAD.n505 PAD.n435 2.24164
R38898 PAD.n572 PAD.n433 2.24164
R38899 PAD.n574 PAD.n435 2.24164
R38900 PAD.n576 PAD.n433 2.24164
R38901 PAD.n501 PAD.n435 2.24164
R38902 PAD.n584 PAD.n433 2.24164
R38903 PAD.n586 PAD.n435 2.24164
R38904 PAD.n588 PAD.n433 2.24164
R38905 PAD.n497 PAD.n435 2.24164
R38906 PAD.n596 PAD.n433 2.24164
R38907 PAD.n598 PAD.n435 2.24164
R38908 PAD.n600 PAD.n433 2.24164
R38909 PAD.n493 PAD.n435 2.24164
R38910 PAD.n608 PAD.n433 2.24164
R38911 PAD.n610 PAD.n435 2.24164
R38912 PAD.n612 PAD.n433 2.24164
R38913 PAD.n489 PAD.n435 2.24164
R38914 PAD.n620 PAD.n433 2.24164
R38915 PAD.n622 PAD.n435 2.24164
R38916 PAD.n624 PAD.n433 2.24164
R38917 PAD.n485 PAD.n435 2.24164
R38918 PAD.n632 PAD.n433 2.24164
R38919 PAD.n634 PAD.n435 2.24164
R38920 PAD.n636 PAD.n433 2.24164
R38921 PAD.n481 PAD.n435 2.24164
R38922 PAD.n644 PAD.n433 2.24164
R38923 PAD.n646 PAD.n435 2.24164
R38924 PAD.n648 PAD.n433 2.24164
R38925 PAD.n477 PAD.n435 2.24164
R38926 PAD.n656 PAD.n433 2.24164
R38927 PAD.n658 PAD.n435 2.24164
R38928 PAD.n660 PAD.n433 2.24164
R38929 PAD.n473 PAD.n435 2.24164
R38930 PAD.n668 PAD.n433 2.24164
R38931 PAD.n670 PAD.n435 2.24164
R38932 PAD.n672 PAD.n433 2.24164
R38933 PAD.n469 PAD.n435 2.24164
R38934 PAD.n680 PAD.n433 2.24164
R38935 PAD.n682 PAD.n435 2.24164
R38936 PAD.n684 PAD.n433 2.24164
R38937 PAD.n465 PAD.n435 2.24164
R38938 PAD.n692 PAD.n433 2.24164
R38939 PAD.n694 PAD.n435 2.24164
R38940 PAD.n696 PAD.n433 2.24164
R38941 PAD.n461 PAD.n435 2.24164
R38942 PAD.n704 PAD.n433 2.24164
R38943 PAD.n706 PAD.n435 2.24164
R38944 PAD.n708 PAD.n433 2.24164
R38945 PAD.n457 PAD.n435 2.24164
R38946 PAD.n716 PAD.n433 2.24164
R38947 PAD.n718 PAD.n435 2.24164
R38948 PAD.n720 PAD.n433 2.24164
R38949 PAD.n453 PAD.n435 2.24164
R38950 PAD.n728 PAD.n433 2.24164
R38951 PAD.n730 PAD.n435 2.24164
R38952 PAD.n732 PAD.n433 2.24164
R38953 PAD.n449 PAD.n435 2.24164
R38954 PAD.n740 PAD.n433 2.24164
R38955 PAD.n742 PAD.n435 2.24164
R38956 PAD.n744 PAD.n433 2.24164
R38957 PAD.n445 PAD.n435 2.24164
R38958 PAD.n752 PAD.n433 2.24164
R38959 PAD.n754 PAD.n435 2.24164
R38960 PAD.n756 PAD.n433 2.24164
R38961 PAD.n441 PAD.n435 2.24164
R38962 PAD.n765 PAD.n433 2.24164
R38963 PAD.n767 PAD.n435 2.24164
R38964 PAD.n769 PAD.n433 2.24164
R38965 PAD.n869 PAD.n828 2.24164
R38966 PAD.n10388 PAD.n823 2.24164
R38967 PAD.n878 PAD.n828 2.24164
R38968 PAD.n10388 PAD.n822 2.24164
R38969 PAD.n882 PAD.n828 2.24164
R38970 PAD.n10388 PAD.n821 2.24164
R38971 PAD.n890 PAD.n828 2.24164
R38972 PAD.n10388 PAD.n820 2.24164
R38973 PAD.n894 PAD.n828 2.24164
R38974 PAD.n10388 PAD.n819 2.24164
R38975 PAD.n902 PAD.n828 2.24164
R38976 PAD.n10388 PAD.n818 2.24164
R38977 PAD.n906 PAD.n828 2.24164
R38978 PAD.n10388 PAD.n817 2.24164
R38979 PAD.n914 PAD.n828 2.24164
R38980 PAD.n10388 PAD.n816 2.24164
R38981 PAD.n918 PAD.n828 2.24164
R38982 PAD.n10388 PAD.n815 2.24164
R38983 PAD.n926 PAD.n828 2.24164
R38984 PAD.n10388 PAD.n814 2.24164
R38985 PAD.n930 PAD.n828 2.24164
R38986 PAD.n10388 PAD.n813 2.24164
R38987 PAD.n938 PAD.n828 2.24164
R38988 PAD.n10388 PAD.n812 2.24164
R38989 PAD.n942 PAD.n828 2.24164
R38990 PAD.n10388 PAD.n811 2.24164
R38991 PAD.n950 PAD.n828 2.24164
R38992 PAD.n10388 PAD.n810 2.24164
R38993 PAD.n954 PAD.n828 2.24164
R38994 PAD.n10388 PAD.n809 2.24164
R38995 PAD.n962 PAD.n828 2.24164
R38996 PAD.n10388 PAD.n808 2.24164
R38997 PAD.n966 PAD.n828 2.24164
R38998 PAD.n10388 PAD.n807 2.24164
R38999 PAD.n974 PAD.n828 2.24164
R39000 PAD.n10388 PAD.n806 2.24164
R39001 PAD.n978 PAD.n828 2.24164
R39002 PAD.n10388 PAD.n805 2.24164
R39003 PAD.n986 PAD.n828 2.24164
R39004 PAD.n10388 PAD.n804 2.24164
R39005 PAD.n990 PAD.n828 2.24164
R39006 PAD.n10388 PAD.n803 2.24164
R39007 PAD.n998 PAD.n828 2.24164
R39008 PAD.n10388 PAD.n802 2.24164
R39009 PAD.n1002 PAD.n828 2.24164
R39010 PAD.n10388 PAD.n801 2.24164
R39011 PAD.n1010 PAD.n828 2.24164
R39012 PAD.n10388 PAD.n800 2.24164
R39013 PAD.n1014 PAD.n828 2.24164
R39014 PAD.n10388 PAD.n799 2.24164
R39015 PAD.n1022 PAD.n828 2.24164
R39016 PAD.n10388 PAD.n798 2.24164
R39017 PAD.n1026 PAD.n828 2.24164
R39018 PAD.n10388 PAD.n797 2.24164
R39019 PAD.n1034 PAD.n828 2.24164
R39020 PAD.n10388 PAD.n796 2.24164
R39021 PAD.n1038 PAD.n828 2.24164
R39022 PAD.n10388 PAD.n795 2.24164
R39023 PAD.n1046 PAD.n828 2.24164
R39024 PAD.n10388 PAD.n794 2.24164
R39025 PAD.n1050 PAD.n828 2.24164
R39026 PAD.n10388 PAD.n793 2.24164
R39027 PAD.n1058 PAD.n828 2.24164
R39028 PAD.n10388 PAD.n792 2.24164
R39029 PAD.n1062 PAD.n828 2.24164
R39030 PAD.n10388 PAD.n791 2.24164
R39031 PAD.n1070 PAD.n828 2.24164
R39032 PAD.n10388 PAD.n790 2.24164
R39033 PAD.n1074 PAD.n828 2.24164
R39034 PAD.n10388 PAD.n789 2.24164
R39035 PAD.n1082 PAD.n828 2.24164
R39036 PAD.n10388 PAD.n788 2.24164
R39037 PAD.n1086 PAD.n828 2.24164
R39038 PAD.n10388 PAD.n787 2.24164
R39039 PAD.n1094 PAD.n828 2.24164
R39040 PAD.n10388 PAD.n786 2.24164
R39041 PAD.n1098 PAD.n828 2.24164
R39042 PAD.n10388 PAD.n785 2.24164
R39043 PAD.n1106 PAD.n828 2.24164
R39044 PAD.n10388 PAD.n784 2.24164
R39045 PAD.n1110 PAD.n828 2.24164
R39046 PAD.n10388 PAD.n783 2.24164
R39047 PAD.n10386 PAD.n828 2.24164
R39048 PAD.n10107 PAD.n1130 2.24164
R39049 PAD.n10109 PAD.n1132 2.24164
R39050 PAD.n10111 PAD.n1130 2.24164
R39051 PAD.n10101 PAD.n1132 2.24164
R39052 PAD.n10119 PAD.n1130 2.24164
R39053 PAD.n10121 PAD.n1132 2.24164
R39054 PAD.n10123 PAD.n1130 2.24164
R39055 PAD.n10097 PAD.n1132 2.24164
R39056 PAD.n10131 PAD.n1130 2.24164
R39057 PAD.n10133 PAD.n1132 2.24164
R39058 PAD.n10135 PAD.n1130 2.24164
R39059 PAD.n10093 PAD.n1132 2.24164
R39060 PAD.n10143 PAD.n1130 2.24164
R39061 PAD.n10145 PAD.n1132 2.24164
R39062 PAD.n10147 PAD.n1130 2.24164
R39063 PAD.n10089 PAD.n1132 2.24164
R39064 PAD.n10155 PAD.n1130 2.24164
R39065 PAD.n10157 PAD.n1132 2.24164
R39066 PAD.n10159 PAD.n1130 2.24164
R39067 PAD.n10085 PAD.n1132 2.24164
R39068 PAD.n10167 PAD.n1130 2.24164
R39069 PAD.n10169 PAD.n1132 2.24164
R39070 PAD.n10171 PAD.n1130 2.24164
R39071 PAD.n10081 PAD.n1132 2.24164
R39072 PAD.n10179 PAD.n1130 2.24164
R39073 PAD.n10181 PAD.n1132 2.24164
R39074 PAD.n10183 PAD.n1130 2.24164
R39075 PAD.n10077 PAD.n1132 2.24164
R39076 PAD.n10191 PAD.n1130 2.24164
R39077 PAD.n10193 PAD.n1132 2.24164
R39078 PAD.n10195 PAD.n1130 2.24164
R39079 PAD.n10073 PAD.n1132 2.24164
R39080 PAD.n10203 PAD.n1130 2.24164
R39081 PAD.n10205 PAD.n1132 2.24164
R39082 PAD.n10207 PAD.n1130 2.24164
R39083 PAD.n10069 PAD.n1132 2.24164
R39084 PAD.n10215 PAD.n1130 2.24164
R39085 PAD.n10217 PAD.n1132 2.24164
R39086 PAD.n10219 PAD.n1130 2.24164
R39087 PAD.n10065 PAD.n1132 2.24164
R39088 PAD.n10227 PAD.n1130 2.24164
R39089 PAD.n10229 PAD.n1132 2.24164
R39090 PAD.n10231 PAD.n1130 2.24164
R39091 PAD.n10061 PAD.n1132 2.24164
R39092 PAD.n10239 PAD.n1130 2.24164
R39093 PAD.n10241 PAD.n1132 2.24164
R39094 PAD.n10243 PAD.n1130 2.24164
R39095 PAD.n10057 PAD.n1132 2.24164
R39096 PAD.n10251 PAD.n1130 2.24164
R39097 PAD.n10253 PAD.n1132 2.24164
R39098 PAD.n10255 PAD.n1130 2.24164
R39099 PAD.n10053 PAD.n1132 2.24164
R39100 PAD.n10263 PAD.n1130 2.24164
R39101 PAD.n10265 PAD.n1132 2.24164
R39102 PAD.n10267 PAD.n1130 2.24164
R39103 PAD.n10049 PAD.n1132 2.24164
R39104 PAD.n10275 PAD.n1130 2.24164
R39105 PAD.n10277 PAD.n1132 2.24164
R39106 PAD.n10279 PAD.n1130 2.24164
R39107 PAD.n10045 PAD.n1132 2.24164
R39108 PAD.n10287 PAD.n1130 2.24164
R39109 PAD.n10289 PAD.n1132 2.24164
R39110 PAD.n10291 PAD.n1130 2.24164
R39111 PAD.n10041 PAD.n1132 2.24164
R39112 PAD.n10299 PAD.n1130 2.24164
R39113 PAD.n10301 PAD.n1132 2.24164
R39114 PAD.n10303 PAD.n1130 2.24164
R39115 PAD.n10037 PAD.n1132 2.24164
R39116 PAD.n10311 PAD.n1130 2.24164
R39117 PAD.n10313 PAD.n1132 2.24164
R39118 PAD.n10315 PAD.n1130 2.24164
R39119 PAD.n10033 PAD.n1132 2.24164
R39120 PAD.n10323 PAD.n1130 2.24164
R39121 PAD.n10325 PAD.n1132 2.24164
R39122 PAD.n10327 PAD.n1130 2.24164
R39123 PAD.n10029 PAD.n1132 2.24164
R39124 PAD.n10335 PAD.n1130 2.24164
R39125 PAD.n10337 PAD.n1132 2.24164
R39126 PAD.n10339 PAD.n1130 2.24164
R39127 PAD.n10025 PAD.n1132 2.24164
R39128 PAD.n10348 PAD.n1130 2.24164
R39129 PAD.n10350 PAD.n1132 2.24164
R39130 PAD.n10352 PAD.n1130 2.24164
R39131 PAD.n1483 PAD.n1482 2.24164
R39132 PAD.n1191 PAD.n1140 2.24164
R39133 PAD.n1483 PAD.n1189 2.24164
R39134 PAD.n1473 PAD.n1140 2.24164
R39135 PAD.n1483 PAD.n1188 2.24164
R39136 PAD.n1197 PAD.n1140 2.24164
R39137 PAD.n1483 PAD.n1187 2.24164
R39138 PAD.n1464 PAD.n1140 2.24164
R39139 PAD.n1483 PAD.n1186 2.24164
R39140 PAD.n1202 PAD.n1140 2.24164
R39141 PAD.n1483 PAD.n1185 2.24164
R39142 PAD.n1455 PAD.n1140 2.24164
R39143 PAD.n1483 PAD.n1184 2.24164
R39144 PAD.n1207 PAD.n1140 2.24164
R39145 PAD.n1483 PAD.n1183 2.24164
R39146 PAD.n1446 PAD.n1140 2.24164
R39147 PAD.n1483 PAD.n1182 2.24164
R39148 PAD.n1212 PAD.n1140 2.24164
R39149 PAD.n1483 PAD.n1181 2.24164
R39150 PAD.n1437 PAD.n1140 2.24164
R39151 PAD.n1483 PAD.n1180 2.24164
R39152 PAD.n1217 PAD.n1140 2.24164
R39153 PAD.n1483 PAD.n1179 2.24164
R39154 PAD.n1428 PAD.n1140 2.24164
R39155 PAD.n1483 PAD.n1178 2.24164
R39156 PAD.n1222 PAD.n1140 2.24164
R39157 PAD.n1483 PAD.n1177 2.24164
R39158 PAD.n1419 PAD.n1140 2.24164
R39159 PAD.n1483 PAD.n1176 2.24164
R39160 PAD.n1227 PAD.n1140 2.24164
R39161 PAD.n1483 PAD.n1175 2.24164
R39162 PAD.n1410 PAD.n1140 2.24164
R39163 PAD.n1483 PAD.n1174 2.24164
R39164 PAD.n1232 PAD.n1140 2.24164
R39165 PAD.n1483 PAD.n1173 2.24164
R39166 PAD.n1401 PAD.n1140 2.24164
R39167 PAD.n1483 PAD.n1172 2.24164
R39168 PAD.n1237 PAD.n1140 2.24164
R39169 PAD.n1483 PAD.n1171 2.24164
R39170 PAD.n1392 PAD.n1140 2.24164
R39171 PAD.n1483 PAD.n1170 2.24164
R39172 PAD.n1242 PAD.n1140 2.24164
R39173 PAD.n1483 PAD.n1169 2.24164
R39174 PAD.n1383 PAD.n1140 2.24164
R39175 PAD.n1483 PAD.n1168 2.24164
R39176 PAD.n1247 PAD.n1140 2.24164
R39177 PAD.n1483 PAD.n1167 2.24164
R39178 PAD.n1374 PAD.n1140 2.24164
R39179 PAD.n1483 PAD.n1166 2.24164
R39180 PAD.n1252 PAD.n1140 2.24164
R39181 PAD.n1483 PAD.n1165 2.24164
R39182 PAD.n1365 PAD.n1140 2.24164
R39183 PAD.n1483 PAD.n1164 2.24164
R39184 PAD.n1257 PAD.n1140 2.24164
R39185 PAD.n1483 PAD.n1163 2.24164
R39186 PAD.n1356 PAD.n1140 2.24164
R39187 PAD.n1483 PAD.n1162 2.24164
R39188 PAD.n1262 PAD.n1140 2.24164
R39189 PAD.n1483 PAD.n1161 2.24164
R39190 PAD.n1347 PAD.n1140 2.24164
R39191 PAD.n1483 PAD.n1160 2.24164
R39192 PAD.n1267 PAD.n1140 2.24164
R39193 PAD.n1483 PAD.n1159 2.24164
R39194 PAD.n1338 PAD.n1140 2.24164
R39195 PAD.n1483 PAD.n1158 2.24164
R39196 PAD.n1272 PAD.n1140 2.24164
R39197 PAD.n1483 PAD.n1157 2.24164
R39198 PAD.n1329 PAD.n1140 2.24164
R39199 PAD.n1483 PAD.n1156 2.24164
R39200 PAD.n1277 PAD.n1140 2.24164
R39201 PAD.n1483 PAD.n1155 2.24164
R39202 PAD.n1320 PAD.n1140 2.24164
R39203 PAD.n1483 PAD.n1154 2.24164
R39204 PAD.n1282 PAD.n1140 2.24164
R39205 PAD.n1483 PAD.n1153 2.24164
R39206 PAD.n1311 PAD.n1140 2.24164
R39207 PAD.n1483 PAD.n1152 2.24164
R39208 PAD.n1287 PAD.n1140 2.24164
R39209 PAD.n1483 PAD.n1151 2.24164
R39210 PAD.n1302 PAD.n1140 2.24164
R39211 PAD.n1483 PAD.n1150 2.24164
R39212 PAD.n1292 PAD.n1140 2.24164
R39213 PAD.n1483 PAD.n1149 2.24164
R39214 PAD.n1577 PAD.n1536 2.24164
R39215 PAD.n9998 PAD.n1530 2.24164
R39216 PAD.n9755 PAD.n1536 2.24164
R39217 PAD.n9998 PAD.n1529 2.24164
R39218 PAD.n9759 PAD.n1536 2.24164
R39219 PAD.n9998 PAD.n1528 2.24164
R39220 PAD.n9767 PAD.n1536 2.24164
R39221 PAD.n9998 PAD.n1527 2.24164
R39222 PAD.n9771 PAD.n1536 2.24164
R39223 PAD.n9998 PAD.n1526 2.24164
R39224 PAD.n9779 PAD.n1536 2.24164
R39225 PAD.n9998 PAD.n1525 2.24164
R39226 PAD.n9783 PAD.n1536 2.24164
R39227 PAD.n9998 PAD.n1524 2.24164
R39228 PAD.n9791 PAD.n1536 2.24164
R39229 PAD.n9998 PAD.n1523 2.24164
R39230 PAD.n9795 PAD.n1536 2.24164
R39231 PAD.n9998 PAD.n1522 2.24164
R39232 PAD.n9803 PAD.n1536 2.24164
R39233 PAD.n9998 PAD.n1521 2.24164
R39234 PAD.n9807 PAD.n1536 2.24164
R39235 PAD.n9998 PAD.n1520 2.24164
R39236 PAD.n9815 PAD.n1536 2.24164
R39237 PAD.n9998 PAD.n1519 2.24164
R39238 PAD.n9819 PAD.n1536 2.24164
R39239 PAD.n9998 PAD.n1518 2.24164
R39240 PAD.n9827 PAD.n1536 2.24164
R39241 PAD.n9998 PAD.n1517 2.24164
R39242 PAD.n9831 PAD.n1536 2.24164
R39243 PAD.n9998 PAD.n1516 2.24164
R39244 PAD.n9839 PAD.n1536 2.24164
R39245 PAD.n9998 PAD.n1515 2.24164
R39246 PAD.n9843 PAD.n1536 2.24164
R39247 PAD.n9998 PAD.n1514 2.24164
R39248 PAD.n9851 PAD.n1536 2.24164
R39249 PAD.n9998 PAD.n1513 2.24164
R39250 PAD.n9855 PAD.n1536 2.24164
R39251 PAD.n9998 PAD.n1512 2.24164
R39252 PAD.n9863 PAD.n1536 2.24164
R39253 PAD.n9998 PAD.n1511 2.24164
R39254 PAD.n9867 PAD.n1536 2.24164
R39255 PAD.n9998 PAD.n1510 2.24164
R39256 PAD.n9875 PAD.n1536 2.24164
R39257 PAD.n9998 PAD.n1509 2.24164
R39258 PAD.n9879 PAD.n1536 2.24164
R39259 PAD.n9998 PAD.n1508 2.24164
R39260 PAD.n9887 PAD.n1536 2.24164
R39261 PAD.n9998 PAD.n1507 2.24164
R39262 PAD.n9891 PAD.n1536 2.24164
R39263 PAD.n9998 PAD.n1506 2.24164
R39264 PAD.n9899 PAD.n1536 2.24164
R39265 PAD.n9998 PAD.n1505 2.24164
R39266 PAD.n9903 PAD.n1536 2.24164
R39267 PAD.n9998 PAD.n1504 2.24164
R39268 PAD.n9911 PAD.n1536 2.24164
R39269 PAD.n9998 PAD.n1503 2.24164
R39270 PAD.n9915 PAD.n1536 2.24164
R39271 PAD.n9998 PAD.n1502 2.24164
R39272 PAD.n9923 PAD.n1536 2.24164
R39273 PAD.n9998 PAD.n1501 2.24164
R39274 PAD.n9927 PAD.n1536 2.24164
R39275 PAD.n9998 PAD.n1500 2.24164
R39276 PAD.n9935 PAD.n1536 2.24164
R39277 PAD.n9998 PAD.n1499 2.24164
R39278 PAD.n9939 PAD.n1536 2.24164
R39279 PAD.n9998 PAD.n1498 2.24164
R39280 PAD.n9947 PAD.n1536 2.24164
R39281 PAD.n9998 PAD.n1497 2.24164
R39282 PAD.n9951 PAD.n1536 2.24164
R39283 PAD.n9998 PAD.n1496 2.24164
R39284 PAD.n9959 PAD.n1536 2.24164
R39285 PAD.n9998 PAD.n1495 2.24164
R39286 PAD.n9963 PAD.n1536 2.24164
R39287 PAD.n9998 PAD.n1494 2.24164
R39288 PAD.n9971 PAD.n1536 2.24164
R39289 PAD.n9998 PAD.n1493 2.24164
R39290 PAD.n9975 PAD.n1536 2.24164
R39291 PAD.n9998 PAD.n1492 2.24164
R39292 PAD.n9983 PAD.n1536 2.24164
R39293 PAD.n9998 PAD.n1491 2.24164
R39294 PAD.n9987 PAD.n1536 2.24164
R39295 PAD.n9998 PAD.n1490 2.24164
R39296 PAD.n9996 PAD.n1536 2.24164
R39297 PAD.n1601 PAD.n1592 2.24164
R39298 PAD.n1928 PAD.n1594 2.24164
R39299 PAD.n1926 PAD.n1592 2.24164
R39300 PAD.n1602 PAD.n1594 2.24164
R39301 PAD.n1918 PAD.n1592 2.24164
R39302 PAD.n1916 PAD.n1594 2.24164
R39303 PAD.n1914 PAD.n1592 2.24164
R39304 PAD.n1607 PAD.n1594 2.24164
R39305 PAD.n1906 PAD.n1592 2.24164
R39306 PAD.n1904 PAD.n1594 2.24164
R39307 PAD.n1902 PAD.n1592 2.24164
R39308 PAD.n1611 PAD.n1594 2.24164
R39309 PAD.n1894 PAD.n1592 2.24164
R39310 PAD.n1892 PAD.n1594 2.24164
R39311 PAD.n1890 PAD.n1592 2.24164
R39312 PAD.n1615 PAD.n1594 2.24164
R39313 PAD.n1882 PAD.n1592 2.24164
R39314 PAD.n1880 PAD.n1594 2.24164
R39315 PAD.n1878 PAD.n1592 2.24164
R39316 PAD.n1619 PAD.n1594 2.24164
R39317 PAD.n1870 PAD.n1592 2.24164
R39318 PAD.n1868 PAD.n1594 2.24164
R39319 PAD.n1866 PAD.n1592 2.24164
R39320 PAD.n1623 PAD.n1594 2.24164
R39321 PAD.n1858 PAD.n1592 2.24164
R39322 PAD.n1856 PAD.n1594 2.24164
R39323 PAD.n1854 PAD.n1592 2.24164
R39324 PAD.n1627 PAD.n1594 2.24164
R39325 PAD.n1846 PAD.n1592 2.24164
R39326 PAD.n1844 PAD.n1594 2.24164
R39327 PAD.n1842 PAD.n1592 2.24164
R39328 PAD.n1631 PAD.n1594 2.24164
R39329 PAD.n1834 PAD.n1592 2.24164
R39330 PAD.n1832 PAD.n1594 2.24164
R39331 PAD.n1830 PAD.n1592 2.24164
R39332 PAD.n1635 PAD.n1594 2.24164
R39333 PAD.n1822 PAD.n1592 2.24164
R39334 PAD.n1820 PAD.n1594 2.24164
R39335 PAD.n1818 PAD.n1592 2.24164
R39336 PAD.n1639 PAD.n1594 2.24164
R39337 PAD.n1810 PAD.n1592 2.24164
R39338 PAD.n1808 PAD.n1594 2.24164
R39339 PAD.n1806 PAD.n1592 2.24164
R39340 PAD.n1643 PAD.n1594 2.24164
R39341 PAD.n1798 PAD.n1592 2.24164
R39342 PAD.n1796 PAD.n1594 2.24164
R39343 PAD.n1794 PAD.n1592 2.24164
R39344 PAD.n1647 PAD.n1594 2.24164
R39345 PAD.n1786 PAD.n1592 2.24164
R39346 PAD.n1784 PAD.n1594 2.24164
R39347 PAD.n1782 PAD.n1592 2.24164
R39348 PAD.n1651 PAD.n1594 2.24164
R39349 PAD.n1774 PAD.n1592 2.24164
R39350 PAD.n1772 PAD.n1594 2.24164
R39351 PAD.n1770 PAD.n1592 2.24164
R39352 PAD.n1655 PAD.n1594 2.24164
R39353 PAD.n1762 PAD.n1592 2.24164
R39354 PAD.n1760 PAD.n1594 2.24164
R39355 PAD.n1758 PAD.n1592 2.24164
R39356 PAD.n1659 PAD.n1594 2.24164
R39357 PAD.n1750 PAD.n1592 2.24164
R39358 PAD.n1748 PAD.n1594 2.24164
R39359 PAD.n1746 PAD.n1592 2.24164
R39360 PAD.n1663 PAD.n1594 2.24164
R39361 PAD.n1738 PAD.n1592 2.24164
R39362 PAD.n1736 PAD.n1594 2.24164
R39363 PAD.n1734 PAD.n1592 2.24164
R39364 PAD.n1667 PAD.n1594 2.24164
R39365 PAD.n1726 PAD.n1592 2.24164
R39366 PAD.n1724 PAD.n1594 2.24164
R39367 PAD.n1722 PAD.n1592 2.24164
R39368 PAD.n1671 PAD.n1594 2.24164
R39369 PAD.n1714 PAD.n1592 2.24164
R39370 PAD.n1712 PAD.n1594 2.24164
R39371 PAD.n1710 PAD.n1592 2.24164
R39372 PAD.n1675 PAD.n1594 2.24164
R39373 PAD.n1702 PAD.n1592 2.24164
R39374 PAD.n1700 PAD.n1594 2.24164
R39375 PAD.n1698 PAD.n1592 2.24164
R39376 PAD.n1679 PAD.n1594 2.24164
R39377 PAD.n1690 PAD.n1592 2.24164
R39378 PAD.n1688 PAD.n1594 2.24164
R39379 PAD.n1686 PAD.n1592 2.24164
R39380 PAD.n2029 PAD.n1988 2.24164
R39381 PAD.n9712 PAD.n1983 2.24164
R39382 PAD.n9469 PAD.n1988 2.24164
R39383 PAD.n9712 PAD.n1982 2.24164
R39384 PAD.n9473 PAD.n1988 2.24164
R39385 PAD.n9712 PAD.n1981 2.24164
R39386 PAD.n9481 PAD.n1988 2.24164
R39387 PAD.n9712 PAD.n1980 2.24164
R39388 PAD.n9485 PAD.n1988 2.24164
R39389 PAD.n9712 PAD.n1979 2.24164
R39390 PAD.n9493 PAD.n1988 2.24164
R39391 PAD.n9712 PAD.n1978 2.24164
R39392 PAD.n9497 PAD.n1988 2.24164
R39393 PAD.n9712 PAD.n1977 2.24164
R39394 PAD.n9505 PAD.n1988 2.24164
R39395 PAD.n9712 PAD.n1976 2.24164
R39396 PAD.n9509 PAD.n1988 2.24164
R39397 PAD.n9712 PAD.n1975 2.24164
R39398 PAD.n9517 PAD.n1988 2.24164
R39399 PAD.n9712 PAD.n1974 2.24164
R39400 PAD.n9521 PAD.n1988 2.24164
R39401 PAD.n9712 PAD.n1973 2.24164
R39402 PAD.n9529 PAD.n1988 2.24164
R39403 PAD.n9712 PAD.n1972 2.24164
R39404 PAD.n9533 PAD.n1988 2.24164
R39405 PAD.n9712 PAD.n1971 2.24164
R39406 PAD.n9541 PAD.n1988 2.24164
R39407 PAD.n9712 PAD.n1970 2.24164
R39408 PAD.n9545 PAD.n1988 2.24164
R39409 PAD.n9712 PAD.n1969 2.24164
R39410 PAD.n9553 PAD.n1988 2.24164
R39411 PAD.n9712 PAD.n1968 2.24164
R39412 PAD.n9557 PAD.n1988 2.24164
R39413 PAD.n9712 PAD.n1967 2.24164
R39414 PAD.n9565 PAD.n1988 2.24164
R39415 PAD.n9712 PAD.n1966 2.24164
R39416 PAD.n9569 PAD.n1988 2.24164
R39417 PAD.n9712 PAD.n1965 2.24164
R39418 PAD.n9577 PAD.n1988 2.24164
R39419 PAD.n9712 PAD.n1964 2.24164
R39420 PAD.n9581 PAD.n1988 2.24164
R39421 PAD.n9712 PAD.n1963 2.24164
R39422 PAD.n9589 PAD.n1988 2.24164
R39423 PAD.n9712 PAD.n1962 2.24164
R39424 PAD.n9593 PAD.n1988 2.24164
R39425 PAD.n9712 PAD.n1961 2.24164
R39426 PAD.n9601 PAD.n1988 2.24164
R39427 PAD.n9712 PAD.n1960 2.24164
R39428 PAD.n9605 PAD.n1988 2.24164
R39429 PAD.n9712 PAD.n1959 2.24164
R39430 PAD.n9613 PAD.n1988 2.24164
R39431 PAD.n9712 PAD.n1958 2.24164
R39432 PAD.n9617 PAD.n1988 2.24164
R39433 PAD.n9712 PAD.n1957 2.24164
R39434 PAD.n9625 PAD.n1988 2.24164
R39435 PAD.n9712 PAD.n1956 2.24164
R39436 PAD.n9629 PAD.n1988 2.24164
R39437 PAD.n9712 PAD.n1955 2.24164
R39438 PAD.n9637 PAD.n1988 2.24164
R39439 PAD.n9712 PAD.n1954 2.24164
R39440 PAD.n9641 PAD.n1988 2.24164
R39441 PAD.n9712 PAD.n1953 2.24164
R39442 PAD.n9649 PAD.n1988 2.24164
R39443 PAD.n9712 PAD.n1952 2.24164
R39444 PAD.n9653 PAD.n1988 2.24164
R39445 PAD.n9712 PAD.n1951 2.24164
R39446 PAD.n9661 PAD.n1988 2.24164
R39447 PAD.n9712 PAD.n1950 2.24164
R39448 PAD.n9665 PAD.n1988 2.24164
R39449 PAD.n9712 PAD.n1949 2.24164
R39450 PAD.n9673 PAD.n1988 2.24164
R39451 PAD.n9712 PAD.n1948 2.24164
R39452 PAD.n9677 PAD.n1988 2.24164
R39453 PAD.n9712 PAD.n1947 2.24164
R39454 PAD.n9685 PAD.n1988 2.24164
R39455 PAD.n9712 PAD.n1946 2.24164
R39456 PAD.n9689 PAD.n1988 2.24164
R39457 PAD.n9712 PAD.n1945 2.24164
R39458 PAD.n9697 PAD.n1988 2.24164
R39459 PAD.n9712 PAD.n1944 2.24164
R39460 PAD.n9701 PAD.n1988 2.24164
R39461 PAD.n9712 PAD.n1943 2.24164
R39462 PAD.n9710 PAD.n1988 2.24164
R39463 PAD.n2132 PAD.n2091 2.24164
R39464 PAD.n9445 PAD.n2087 2.24164
R39465 PAD.n9203 PAD.n2091 2.24164
R39466 PAD.n9445 PAD.n2086 2.24164
R39467 PAD.n9207 PAD.n2091 2.24164
R39468 PAD.n9445 PAD.n2085 2.24164
R39469 PAD.n9215 PAD.n2091 2.24164
R39470 PAD.n9445 PAD.n2084 2.24164
R39471 PAD.n9219 PAD.n2091 2.24164
R39472 PAD.n9445 PAD.n2083 2.24164
R39473 PAD.n9227 PAD.n2091 2.24164
R39474 PAD.n9445 PAD.n2082 2.24164
R39475 PAD.n9231 PAD.n2091 2.24164
R39476 PAD.n9445 PAD.n2081 2.24164
R39477 PAD.n9239 PAD.n2091 2.24164
R39478 PAD.n9445 PAD.n2080 2.24164
R39479 PAD.n9243 PAD.n2091 2.24164
R39480 PAD.n9445 PAD.n2079 2.24164
R39481 PAD.n9251 PAD.n2091 2.24164
R39482 PAD.n9445 PAD.n2078 2.24164
R39483 PAD.n9255 PAD.n2091 2.24164
R39484 PAD.n9445 PAD.n2077 2.24164
R39485 PAD.n9263 PAD.n2091 2.24164
R39486 PAD.n9445 PAD.n2076 2.24164
R39487 PAD.n9267 PAD.n2091 2.24164
R39488 PAD.n9445 PAD.n2075 2.24164
R39489 PAD.n9275 PAD.n2091 2.24164
R39490 PAD.n9445 PAD.n2074 2.24164
R39491 PAD.n9279 PAD.n2091 2.24164
R39492 PAD.n9445 PAD.n2073 2.24164
R39493 PAD.n9287 PAD.n2091 2.24164
R39494 PAD.n9445 PAD.n2072 2.24164
R39495 PAD.n9291 PAD.n2091 2.24164
R39496 PAD.n9445 PAD.n2071 2.24164
R39497 PAD.n9299 PAD.n2091 2.24164
R39498 PAD.n9445 PAD.n2070 2.24164
R39499 PAD.n9303 PAD.n2091 2.24164
R39500 PAD.n9445 PAD.n2069 2.24164
R39501 PAD.n9311 PAD.n2091 2.24164
R39502 PAD.n9445 PAD.n2068 2.24164
R39503 PAD.n9315 PAD.n2091 2.24164
R39504 PAD.n9445 PAD.n2067 2.24164
R39505 PAD.n9323 PAD.n2091 2.24164
R39506 PAD.n9445 PAD.n2066 2.24164
R39507 PAD.n9327 PAD.n2091 2.24164
R39508 PAD.n9445 PAD.n2065 2.24164
R39509 PAD.n9335 PAD.n2091 2.24164
R39510 PAD.n9445 PAD.n2064 2.24164
R39511 PAD.n9339 PAD.n2091 2.24164
R39512 PAD.n9445 PAD.n2063 2.24164
R39513 PAD.n9347 PAD.n2091 2.24164
R39514 PAD.n9445 PAD.n2062 2.24164
R39515 PAD.n9351 PAD.n2091 2.24164
R39516 PAD.n9445 PAD.n2061 2.24164
R39517 PAD.n9359 PAD.n2091 2.24164
R39518 PAD.n9445 PAD.n2060 2.24164
R39519 PAD.n9363 PAD.n2091 2.24164
R39520 PAD.n9445 PAD.n2059 2.24164
R39521 PAD.n9371 PAD.n2091 2.24164
R39522 PAD.n9445 PAD.n2058 2.24164
R39523 PAD.n9375 PAD.n2091 2.24164
R39524 PAD.n9445 PAD.n2057 2.24164
R39525 PAD.n9383 PAD.n2091 2.24164
R39526 PAD.n9445 PAD.n2056 2.24164
R39527 PAD.n9387 PAD.n2091 2.24164
R39528 PAD.n9445 PAD.n2055 2.24164
R39529 PAD.n9395 PAD.n2091 2.24164
R39530 PAD.n9445 PAD.n2054 2.24164
R39531 PAD.n9399 PAD.n2091 2.24164
R39532 PAD.n9445 PAD.n2053 2.24164
R39533 PAD.n9407 PAD.n2091 2.24164
R39534 PAD.n9445 PAD.n2052 2.24164
R39535 PAD.n9411 PAD.n2091 2.24164
R39536 PAD.n9445 PAD.n2051 2.24164
R39537 PAD.n9419 PAD.n2091 2.24164
R39538 PAD.n9445 PAD.n2050 2.24164
R39539 PAD.n9423 PAD.n2091 2.24164
R39540 PAD.n9445 PAD.n2049 2.24164
R39541 PAD.n9431 PAD.n2091 2.24164
R39542 PAD.n9445 PAD.n2048 2.24164
R39543 PAD.n9435 PAD.n2091 2.24164
R39544 PAD.n9445 PAD.n2047 2.24164
R39545 PAD.n9443 PAD.n2091 2.24164
R39546 PAD.n2153 PAD.n2146 2.24164
R39547 PAD.n2479 PAD.n2139 2.24164
R39548 PAD.n2477 PAD.n2146 2.24164
R39549 PAD.n2154 PAD.n2139 2.24164
R39550 PAD.n2469 PAD.n2146 2.24164
R39551 PAD.n2467 PAD.n2139 2.24164
R39552 PAD.n2465 PAD.n2146 2.24164
R39553 PAD.n2159 PAD.n2139 2.24164
R39554 PAD.n2457 PAD.n2146 2.24164
R39555 PAD.n2455 PAD.n2139 2.24164
R39556 PAD.n2453 PAD.n2146 2.24164
R39557 PAD.n2163 PAD.n2139 2.24164
R39558 PAD.n2445 PAD.n2146 2.24164
R39559 PAD.n2443 PAD.n2139 2.24164
R39560 PAD.n2441 PAD.n2146 2.24164
R39561 PAD.n2167 PAD.n2139 2.24164
R39562 PAD.n2433 PAD.n2146 2.24164
R39563 PAD.n2431 PAD.n2139 2.24164
R39564 PAD.n2429 PAD.n2146 2.24164
R39565 PAD.n2171 PAD.n2139 2.24164
R39566 PAD.n2421 PAD.n2146 2.24164
R39567 PAD.n2419 PAD.n2139 2.24164
R39568 PAD.n2417 PAD.n2146 2.24164
R39569 PAD.n2175 PAD.n2139 2.24164
R39570 PAD.n2409 PAD.n2146 2.24164
R39571 PAD.n2407 PAD.n2139 2.24164
R39572 PAD.n2405 PAD.n2146 2.24164
R39573 PAD.n2179 PAD.n2139 2.24164
R39574 PAD.n2397 PAD.n2146 2.24164
R39575 PAD.n2395 PAD.n2139 2.24164
R39576 PAD.n2393 PAD.n2146 2.24164
R39577 PAD.n2183 PAD.n2139 2.24164
R39578 PAD.n2385 PAD.n2146 2.24164
R39579 PAD.n2383 PAD.n2139 2.24164
R39580 PAD.n2381 PAD.n2146 2.24164
R39581 PAD.n2187 PAD.n2139 2.24164
R39582 PAD.n2373 PAD.n2146 2.24164
R39583 PAD.n2371 PAD.n2139 2.24164
R39584 PAD.n2369 PAD.n2146 2.24164
R39585 PAD.n2191 PAD.n2139 2.24164
R39586 PAD.n2361 PAD.n2146 2.24164
R39587 PAD.n2359 PAD.n2139 2.24164
R39588 PAD.n2357 PAD.n2146 2.24164
R39589 PAD.n2195 PAD.n2139 2.24164
R39590 PAD.n2349 PAD.n2146 2.24164
R39591 PAD.n2347 PAD.n2139 2.24164
R39592 PAD.n2345 PAD.n2146 2.24164
R39593 PAD.n2199 PAD.n2139 2.24164
R39594 PAD.n2337 PAD.n2146 2.24164
R39595 PAD.n2335 PAD.n2139 2.24164
R39596 PAD.n2333 PAD.n2146 2.24164
R39597 PAD.n2203 PAD.n2139 2.24164
R39598 PAD.n2325 PAD.n2146 2.24164
R39599 PAD.n2323 PAD.n2139 2.24164
R39600 PAD.n2321 PAD.n2146 2.24164
R39601 PAD.n2207 PAD.n2139 2.24164
R39602 PAD.n2313 PAD.n2146 2.24164
R39603 PAD.n2311 PAD.n2139 2.24164
R39604 PAD.n2309 PAD.n2146 2.24164
R39605 PAD.n2211 PAD.n2139 2.24164
R39606 PAD.n2301 PAD.n2146 2.24164
R39607 PAD.n2299 PAD.n2139 2.24164
R39608 PAD.n2297 PAD.n2146 2.24164
R39609 PAD.n2215 PAD.n2139 2.24164
R39610 PAD.n2289 PAD.n2146 2.24164
R39611 PAD.n2287 PAD.n2139 2.24164
R39612 PAD.n2285 PAD.n2146 2.24164
R39613 PAD.n2219 PAD.n2139 2.24164
R39614 PAD.n2277 PAD.n2146 2.24164
R39615 PAD.n2275 PAD.n2139 2.24164
R39616 PAD.n2273 PAD.n2146 2.24164
R39617 PAD.n2223 PAD.n2139 2.24164
R39618 PAD.n2265 PAD.n2146 2.24164
R39619 PAD.n2263 PAD.n2139 2.24164
R39620 PAD.n2261 PAD.n2146 2.24164
R39621 PAD.n2227 PAD.n2139 2.24164
R39622 PAD.n2253 PAD.n2146 2.24164
R39623 PAD.n2251 PAD.n2139 2.24164
R39624 PAD.n2249 PAD.n2146 2.24164
R39625 PAD.n2231 PAD.n2139 2.24164
R39626 PAD.n2241 PAD.n2146 2.24164
R39627 PAD.n2239 PAD.n2139 2.24164
R39628 PAD.n2237 PAD.n2146 2.24164
R39629 PAD.n2500 PAD.n2494 2.24164
R39630 PAD.n2826 PAD.n2487 2.24164
R39631 PAD.n2824 PAD.n2494 2.24164
R39632 PAD.n2501 PAD.n2487 2.24164
R39633 PAD.n2816 PAD.n2494 2.24164
R39634 PAD.n2814 PAD.n2487 2.24164
R39635 PAD.n2812 PAD.n2494 2.24164
R39636 PAD.n2506 PAD.n2487 2.24164
R39637 PAD.n2804 PAD.n2494 2.24164
R39638 PAD.n2802 PAD.n2487 2.24164
R39639 PAD.n2800 PAD.n2494 2.24164
R39640 PAD.n2510 PAD.n2487 2.24164
R39641 PAD.n2792 PAD.n2494 2.24164
R39642 PAD.n2790 PAD.n2487 2.24164
R39643 PAD.n2788 PAD.n2494 2.24164
R39644 PAD.n2514 PAD.n2487 2.24164
R39645 PAD.n2780 PAD.n2494 2.24164
R39646 PAD.n2778 PAD.n2487 2.24164
R39647 PAD.n2776 PAD.n2494 2.24164
R39648 PAD.n2518 PAD.n2487 2.24164
R39649 PAD.n2768 PAD.n2494 2.24164
R39650 PAD.n2766 PAD.n2487 2.24164
R39651 PAD.n2764 PAD.n2494 2.24164
R39652 PAD.n2522 PAD.n2487 2.24164
R39653 PAD.n2756 PAD.n2494 2.24164
R39654 PAD.n2754 PAD.n2487 2.24164
R39655 PAD.n2752 PAD.n2494 2.24164
R39656 PAD.n2526 PAD.n2487 2.24164
R39657 PAD.n2744 PAD.n2494 2.24164
R39658 PAD.n2742 PAD.n2487 2.24164
R39659 PAD.n2740 PAD.n2494 2.24164
R39660 PAD.n2530 PAD.n2487 2.24164
R39661 PAD.n2732 PAD.n2494 2.24164
R39662 PAD.n2730 PAD.n2487 2.24164
R39663 PAD.n2728 PAD.n2494 2.24164
R39664 PAD.n2534 PAD.n2487 2.24164
R39665 PAD.n2720 PAD.n2494 2.24164
R39666 PAD.n2718 PAD.n2487 2.24164
R39667 PAD.n2716 PAD.n2494 2.24164
R39668 PAD.n2538 PAD.n2487 2.24164
R39669 PAD.n2708 PAD.n2494 2.24164
R39670 PAD.n2706 PAD.n2487 2.24164
R39671 PAD.n2704 PAD.n2494 2.24164
R39672 PAD.n2542 PAD.n2487 2.24164
R39673 PAD.n2696 PAD.n2494 2.24164
R39674 PAD.n2694 PAD.n2487 2.24164
R39675 PAD.n2692 PAD.n2494 2.24164
R39676 PAD.n2546 PAD.n2487 2.24164
R39677 PAD.n2684 PAD.n2494 2.24164
R39678 PAD.n2682 PAD.n2487 2.24164
R39679 PAD.n2680 PAD.n2494 2.24164
R39680 PAD.n2550 PAD.n2487 2.24164
R39681 PAD.n2672 PAD.n2494 2.24164
R39682 PAD.n2670 PAD.n2487 2.24164
R39683 PAD.n2668 PAD.n2494 2.24164
R39684 PAD.n2554 PAD.n2487 2.24164
R39685 PAD.n2660 PAD.n2494 2.24164
R39686 PAD.n2658 PAD.n2487 2.24164
R39687 PAD.n2656 PAD.n2494 2.24164
R39688 PAD.n2558 PAD.n2487 2.24164
R39689 PAD.n2648 PAD.n2494 2.24164
R39690 PAD.n2646 PAD.n2487 2.24164
R39691 PAD.n2644 PAD.n2494 2.24164
R39692 PAD.n2562 PAD.n2487 2.24164
R39693 PAD.n2636 PAD.n2494 2.24164
R39694 PAD.n2634 PAD.n2487 2.24164
R39695 PAD.n2632 PAD.n2494 2.24164
R39696 PAD.n2566 PAD.n2487 2.24164
R39697 PAD.n2624 PAD.n2494 2.24164
R39698 PAD.n2622 PAD.n2487 2.24164
R39699 PAD.n2620 PAD.n2494 2.24164
R39700 PAD.n2570 PAD.n2487 2.24164
R39701 PAD.n2612 PAD.n2494 2.24164
R39702 PAD.n2610 PAD.n2487 2.24164
R39703 PAD.n2608 PAD.n2494 2.24164
R39704 PAD.n2574 PAD.n2487 2.24164
R39705 PAD.n2600 PAD.n2494 2.24164
R39706 PAD.n2598 PAD.n2487 2.24164
R39707 PAD.n2596 PAD.n2494 2.24164
R39708 PAD.n2578 PAD.n2487 2.24164
R39709 PAD.n2588 PAD.n2494 2.24164
R39710 PAD.n2586 PAD.n2487 2.24164
R39711 PAD.n2584 PAD.n2494 2.24164
R39712 PAD.n9116 PAD.n2879 2.24164
R39713 PAD.n9140 PAD.n2875 2.24164
R39714 PAD.n8840 PAD.n2879 2.24164
R39715 PAD.n9140 PAD.n2874 2.24164
R39716 PAD.n9109 PAD.n2879 2.24164
R39717 PAD.n9140 PAD.n2873 2.24164
R39718 PAD.n8845 PAD.n2879 2.24164
R39719 PAD.n9140 PAD.n2872 2.24164
R39720 PAD.n9100 PAD.n2879 2.24164
R39721 PAD.n9140 PAD.n2871 2.24164
R39722 PAD.n8850 PAD.n2879 2.24164
R39723 PAD.n9140 PAD.n2870 2.24164
R39724 PAD.n9091 PAD.n2879 2.24164
R39725 PAD.n9140 PAD.n2869 2.24164
R39726 PAD.n8855 PAD.n2879 2.24164
R39727 PAD.n9140 PAD.n2868 2.24164
R39728 PAD.n9082 PAD.n2879 2.24164
R39729 PAD.n9140 PAD.n2867 2.24164
R39730 PAD.n8860 PAD.n2879 2.24164
R39731 PAD.n9140 PAD.n2866 2.24164
R39732 PAD.n9073 PAD.n2879 2.24164
R39733 PAD.n9140 PAD.n2865 2.24164
R39734 PAD.n8865 PAD.n2879 2.24164
R39735 PAD.n9140 PAD.n2864 2.24164
R39736 PAD.n9064 PAD.n2879 2.24164
R39737 PAD.n9140 PAD.n2863 2.24164
R39738 PAD.n8870 PAD.n2879 2.24164
R39739 PAD.n9140 PAD.n2862 2.24164
R39740 PAD.n9055 PAD.n2879 2.24164
R39741 PAD.n9140 PAD.n2861 2.24164
R39742 PAD.n8875 PAD.n2879 2.24164
R39743 PAD.n9140 PAD.n2860 2.24164
R39744 PAD.n9046 PAD.n2879 2.24164
R39745 PAD.n9140 PAD.n2859 2.24164
R39746 PAD.n8880 PAD.n2879 2.24164
R39747 PAD.n9140 PAD.n2858 2.24164
R39748 PAD.n9037 PAD.n2879 2.24164
R39749 PAD.n9140 PAD.n2857 2.24164
R39750 PAD.n8885 PAD.n2879 2.24164
R39751 PAD.n9140 PAD.n2856 2.24164
R39752 PAD.n9028 PAD.n2879 2.24164
R39753 PAD.n9140 PAD.n2855 2.24164
R39754 PAD.n8890 PAD.n2879 2.24164
R39755 PAD.n9140 PAD.n2854 2.24164
R39756 PAD.n9019 PAD.n2879 2.24164
R39757 PAD.n9140 PAD.n2853 2.24164
R39758 PAD.n8895 PAD.n2879 2.24164
R39759 PAD.n9140 PAD.n2852 2.24164
R39760 PAD.n9010 PAD.n2879 2.24164
R39761 PAD.n9140 PAD.n2851 2.24164
R39762 PAD.n8900 PAD.n2879 2.24164
R39763 PAD.n9140 PAD.n2850 2.24164
R39764 PAD.n9001 PAD.n2879 2.24164
R39765 PAD.n9140 PAD.n2849 2.24164
R39766 PAD.n8905 PAD.n2879 2.24164
R39767 PAD.n9140 PAD.n2848 2.24164
R39768 PAD.n8992 PAD.n2879 2.24164
R39769 PAD.n9140 PAD.n2847 2.24164
R39770 PAD.n8910 PAD.n2879 2.24164
R39771 PAD.n9140 PAD.n2846 2.24164
R39772 PAD.n8983 PAD.n2879 2.24164
R39773 PAD.n9140 PAD.n2845 2.24164
R39774 PAD.n8915 PAD.n2879 2.24164
R39775 PAD.n9140 PAD.n2844 2.24164
R39776 PAD.n8974 PAD.n2879 2.24164
R39777 PAD.n9140 PAD.n2843 2.24164
R39778 PAD.n8920 PAD.n2879 2.24164
R39779 PAD.n9140 PAD.n2842 2.24164
R39780 PAD.n8965 PAD.n2879 2.24164
R39781 PAD.n9140 PAD.n2841 2.24164
R39782 PAD.n8925 PAD.n2879 2.24164
R39783 PAD.n9140 PAD.n2840 2.24164
R39784 PAD.n8956 PAD.n2879 2.24164
R39785 PAD.n9140 PAD.n2839 2.24164
R39786 PAD.n8930 PAD.n2879 2.24164
R39787 PAD.n9140 PAD.n2838 2.24164
R39788 PAD.n8947 PAD.n2879 2.24164
R39789 PAD.n9140 PAD.n2837 2.24164
R39790 PAD.n8935 PAD.n2879 2.24164
R39791 PAD.n9140 PAD.n2836 2.24164
R39792 PAD.n8938 PAD.n2879 2.24164
R39793 PAD.n9140 PAD.n2835 2.24164
R39794 PAD.n9138 PAD.n2879 2.24164
R39795 PAD.n8821 PAD.n8820 2.24164
R39796 PAD.n8812 PAD.n2891 2.24164
R39797 PAD.n8821 PAD.n2945 2.24164
R39798 PAD.n8809 PAD.n2891 2.24164
R39799 PAD.n8821 PAD.n2944 2.24164
R39800 PAD.n8801 PAD.n2891 2.24164
R39801 PAD.n8821 PAD.n2943 2.24164
R39802 PAD.n8797 PAD.n2891 2.24164
R39803 PAD.n8821 PAD.n2942 2.24164
R39804 PAD.n8789 PAD.n2891 2.24164
R39805 PAD.n8821 PAD.n2941 2.24164
R39806 PAD.n8785 PAD.n2891 2.24164
R39807 PAD.n8821 PAD.n2940 2.24164
R39808 PAD.n8777 PAD.n2891 2.24164
R39809 PAD.n8821 PAD.n2939 2.24164
R39810 PAD.n8773 PAD.n2891 2.24164
R39811 PAD.n8821 PAD.n2938 2.24164
R39812 PAD.n8765 PAD.n2891 2.24164
R39813 PAD.n8821 PAD.n2937 2.24164
R39814 PAD.n8761 PAD.n2891 2.24164
R39815 PAD.n8821 PAD.n2936 2.24164
R39816 PAD.n8753 PAD.n2891 2.24164
R39817 PAD.n8821 PAD.n2935 2.24164
R39818 PAD.n8749 PAD.n2891 2.24164
R39819 PAD.n8821 PAD.n2934 2.24164
R39820 PAD.n8741 PAD.n2891 2.24164
R39821 PAD.n8821 PAD.n2933 2.24164
R39822 PAD.n8737 PAD.n2891 2.24164
R39823 PAD.n8821 PAD.n2932 2.24164
R39824 PAD.n8729 PAD.n2891 2.24164
R39825 PAD.n8821 PAD.n2931 2.24164
R39826 PAD.n8725 PAD.n2891 2.24164
R39827 PAD.n8821 PAD.n2930 2.24164
R39828 PAD.n8717 PAD.n2891 2.24164
R39829 PAD.n8821 PAD.n2929 2.24164
R39830 PAD.n8713 PAD.n2891 2.24164
R39831 PAD.n8821 PAD.n2928 2.24164
R39832 PAD.n8705 PAD.n2891 2.24164
R39833 PAD.n8821 PAD.n2927 2.24164
R39834 PAD.n8701 PAD.n2891 2.24164
R39835 PAD.n8821 PAD.n2926 2.24164
R39836 PAD.n8693 PAD.n2891 2.24164
R39837 PAD.n8821 PAD.n2925 2.24164
R39838 PAD.n8689 PAD.n2891 2.24164
R39839 PAD.n8821 PAD.n2924 2.24164
R39840 PAD.n8681 PAD.n2891 2.24164
R39841 PAD.n8821 PAD.n2923 2.24164
R39842 PAD.n8677 PAD.n2891 2.24164
R39843 PAD.n8821 PAD.n2922 2.24164
R39844 PAD.n8669 PAD.n2891 2.24164
R39845 PAD.n8821 PAD.n2921 2.24164
R39846 PAD.n8665 PAD.n2891 2.24164
R39847 PAD.n8821 PAD.n2920 2.24164
R39848 PAD.n8657 PAD.n2891 2.24164
R39849 PAD.n8821 PAD.n2919 2.24164
R39850 PAD.n8653 PAD.n2891 2.24164
R39851 PAD.n8821 PAD.n2918 2.24164
R39852 PAD.n8645 PAD.n2891 2.24164
R39853 PAD.n8821 PAD.n2917 2.24164
R39854 PAD.n8641 PAD.n2891 2.24164
R39855 PAD.n8821 PAD.n2916 2.24164
R39856 PAD.n8633 PAD.n2891 2.24164
R39857 PAD.n8821 PAD.n2915 2.24164
R39858 PAD.n8629 PAD.n2891 2.24164
R39859 PAD.n8821 PAD.n2914 2.24164
R39860 PAD.n8621 PAD.n2891 2.24164
R39861 PAD.n8821 PAD.n2913 2.24164
R39862 PAD.n8617 PAD.n2891 2.24164
R39863 PAD.n8821 PAD.n2912 2.24164
R39864 PAD.n8609 PAD.n2891 2.24164
R39865 PAD.n8821 PAD.n2911 2.24164
R39866 PAD.n8605 PAD.n2891 2.24164
R39867 PAD.n8821 PAD.n2910 2.24164
R39868 PAD.n8597 PAD.n2891 2.24164
R39869 PAD.n8821 PAD.n2909 2.24164
R39870 PAD.n8593 PAD.n2891 2.24164
R39871 PAD.n8821 PAD.n2908 2.24164
R39872 PAD.n8585 PAD.n2891 2.24164
R39873 PAD.n8821 PAD.n2907 2.24164
R39874 PAD.n8581 PAD.n2891 2.24164
R39875 PAD.n8821 PAD.n2906 2.24164
R39876 PAD.n8573 PAD.n2891 2.24164
R39877 PAD.n8821 PAD.n2905 2.24164
R39878 PAD.n3038 PAD.n2997 2.24164
R39879 PAD.n8517 PAD.n2993 2.24164
R39880 PAD.n3047 PAD.n2997 2.24164
R39881 PAD.n8517 PAD.n2992 2.24164
R39882 PAD.n3051 PAD.n2997 2.24164
R39883 PAD.n8517 PAD.n2991 2.24164
R39884 PAD.n3059 PAD.n2997 2.24164
R39885 PAD.n8517 PAD.n2990 2.24164
R39886 PAD.n3063 PAD.n2997 2.24164
R39887 PAD.n8517 PAD.n2989 2.24164
R39888 PAD.n3071 PAD.n2997 2.24164
R39889 PAD.n8517 PAD.n2988 2.24164
R39890 PAD.n3075 PAD.n2997 2.24164
R39891 PAD.n8517 PAD.n2987 2.24164
R39892 PAD.n3083 PAD.n2997 2.24164
R39893 PAD.n8517 PAD.n2986 2.24164
R39894 PAD.n3087 PAD.n2997 2.24164
R39895 PAD.n8517 PAD.n2985 2.24164
R39896 PAD.n3095 PAD.n2997 2.24164
R39897 PAD.n8517 PAD.n2984 2.24164
R39898 PAD.n3099 PAD.n2997 2.24164
R39899 PAD.n8517 PAD.n2983 2.24164
R39900 PAD.n3107 PAD.n2997 2.24164
R39901 PAD.n8517 PAD.n2982 2.24164
R39902 PAD.n3111 PAD.n2997 2.24164
R39903 PAD.n8517 PAD.n2981 2.24164
R39904 PAD.n3119 PAD.n2997 2.24164
R39905 PAD.n8517 PAD.n2980 2.24164
R39906 PAD.n3123 PAD.n2997 2.24164
R39907 PAD.n8517 PAD.n2979 2.24164
R39908 PAD.n3131 PAD.n2997 2.24164
R39909 PAD.n8517 PAD.n2978 2.24164
R39910 PAD.n3135 PAD.n2997 2.24164
R39911 PAD.n8517 PAD.n2977 2.24164
R39912 PAD.n3143 PAD.n2997 2.24164
R39913 PAD.n8517 PAD.n2976 2.24164
R39914 PAD.n3147 PAD.n2997 2.24164
R39915 PAD.n8517 PAD.n2975 2.24164
R39916 PAD.n3155 PAD.n2997 2.24164
R39917 PAD.n8517 PAD.n2974 2.24164
R39918 PAD.n3159 PAD.n2997 2.24164
R39919 PAD.n8517 PAD.n2973 2.24164
R39920 PAD.n3167 PAD.n2997 2.24164
R39921 PAD.n8517 PAD.n2972 2.24164
R39922 PAD.n3171 PAD.n2997 2.24164
R39923 PAD.n8517 PAD.n2971 2.24164
R39924 PAD.n3179 PAD.n2997 2.24164
R39925 PAD.n8517 PAD.n2970 2.24164
R39926 PAD.n3183 PAD.n2997 2.24164
R39927 PAD.n8517 PAD.n2969 2.24164
R39928 PAD.n3191 PAD.n2997 2.24164
R39929 PAD.n8517 PAD.n2968 2.24164
R39930 PAD.n3195 PAD.n2997 2.24164
R39931 PAD.n8517 PAD.n2967 2.24164
R39932 PAD.n3203 PAD.n2997 2.24164
R39933 PAD.n8517 PAD.n2966 2.24164
R39934 PAD.n3207 PAD.n2997 2.24164
R39935 PAD.n8517 PAD.n2965 2.24164
R39936 PAD.n3215 PAD.n2997 2.24164
R39937 PAD.n8517 PAD.n2964 2.24164
R39938 PAD.n3219 PAD.n2997 2.24164
R39939 PAD.n8517 PAD.n2963 2.24164
R39940 PAD.n3227 PAD.n2997 2.24164
R39941 PAD.n8517 PAD.n2962 2.24164
R39942 PAD.n3231 PAD.n2997 2.24164
R39943 PAD.n8517 PAD.n2961 2.24164
R39944 PAD.n3239 PAD.n2997 2.24164
R39945 PAD.n8517 PAD.n2960 2.24164
R39946 PAD.n3243 PAD.n2997 2.24164
R39947 PAD.n8517 PAD.n2959 2.24164
R39948 PAD.n3251 PAD.n2997 2.24164
R39949 PAD.n8517 PAD.n2958 2.24164
R39950 PAD.n3255 PAD.n2997 2.24164
R39951 PAD.n8517 PAD.n2957 2.24164
R39952 PAD.n3263 PAD.n2997 2.24164
R39953 PAD.n8517 PAD.n2956 2.24164
R39954 PAD.n3267 PAD.n2997 2.24164
R39955 PAD.n8517 PAD.n2955 2.24164
R39956 PAD.n3275 PAD.n2997 2.24164
R39957 PAD.n8517 PAD.n2954 2.24164
R39958 PAD.n3279 PAD.n2997 2.24164
R39959 PAD.n8517 PAD.n2953 2.24164
R39960 PAD.n8515 PAD.n2997 2.24164
R39961 PAD.n3383 PAD.n3342 2.24164
R39962 PAD.n8492 PAD.n3337 2.24164
R39963 PAD.n3392 PAD.n3342 2.24164
R39964 PAD.n8492 PAD.n3336 2.24164
R39965 PAD.n3396 PAD.n3342 2.24164
R39966 PAD.n8492 PAD.n3335 2.24164
R39967 PAD.n3404 PAD.n3342 2.24164
R39968 PAD.n8492 PAD.n3334 2.24164
R39969 PAD.n3408 PAD.n3342 2.24164
R39970 PAD.n8492 PAD.n3333 2.24164
R39971 PAD.n3416 PAD.n3342 2.24164
R39972 PAD.n8492 PAD.n3332 2.24164
R39973 PAD.n3420 PAD.n3342 2.24164
R39974 PAD.n8492 PAD.n3331 2.24164
R39975 PAD.n3428 PAD.n3342 2.24164
R39976 PAD.n8492 PAD.n3330 2.24164
R39977 PAD.n3432 PAD.n3342 2.24164
R39978 PAD.n8492 PAD.n3329 2.24164
R39979 PAD.n3440 PAD.n3342 2.24164
R39980 PAD.n8492 PAD.n3328 2.24164
R39981 PAD.n3444 PAD.n3342 2.24164
R39982 PAD.n8492 PAD.n3327 2.24164
R39983 PAD.n3452 PAD.n3342 2.24164
R39984 PAD.n8492 PAD.n3326 2.24164
R39985 PAD.n3456 PAD.n3342 2.24164
R39986 PAD.n8492 PAD.n3325 2.24164
R39987 PAD.n3464 PAD.n3342 2.24164
R39988 PAD.n8492 PAD.n3324 2.24164
R39989 PAD.n3468 PAD.n3342 2.24164
R39990 PAD.n8492 PAD.n3323 2.24164
R39991 PAD.n3476 PAD.n3342 2.24164
R39992 PAD.n8492 PAD.n3322 2.24164
R39993 PAD.n3480 PAD.n3342 2.24164
R39994 PAD.n8492 PAD.n3321 2.24164
R39995 PAD.n3488 PAD.n3342 2.24164
R39996 PAD.n8492 PAD.n3320 2.24164
R39997 PAD.n3492 PAD.n3342 2.24164
R39998 PAD.n8492 PAD.n3319 2.24164
R39999 PAD.n3500 PAD.n3342 2.24164
R40000 PAD.n8492 PAD.n3318 2.24164
R40001 PAD.n3504 PAD.n3342 2.24164
R40002 PAD.n8492 PAD.n3317 2.24164
R40003 PAD.n3512 PAD.n3342 2.24164
R40004 PAD.n8492 PAD.n3316 2.24164
R40005 PAD.n3516 PAD.n3342 2.24164
R40006 PAD.n8492 PAD.n3315 2.24164
R40007 PAD.n3524 PAD.n3342 2.24164
R40008 PAD.n8492 PAD.n3314 2.24164
R40009 PAD.n3528 PAD.n3342 2.24164
R40010 PAD.n8492 PAD.n3313 2.24164
R40011 PAD.n3536 PAD.n3342 2.24164
R40012 PAD.n8492 PAD.n3312 2.24164
R40013 PAD.n3540 PAD.n3342 2.24164
R40014 PAD.n8492 PAD.n3311 2.24164
R40015 PAD.n3548 PAD.n3342 2.24164
R40016 PAD.n8492 PAD.n3310 2.24164
R40017 PAD.n3552 PAD.n3342 2.24164
R40018 PAD.n8492 PAD.n3309 2.24164
R40019 PAD.n3560 PAD.n3342 2.24164
R40020 PAD.n8492 PAD.n3308 2.24164
R40021 PAD.n3564 PAD.n3342 2.24164
R40022 PAD.n8492 PAD.n3307 2.24164
R40023 PAD.n3572 PAD.n3342 2.24164
R40024 PAD.n8492 PAD.n3306 2.24164
R40025 PAD.n3576 PAD.n3342 2.24164
R40026 PAD.n8492 PAD.n3305 2.24164
R40027 PAD.n3584 PAD.n3342 2.24164
R40028 PAD.n8492 PAD.n3304 2.24164
R40029 PAD.n3588 PAD.n3342 2.24164
R40030 PAD.n8492 PAD.n3303 2.24164
R40031 PAD.n3596 PAD.n3342 2.24164
R40032 PAD.n8492 PAD.n3302 2.24164
R40033 PAD.n3600 PAD.n3342 2.24164
R40034 PAD.n8492 PAD.n3301 2.24164
R40035 PAD.n3608 PAD.n3342 2.24164
R40036 PAD.n8492 PAD.n3300 2.24164
R40037 PAD.n3612 PAD.n3342 2.24164
R40038 PAD.n8492 PAD.n3299 2.24164
R40039 PAD.n3620 PAD.n3342 2.24164
R40040 PAD.n8492 PAD.n3298 2.24164
R40041 PAD.n3624 PAD.n3342 2.24164
R40042 PAD.n8492 PAD.n3297 2.24164
R40043 PAD.n8490 PAD.n3342 2.24164
R40044 PAD.n3728 PAD.n3687 2.24164
R40045 PAD.n8468 PAD.n3682 2.24164
R40046 PAD.n3737 PAD.n3687 2.24164
R40047 PAD.n8468 PAD.n3681 2.24164
R40048 PAD.n3741 PAD.n3687 2.24164
R40049 PAD.n8468 PAD.n3680 2.24164
R40050 PAD.n3749 PAD.n3687 2.24164
R40051 PAD.n8468 PAD.n3679 2.24164
R40052 PAD.n3753 PAD.n3687 2.24164
R40053 PAD.n8468 PAD.n3678 2.24164
R40054 PAD.n3761 PAD.n3687 2.24164
R40055 PAD.n8468 PAD.n3677 2.24164
R40056 PAD.n3765 PAD.n3687 2.24164
R40057 PAD.n8468 PAD.n3676 2.24164
R40058 PAD.n3773 PAD.n3687 2.24164
R40059 PAD.n8468 PAD.n3675 2.24164
R40060 PAD.n3777 PAD.n3687 2.24164
R40061 PAD.n8468 PAD.n3674 2.24164
R40062 PAD.n3785 PAD.n3687 2.24164
R40063 PAD.n8468 PAD.n3673 2.24164
R40064 PAD.n3789 PAD.n3687 2.24164
R40065 PAD.n8468 PAD.n3672 2.24164
R40066 PAD.n3797 PAD.n3687 2.24164
R40067 PAD.n8468 PAD.n3671 2.24164
R40068 PAD.n3801 PAD.n3687 2.24164
R40069 PAD.n8468 PAD.n3670 2.24164
R40070 PAD.n3809 PAD.n3687 2.24164
R40071 PAD.n8468 PAD.n3669 2.24164
R40072 PAD.n3813 PAD.n3687 2.24164
R40073 PAD.n8468 PAD.n3668 2.24164
R40074 PAD.n3821 PAD.n3687 2.24164
R40075 PAD.n8468 PAD.n3667 2.24164
R40076 PAD.n3825 PAD.n3687 2.24164
R40077 PAD.n8468 PAD.n3666 2.24164
R40078 PAD.n3833 PAD.n3687 2.24164
R40079 PAD.n8468 PAD.n3665 2.24164
R40080 PAD.n3837 PAD.n3687 2.24164
R40081 PAD.n8468 PAD.n3664 2.24164
R40082 PAD.n3845 PAD.n3687 2.24164
R40083 PAD.n8468 PAD.n3663 2.24164
R40084 PAD.n3849 PAD.n3687 2.24164
R40085 PAD.n8468 PAD.n3662 2.24164
R40086 PAD.n3857 PAD.n3687 2.24164
R40087 PAD.n8468 PAD.n3661 2.24164
R40088 PAD.n3861 PAD.n3687 2.24164
R40089 PAD.n8468 PAD.n3660 2.24164
R40090 PAD.n3869 PAD.n3687 2.24164
R40091 PAD.n8468 PAD.n3659 2.24164
R40092 PAD.n3873 PAD.n3687 2.24164
R40093 PAD.n8468 PAD.n3658 2.24164
R40094 PAD.n3881 PAD.n3687 2.24164
R40095 PAD.n8468 PAD.n3657 2.24164
R40096 PAD.n3885 PAD.n3687 2.24164
R40097 PAD.n8468 PAD.n3656 2.24164
R40098 PAD.n3893 PAD.n3687 2.24164
R40099 PAD.n8468 PAD.n3655 2.24164
R40100 PAD.n3897 PAD.n3687 2.24164
R40101 PAD.n8468 PAD.n3654 2.24164
R40102 PAD.n3905 PAD.n3687 2.24164
R40103 PAD.n8468 PAD.n3653 2.24164
R40104 PAD.n3909 PAD.n3687 2.24164
R40105 PAD.n8468 PAD.n3652 2.24164
R40106 PAD.n3917 PAD.n3687 2.24164
R40107 PAD.n8468 PAD.n3651 2.24164
R40108 PAD.n3921 PAD.n3687 2.24164
R40109 PAD.n8468 PAD.n3650 2.24164
R40110 PAD.n3929 PAD.n3687 2.24164
R40111 PAD.n8468 PAD.n3649 2.24164
R40112 PAD.n3933 PAD.n3687 2.24164
R40113 PAD.n8468 PAD.n3648 2.24164
R40114 PAD.n3941 PAD.n3687 2.24164
R40115 PAD.n8468 PAD.n3647 2.24164
R40116 PAD.n3945 PAD.n3687 2.24164
R40117 PAD.n8468 PAD.n3646 2.24164
R40118 PAD.n3953 PAD.n3687 2.24164
R40119 PAD.n8468 PAD.n3645 2.24164
R40120 PAD.n3957 PAD.n3687 2.24164
R40121 PAD.n8468 PAD.n3644 2.24164
R40122 PAD.n3965 PAD.n3687 2.24164
R40123 PAD.n8468 PAD.n3643 2.24164
R40124 PAD.n3969 PAD.n3687 2.24164
R40125 PAD.n8468 PAD.n3642 2.24164
R40126 PAD.n8466 PAD.n3687 2.24164
R40127 PAD.n4069 PAD.n4028 2.24164
R40128 PAD.n8444 PAD.n4024 2.24164
R40129 PAD.n4078 PAD.n4028 2.24164
R40130 PAD.n8444 PAD.n4023 2.24164
R40131 PAD.n4082 PAD.n4028 2.24164
R40132 PAD.n8444 PAD.n4022 2.24164
R40133 PAD.n4090 PAD.n4028 2.24164
R40134 PAD.n8444 PAD.n4021 2.24164
R40135 PAD.n4094 PAD.n4028 2.24164
R40136 PAD.n8444 PAD.n4020 2.24164
R40137 PAD.n4102 PAD.n4028 2.24164
R40138 PAD.n8444 PAD.n4019 2.24164
R40139 PAD.n4106 PAD.n4028 2.24164
R40140 PAD.n8444 PAD.n4018 2.24164
R40141 PAD.n4114 PAD.n4028 2.24164
R40142 PAD.n8444 PAD.n4017 2.24164
R40143 PAD.n4118 PAD.n4028 2.24164
R40144 PAD.n8444 PAD.n4016 2.24164
R40145 PAD.n4126 PAD.n4028 2.24164
R40146 PAD.n8444 PAD.n4015 2.24164
R40147 PAD.n4130 PAD.n4028 2.24164
R40148 PAD.n8444 PAD.n4014 2.24164
R40149 PAD.n4138 PAD.n4028 2.24164
R40150 PAD.n8444 PAD.n4013 2.24164
R40151 PAD.n4142 PAD.n4028 2.24164
R40152 PAD.n8444 PAD.n4012 2.24164
R40153 PAD.n4150 PAD.n4028 2.24164
R40154 PAD.n8444 PAD.n4011 2.24164
R40155 PAD.n4154 PAD.n4028 2.24164
R40156 PAD.n8444 PAD.n4010 2.24164
R40157 PAD.n4162 PAD.n4028 2.24164
R40158 PAD.n8444 PAD.n4009 2.24164
R40159 PAD.n4166 PAD.n4028 2.24164
R40160 PAD.n8444 PAD.n4008 2.24164
R40161 PAD.n4174 PAD.n4028 2.24164
R40162 PAD.n8444 PAD.n4007 2.24164
R40163 PAD.n4178 PAD.n4028 2.24164
R40164 PAD.n8444 PAD.n4006 2.24164
R40165 PAD.n4186 PAD.n4028 2.24164
R40166 PAD.n8444 PAD.n4005 2.24164
R40167 PAD.n4190 PAD.n4028 2.24164
R40168 PAD.n8444 PAD.n4004 2.24164
R40169 PAD.n4198 PAD.n4028 2.24164
R40170 PAD.n8444 PAD.n4003 2.24164
R40171 PAD.n4202 PAD.n4028 2.24164
R40172 PAD.n8444 PAD.n4002 2.24164
R40173 PAD.n4210 PAD.n4028 2.24164
R40174 PAD.n8444 PAD.n4001 2.24164
R40175 PAD.n4214 PAD.n4028 2.24164
R40176 PAD.n8444 PAD.n4000 2.24164
R40177 PAD.n4222 PAD.n4028 2.24164
R40178 PAD.n8444 PAD.n3999 2.24164
R40179 PAD.n4226 PAD.n4028 2.24164
R40180 PAD.n8444 PAD.n3998 2.24164
R40181 PAD.n4234 PAD.n4028 2.24164
R40182 PAD.n8444 PAD.n3997 2.24164
R40183 PAD.n4238 PAD.n4028 2.24164
R40184 PAD.n8444 PAD.n3996 2.24164
R40185 PAD.n4246 PAD.n4028 2.24164
R40186 PAD.n8444 PAD.n3995 2.24164
R40187 PAD.n4250 PAD.n4028 2.24164
R40188 PAD.n8444 PAD.n3994 2.24164
R40189 PAD.n4258 PAD.n4028 2.24164
R40190 PAD.n8444 PAD.n3993 2.24164
R40191 PAD.n4262 PAD.n4028 2.24164
R40192 PAD.n8444 PAD.n3992 2.24164
R40193 PAD.n4270 PAD.n4028 2.24164
R40194 PAD.n8444 PAD.n3991 2.24164
R40195 PAD.n4274 PAD.n4028 2.24164
R40196 PAD.n8444 PAD.n3990 2.24164
R40197 PAD.n4282 PAD.n4028 2.24164
R40198 PAD.n8444 PAD.n3989 2.24164
R40199 PAD.n4286 PAD.n4028 2.24164
R40200 PAD.n8444 PAD.n3988 2.24164
R40201 PAD.n4294 PAD.n4028 2.24164
R40202 PAD.n8444 PAD.n3987 2.24164
R40203 PAD.n4298 PAD.n4028 2.24164
R40204 PAD.n8444 PAD.n3986 2.24164
R40205 PAD.n4306 PAD.n4028 2.24164
R40206 PAD.n8444 PAD.n3985 2.24164
R40207 PAD.n4310 PAD.n4028 2.24164
R40208 PAD.n8444 PAD.n3984 2.24164
R40209 PAD.n8442 PAD.n4028 2.24164
R40210 PAD.n4421 PAD.n4331 2.24164
R40211 PAD.n4423 PAD.n4333 2.24164
R40212 PAD.n4425 PAD.n4331 2.24164
R40213 PAD.n4415 PAD.n4333 2.24164
R40214 PAD.n4433 PAD.n4331 2.24164
R40215 PAD.n4435 PAD.n4333 2.24164
R40216 PAD.n4437 PAD.n4331 2.24164
R40217 PAD.n4411 PAD.n4333 2.24164
R40218 PAD.n4445 PAD.n4331 2.24164
R40219 PAD.n4447 PAD.n4333 2.24164
R40220 PAD.n4449 PAD.n4331 2.24164
R40221 PAD.n4407 PAD.n4333 2.24164
R40222 PAD.n4457 PAD.n4331 2.24164
R40223 PAD.n4459 PAD.n4333 2.24164
R40224 PAD.n4461 PAD.n4331 2.24164
R40225 PAD.n4403 PAD.n4333 2.24164
R40226 PAD.n4469 PAD.n4331 2.24164
R40227 PAD.n4471 PAD.n4333 2.24164
R40228 PAD.n4473 PAD.n4331 2.24164
R40229 PAD.n4399 PAD.n4333 2.24164
R40230 PAD.n4481 PAD.n4331 2.24164
R40231 PAD.n4483 PAD.n4333 2.24164
R40232 PAD.n4485 PAD.n4331 2.24164
R40233 PAD.n4395 PAD.n4333 2.24164
R40234 PAD.n4493 PAD.n4331 2.24164
R40235 PAD.n4495 PAD.n4333 2.24164
R40236 PAD.n4497 PAD.n4331 2.24164
R40237 PAD.n4391 PAD.n4333 2.24164
R40238 PAD.n4505 PAD.n4331 2.24164
R40239 PAD.n4507 PAD.n4333 2.24164
R40240 PAD.n4509 PAD.n4331 2.24164
R40241 PAD.n4387 PAD.n4333 2.24164
R40242 PAD.n4517 PAD.n4331 2.24164
R40243 PAD.n4519 PAD.n4333 2.24164
R40244 PAD.n4521 PAD.n4331 2.24164
R40245 PAD.n4383 PAD.n4333 2.24164
R40246 PAD.n4529 PAD.n4331 2.24164
R40247 PAD.n4531 PAD.n4333 2.24164
R40248 PAD.n4533 PAD.n4331 2.24164
R40249 PAD.n4379 PAD.n4333 2.24164
R40250 PAD.n4541 PAD.n4331 2.24164
R40251 PAD.n4543 PAD.n4333 2.24164
R40252 PAD.n4545 PAD.n4331 2.24164
R40253 PAD.n4375 PAD.n4333 2.24164
R40254 PAD.n4553 PAD.n4331 2.24164
R40255 PAD.n4555 PAD.n4333 2.24164
R40256 PAD.n4557 PAD.n4331 2.24164
R40257 PAD.n4371 PAD.n4333 2.24164
R40258 PAD.n4565 PAD.n4331 2.24164
R40259 PAD.n4567 PAD.n4333 2.24164
R40260 PAD.n4569 PAD.n4331 2.24164
R40261 PAD.n4367 PAD.n4333 2.24164
R40262 PAD.n4577 PAD.n4331 2.24164
R40263 PAD.n4579 PAD.n4333 2.24164
R40264 PAD.n4581 PAD.n4331 2.24164
R40265 PAD.n4363 PAD.n4333 2.24164
R40266 PAD.n4589 PAD.n4331 2.24164
R40267 PAD.n4591 PAD.n4333 2.24164
R40268 PAD.n4593 PAD.n4331 2.24164
R40269 PAD.n4359 PAD.n4333 2.24164
R40270 PAD.n4601 PAD.n4331 2.24164
R40271 PAD.n4603 PAD.n4333 2.24164
R40272 PAD.n4605 PAD.n4331 2.24164
R40273 PAD.n4355 PAD.n4333 2.24164
R40274 PAD.n4613 PAD.n4331 2.24164
R40275 PAD.n4615 PAD.n4333 2.24164
R40276 PAD.n4617 PAD.n4331 2.24164
R40277 PAD.n4351 PAD.n4333 2.24164
R40278 PAD.n4625 PAD.n4331 2.24164
R40279 PAD.n4627 PAD.n4333 2.24164
R40280 PAD.n4629 PAD.n4331 2.24164
R40281 PAD.n4347 PAD.n4333 2.24164
R40282 PAD.n4637 PAD.n4331 2.24164
R40283 PAD.n4639 PAD.n4333 2.24164
R40284 PAD.n4641 PAD.n4331 2.24164
R40285 PAD.n4343 PAD.n4333 2.24164
R40286 PAD.n4649 PAD.n4331 2.24164
R40287 PAD.n4651 PAD.n4333 2.24164
R40288 PAD.n4653 PAD.n4331 2.24164
R40289 PAD.n4339 PAD.n4333 2.24164
R40290 PAD.n4662 PAD.n4331 2.24164
R40291 PAD.n4664 PAD.n4333 2.24164
R40292 PAD.n4666 PAD.n4331 2.24164
R40293 PAD.n8397 PAD.n8396 2.24164
R40294 PAD.n4726 PAD.n4673 2.24164
R40295 PAD.n8397 PAD.n4723 2.24164
R40296 PAD.n8387 PAD.n4673 2.24164
R40297 PAD.n8397 PAD.n4722 2.24164
R40298 PAD.n4732 PAD.n4673 2.24164
R40299 PAD.n8397 PAD.n4721 2.24164
R40300 PAD.n8378 PAD.n4673 2.24164
R40301 PAD.n8397 PAD.n4720 2.24164
R40302 PAD.n4737 PAD.n4673 2.24164
R40303 PAD.n8397 PAD.n4719 2.24164
R40304 PAD.n8369 PAD.n4673 2.24164
R40305 PAD.n8397 PAD.n4718 2.24164
R40306 PAD.n4742 PAD.n4673 2.24164
R40307 PAD.n8397 PAD.n4717 2.24164
R40308 PAD.n8360 PAD.n4673 2.24164
R40309 PAD.n8397 PAD.n4716 2.24164
R40310 PAD.n4747 PAD.n4673 2.24164
R40311 PAD.n8397 PAD.n4715 2.24164
R40312 PAD.n8351 PAD.n4673 2.24164
R40313 PAD.n8397 PAD.n4714 2.24164
R40314 PAD.n4752 PAD.n4673 2.24164
R40315 PAD.n8397 PAD.n4713 2.24164
R40316 PAD.n8342 PAD.n4673 2.24164
R40317 PAD.n8397 PAD.n4712 2.24164
R40318 PAD.n4757 PAD.n4673 2.24164
R40319 PAD.n8397 PAD.n4711 2.24164
R40320 PAD.n8333 PAD.n4673 2.24164
R40321 PAD.n8397 PAD.n4710 2.24164
R40322 PAD.n4762 PAD.n4673 2.24164
R40323 PAD.n8397 PAD.n4709 2.24164
R40324 PAD.n8324 PAD.n4673 2.24164
R40325 PAD.n8397 PAD.n4708 2.24164
R40326 PAD.n4767 PAD.n4673 2.24164
R40327 PAD.n8397 PAD.n4707 2.24164
R40328 PAD.n8315 PAD.n4673 2.24164
R40329 PAD.n8397 PAD.n4706 2.24164
R40330 PAD.n4772 PAD.n4673 2.24164
R40331 PAD.n8397 PAD.n4705 2.24164
R40332 PAD.n8306 PAD.n4673 2.24164
R40333 PAD.n8397 PAD.n4704 2.24164
R40334 PAD.n4777 PAD.n4673 2.24164
R40335 PAD.n8397 PAD.n4703 2.24164
R40336 PAD.n8297 PAD.n4673 2.24164
R40337 PAD.n8397 PAD.n4702 2.24164
R40338 PAD.n4782 PAD.n4673 2.24164
R40339 PAD.n8397 PAD.n4701 2.24164
R40340 PAD.n8288 PAD.n4673 2.24164
R40341 PAD.n8397 PAD.n4700 2.24164
R40342 PAD.n4787 PAD.n4673 2.24164
R40343 PAD.n8397 PAD.n4699 2.24164
R40344 PAD.n8279 PAD.n4673 2.24164
R40345 PAD.n8397 PAD.n4698 2.24164
R40346 PAD.n4792 PAD.n4673 2.24164
R40347 PAD.n8397 PAD.n4697 2.24164
R40348 PAD.n8270 PAD.n4673 2.24164
R40349 PAD.n8397 PAD.n4696 2.24164
R40350 PAD.n4797 PAD.n4673 2.24164
R40351 PAD.n8397 PAD.n4695 2.24164
R40352 PAD.n8261 PAD.n4673 2.24164
R40353 PAD.n8397 PAD.n4694 2.24164
R40354 PAD.n4802 PAD.n4673 2.24164
R40355 PAD.n8397 PAD.n4693 2.24164
R40356 PAD.n8252 PAD.n4673 2.24164
R40357 PAD.n8397 PAD.n4692 2.24164
R40358 PAD.n4807 PAD.n4673 2.24164
R40359 PAD.n8397 PAD.n4691 2.24164
R40360 PAD.n8243 PAD.n4673 2.24164
R40361 PAD.n8397 PAD.n4690 2.24164
R40362 PAD.n4812 PAD.n4673 2.24164
R40363 PAD.n8397 PAD.n4689 2.24164
R40364 PAD.n8234 PAD.n4673 2.24164
R40365 PAD.n8397 PAD.n4688 2.24164
R40366 PAD.n4817 PAD.n4673 2.24164
R40367 PAD.n8397 PAD.n4687 2.24164
R40368 PAD.n8225 PAD.n4673 2.24164
R40369 PAD.n8397 PAD.n4686 2.24164
R40370 PAD.n4822 PAD.n4673 2.24164
R40371 PAD.n8397 PAD.n4685 2.24164
R40372 PAD.n8216 PAD.n4673 2.24164
R40373 PAD.n8397 PAD.n4684 2.24164
R40374 PAD.n4827 PAD.n4673 2.24164
R40375 PAD.n8397 PAD.n4683 2.24164
R40376 PAD.n4849 PAD.n4840 2.24164
R40377 PAD.n5175 PAD.n4843 2.24164
R40378 PAD.n5173 PAD.n4840 2.24164
R40379 PAD.n4850 PAD.n4843 2.24164
R40380 PAD.n5165 PAD.n4840 2.24164
R40381 PAD.n5163 PAD.n4843 2.24164
R40382 PAD.n5161 PAD.n4840 2.24164
R40383 PAD.n4855 PAD.n4843 2.24164
R40384 PAD.n5153 PAD.n4840 2.24164
R40385 PAD.n5151 PAD.n4843 2.24164
R40386 PAD.n5149 PAD.n4840 2.24164
R40387 PAD.n4859 PAD.n4843 2.24164
R40388 PAD.n5141 PAD.n4840 2.24164
R40389 PAD.n5139 PAD.n4843 2.24164
R40390 PAD.n5137 PAD.n4840 2.24164
R40391 PAD.n4863 PAD.n4843 2.24164
R40392 PAD.n5129 PAD.n4840 2.24164
R40393 PAD.n5127 PAD.n4843 2.24164
R40394 PAD.n5125 PAD.n4840 2.24164
R40395 PAD.n4867 PAD.n4843 2.24164
R40396 PAD.n5117 PAD.n4840 2.24164
R40397 PAD.n5115 PAD.n4843 2.24164
R40398 PAD.n5113 PAD.n4840 2.24164
R40399 PAD.n4871 PAD.n4843 2.24164
R40400 PAD.n5105 PAD.n4840 2.24164
R40401 PAD.n5103 PAD.n4843 2.24164
R40402 PAD.n5101 PAD.n4840 2.24164
R40403 PAD.n4875 PAD.n4843 2.24164
R40404 PAD.n5093 PAD.n4840 2.24164
R40405 PAD.n5091 PAD.n4843 2.24164
R40406 PAD.n5089 PAD.n4840 2.24164
R40407 PAD.n4879 PAD.n4843 2.24164
R40408 PAD.n5081 PAD.n4840 2.24164
R40409 PAD.n5079 PAD.n4843 2.24164
R40410 PAD.n5077 PAD.n4840 2.24164
R40411 PAD.n4883 PAD.n4843 2.24164
R40412 PAD.n5069 PAD.n4840 2.24164
R40413 PAD.n5067 PAD.n4843 2.24164
R40414 PAD.n5065 PAD.n4840 2.24164
R40415 PAD.n4887 PAD.n4843 2.24164
R40416 PAD.n5057 PAD.n4840 2.24164
R40417 PAD.n5055 PAD.n4843 2.24164
R40418 PAD.n5053 PAD.n4840 2.24164
R40419 PAD.n4891 PAD.n4843 2.24164
R40420 PAD.n5045 PAD.n4840 2.24164
R40421 PAD.n5043 PAD.n4843 2.24164
R40422 PAD.n5041 PAD.n4840 2.24164
R40423 PAD.n4895 PAD.n4843 2.24164
R40424 PAD.n5033 PAD.n4840 2.24164
R40425 PAD.n5031 PAD.n4843 2.24164
R40426 PAD.n5029 PAD.n4840 2.24164
R40427 PAD.n4899 PAD.n4843 2.24164
R40428 PAD.n5021 PAD.n4840 2.24164
R40429 PAD.n5019 PAD.n4843 2.24164
R40430 PAD.n5017 PAD.n4840 2.24164
R40431 PAD.n4903 PAD.n4843 2.24164
R40432 PAD.n5009 PAD.n4840 2.24164
R40433 PAD.n5007 PAD.n4843 2.24164
R40434 PAD.n5005 PAD.n4840 2.24164
R40435 PAD.n4907 PAD.n4843 2.24164
R40436 PAD.n4997 PAD.n4840 2.24164
R40437 PAD.n4995 PAD.n4843 2.24164
R40438 PAD.n4993 PAD.n4840 2.24164
R40439 PAD.n4911 PAD.n4843 2.24164
R40440 PAD.n4985 PAD.n4840 2.24164
R40441 PAD.n4983 PAD.n4843 2.24164
R40442 PAD.n4981 PAD.n4840 2.24164
R40443 PAD.n4915 PAD.n4843 2.24164
R40444 PAD.n4973 PAD.n4840 2.24164
R40445 PAD.n4971 PAD.n4843 2.24164
R40446 PAD.n4969 PAD.n4840 2.24164
R40447 PAD.n4919 PAD.n4843 2.24164
R40448 PAD.n4961 PAD.n4840 2.24164
R40449 PAD.n4959 PAD.n4843 2.24164
R40450 PAD.n4957 PAD.n4840 2.24164
R40451 PAD.n4923 PAD.n4843 2.24164
R40452 PAD.n4949 PAD.n4840 2.24164
R40453 PAD.n4947 PAD.n4843 2.24164
R40454 PAD.n4945 PAD.n4840 2.24164
R40455 PAD.n4927 PAD.n4843 2.24164
R40456 PAD.n4937 PAD.n4840 2.24164
R40457 PAD.n4935 PAD.n4843 2.24164
R40458 PAD.n4933 PAD.n4840 2.24164
R40459 PAD.n8163 PAD.n8162 2.24164
R40460 PAD.n7872 PAD.n5183 2.24164
R40461 PAD.n8163 PAD.n7870 2.24164
R40462 PAD.n8153 PAD.n5183 2.24164
R40463 PAD.n8163 PAD.n7869 2.24164
R40464 PAD.n7878 PAD.n5183 2.24164
R40465 PAD.n8163 PAD.n7868 2.24164
R40466 PAD.n8144 PAD.n5183 2.24164
R40467 PAD.n8163 PAD.n7867 2.24164
R40468 PAD.n7883 PAD.n5183 2.24164
R40469 PAD.n8163 PAD.n7866 2.24164
R40470 PAD.n8135 PAD.n5183 2.24164
R40471 PAD.n8163 PAD.n7865 2.24164
R40472 PAD.n7888 PAD.n5183 2.24164
R40473 PAD.n8163 PAD.n7864 2.24164
R40474 PAD.n8126 PAD.n5183 2.24164
R40475 PAD.n8163 PAD.n7863 2.24164
R40476 PAD.n7893 PAD.n5183 2.24164
R40477 PAD.n8163 PAD.n7862 2.24164
R40478 PAD.n8117 PAD.n5183 2.24164
R40479 PAD.n8163 PAD.n7861 2.24164
R40480 PAD.n7898 PAD.n5183 2.24164
R40481 PAD.n8163 PAD.n7860 2.24164
R40482 PAD.n8108 PAD.n5183 2.24164
R40483 PAD.n8163 PAD.n7859 2.24164
R40484 PAD.n7903 PAD.n5183 2.24164
R40485 PAD.n8163 PAD.n7858 2.24164
R40486 PAD.n8099 PAD.n5183 2.24164
R40487 PAD.n8163 PAD.n7857 2.24164
R40488 PAD.n7908 PAD.n5183 2.24164
R40489 PAD.n8163 PAD.n7856 2.24164
R40490 PAD.n8090 PAD.n5183 2.24164
R40491 PAD.n8163 PAD.n7855 2.24164
R40492 PAD.n7913 PAD.n5183 2.24164
R40493 PAD.n8163 PAD.n7854 2.24164
R40494 PAD.n8081 PAD.n5183 2.24164
R40495 PAD.n8163 PAD.n7853 2.24164
R40496 PAD.n7918 PAD.n5183 2.24164
R40497 PAD.n8163 PAD.n7852 2.24164
R40498 PAD.n8072 PAD.n5183 2.24164
R40499 PAD.n8163 PAD.n7851 2.24164
R40500 PAD.n7923 PAD.n5183 2.24164
R40501 PAD.n8163 PAD.n7850 2.24164
R40502 PAD.n8063 PAD.n5183 2.24164
R40503 PAD.n8163 PAD.n7849 2.24164
R40504 PAD.n7928 PAD.n5183 2.24164
R40505 PAD.n8163 PAD.n7848 2.24164
R40506 PAD.n8054 PAD.n5183 2.24164
R40507 PAD.n8163 PAD.n7847 2.24164
R40508 PAD.n7933 PAD.n5183 2.24164
R40509 PAD.n8163 PAD.n7846 2.24164
R40510 PAD.n8045 PAD.n5183 2.24164
R40511 PAD.n8163 PAD.n7845 2.24164
R40512 PAD.n7938 PAD.n5183 2.24164
R40513 PAD.n8163 PAD.n7844 2.24164
R40514 PAD.n8036 PAD.n5183 2.24164
R40515 PAD.n8163 PAD.n7843 2.24164
R40516 PAD.n7943 PAD.n5183 2.24164
R40517 PAD.n8163 PAD.n7842 2.24164
R40518 PAD.n8027 PAD.n5183 2.24164
R40519 PAD.n8163 PAD.n7841 2.24164
R40520 PAD.n7948 PAD.n5183 2.24164
R40521 PAD.n8163 PAD.n7840 2.24164
R40522 PAD.n8018 PAD.n5183 2.24164
R40523 PAD.n8163 PAD.n7839 2.24164
R40524 PAD.n7953 PAD.n5183 2.24164
R40525 PAD.n8163 PAD.n7838 2.24164
R40526 PAD.n8009 PAD.n5183 2.24164
R40527 PAD.n8163 PAD.n7837 2.24164
R40528 PAD.n7958 PAD.n5183 2.24164
R40529 PAD.n8163 PAD.n7836 2.24164
R40530 PAD.n8000 PAD.n5183 2.24164
R40531 PAD.n8163 PAD.n7835 2.24164
R40532 PAD.n7963 PAD.n5183 2.24164
R40533 PAD.n8163 PAD.n7834 2.24164
R40534 PAD.n7991 PAD.n5183 2.24164
R40535 PAD.n8163 PAD.n7833 2.24164
R40536 PAD.n7968 PAD.n5183 2.24164
R40537 PAD.n8163 PAD.n7832 2.24164
R40538 PAD.n7982 PAD.n5183 2.24164
R40539 PAD.n8163 PAD.n7831 2.24164
R40540 PAD.n7975 PAD.n5183 2.24164
R40541 PAD.n8163 PAD.n7830 2.24164
R40542 PAD.n5213 PAD.n5204 2.24164
R40543 PAD.n5539 PAD.n5197 2.24164
R40544 PAD.n5537 PAD.n5204 2.24164
R40545 PAD.n5214 PAD.n5197 2.24164
R40546 PAD.n5529 PAD.n5204 2.24164
R40547 PAD.n5527 PAD.n5197 2.24164
R40548 PAD.n5525 PAD.n5204 2.24164
R40549 PAD.n5219 PAD.n5197 2.24164
R40550 PAD.n5517 PAD.n5204 2.24164
R40551 PAD.n5515 PAD.n5197 2.24164
R40552 PAD.n5513 PAD.n5204 2.24164
R40553 PAD.n5223 PAD.n5197 2.24164
R40554 PAD.n5505 PAD.n5204 2.24164
R40555 PAD.n5503 PAD.n5197 2.24164
R40556 PAD.n5501 PAD.n5204 2.24164
R40557 PAD.n5227 PAD.n5197 2.24164
R40558 PAD.n5493 PAD.n5204 2.24164
R40559 PAD.n5491 PAD.n5197 2.24164
R40560 PAD.n5489 PAD.n5204 2.24164
R40561 PAD.n5231 PAD.n5197 2.24164
R40562 PAD.n5481 PAD.n5204 2.24164
R40563 PAD.n5479 PAD.n5197 2.24164
R40564 PAD.n5477 PAD.n5204 2.24164
R40565 PAD.n5235 PAD.n5197 2.24164
R40566 PAD.n5469 PAD.n5204 2.24164
R40567 PAD.n5467 PAD.n5197 2.24164
R40568 PAD.n5465 PAD.n5204 2.24164
R40569 PAD.n5239 PAD.n5197 2.24164
R40570 PAD.n5457 PAD.n5204 2.24164
R40571 PAD.n5455 PAD.n5197 2.24164
R40572 PAD.n5453 PAD.n5204 2.24164
R40573 PAD.n5243 PAD.n5197 2.24164
R40574 PAD.n5445 PAD.n5204 2.24164
R40575 PAD.n5443 PAD.n5197 2.24164
R40576 PAD.n5441 PAD.n5204 2.24164
R40577 PAD.n5247 PAD.n5197 2.24164
R40578 PAD.n5433 PAD.n5204 2.24164
R40579 PAD.n5431 PAD.n5197 2.24164
R40580 PAD.n5429 PAD.n5204 2.24164
R40581 PAD.n5251 PAD.n5197 2.24164
R40582 PAD.n5421 PAD.n5204 2.24164
R40583 PAD.n5419 PAD.n5197 2.24164
R40584 PAD.n5417 PAD.n5204 2.24164
R40585 PAD.n5255 PAD.n5197 2.24164
R40586 PAD.n5409 PAD.n5204 2.24164
R40587 PAD.n5407 PAD.n5197 2.24164
R40588 PAD.n5405 PAD.n5204 2.24164
R40589 PAD.n5259 PAD.n5197 2.24164
R40590 PAD.n5397 PAD.n5204 2.24164
R40591 PAD.n5395 PAD.n5197 2.24164
R40592 PAD.n5393 PAD.n5204 2.24164
R40593 PAD.n5263 PAD.n5197 2.24164
R40594 PAD.n5385 PAD.n5204 2.24164
R40595 PAD.n5383 PAD.n5197 2.24164
R40596 PAD.n5381 PAD.n5204 2.24164
R40597 PAD.n5267 PAD.n5197 2.24164
R40598 PAD.n5373 PAD.n5204 2.24164
R40599 PAD.n5371 PAD.n5197 2.24164
R40600 PAD.n5369 PAD.n5204 2.24164
R40601 PAD.n5271 PAD.n5197 2.24164
R40602 PAD.n5361 PAD.n5204 2.24164
R40603 PAD.n5359 PAD.n5197 2.24164
R40604 PAD.n5357 PAD.n5204 2.24164
R40605 PAD.n5275 PAD.n5197 2.24164
R40606 PAD.n5349 PAD.n5204 2.24164
R40607 PAD.n5347 PAD.n5197 2.24164
R40608 PAD.n5345 PAD.n5204 2.24164
R40609 PAD.n5279 PAD.n5197 2.24164
R40610 PAD.n5337 PAD.n5204 2.24164
R40611 PAD.n5335 PAD.n5197 2.24164
R40612 PAD.n5333 PAD.n5204 2.24164
R40613 PAD.n5283 PAD.n5197 2.24164
R40614 PAD.n5325 PAD.n5204 2.24164
R40615 PAD.n5323 PAD.n5197 2.24164
R40616 PAD.n5321 PAD.n5204 2.24164
R40617 PAD.n5287 PAD.n5197 2.24164
R40618 PAD.n5313 PAD.n5204 2.24164
R40619 PAD.n5311 PAD.n5197 2.24164
R40620 PAD.n5309 PAD.n5204 2.24164
R40621 PAD.n5291 PAD.n5197 2.24164
R40622 PAD.n5301 PAD.n5204 2.24164
R40623 PAD.n5299 PAD.n5197 2.24164
R40624 PAD.n5297 PAD.n5204 2.24164
R40625 PAD.n7520 PAD.n7519 2.24164
R40626 PAD.n7511 PAD.n7207 2.24164
R40627 PAD.n7520 PAD.n7199 2.24164
R40628 PAD.n7508 PAD.n7207 2.24164
R40629 PAD.n7520 PAD.n7198 2.24164
R40630 PAD.n7500 PAD.n7207 2.24164
R40631 PAD.n7520 PAD.n7197 2.24164
R40632 PAD.n7496 PAD.n7207 2.24164
R40633 PAD.n7520 PAD.n7196 2.24164
R40634 PAD.n7488 PAD.n7207 2.24164
R40635 PAD.n7520 PAD.n7195 2.24164
R40636 PAD.n7484 PAD.n7207 2.24164
R40637 PAD.n7520 PAD.n7194 2.24164
R40638 PAD.n7476 PAD.n7207 2.24164
R40639 PAD.n7520 PAD.n7193 2.24164
R40640 PAD.n7472 PAD.n7207 2.24164
R40641 PAD.n7520 PAD.n7192 2.24164
R40642 PAD.n7464 PAD.n7207 2.24164
R40643 PAD.n7520 PAD.n7191 2.24164
R40644 PAD.n7460 PAD.n7207 2.24164
R40645 PAD.n7520 PAD.n7190 2.24164
R40646 PAD.n7452 PAD.n7207 2.24164
R40647 PAD.n7520 PAD.n7189 2.24164
R40648 PAD.n7448 PAD.n7207 2.24164
R40649 PAD.n7520 PAD.n7188 2.24164
R40650 PAD.n7440 PAD.n7207 2.24164
R40651 PAD.n7520 PAD.n7187 2.24164
R40652 PAD.n7436 PAD.n7207 2.24164
R40653 PAD.n7520 PAD.n7186 2.24164
R40654 PAD.n7428 PAD.n7207 2.24164
R40655 PAD.n7520 PAD.n7185 2.24164
R40656 PAD.n7424 PAD.n7207 2.24164
R40657 PAD.n7520 PAD.n7184 2.24164
R40658 PAD.n7416 PAD.n7207 2.24164
R40659 PAD.n7520 PAD.n7183 2.24164
R40660 PAD.n7412 PAD.n7207 2.24164
R40661 PAD.n7520 PAD.n7182 2.24164
R40662 PAD.n7404 PAD.n7207 2.24164
R40663 PAD.n7520 PAD.n7181 2.24164
R40664 PAD.n7400 PAD.n7207 2.24164
R40665 PAD.n7520 PAD.n7180 2.24164
R40666 PAD.n7392 PAD.n7207 2.24164
R40667 PAD.n7520 PAD.n7179 2.24164
R40668 PAD.n7388 PAD.n7207 2.24164
R40669 PAD.n7520 PAD.n7178 2.24164
R40670 PAD.n7380 PAD.n7207 2.24164
R40671 PAD.n7520 PAD.n7177 2.24164
R40672 PAD.n7376 PAD.n7207 2.24164
R40673 PAD.n7520 PAD.n7176 2.24164
R40674 PAD.n7368 PAD.n7207 2.24164
R40675 PAD.n7520 PAD.n7175 2.24164
R40676 PAD.n7364 PAD.n7207 2.24164
R40677 PAD.n7520 PAD.n7174 2.24164
R40678 PAD.n7356 PAD.n7207 2.24164
R40679 PAD.n7520 PAD.n7173 2.24164
R40680 PAD.n7352 PAD.n7207 2.24164
R40681 PAD.n7520 PAD.n7172 2.24164
R40682 PAD.n7344 PAD.n7207 2.24164
R40683 PAD.n7520 PAD.n7171 2.24164
R40684 PAD.n7340 PAD.n7207 2.24164
R40685 PAD.n7520 PAD.n7170 2.24164
R40686 PAD.n7332 PAD.n7207 2.24164
R40687 PAD.n7520 PAD.n7169 2.24164
R40688 PAD.n7328 PAD.n7207 2.24164
R40689 PAD.n7520 PAD.n7168 2.24164
R40690 PAD.n7320 PAD.n7207 2.24164
R40691 PAD.n7520 PAD.n7167 2.24164
R40692 PAD.n7316 PAD.n7207 2.24164
R40693 PAD.n7520 PAD.n7166 2.24164
R40694 PAD.n7308 PAD.n7207 2.24164
R40695 PAD.n7520 PAD.n7165 2.24164
R40696 PAD.n7304 PAD.n7207 2.24164
R40697 PAD.n7520 PAD.n7164 2.24164
R40698 PAD.n7296 PAD.n7207 2.24164
R40699 PAD.n7520 PAD.n7163 2.24164
R40700 PAD.n7292 PAD.n7207 2.24164
R40701 PAD.n7520 PAD.n7162 2.24164
R40702 PAD.n7284 PAD.n7207 2.24164
R40703 PAD.n7520 PAD.n7161 2.24164
R40704 PAD.n7280 PAD.n7207 2.24164
R40705 PAD.n7520 PAD.n7160 2.24164
R40706 PAD.n7272 PAD.n7207 2.24164
R40707 PAD.n7520 PAD.n7159 2.24164
R40708 PAD.n7782 PAD.n7781 2.24164
R40709 PAD.n7773 PAD.n7105 2.24164
R40710 PAD.n7782 PAD.n7102 2.24164
R40711 PAD.n7770 PAD.n7105 2.24164
R40712 PAD.n7782 PAD.n7101 2.24164
R40713 PAD.n7762 PAD.n7105 2.24164
R40714 PAD.n7782 PAD.n7100 2.24164
R40715 PAD.n7758 PAD.n7105 2.24164
R40716 PAD.n7782 PAD.n7099 2.24164
R40717 PAD.n7750 PAD.n7105 2.24164
R40718 PAD.n7782 PAD.n7098 2.24164
R40719 PAD.n7746 PAD.n7105 2.24164
R40720 PAD.n7782 PAD.n7097 2.24164
R40721 PAD.n7738 PAD.n7105 2.24164
R40722 PAD.n7782 PAD.n7096 2.24164
R40723 PAD.n7734 PAD.n7105 2.24164
R40724 PAD.n7782 PAD.n7095 2.24164
R40725 PAD.n7726 PAD.n7105 2.24164
R40726 PAD.n7782 PAD.n7094 2.24164
R40727 PAD.n7722 PAD.n7105 2.24164
R40728 PAD.n7782 PAD.n7093 2.24164
R40729 PAD.n7714 PAD.n7105 2.24164
R40730 PAD.n7782 PAD.n7092 2.24164
R40731 PAD.n7710 PAD.n7105 2.24164
R40732 PAD.n7782 PAD.n7091 2.24164
R40733 PAD.n7702 PAD.n7105 2.24164
R40734 PAD.n7782 PAD.n7090 2.24164
R40735 PAD.n7698 PAD.n7105 2.24164
R40736 PAD.n7782 PAD.n7089 2.24164
R40737 PAD.n7690 PAD.n7105 2.24164
R40738 PAD.n7782 PAD.n7088 2.24164
R40739 PAD.n7686 PAD.n7105 2.24164
R40740 PAD.n7782 PAD.n7087 2.24164
R40741 PAD.n7678 PAD.n7105 2.24164
R40742 PAD.n7782 PAD.n7086 2.24164
R40743 PAD.n7674 PAD.n7105 2.24164
R40744 PAD.n7782 PAD.n7085 2.24164
R40745 PAD.n7666 PAD.n7105 2.24164
R40746 PAD.n7782 PAD.n7084 2.24164
R40747 PAD.n7662 PAD.n7105 2.24164
R40748 PAD.n7782 PAD.n7083 2.24164
R40749 PAD.n7654 PAD.n7105 2.24164
R40750 PAD.n7782 PAD.n7082 2.24164
R40751 PAD.n7650 PAD.n7105 2.24164
R40752 PAD.n7782 PAD.n7081 2.24164
R40753 PAD.n7642 PAD.n7105 2.24164
R40754 PAD.n7782 PAD.n7080 2.24164
R40755 PAD.n7638 PAD.n7105 2.24164
R40756 PAD.n7782 PAD.n7079 2.24164
R40757 PAD.n7630 PAD.n7105 2.24164
R40758 PAD.n7782 PAD.n7078 2.24164
R40759 PAD.n7626 PAD.n7105 2.24164
R40760 PAD.n7782 PAD.n7077 2.24164
R40761 PAD.n7618 PAD.n7105 2.24164
R40762 PAD.n7782 PAD.n7076 2.24164
R40763 PAD.n7614 PAD.n7105 2.24164
R40764 PAD.n7782 PAD.n7075 2.24164
R40765 PAD.n7606 PAD.n7105 2.24164
R40766 PAD.n7782 PAD.n7074 2.24164
R40767 PAD.n7602 PAD.n7105 2.24164
R40768 PAD.n7782 PAD.n7073 2.24164
R40769 PAD.n7594 PAD.n7105 2.24164
R40770 PAD.n7782 PAD.n7072 2.24164
R40771 PAD.n7590 PAD.n7105 2.24164
R40772 PAD.n7782 PAD.n7071 2.24164
R40773 PAD.n7582 PAD.n7105 2.24164
R40774 PAD.n7782 PAD.n7070 2.24164
R40775 PAD.n7578 PAD.n7105 2.24164
R40776 PAD.n7782 PAD.n7069 2.24164
R40777 PAD.n7570 PAD.n7105 2.24164
R40778 PAD.n7782 PAD.n7068 2.24164
R40779 PAD.n7566 PAD.n7105 2.24164
R40780 PAD.n7782 PAD.n7067 2.24164
R40781 PAD.n7558 PAD.n7105 2.24164
R40782 PAD.n7782 PAD.n7066 2.24164
R40783 PAD.n7554 PAD.n7105 2.24164
R40784 PAD.n7782 PAD.n7065 2.24164
R40785 PAD.n7546 PAD.n7105 2.24164
R40786 PAD.n7782 PAD.n7064 2.24164
R40787 PAD.n7542 PAD.n7105 2.24164
R40788 PAD.n7782 PAD.n7063 2.24164
R40789 PAD.n7534 PAD.n7105 2.24164
R40790 PAD.n7782 PAD.n7062 2.24164
R40791 PAD.n6721 PAD.n6712 2.24164
R40792 PAD.n7047 PAD.n6713 2.24164
R40793 PAD.n7045 PAD.n6712 2.24164
R40794 PAD.n6722 PAD.n6713 2.24164
R40795 PAD.n7037 PAD.n6712 2.24164
R40796 PAD.n7035 PAD.n6713 2.24164
R40797 PAD.n7033 PAD.n6712 2.24164
R40798 PAD.n6727 PAD.n6713 2.24164
R40799 PAD.n7025 PAD.n6712 2.24164
R40800 PAD.n7023 PAD.n6713 2.24164
R40801 PAD.n7021 PAD.n6712 2.24164
R40802 PAD.n6731 PAD.n6713 2.24164
R40803 PAD.n7013 PAD.n6712 2.24164
R40804 PAD.n7011 PAD.n6713 2.24164
R40805 PAD.n7009 PAD.n6712 2.24164
R40806 PAD.n6735 PAD.n6713 2.24164
R40807 PAD.n7001 PAD.n6712 2.24164
R40808 PAD.n6999 PAD.n6713 2.24164
R40809 PAD.n6997 PAD.n6712 2.24164
R40810 PAD.n6739 PAD.n6713 2.24164
R40811 PAD.n6989 PAD.n6712 2.24164
R40812 PAD.n6987 PAD.n6713 2.24164
R40813 PAD.n6985 PAD.n6712 2.24164
R40814 PAD.n6743 PAD.n6713 2.24164
R40815 PAD.n6977 PAD.n6712 2.24164
R40816 PAD.n6975 PAD.n6713 2.24164
R40817 PAD.n6973 PAD.n6712 2.24164
R40818 PAD.n6747 PAD.n6713 2.24164
R40819 PAD.n6965 PAD.n6712 2.24164
R40820 PAD.n6963 PAD.n6713 2.24164
R40821 PAD.n6961 PAD.n6712 2.24164
R40822 PAD.n6751 PAD.n6713 2.24164
R40823 PAD.n6953 PAD.n6712 2.24164
R40824 PAD.n6951 PAD.n6713 2.24164
R40825 PAD.n6949 PAD.n6712 2.24164
R40826 PAD.n6755 PAD.n6713 2.24164
R40827 PAD.n6941 PAD.n6712 2.24164
R40828 PAD.n6939 PAD.n6713 2.24164
R40829 PAD.n6937 PAD.n6712 2.24164
R40830 PAD.n6759 PAD.n6713 2.24164
R40831 PAD.n6929 PAD.n6712 2.24164
R40832 PAD.n6927 PAD.n6713 2.24164
R40833 PAD.n6925 PAD.n6712 2.24164
R40834 PAD.n6763 PAD.n6713 2.24164
R40835 PAD.n6917 PAD.n6712 2.24164
R40836 PAD.n6915 PAD.n6713 2.24164
R40837 PAD.n6913 PAD.n6712 2.24164
R40838 PAD.n6767 PAD.n6713 2.24164
R40839 PAD.n6905 PAD.n6712 2.24164
R40840 PAD.n6903 PAD.n6713 2.24164
R40841 PAD.n6901 PAD.n6712 2.24164
R40842 PAD.n6771 PAD.n6713 2.24164
R40843 PAD.n6893 PAD.n6712 2.24164
R40844 PAD.n6891 PAD.n6713 2.24164
R40845 PAD.n6889 PAD.n6712 2.24164
R40846 PAD.n6775 PAD.n6713 2.24164
R40847 PAD.n6881 PAD.n6712 2.24164
R40848 PAD.n6879 PAD.n6713 2.24164
R40849 PAD.n6877 PAD.n6712 2.24164
R40850 PAD.n6779 PAD.n6713 2.24164
R40851 PAD.n6869 PAD.n6712 2.24164
R40852 PAD.n6867 PAD.n6713 2.24164
R40853 PAD.n6865 PAD.n6712 2.24164
R40854 PAD.n6783 PAD.n6713 2.24164
R40855 PAD.n6857 PAD.n6712 2.24164
R40856 PAD.n6855 PAD.n6713 2.24164
R40857 PAD.n6853 PAD.n6712 2.24164
R40858 PAD.n6787 PAD.n6713 2.24164
R40859 PAD.n6845 PAD.n6712 2.24164
R40860 PAD.n6843 PAD.n6713 2.24164
R40861 PAD.n6841 PAD.n6712 2.24164
R40862 PAD.n6791 PAD.n6713 2.24164
R40863 PAD.n6833 PAD.n6712 2.24164
R40864 PAD.n6831 PAD.n6713 2.24164
R40865 PAD.n6829 PAD.n6712 2.24164
R40866 PAD.n6795 PAD.n6713 2.24164
R40867 PAD.n6821 PAD.n6712 2.24164
R40868 PAD.n6819 PAD.n6713 2.24164
R40869 PAD.n6817 PAD.n6712 2.24164
R40870 PAD.n6799 PAD.n6713 2.24164
R40871 PAD.n6809 PAD.n6712 2.24164
R40872 PAD.n6807 PAD.n6713 2.24164
R40873 PAD.n6805 PAD.n6712 2.24164
R40874 PAD.n5894 PAD.n5893 2.24164
R40875 PAD.n5603 PAD.n5551 2.24164
R40876 PAD.n5894 PAD.n5601 2.24164
R40877 PAD.n5884 PAD.n5551 2.24164
R40878 PAD.n5894 PAD.n5600 2.24164
R40879 PAD.n5609 PAD.n5551 2.24164
R40880 PAD.n5894 PAD.n5599 2.24164
R40881 PAD.n5875 PAD.n5551 2.24164
R40882 PAD.n5894 PAD.n5598 2.24164
R40883 PAD.n5614 PAD.n5551 2.24164
R40884 PAD.n5894 PAD.n5597 2.24164
R40885 PAD.n5866 PAD.n5551 2.24164
R40886 PAD.n5894 PAD.n5596 2.24164
R40887 PAD.n5619 PAD.n5551 2.24164
R40888 PAD.n5894 PAD.n5595 2.24164
R40889 PAD.n5857 PAD.n5551 2.24164
R40890 PAD.n5894 PAD.n5594 2.24164
R40891 PAD.n5624 PAD.n5551 2.24164
R40892 PAD.n5894 PAD.n5593 2.24164
R40893 PAD.n5848 PAD.n5551 2.24164
R40894 PAD.n5894 PAD.n5592 2.24164
R40895 PAD.n5629 PAD.n5551 2.24164
R40896 PAD.n5894 PAD.n5591 2.24164
R40897 PAD.n5839 PAD.n5551 2.24164
R40898 PAD.n5894 PAD.n5590 2.24164
R40899 PAD.n5634 PAD.n5551 2.24164
R40900 PAD.n5894 PAD.n5589 2.24164
R40901 PAD.n5830 PAD.n5551 2.24164
R40902 PAD.n5894 PAD.n5588 2.24164
R40903 PAD.n5639 PAD.n5551 2.24164
R40904 PAD.n5894 PAD.n5587 2.24164
R40905 PAD.n5821 PAD.n5551 2.24164
R40906 PAD.n5894 PAD.n5586 2.24164
R40907 PAD.n5644 PAD.n5551 2.24164
R40908 PAD.n5894 PAD.n5585 2.24164
R40909 PAD.n5812 PAD.n5551 2.24164
R40910 PAD.n5894 PAD.n5584 2.24164
R40911 PAD.n5649 PAD.n5551 2.24164
R40912 PAD.n5894 PAD.n5583 2.24164
R40913 PAD.n5803 PAD.n5551 2.24164
R40914 PAD.n5894 PAD.n5582 2.24164
R40915 PAD.n5654 PAD.n5551 2.24164
R40916 PAD.n5894 PAD.n5581 2.24164
R40917 PAD.n5794 PAD.n5551 2.24164
R40918 PAD.n5894 PAD.n5580 2.24164
R40919 PAD.n5659 PAD.n5551 2.24164
R40920 PAD.n5894 PAD.n5579 2.24164
R40921 PAD.n5785 PAD.n5551 2.24164
R40922 PAD.n5894 PAD.n5578 2.24164
R40923 PAD.n5664 PAD.n5551 2.24164
R40924 PAD.n5894 PAD.n5577 2.24164
R40925 PAD.n5776 PAD.n5551 2.24164
R40926 PAD.n5894 PAD.n5576 2.24164
R40927 PAD.n5669 PAD.n5551 2.24164
R40928 PAD.n5894 PAD.n5575 2.24164
R40929 PAD.n5767 PAD.n5551 2.24164
R40930 PAD.n5894 PAD.n5574 2.24164
R40931 PAD.n5674 PAD.n5551 2.24164
R40932 PAD.n5894 PAD.n5573 2.24164
R40933 PAD.n5758 PAD.n5551 2.24164
R40934 PAD.n5894 PAD.n5572 2.24164
R40935 PAD.n5679 PAD.n5551 2.24164
R40936 PAD.n5894 PAD.n5571 2.24164
R40937 PAD.n5749 PAD.n5551 2.24164
R40938 PAD.n5894 PAD.n5570 2.24164
R40939 PAD.n5684 PAD.n5551 2.24164
R40940 PAD.n5894 PAD.n5569 2.24164
R40941 PAD.n5740 PAD.n5551 2.24164
R40942 PAD.n5894 PAD.n5568 2.24164
R40943 PAD.n5689 PAD.n5551 2.24164
R40944 PAD.n5894 PAD.n5567 2.24164
R40945 PAD.n5731 PAD.n5551 2.24164
R40946 PAD.n5894 PAD.n5566 2.24164
R40947 PAD.n5694 PAD.n5551 2.24164
R40948 PAD.n5894 PAD.n5565 2.24164
R40949 PAD.n5722 PAD.n5551 2.24164
R40950 PAD.n5894 PAD.n5564 2.24164
R40951 PAD.n5699 PAD.n5551 2.24164
R40952 PAD.n5894 PAD.n5563 2.24164
R40953 PAD.n5713 PAD.n5551 2.24164
R40954 PAD.n5894 PAD.n5562 2.24164
R40955 PAD.n5706 PAD.n5551 2.24164
R40956 PAD.n5894 PAD.n5561 2.24164
R40957 PAD.n6678 PAD.n5902 2.24164
R40958 PAD.n6689 PAD.n5906 2.24164
R40959 PAD.n6678 PAD.n6397 2.24164
R40960 PAD.n6689 PAD.n5907 2.24164
R40961 PAD.n6678 PAD.n6398 2.24164
R40962 PAD.n6689 PAD.n5908 2.24164
R40963 PAD.n6678 PAD.n6399 2.24164
R40964 PAD.n6689 PAD.n5909 2.24164
R40965 PAD.n6678 PAD.n6400 2.24164
R40966 PAD.n6689 PAD.n5910 2.24164
R40967 PAD.n6678 PAD.n6401 2.24164
R40968 PAD.n6689 PAD.n5911 2.24164
R40969 PAD.n6678 PAD.n6402 2.24164
R40970 PAD.n6689 PAD.n5912 2.24164
R40971 PAD.n6678 PAD.n6403 2.24164
R40972 PAD.n6689 PAD.n5913 2.24164
R40973 PAD.n6678 PAD.n6404 2.24164
R40974 PAD.n6689 PAD.n5914 2.24164
R40975 PAD.n6678 PAD.n6405 2.24164
R40976 PAD.n6689 PAD.n5915 2.24164
R40977 PAD.n6678 PAD.n6406 2.24164
R40978 PAD.n6689 PAD.n5916 2.24164
R40979 PAD.n6678 PAD.n6407 2.24164
R40980 PAD.n6689 PAD.n5917 2.24164
R40981 PAD.n6678 PAD.n6408 2.24164
R40982 PAD.n6689 PAD.n5918 2.24164
R40983 PAD.n6678 PAD.n6409 2.24164
R40984 PAD.n6689 PAD.n5919 2.24164
R40985 PAD.n6678 PAD.n6410 2.24164
R40986 PAD.n6689 PAD.n5920 2.24164
R40987 PAD.n6678 PAD.n6411 2.24164
R40988 PAD.n6689 PAD.n5921 2.24164
R40989 PAD.n6678 PAD.n6412 2.24164
R40990 PAD.n6689 PAD.n5922 2.24164
R40991 PAD.n6678 PAD.n6413 2.24164
R40992 PAD.n6689 PAD.n5923 2.24164
R40993 PAD.n6678 PAD.n6414 2.24164
R40994 PAD.n6689 PAD.n5924 2.24164
R40995 PAD.n6678 PAD.n6415 2.24164
R40996 PAD.n6689 PAD.n5925 2.24164
R40997 PAD.n6678 PAD.n6416 2.24164
R40998 PAD.n6689 PAD.n5926 2.24164
R40999 PAD.n6678 PAD.n6417 2.24164
R41000 PAD.n6689 PAD.n5927 2.24164
R41001 PAD.n6678 PAD.n6418 2.24164
R41002 PAD.n6689 PAD.n5928 2.24164
R41003 PAD.n6678 PAD.n6419 2.24164
R41004 PAD.n6689 PAD.n5929 2.24164
R41005 PAD.n6678 PAD.n6420 2.24164
R41006 PAD.n6689 PAD.n5930 2.24164
R41007 PAD.n6678 PAD.n6421 2.24164
R41008 PAD.n6689 PAD.n5931 2.24164
R41009 PAD.n6678 PAD.n6422 2.24164
R41010 PAD.n6689 PAD.n5932 2.24164
R41011 PAD.n6678 PAD.n6423 2.24164
R41012 PAD.n6689 PAD.n5933 2.24164
R41013 PAD.n6678 PAD.n6424 2.24164
R41014 PAD.n6689 PAD.n5934 2.24164
R41015 PAD.n6678 PAD.n6425 2.24164
R41016 PAD.n6689 PAD.n5935 2.24164
R41017 PAD.n6678 PAD.n6426 2.24164
R41018 PAD.n6689 PAD.n5936 2.24164
R41019 PAD.n6678 PAD.n6427 2.24164
R41020 PAD.n6689 PAD.n5937 2.24164
R41021 PAD.n6678 PAD.n6428 2.24164
R41022 PAD.n6689 PAD.n5938 2.24164
R41023 PAD.n6678 PAD.n6429 2.24164
R41024 PAD.n6689 PAD.n5939 2.24164
R41025 PAD.n6678 PAD.n6430 2.24164
R41026 PAD.n6689 PAD.n5940 2.24164
R41027 PAD.n6678 PAD.n6431 2.24164
R41028 PAD.n6689 PAD.n5941 2.24164
R41029 PAD.n6678 PAD.n6432 2.24164
R41030 PAD.n6689 PAD.n5942 2.24164
R41031 PAD.n6678 PAD.n6433 2.24164
R41032 PAD.n6689 PAD.n5943 2.24164
R41033 PAD.n6678 PAD.n6434 2.24164
R41034 PAD.n6689 PAD.n5944 2.24164
R41035 PAD.n6678 PAD.n6435 2.24164
R41036 PAD.n6689 PAD.n5945 2.24164
R41037 PAD.n6678 PAD.n6677 2.24164
R41038 PAD.n6689 PAD.n5946 2.24164
R41039 PAD.n6678 PAD.n5947 2.24164
R41040 PAD.n11518 PAD.n10745 1.1255
R41041 PAD.n11520 PAD.n11519 1.1255
R41042 PAD.n11089 PAD.n10744 1.1255
R41043 PAD.n10751 PAD.n10746 1.1255
R41044 PAD.n17 PAD.n15 1.1255
R41045 PAD.n11537 PAD.n11536 1.1255
R41046 PAD.n10725 PAD.n10724 1.1255
R41047 PAD.n10723 PAD.n369 1.1255
R41048 PAD.n10722 PAD.n10721 1.1255
R41049 PAD.n371 PAD.n370 1.1255
R41050 PAD.n10699 PAD.n10698 1.1255
R41051 PAD.n10412 PAD.n428 1.1255
R41052 PAD.n10411 PAD.n10410 1.1255
R41053 PAD.n10395 PAD.n10394 1.1255
R41054 PAD.n10393 PAD.n778 1.1255
R41055 PAD.n10392 PAD.n10391 1.1255
R41056 PAD.n10369 PAD.n1123 1.1255
R41057 PAD.n10371 PAD.n10370 1.1255
R41058 PAD.n10368 PAD.n1122 1.1255
R41059 PAD.n10365 PAD.n10364 1.1255
R41060 PAD.n1126 PAD.n1125 1.1255
R41061 PAD.n10014 PAD.n10013 1.1255
R41062 PAD.n10011 PAD.n10010 1.1255
R41063 PAD.n1147 PAD.n1146 1.1255
R41064 PAD.n1583 PAD.n1582 1.1255
R41065 PAD.n9747 PAD.n1584 1.1255
R41066 PAD.n9727 PAD.n1581 1.1255
R41067 PAD.n9728 PAD.n1597 1.1255
R41068 PAD.n9730 PAD.n9729 1.1255
R41069 PAD.n9725 PAD.n9724 1.1255
R41070 PAD.n1934 PAD.n1933 1.1255
R41071 PAD.n9461 PAD.n2034 1.1255
R41072 PAD.n9192 PAD.n2033 1.1255
R41073 PAD.n9193 PAD.n2036 1.1255
R41074 PAD.n9195 PAD.n9194 1.1255
R41075 PAD.n9191 PAD.n2137 1.1255
R41076 PAD.n9169 PAD.n2136 1.1255
R41077 PAD.n9170 PAD.n2149 1.1255
R41078 PAD.n9173 PAD.n9172 1.1255
R41079 PAD.n9166 PAD.n9165 1.1255
R41080 PAD.n2485 PAD.n2484 1.1255
R41081 PAD.n9149 PAD.n9148 1.1255
R41082 PAD.n9146 PAD.n9145 1.1255
R41083 PAD.n2832 PAD.n2831 1.1255
R41084 PAD.n9123 PAD.n9122 1.1255
R41085 PAD.n9126 PAD.n9125 1.1255
R41086 PAD.n8836 PAD.n2886 1.1255
R41087 PAD.n8835 PAD.n8834 1.1255
R41088 PAD.n8525 PAD.n8524 1.1255
R41089 PAD.n8523 PAD.n2948 1.1255
R41090 PAD.n8522 PAD.n8521 1.1255
R41091 PAD.n8498 PAD.n3292 1.1255
R41092 PAD.n8500 PAD.n8499 1.1255
R41093 PAD.n8497 PAD.n3291 1.1255
R41094 PAD.n8496 PAD.n8495 1.1255
R41095 PAD.n8476 PAD.n8475 1.1255
R41096 PAD.n8474 PAD.n3635 1.1255
R41097 PAD.n8472 PAD.n8471 1.1255
R41098 PAD.n8451 PAD.n8450 1.1255
R41099 PAD.n8449 PAD.n3979 1.1255
R41100 PAD.n8448 PAD.n8447 1.1255
R41101 PAD.n8426 PAD.n4324 1.1255
R41102 PAD.n8428 PAD.n8427 1.1255
R41103 PAD.n8425 PAD.n4323 1.1255
R41104 PAD.n8423 PAD.n8422 1.1255
R41105 PAD.n4327 PAD.n4326 1.1255
R41106 PAD.n8405 PAD.n8404 1.1255
R41107 PAD.n8403 PAD.n4675 1.1255
R41108 PAD.n8401 PAD.n8400 1.1255
R41109 PAD.n4678 PAD.n4677 1.1255
R41110 PAD.n8192 PAD.n8191 1.1255
R41111 PAD.n8189 PAD.n8188 1.1255
R41112 PAD.n5181 PAD.n5180 1.1255
R41113 PAD.n8172 PAD.n8171 1.1255
R41114 PAD.n8169 PAD.n8168 1.1255
R41115 PAD.n5195 PAD.n5194 1.1255
R41116 PAD.n7814 PAD.n7813 1.1255
R41117 PAD.n7817 PAD.n7816 1.1255
R41118 PAD.n5209 PAD.n5207 1.1255
R41119 PAD.n7226 PAD.n7225 1.1255
R41120 PAD.n7227 PAD.n7208 1.1255
R41121 PAD.n7220 PAD.n7219 1.1255
R41122 PAD.n7211 PAD.n7210 1.1255
R41123 PAD.n7213 PAD.n7212 1.1255
R41124 PAD.n7786 PAD.n7785 1.1255
R41125 PAD.n7787 PAD.n6717 1.1255
R41126 PAD.n7789 PAD.n7788 1.1255
R41127 PAD.n7054 PAD.n7053 1.1255
R41128 PAD.n5548 PAD.n5546 1.1255
R41129 PAD.n7805 PAD.n7804 1.1255
R41130 PAD.n6697 PAD.n5544 1.1255
R41131 PAD.n6696 PAD.n6695 1.1255
R41132 PAD.n6694 PAD.n5896 1.1255
R41133 PAD.n6394 PAD.n5897 1.1255
R41134 PAD.n6393 PAD.n6392 1.1255
R41135 PAD.n6391 PAD.n5955 1.1255
R41136 PAD.n5970 PAD.n5955 1.1255
R41137 PAD.n6393 PAD.n5954 1.1255
R41138 PAD.n6395 PAD.n6394 1.1255
R41139 PAD.n6681 PAD.n5896 1.1255
R41140 PAD.n6696 PAD.n5895 1.1255
R41141 PAD.n6698 PAD.n6697 1.1255
R41142 PAD.n7804 PAD.n7803 1.1255
R41143 PAD.n5550 PAD.n5548 1.1255
R41144 PAD.n7053 PAD.n7052 1.1255
R41145 PAD.n7790 PAD.n7789 1.1255
R41146 PAD.n6717 PAD.n6715 1.1255
R41147 PAD.n7785 PAD.n7784 1.1255
R41148 PAD.n7214 PAD.n7213 1.1255
R41149 PAD.n7217 PAD.n7211 1.1255
R41150 PAD.n7219 PAD.n7218 1.1255
R41151 PAD.n7208 PAD.n7202 1.1255
R41152 PAD.n7225 PAD.n7224 1.1255
R41153 PAD.n5207 PAD.n5205 1.1255
R41154 PAD.n7818 PAD.n7817 1.1255
R41155 PAD.n7813 PAD.n5196 1.1255
R41156 PAD.n8166 PAD.n5195 1.1255
R41157 PAD.n8168 PAD.n8167 1.1255
R41158 PAD.n8173 PAD.n8172 1.1255
R41159 PAD.n5182 PAD.n5181 1.1255
R41160 PAD.n8188 PAD.n8187 1.1255
R41161 PAD.n8193 PAD.n8192 1.1255
R41162 PAD.n4680 PAD.n4678 1.1255
R41163 PAD.n8400 PAD.n8399 1.1255
R41164 PAD.n4675 PAD.n4674 1.1255
R41165 PAD.n8406 PAD.n8405 1.1255
R41166 PAD.n4329 PAD.n4327 1.1255
R41167 PAD.n8422 PAD.n8421 1.1255
R41168 PAD.n4323 PAD.n4320 1.1255
R41169 PAD.n8429 PAD.n8428 1.1255
R41170 PAD.n4324 PAD.n4322 1.1255
R41171 PAD.n8447 PAD.n8446 1.1255
R41172 PAD.n3979 PAD.n3978 1.1255
R41173 PAD.n8452 PAD.n8451 1.1255
R41174 PAD.n8471 PAD.n8470 1.1255
R41175 PAD.n3635 PAD.n3634 1.1255
R41176 PAD.n8477 PAD.n8476 1.1255
R41177 PAD.n8495 PAD.n8494 1.1255
R41178 PAD.n3291 PAD.n3288 1.1255
R41179 PAD.n8501 PAD.n8500 1.1255
R41180 PAD.n3292 PAD.n3290 1.1255
R41181 PAD.n8521 PAD.n8520 1.1255
R41182 PAD.n2948 PAD.n2947 1.1255
R41183 PAD.n8526 PAD.n8525 1.1255
R41184 PAD.n8834 PAD.n8833 1.1255
R41185 PAD.n2886 PAD.n2884 1.1255
R41186 PAD.n9127 PAD.n9126 1.1255
R41187 PAD.n9122 PAD.n9121 1.1255
R41188 PAD.n2833 PAD.n2832 1.1255
R41189 PAD.n9145 PAD.n9144 1.1255
R41190 PAD.n9150 PAD.n9149 1.1255
R41191 PAD.n2486 PAD.n2485 1.1255
R41192 PAD.n9165 PAD.n9164 1.1255
R41193 PAD.n9174 PAD.n9173 1.1255
R41194 PAD.n2149 PAD.n2138 1.1255
R41195 PAD.n9188 PAD.n2136 1.1255
R41196 PAD.n9191 PAD.n9190 1.1255
R41197 PAD.n9195 PAD.n2035 1.1255
R41198 PAD.n9457 PAD.n2036 1.1255
R41199 PAD.n9458 PAD.n2033 1.1255
R41200 PAD.n9461 PAD.n9460 1.1255
R41201 PAD.n1935 PAD.n1934 1.1255
R41202 PAD.n9724 PAD.n9723 1.1255
R41203 PAD.n9731 PAD.n9730 1.1255
R41204 PAD.n1597 PAD.n1585 1.1255
R41205 PAD.n9743 PAD.n1581 1.1255
R41206 PAD.n9747 PAD.n9746 1.1255
R41207 PAD.n9745 PAD.n1582 1.1255
R41208 PAD.n1148 PAD.n1147 1.1255
R41209 PAD.n10010 PAD.n10009 1.1255
R41210 PAD.n10015 PAD.n10014 1.1255
R41211 PAD.n1128 PAD.n1126 1.1255
R41212 PAD.n10364 PAD.n10363 1.1255
R41213 PAD.n1122 PAD.n1119 1.1255
R41214 PAD.n10372 PAD.n10371 1.1255
R41215 PAD.n1123 PAD.n1121 1.1255
R41216 PAD.n10391 PAD.n10390 1.1255
R41217 PAD.n778 PAD.n777 1.1255
R41218 PAD.n10396 PAD.n10395 1.1255
R41219 PAD.n10410 PAD.n10409 1.1255
R41220 PAD.n428 PAD.n426 1.1255
R41221 PAD.n10700 PAD.n10699 1.1255
R41222 PAD.n372 PAD.n371 1.1255
R41223 PAD.n10721 PAD.n10720 1.1255
R41224 PAD.n369 PAD.n368 1.1255
R41225 PAD.n10726 PAD.n10725 1.1255
R41226 PAD.n11536 PAD.n11535 1.1255
R41227 PAD.n19 PAD.n17 1.1255
R41228 PAD.n10752 PAD.n10751 1.1255
R41229 PAD.n10744 PAD.n10742 1.1255
R41230 PAD.n11521 PAD.n11520 1.1255
R41231 PAD.n10745 PAD.n10743 1.1255
R41232 PAD.n5971 PAD.n5970 1.1255
R41233 PAD.n5954 PAD.n5903 1.1255
R41234 PAD.n6396 PAD.n6395 1.1255
R41235 PAD.n6682 PAD.n6681 1.1255
R41236 PAD.n6679 PAD.n5895 1.1255
R41237 PAD.n6699 PAD.n6698 1.1255
R41238 PAD.n7803 PAD.n7802 1.1255
R41239 PAD.n5552 PAD.n5550 1.1255
R41240 PAD.n7052 PAD.n6712 1.1255
R41241 PAD.n7791 PAD.n7790 1.1255
R41242 PAD.n7060 PAD.n6715 1.1255
R41243 PAD.n7784 PAD.n7783 1.1255
R41244 PAD.n7214 PAD.n7103 1.1255
R41245 PAD.n7217 PAD.n7216 1.1255
R41246 PAD.n7218 PAD.n7158 1.1255
R41247 PAD.n7202 PAD.n7200 1.1255
R41248 PAD.n7224 PAD.n7223 1.1255
R41249 PAD.n7221 PAD.n5205 1.1255
R41250 PAD.n7819 PAD.n7818 1.1255
R41251 PAD.n7829 PAD.n5196 1.1255
R41252 PAD.n8166 PAD.n8165 1.1255
R41253 PAD.n8167 PAD.n5190 1.1255
R41254 PAD.n8174 PAD.n8173 1.1255
R41255 PAD.n8184 PAD.n5182 1.1255
R41256 PAD.n8187 PAD.n8186 1.1255
R41257 PAD.n8194 PAD.n8193 1.1255
R41258 PAD.n4841 PAD.n4680 1.1255
R41259 PAD.n8399 PAD.n8398 1.1255
R41260 PAD.n4724 PAD.n4674 1.1255
R41261 PAD.n8407 PAD.n8406 1.1255
R41262 PAD.n8409 PAD.n4329 1.1255
R41263 PAD.n8421 PAD.n8420 1.1255
R41264 PAD.n4332 PAD.n4320 1.1255
R41265 PAD.n8430 PAD.n8429 1.1255
R41266 PAD.n4322 PAD.n4321 1.1255
R41267 PAD.n8446 PAD.n8445 1.1255
R41268 PAD.n3978 PAD.n3977 1.1255
R41269 PAD.n8453 PAD.n8452 1.1255
R41270 PAD.n8470 PAD.n8469 1.1255
R41271 PAD.n3634 PAD.n3633 1.1255
R41272 PAD.n8478 PAD.n8477 1.1255
R41273 PAD.n8494 PAD.n8493 1.1255
R41274 PAD.n3288 PAD.n3287 1.1255
R41275 PAD.n8502 PAD.n8501 1.1255
R41276 PAD.n3290 PAD.n3289 1.1255
R41277 PAD.n8520 PAD.n8519 1.1255
R41278 PAD.n2947 PAD.n2904 1.1255
R41279 PAD.n8527 PAD.n8526 1.1255
R41280 PAD.n8833 PAD.n8832 1.1255
R41281 PAD.n2892 PAD.n2884 1.1255
R41282 PAD.n9128 PAD.n9127 1.1255
R41283 PAD.n9121 PAD.n2834 1.1255
R41284 PAD.n9141 PAD.n2833 1.1255
R41285 PAD.n9144 PAD.n9143 1.1255
R41286 PAD.n9151 PAD.n9150 1.1255
R41287 PAD.n9161 PAD.n2486 1.1255
R41288 PAD.n9164 PAD.n9163 1.1255
R41289 PAD.n9175 PAD.n9174 1.1255
R41290 PAD.n9185 PAD.n2138 1.1255
R41291 PAD.n9188 PAD.n9187 1.1255
R41292 PAD.n9190 PAD.n2046 1.1255
R41293 PAD.n2089 PAD.n2035 1.1255
R41294 PAD.n9457 PAD.n9456 1.1255
R41295 PAD.n9458 PAD.n1942 1.1255
R41296 PAD.n9460 PAD.n1986 1.1255
R41297 PAD.n1936 PAD.n1935 1.1255
R41298 PAD.n9723 PAD.n9722 1.1255
R41299 PAD.n9732 PAD.n9731 1.1255
R41300 PAD.n1593 PAD.n1585 1.1255
R41301 PAD.n9743 PAD.n9742 1.1255
R41302 PAD.n9746 PAD.n1489 1.1255
R41303 PAD.n9745 PAD.n1534 1.1255
R41304 PAD.n1532 PAD.n1148 1.1255
R41305 PAD.n10009 PAD.n10008 1.1255
R41306 PAD.n10016 PAD.n10015 1.1255
R41307 PAD.n1141 PAD.n1128 1.1255
R41308 PAD.n10363 PAD.n10362 1.1255
R41309 PAD.n1131 PAD.n1119 1.1255
R41310 PAD.n10373 PAD.n10372 1.1255
R41311 PAD.n1121 PAD.n1120 1.1255
R41312 PAD.n10390 PAD.n10389 1.1255
R41313 PAD.n777 PAD.n776 1.1255
R41314 PAD.n10397 PAD.n10396 1.1255
R41315 PAD.n10409 PAD.n10408 1.1255
R41316 PAD.n434 PAD.n426 1.1255
R41317 PAD.n10701 PAD.n10700 1.1255
R41318 PAD.n418 PAD.n372 1.1255
R41319 PAD.n10720 PAD.n10719 1.1255
R41320 PAD.n10717 PAD.n368 1.1255
R41321 PAD.n10727 PAD.n10726 1.1255
R41322 PAD.n11535 PAD.n11534 1.1255
R41323 PAD.n11533 PAD.n19 1.1255
R41324 PAD.n10753 PAD.n10752 1.1255
R41325 PAD.n10742 PAD.n10740 1.1255
R41326 PAD.n11522 PAD.n11521 1.1255
R41327 PAD.n11500 PAD.n10743 1.1255
R41328 PAD.n4 PAD.t5 0.9641
R41329 PAD.n7 PAD.t3 0.9641
R41330 PAD.n2 PAD.t21 0.9641
R41331 PAD.n11506 PAD.n11505 0.902975
R41332 PAD.n6376 PAD.n6375 0.902975
R41333 PAD.n11498 PAD.n11156 0.9005
R41334 PAD.n11497 PAD.n11154 0.9005
R41335 PAD.n11496 PAD.n11158 0.9005
R41336 PAD.n11305 PAD.n11153 0.9005
R41337 PAD.n11492 PAD.n11160 0.9005
R41338 PAD.n11491 PAD.n11152 0.9005
R41339 PAD.n11490 PAD.n11162 0.9005
R41340 PAD.n11307 PAD.n11151 0.9005
R41341 PAD.n11486 PAD.n11164 0.9005
R41342 PAD.n11485 PAD.n11150 0.9005
R41343 PAD.n11484 PAD.n11166 0.9005
R41344 PAD.n11309 PAD.n11149 0.9005
R41345 PAD.n11480 PAD.n11168 0.9005
R41346 PAD.n11479 PAD.n11148 0.9005
R41347 PAD.n11478 PAD.n11170 0.9005
R41348 PAD.n11311 PAD.n11147 0.9005
R41349 PAD.n11474 PAD.n11172 0.9005
R41350 PAD.n11473 PAD.n11146 0.9005
R41351 PAD.n11472 PAD.n11174 0.9005
R41352 PAD.n11313 PAD.n11145 0.9005
R41353 PAD.n11468 PAD.n11176 0.9005
R41354 PAD.n11467 PAD.n11144 0.9005
R41355 PAD.n11466 PAD.n11178 0.9005
R41356 PAD.n11315 PAD.n11143 0.9005
R41357 PAD.n11462 PAD.n11180 0.9005
R41358 PAD.n11461 PAD.n11142 0.9005
R41359 PAD.n11460 PAD.n11182 0.9005
R41360 PAD.n11317 PAD.n11141 0.9005
R41361 PAD.n11456 PAD.n11184 0.9005
R41362 PAD.n11455 PAD.n11140 0.9005
R41363 PAD.n11454 PAD.n11186 0.9005
R41364 PAD.n11319 PAD.n11139 0.9005
R41365 PAD.n11450 PAD.n11188 0.9005
R41366 PAD.n11449 PAD.n11138 0.9005
R41367 PAD.n11448 PAD.n11190 0.9005
R41368 PAD.n11321 PAD.n11137 0.9005
R41369 PAD.n11444 PAD.n11192 0.9005
R41370 PAD.n11443 PAD.n11136 0.9005
R41371 PAD.n11442 PAD.n11194 0.9005
R41372 PAD.n11323 PAD.n11135 0.9005
R41373 PAD.n11438 PAD.n11196 0.9005
R41374 PAD.n11437 PAD.n11134 0.9005
R41375 PAD.n11436 PAD.n11198 0.9005
R41376 PAD.n11325 PAD.n11133 0.9005
R41377 PAD.n11432 PAD.n11200 0.9005
R41378 PAD.n11431 PAD.n11132 0.9005
R41379 PAD.n11430 PAD.n11202 0.9005
R41380 PAD.n11327 PAD.n11131 0.9005
R41381 PAD.n11426 PAD.n11204 0.9005
R41382 PAD.n11425 PAD.n11130 0.9005
R41383 PAD.n11424 PAD.n11206 0.9005
R41384 PAD.n11329 PAD.n11129 0.9005
R41385 PAD.n11420 PAD.n11208 0.9005
R41386 PAD.n11419 PAD.n11128 0.9005
R41387 PAD.n11418 PAD.n11210 0.9005
R41388 PAD.n11331 PAD.n11127 0.9005
R41389 PAD.n11414 PAD.n11212 0.9005
R41390 PAD.n11413 PAD.n11126 0.9005
R41391 PAD.n11412 PAD.n11214 0.9005
R41392 PAD.n11333 PAD.n11125 0.9005
R41393 PAD.n11408 PAD.n11216 0.9005
R41394 PAD.n11407 PAD.n11124 0.9005
R41395 PAD.n11406 PAD.n11218 0.9005
R41396 PAD.n11335 PAD.n11123 0.9005
R41397 PAD.n11402 PAD.n11220 0.9005
R41398 PAD.n11401 PAD.n11122 0.9005
R41399 PAD.n11400 PAD.n11222 0.9005
R41400 PAD.n11337 PAD.n11121 0.9005
R41401 PAD.n11396 PAD.n11224 0.9005
R41402 PAD.n11395 PAD.n11120 0.9005
R41403 PAD.n11394 PAD.n11226 0.9005
R41404 PAD.n11339 PAD.n11119 0.9005
R41405 PAD.n11390 PAD.n11228 0.9005
R41406 PAD.n11389 PAD.n11118 0.9005
R41407 PAD.n11388 PAD.n11230 0.9005
R41408 PAD.n11341 PAD.n11117 0.9005
R41409 PAD.n11384 PAD.n11232 0.9005
R41410 PAD.n11383 PAD.n11116 0.9005
R41411 PAD.n11382 PAD.n11234 0.9005
R41412 PAD.n11343 PAD.n11115 0.9005
R41413 PAD.n11378 PAD.n11236 0.9005
R41414 PAD.n11377 PAD.n11114 0.9005
R41415 PAD.n11376 PAD.n11238 0.9005
R41416 PAD.n11345 PAD.n11113 0.9005
R41417 PAD.n11372 PAD.n11240 0.9005
R41418 PAD.n11371 PAD.n11112 0.9005
R41419 PAD.n11370 PAD.n11242 0.9005
R41420 PAD.n11347 PAD.n11111 0.9005
R41421 PAD.n11366 PAD.n11244 0.9005
R41422 PAD.n11365 PAD.n11110 0.9005
R41423 PAD.n11364 PAD.n11246 0.9005
R41424 PAD.n11349 PAD.n11109 0.9005
R41425 PAD.n11360 PAD.n11248 0.9005
R41426 PAD.n11359 PAD.n11108 0.9005
R41427 PAD.n11358 PAD.n11250 0.9005
R41428 PAD.n11351 PAD.n11107 0.9005
R41429 PAD.n11354 PAD.n11252 0.9005
R41430 PAD.n11353 PAD.n11106 0.9005
R41431 PAD.n11508 PAD.n11506 0.9005
R41432 PAD.n11497 PAD.n11304 0.9005
R41433 PAD.n11496 PAD.n11495 0.9005
R41434 PAD.n11494 PAD.n11305 0.9005
R41435 PAD.n11493 PAD.n11492 0.9005
R41436 PAD.n11491 PAD.n11306 0.9005
R41437 PAD.n11490 PAD.n11489 0.9005
R41438 PAD.n11488 PAD.n11307 0.9005
R41439 PAD.n11487 PAD.n11486 0.9005
R41440 PAD.n11485 PAD.n11308 0.9005
R41441 PAD.n11484 PAD.n11483 0.9005
R41442 PAD.n11482 PAD.n11309 0.9005
R41443 PAD.n11481 PAD.n11480 0.9005
R41444 PAD.n11479 PAD.n11310 0.9005
R41445 PAD.n11478 PAD.n11477 0.9005
R41446 PAD.n11476 PAD.n11311 0.9005
R41447 PAD.n11475 PAD.n11474 0.9005
R41448 PAD.n11473 PAD.n11312 0.9005
R41449 PAD.n11472 PAD.n11471 0.9005
R41450 PAD.n11470 PAD.n11313 0.9005
R41451 PAD.n11469 PAD.n11468 0.9005
R41452 PAD.n11467 PAD.n11314 0.9005
R41453 PAD.n11466 PAD.n11465 0.9005
R41454 PAD.n11464 PAD.n11315 0.9005
R41455 PAD.n11463 PAD.n11462 0.9005
R41456 PAD.n11461 PAD.n11316 0.9005
R41457 PAD.n11460 PAD.n11459 0.9005
R41458 PAD.n11458 PAD.n11317 0.9005
R41459 PAD.n11457 PAD.n11456 0.9005
R41460 PAD.n11455 PAD.n11318 0.9005
R41461 PAD.n11454 PAD.n11453 0.9005
R41462 PAD.n11452 PAD.n11319 0.9005
R41463 PAD.n11451 PAD.n11450 0.9005
R41464 PAD.n11449 PAD.n11320 0.9005
R41465 PAD.n11448 PAD.n11447 0.9005
R41466 PAD.n11446 PAD.n11321 0.9005
R41467 PAD.n11445 PAD.n11444 0.9005
R41468 PAD.n11443 PAD.n11322 0.9005
R41469 PAD.n11442 PAD.n11441 0.9005
R41470 PAD.n11440 PAD.n11323 0.9005
R41471 PAD.n11439 PAD.n11438 0.9005
R41472 PAD.n11437 PAD.n11324 0.9005
R41473 PAD.n11436 PAD.n11435 0.9005
R41474 PAD.n11434 PAD.n11325 0.9005
R41475 PAD.n11433 PAD.n11432 0.9005
R41476 PAD.n11431 PAD.n11326 0.9005
R41477 PAD.n11430 PAD.n11429 0.9005
R41478 PAD.n11428 PAD.n11327 0.9005
R41479 PAD.n11427 PAD.n11426 0.9005
R41480 PAD.n11425 PAD.n11328 0.9005
R41481 PAD.n11424 PAD.n11423 0.9005
R41482 PAD.n11422 PAD.n11329 0.9005
R41483 PAD.n11421 PAD.n11420 0.9005
R41484 PAD.n11419 PAD.n11330 0.9005
R41485 PAD.n11418 PAD.n11417 0.9005
R41486 PAD.n11416 PAD.n11331 0.9005
R41487 PAD.n11415 PAD.n11414 0.9005
R41488 PAD.n11413 PAD.n11332 0.9005
R41489 PAD.n11412 PAD.n11411 0.9005
R41490 PAD.n11410 PAD.n11333 0.9005
R41491 PAD.n11409 PAD.n11408 0.9005
R41492 PAD.n11407 PAD.n11334 0.9005
R41493 PAD.n11406 PAD.n11405 0.9005
R41494 PAD.n11404 PAD.n11335 0.9005
R41495 PAD.n11403 PAD.n11402 0.9005
R41496 PAD.n11401 PAD.n11336 0.9005
R41497 PAD.n11400 PAD.n11399 0.9005
R41498 PAD.n11398 PAD.n11337 0.9005
R41499 PAD.n11397 PAD.n11396 0.9005
R41500 PAD.n11395 PAD.n11338 0.9005
R41501 PAD.n11394 PAD.n11393 0.9005
R41502 PAD.n11392 PAD.n11339 0.9005
R41503 PAD.n11391 PAD.n11390 0.9005
R41504 PAD.n11389 PAD.n11340 0.9005
R41505 PAD.n11388 PAD.n11387 0.9005
R41506 PAD.n11386 PAD.n11341 0.9005
R41507 PAD.n11385 PAD.n11384 0.9005
R41508 PAD.n11383 PAD.n11342 0.9005
R41509 PAD.n11382 PAD.n11381 0.9005
R41510 PAD.n11380 PAD.n11343 0.9005
R41511 PAD.n11379 PAD.n11378 0.9005
R41512 PAD.n11377 PAD.n11344 0.9005
R41513 PAD.n11376 PAD.n11375 0.9005
R41514 PAD.n11374 PAD.n11345 0.9005
R41515 PAD.n11373 PAD.n11372 0.9005
R41516 PAD.n11371 PAD.n11346 0.9005
R41517 PAD.n11370 PAD.n11369 0.9005
R41518 PAD.n11368 PAD.n11347 0.9005
R41519 PAD.n11367 PAD.n11366 0.9005
R41520 PAD.n11365 PAD.n11348 0.9005
R41521 PAD.n11364 PAD.n11363 0.9005
R41522 PAD.n11362 PAD.n11349 0.9005
R41523 PAD.n11361 PAD.n11360 0.9005
R41524 PAD.n11359 PAD.n11350 0.9005
R41525 PAD.n11358 PAD.n11357 0.9005
R41526 PAD.n11356 PAD.n11351 0.9005
R41527 PAD.n11355 PAD.n11354 0.9005
R41528 PAD.n11353 PAD.n11352 0.9005
R41529 PAD.n11499 PAD.n11498 0.9005
R41530 PAD.n6226 PAD.n6225 0.9005
R41531 PAD.n6227 PAD.n6224 0.9005
R41532 PAD.n6229 PAD.n6228 0.9005
R41533 PAD.n6230 PAD.n6223 0.9005
R41534 PAD.n6232 PAD.n6231 0.9005
R41535 PAD.n6233 PAD.n6222 0.9005
R41536 PAD.n6235 PAD.n6234 0.9005
R41537 PAD.n6236 PAD.n6221 0.9005
R41538 PAD.n6238 PAD.n6237 0.9005
R41539 PAD.n6239 PAD.n6220 0.9005
R41540 PAD.n6241 PAD.n6240 0.9005
R41541 PAD.n6242 PAD.n6219 0.9005
R41542 PAD.n6244 PAD.n6243 0.9005
R41543 PAD.n6245 PAD.n6218 0.9005
R41544 PAD.n6247 PAD.n6246 0.9005
R41545 PAD.n6248 PAD.n6217 0.9005
R41546 PAD.n6250 PAD.n6249 0.9005
R41547 PAD.n6251 PAD.n6216 0.9005
R41548 PAD.n6253 PAD.n6252 0.9005
R41549 PAD.n6254 PAD.n6215 0.9005
R41550 PAD.n6256 PAD.n6255 0.9005
R41551 PAD.n6257 PAD.n6214 0.9005
R41552 PAD.n6259 PAD.n6258 0.9005
R41553 PAD.n6260 PAD.n6213 0.9005
R41554 PAD.n6262 PAD.n6261 0.9005
R41555 PAD.n6263 PAD.n6212 0.9005
R41556 PAD.n6265 PAD.n6264 0.9005
R41557 PAD.n6266 PAD.n6211 0.9005
R41558 PAD.n6268 PAD.n6267 0.9005
R41559 PAD.n6269 PAD.n6210 0.9005
R41560 PAD.n6271 PAD.n6270 0.9005
R41561 PAD.n6272 PAD.n6209 0.9005
R41562 PAD.n6274 PAD.n6273 0.9005
R41563 PAD.n6275 PAD.n6208 0.9005
R41564 PAD.n6277 PAD.n6276 0.9005
R41565 PAD.n6278 PAD.n6207 0.9005
R41566 PAD.n6280 PAD.n6279 0.9005
R41567 PAD.n6281 PAD.n6206 0.9005
R41568 PAD.n6283 PAD.n6282 0.9005
R41569 PAD.n6284 PAD.n6205 0.9005
R41570 PAD.n6286 PAD.n6285 0.9005
R41571 PAD.n6287 PAD.n6204 0.9005
R41572 PAD.n6289 PAD.n6288 0.9005
R41573 PAD.n6290 PAD.n6203 0.9005
R41574 PAD.n6292 PAD.n6291 0.9005
R41575 PAD.n6293 PAD.n6202 0.9005
R41576 PAD.n6295 PAD.n6294 0.9005
R41577 PAD.n6296 PAD.n6201 0.9005
R41578 PAD.n6298 PAD.n6297 0.9005
R41579 PAD.n6299 PAD.n6200 0.9005
R41580 PAD.n6301 PAD.n6300 0.9005
R41581 PAD.n6302 PAD.n6199 0.9005
R41582 PAD.n6304 PAD.n6303 0.9005
R41583 PAD.n6305 PAD.n6198 0.9005
R41584 PAD.n6307 PAD.n6306 0.9005
R41585 PAD.n6308 PAD.n6197 0.9005
R41586 PAD.n6310 PAD.n6309 0.9005
R41587 PAD.n6311 PAD.n6196 0.9005
R41588 PAD.n6313 PAD.n6312 0.9005
R41589 PAD.n6314 PAD.n6195 0.9005
R41590 PAD.n6316 PAD.n6315 0.9005
R41591 PAD.n6317 PAD.n6194 0.9005
R41592 PAD.n6319 PAD.n6318 0.9005
R41593 PAD.n6320 PAD.n6193 0.9005
R41594 PAD.n6322 PAD.n6321 0.9005
R41595 PAD.n6323 PAD.n6192 0.9005
R41596 PAD.n6325 PAD.n6324 0.9005
R41597 PAD.n6326 PAD.n6191 0.9005
R41598 PAD.n6328 PAD.n6327 0.9005
R41599 PAD.n6329 PAD.n6190 0.9005
R41600 PAD.n6331 PAD.n6330 0.9005
R41601 PAD.n6332 PAD.n6189 0.9005
R41602 PAD.n6334 PAD.n6333 0.9005
R41603 PAD.n6335 PAD.n6188 0.9005
R41604 PAD.n6337 PAD.n6336 0.9005
R41605 PAD.n6338 PAD.n6187 0.9005
R41606 PAD.n6340 PAD.n6339 0.9005
R41607 PAD.n6341 PAD.n6186 0.9005
R41608 PAD.n6343 PAD.n6342 0.9005
R41609 PAD.n6344 PAD.n6185 0.9005
R41610 PAD.n6346 PAD.n6345 0.9005
R41611 PAD.n6347 PAD.n6184 0.9005
R41612 PAD.n6349 PAD.n6348 0.9005
R41613 PAD.n6350 PAD.n6183 0.9005
R41614 PAD.n6352 PAD.n6351 0.9005
R41615 PAD.n6353 PAD.n6182 0.9005
R41616 PAD.n6355 PAD.n6354 0.9005
R41617 PAD.n6356 PAD.n6181 0.9005
R41618 PAD.n6358 PAD.n6357 0.9005
R41619 PAD.n6359 PAD.n6180 0.9005
R41620 PAD.n6361 PAD.n6360 0.9005
R41621 PAD.n6362 PAD.n6179 0.9005
R41622 PAD.n6364 PAD.n6363 0.9005
R41623 PAD.n6365 PAD.n6178 0.9005
R41624 PAD.n6367 PAD.n6366 0.9005
R41625 PAD.n6368 PAD.n6177 0.9005
R41626 PAD.n6370 PAD.n6369 0.9005
R41627 PAD.n6371 PAD.n5978 0.9005
R41628 PAD.n6370 PAD.n6032 0.9005
R41629 PAD.n6226 PAD.n6034 0.9005
R41630 PAD.n6227 PAD.n6030 0.9005
R41631 PAD.n6228 PAD.n6037 0.9005
R41632 PAD.n6223 PAD.n6029 0.9005
R41633 PAD.n6232 PAD.n6040 0.9005
R41634 PAD.n6233 PAD.n6028 0.9005
R41635 PAD.n6234 PAD.n6043 0.9005
R41636 PAD.n6221 PAD.n6027 0.9005
R41637 PAD.n6238 PAD.n6046 0.9005
R41638 PAD.n6239 PAD.n6026 0.9005
R41639 PAD.n6240 PAD.n6049 0.9005
R41640 PAD.n6219 PAD.n6025 0.9005
R41641 PAD.n6244 PAD.n6052 0.9005
R41642 PAD.n6245 PAD.n6024 0.9005
R41643 PAD.n6246 PAD.n6055 0.9005
R41644 PAD.n6217 PAD.n6023 0.9005
R41645 PAD.n6250 PAD.n6058 0.9005
R41646 PAD.n6251 PAD.n6022 0.9005
R41647 PAD.n6252 PAD.n6061 0.9005
R41648 PAD.n6215 PAD.n6021 0.9005
R41649 PAD.n6256 PAD.n6064 0.9005
R41650 PAD.n6257 PAD.n6020 0.9005
R41651 PAD.n6258 PAD.n6067 0.9005
R41652 PAD.n6213 PAD.n6019 0.9005
R41653 PAD.n6262 PAD.n6070 0.9005
R41654 PAD.n6263 PAD.n6018 0.9005
R41655 PAD.n6264 PAD.n6073 0.9005
R41656 PAD.n6211 PAD.n6017 0.9005
R41657 PAD.n6268 PAD.n6076 0.9005
R41658 PAD.n6269 PAD.n6016 0.9005
R41659 PAD.n6270 PAD.n6079 0.9005
R41660 PAD.n6209 PAD.n6015 0.9005
R41661 PAD.n6274 PAD.n6082 0.9005
R41662 PAD.n6275 PAD.n6014 0.9005
R41663 PAD.n6276 PAD.n6085 0.9005
R41664 PAD.n6207 PAD.n6013 0.9005
R41665 PAD.n6280 PAD.n6088 0.9005
R41666 PAD.n6281 PAD.n6012 0.9005
R41667 PAD.n6282 PAD.n6091 0.9005
R41668 PAD.n6205 PAD.n6011 0.9005
R41669 PAD.n6286 PAD.n6094 0.9005
R41670 PAD.n6287 PAD.n6010 0.9005
R41671 PAD.n6288 PAD.n6097 0.9005
R41672 PAD.n6203 PAD.n6009 0.9005
R41673 PAD.n6292 PAD.n6100 0.9005
R41674 PAD.n6293 PAD.n6008 0.9005
R41675 PAD.n6294 PAD.n6103 0.9005
R41676 PAD.n6201 PAD.n6007 0.9005
R41677 PAD.n6298 PAD.n6106 0.9005
R41678 PAD.n6299 PAD.n6006 0.9005
R41679 PAD.n6300 PAD.n6109 0.9005
R41680 PAD.n6199 PAD.n6005 0.9005
R41681 PAD.n6304 PAD.n6112 0.9005
R41682 PAD.n6305 PAD.n6004 0.9005
R41683 PAD.n6306 PAD.n6115 0.9005
R41684 PAD.n6197 PAD.n6003 0.9005
R41685 PAD.n6310 PAD.n6118 0.9005
R41686 PAD.n6311 PAD.n6002 0.9005
R41687 PAD.n6312 PAD.n6121 0.9005
R41688 PAD.n6195 PAD.n6001 0.9005
R41689 PAD.n6316 PAD.n6124 0.9005
R41690 PAD.n6317 PAD.n6000 0.9005
R41691 PAD.n6318 PAD.n6127 0.9005
R41692 PAD.n6193 PAD.n5999 0.9005
R41693 PAD.n6322 PAD.n6130 0.9005
R41694 PAD.n6323 PAD.n5998 0.9005
R41695 PAD.n6324 PAD.n6133 0.9005
R41696 PAD.n6191 PAD.n5997 0.9005
R41697 PAD.n6328 PAD.n6136 0.9005
R41698 PAD.n6329 PAD.n5996 0.9005
R41699 PAD.n6330 PAD.n6139 0.9005
R41700 PAD.n6189 PAD.n5995 0.9005
R41701 PAD.n6334 PAD.n6142 0.9005
R41702 PAD.n6335 PAD.n5994 0.9005
R41703 PAD.n6336 PAD.n6145 0.9005
R41704 PAD.n6187 PAD.n5993 0.9005
R41705 PAD.n6340 PAD.n6148 0.9005
R41706 PAD.n6341 PAD.n5992 0.9005
R41707 PAD.n6342 PAD.n6151 0.9005
R41708 PAD.n6185 PAD.n5991 0.9005
R41709 PAD.n6346 PAD.n6154 0.9005
R41710 PAD.n6347 PAD.n5990 0.9005
R41711 PAD.n6348 PAD.n6157 0.9005
R41712 PAD.n6183 PAD.n5989 0.9005
R41713 PAD.n6352 PAD.n6160 0.9005
R41714 PAD.n6353 PAD.n5988 0.9005
R41715 PAD.n6354 PAD.n6163 0.9005
R41716 PAD.n6181 PAD.n5987 0.9005
R41717 PAD.n6358 PAD.n6166 0.9005
R41718 PAD.n6359 PAD.n5986 0.9005
R41719 PAD.n6360 PAD.n6169 0.9005
R41720 PAD.n6179 PAD.n5985 0.9005
R41721 PAD.n6364 PAD.n6172 0.9005
R41722 PAD.n6365 PAD.n5984 0.9005
R41723 PAD.n6366 PAD.n6175 0.9005
R41724 PAD.n6177 PAD.n5983 0.9005
R41725 PAD.n6372 PAD.n6371 0.9005
R41726 PAD.n6375 PAD.n6374 0.9005
R41727 PAD.n7809 PAD.n7808 0.87242
R41728 PAD.n11540 PAD.n11539 0.87242
R41729 PAD.n7810 PAD.n7809 0.79382
R41730 PAD.n3636 PAD.n10 0.79382
R41731 PAD.n11541 PAD.n11 0.79382
R41732 PAD.n11540 PAD.n12 0.79382
R41733 PAD.n11512 PAD.n11090 0.761105
R41734 PAD.n6385 PAD.n5956 0.758684
R41735 PAD.n11104 PAD.n11093 0.7505
R41736 PAD.n11515 PAD.n11514 0.7505
R41737 PAD.n11102 PAD.n11101 0.7505
R41738 PAD.n11516 PAD.n11515 0.7505
R41739 PAD.n11093 PAD.n11091 0.7505
R41740 PAD.n6389 PAD.n6388 0.7505
R41741 PAD.n5959 PAD.n5957 0.7505
R41742 PAD.n5969 PAD.n5959 0.7505
R41743 PAD.n6388 PAD.n6387 0.7505
R41744 PAD.n5968 PAD.n5967 0.7505
R41745 PAD.n10366 PAD.n13 0.408955
R41746 PAD.n9171 PAD.n9168 0.408955
R41747 PAD.n7812 PAD.n7811 0.408955
R41748 PAD.n8473 PAD.n3637 0.408866
R41749 PAD.n11517 PAD.n11090 0.384314
R41750 PAD.n6390 PAD.n5956 0.38336
R41751 PAD.n6 PAD.n5 0.204443
R41752 PAD.n1 PAD.n0 0.199354
R41753 PAD.n9 PAD.n3 0.102972
R41754 PAD PAD.n9 0.0996761
R41755 PAD PAD.n11542 0.09545
R41756 PAD.n1 PAD 0.0811609
R41757 PAD.n8 PAD 0.0811609
R41758 PAD.n7809 PAD.n10 0.0791
R41759 PAD.n11541 PAD.n11540 0.0791
R41760 PAD.n9 PAD.n8 0.0751609
R41761 PAD.n3 PAD 0.0548109
R41762 PAD.n6 PAD 0.0548109
R41763 PAD.n5 PAD 0.0548109
R41764 PAD.n3636 PAD.n11 0.0433318
R41765 PAD.n11542 PAD.n10 0.03995
R41766 PAD.n11542 PAD.n11541 0.03965
R41767 PAD.n7517 PAD.n7209 0.0380882
R41768 PAD.n7513 PAD.n7209 0.0380882
R41769 PAD.n7513 PAD.n7510 0.0380882
R41770 PAD.n7510 PAD.n7506 0.0380882
R41771 PAD.n7506 PAD.n7229 0.0380882
R41772 PAD.n7502 PAD.n7229 0.0380882
R41773 PAD.n7502 PAD.n7498 0.0380882
R41774 PAD.n7498 PAD.n7494 0.0380882
R41775 PAD.n7494 PAD.n7231 0.0380882
R41776 PAD.n7490 PAD.n7231 0.0380882
R41777 PAD.n7490 PAD.n7486 0.0380882
R41778 PAD.n7486 PAD.n7482 0.0380882
R41779 PAD.n7482 PAD.n7233 0.0380882
R41780 PAD.n7478 PAD.n7233 0.0380882
R41781 PAD.n7478 PAD.n7474 0.0380882
R41782 PAD.n7474 PAD.n7470 0.0380882
R41783 PAD.n7470 PAD.n7235 0.0380882
R41784 PAD.n7466 PAD.n7235 0.0380882
R41785 PAD.n7466 PAD.n7462 0.0380882
R41786 PAD.n7462 PAD.n7458 0.0380882
R41787 PAD.n7458 PAD.n7237 0.0380882
R41788 PAD.n7454 PAD.n7237 0.0380882
R41789 PAD.n7454 PAD.n7450 0.0380882
R41790 PAD.n7450 PAD.n7446 0.0380882
R41791 PAD.n7446 PAD.n7239 0.0380882
R41792 PAD.n7442 PAD.n7239 0.0380882
R41793 PAD.n7442 PAD.n7438 0.0380882
R41794 PAD.n7438 PAD.n7434 0.0380882
R41795 PAD.n7434 PAD.n7241 0.0380882
R41796 PAD.n7430 PAD.n7241 0.0380882
R41797 PAD.n7430 PAD.n7426 0.0380882
R41798 PAD.n7426 PAD.n7422 0.0380882
R41799 PAD.n7422 PAD.n7243 0.0380882
R41800 PAD.n7418 PAD.n7243 0.0380882
R41801 PAD.n7418 PAD.n7414 0.0380882
R41802 PAD.n7414 PAD.n7410 0.0380882
R41803 PAD.n7410 PAD.n7245 0.0380882
R41804 PAD.n7406 PAD.n7245 0.0380882
R41805 PAD.n7406 PAD.n7402 0.0380882
R41806 PAD.n7402 PAD.n7398 0.0380882
R41807 PAD.n7398 PAD.n7247 0.0380882
R41808 PAD.n7394 PAD.n7247 0.0380882
R41809 PAD.n7394 PAD.n7390 0.0380882
R41810 PAD.n7390 PAD.n7386 0.0380882
R41811 PAD.n7386 PAD.n7249 0.0380882
R41812 PAD.n7382 PAD.n7249 0.0380882
R41813 PAD.n7382 PAD.n7378 0.0380882
R41814 PAD.n7378 PAD.n7374 0.0380882
R41815 PAD.n7374 PAD.n7251 0.0380882
R41816 PAD.n7370 PAD.n7251 0.0380882
R41817 PAD.n7370 PAD.n7366 0.0380882
R41818 PAD.n7366 PAD.n7362 0.0380882
R41819 PAD.n7362 PAD.n7253 0.0380882
R41820 PAD.n7358 PAD.n7253 0.0380882
R41821 PAD.n7358 PAD.n7354 0.0380882
R41822 PAD.n7354 PAD.n7350 0.0380882
R41823 PAD.n7350 PAD.n7255 0.0380882
R41824 PAD.n7346 PAD.n7255 0.0380882
R41825 PAD.n7346 PAD.n7342 0.0380882
R41826 PAD.n7342 PAD.n7338 0.0380882
R41827 PAD.n7338 PAD.n7257 0.0380882
R41828 PAD.n7334 PAD.n7257 0.0380882
R41829 PAD.n7334 PAD.n7330 0.0380882
R41830 PAD.n7330 PAD.n7326 0.0380882
R41831 PAD.n7326 PAD.n7259 0.0380882
R41832 PAD.n7322 PAD.n7259 0.0380882
R41833 PAD.n7322 PAD.n7318 0.0380882
R41834 PAD.n7318 PAD.n7314 0.0380882
R41835 PAD.n7314 PAD.n7261 0.0380882
R41836 PAD.n7310 PAD.n7261 0.0380882
R41837 PAD.n7310 PAD.n7306 0.0380882
R41838 PAD.n7306 PAD.n7302 0.0380882
R41839 PAD.n7302 PAD.n7263 0.0380882
R41840 PAD.n7298 PAD.n7263 0.0380882
R41841 PAD.n7298 PAD.n7294 0.0380882
R41842 PAD.n7294 PAD.n7290 0.0380882
R41843 PAD.n7290 PAD.n7265 0.0380882
R41844 PAD.n7286 PAD.n7265 0.0380882
R41845 PAD.n7286 PAD.n7282 0.0380882
R41846 PAD.n7282 PAD.n7278 0.0380882
R41847 PAD.n7278 PAD.n7267 0.0380882
R41848 PAD.n7274 PAD.n7267 0.0380882
R41849 PAD.n7274 PAD.n7270 0.0380882
R41850 PAD.n7516 PAD.n7515 0.0380882
R41851 PAD.n7515 PAD.n7514 0.0380882
R41852 PAD.n7514 PAD.n7228 0.0380882
R41853 PAD.n7505 PAD.n7228 0.0380882
R41854 PAD.n7505 PAD.n7504 0.0380882
R41855 PAD.n7504 PAD.n7503 0.0380882
R41856 PAD.n7503 PAD.n7230 0.0380882
R41857 PAD.n7493 PAD.n7230 0.0380882
R41858 PAD.n7493 PAD.n7492 0.0380882
R41859 PAD.n7492 PAD.n7491 0.0380882
R41860 PAD.n7491 PAD.n7232 0.0380882
R41861 PAD.n7481 PAD.n7232 0.0380882
R41862 PAD.n7481 PAD.n7480 0.0380882
R41863 PAD.n7480 PAD.n7479 0.0380882
R41864 PAD.n7479 PAD.n7234 0.0380882
R41865 PAD.n7469 PAD.n7234 0.0380882
R41866 PAD.n7469 PAD.n7468 0.0380882
R41867 PAD.n7468 PAD.n7467 0.0380882
R41868 PAD.n7467 PAD.n7236 0.0380882
R41869 PAD.n7457 PAD.n7236 0.0380882
R41870 PAD.n7457 PAD.n7456 0.0380882
R41871 PAD.n7456 PAD.n7455 0.0380882
R41872 PAD.n7455 PAD.n7238 0.0380882
R41873 PAD.n7445 PAD.n7238 0.0380882
R41874 PAD.n7445 PAD.n7444 0.0380882
R41875 PAD.n7444 PAD.n7443 0.0380882
R41876 PAD.n7443 PAD.n7240 0.0380882
R41877 PAD.n7433 PAD.n7240 0.0380882
R41878 PAD.n7433 PAD.n7432 0.0380882
R41879 PAD.n7432 PAD.n7431 0.0380882
R41880 PAD.n7431 PAD.n7242 0.0380882
R41881 PAD.n7421 PAD.n7242 0.0380882
R41882 PAD.n7421 PAD.n7420 0.0380882
R41883 PAD.n7420 PAD.n7419 0.0380882
R41884 PAD.n7419 PAD.n7244 0.0380882
R41885 PAD.n7409 PAD.n7244 0.0380882
R41886 PAD.n7409 PAD.n7408 0.0380882
R41887 PAD.n7408 PAD.n7407 0.0380882
R41888 PAD.n7407 PAD.n7246 0.0380882
R41889 PAD.n7397 PAD.n7246 0.0380882
R41890 PAD.n7397 PAD.n7396 0.0380882
R41891 PAD.n7396 PAD.n7395 0.0380882
R41892 PAD.n7395 PAD.n7248 0.0380882
R41893 PAD.n7385 PAD.n7248 0.0380882
R41894 PAD.n7385 PAD.n7384 0.0380882
R41895 PAD.n7384 PAD.n7383 0.0380882
R41896 PAD.n7383 PAD.n7250 0.0380882
R41897 PAD.n7373 PAD.n7250 0.0380882
R41898 PAD.n7373 PAD.n7372 0.0380882
R41899 PAD.n7372 PAD.n7371 0.0380882
R41900 PAD.n7371 PAD.n7252 0.0380882
R41901 PAD.n7361 PAD.n7252 0.0380882
R41902 PAD.n7361 PAD.n7360 0.0380882
R41903 PAD.n7360 PAD.n7359 0.0380882
R41904 PAD.n7359 PAD.n7254 0.0380882
R41905 PAD.n7349 PAD.n7254 0.0380882
R41906 PAD.n7349 PAD.n7348 0.0380882
R41907 PAD.n7348 PAD.n7347 0.0380882
R41908 PAD.n7347 PAD.n7256 0.0380882
R41909 PAD.n7337 PAD.n7256 0.0380882
R41910 PAD.n7337 PAD.n7336 0.0380882
R41911 PAD.n7336 PAD.n7335 0.0380882
R41912 PAD.n7335 PAD.n7258 0.0380882
R41913 PAD.n7325 PAD.n7258 0.0380882
R41914 PAD.n7325 PAD.n7324 0.0380882
R41915 PAD.n7324 PAD.n7323 0.0380882
R41916 PAD.n7323 PAD.n7260 0.0380882
R41917 PAD.n7313 PAD.n7260 0.0380882
R41918 PAD.n7313 PAD.n7312 0.0380882
R41919 PAD.n7312 PAD.n7311 0.0380882
R41920 PAD.n7311 PAD.n7262 0.0380882
R41921 PAD.n7301 PAD.n7262 0.0380882
R41922 PAD.n7301 PAD.n7300 0.0380882
R41923 PAD.n7300 PAD.n7299 0.0380882
R41924 PAD.n7299 PAD.n7264 0.0380882
R41925 PAD.n7289 PAD.n7264 0.0380882
R41926 PAD.n7289 PAD.n7288 0.0380882
R41927 PAD.n7288 PAD.n7287 0.0380882
R41928 PAD.n7287 PAD.n7266 0.0380882
R41929 PAD.n7277 PAD.n7266 0.0380882
R41930 PAD.n7277 PAD.n7276 0.0380882
R41931 PAD.n7276 PAD.n7275 0.0380882
R41932 PAD.n7275 PAD.n7268 0.0380882
R41933 PAD.n121 PAD.n120 0.0380882
R41934 PAD.n122 PAD.n121 0.0380882
R41935 PAD.n122 PAD.n115 0.0380882
R41936 PAD.n132 PAD.n115 0.0380882
R41937 PAD.n133 PAD.n132 0.0380882
R41938 PAD.n134 PAD.n133 0.0380882
R41939 PAD.n134 PAD.n113 0.0380882
R41940 PAD.n144 PAD.n113 0.0380882
R41941 PAD.n145 PAD.n144 0.0380882
R41942 PAD.n146 PAD.n145 0.0380882
R41943 PAD.n146 PAD.n111 0.0380882
R41944 PAD.n156 PAD.n111 0.0380882
R41945 PAD.n157 PAD.n156 0.0380882
R41946 PAD.n158 PAD.n157 0.0380882
R41947 PAD.n158 PAD.n109 0.0380882
R41948 PAD.n168 PAD.n109 0.0380882
R41949 PAD.n169 PAD.n168 0.0380882
R41950 PAD.n170 PAD.n169 0.0380882
R41951 PAD.n170 PAD.n107 0.0380882
R41952 PAD.n180 PAD.n107 0.0380882
R41953 PAD.n181 PAD.n180 0.0380882
R41954 PAD.n182 PAD.n181 0.0380882
R41955 PAD.n182 PAD.n105 0.0380882
R41956 PAD.n192 PAD.n105 0.0380882
R41957 PAD.n193 PAD.n192 0.0380882
R41958 PAD.n194 PAD.n193 0.0380882
R41959 PAD.n194 PAD.n103 0.0380882
R41960 PAD.n204 PAD.n103 0.0380882
R41961 PAD.n205 PAD.n204 0.0380882
R41962 PAD.n206 PAD.n205 0.0380882
R41963 PAD.n206 PAD.n101 0.0380882
R41964 PAD.n216 PAD.n101 0.0380882
R41965 PAD.n217 PAD.n216 0.0380882
R41966 PAD.n218 PAD.n217 0.0380882
R41967 PAD.n218 PAD.n99 0.0380882
R41968 PAD.n228 PAD.n99 0.0380882
R41969 PAD.n229 PAD.n228 0.0380882
R41970 PAD.n230 PAD.n229 0.0380882
R41971 PAD.n230 PAD.n97 0.0380882
R41972 PAD.n240 PAD.n97 0.0380882
R41973 PAD.n241 PAD.n240 0.0380882
R41974 PAD.n242 PAD.n241 0.0380882
R41975 PAD.n242 PAD.n95 0.0380882
R41976 PAD.n252 PAD.n95 0.0380882
R41977 PAD.n253 PAD.n252 0.0380882
R41978 PAD.n254 PAD.n253 0.0380882
R41979 PAD.n254 PAD.n93 0.0380882
R41980 PAD.n264 PAD.n93 0.0380882
R41981 PAD.n265 PAD.n264 0.0380882
R41982 PAD.n266 PAD.n265 0.0380882
R41983 PAD.n266 PAD.n91 0.0380882
R41984 PAD.n276 PAD.n91 0.0380882
R41985 PAD.n277 PAD.n276 0.0380882
R41986 PAD.n278 PAD.n277 0.0380882
R41987 PAD.n278 PAD.n89 0.0380882
R41988 PAD.n288 PAD.n89 0.0380882
R41989 PAD.n289 PAD.n288 0.0380882
R41990 PAD.n290 PAD.n289 0.0380882
R41991 PAD.n290 PAD.n87 0.0380882
R41992 PAD.n300 PAD.n87 0.0380882
R41993 PAD.n301 PAD.n300 0.0380882
R41994 PAD.n302 PAD.n301 0.0380882
R41995 PAD.n302 PAD.n85 0.0380882
R41996 PAD.n312 PAD.n85 0.0380882
R41997 PAD.n313 PAD.n312 0.0380882
R41998 PAD.n314 PAD.n313 0.0380882
R41999 PAD.n314 PAD.n83 0.0380882
R42000 PAD.n324 PAD.n83 0.0380882
R42001 PAD.n325 PAD.n324 0.0380882
R42002 PAD.n326 PAD.n325 0.0380882
R42003 PAD.n326 PAD.n81 0.0380882
R42004 PAD.n336 PAD.n81 0.0380882
R42005 PAD.n337 PAD.n336 0.0380882
R42006 PAD.n338 PAD.n337 0.0380882
R42007 PAD.n338 PAD.n79 0.0380882
R42008 PAD.n348 PAD.n79 0.0380882
R42009 PAD.n349 PAD.n348 0.0380882
R42010 PAD.n350 PAD.n349 0.0380882
R42011 PAD.n350 PAD.n77 0.0380882
R42012 PAD.n360 PAD.n77 0.0380882
R42013 PAD.n361 PAD.n360 0.0380882
R42014 PAD.n362 PAD.n361 0.0380882
R42015 PAD.n362 PAD.n26 0.0380882
R42016 PAD.n10695 PAD.n10694 0.0380882
R42017 PAD.n10694 PAD.n10691 0.0380882
R42018 PAD.n10691 PAD.n10414 0.0380882
R42019 PAD.n10687 PAD.n10414 0.0380882
R42020 PAD.n10687 PAD.n10683 0.0380882
R42021 PAD.n10683 PAD.n10682 0.0380882
R42022 PAD.n10682 PAD.n10419 0.0380882
R42023 PAD.n10678 PAD.n10419 0.0380882
R42024 PAD.n10678 PAD.n10674 0.0380882
R42025 PAD.n10674 PAD.n10673 0.0380882
R42026 PAD.n10673 PAD.n10424 0.0380882
R42027 PAD.n10669 PAD.n10424 0.0380882
R42028 PAD.n10669 PAD.n10665 0.0380882
R42029 PAD.n10665 PAD.n10664 0.0380882
R42030 PAD.n10664 PAD.n10429 0.0380882
R42031 PAD.n10660 PAD.n10429 0.0380882
R42032 PAD.n10660 PAD.n10656 0.0380882
R42033 PAD.n10656 PAD.n10655 0.0380882
R42034 PAD.n10655 PAD.n10434 0.0380882
R42035 PAD.n10651 PAD.n10434 0.0380882
R42036 PAD.n10651 PAD.n10647 0.0380882
R42037 PAD.n10647 PAD.n10646 0.0380882
R42038 PAD.n10646 PAD.n10439 0.0380882
R42039 PAD.n10642 PAD.n10439 0.0380882
R42040 PAD.n10642 PAD.n10638 0.0380882
R42041 PAD.n10638 PAD.n10637 0.0380882
R42042 PAD.n10637 PAD.n10444 0.0380882
R42043 PAD.n10633 PAD.n10444 0.0380882
R42044 PAD.n10633 PAD.n10629 0.0380882
R42045 PAD.n10629 PAD.n10628 0.0380882
R42046 PAD.n10628 PAD.n10449 0.0380882
R42047 PAD.n10624 PAD.n10449 0.0380882
R42048 PAD.n10624 PAD.n10620 0.0380882
R42049 PAD.n10620 PAD.n10619 0.0380882
R42050 PAD.n10619 PAD.n10454 0.0380882
R42051 PAD.n10615 PAD.n10454 0.0380882
R42052 PAD.n10615 PAD.n10611 0.0380882
R42053 PAD.n10611 PAD.n10610 0.0380882
R42054 PAD.n10610 PAD.n10459 0.0380882
R42055 PAD.n10606 PAD.n10459 0.0380882
R42056 PAD.n10606 PAD.n10602 0.0380882
R42057 PAD.n10602 PAD.n10601 0.0380882
R42058 PAD.n10601 PAD.n10464 0.0380882
R42059 PAD.n10597 PAD.n10464 0.0380882
R42060 PAD.n10597 PAD.n10593 0.0380882
R42061 PAD.n10593 PAD.n10592 0.0380882
R42062 PAD.n10592 PAD.n10469 0.0380882
R42063 PAD.n10588 PAD.n10469 0.0380882
R42064 PAD.n10588 PAD.n10584 0.0380882
R42065 PAD.n10584 PAD.n10583 0.0380882
R42066 PAD.n10583 PAD.n10474 0.0380882
R42067 PAD.n10579 PAD.n10474 0.0380882
R42068 PAD.n10579 PAD.n10575 0.0380882
R42069 PAD.n10575 PAD.n10574 0.0380882
R42070 PAD.n10574 PAD.n10479 0.0380882
R42071 PAD.n10570 PAD.n10479 0.0380882
R42072 PAD.n10570 PAD.n10566 0.0380882
R42073 PAD.n10566 PAD.n10565 0.0380882
R42074 PAD.n10565 PAD.n10484 0.0380882
R42075 PAD.n10561 PAD.n10484 0.0380882
R42076 PAD.n10561 PAD.n10557 0.0380882
R42077 PAD.n10557 PAD.n10556 0.0380882
R42078 PAD.n10556 PAD.n10489 0.0380882
R42079 PAD.n10552 PAD.n10489 0.0380882
R42080 PAD.n10552 PAD.n10548 0.0380882
R42081 PAD.n10548 PAD.n10547 0.0380882
R42082 PAD.n10547 PAD.n10494 0.0380882
R42083 PAD.n10543 PAD.n10494 0.0380882
R42084 PAD.n10543 PAD.n10539 0.0380882
R42085 PAD.n10539 PAD.n10538 0.0380882
R42086 PAD.n10538 PAD.n10499 0.0380882
R42087 PAD.n10534 PAD.n10499 0.0380882
R42088 PAD.n10534 PAD.n10530 0.0380882
R42089 PAD.n10530 PAD.n10529 0.0380882
R42090 PAD.n10529 PAD.n10504 0.0380882
R42091 PAD.n10525 PAD.n10504 0.0380882
R42092 PAD.n10525 PAD.n10521 0.0380882
R42093 PAD.n10521 PAD.n10520 0.0380882
R42094 PAD.n10520 PAD.n10509 0.0380882
R42095 PAD.n10516 PAD.n10509 0.0380882
R42096 PAD.n10516 PAD.n420 0.0380882
R42097 PAD.n10712 PAD.n420 0.0380882
R42098 PAD.n10712 PAD.n416 0.0380882
R42099 PAD.n10696 PAD.n10413 0.0380882
R42100 PAD.n10690 PAD.n10413 0.0380882
R42101 PAD.n10690 PAD.n10689 0.0380882
R42102 PAD.n10689 PAD.n10688 0.0380882
R42103 PAD.n10688 PAD.n10418 0.0380882
R42104 PAD.n10681 PAD.n10418 0.0380882
R42105 PAD.n10681 PAD.n10680 0.0380882
R42106 PAD.n10680 PAD.n10679 0.0380882
R42107 PAD.n10679 PAD.n10423 0.0380882
R42108 PAD.n10672 PAD.n10423 0.0380882
R42109 PAD.n10672 PAD.n10671 0.0380882
R42110 PAD.n10671 PAD.n10670 0.0380882
R42111 PAD.n10670 PAD.n10428 0.0380882
R42112 PAD.n10663 PAD.n10428 0.0380882
R42113 PAD.n10663 PAD.n10662 0.0380882
R42114 PAD.n10662 PAD.n10661 0.0380882
R42115 PAD.n10661 PAD.n10433 0.0380882
R42116 PAD.n10654 PAD.n10433 0.0380882
R42117 PAD.n10654 PAD.n10653 0.0380882
R42118 PAD.n10653 PAD.n10652 0.0380882
R42119 PAD.n10652 PAD.n10438 0.0380882
R42120 PAD.n10645 PAD.n10438 0.0380882
R42121 PAD.n10645 PAD.n10644 0.0380882
R42122 PAD.n10644 PAD.n10643 0.0380882
R42123 PAD.n10643 PAD.n10443 0.0380882
R42124 PAD.n10636 PAD.n10443 0.0380882
R42125 PAD.n10636 PAD.n10635 0.0380882
R42126 PAD.n10635 PAD.n10634 0.0380882
R42127 PAD.n10634 PAD.n10448 0.0380882
R42128 PAD.n10627 PAD.n10448 0.0380882
R42129 PAD.n10627 PAD.n10626 0.0380882
R42130 PAD.n10626 PAD.n10625 0.0380882
R42131 PAD.n10625 PAD.n10453 0.0380882
R42132 PAD.n10618 PAD.n10453 0.0380882
R42133 PAD.n10618 PAD.n10617 0.0380882
R42134 PAD.n10617 PAD.n10616 0.0380882
R42135 PAD.n10616 PAD.n10458 0.0380882
R42136 PAD.n10609 PAD.n10458 0.0380882
R42137 PAD.n10609 PAD.n10608 0.0380882
R42138 PAD.n10608 PAD.n10607 0.0380882
R42139 PAD.n10607 PAD.n10463 0.0380882
R42140 PAD.n10600 PAD.n10463 0.0380882
R42141 PAD.n10600 PAD.n10599 0.0380882
R42142 PAD.n10599 PAD.n10598 0.0380882
R42143 PAD.n10598 PAD.n10468 0.0380882
R42144 PAD.n10591 PAD.n10468 0.0380882
R42145 PAD.n10591 PAD.n10590 0.0380882
R42146 PAD.n10590 PAD.n10589 0.0380882
R42147 PAD.n10589 PAD.n10473 0.0380882
R42148 PAD.n10582 PAD.n10473 0.0380882
R42149 PAD.n10582 PAD.n10581 0.0380882
R42150 PAD.n10581 PAD.n10580 0.0380882
R42151 PAD.n10580 PAD.n10478 0.0380882
R42152 PAD.n10573 PAD.n10478 0.0380882
R42153 PAD.n10573 PAD.n10572 0.0380882
R42154 PAD.n10572 PAD.n10571 0.0380882
R42155 PAD.n10571 PAD.n10483 0.0380882
R42156 PAD.n10564 PAD.n10483 0.0380882
R42157 PAD.n10564 PAD.n10563 0.0380882
R42158 PAD.n10563 PAD.n10562 0.0380882
R42159 PAD.n10562 PAD.n10488 0.0380882
R42160 PAD.n10555 PAD.n10488 0.0380882
R42161 PAD.n10555 PAD.n10554 0.0380882
R42162 PAD.n10554 PAD.n10553 0.0380882
R42163 PAD.n10553 PAD.n10493 0.0380882
R42164 PAD.n10546 PAD.n10493 0.0380882
R42165 PAD.n10546 PAD.n10545 0.0380882
R42166 PAD.n10545 PAD.n10544 0.0380882
R42167 PAD.n10544 PAD.n10498 0.0380882
R42168 PAD.n10537 PAD.n10498 0.0380882
R42169 PAD.n10537 PAD.n10536 0.0380882
R42170 PAD.n10536 PAD.n10535 0.0380882
R42171 PAD.n10535 PAD.n10503 0.0380882
R42172 PAD.n10528 PAD.n10503 0.0380882
R42173 PAD.n10528 PAD.n10527 0.0380882
R42174 PAD.n10527 PAD.n10526 0.0380882
R42175 PAD.n10526 PAD.n10508 0.0380882
R42176 PAD.n10519 PAD.n10508 0.0380882
R42177 PAD.n10519 PAD.n10518 0.0380882
R42178 PAD.n10518 PAD.n10517 0.0380882
R42179 PAD.n10517 PAD.n421 0.0380882
R42180 PAD.n10711 PAD.n421 0.0380882
R42181 PAD.n10711 PAD.n10710 0.0380882
R42182 PAD.n522 PAD.n520 0.0380882
R42183 PAD.n530 PAD.n520 0.0380882
R42184 PAD.n530 PAD.n518 0.0380882
R42185 PAD.n534 PAD.n518 0.0380882
R42186 PAD.n534 PAD.n516 0.0380882
R42187 PAD.n542 PAD.n516 0.0380882
R42188 PAD.n542 PAD.n514 0.0380882
R42189 PAD.n546 PAD.n514 0.0380882
R42190 PAD.n546 PAD.n512 0.0380882
R42191 PAD.n554 PAD.n512 0.0380882
R42192 PAD.n554 PAD.n510 0.0380882
R42193 PAD.n558 PAD.n510 0.0380882
R42194 PAD.n558 PAD.n508 0.0380882
R42195 PAD.n566 PAD.n508 0.0380882
R42196 PAD.n566 PAD.n506 0.0380882
R42197 PAD.n570 PAD.n506 0.0380882
R42198 PAD.n570 PAD.n504 0.0380882
R42199 PAD.n578 PAD.n504 0.0380882
R42200 PAD.n578 PAD.n502 0.0380882
R42201 PAD.n582 PAD.n502 0.0380882
R42202 PAD.n582 PAD.n500 0.0380882
R42203 PAD.n590 PAD.n500 0.0380882
R42204 PAD.n590 PAD.n498 0.0380882
R42205 PAD.n594 PAD.n498 0.0380882
R42206 PAD.n594 PAD.n496 0.0380882
R42207 PAD.n602 PAD.n496 0.0380882
R42208 PAD.n602 PAD.n494 0.0380882
R42209 PAD.n606 PAD.n494 0.0380882
R42210 PAD.n606 PAD.n492 0.0380882
R42211 PAD.n614 PAD.n492 0.0380882
R42212 PAD.n614 PAD.n490 0.0380882
R42213 PAD.n618 PAD.n490 0.0380882
R42214 PAD.n618 PAD.n488 0.0380882
R42215 PAD.n626 PAD.n488 0.0380882
R42216 PAD.n626 PAD.n486 0.0380882
R42217 PAD.n630 PAD.n486 0.0380882
R42218 PAD.n630 PAD.n484 0.0380882
R42219 PAD.n638 PAD.n484 0.0380882
R42220 PAD.n638 PAD.n482 0.0380882
R42221 PAD.n642 PAD.n482 0.0380882
R42222 PAD.n642 PAD.n480 0.0380882
R42223 PAD.n650 PAD.n480 0.0380882
R42224 PAD.n650 PAD.n478 0.0380882
R42225 PAD.n654 PAD.n478 0.0380882
R42226 PAD.n654 PAD.n476 0.0380882
R42227 PAD.n662 PAD.n476 0.0380882
R42228 PAD.n662 PAD.n474 0.0380882
R42229 PAD.n666 PAD.n474 0.0380882
R42230 PAD.n666 PAD.n472 0.0380882
R42231 PAD.n674 PAD.n472 0.0380882
R42232 PAD.n674 PAD.n470 0.0380882
R42233 PAD.n678 PAD.n470 0.0380882
R42234 PAD.n678 PAD.n468 0.0380882
R42235 PAD.n686 PAD.n468 0.0380882
R42236 PAD.n686 PAD.n466 0.0380882
R42237 PAD.n690 PAD.n466 0.0380882
R42238 PAD.n690 PAD.n464 0.0380882
R42239 PAD.n698 PAD.n464 0.0380882
R42240 PAD.n698 PAD.n462 0.0380882
R42241 PAD.n702 PAD.n462 0.0380882
R42242 PAD.n702 PAD.n460 0.0380882
R42243 PAD.n710 PAD.n460 0.0380882
R42244 PAD.n710 PAD.n458 0.0380882
R42245 PAD.n714 PAD.n458 0.0380882
R42246 PAD.n714 PAD.n456 0.0380882
R42247 PAD.n722 PAD.n456 0.0380882
R42248 PAD.n722 PAD.n454 0.0380882
R42249 PAD.n726 PAD.n454 0.0380882
R42250 PAD.n726 PAD.n452 0.0380882
R42251 PAD.n734 PAD.n452 0.0380882
R42252 PAD.n734 PAD.n450 0.0380882
R42253 PAD.n738 PAD.n450 0.0380882
R42254 PAD.n738 PAD.n448 0.0380882
R42255 PAD.n746 PAD.n448 0.0380882
R42256 PAD.n746 PAD.n446 0.0380882
R42257 PAD.n750 PAD.n446 0.0380882
R42258 PAD.n750 PAD.n444 0.0380882
R42259 PAD.n758 PAD.n444 0.0380882
R42260 PAD.n758 PAD.n442 0.0380882
R42261 PAD.n763 PAD.n442 0.0380882
R42262 PAD.n763 PAD.n440 0.0380882
R42263 PAD.n440 PAD.n439 0.0380882
R42264 PAD.n771 PAD.n439 0.0380882
R42265 PAD.n521 PAD.n519 0.0380882
R42266 PAD.n531 PAD.n519 0.0380882
R42267 PAD.n532 PAD.n531 0.0380882
R42268 PAD.n533 PAD.n532 0.0380882
R42269 PAD.n533 PAD.n515 0.0380882
R42270 PAD.n543 PAD.n515 0.0380882
R42271 PAD.n544 PAD.n543 0.0380882
R42272 PAD.n545 PAD.n544 0.0380882
R42273 PAD.n545 PAD.n511 0.0380882
R42274 PAD.n555 PAD.n511 0.0380882
R42275 PAD.n556 PAD.n555 0.0380882
R42276 PAD.n557 PAD.n556 0.0380882
R42277 PAD.n557 PAD.n507 0.0380882
R42278 PAD.n567 PAD.n507 0.0380882
R42279 PAD.n568 PAD.n567 0.0380882
R42280 PAD.n569 PAD.n568 0.0380882
R42281 PAD.n569 PAD.n503 0.0380882
R42282 PAD.n579 PAD.n503 0.0380882
R42283 PAD.n580 PAD.n579 0.0380882
R42284 PAD.n581 PAD.n580 0.0380882
R42285 PAD.n581 PAD.n499 0.0380882
R42286 PAD.n591 PAD.n499 0.0380882
R42287 PAD.n592 PAD.n591 0.0380882
R42288 PAD.n593 PAD.n592 0.0380882
R42289 PAD.n593 PAD.n495 0.0380882
R42290 PAD.n603 PAD.n495 0.0380882
R42291 PAD.n604 PAD.n603 0.0380882
R42292 PAD.n605 PAD.n604 0.0380882
R42293 PAD.n605 PAD.n491 0.0380882
R42294 PAD.n615 PAD.n491 0.0380882
R42295 PAD.n616 PAD.n615 0.0380882
R42296 PAD.n617 PAD.n616 0.0380882
R42297 PAD.n617 PAD.n487 0.0380882
R42298 PAD.n627 PAD.n487 0.0380882
R42299 PAD.n628 PAD.n627 0.0380882
R42300 PAD.n629 PAD.n628 0.0380882
R42301 PAD.n629 PAD.n483 0.0380882
R42302 PAD.n639 PAD.n483 0.0380882
R42303 PAD.n640 PAD.n639 0.0380882
R42304 PAD.n641 PAD.n640 0.0380882
R42305 PAD.n641 PAD.n479 0.0380882
R42306 PAD.n651 PAD.n479 0.0380882
R42307 PAD.n652 PAD.n651 0.0380882
R42308 PAD.n653 PAD.n652 0.0380882
R42309 PAD.n653 PAD.n475 0.0380882
R42310 PAD.n663 PAD.n475 0.0380882
R42311 PAD.n664 PAD.n663 0.0380882
R42312 PAD.n665 PAD.n664 0.0380882
R42313 PAD.n665 PAD.n471 0.0380882
R42314 PAD.n675 PAD.n471 0.0380882
R42315 PAD.n676 PAD.n675 0.0380882
R42316 PAD.n677 PAD.n676 0.0380882
R42317 PAD.n677 PAD.n467 0.0380882
R42318 PAD.n687 PAD.n467 0.0380882
R42319 PAD.n688 PAD.n687 0.0380882
R42320 PAD.n689 PAD.n688 0.0380882
R42321 PAD.n689 PAD.n463 0.0380882
R42322 PAD.n699 PAD.n463 0.0380882
R42323 PAD.n700 PAD.n699 0.0380882
R42324 PAD.n701 PAD.n700 0.0380882
R42325 PAD.n701 PAD.n459 0.0380882
R42326 PAD.n711 PAD.n459 0.0380882
R42327 PAD.n712 PAD.n711 0.0380882
R42328 PAD.n713 PAD.n712 0.0380882
R42329 PAD.n713 PAD.n455 0.0380882
R42330 PAD.n723 PAD.n455 0.0380882
R42331 PAD.n724 PAD.n723 0.0380882
R42332 PAD.n725 PAD.n724 0.0380882
R42333 PAD.n725 PAD.n451 0.0380882
R42334 PAD.n735 PAD.n451 0.0380882
R42335 PAD.n736 PAD.n735 0.0380882
R42336 PAD.n737 PAD.n736 0.0380882
R42337 PAD.n737 PAD.n447 0.0380882
R42338 PAD.n747 PAD.n447 0.0380882
R42339 PAD.n748 PAD.n747 0.0380882
R42340 PAD.n749 PAD.n748 0.0380882
R42341 PAD.n749 PAD.n443 0.0380882
R42342 PAD.n759 PAD.n443 0.0380882
R42343 PAD.n760 PAD.n759 0.0380882
R42344 PAD.n762 PAD.n760 0.0380882
R42345 PAD.n762 PAD.n761 0.0380882
R42346 PAD.n761 PAD.n438 0.0380882
R42347 PAD.n772 PAD.n438 0.0380882
R42348 PAD.n872 PAD.n871 0.0380882
R42349 PAD.n876 PAD.n871 0.0380882
R42350 PAD.n880 PAD.n876 0.0380882
R42351 PAD.n884 PAD.n880 0.0380882
R42352 PAD.n884 PAD.n867 0.0380882
R42353 PAD.n888 PAD.n867 0.0380882
R42354 PAD.n892 PAD.n888 0.0380882
R42355 PAD.n896 PAD.n892 0.0380882
R42356 PAD.n896 PAD.n865 0.0380882
R42357 PAD.n900 PAD.n865 0.0380882
R42358 PAD.n904 PAD.n900 0.0380882
R42359 PAD.n908 PAD.n904 0.0380882
R42360 PAD.n908 PAD.n863 0.0380882
R42361 PAD.n912 PAD.n863 0.0380882
R42362 PAD.n916 PAD.n912 0.0380882
R42363 PAD.n920 PAD.n916 0.0380882
R42364 PAD.n920 PAD.n861 0.0380882
R42365 PAD.n924 PAD.n861 0.0380882
R42366 PAD.n928 PAD.n924 0.0380882
R42367 PAD.n932 PAD.n928 0.0380882
R42368 PAD.n932 PAD.n859 0.0380882
R42369 PAD.n936 PAD.n859 0.0380882
R42370 PAD.n940 PAD.n936 0.0380882
R42371 PAD.n944 PAD.n940 0.0380882
R42372 PAD.n944 PAD.n857 0.0380882
R42373 PAD.n948 PAD.n857 0.0380882
R42374 PAD.n952 PAD.n948 0.0380882
R42375 PAD.n956 PAD.n952 0.0380882
R42376 PAD.n956 PAD.n855 0.0380882
R42377 PAD.n960 PAD.n855 0.0380882
R42378 PAD.n964 PAD.n960 0.0380882
R42379 PAD.n968 PAD.n964 0.0380882
R42380 PAD.n968 PAD.n853 0.0380882
R42381 PAD.n972 PAD.n853 0.0380882
R42382 PAD.n976 PAD.n972 0.0380882
R42383 PAD.n980 PAD.n976 0.0380882
R42384 PAD.n980 PAD.n851 0.0380882
R42385 PAD.n984 PAD.n851 0.0380882
R42386 PAD.n988 PAD.n984 0.0380882
R42387 PAD.n992 PAD.n988 0.0380882
R42388 PAD.n992 PAD.n849 0.0380882
R42389 PAD.n996 PAD.n849 0.0380882
R42390 PAD.n1000 PAD.n996 0.0380882
R42391 PAD.n1004 PAD.n1000 0.0380882
R42392 PAD.n1004 PAD.n847 0.0380882
R42393 PAD.n1008 PAD.n847 0.0380882
R42394 PAD.n1012 PAD.n1008 0.0380882
R42395 PAD.n1016 PAD.n1012 0.0380882
R42396 PAD.n1016 PAD.n845 0.0380882
R42397 PAD.n1020 PAD.n845 0.0380882
R42398 PAD.n1024 PAD.n1020 0.0380882
R42399 PAD.n1028 PAD.n1024 0.0380882
R42400 PAD.n1028 PAD.n843 0.0380882
R42401 PAD.n1032 PAD.n843 0.0380882
R42402 PAD.n1036 PAD.n1032 0.0380882
R42403 PAD.n1040 PAD.n1036 0.0380882
R42404 PAD.n1040 PAD.n841 0.0380882
R42405 PAD.n1044 PAD.n841 0.0380882
R42406 PAD.n1048 PAD.n1044 0.0380882
R42407 PAD.n1052 PAD.n1048 0.0380882
R42408 PAD.n1052 PAD.n839 0.0380882
R42409 PAD.n1056 PAD.n839 0.0380882
R42410 PAD.n1060 PAD.n1056 0.0380882
R42411 PAD.n1064 PAD.n1060 0.0380882
R42412 PAD.n1064 PAD.n837 0.0380882
R42413 PAD.n1068 PAD.n837 0.0380882
R42414 PAD.n1072 PAD.n1068 0.0380882
R42415 PAD.n1076 PAD.n1072 0.0380882
R42416 PAD.n1076 PAD.n835 0.0380882
R42417 PAD.n1080 PAD.n835 0.0380882
R42418 PAD.n1084 PAD.n1080 0.0380882
R42419 PAD.n1088 PAD.n1084 0.0380882
R42420 PAD.n1088 PAD.n833 0.0380882
R42421 PAD.n1092 PAD.n833 0.0380882
R42422 PAD.n1096 PAD.n1092 0.0380882
R42423 PAD.n1100 PAD.n1096 0.0380882
R42424 PAD.n1100 PAD.n831 0.0380882
R42425 PAD.n1104 PAD.n831 0.0380882
R42426 PAD.n1108 PAD.n1104 0.0380882
R42427 PAD.n1112 PAD.n1108 0.0380882
R42428 PAD.n1112 PAD.n829 0.0380882
R42429 PAD.n10384 PAD.n829 0.0380882
R42430 PAD.n10384 PAD.n826 0.0380882
R42431 PAD.n874 PAD.n873 0.0380882
R42432 PAD.n875 PAD.n874 0.0380882
R42433 PAD.n875 PAD.n868 0.0380882
R42434 PAD.n885 PAD.n868 0.0380882
R42435 PAD.n886 PAD.n885 0.0380882
R42436 PAD.n887 PAD.n886 0.0380882
R42437 PAD.n887 PAD.n866 0.0380882
R42438 PAD.n897 PAD.n866 0.0380882
R42439 PAD.n898 PAD.n897 0.0380882
R42440 PAD.n899 PAD.n898 0.0380882
R42441 PAD.n899 PAD.n864 0.0380882
R42442 PAD.n909 PAD.n864 0.0380882
R42443 PAD.n910 PAD.n909 0.0380882
R42444 PAD.n911 PAD.n910 0.0380882
R42445 PAD.n911 PAD.n862 0.0380882
R42446 PAD.n921 PAD.n862 0.0380882
R42447 PAD.n922 PAD.n921 0.0380882
R42448 PAD.n923 PAD.n922 0.0380882
R42449 PAD.n923 PAD.n860 0.0380882
R42450 PAD.n933 PAD.n860 0.0380882
R42451 PAD.n934 PAD.n933 0.0380882
R42452 PAD.n935 PAD.n934 0.0380882
R42453 PAD.n935 PAD.n858 0.0380882
R42454 PAD.n945 PAD.n858 0.0380882
R42455 PAD.n946 PAD.n945 0.0380882
R42456 PAD.n947 PAD.n946 0.0380882
R42457 PAD.n947 PAD.n856 0.0380882
R42458 PAD.n957 PAD.n856 0.0380882
R42459 PAD.n958 PAD.n957 0.0380882
R42460 PAD.n959 PAD.n958 0.0380882
R42461 PAD.n959 PAD.n854 0.0380882
R42462 PAD.n969 PAD.n854 0.0380882
R42463 PAD.n970 PAD.n969 0.0380882
R42464 PAD.n971 PAD.n970 0.0380882
R42465 PAD.n971 PAD.n852 0.0380882
R42466 PAD.n981 PAD.n852 0.0380882
R42467 PAD.n982 PAD.n981 0.0380882
R42468 PAD.n983 PAD.n982 0.0380882
R42469 PAD.n983 PAD.n850 0.0380882
R42470 PAD.n993 PAD.n850 0.0380882
R42471 PAD.n994 PAD.n993 0.0380882
R42472 PAD.n995 PAD.n994 0.0380882
R42473 PAD.n995 PAD.n848 0.0380882
R42474 PAD.n1005 PAD.n848 0.0380882
R42475 PAD.n1006 PAD.n1005 0.0380882
R42476 PAD.n1007 PAD.n1006 0.0380882
R42477 PAD.n1007 PAD.n846 0.0380882
R42478 PAD.n1017 PAD.n846 0.0380882
R42479 PAD.n1018 PAD.n1017 0.0380882
R42480 PAD.n1019 PAD.n1018 0.0380882
R42481 PAD.n1019 PAD.n844 0.0380882
R42482 PAD.n1029 PAD.n844 0.0380882
R42483 PAD.n1030 PAD.n1029 0.0380882
R42484 PAD.n1031 PAD.n1030 0.0380882
R42485 PAD.n1031 PAD.n842 0.0380882
R42486 PAD.n1041 PAD.n842 0.0380882
R42487 PAD.n1042 PAD.n1041 0.0380882
R42488 PAD.n1043 PAD.n1042 0.0380882
R42489 PAD.n1043 PAD.n840 0.0380882
R42490 PAD.n1053 PAD.n840 0.0380882
R42491 PAD.n1054 PAD.n1053 0.0380882
R42492 PAD.n1055 PAD.n1054 0.0380882
R42493 PAD.n1055 PAD.n838 0.0380882
R42494 PAD.n1065 PAD.n838 0.0380882
R42495 PAD.n1066 PAD.n1065 0.0380882
R42496 PAD.n1067 PAD.n1066 0.0380882
R42497 PAD.n1067 PAD.n836 0.0380882
R42498 PAD.n1077 PAD.n836 0.0380882
R42499 PAD.n1078 PAD.n1077 0.0380882
R42500 PAD.n1079 PAD.n1078 0.0380882
R42501 PAD.n1079 PAD.n834 0.0380882
R42502 PAD.n1089 PAD.n834 0.0380882
R42503 PAD.n1090 PAD.n1089 0.0380882
R42504 PAD.n1091 PAD.n1090 0.0380882
R42505 PAD.n1091 PAD.n832 0.0380882
R42506 PAD.n1101 PAD.n832 0.0380882
R42507 PAD.n1102 PAD.n1101 0.0380882
R42508 PAD.n1103 PAD.n1102 0.0380882
R42509 PAD.n1103 PAD.n830 0.0380882
R42510 PAD.n1113 PAD.n830 0.0380882
R42511 PAD.n1114 PAD.n1113 0.0380882
R42512 PAD.n10383 PAD.n1114 0.0380882
R42513 PAD.n10383 PAD.n10382 0.0380882
R42514 PAD.n10105 PAD.n10104 0.0380882
R42515 PAD.n10113 PAD.n10104 0.0380882
R42516 PAD.n10113 PAD.n10102 0.0380882
R42517 PAD.n10117 PAD.n10102 0.0380882
R42518 PAD.n10117 PAD.n10100 0.0380882
R42519 PAD.n10125 PAD.n10100 0.0380882
R42520 PAD.n10125 PAD.n10098 0.0380882
R42521 PAD.n10129 PAD.n10098 0.0380882
R42522 PAD.n10129 PAD.n10096 0.0380882
R42523 PAD.n10137 PAD.n10096 0.0380882
R42524 PAD.n10137 PAD.n10094 0.0380882
R42525 PAD.n10141 PAD.n10094 0.0380882
R42526 PAD.n10141 PAD.n10092 0.0380882
R42527 PAD.n10149 PAD.n10092 0.0380882
R42528 PAD.n10149 PAD.n10090 0.0380882
R42529 PAD.n10153 PAD.n10090 0.0380882
R42530 PAD.n10153 PAD.n10088 0.0380882
R42531 PAD.n10161 PAD.n10088 0.0380882
R42532 PAD.n10161 PAD.n10086 0.0380882
R42533 PAD.n10165 PAD.n10086 0.0380882
R42534 PAD.n10165 PAD.n10084 0.0380882
R42535 PAD.n10173 PAD.n10084 0.0380882
R42536 PAD.n10173 PAD.n10082 0.0380882
R42537 PAD.n10177 PAD.n10082 0.0380882
R42538 PAD.n10177 PAD.n10080 0.0380882
R42539 PAD.n10185 PAD.n10080 0.0380882
R42540 PAD.n10185 PAD.n10078 0.0380882
R42541 PAD.n10189 PAD.n10078 0.0380882
R42542 PAD.n10189 PAD.n10076 0.0380882
R42543 PAD.n10197 PAD.n10076 0.0380882
R42544 PAD.n10197 PAD.n10074 0.0380882
R42545 PAD.n10201 PAD.n10074 0.0380882
R42546 PAD.n10201 PAD.n10072 0.0380882
R42547 PAD.n10209 PAD.n10072 0.0380882
R42548 PAD.n10209 PAD.n10070 0.0380882
R42549 PAD.n10213 PAD.n10070 0.0380882
R42550 PAD.n10213 PAD.n10068 0.0380882
R42551 PAD.n10221 PAD.n10068 0.0380882
R42552 PAD.n10221 PAD.n10066 0.0380882
R42553 PAD.n10225 PAD.n10066 0.0380882
R42554 PAD.n10225 PAD.n10064 0.0380882
R42555 PAD.n10233 PAD.n10064 0.0380882
R42556 PAD.n10233 PAD.n10062 0.0380882
R42557 PAD.n10237 PAD.n10062 0.0380882
R42558 PAD.n10237 PAD.n10060 0.0380882
R42559 PAD.n10245 PAD.n10060 0.0380882
R42560 PAD.n10245 PAD.n10058 0.0380882
R42561 PAD.n10249 PAD.n10058 0.0380882
R42562 PAD.n10249 PAD.n10056 0.0380882
R42563 PAD.n10257 PAD.n10056 0.0380882
R42564 PAD.n10257 PAD.n10054 0.0380882
R42565 PAD.n10261 PAD.n10054 0.0380882
R42566 PAD.n10261 PAD.n10052 0.0380882
R42567 PAD.n10269 PAD.n10052 0.0380882
R42568 PAD.n10269 PAD.n10050 0.0380882
R42569 PAD.n10273 PAD.n10050 0.0380882
R42570 PAD.n10273 PAD.n10048 0.0380882
R42571 PAD.n10281 PAD.n10048 0.0380882
R42572 PAD.n10281 PAD.n10046 0.0380882
R42573 PAD.n10285 PAD.n10046 0.0380882
R42574 PAD.n10285 PAD.n10044 0.0380882
R42575 PAD.n10293 PAD.n10044 0.0380882
R42576 PAD.n10293 PAD.n10042 0.0380882
R42577 PAD.n10297 PAD.n10042 0.0380882
R42578 PAD.n10297 PAD.n10040 0.0380882
R42579 PAD.n10305 PAD.n10040 0.0380882
R42580 PAD.n10305 PAD.n10038 0.0380882
R42581 PAD.n10309 PAD.n10038 0.0380882
R42582 PAD.n10309 PAD.n10036 0.0380882
R42583 PAD.n10317 PAD.n10036 0.0380882
R42584 PAD.n10317 PAD.n10034 0.0380882
R42585 PAD.n10321 PAD.n10034 0.0380882
R42586 PAD.n10321 PAD.n10032 0.0380882
R42587 PAD.n10329 PAD.n10032 0.0380882
R42588 PAD.n10329 PAD.n10030 0.0380882
R42589 PAD.n10333 PAD.n10030 0.0380882
R42590 PAD.n10333 PAD.n10028 0.0380882
R42591 PAD.n10341 PAD.n10028 0.0380882
R42592 PAD.n10341 PAD.n10026 0.0380882
R42593 PAD.n10346 PAD.n10026 0.0380882
R42594 PAD.n10346 PAD.n10024 0.0380882
R42595 PAD.n10024 PAD.n10023 0.0380882
R42596 PAD.n10354 PAD.n10023 0.0380882
R42597 PAD.n10103 PAD.n1124 0.0380882
R42598 PAD.n10114 PAD.n10103 0.0380882
R42599 PAD.n10115 PAD.n10114 0.0380882
R42600 PAD.n10116 PAD.n10115 0.0380882
R42601 PAD.n10116 PAD.n10099 0.0380882
R42602 PAD.n10126 PAD.n10099 0.0380882
R42603 PAD.n10127 PAD.n10126 0.0380882
R42604 PAD.n10128 PAD.n10127 0.0380882
R42605 PAD.n10128 PAD.n10095 0.0380882
R42606 PAD.n10138 PAD.n10095 0.0380882
R42607 PAD.n10139 PAD.n10138 0.0380882
R42608 PAD.n10140 PAD.n10139 0.0380882
R42609 PAD.n10140 PAD.n10091 0.0380882
R42610 PAD.n10150 PAD.n10091 0.0380882
R42611 PAD.n10151 PAD.n10150 0.0380882
R42612 PAD.n10152 PAD.n10151 0.0380882
R42613 PAD.n10152 PAD.n10087 0.0380882
R42614 PAD.n10162 PAD.n10087 0.0380882
R42615 PAD.n10163 PAD.n10162 0.0380882
R42616 PAD.n10164 PAD.n10163 0.0380882
R42617 PAD.n10164 PAD.n10083 0.0380882
R42618 PAD.n10174 PAD.n10083 0.0380882
R42619 PAD.n10175 PAD.n10174 0.0380882
R42620 PAD.n10176 PAD.n10175 0.0380882
R42621 PAD.n10176 PAD.n10079 0.0380882
R42622 PAD.n10186 PAD.n10079 0.0380882
R42623 PAD.n10187 PAD.n10186 0.0380882
R42624 PAD.n10188 PAD.n10187 0.0380882
R42625 PAD.n10188 PAD.n10075 0.0380882
R42626 PAD.n10198 PAD.n10075 0.0380882
R42627 PAD.n10199 PAD.n10198 0.0380882
R42628 PAD.n10200 PAD.n10199 0.0380882
R42629 PAD.n10200 PAD.n10071 0.0380882
R42630 PAD.n10210 PAD.n10071 0.0380882
R42631 PAD.n10211 PAD.n10210 0.0380882
R42632 PAD.n10212 PAD.n10211 0.0380882
R42633 PAD.n10212 PAD.n10067 0.0380882
R42634 PAD.n10222 PAD.n10067 0.0380882
R42635 PAD.n10223 PAD.n10222 0.0380882
R42636 PAD.n10224 PAD.n10223 0.0380882
R42637 PAD.n10224 PAD.n10063 0.0380882
R42638 PAD.n10234 PAD.n10063 0.0380882
R42639 PAD.n10235 PAD.n10234 0.0380882
R42640 PAD.n10236 PAD.n10235 0.0380882
R42641 PAD.n10236 PAD.n10059 0.0380882
R42642 PAD.n10246 PAD.n10059 0.0380882
R42643 PAD.n10247 PAD.n10246 0.0380882
R42644 PAD.n10248 PAD.n10247 0.0380882
R42645 PAD.n10248 PAD.n10055 0.0380882
R42646 PAD.n10258 PAD.n10055 0.0380882
R42647 PAD.n10259 PAD.n10258 0.0380882
R42648 PAD.n10260 PAD.n10259 0.0380882
R42649 PAD.n10260 PAD.n10051 0.0380882
R42650 PAD.n10270 PAD.n10051 0.0380882
R42651 PAD.n10271 PAD.n10270 0.0380882
R42652 PAD.n10272 PAD.n10271 0.0380882
R42653 PAD.n10272 PAD.n10047 0.0380882
R42654 PAD.n10282 PAD.n10047 0.0380882
R42655 PAD.n10283 PAD.n10282 0.0380882
R42656 PAD.n10284 PAD.n10283 0.0380882
R42657 PAD.n10284 PAD.n10043 0.0380882
R42658 PAD.n10294 PAD.n10043 0.0380882
R42659 PAD.n10295 PAD.n10294 0.0380882
R42660 PAD.n10296 PAD.n10295 0.0380882
R42661 PAD.n10296 PAD.n10039 0.0380882
R42662 PAD.n10306 PAD.n10039 0.0380882
R42663 PAD.n10307 PAD.n10306 0.0380882
R42664 PAD.n10308 PAD.n10307 0.0380882
R42665 PAD.n10308 PAD.n10035 0.0380882
R42666 PAD.n10318 PAD.n10035 0.0380882
R42667 PAD.n10319 PAD.n10318 0.0380882
R42668 PAD.n10320 PAD.n10319 0.0380882
R42669 PAD.n10320 PAD.n10031 0.0380882
R42670 PAD.n10330 PAD.n10031 0.0380882
R42671 PAD.n10331 PAD.n10330 0.0380882
R42672 PAD.n10332 PAD.n10331 0.0380882
R42673 PAD.n10332 PAD.n10027 0.0380882
R42674 PAD.n10342 PAD.n10027 0.0380882
R42675 PAD.n10343 PAD.n10342 0.0380882
R42676 PAD.n10345 PAD.n10343 0.0380882
R42677 PAD.n10345 PAD.n10344 0.0380882
R42678 PAD.n10344 PAD.n10022 0.0380882
R42679 PAD.n10355 PAD.n10022 0.0380882
R42680 PAD.n1480 PAD.n1479 0.0380882
R42681 PAD.n1479 PAD.n1193 0.0380882
R42682 PAD.n1475 PAD.n1193 0.0380882
R42683 PAD.n1475 PAD.n1471 0.0380882
R42684 PAD.n1471 PAD.n1470 0.0380882
R42685 PAD.n1470 PAD.n1195 0.0380882
R42686 PAD.n1466 PAD.n1195 0.0380882
R42687 PAD.n1466 PAD.n1462 0.0380882
R42688 PAD.n1462 PAD.n1461 0.0380882
R42689 PAD.n1461 PAD.n1200 0.0380882
R42690 PAD.n1457 PAD.n1200 0.0380882
R42691 PAD.n1457 PAD.n1453 0.0380882
R42692 PAD.n1453 PAD.n1452 0.0380882
R42693 PAD.n1452 PAD.n1205 0.0380882
R42694 PAD.n1448 PAD.n1205 0.0380882
R42695 PAD.n1448 PAD.n1444 0.0380882
R42696 PAD.n1444 PAD.n1443 0.0380882
R42697 PAD.n1443 PAD.n1210 0.0380882
R42698 PAD.n1439 PAD.n1210 0.0380882
R42699 PAD.n1439 PAD.n1435 0.0380882
R42700 PAD.n1435 PAD.n1434 0.0380882
R42701 PAD.n1434 PAD.n1215 0.0380882
R42702 PAD.n1430 PAD.n1215 0.0380882
R42703 PAD.n1430 PAD.n1426 0.0380882
R42704 PAD.n1426 PAD.n1425 0.0380882
R42705 PAD.n1425 PAD.n1220 0.0380882
R42706 PAD.n1421 PAD.n1220 0.0380882
R42707 PAD.n1421 PAD.n1417 0.0380882
R42708 PAD.n1417 PAD.n1416 0.0380882
R42709 PAD.n1416 PAD.n1225 0.0380882
R42710 PAD.n1412 PAD.n1225 0.0380882
R42711 PAD.n1412 PAD.n1408 0.0380882
R42712 PAD.n1408 PAD.n1407 0.0380882
R42713 PAD.n1407 PAD.n1230 0.0380882
R42714 PAD.n1403 PAD.n1230 0.0380882
R42715 PAD.n1403 PAD.n1399 0.0380882
R42716 PAD.n1399 PAD.n1398 0.0380882
R42717 PAD.n1398 PAD.n1235 0.0380882
R42718 PAD.n1394 PAD.n1235 0.0380882
R42719 PAD.n1394 PAD.n1390 0.0380882
R42720 PAD.n1390 PAD.n1389 0.0380882
R42721 PAD.n1389 PAD.n1240 0.0380882
R42722 PAD.n1385 PAD.n1240 0.0380882
R42723 PAD.n1385 PAD.n1381 0.0380882
R42724 PAD.n1381 PAD.n1380 0.0380882
R42725 PAD.n1380 PAD.n1245 0.0380882
R42726 PAD.n1376 PAD.n1245 0.0380882
R42727 PAD.n1376 PAD.n1372 0.0380882
R42728 PAD.n1372 PAD.n1371 0.0380882
R42729 PAD.n1371 PAD.n1250 0.0380882
R42730 PAD.n1367 PAD.n1250 0.0380882
R42731 PAD.n1367 PAD.n1363 0.0380882
R42732 PAD.n1363 PAD.n1362 0.0380882
R42733 PAD.n1362 PAD.n1255 0.0380882
R42734 PAD.n1358 PAD.n1255 0.0380882
R42735 PAD.n1358 PAD.n1354 0.0380882
R42736 PAD.n1354 PAD.n1353 0.0380882
R42737 PAD.n1353 PAD.n1260 0.0380882
R42738 PAD.n1349 PAD.n1260 0.0380882
R42739 PAD.n1349 PAD.n1345 0.0380882
R42740 PAD.n1345 PAD.n1344 0.0380882
R42741 PAD.n1344 PAD.n1265 0.0380882
R42742 PAD.n1340 PAD.n1265 0.0380882
R42743 PAD.n1340 PAD.n1336 0.0380882
R42744 PAD.n1336 PAD.n1335 0.0380882
R42745 PAD.n1335 PAD.n1270 0.0380882
R42746 PAD.n1331 PAD.n1270 0.0380882
R42747 PAD.n1331 PAD.n1327 0.0380882
R42748 PAD.n1327 PAD.n1326 0.0380882
R42749 PAD.n1326 PAD.n1275 0.0380882
R42750 PAD.n1322 PAD.n1275 0.0380882
R42751 PAD.n1322 PAD.n1318 0.0380882
R42752 PAD.n1318 PAD.n1317 0.0380882
R42753 PAD.n1317 PAD.n1280 0.0380882
R42754 PAD.n1313 PAD.n1280 0.0380882
R42755 PAD.n1313 PAD.n1309 0.0380882
R42756 PAD.n1309 PAD.n1308 0.0380882
R42757 PAD.n1308 PAD.n1285 0.0380882
R42758 PAD.n1304 PAD.n1285 0.0380882
R42759 PAD.n1304 PAD.n1300 0.0380882
R42760 PAD.n1300 PAD.n1299 0.0380882
R42761 PAD.n1299 PAD.n1290 0.0380882
R42762 PAD.n1295 PAD.n1290 0.0380882
R42763 PAD.n1478 PAD.n1145 0.0380882
R42764 PAD.n1478 PAD.n1477 0.0380882
R42765 PAD.n1477 PAD.n1476 0.0380882
R42766 PAD.n1476 PAD.n1194 0.0380882
R42767 PAD.n1469 PAD.n1194 0.0380882
R42768 PAD.n1469 PAD.n1468 0.0380882
R42769 PAD.n1468 PAD.n1467 0.0380882
R42770 PAD.n1467 PAD.n1199 0.0380882
R42771 PAD.n1460 PAD.n1199 0.0380882
R42772 PAD.n1460 PAD.n1459 0.0380882
R42773 PAD.n1459 PAD.n1458 0.0380882
R42774 PAD.n1458 PAD.n1204 0.0380882
R42775 PAD.n1451 PAD.n1204 0.0380882
R42776 PAD.n1451 PAD.n1450 0.0380882
R42777 PAD.n1450 PAD.n1449 0.0380882
R42778 PAD.n1449 PAD.n1209 0.0380882
R42779 PAD.n1442 PAD.n1209 0.0380882
R42780 PAD.n1442 PAD.n1441 0.0380882
R42781 PAD.n1441 PAD.n1440 0.0380882
R42782 PAD.n1440 PAD.n1214 0.0380882
R42783 PAD.n1433 PAD.n1214 0.0380882
R42784 PAD.n1433 PAD.n1432 0.0380882
R42785 PAD.n1432 PAD.n1431 0.0380882
R42786 PAD.n1431 PAD.n1219 0.0380882
R42787 PAD.n1424 PAD.n1219 0.0380882
R42788 PAD.n1424 PAD.n1423 0.0380882
R42789 PAD.n1423 PAD.n1422 0.0380882
R42790 PAD.n1422 PAD.n1224 0.0380882
R42791 PAD.n1415 PAD.n1224 0.0380882
R42792 PAD.n1415 PAD.n1414 0.0380882
R42793 PAD.n1414 PAD.n1413 0.0380882
R42794 PAD.n1413 PAD.n1229 0.0380882
R42795 PAD.n1406 PAD.n1229 0.0380882
R42796 PAD.n1406 PAD.n1405 0.0380882
R42797 PAD.n1405 PAD.n1404 0.0380882
R42798 PAD.n1404 PAD.n1234 0.0380882
R42799 PAD.n1397 PAD.n1234 0.0380882
R42800 PAD.n1397 PAD.n1396 0.0380882
R42801 PAD.n1396 PAD.n1395 0.0380882
R42802 PAD.n1395 PAD.n1239 0.0380882
R42803 PAD.n1388 PAD.n1239 0.0380882
R42804 PAD.n1388 PAD.n1387 0.0380882
R42805 PAD.n1387 PAD.n1386 0.0380882
R42806 PAD.n1386 PAD.n1244 0.0380882
R42807 PAD.n1379 PAD.n1244 0.0380882
R42808 PAD.n1379 PAD.n1378 0.0380882
R42809 PAD.n1378 PAD.n1377 0.0380882
R42810 PAD.n1377 PAD.n1249 0.0380882
R42811 PAD.n1370 PAD.n1249 0.0380882
R42812 PAD.n1370 PAD.n1369 0.0380882
R42813 PAD.n1369 PAD.n1368 0.0380882
R42814 PAD.n1368 PAD.n1254 0.0380882
R42815 PAD.n1361 PAD.n1254 0.0380882
R42816 PAD.n1361 PAD.n1360 0.0380882
R42817 PAD.n1360 PAD.n1359 0.0380882
R42818 PAD.n1359 PAD.n1259 0.0380882
R42819 PAD.n1352 PAD.n1259 0.0380882
R42820 PAD.n1352 PAD.n1351 0.0380882
R42821 PAD.n1351 PAD.n1350 0.0380882
R42822 PAD.n1350 PAD.n1264 0.0380882
R42823 PAD.n1343 PAD.n1264 0.0380882
R42824 PAD.n1343 PAD.n1342 0.0380882
R42825 PAD.n1342 PAD.n1341 0.0380882
R42826 PAD.n1341 PAD.n1269 0.0380882
R42827 PAD.n1334 PAD.n1269 0.0380882
R42828 PAD.n1334 PAD.n1333 0.0380882
R42829 PAD.n1333 PAD.n1332 0.0380882
R42830 PAD.n1332 PAD.n1274 0.0380882
R42831 PAD.n1325 PAD.n1274 0.0380882
R42832 PAD.n1325 PAD.n1324 0.0380882
R42833 PAD.n1324 PAD.n1323 0.0380882
R42834 PAD.n1323 PAD.n1279 0.0380882
R42835 PAD.n1316 PAD.n1279 0.0380882
R42836 PAD.n1316 PAD.n1315 0.0380882
R42837 PAD.n1315 PAD.n1314 0.0380882
R42838 PAD.n1314 PAD.n1284 0.0380882
R42839 PAD.n1307 PAD.n1284 0.0380882
R42840 PAD.n1307 PAD.n1306 0.0380882
R42841 PAD.n1306 PAD.n1305 0.0380882
R42842 PAD.n1305 PAD.n1289 0.0380882
R42843 PAD.n1298 PAD.n1289 0.0380882
R42844 PAD.n1298 PAD.n1297 0.0380882
R42845 PAD.n1297 PAD.n1296 0.0380882
R42846 PAD.n9749 PAD.n1579 0.0380882
R42847 PAD.n9753 PAD.n1579 0.0380882
R42848 PAD.n9757 PAD.n9753 0.0380882
R42849 PAD.n9761 PAD.n9757 0.0380882
R42850 PAD.n9761 PAD.n1575 0.0380882
R42851 PAD.n9765 PAD.n1575 0.0380882
R42852 PAD.n9769 PAD.n9765 0.0380882
R42853 PAD.n9773 PAD.n9769 0.0380882
R42854 PAD.n9773 PAD.n1573 0.0380882
R42855 PAD.n9777 PAD.n1573 0.0380882
R42856 PAD.n9781 PAD.n9777 0.0380882
R42857 PAD.n9785 PAD.n9781 0.0380882
R42858 PAD.n9785 PAD.n1571 0.0380882
R42859 PAD.n9789 PAD.n1571 0.0380882
R42860 PAD.n9793 PAD.n9789 0.0380882
R42861 PAD.n9797 PAD.n9793 0.0380882
R42862 PAD.n9797 PAD.n1569 0.0380882
R42863 PAD.n9801 PAD.n1569 0.0380882
R42864 PAD.n9805 PAD.n9801 0.0380882
R42865 PAD.n9809 PAD.n9805 0.0380882
R42866 PAD.n9809 PAD.n1567 0.0380882
R42867 PAD.n9813 PAD.n1567 0.0380882
R42868 PAD.n9817 PAD.n9813 0.0380882
R42869 PAD.n9821 PAD.n9817 0.0380882
R42870 PAD.n9821 PAD.n1565 0.0380882
R42871 PAD.n9825 PAD.n1565 0.0380882
R42872 PAD.n9829 PAD.n9825 0.0380882
R42873 PAD.n9833 PAD.n9829 0.0380882
R42874 PAD.n9833 PAD.n1563 0.0380882
R42875 PAD.n9837 PAD.n1563 0.0380882
R42876 PAD.n9841 PAD.n9837 0.0380882
R42877 PAD.n9845 PAD.n9841 0.0380882
R42878 PAD.n9845 PAD.n1561 0.0380882
R42879 PAD.n9849 PAD.n1561 0.0380882
R42880 PAD.n9853 PAD.n9849 0.0380882
R42881 PAD.n9857 PAD.n9853 0.0380882
R42882 PAD.n9857 PAD.n1559 0.0380882
R42883 PAD.n9861 PAD.n1559 0.0380882
R42884 PAD.n9865 PAD.n9861 0.0380882
R42885 PAD.n9869 PAD.n9865 0.0380882
R42886 PAD.n9869 PAD.n1557 0.0380882
R42887 PAD.n9873 PAD.n1557 0.0380882
R42888 PAD.n9877 PAD.n9873 0.0380882
R42889 PAD.n9881 PAD.n9877 0.0380882
R42890 PAD.n9881 PAD.n1555 0.0380882
R42891 PAD.n9885 PAD.n1555 0.0380882
R42892 PAD.n9889 PAD.n9885 0.0380882
R42893 PAD.n9893 PAD.n9889 0.0380882
R42894 PAD.n9893 PAD.n1553 0.0380882
R42895 PAD.n9897 PAD.n1553 0.0380882
R42896 PAD.n9901 PAD.n9897 0.0380882
R42897 PAD.n9905 PAD.n9901 0.0380882
R42898 PAD.n9905 PAD.n1551 0.0380882
R42899 PAD.n9909 PAD.n1551 0.0380882
R42900 PAD.n9913 PAD.n9909 0.0380882
R42901 PAD.n9917 PAD.n9913 0.0380882
R42902 PAD.n9917 PAD.n1549 0.0380882
R42903 PAD.n9921 PAD.n1549 0.0380882
R42904 PAD.n9925 PAD.n9921 0.0380882
R42905 PAD.n9929 PAD.n9925 0.0380882
R42906 PAD.n9929 PAD.n1547 0.0380882
R42907 PAD.n9933 PAD.n1547 0.0380882
R42908 PAD.n9937 PAD.n9933 0.0380882
R42909 PAD.n9941 PAD.n9937 0.0380882
R42910 PAD.n9941 PAD.n1545 0.0380882
R42911 PAD.n9945 PAD.n1545 0.0380882
R42912 PAD.n9949 PAD.n9945 0.0380882
R42913 PAD.n9953 PAD.n9949 0.0380882
R42914 PAD.n9953 PAD.n1543 0.0380882
R42915 PAD.n9957 PAD.n1543 0.0380882
R42916 PAD.n9961 PAD.n9957 0.0380882
R42917 PAD.n9965 PAD.n9961 0.0380882
R42918 PAD.n9965 PAD.n1541 0.0380882
R42919 PAD.n9969 PAD.n1541 0.0380882
R42920 PAD.n9973 PAD.n9969 0.0380882
R42921 PAD.n9977 PAD.n9973 0.0380882
R42922 PAD.n9977 PAD.n1539 0.0380882
R42923 PAD.n9981 PAD.n1539 0.0380882
R42924 PAD.n9985 PAD.n9981 0.0380882
R42925 PAD.n9989 PAD.n9985 0.0380882
R42926 PAD.n9989 PAD.n1537 0.0380882
R42927 PAD.n9994 PAD.n1537 0.0380882
R42928 PAD.n9994 PAD.n1535 0.0380882
R42929 PAD.n9751 PAD.n9750 0.0380882
R42930 PAD.n9752 PAD.n9751 0.0380882
R42931 PAD.n9752 PAD.n1576 0.0380882
R42932 PAD.n9762 PAD.n1576 0.0380882
R42933 PAD.n9763 PAD.n9762 0.0380882
R42934 PAD.n9764 PAD.n9763 0.0380882
R42935 PAD.n9764 PAD.n1574 0.0380882
R42936 PAD.n9774 PAD.n1574 0.0380882
R42937 PAD.n9775 PAD.n9774 0.0380882
R42938 PAD.n9776 PAD.n9775 0.0380882
R42939 PAD.n9776 PAD.n1572 0.0380882
R42940 PAD.n9786 PAD.n1572 0.0380882
R42941 PAD.n9787 PAD.n9786 0.0380882
R42942 PAD.n9788 PAD.n9787 0.0380882
R42943 PAD.n9788 PAD.n1570 0.0380882
R42944 PAD.n9798 PAD.n1570 0.0380882
R42945 PAD.n9799 PAD.n9798 0.0380882
R42946 PAD.n9800 PAD.n9799 0.0380882
R42947 PAD.n9800 PAD.n1568 0.0380882
R42948 PAD.n9810 PAD.n1568 0.0380882
R42949 PAD.n9811 PAD.n9810 0.0380882
R42950 PAD.n9812 PAD.n9811 0.0380882
R42951 PAD.n9812 PAD.n1566 0.0380882
R42952 PAD.n9822 PAD.n1566 0.0380882
R42953 PAD.n9823 PAD.n9822 0.0380882
R42954 PAD.n9824 PAD.n9823 0.0380882
R42955 PAD.n9824 PAD.n1564 0.0380882
R42956 PAD.n9834 PAD.n1564 0.0380882
R42957 PAD.n9835 PAD.n9834 0.0380882
R42958 PAD.n9836 PAD.n9835 0.0380882
R42959 PAD.n9836 PAD.n1562 0.0380882
R42960 PAD.n9846 PAD.n1562 0.0380882
R42961 PAD.n9847 PAD.n9846 0.0380882
R42962 PAD.n9848 PAD.n9847 0.0380882
R42963 PAD.n9848 PAD.n1560 0.0380882
R42964 PAD.n9858 PAD.n1560 0.0380882
R42965 PAD.n9859 PAD.n9858 0.0380882
R42966 PAD.n9860 PAD.n9859 0.0380882
R42967 PAD.n9860 PAD.n1558 0.0380882
R42968 PAD.n9870 PAD.n1558 0.0380882
R42969 PAD.n9871 PAD.n9870 0.0380882
R42970 PAD.n9872 PAD.n9871 0.0380882
R42971 PAD.n9872 PAD.n1556 0.0380882
R42972 PAD.n9882 PAD.n1556 0.0380882
R42973 PAD.n9883 PAD.n9882 0.0380882
R42974 PAD.n9884 PAD.n9883 0.0380882
R42975 PAD.n9884 PAD.n1554 0.0380882
R42976 PAD.n9894 PAD.n1554 0.0380882
R42977 PAD.n9895 PAD.n9894 0.0380882
R42978 PAD.n9896 PAD.n9895 0.0380882
R42979 PAD.n9896 PAD.n1552 0.0380882
R42980 PAD.n9906 PAD.n1552 0.0380882
R42981 PAD.n9907 PAD.n9906 0.0380882
R42982 PAD.n9908 PAD.n9907 0.0380882
R42983 PAD.n9908 PAD.n1550 0.0380882
R42984 PAD.n9918 PAD.n1550 0.0380882
R42985 PAD.n9919 PAD.n9918 0.0380882
R42986 PAD.n9920 PAD.n9919 0.0380882
R42987 PAD.n9920 PAD.n1548 0.0380882
R42988 PAD.n9930 PAD.n1548 0.0380882
R42989 PAD.n9931 PAD.n9930 0.0380882
R42990 PAD.n9932 PAD.n9931 0.0380882
R42991 PAD.n9932 PAD.n1546 0.0380882
R42992 PAD.n9942 PAD.n1546 0.0380882
R42993 PAD.n9943 PAD.n9942 0.0380882
R42994 PAD.n9944 PAD.n9943 0.0380882
R42995 PAD.n9944 PAD.n1544 0.0380882
R42996 PAD.n9954 PAD.n1544 0.0380882
R42997 PAD.n9955 PAD.n9954 0.0380882
R42998 PAD.n9956 PAD.n9955 0.0380882
R42999 PAD.n9956 PAD.n1542 0.0380882
R43000 PAD.n9966 PAD.n1542 0.0380882
R43001 PAD.n9967 PAD.n9966 0.0380882
R43002 PAD.n9968 PAD.n9967 0.0380882
R43003 PAD.n9968 PAD.n1540 0.0380882
R43004 PAD.n9978 PAD.n1540 0.0380882
R43005 PAD.n9979 PAD.n9978 0.0380882
R43006 PAD.n9980 PAD.n9979 0.0380882
R43007 PAD.n9980 PAD.n1538 0.0380882
R43008 PAD.n9990 PAD.n1538 0.0380882
R43009 PAD.n9991 PAD.n9990 0.0380882
R43010 PAD.n9993 PAD.n9991 0.0380882
R43011 PAD.n9993 PAD.n9992 0.0380882
R43012 PAD.n1931 PAD.n1930 0.0380882
R43013 PAD.n1930 PAD.n1600 0.0380882
R43014 PAD.n1924 PAD.n1600 0.0380882
R43015 PAD.n1924 PAD.n1603 0.0380882
R43016 PAD.n1920 PAD.n1603 0.0380882
R43017 PAD.n1920 PAD.n1606 0.0380882
R43018 PAD.n1912 PAD.n1606 0.0380882
R43019 PAD.n1912 PAD.n1608 0.0380882
R43020 PAD.n1908 PAD.n1608 0.0380882
R43021 PAD.n1908 PAD.n1610 0.0380882
R43022 PAD.n1900 PAD.n1610 0.0380882
R43023 PAD.n1900 PAD.n1612 0.0380882
R43024 PAD.n1896 PAD.n1612 0.0380882
R43025 PAD.n1896 PAD.n1614 0.0380882
R43026 PAD.n1888 PAD.n1614 0.0380882
R43027 PAD.n1888 PAD.n1616 0.0380882
R43028 PAD.n1884 PAD.n1616 0.0380882
R43029 PAD.n1884 PAD.n1618 0.0380882
R43030 PAD.n1876 PAD.n1618 0.0380882
R43031 PAD.n1876 PAD.n1620 0.0380882
R43032 PAD.n1872 PAD.n1620 0.0380882
R43033 PAD.n1872 PAD.n1622 0.0380882
R43034 PAD.n1864 PAD.n1622 0.0380882
R43035 PAD.n1864 PAD.n1624 0.0380882
R43036 PAD.n1860 PAD.n1624 0.0380882
R43037 PAD.n1860 PAD.n1626 0.0380882
R43038 PAD.n1852 PAD.n1626 0.0380882
R43039 PAD.n1852 PAD.n1628 0.0380882
R43040 PAD.n1848 PAD.n1628 0.0380882
R43041 PAD.n1848 PAD.n1630 0.0380882
R43042 PAD.n1840 PAD.n1630 0.0380882
R43043 PAD.n1840 PAD.n1632 0.0380882
R43044 PAD.n1836 PAD.n1632 0.0380882
R43045 PAD.n1836 PAD.n1634 0.0380882
R43046 PAD.n1828 PAD.n1634 0.0380882
R43047 PAD.n1828 PAD.n1636 0.0380882
R43048 PAD.n1824 PAD.n1636 0.0380882
R43049 PAD.n1824 PAD.n1638 0.0380882
R43050 PAD.n1816 PAD.n1638 0.0380882
R43051 PAD.n1816 PAD.n1640 0.0380882
R43052 PAD.n1812 PAD.n1640 0.0380882
R43053 PAD.n1812 PAD.n1642 0.0380882
R43054 PAD.n1804 PAD.n1642 0.0380882
R43055 PAD.n1804 PAD.n1644 0.0380882
R43056 PAD.n1800 PAD.n1644 0.0380882
R43057 PAD.n1800 PAD.n1646 0.0380882
R43058 PAD.n1792 PAD.n1646 0.0380882
R43059 PAD.n1792 PAD.n1648 0.0380882
R43060 PAD.n1788 PAD.n1648 0.0380882
R43061 PAD.n1788 PAD.n1650 0.0380882
R43062 PAD.n1780 PAD.n1650 0.0380882
R43063 PAD.n1780 PAD.n1652 0.0380882
R43064 PAD.n1776 PAD.n1652 0.0380882
R43065 PAD.n1776 PAD.n1654 0.0380882
R43066 PAD.n1768 PAD.n1654 0.0380882
R43067 PAD.n1768 PAD.n1656 0.0380882
R43068 PAD.n1764 PAD.n1656 0.0380882
R43069 PAD.n1764 PAD.n1658 0.0380882
R43070 PAD.n1756 PAD.n1658 0.0380882
R43071 PAD.n1756 PAD.n1660 0.0380882
R43072 PAD.n1752 PAD.n1660 0.0380882
R43073 PAD.n1752 PAD.n1662 0.0380882
R43074 PAD.n1744 PAD.n1662 0.0380882
R43075 PAD.n1744 PAD.n1664 0.0380882
R43076 PAD.n1740 PAD.n1664 0.0380882
R43077 PAD.n1740 PAD.n1666 0.0380882
R43078 PAD.n1732 PAD.n1666 0.0380882
R43079 PAD.n1732 PAD.n1668 0.0380882
R43080 PAD.n1728 PAD.n1668 0.0380882
R43081 PAD.n1728 PAD.n1670 0.0380882
R43082 PAD.n1720 PAD.n1670 0.0380882
R43083 PAD.n1720 PAD.n1672 0.0380882
R43084 PAD.n1716 PAD.n1672 0.0380882
R43085 PAD.n1716 PAD.n1674 0.0380882
R43086 PAD.n1708 PAD.n1674 0.0380882
R43087 PAD.n1708 PAD.n1676 0.0380882
R43088 PAD.n1704 PAD.n1676 0.0380882
R43089 PAD.n1704 PAD.n1678 0.0380882
R43090 PAD.n1696 PAD.n1678 0.0380882
R43091 PAD.n1696 PAD.n1680 0.0380882
R43092 PAD.n1692 PAD.n1680 0.0380882
R43093 PAD.n1692 PAD.n1682 0.0380882
R43094 PAD.n1684 PAD.n1682 0.0380882
R43095 PAD.n1932 PAD.n1598 0.0380882
R43096 PAD.n1604 PAD.n1598 0.0380882
R43097 PAD.n1923 PAD.n1604 0.0380882
R43098 PAD.n1923 PAD.n1922 0.0380882
R43099 PAD.n1922 PAD.n1921 0.0380882
R43100 PAD.n1921 PAD.n1605 0.0380882
R43101 PAD.n1911 PAD.n1605 0.0380882
R43102 PAD.n1911 PAD.n1910 0.0380882
R43103 PAD.n1910 PAD.n1909 0.0380882
R43104 PAD.n1909 PAD.n1609 0.0380882
R43105 PAD.n1899 PAD.n1609 0.0380882
R43106 PAD.n1899 PAD.n1898 0.0380882
R43107 PAD.n1898 PAD.n1897 0.0380882
R43108 PAD.n1897 PAD.n1613 0.0380882
R43109 PAD.n1887 PAD.n1613 0.0380882
R43110 PAD.n1887 PAD.n1886 0.0380882
R43111 PAD.n1886 PAD.n1885 0.0380882
R43112 PAD.n1885 PAD.n1617 0.0380882
R43113 PAD.n1875 PAD.n1617 0.0380882
R43114 PAD.n1875 PAD.n1874 0.0380882
R43115 PAD.n1874 PAD.n1873 0.0380882
R43116 PAD.n1873 PAD.n1621 0.0380882
R43117 PAD.n1863 PAD.n1621 0.0380882
R43118 PAD.n1863 PAD.n1862 0.0380882
R43119 PAD.n1862 PAD.n1861 0.0380882
R43120 PAD.n1861 PAD.n1625 0.0380882
R43121 PAD.n1851 PAD.n1625 0.0380882
R43122 PAD.n1851 PAD.n1850 0.0380882
R43123 PAD.n1850 PAD.n1849 0.0380882
R43124 PAD.n1849 PAD.n1629 0.0380882
R43125 PAD.n1839 PAD.n1629 0.0380882
R43126 PAD.n1839 PAD.n1838 0.0380882
R43127 PAD.n1838 PAD.n1837 0.0380882
R43128 PAD.n1837 PAD.n1633 0.0380882
R43129 PAD.n1827 PAD.n1633 0.0380882
R43130 PAD.n1827 PAD.n1826 0.0380882
R43131 PAD.n1826 PAD.n1825 0.0380882
R43132 PAD.n1825 PAD.n1637 0.0380882
R43133 PAD.n1815 PAD.n1637 0.0380882
R43134 PAD.n1815 PAD.n1814 0.0380882
R43135 PAD.n1814 PAD.n1813 0.0380882
R43136 PAD.n1813 PAD.n1641 0.0380882
R43137 PAD.n1803 PAD.n1641 0.0380882
R43138 PAD.n1803 PAD.n1802 0.0380882
R43139 PAD.n1802 PAD.n1801 0.0380882
R43140 PAD.n1801 PAD.n1645 0.0380882
R43141 PAD.n1791 PAD.n1645 0.0380882
R43142 PAD.n1791 PAD.n1790 0.0380882
R43143 PAD.n1790 PAD.n1789 0.0380882
R43144 PAD.n1789 PAD.n1649 0.0380882
R43145 PAD.n1779 PAD.n1649 0.0380882
R43146 PAD.n1779 PAD.n1778 0.0380882
R43147 PAD.n1778 PAD.n1777 0.0380882
R43148 PAD.n1777 PAD.n1653 0.0380882
R43149 PAD.n1767 PAD.n1653 0.0380882
R43150 PAD.n1767 PAD.n1766 0.0380882
R43151 PAD.n1766 PAD.n1765 0.0380882
R43152 PAD.n1765 PAD.n1657 0.0380882
R43153 PAD.n1755 PAD.n1657 0.0380882
R43154 PAD.n1755 PAD.n1754 0.0380882
R43155 PAD.n1754 PAD.n1753 0.0380882
R43156 PAD.n1753 PAD.n1661 0.0380882
R43157 PAD.n1743 PAD.n1661 0.0380882
R43158 PAD.n1743 PAD.n1742 0.0380882
R43159 PAD.n1742 PAD.n1741 0.0380882
R43160 PAD.n1741 PAD.n1665 0.0380882
R43161 PAD.n1731 PAD.n1665 0.0380882
R43162 PAD.n1731 PAD.n1730 0.0380882
R43163 PAD.n1730 PAD.n1729 0.0380882
R43164 PAD.n1729 PAD.n1669 0.0380882
R43165 PAD.n1719 PAD.n1669 0.0380882
R43166 PAD.n1719 PAD.n1718 0.0380882
R43167 PAD.n1718 PAD.n1717 0.0380882
R43168 PAD.n1717 PAD.n1673 0.0380882
R43169 PAD.n1707 PAD.n1673 0.0380882
R43170 PAD.n1707 PAD.n1706 0.0380882
R43171 PAD.n1706 PAD.n1705 0.0380882
R43172 PAD.n1705 PAD.n1677 0.0380882
R43173 PAD.n1695 PAD.n1677 0.0380882
R43174 PAD.n1695 PAD.n1694 0.0380882
R43175 PAD.n1694 PAD.n1693 0.0380882
R43176 PAD.n1693 PAD.n1681 0.0380882
R43177 PAD.n1683 PAD.n1681 0.0380882
R43178 PAD.n9463 PAD.n2031 0.0380882
R43179 PAD.n9467 PAD.n2031 0.0380882
R43180 PAD.n9471 PAD.n9467 0.0380882
R43181 PAD.n9475 PAD.n9471 0.0380882
R43182 PAD.n9475 PAD.n2027 0.0380882
R43183 PAD.n9479 PAD.n2027 0.0380882
R43184 PAD.n9483 PAD.n9479 0.0380882
R43185 PAD.n9487 PAD.n9483 0.0380882
R43186 PAD.n9487 PAD.n2025 0.0380882
R43187 PAD.n9491 PAD.n2025 0.0380882
R43188 PAD.n9495 PAD.n9491 0.0380882
R43189 PAD.n9499 PAD.n9495 0.0380882
R43190 PAD.n9499 PAD.n2023 0.0380882
R43191 PAD.n9503 PAD.n2023 0.0380882
R43192 PAD.n9507 PAD.n9503 0.0380882
R43193 PAD.n9511 PAD.n9507 0.0380882
R43194 PAD.n9511 PAD.n2021 0.0380882
R43195 PAD.n9515 PAD.n2021 0.0380882
R43196 PAD.n9519 PAD.n9515 0.0380882
R43197 PAD.n9523 PAD.n9519 0.0380882
R43198 PAD.n9523 PAD.n2019 0.0380882
R43199 PAD.n9527 PAD.n2019 0.0380882
R43200 PAD.n9531 PAD.n9527 0.0380882
R43201 PAD.n9535 PAD.n9531 0.0380882
R43202 PAD.n9535 PAD.n2017 0.0380882
R43203 PAD.n9539 PAD.n2017 0.0380882
R43204 PAD.n9543 PAD.n9539 0.0380882
R43205 PAD.n9547 PAD.n9543 0.0380882
R43206 PAD.n9547 PAD.n2015 0.0380882
R43207 PAD.n9551 PAD.n2015 0.0380882
R43208 PAD.n9555 PAD.n9551 0.0380882
R43209 PAD.n9559 PAD.n9555 0.0380882
R43210 PAD.n9559 PAD.n2013 0.0380882
R43211 PAD.n9563 PAD.n2013 0.0380882
R43212 PAD.n9567 PAD.n9563 0.0380882
R43213 PAD.n9571 PAD.n9567 0.0380882
R43214 PAD.n9571 PAD.n2011 0.0380882
R43215 PAD.n9575 PAD.n2011 0.0380882
R43216 PAD.n9579 PAD.n9575 0.0380882
R43217 PAD.n9583 PAD.n9579 0.0380882
R43218 PAD.n9583 PAD.n2009 0.0380882
R43219 PAD.n9587 PAD.n2009 0.0380882
R43220 PAD.n9591 PAD.n9587 0.0380882
R43221 PAD.n9595 PAD.n9591 0.0380882
R43222 PAD.n9595 PAD.n2007 0.0380882
R43223 PAD.n9599 PAD.n2007 0.0380882
R43224 PAD.n9603 PAD.n9599 0.0380882
R43225 PAD.n9607 PAD.n9603 0.0380882
R43226 PAD.n9607 PAD.n2005 0.0380882
R43227 PAD.n9611 PAD.n2005 0.0380882
R43228 PAD.n9615 PAD.n9611 0.0380882
R43229 PAD.n9619 PAD.n9615 0.0380882
R43230 PAD.n9619 PAD.n2003 0.0380882
R43231 PAD.n9623 PAD.n2003 0.0380882
R43232 PAD.n9627 PAD.n9623 0.0380882
R43233 PAD.n9631 PAD.n9627 0.0380882
R43234 PAD.n9631 PAD.n2001 0.0380882
R43235 PAD.n9635 PAD.n2001 0.0380882
R43236 PAD.n9639 PAD.n9635 0.0380882
R43237 PAD.n9643 PAD.n9639 0.0380882
R43238 PAD.n9643 PAD.n1999 0.0380882
R43239 PAD.n9647 PAD.n1999 0.0380882
R43240 PAD.n9651 PAD.n9647 0.0380882
R43241 PAD.n9655 PAD.n9651 0.0380882
R43242 PAD.n9655 PAD.n1997 0.0380882
R43243 PAD.n9659 PAD.n1997 0.0380882
R43244 PAD.n9663 PAD.n9659 0.0380882
R43245 PAD.n9667 PAD.n9663 0.0380882
R43246 PAD.n9667 PAD.n1995 0.0380882
R43247 PAD.n9671 PAD.n1995 0.0380882
R43248 PAD.n9675 PAD.n9671 0.0380882
R43249 PAD.n9679 PAD.n9675 0.0380882
R43250 PAD.n9679 PAD.n1993 0.0380882
R43251 PAD.n9683 PAD.n1993 0.0380882
R43252 PAD.n9687 PAD.n9683 0.0380882
R43253 PAD.n9691 PAD.n9687 0.0380882
R43254 PAD.n9691 PAD.n1991 0.0380882
R43255 PAD.n9695 PAD.n1991 0.0380882
R43256 PAD.n9699 PAD.n9695 0.0380882
R43257 PAD.n9703 PAD.n9699 0.0380882
R43258 PAD.n9703 PAD.n1989 0.0380882
R43259 PAD.n9708 PAD.n1989 0.0380882
R43260 PAD.n9708 PAD.n1987 0.0380882
R43261 PAD.n9465 PAD.n9464 0.0380882
R43262 PAD.n9466 PAD.n9465 0.0380882
R43263 PAD.n9466 PAD.n2028 0.0380882
R43264 PAD.n9476 PAD.n2028 0.0380882
R43265 PAD.n9477 PAD.n9476 0.0380882
R43266 PAD.n9478 PAD.n9477 0.0380882
R43267 PAD.n9478 PAD.n2026 0.0380882
R43268 PAD.n9488 PAD.n2026 0.0380882
R43269 PAD.n9489 PAD.n9488 0.0380882
R43270 PAD.n9490 PAD.n9489 0.0380882
R43271 PAD.n9490 PAD.n2024 0.0380882
R43272 PAD.n9500 PAD.n2024 0.0380882
R43273 PAD.n9501 PAD.n9500 0.0380882
R43274 PAD.n9502 PAD.n9501 0.0380882
R43275 PAD.n9502 PAD.n2022 0.0380882
R43276 PAD.n9512 PAD.n2022 0.0380882
R43277 PAD.n9513 PAD.n9512 0.0380882
R43278 PAD.n9514 PAD.n9513 0.0380882
R43279 PAD.n9514 PAD.n2020 0.0380882
R43280 PAD.n9524 PAD.n2020 0.0380882
R43281 PAD.n9525 PAD.n9524 0.0380882
R43282 PAD.n9526 PAD.n9525 0.0380882
R43283 PAD.n9526 PAD.n2018 0.0380882
R43284 PAD.n9536 PAD.n2018 0.0380882
R43285 PAD.n9537 PAD.n9536 0.0380882
R43286 PAD.n9538 PAD.n9537 0.0380882
R43287 PAD.n9538 PAD.n2016 0.0380882
R43288 PAD.n9548 PAD.n2016 0.0380882
R43289 PAD.n9549 PAD.n9548 0.0380882
R43290 PAD.n9550 PAD.n9549 0.0380882
R43291 PAD.n9550 PAD.n2014 0.0380882
R43292 PAD.n9560 PAD.n2014 0.0380882
R43293 PAD.n9561 PAD.n9560 0.0380882
R43294 PAD.n9562 PAD.n9561 0.0380882
R43295 PAD.n9562 PAD.n2012 0.0380882
R43296 PAD.n9572 PAD.n2012 0.0380882
R43297 PAD.n9573 PAD.n9572 0.0380882
R43298 PAD.n9574 PAD.n9573 0.0380882
R43299 PAD.n9574 PAD.n2010 0.0380882
R43300 PAD.n9584 PAD.n2010 0.0380882
R43301 PAD.n9585 PAD.n9584 0.0380882
R43302 PAD.n9586 PAD.n9585 0.0380882
R43303 PAD.n9586 PAD.n2008 0.0380882
R43304 PAD.n9596 PAD.n2008 0.0380882
R43305 PAD.n9597 PAD.n9596 0.0380882
R43306 PAD.n9598 PAD.n9597 0.0380882
R43307 PAD.n9598 PAD.n2006 0.0380882
R43308 PAD.n9608 PAD.n2006 0.0380882
R43309 PAD.n9609 PAD.n9608 0.0380882
R43310 PAD.n9610 PAD.n9609 0.0380882
R43311 PAD.n9610 PAD.n2004 0.0380882
R43312 PAD.n9620 PAD.n2004 0.0380882
R43313 PAD.n9621 PAD.n9620 0.0380882
R43314 PAD.n9622 PAD.n9621 0.0380882
R43315 PAD.n9622 PAD.n2002 0.0380882
R43316 PAD.n9632 PAD.n2002 0.0380882
R43317 PAD.n9633 PAD.n9632 0.0380882
R43318 PAD.n9634 PAD.n9633 0.0380882
R43319 PAD.n9634 PAD.n2000 0.0380882
R43320 PAD.n9644 PAD.n2000 0.0380882
R43321 PAD.n9645 PAD.n9644 0.0380882
R43322 PAD.n9646 PAD.n9645 0.0380882
R43323 PAD.n9646 PAD.n1998 0.0380882
R43324 PAD.n9656 PAD.n1998 0.0380882
R43325 PAD.n9657 PAD.n9656 0.0380882
R43326 PAD.n9658 PAD.n9657 0.0380882
R43327 PAD.n9658 PAD.n1996 0.0380882
R43328 PAD.n9668 PAD.n1996 0.0380882
R43329 PAD.n9669 PAD.n9668 0.0380882
R43330 PAD.n9670 PAD.n9669 0.0380882
R43331 PAD.n9670 PAD.n1994 0.0380882
R43332 PAD.n9680 PAD.n1994 0.0380882
R43333 PAD.n9681 PAD.n9680 0.0380882
R43334 PAD.n9682 PAD.n9681 0.0380882
R43335 PAD.n9682 PAD.n1992 0.0380882
R43336 PAD.n9692 PAD.n1992 0.0380882
R43337 PAD.n9693 PAD.n9692 0.0380882
R43338 PAD.n9694 PAD.n9693 0.0380882
R43339 PAD.n9694 PAD.n1990 0.0380882
R43340 PAD.n9704 PAD.n1990 0.0380882
R43341 PAD.n9705 PAD.n9704 0.0380882
R43342 PAD.n9707 PAD.n9705 0.0380882
R43343 PAD.n9707 PAD.n9706 0.0380882
R43344 PAD.n9197 PAD.n2134 0.0380882
R43345 PAD.n9201 PAD.n2134 0.0380882
R43346 PAD.n9205 PAD.n9201 0.0380882
R43347 PAD.n9209 PAD.n9205 0.0380882
R43348 PAD.n9209 PAD.n2130 0.0380882
R43349 PAD.n9213 PAD.n2130 0.0380882
R43350 PAD.n9217 PAD.n9213 0.0380882
R43351 PAD.n9221 PAD.n9217 0.0380882
R43352 PAD.n9221 PAD.n2128 0.0380882
R43353 PAD.n9225 PAD.n2128 0.0380882
R43354 PAD.n9229 PAD.n9225 0.0380882
R43355 PAD.n9233 PAD.n9229 0.0380882
R43356 PAD.n9233 PAD.n2126 0.0380882
R43357 PAD.n9237 PAD.n2126 0.0380882
R43358 PAD.n9241 PAD.n9237 0.0380882
R43359 PAD.n9245 PAD.n9241 0.0380882
R43360 PAD.n9245 PAD.n2124 0.0380882
R43361 PAD.n9249 PAD.n2124 0.0380882
R43362 PAD.n9253 PAD.n9249 0.0380882
R43363 PAD.n9257 PAD.n9253 0.0380882
R43364 PAD.n9257 PAD.n2122 0.0380882
R43365 PAD.n9261 PAD.n2122 0.0380882
R43366 PAD.n9265 PAD.n9261 0.0380882
R43367 PAD.n9269 PAD.n9265 0.0380882
R43368 PAD.n9269 PAD.n2120 0.0380882
R43369 PAD.n9273 PAD.n2120 0.0380882
R43370 PAD.n9277 PAD.n9273 0.0380882
R43371 PAD.n9281 PAD.n9277 0.0380882
R43372 PAD.n9281 PAD.n2118 0.0380882
R43373 PAD.n9285 PAD.n2118 0.0380882
R43374 PAD.n9289 PAD.n9285 0.0380882
R43375 PAD.n9293 PAD.n9289 0.0380882
R43376 PAD.n9293 PAD.n2116 0.0380882
R43377 PAD.n9297 PAD.n2116 0.0380882
R43378 PAD.n9301 PAD.n9297 0.0380882
R43379 PAD.n9305 PAD.n9301 0.0380882
R43380 PAD.n9305 PAD.n2114 0.0380882
R43381 PAD.n9309 PAD.n2114 0.0380882
R43382 PAD.n9313 PAD.n9309 0.0380882
R43383 PAD.n9317 PAD.n9313 0.0380882
R43384 PAD.n9317 PAD.n2112 0.0380882
R43385 PAD.n9321 PAD.n2112 0.0380882
R43386 PAD.n9325 PAD.n9321 0.0380882
R43387 PAD.n9329 PAD.n9325 0.0380882
R43388 PAD.n9329 PAD.n2110 0.0380882
R43389 PAD.n9333 PAD.n2110 0.0380882
R43390 PAD.n9337 PAD.n9333 0.0380882
R43391 PAD.n9341 PAD.n9337 0.0380882
R43392 PAD.n9341 PAD.n2108 0.0380882
R43393 PAD.n9345 PAD.n2108 0.0380882
R43394 PAD.n9349 PAD.n9345 0.0380882
R43395 PAD.n9353 PAD.n9349 0.0380882
R43396 PAD.n9353 PAD.n2106 0.0380882
R43397 PAD.n9357 PAD.n2106 0.0380882
R43398 PAD.n9361 PAD.n9357 0.0380882
R43399 PAD.n9365 PAD.n9361 0.0380882
R43400 PAD.n9365 PAD.n2104 0.0380882
R43401 PAD.n9369 PAD.n2104 0.0380882
R43402 PAD.n9373 PAD.n9369 0.0380882
R43403 PAD.n9377 PAD.n9373 0.0380882
R43404 PAD.n9377 PAD.n2102 0.0380882
R43405 PAD.n9381 PAD.n2102 0.0380882
R43406 PAD.n9385 PAD.n9381 0.0380882
R43407 PAD.n9389 PAD.n9385 0.0380882
R43408 PAD.n9389 PAD.n2100 0.0380882
R43409 PAD.n9393 PAD.n2100 0.0380882
R43410 PAD.n9397 PAD.n9393 0.0380882
R43411 PAD.n9401 PAD.n9397 0.0380882
R43412 PAD.n9401 PAD.n2098 0.0380882
R43413 PAD.n9405 PAD.n2098 0.0380882
R43414 PAD.n9409 PAD.n9405 0.0380882
R43415 PAD.n9413 PAD.n9409 0.0380882
R43416 PAD.n9413 PAD.n2096 0.0380882
R43417 PAD.n9417 PAD.n2096 0.0380882
R43418 PAD.n9421 PAD.n9417 0.0380882
R43419 PAD.n9425 PAD.n9421 0.0380882
R43420 PAD.n9425 PAD.n2094 0.0380882
R43421 PAD.n9429 PAD.n2094 0.0380882
R43422 PAD.n9433 PAD.n9429 0.0380882
R43423 PAD.n9437 PAD.n9433 0.0380882
R43424 PAD.n9437 PAD.n2092 0.0380882
R43425 PAD.n9441 PAD.n2092 0.0380882
R43426 PAD.n9441 PAD.n2090 0.0380882
R43427 PAD.n9199 PAD.n9198 0.0380882
R43428 PAD.n9200 PAD.n9199 0.0380882
R43429 PAD.n9200 PAD.n2131 0.0380882
R43430 PAD.n9210 PAD.n2131 0.0380882
R43431 PAD.n9211 PAD.n9210 0.0380882
R43432 PAD.n9212 PAD.n9211 0.0380882
R43433 PAD.n9212 PAD.n2129 0.0380882
R43434 PAD.n9222 PAD.n2129 0.0380882
R43435 PAD.n9223 PAD.n9222 0.0380882
R43436 PAD.n9224 PAD.n9223 0.0380882
R43437 PAD.n9224 PAD.n2127 0.0380882
R43438 PAD.n9234 PAD.n2127 0.0380882
R43439 PAD.n9235 PAD.n9234 0.0380882
R43440 PAD.n9236 PAD.n9235 0.0380882
R43441 PAD.n9236 PAD.n2125 0.0380882
R43442 PAD.n9246 PAD.n2125 0.0380882
R43443 PAD.n9247 PAD.n9246 0.0380882
R43444 PAD.n9248 PAD.n9247 0.0380882
R43445 PAD.n9248 PAD.n2123 0.0380882
R43446 PAD.n9258 PAD.n2123 0.0380882
R43447 PAD.n9259 PAD.n9258 0.0380882
R43448 PAD.n9260 PAD.n9259 0.0380882
R43449 PAD.n9260 PAD.n2121 0.0380882
R43450 PAD.n9270 PAD.n2121 0.0380882
R43451 PAD.n9271 PAD.n9270 0.0380882
R43452 PAD.n9272 PAD.n9271 0.0380882
R43453 PAD.n9272 PAD.n2119 0.0380882
R43454 PAD.n9282 PAD.n2119 0.0380882
R43455 PAD.n9283 PAD.n9282 0.0380882
R43456 PAD.n9284 PAD.n9283 0.0380882
R43457 PAD.n9284 PAD.n2117 0.0380882
R43458 PAD.n9294 PAD.n2117 0.0380882
R43459 PAD.n9295 PAD.n9294 0.0380882
R43460 PAD.n9296 PAD.n9295 0.0380882
R43461 PAD.n9296 PAD.n2115 0.0380882
R43462 PAD.n9306 PAD.n2115 0.0380882
R43463 PAD.n9307 PAD.n9306 0.0380882
R43464 PAD.n9308 PAD.n9307 0.0380882
R43465 PAD.n9308 PAD.n2113 0.0380882
R43466 PAD.n9318 PAD.n2113 0.0380882
R43467 PAD.n9319 PAD.n9318 0.0380882
R43468 PAD.n9320 PAD.n9319 0.0380882
R43469 PAD.n9320 PAD.n2111 0.0380882
R43470 PAD.n9330 PAD.n2111 0.0380882
R43471 PAD.n9331 PAD.n9330 0.0380882
R43472 PAD.n9332 PAD.n9331 0.0380882
R43473 PAD.n9332 PAD.n2109 0.0380882
R43474 PAD.n9342 PAD.n2109 0.0380882
R43475 PAD.n9343 PAD.n9342 0.0380882
R43476 PAD.n9344 PAD.n9343 0.0380882
R43477 PAD.n9344 PAD.n2107 0.0380882
R43478 PAD.n9354 PAD.n2107 0.0380882
R43479 PAD.n9355 PAD.n9354 0.0380882
R43480 PAD.n9356 PAD.n9355 0.0380882
R43481 PAD.n9356 PAD.n2105 0.0380882
R43482 PAD.n9366 PAD.n2105 0.0380882
R43483 PAD.n9367 PAD.n9366 0.0380882
R43484 PAD.n9368 PAD.n9367 0.0380882
R43485 PAD.n9368 PAD.n2103 0.0380882
R43486 PAD.n9378 PAD.n2103 0.0380882
R43487 PAD.n9379 PAD.n9378 0.0380882
R43488 PAD.n9380 PAD.n9379 0.0380882
R43489 PAD.n9380 PAD.n2101 0.0380882
R43490 PAD.n9390 PAD.n2101 0.0380882
R43491 PAD.n9391 PAD.n9390 0.0380882
R43492 PAD.n9392 PAD.n9391 0.0380882
R43493 PAD.n9392 PAD.n2099 0.0380882
R43494 PAD.n9402 PAD.n2099 0.0380882
R43495 PAD.n9403 PAD.n9402 0.0380882
R43496 PAD.n9404 PAD.n9403 0.0380882
R43497 PAD.n9404 PAD.n2097 0.0380882
R43498 PAD.n9414 PAD.n2097 0.0380882
R43499 PAD.n9415 PAD.n9414 0.0380882
R43500 PAD.n9416 PAD.n9415 0.0380882
R43501 PAD.n9416 PAD.n2095 0.0380882
R43502 PAD.n9426 PAD.n2095 0.0380882
R43503 PAD.n9427 PAD.n9426 0.0380882
R43504 PAD.n9428 PAD.n9427 0.0380882
R43505 PAD.n9428 PAD.n2093 0.0380882
R43506 PAD.n9438 PAD.n2093 0.0380882
R43507 PAD.n9439 PAD.n9438 0.0380882
R43508 PAD.n9440 PAD.n9439 0.0380882
R43509 PAD.n9440 PAD.n2040 0.0380882
R43510 PAD.n2482 PAD.n2481 0.0380882
R43511 PAD.n2481 PAD.n2152 0.0380882
R43512 PAD.n2475 PAD.n2152 0.0380882
R43513 PAD.n2475 PAD.n2155 0.0380882
R43514 PAD.n2471 PAD.n2155 0.0380882
R43515 PAD.n2471 PAD.n2158 0.0380882
R43516 PAD.n2463 PAD.n2158 0.0380882
R43517 PAD.n2463 PAD.n2160 0.0380882
R43518 PAD.n2459 PAD.n2160 0.0380882
R43519 PAD.n2459 PAD.n2162 0.0380882
R43520 PAD.n2451 PAD.n2162 0.0380882
R43521 PAD.n2451 PAD.n2164 0.0380882
R43522 PAD.n2447 PAD.n2164 0.0380882
R43523 PAD.n2447 PAD.n2166 0.0380882
R43524 PAD.n2439 PAD.n2166 0.0380882
R43525 PAD.n2439 PAD.n2168 0.0380882
R43526 PAD.n2435 PAD.n2168 0.0380882
R43527 PAD.n2435 PAD.n2170 0.0380882
R43528 PAD.n2427 PAD.n2170 0.0380882
R43529 PAD.n2427 PAD.n2172 0.0380882
R43530 PAD.n2423 PAD.n2172 0.0380882
R43531 PAD.n2423 PAD.n2174 0.0380882
R43532 PAD.n2415 PAD.n2174 0.0380882
R43533 PAD.n2415 PAD.n2176 0.0380882
R43534 PAD.n2411 PAD.n2176 0.0380882
R43535 PAD.n2411 PAD.n2178 0.0380882
R43536 PAD.n2403 PAD.n2178 0.0380882
R43537 PAD.n2403 PAD.n2180 0.0380882
R43538 PAD.n2399 PAD.n2180 0.0380882
R43539 PAD.n2399 PAD.n2182 0.0380882
R43540 PAD.n2391 PAD.n2182 0.0380882
R43541 PAD.n2391 PAD.n2184 0.0380882
R43542 PAD.n2387 PAD.n2184 0.0380882
R43543 PAD.n2387 PAD.n2186 0.0380882
R43544 PAD.n2379 PAD.n2186 0.0380882
R43545 PAD.n2379 PAD.n2188 0.0380882
R43546 PAD.n2375 PAD.n2188 0.0380882
R43547 PAD.n2375 PAD.n2190 0.0380882
R43548 PAD.n2367 PAD.n2190 0.0380882
R43549 PAD.n2367 PAD.n2192 0.0380882
R43550 PAD.n2363 PAD.n2192 0.0380882
R43551 PAD.n2363 PAD.n2194 0.0380882
R43552 PAD.n2355 PAD.n2194 0.0380882
R43553 PAD.n2355 PAD.n2196 0.0380882
R43554 PAD.n2351 PAD.n2196 0.0380882
R43555 PAD.n2351 PAD.n2198 0.0380882
R43556 PAD.n2343 PAD.n2198 0.0380882
R43557 PAD.n2343 PAD.n2200 0.0380882
R43558 PAD.n2339 PAD.n2200 0.0380882
R43559 PAD.n2339 PAD.n2202 0.0380882
R43560 PAD.n2331 PAD.n2202 0.0380882
R43561 PAD.n2331 PAD.n2204 0.0380882
R43562 PAD.n2327 PAD.n2204 0.0380882
R43563 PAD.n2327 PAD.n2206 0.0380882
R43564 PAD.n2319 PAD.n2206 0.0380882
R43565 PAD.n2319 PAD.n2208 0.0380882
R43566 PAD.n2315 PAD.n2208 0.0380882
R43567 PAD.n2315 PAD.n2210 0.0380882
R43568 PAD.n2307 PAD.n2210 0.0380882
R43569 PAD.n2307 PAD.n2212 0.0380882
R43570 PAD.n2303 PAD.n2212 0.0380882
R43571 PAD.n2303 PAD.n2214 0.0380882
R43572 PAD.n2295 PAD.n2214 0.0380882
R43573 PAD.n2295 PAD.n2216 0.0380882
R43574 PAD.n2291 PAD.n2216 0.0380882
R43575 PAD.n2291 PAD.n2218 0.0380882
R43576 PAD.n2283 PAD.n2218 0.0380882
R43577 PAD.n2283 PAD.n2220 0.0380882
R43578 PAD.n2279 PAD.n2220 0.0380882
R43579 PAD.n2279 PAD.n2222 0.0380882
R43580 PAD.n2271 PAD.n2222 0.0380882
R43581 PAD.n2271 PAD.n2224 0.0380882
R43582 PAD.n2267 PAD.n2224 0.0380882
R43583 PAD.n2267 PAD.n2226 0.0380882
R43584 PAD.n2259 PAD.n2226 0.0380882
R43585 PAD.n2259 PAD.n2228 0.0380882
R43586 PAD.n2255 PAD.n2228 0.0380882
R43587 PAD.n2255 PAD.n2230 0.0380882
R43588 PAD.n2247 PAD.n2230 0.0380882
R43589 PAD.n2247 PAD.n2232 0.0380882
R43590 PAD.n2243 PAD.n2232 0.0380882
R43591 PAD.n2243 PAD.n2234 0.0380882
R43592 PAD.n2235 PAD.n2234 0.0380882
R43593 PAD.n2483 PAD.n2150 0.0380882
R43594 PAD.n2156 PAD.n2150 0.0380882
R43595 PAD.n2474 PAD.n2156 0.0380882
R43596 PAD.n2474 PAD.n2473 0.0380882
R43597 PAD.n2473 PAD.n2472 0.0380882
R43598 PAD.n2472 PAD.n2157 0.0380882
R43599 PAD.n2462 PAD.n2157 0.0380882
R43600 PAD.n2462 PAD.n2461 0.0380882
R43601 PAD.n2461 PAD.n2460 0.0380882
R43602 PAD.n2460 PAD.n2161 0.0380882
R43603 PAD.n2450 PAD.n2161 0.0380882
R43604 PAD.n2450 PAD.n2449 0.0380882
R43605 PAD.n2449 PAD.n2448 0.0380882
R43606 PAD.n2448 PAD.n2165 0.0380882
R43607 PAD.n2438 PAD.n2165 0.0380882
R43608 PAD.n2438 PAD.n2437 0.0380882
R43609 PAD.n2437 PAD.n2436 0.0380882
R43610 PAD.n2436 PAD.n2169 0.0380882
R43611 PAD.n2426 PAD.n2169 0.0380882
R43612 PAD.n2426 PAD.n2425 0.0380882
R43613 PAD.n2425 PAD.n2424 0.0380882
R43614 PAD.n2424 PAD.n2173 0.0380882
R43615 PAD.n2414 PAD.n2173 0.0380882
R43616 PAD.n2414 PAD.n2413 0.0380882
R43617 PAD.n2413 PAD.n2412 0.0380882
R43618 PAD.n2412 PAD.n2177 0.0380882
R43619 PAD.n2402 PAD.n2177 0.0380882
R43620 PAD.n2402 PAD.n2401 0.0380882
R43621 PAD.n2401 PAD.n2400 0.0380882
R43622 PAD.n2400 PAD.n2181 0.0380882
R43623 PAD.n2390 PAD.n2181 0.0380882
R43624 PAD.n2390 PAD.n2389 0.0380882
R43625 PAD.n2389 PAD.n2388 0.0380882
R43626 PAD.n2388 PAD.n2185 0.0380882
R43627 PAD.n2378 PAD.n2185 0.0380882
R43628 PAD.n2378 PAD.n2377 0.0380882
R43629 PAD.n2377 PAD.n2376 0.0380882
R43630 PAD.n2376 PAD.n2189 0.0380882
R43631 PAD.n2366 PAD.n2189 0.0380882
R43632 PAD.n2366 PAD.n2365 0.0380882
R43633 PAD.n2365 PAD.n2364 0.0380882
R43634 PAD.n2364 PAD.n2193 0.0380882
R43635 PAD.n2354 PAD.n2193 0.0380882
R43636 PAD.n2354 PAD.n2353 0.0380882
R43637 PAD.n2353 PAD.n2352 0.0380882
R43638 PAD.n2352 PAD.n2197 0.0380882
R43639 PAD.n2342 PAD.n2197 0.0380882
R43640 PAD.n2342 PAD.n2341 0.0380882
R43641 PAD.n2341 PAD.n2340 0.0380882
R43642 PAD.n2340 PAD.n2201 0.0380882
R43643 PAD.n2330 PAD.n2201 0.0380882
R43644 PAD.n2330 PAD.n2329 0.0380882
R43645 PAD.n2329 PAD.n2328 0.0380882
R43646 PAD.n2328 PAD.n2205 0.0380882
R43647 PAD.n2318 PAD.n2205 0.0380882
R43648 PAD.n2318 PAD.n2317 0.0380882
R43649 PAD.n2317 PAD.n2316 0.0380882
R43650 PAD.n2316 PAD.n2209 0.0380882
R43651 PAD.n2306 PAD.n2209 0.0380882
R43652 PAD.n2306 PAD.n2305 0.0380882
R43653 PAD.n2305 PAD.n2304 0.0380882
R43654 PAD.n2304 PAD.n2213 0.0380882
R43655 PAD.n2294 PAD.n2213 0.0380882
R43656 PAD.n2294 PAD.n2293 0.0380882
R43657 PAD.n2293 PAD.n2292 0.0380882
R43658 PAD.n2292 PAD.n2217 0.0380882
R43659 PAD.n2282 PAD.n2217 0.0380882
R43660 PAD.n2282 PAD.n2281 0.0380882
R43661 PAD.n2281 PAD.n2280 0.0380882
R43662 PAD.n2280 PAD.n2221 0.0380882
R43663 PAD.n2270 PAD.n2221 0.0380882
R43664 PAD.n2270 PAD.n2269 0.0380882
R43665 PAD.n2269 PAD.n2268 0.0380882
R43666 PAD.n2268 PAD.n2225 0.0380882
R43667 PAD.n2258 PAD.n2225 0.0380882
R43668 PAD.n2258 PAD.n2257 0.0380882
R43669 PAD.n2257 PAD.n2256 0.0380882
R43670 PAD.n2256 PAD.n2229 0.0380882
R43671 PAD.n2246 PAD.n2229 0.0380882
R43672 PAD.n2246 PAD.n2245 0.0380882
R43673 PAD.n2245 PAD.n2244 0.0380882
R43674 PAD.n2244 PAD.n2233 0.0380882
R43675 PAD.n2233 PAD.n2142 0.0380882
R43676 PAD.n2829 PAD.n2828 0.0380882
R43677 PAD.n2828 PAD.n2499 0.0380882
R43678 PAD.n2822 PAD.n2499 0.0380882
R43679 PAD.n2822 PAD.n2502 0.0380882
R43680 PAD.n2818 PAD.n2502 0.0380882
R43681 PAD.n2818 PAD.n2505 0.0380882
R43682 PAD.n2810 PAD.n2505 0.0380882
R43683 PAD.n2810 PAD.n2507 0.0380882
R43684 PAD.n2806 PAD.n2507 0.0380882
R43685 PAD.n2806 PAD.n2509 0.0380882
R43686 PAD.n2798 PAD.n2509 0.0380882
R43687 PAD.n2798 PAD.n2511 0.0380882
R43688 PAD.n2794 PAD.n2511 0.0380882
R43689 PAD.n2794 PAD.n2513 0.0380882
R43690 PAD.n2786 PAD.n2513 0.0380882
R43691 PAD.n2786 PAD.n2515 0.0380882
R43692 PAD.n2782 PAD.n2515 0.0380882
R43693 PAD.n2782 PAD.n2517 0.0380882
R43694 PAD.n2774 PAD.n2517 0.0380882
R43695 PAD.n2774 PAD.n2519 0.0380882
R43696 PAD.n2770 PAD.n2519 0.0380882
R43697 PAD.n2770 PAD.n2521 0.0380882
R43698 PAD.n2762 PAD.n2521 0.0380882
R43699 PAD.n2762 PAD.n2523 0.0380882
R43700 PAD.n2758 PAD.n2523 0.0380882
R43701 PAD.n2758 PAD.n2525 0.0380882
R43702 PAD.n2750 PAD.n2525 0.0380882
R43703 PAD.n2750 PAD.n2527 0.0380882
R43704 PAD.n2746 PAD.n2527 0.0380882
R43705 PAD.n2746 PAD.n2529 0.0380882
R43706 PAD.n2738 PAD.n2529 0.0380882
R43707 PAD.n2738 PAD.n2531 0.0380882
R43708 PAD.n2734 PAD.n2531 0.0380882
R43709 PAD.n2734 PAD.n2533 0.0380882
R43710 PAD.n2726 PAD.n2533 0.0380882
R43711 PAD.n2726 PAD.n2535 0.0380882
R43712 PAD.n2722 PAD.n2535 0.0380882
R43713 PAD.n2722 PAD.n2537 0.0380882
R43714 PAD.n2714 PAD.n2537 0.0380882
R43715 PAD.n2714 PAD.n2539 0.0380882
R43716 PAD.n2710 PAD.n2539 0.0380882
R43717 PAD.n2710 PAD.n2541 0.0380882
R43718 PAD.n2702 PAD.n2541 0.0380882
R43719 PAD.n2702 PAD.n2543 0.0380882
R43720 PAD.n2698 PAD.n2543 0.0380882
R43721 PAD.n2698 PAD.n2545 0.0380882
R43722 PAD.n2690 PAD.n2545 0.0380882
R43723 PAD.n2690 PAD.n2547 0.0380882
R43724 PAD.n2686 PAD.n2547 0.0380882
R43725 PAD.n2686 PAD.n2549 0.0380882
R43726 PAD.n2678 PAD.n2549 0.0380882
R43727 PAD.n2678 PAD.n2551 0.0380882
R43728 PAD.n2674 PAD.n2551 0.0380882
R43729 PAD.n2674 PAD.n2553 0.0380882
R43730 PAD.n2666 PAD.n2553 0.0380882
R43731 PAD.n2666 PAD.n2555 0.0380882
R43732 PAD.n2662 PAD.n2555 0.0380882
R43733 PAD.n2662 PAD.n2557 0.0380882
R43734 PAD.n2654 PAD.n2557 0.0380882
R43735 PAD.n2654 PAD.n2559 0.0380882
R43736 PAD.n2650 PAD.n2559 0.0380882
R43737 PAD.n2650 PAD.n2561 0.0380882
R43738 PAD.n2642 PAD.n2561 0.0380882
R43739 PAD.n2642 PAD.n2563 0.0380882
R43740 PAD.n2638 PAD.n2563 0.0380882
R43741 PAD.n2638 PAD.n2565 0.0380882
R43742 PAD.n2630 PAD.n2565 0.0380882
R43743 PAD.n2630 PAD.n2567 0.0380882
R43744 PAD.n2626 PAD.n2567 0.0380882
R43745 PAD.n2626 PAD.n2569 0.0380882
R43746 PAD.n2618 PAD.n2569 0.0380882
R43747 PAD.n2618 PAD.n2571 0.0380882
R43748 PAD.n2614 PAD.n2571 0.0380882
R43749 PAD.n2614 PAD.n2573 0.0380882
R43750 PAD.n2606 PAD.n2573 0.0380882
R43751 PAD.n2606 PAD.n2575 0.0380882
R43752 PAD.n2602 PAD.n2575 0.0380882
R43753 PAD.n2602 PAD.n2577 0.0380882
R43754 PAD.n2594 PAD.n2577 0.0380882
R43755 PAD.n2594 PAD.n2579 0.0380882
R43756 PAD.n2590 PAD.n2579 0.0380882
R43757 PAD.n2590 PAD.n2581 0.0380882
R43758 PAD.n2582 PAD.n2581 0.0380882
R43759 PAD.n2830 PAD.n2497 0.0380882
R43760 PAD.n2503 PAD.n2497 0.0380882
R43761 PAD.n2821 PAD.n2503 0.0380882
R43762 PAD.n2821 PAD.n2820 0.0380882
R43763 PAD.n2820 PAD.n2819 0.0380882
R43764 PAD.n2819 PAD.n2504 0.0380882
R43765 PAD.n2809 PAD.n2504 0.0380882
R43766 PAD.n2809 PAD.n2808 0.0380882
R43767 PAD.n2808 PAD.n2807 0.0380882
R43768 PAD.n2807 PAD.n2508 0.0380882
R43769 PAD.n2797 PAD.n2508 0.0380882
R43770 PAD.n2797 PAD.n2796 0.0380882
R43771 PAD.n2796 PAD.n2795 0.0380882
R43772 PAD.n2795 PAD.n2512 0.0380882
R43773 PAD.n2785 PAD.n2512 0.0380882
R43774 PAD.n2785 PAD.n2784 0.0380882
R43775 PAD.n2784 PAD.n2783 0.0380882
R43776 PAD.n2783 PAD.n2516 0.0380882
R43777 PAD.n2773 PAD.n2516 0.0380882
R43778 PAD.n2773 PAD.n2772 0.0380882
R43779 PAD.n2772 PAD.n2771 0.0380882
R43780 PAD.n2771 PAD.n2520 0.0380882
R43781 PAD.n2761 PAD.n2520 0.0380882
R43782 PAD.n2761 PAD.n2760 0.0380882
R43783 PAD.n2760 PAD.n2759 0.0380882
R43784 PAD.n2759 PAD.n2524 0.0380882
R43785 PAD.n2749 PAD.n2524 0.0380882
R43786 PAD.n2749 PAD.n2748 0.0380882
R43787 PAD.n2748 PAD.n2747 0.0380882
R43788 PAD.n2747 PAD.n2528 0.0380882
R43789 PAD.n2737 PAD.n2528 0.0380882
R43790 PAD.n2737 PAD.n2736 0.0380882
R43791 PAD.n2736 PAD.n2735 0.0380882
R43792 PAD.n2735 PAD.n2532 0.0380882
R43793 PAD.n2725 PAD.n2532 0.0380882
R43794 PAD.n2725 PAD.n2724 0.0380882
R43795 PAD.n2724 PAD.n2723 0.0380882
R43796 PAD.n2723 PAD.n2536 0.0380882
R43797 PAD.n2713 PAD.n2536 0.0380882
R43798 PAD.n2713 PAD.n2712 0.0380882
R43799 PAD.n2712 PAD.n2711 0.0380882
R43800 PAD.n2711 PAD.n2540 0.0380882
R43801 PAD.n2701 PAD.n2540 0.0380882
R43802 PAD.n2701 PAD.n2700 0.0380882
R43803 PAD.n2700 PAD.n2699 0.0380882
R43804 PAD.n2699 PAD.n2544 0.0380882
R43805 PAD.n2689 PAD.n2544 0.0380882
R43806 PAD.n2689 PAD.n2688 0.0380882
R43807 PAD.n2688 PAD.n2687 0.0380882
R43808 PAD.n2687 PAD.n2548 0.0380882
R43809 PAD.n2677 PAD.n2548 0.0380882
R43810 PAD.n2677 PAD.n2676 0.0380882
R43811 PAD.n2676 PAD.n2675 0.0380882
R43812 PAD.n2675 PAD.n2552 0.0380882
R43813 PAD.n2665 PAD.n2552 0.0380882
R43814 PAD.n2665 PAD.n2664 0.0380882
R43815 PAD.n2664 PAD.n2663 0.0380882
R43816 PAD.n2663 PAD.n2556 0.0380882
R43817 PAD.n2653 PAD.n2556 0.0380882
R43818 PAD.n2653 PAD.n2652 0.0380882
R43819 PAD.n2652 PAD.n2651 0.0380882
R43820 PAD.n2651 PAD.n2560 0.0380882
R43821 PAD.n2641 PAD.n2560 0.0380882
R43822 PAD.n2641 PAD.n2640 0.0380882
R43823 PAD.n2640 PAD.n2639 0.0380882
R43824 PAD.n2639 PAD.n2564 0.0380882
R43825 PAD.n2629 PAD.n2564 0.0380882
R43826 PAD.n2629 PAD.n2628 0.0380882
R43827 PAD.n2628 PAD.n2627 0.0380882
R43828 PAD.n2627 PAD.n2568 0.0380882
R43829 PAD.n2617 PAD.n2568 0.0380882
R43830 PAD.n2617 PAD.n2616 0.0380882
R43831 PAD.n2616 PAD.n2615 0.0380882
R43832 PAD.n2615 PAD.n2572 0.0380882
R43833 PAD.n2605 PAD.n2572 0.0380882
R43834 PAD.n2605 PAD.n2604 0.0380882
R43835 PAD.n2604 PAD.n2603 0.0380882
R43836 PAD.n2603 PAD.n2576 0.0380882
R43837 PAD.n2593 PAD.n2576 0.0380882
R43838 PAD.n2593 PAD.n2592 0.0380882
R43839 PAD.n2592 PAD.n2591 0.0380882
R43840 PAD.n2591 PAD.n2580 0.0380882
R43841 PAD.n2580 PAD.n2490 0.0380882
R43842 PAD.n9119 PAD.n9118 0.0380882
R43843 PAD.n9118 PAD.n9115 0.0380882
R43844 PAD.n9115 PAD.n8838 0.0380882
R43845 PAD.n9111 PAD.n8838 0.0380882
R43846 PAD.n9111 PAD.n9107 0.0380882
R43847 PAD.n9107 PAD.n9106 0.0380882
R43848 PAD.n9106 PAD.n8843 0.0380882
R43849 PAD.n9102 PAD.n8843 0.0380882
R43850 PAD.n9102 PAD.n9098 0.0380882
R43851 PAD.n9098 PAD.n9097 0.0380882
R43852 PAD.n9097 PAD.n8848 0.0380882
R43853 PAD.n9093 PAD.n8848 0.0380882
R43854 PAD.n9093 PAD.n9089 0.0380882
R43855 PAD.n9089 PAD.n9088 0.0380882
R43856 PAD.n9088 PAD.n8853 0.0380882
R43857 PAD.n9084 PAD.n8853 0.0380882
R43858 PAD.n9084 PAD.n9080 0.0380882
R43859 PAD.n9080 PAD.n9079 0.0380882
R43860 PAD.n9079 PAD.n8858 0.0380882
R43861 PAD.n9075 PAD.n8858 0.0380882
R43862 PAD.n9075 PAD.n9071 0.0380882
R43863 PAD.n9071 PAD.n9070 0.0380882
R43864 PAD.n9070 PAD.n8863 0.0380882
R43865 PAD.n9066 PAD.n8863 0.0380882
R43866 PAD.n9066 PAD.n9062 0.0380882
R43867 PAD.n9062 PAD.n9061 0.0380882
R43868 PAD.n9061 PAD.n8868 0.0380882
R43869 PAD.n9057 PAD.n8868 0.0380882
R43870 PAD.n9057 PAD.n9053 0.0380882
R43871 PAD.n9053 PAD.n9052 0.0380882
R43872 PAD.n9052 PAD.n8873 0.0380882
R43873 PAD.n9048 PAD.n8873 0.0380882
R43874 PAD.n9048 PAD.n9044 0.0380882
R43875 PAD.n9044 PAD.n9043 0.0380882
R43876 PAD.n9043 PAD.n8878 0.0380882
R43877 PAD.n9039 PAD.n8878 0.0380882
R43878 PAD.n9039 PAD.n9035 0.0380882
R43879 PAD.n9035 PAD.n9034 0.0380882
R43880 PAD.n9034 PAD.n8883 0.0380882
R43881 PAD.n9030 PAD.n8883 0.0380882
R43882 PAD.n9030 PAD.n9026 0.0380882
R43883 PAD.n9026 PAD.n9025 0.0380882
R43884 PAD.n9025 PAD.n8888 0.0380882
R43885 PAD.n9021 PAD.n8888 0.0380882
R43886 PAD.n9021 PAD.n9017 0.0380882
R43887 PAD.n9017 PAD.n9016 0.0380882
R43888 PAD.n9016 PAD.n8893 0.0380882
R43889 PAD.n9012 PAD.n8893 0.0380882
R43890 PAD.n9012 PAD.n9008 0.0380882
R43891 PAD.n9008 PAD.n9007 0.0380882
R43892 PAD.n9007 PAD.n8898 0.0380882
R43893 PAD.n9003 PAD.n8898 0.0380882
R43894 PAD.n9003 PAD.n8999 0.0380882
R43895 PAD.n8999 PAD.n8998 0.0380882
R43896 PAD.n8998 PAD.n8903 0.0380882
R43897 PAD.n8994 PAD.n8903 0.0380882
R43898 PAD.n8994 PAD.n8990 0.0380882
R43899 PAD.n8990 PAD.n8989 0.0380882
R43900 PAD.n8989 PAD.n8908 0.0380882
R43901 PAD.n8985 PAD.n8908 0.0380882
R43902 PAD.n8985 PAD.n8981 0.0380882
R43903 PAD.n8981 PAD.n8980 0.0380882
R43904 PAD.n8980 PAD.n8913 0.0380882
R43905 PAD.n8976 PAD.n8913 0.0380882
R43906 PAD.n8976 PAD.n8972 0.0380882
R43907 PAD.n8972 PAD.n8971 0.0380882
R43908 PAD.n8971 PAD.n8918 0.0380882
R43909 PAD.n8967 PAD.n8918 0.0380882
R43910 PAD.n8967 PAD.n8963 0.0380882
R43911 PAD.n8963 PAD.n8962 0.0380882
R43912 PAD.n8962 PAD.n8923 0.0380882
R43913 PAD.n8958 PAD.n8923 0.0380882
R43914 PAD.n8958 PAD.n8954 0.0380882
R43915 PAD.n8954 PAD.n8953 0.0380882
R43916 PAD.n8953 PAD.n8928 0.0380882
R43917 PAD.n8949 PAD.n8928 0.0380882
R43918 PAD.n8949 PAD.n8945 0.0380882
R43919 PAD.n8945 PAD.n8944 0.0380882
R43920 PAD.n8944 PAD.n8933 0.0380882
R43921 PAD.n8940 PAD.n8933 0.0380882
R43922 PAD.n8940 PAD.n2880 0.0380882
R43923 PAD.n9136 PAD.n2880 0.0380882
R43924 PAD.n9136 PAD.n2877 0.0380882
R43925 PAD.n9120 PAD.n8837 0.0380882
R43926 PAD.n9114 PAD.n8837 0.0380882
R43927 PAD.n9114 PAD.n9113 0.0380882
R43928 PAD.n9113 PAD.n9112 0.0380882
R43929 PAD.n9112 PAD.n8842 0.0380882
R43930 PAD.n9105 PAD.n8842 0.0380882
R43931 PAD.n9105 PAD.n9104 0.0380882
R43932 PAD.n9104 PAD.n9103 0.0380882
R43933 PAD.n9103 PAD.n8847 0.0380882
R43934 PAD.n9096 PAD.n8847 0.0380882
R43935 PAD.n9096 PAD.n9095 0.0380882
R43936 PAD.n9095 PAD.n9094 0.0380882
R43937 PAD.n9094 PAD.n8852 0.0380882
R43938 PAD.n9087 PAD.n8852 0.0380882
R43939 PAD.n9087 PAD.n9086 0.0380882
R43940 PAD.n9086 PAD.n9085 0.0380882
R43941 PAD.n9085 PAD.n8857 0.0380882
R43942 PAD.n9078 PAD.n8857 0.0380882
R43943 PAD.n9078 PAD.n9077 0.0380882
R43944 PAD.n9077 PAD.n9076 0.0380882
R43945 PAD.n9076 PAD.n8862 0.0380882
R43946 PAD.n9069 PAD.n8862 0.0380882
R43947 PAD.n9069 PAD.n9068 0.0380882
R43948 PAD.n9068 PAD.n9067 0.0380882
R43949 PAD.n9067 PAD.n8867 0.0380882
R43950 PAD.n9060 PAD.n8867 0.0380882
R43951 PAD.n9060 PAD.n9059 0.0380882
R43952 PAD.n9059 PAD.n9058 0.0380882
R43953 PAD.n9058 PAD.n8872 0.0380882
R43954 PAD.n9051 PAD.n8872 0.0380882
R43955 PAD.n9051 PAD.n9050 0.0380882
R43956 PAD.n9050 PAD.n9049 0.0380882
R43957 PAD.n9049 PAD.n8877 0.0380882
R43958 PAD.n9042 PAD.n8877 0.0380882
R43959 PAD.n9042 PAD.n9041 0.0380882
R43960 PAD.n9041 PAD.n9040 0.0380882
R43961 PAD.n9040 PAD.n8882 0.0380882
R43962 PAD.n9033 PAD.n8882 0.0380882
R43963 PAD.n9033 PAD.n9032 0.0380882
R43964 PAD.n9032 PAD.n9031 0.0380882
R43965 PAD.n9031 PAD.n8887 0.0380882
R43966 PAD.n9024 PAD.n8887 0.0380882
R43967 PAD.n9024 PAD.n9023 0.0380882
R43968 PAD.n9023 PAD.n9022 0.0380882
R43969 PAD.n9022 PAD.n8892 0.0380882
R43970 PAD.n9015 PAD.n8892 0.0380882
R43971 PAD.n9015 PAD.n9014 0.0380882
R43972 PAD.n9014 PAD.n9013 0.0380882
R43973 PAD.n9013 PAD.n8897 0.0380882
R43974 PAD.n9006 PAD.n8897 0.0380882
R43975 PAD.n9006 PAD.n9005 0.0380882
R43976 PAD.n9005 PAD.n9004 0.0380882
R43977 PAD.n9004 PAD.n8902 0.0380882
R43978 PAD.n8997 PAD.n8902 0.0380882
R43979 PAD.n8997 PAD.n8996 0.0380882
R43980 PAD.n8996 PAD.n8995 0.0380882
R43981 PAD.n8995 PAD.n8907 0.0380882
R43982 PAD.n8988 PAD.n8907 0.0380882
R43983 PAD.n8988 PAD.n8987 0.0380882
R43984 PAD.n8987 PAD.n8986 0.0380882
R43985 PAD.n8986 PAD.n8912 0.0380882
R43986 PAD.n8979 PAD.n8912 0.0380882
R43987 PAD.n8979 PAD.n8978 0.0380882
R43988 PAD.n8978 PAD.n8977 0.0380882
R43989 PAD.n8977 PAD.n8917 0.0380882
R43990 PAD.n8970 PAD.n8917 0.0380882
R43991 PAD.n8970 PAD.n8969 0.0380882
R43992 PAD.n8969 PAD.n8968 0.0380882
R43993 PAD.n8968 PAD.n8922 0.0380882
R43994 PAD.n8961 PAD.n8922 0.0380882
R43995 PAD.n8961 PAD.n8960 0.0380882
R43996 PAD.n8960 PAD.n8959 0.0380882
R43997 PAD.n8959 PAD.n8927 0.0380882
R43998 PAD.n8952 PAD.n8927 0.0380882
R43999 PAD.n8952 PAD.n8951 0.0380882
R44000 PAD.n8951 PAD.n8950 0.0380882
R44001 PAD.n8950 PAD.n8932 0.0380882
R44002 PAD.n8943 PAD.n8932 0.0380882
R44003 PAD.n8943 PAD.n8942 0.0380882
R44004 PAD.n8942 PAD.n8941 0.0380882
R44005 PAD.n8941 PAD.n2881 0.0380882
R44006 PAD.n9135 PAD.n2881 0.0380882
R44007 PAD.n9135 PAD.n9134 0.0380882
R44008 PAD.n8818 PAD.n8529 0.0380882
R44009 PAD.n8814 PAD.n8529 0.0380882
R44010 PAD.n8814 PAD.n8811 0.0380882
R44011 PAD.n8811 PAD.n8807 0.0380882
R44012 PAD.n8807 PAD.n8531 0.0380882
R44013 PAD.n8803 PAD.n8531 0.0380882
R44014 PAD.n8803 PAD.n8799 0.0380882
R44015 PAD.n8799 PAD.n8795 0.0380882
R44016 PAD.n8795 PAD.n8533 0.0380882
R44017 PAD.n8791 PAD.n8533 0.0380882
R44018 PAD.n8791 PAD.n8787 0.0380882
R44019 PAD.n8787 PAD.n8783 0.0380882
R44020 PAD.n8783 PAD.n8535 0.0380882
R44021 PAD.n8779 PAD.n8535 0.0380882
R44022 PAD.n8779 PAD.n8775 0.0380882
R44023 PAD.n8775 PAD.n8771 0.0380882
R44024 PAD.n8771 PAD.n8537 0.0380882
R44025 PAD.n8767 PAD.n8537 0.0380882
R44026 PAD.n8767 PAD.n8763 0.0380882
R44027 PAD.n8763 PAD.n8759 0.0380882
R44028 PAD.n8759 PAD.n8539 0.0380882
R44029 PAD.n8755 PAD.n8539 0.0380882
R44030 PAD.n8755 PAD.n8751 0.0380882
R44031 PAD.n8751 PAD.n8747 0.0380882
R44032 PAD.n8747 PAD.n8541 0.0380882
R44033 PAD.n8743 PAD.n8541 0.0380882
R44034 PAD.n8743 PAD.n8739 0.0380882
R44035 PAD.n8739 PAD.n8735 0.0380882
R44036 PAD.n8735 PAD.n8543 0.0380882
R44037 PAD.n8731 PAD.n8543 0.0380882
R44038 PAD.n8731 PAD.n8727 0.0380882
R44039 PAD.n8727 PAD.n8723 0.0380882
R44040 PAD.n8723 PAD.n8545 0.0380882
R44041 PAD.n8719 PAD.n8545 0.0380882
R44042 PAD.n8719 PAD.n8715 0.0380882
R44043 PAD.n8715 PAD.n8711 0.0380882
R44044 PAD.n8711 PAD.n8547 0.0380882
R44045 PAD.n8707 PAD.n8547 0.0380882
R44046 PAD.n8707 PAD.n8703 0.0380882
R44047 PAD.n8703 PAD.n8699 0.0380882
R44048 PAD.n8699 PAD.n8549 0.0380882
R44049 PAD.n8695 PAD.n8549 0.0380882
R44050 PAD.n8695 PAD.n8691 0.0380882
R44051 PAD.n8691 PAD.n8687 0.0380882
R44052 PAD.n8687 PAD.n8551 0.0380882
R44053 PAD.n8683 PAD.n8551 0.0380882
R44054 PAD.n8683 PAD.n8679 0.0380882
R44055 PAD.n8679 PAD.n8675 0.0380882
R44056 PAD.n8675 PAD.n8553 0.0380882
R44057 PAD.n8671 PAD.n8553 0.0380882
R44058 PAD.n8671 PAD.n8667 0.0380882
R44059 PAD.n8667 PAD.n8663 0.0380882
R44060 PAD.n8663 PAD.n8555 0.0380882
R44061 PAD.n8659 PAD.n8555 0.0380882
R44062 PAD.n8659 PAD.n8655 0.0380882
R44063 PAD.n8655 PAD.n8651 0.0380882
R44064 PAD.n8651 PAD.n8557 0.0380882
R44065 PAD.n8647 PAD.n8557 0.0380882
R44066 PAD.n8647 PAD.n8643 0.0380882
R44067 PAD.n8643 PAD.n8639 0.0380882
R44068 PAD.n8639 PAD.n8559 0.0380882
R44069 PAD.n8635 PAD.n8559 0.0380882
R44070 PAD.n8635 PAD.n8631 0.0380882
R44071 PAD.n8631 PAD.n8627 0.0380882
R44072 PAD.n8627 PAD.n8561 0.0380882
R44073 PAD.n8623 PAD.n8561 0.0380882
R44074 PAD.n8623 PAD.n8619 0.0380882
R44075 PAD.n8619 PAD.n8615 0.0380882
R44076 PAD.n8615 PAD.n8563 0.0380882
R44077 PAD.n8611 PAD.n8563 0.0380882
R44078 PAD.n8611 PAD.n8607 0.0380882
R44079 PAD.n8607 PAD.n8603 0.0380882
R44080 PAD.n8603 PAD.n8565 0.0380882
R44081 PAD.n8599 PAD.n8565 0.0380882
R44082 PAD.n8599 PAD.n8595 0.0380882
R44083 PAD.n8595 PAD.n8591 0.0380882
R44084 PAD.n8591 PAD.n8567 0.0380882
R44085 PAD.n8587 PAD.n8567 0.0380882
R44086 PAD.n8587 PAD.n8583 0.0380882
R44087 PAD.n8583 PAD.n8579 0.0380882
R44088 PAD.n8579 PAD.n8569 0.0380882
R44089 PAD.n8575 PAD.n8569 0.0380882
R44090 PAD.n8575 PAD.n8571 0.0380882
R44091 PAD.n8817 PAD.n8816 0.0380882
R44092 PAD.n8816 PAD.n8815 0.0380882
R44093 PAD.n8815 PAD.n8530 0.0380882
R44094 PAD.n8806 PAD.n8530 0.0380882
R44095 PAD.n8806 PAD.n8805 0.0380882
R44096 PAD.n8805 PAD.n8804 0.0380882
R44097 PAD.n8804 PAD.n8532 0.0380882
R44098 PAD.n8794 PAD.n8532 0.0380882
R44099 PAD.n8794 PAD.n8793 0.0380882
R44100 PAD.n8793 PAD.n8792 0.0380882
R44101 PAD.n8792 PAD.n8534 0.0380882
R44102 PAD.n8782 PAD.n8534 0.0380882
R44103 PAD.n8782 PAD.n8781 0.0380882
R44104 PAD.n8781 PAD.n8780 0.0380882
R44105 PAD.n8780 PAD.n8536 0.0380882
R44106 PAD.n8770 PAD.n8536 0.0380882
R44107 PAD.n8770 PAD.n8769 0.0380882
R44108 PAD.n8769 PAD.n8768 0.0380882
R44109 PAD.n8768 PAD.n8538 0.0380882
R44110 PAD.n8758 PAD.n8538 0.0380882
R44111 PAD.n8758 PAD.n8757 0.0380882
R44112 PAD.n8757 PAD.n8756 0.0380882
R44113 PAD.n8756 PAD.n8540 0.0380882
R44114 PAD.n8746 PAD.n8540 0.0380882
R44115 PAD.n8746 PAD.n8745 0.0380882
R44116 PAD.n8745 PAD.n8744 0.0380882
R44117 PAD.n8744 PAD.n8542 0.0380882
R44118 PAD.n8734 PAD.n8542 0.0380882
R44119 PAD.n8734 PAD.n8733 0.0380882
R44120 PAD.n8733 PAD.n8732 0.0380882
R44121 PAD.n8732 PAD.n8544 0.0380882
R44122 PAD.n8722 PAD.n8544 0.0380882
R44123 PAD.n8722 PAD.n8721 0.0380882
R44124 PAD.n8721 PAD.n8720 0.0380882
R44125 PAD.n8720 PAD.n8546 0.0380882
R44126 PAD.n8710 PAD.n8546 0.0380882
R44127 PAD.n8710 PAD.n8709 0.0380882
R44128 PAD.n8709 PAD.n8708 0.0380882
R44129 PAD.n8708 PAD.n8548 0.0380882
R44130 PAD.n8698 PAD.n8548 0.0380882
R44131 PAD.n8698 PAD.n8697 0.0380882
R44132 PAD.n8697 PAD.n8696 0.0380882
R44133 PAD.n8696 PAD.n8550 0.0380882
R44134 PAD.n8686 PAD.n8550 0.0380882
R44135 PAD.n8686 PAD.n8685 0.0380882
R44136 PAD.n8685 PAD.n8684 0.0380882
R44137 PAD.n8684 PAD.n8552 0.0380882
R44138 PAD.n8674 PAD.n8552 0.0380882
R44139 PAD.n8674 PAD.n8673 0.0380882
R44140 PAD.n8673 PAD.n8672 0.0380882
R44141 PAD.n8672 PAD.n8554 0.0380882
R44142 PAD.n8662 PAD.n8554 0.0380882
R44143 PAD.n8662 PAD.n8661 0.0380882
R44144 PAD.n8661 PAD.n8660 0.0380882
R44145 PAD.n8660 PAD.n8556 0.0380882
R44146 PAD.n8650 PAD.n8556 0.0380882
R44147 PAD.n8650 PAD.n8649 0.0380882
R44148 PAD.n8649 PAD.n8648 0.0380882
R44149 PAD.n8648 PAD.n8558 0.0380882
R44150 PAD.n8638 PAD.n8558 0.0380882
R44151 PAD.n8638 PAD.n8637 0.0380882
R44152 PAD.n8637 PAD.n8636 0.0380882
R44153 PAD.n8636 PAD.n8560 0.0380882
R44154 PAD.n8626 PAD.n8560 0.0380882
R44155 PAD.n8626 PAD.n8625 0.0380882
R44156 PAD.n8625 PAD.n8624 0.0380882
R44157 PAD.n8624 PAD.n8562 0.0380882
R44158 PAD.n8614 PAD.n8562 0.0380882
R44159 PAD.n8614 PAD.n8613 0.0380882
R44160 PAD.n8613 PAD.n8612 0.0380882
R44161 PAD.n8612 PAD.n8564 0.0380882
R44162 PAD.n8602 PAD.n8564 0.0380882
R44163 PAD.n8602 PAD.n8601 0.0380882
R44164 PAD.n8601 PAD.n8600 0.0380882
R44165 PAD.n8600 PAD.n8566 0.0380882
R44166 PAD.n8590 PAD.n8566 0.0380882
R44167 PAD.n8590 PAD.n8589 0.0380882
R44168 PAD.n8589 PAD.n8588 0.0380882
R44169 PAD.n8588 PAD.n8568 0.0380882
R44170 PAD.n8578 PAD.n8568 0.0380882
R44171 PAD.n8578 PAD.n8577 0.0380882
R44172 PAD.n8577 PAD.n8576 0.0380882
R44173 PAD.n8576 PAD.n2898 0.0380882
R44174 PAD.n3041 PAD.n3040 0.0380882
R44175 PAD.n3045 PAD.n3040 0.0380882
R44176 PAD.n3049 PAD.n3045 0.0380882
R44177 PAD.n3053 PAD.n3049 0.0380882
R44178 PAD.n3053 PAD.n3036 0.0380882
R44179 PAD.n3057 PAD.n3036 0.0380882
R44180 PAD.n3061 PAD.n3057 0.0380882
R44181 PAD.n3065 PAD.n3061 0.0380882
R44182 PAD.n3065 PAD.n3034 0.0380882
R44183 PAD.n3069 PAD.n3034 0.0380882
R44184 PAD.n3073 PAD.n3069 0.0380882
R44185 PAD.n3077 PAD.n3073 0.0380882
R44186 PAD.n3077 PAD.n3032 0.0380882
R44187 PAD.n3081 PAD.n3032 0.0380882
R44188 PAD.n3085 PAD.n3081 0.0380882
R44189 PAD.n3089 PAD.n3085 0.0380882
R44190 PAD.n3089 PAD.n3030 0.0380882
R44191 PAD.n3093 PAD.n3030 0.0380882
R44192 PAD.n3097 PAD.n3093 0.0380882
R44193 PAD.n3101 PAD.n3097 0.0380882
R44194 PAD.n3101 PAD.n3028 0.0380882
R44195 PAD.n3105 PAD.n3028 0.0380882
R44196 PAD.n3109 PAD.n3105 0.0380882
R44197 PAD.n3113 PAD.n3109 0.0380882
R44198 PAD.n3113 PAD.n3026 0.0380882
R44199 PAD.n3117 PAD.n3026 0.0380882
R44200 PAD.n3121 PAD.n3117 0.0380882
R44201 PAD.n3125 PAD.n3121 0.0380882
R44202 PAD.n3125 PAD.n3024 0.0380882
R44203 PAD.n3129 PAD.n3024 0.0380882
R44204 PAD.n3133 PAD.n3129 0.0380882
R44205 PAD.n3137 PAD.n3133 0.0380882
R44206 PAD.n3137 PAD.n3022 0.0380882
R44207 PAD.n3141 PAD.n3022 0.0380882
R44208 PAD.n3145 PAD.n3141 0.0380882
R44209 PAD.n3149 PAD.n3145 0.0380882
R44210 PAD.n3149 PAD.n3020 0.0380882
R44211 PAD.n3153 PAD.n3020 0.0380882
R44212 PAD.n3157 PAD.n3153 0.0380882
R44213 PAD.n3161 PAD.n3157 0.0380882
R44214 PAD.n3161 PAD.n3018 0.0380882
R44215 PAD.n3165 PAD.n3018 0.0380882
R44216 PAD.n3169 PAD.n3165 0.0380882
R44217 PAD.n3173 PAD.n3169 0.0380882
R44218 PAD.n3173 PAD.n3016 0.0380882
R44219 PAD.n3177 PAD.n3016 0.0380882
R44220 PAD.n3181 PAD.n3177 0.0380882
R44221 PAD.n3185 PAD.n3181 0.0380882
R44222 PAD.n3185 PAD.n3014 0.0380882
R44223 PAD.n3189 PAD.n3014 0.0380882
R44224 PAD.n3193 PAD.n3189 0.0380882
R44225 PAD.n3197 PAD.n3193 0.0380882
R44226 PAD.n3197 PAD.n3012 0.0380882
R44227 PAD.n3201 PAD.n3012 0.0380882
R44228 PAD.n3205 PAD.n3201 0.0380882
R44229 PAD.n3209 PAD.n3205 0.0380882
R44230 PAD.n3209 PAD.n3010 0.0380882
R44231 PAD.n3213 PAD.n3010 0.0380882
R44232 PAD.n3217 PAD.n3213 0.0380882
R44233 PAD.n3221 PAD.n3217 0.0380882
R44234 PAD.n3221 PAD.n3008 0.0380882
R44235 PAD.n3225 PAD.n3008 0.0380882
R44236 PAD.n3229 PAD.n3225 0.0380882
R44237 PAD.n3233 PAD.n3229 0.0380882
R44238 PAD.n3233 PAD.n3006 0.0380882
R44239 PAD.n3237 PAD.n3006 0.0380882
R44240 PAD.n3241 PAD.n3237 0.0380882
R44241 PAD.n3245 PAD.n3241 0.0380882
R44242 PAD.n3245 PAD.n3004 0.0380882
R44243 PAD.n3249 PAD.n3004 0.0380882
R44244 PAD.n3253 PAD.n3249 0.0380882
R44245 PAD.n3257 PAD.n3253 0.0380882
R44246 PAD.n3257 PAD.n3002 0.0380882
R44247 PAD.n3261 PAD.n3002 0.0380882
R44248 PAD.n3265 PAD.n3261 0.0380882
R44249 PAD.n3269 PAD.n3265 0.0380882
R44250 PAD.n3269 PAD.n3000 0.0380882
R44251 PAD.n3273 PAD.n3000 0.0380882
R44252 PAD.n3277 PAD.n3273 0.0380882
R44253 PAD.n3281 PAD.n3277 0.0380882
R44254 PAD.n3281 PAD.n2998 0.0380882
R44255 PAD.n8513 PAD.n2998 0.0380882
R44256 PAD.n8513 PAD.n2995 0.0380882
R44257 PAD.n3043 PAD.n3042 0.0380882
R44258 PAD.n3044 PAD.n3043 0.0380882
R44259 PAD.n3044 PAD.n3037 0.0380882
R44260 PAD.n3054 PAD.n3037 0.0380882
R44261 PAD.n3055 PAD.n3054 0.0380882
R44262 PAD.n3056 PAD.n3055 0.0380882
R44263 PAD.n3056 PAD.n3035 0.0380882
R44264 PAD.n3066 PAD.n3035 0.0380882
R44265 PAD.n3067 PAD.n3066 0.0380882
R44266 PAD.n3068 PAD.n3067 0.0380882
R44267 PAD.n3068 PAD.n3033 0.0380882
R44268 PAD.n3078 PAD.n3033 0.0380882
R44269 PAD.n3079 PAD.n3078 0.0380882
R44270 PAD.n3080 PAD.n3079 0.0380882
R44271 PAD.n3080 PAD.n3031 0.0380882
R44272 PAD.n3090 PAD.n3031 0.0380882
R44273 PAD.n3091 PAD.n3090 0.0380882
R44274 PAD.n3092 PAD.n3091 0.0380882
R44275 PAD.n3092 PAD.n3029 0.0380882
R44276 PAD.n3102 PAD.n3029 0.0380882
R44277 PAD.n3103 PAD.n3102 0.0380882
R44278 PAD.n3104 PAD.n3103 0.0380882
R44279 PAD.n3104 PAD.n3027 0.0380882
R44280 PAD.n3114 PAD.n3027 0.0380882
R44281 PAD.n3115 PAD.n3114 0.0380882
R44282 PAD.n3116 PAD.n3115 0.0380882
R44283 PAD.n3116 PAD.n3025 0.0380882
R44284 PAD.n3126 PAD.n3025 0.0380882
R44285 PAD.n3127 PAD.n3126 0.0380882
R44286 PAD.n3128 PAD.n3127 0.0380882
R44287 PAD.n3128 PAD.n3023 0.0380882
R44288 PAD.n3138 PAD.n3023 0.0380882
R44289 PAD.n3139 PAD.n3138 0.0380882
R44290 PAD.n3140 PAD.n3139 0.0380882
R44291 PAD.n3140 PAD.n3021 0.0380882
R44292 PAD.n3150 PAD.n3021 0.0380882
R44293 PAD.n3151 PAD.n3150 0.0380882
R44294 PAD.n3152 PAD.n3151 0.0380882
R44295 PAD.n3152 PAD.n3019 0.0380882
R44296 PAD.n3162 PAD.n3019 0.0380882
R44297 PAD.n3163 PAD.n3162 0.0380882
R44298 PAD.n3164 PAD.n3163 0.0380882
R44299 PAD.n3164 PAD.n3017 0.0380882
R44300 PAD.n3174 PAD.n3017 0.0380882
R44301 PAD.n3175 PAD.n3174 0.0380882
R44302 PAD.n3176 PAD.n3175 0.0380882
R44303 PAD.n3176 PAD.n3015 0.0380882
R44304 PAD.n3186 PAD.n3015 0.0380882
R44305 PAD.n3187 PAD.n3186 0.0380882
R44306 PAD.n3188 PAD.n3187 0.0380882
R44307 PAD.n3188 PAD.n3013 0.0380882
R44308 PAD.n3198 PAD.n3013 0.0380882
R44309 PAD.n3199 PAD.n3198 0.0380882
R44310 PAD.n3200 PAD.n3199 0.0380882
R44311 PAD.n3200 PAD.n3011 0.0380882
R44312 PAD.n3210 PAD.n3011 0.0380882
R44313 PAD.n3211 PAD.n3210 0.0380882
R44314 PAD.n3212 PAD.n3211 0.0380882
R44315 PAD.n3212 PAD.n3009 0.0380882
R44316 PAD.n3222 PAD.n3009 0.0380882
R44317 PAD.n3223 PAD.n3222 0.0380882
R44318 PAD.n3224 PAD.n3223 0.0380882
R44319 PAD.n3224 PAD.n3007 0.0380882
R44320 PAD.n3234 PAD.n3007 0.0380882
R44321 PAD.n3235 PAD.n3234 0.0380882
R44322 PAD.n3236 PAD.n3235 0.0380882
R44323 PAD.n3236 PAD.n3005 0.0380882
R44324 PAD.n3246 PAD.n3005 0.0380882
R44325 PAD.n3247 PAD.n3246 0.0380882
R44326 PAD.n3248 PAD.n3247 0.0380882
R44327 PAD.n3248 PAD.n3003 0.0380882
R44328 PAD.n3258 PAD.n3003 0.0380882
R44329 PAD.n3259 PAD.n3258 0.0380882
R44330 PAD.n3260 PAD.n3259 0.0380882
R44331 PAD.n3260 PAD.n3001 0.0380882
R44332 PAD.n3270 PAD.n3001 0.0380882
R44333 PAD.n3271 PAD.n3270 0.0380882
R44334 PAD.n3272 PAD.n3271 0.0380882
R44335 PAD.n3272 PAD.n2999 0.0380882
R44336 PAD.n3282 PAD.n2999 0.0380882
R44337 PAD.n3283 PAD.n3282 0.0380882
R44338 PAD.n8512 PAD.n3283 0.0380882
R44339 PAD.n8512 PAD.n8511 0.0380882
R44340 PAD.n3386 PAD.n3385 0.0380882
R44341 PAD.n3390 PAD.n3385 0.0380882
R44342 PAD.n3394 PAD.n3390 0.0380882
R44343 PAD.n3398 PAD.n3394 0.0380882
R44344 PAD.n3398 PAD.n3381 0.0380882
R44345 PAD.n3402 PAD.n3381 0.0380882
R44346 PAD.n3406 PAD.n3402 0.0380882
R44347 PAD.n3410 PAD.n3406 0.0380882
R44348 PAD.n3410 PAD.n3379 0.0380882
R44349 PAD.n3414 PAD.n3379 0.0380882
R44350 PAD.n3418 PAD.n3414 0.0380882
R44351 PAD.n3422 PAD.n3418 0.0380882
R44352 PAD.n3422 PAD.n3377 0.0380882
R44353 PAD.n3426 PAD.n3377 0.0380882
R44354 PAD.n3430 PAD.n3426 0.0380882
R44355 PAD.n3434 PAD.n3430 0.0380882
R44356 PAD.n3434 PAD.n3375 0.0380882
R44357 PAD.n3438 PAD.n3375 0.0380882
R44358 PAD.n3442 PAD.n3438 0.0380882
R44359 PAD.n3446 PAD.n3442 0.0380882
R44360 PAD.n3446 PAD.n3373 0.0380882
R44361 PAD.n3450 PAD.n3373 0.0380882
R44362 PAD.n3454 PAD.n3450 0.0380882
R44363 PAD.n3458 PAD.n3454 0.0380882
R44364 PAD.n3458 PAD.n3371 0.0380882
R44365 PAD.n3462 PAD.n3371 0.0380882
R44366 PAD.n3466 PAD.n3462 0.0380882
R44367 PAD.n3470 PAD.n3466 0.0380882
R44368 PAD.n3470 PAD.n3369 0.0380882
R44369 PAD.n3474 PAD.n3369 0.0380882
R44370 PAD.n3478 PAD.n3474 0.0380882
R44371 PAD.n3482 PAD.n3478 0.0380882
R44372 PAD.n3482 PAD.n3367 0.0380882
R44373 PAD.n3486 PAD.n3367 0.0380882
R44374 PAD.n3490 PAD.n3486 0.0380882
R44375 PAD.n3494 PAD.n3490 0.0380882
R44376 PAD.n3494 PAD.n3365 0.0380882
R44377 PAD.n3498 PAD.n3365 0.0380882
R44378 PAD.n3502 PAD.n3498 0.0380882
R44379 PAD.n3506 PAD.n3502 0.0380882
R44380 PAD.n3506 PAD.n3363 0.0380882
R44381 PAD.n3510 PAD.n3363 0.0380882
R44382 PAD.n3514 PAD.n3510 0.0380882
R44383 PAD.n3518 PAD.n3514 0.0380882
R44384 PAD.n3518 PAD.n3361 0.0380882
R44385 PAD.n3522 PAD.n3361 0.0380882
R44386 PAD.n3526 PAD.n3522 0.0380882
R44387 PAD.n3530 PAD.n3526 0.0380882
R44388 PAD.n3530 PAD.n3359 0.0380882
R44389 PAD.n3534 PAD.n3359 0.0380882
R44390 PAD.n3538 PAD.n3534 0.0380882
R44391 PAD.n3542 PAD.n3538 0.0380882
R44392 PAD.n3542 PAD.n3357 0.0380882
R44393 PAD.n3546 PAD.n3357 0.0380882
R44394 PAD.n3550 PAD.n3546 0.0380882
R44395 PAD.n3554 PAD.n3550 0.0380882
R44396 PAD.n3554 PAD.n3355 0.0380882
R44397 PAD.n3558 PAD.n3355 0.0380882
R44398 PAD.n3562 PAD.n3558 0.0380882
R44399 PAD.n3566 PAD.n3562 0.0380882
R44400 PAD.n3566 PAD.n3353 0.0380882
R44401 PAD.n3570 PAD.n3353 0.0380882
R44402 PAD.n3574 PAD.n3570 0.0380882
R44403 PAD.n3578 PAD.n3574 0.0380882
R44404 PAD.n3578 PAD.n3351 0.0380882
R44405 PAD.n3582 PAD.n3351 0.0380882
R44406 PAD.n3586 PAD.n3582 0.0380882
R44407 PAD.n3590 PAD.n3586 0.0380882
R44408 PAD.n3590 PAD.n3349 0.0380882
R44409 PAD.n3594 PAD.n3349 0.0380882
R44410 PAD.n3598 PAD.n3594 0.0380882
R44411 PAD.n3602 PAD.n3598 0.0380882
R44412 PAD.n3602 PAD.n3347 0.0380882
R44413 PAD.n3606 PAD.n3347 0.0380882
R44414 PAD.n3610 PAD.n3606 0.0380882
R44415 PAD.n3614 PAD.n3610 0.0380882
R44416 PAD.n3614 PAD.n3345 0.0380882
R44417 PAD.n3618 PAD.n3345 0.0380882
R44418 PAD.n3622 PAD.n3618 0.0380882
R44419 PAD.n3626 PAD.n3622 0.0380882
R44420 PAD.n3626 PAD.n3343 0.0380882
R44421 PAD.n8488 PAD.n3343 0.0380882
R44422 PAD.n8488 PAD.n3340 0.0380882
R44423 PAD.n3388 PAD.n3387 0.0380882
R44424 PAD.n3389 PAD.n3388 0.0380882
R44425 PAD.n3389 PAD.n3382 0.0380882
R44426 PAD.n3399 PAD.n3382 0.0380882
R44427 PAD.n3400 PAD.n3399 0.0380882
R44428 PAD.n3401 PAD.n3400 0.0380882
R44429 PAD.n3401 PAD.n3380 0.0380882
R44430 PAD.n3411 PAD.n3380 0.0380882
R44431 PAD.n3412 PAD.n3411 0.0380882
R44432 PAD.n3413 PAD.n3412 0.0380882
R44433 PAD.n3413 PAD.n3378 0.0380882
R44434 PAD.n3423 PAD.n3378 0.0380882
R44435 PAD.n3424 PAD.n3423 0.0380882
R44436 PAD.n3425 PAD.n3424 0.0380882
R44437 PAD.n3425 PAD.n3376 0.0380882
R44438 PAD.n3435 PAD.n3376 0.0380882
R44439 PAD.n3436 PAD.n3435 0.0380882
R44440 PAD.n3437 PAD.n3436 0.0380882
R44441 PAD.n3437 PAD.n3374 0.0380882
R44442 PAD.n3447 PAD.n3374 0.0380882
R44443 PAD.n3448 PAD.n3447 0.0380882
R44444 PAD.n3449 PAD.n3448 0.0380882
R44445 PAD.n3449 PAD.n3372 0.0380882
R44446 PAD.n3459 PAD.n3372 0.0380882
R44447 PAD.n3460 PAD.n3459 0.0380882
R44448 PAD.n3461 PAD.n3460 0.0380882
R44449 PAD.n3461 PAD.n3370 0.0380882
R44450 PAD.n3471 PAD.n3370 0.0380882
R44451 PAD.n3472 PAD.n3471 0.0380882
R44452 PAD.n3473 PAD.n3472 0.0380882
R44453 PAD.n3473 PAD.n3368 0.0380882
R44454 PAD.n3483 PAD.n3368 0.0380882
R44455 PAD.n3484 PAD.n3483 0.0380882
R44456 PAD.n3485 PAD.n3484 0.0380882
R44457 PAD.n3485 PAD.n3366 0.0380882
R44458 PAD.n3495 PAD.n3366 0.0380882
R44459 PAD.n3496 PAD.n3495 0.0380882
R44460 PAD.n3497 PAD.n3496 0.0380882
R44461 PAD.n3497 PAD.n3364 0.0380882
R44462 PAD.n3507 PAD.n3364 0.0380882
R44463 PAD.n3508 PAD.n3507 0.0380882
R44464 PAD.n3509 PAD.n3508 0.0380882
R44465 PAD.n3509 PAD.n3362 0.0380882
R44466 PAD.n3519 PAD.n3362 0.0380882
R44467 PAD.n3520 PAD.n3519 0.0380882
R44468 PAD.n3521 PAD.n3520 0.0380882
R44469 PAD.n3521 PAD.n3360 0.0380882
R44470 PAD.n3531 PAD.n3360 0.0380882
R44471 PAD.n3532 PAD.n3531 0.0380882
R44472 PAD.n3533 PAD.n3532 0.0380882
R44473 PAD.n3533 PAD.n3358 0.0380882
R44474 PAD.n3543 PAD.n3358 0.0380882
R44475 PAD.n3544 PAD.n3543 0.0380882
R44476 PAD.n3545 PAD.n3544 0.0380882
R44477 PAD.n3545 PAD.n3356 0.0380882
R44478 PAD.n3555 PAD.n3356 0.0380882
R44479 PAD.n3556 PAD.n3555 0.0380882
R44480 PAD.n3557 PAD.n3556 0.0380882
R44481 PAD.n3557 PAD.n3354 0.0380882
R44482 PAD.n3567 PAD.n3354 0.0380882
R44483 PAD.n3568 PAD.n3567 0.0380882
R44484 PAD.n3569 PAD.n3568 0.0380882
R44485 PAD.n3569 PAD.n3352 0.0380882
R44486 PAD.n3579 PAD.n3352 0.0380882
R44487 PAD.n3580 PAD.n3579 0.0380882
R44488 PAD.n3581 PAD.n3580 0.0380882
R44489 PAD.n3581 PAD.n3350 0.0380882
R44490 PAD.n3591 PAD.n3350 0.0380882
R44491 PAD.n3592 PAD.n3591 0.0380882
R44492 PAD.n3593 PAD.n3592 0.0380882
R44493 PAD.n3593 PAD.n3348 0.0380882
R44494 PAD.n3603 PAD.n3348 0.0380882
R44495 PAD.n3604 PAD.n3603 0.0380882
R44496 PAD.n3605 PAD.n3604 0.0380882
R44497 PAD.n3605 PAD.n3346 0.0380882
R44498 PAD.n3615 PAD.n3346 0.0380882
R44499 PAD.n3616 PAD.n3615 0.0380882
R44500 PAD.n3617 PAD.n3616 0.0380882
R44501 PAD.n3617 PAD.n3344 0.0380882
R44502 PAD.n3627 PAD.n3344 0.0380882
R44503 PAD.n3628 PAD.n3627 0.0380882
R44504 PAD.n8487 PAD.n3628 0.0380882
R44505 PAD.n8487 PAD.n8486 0.0380882
R44506 PAD.n3731 PAD.n3730 0.0380882
R44507 PAD.n3735 PAD.n3730 0.0380882
R44508 PAD.n3739 PAD.n3735 0.0380882
R44509 PAD.n3743 PAD.n3739 0.0380882
R44510 PAD.n3743 PAD.n3726 0.0380882
R44511 PAD.n3747 PAD.n3726 0.0380882
R44512 PAD.n3751 PAD.n3747 0.0380882
R44513 PAD.n3755 PAD.n3751 0.0380882
R44514 PAD.n3755 PAD.n3724 0.0380882
R44515 PAD.n3759 PAD.n3724 0.0380882
R44516 PAD.n3763 PAD.n3759 0.0380882
R44517 PAD.n3767 PAD.n3763 0.0380882
R44518 PAD.n3767 PAD.n3722 0.0380882
R44519 PAD.n3771 PAD.n3722 0.0380882
R44520 PAD.n3775 PAD.n3771 0.0380882
R44521 PAD.n3779 PAD.n3775 0.0380882
R44522 PAD.n3779 PAD.n3720 0.0380882
R44523 PAD.n3783 PAD.n3720 0.0380882
R44524 PAD.n3787 PAD.n3783 0.0380882
R44525 PAD.n3791 PAD.n3787 0.0380882
R44526 PAD.n3791 PAD.n3718 0.0380882
R44527 PAD.n3795 PAD.n3718 0.0380882
R44528 PAD.n3799 PAD.n3795 0.0380882
R44529 PAD.n3803 PAD.n3799 0.0380882
R44530 PAD.n3803 PAD.n3716 0.0380882
R44531 PAD.n3807 PAD.n3716 0.0380882
R44532 PAD.n3811 PAD.n3807 0.0380882
R44533 PAD.n3815 PAD.n3811 0.0380882
R44534 PAD.n3815 PAD.n3714 0.0380882
R44535 PAD.n3819 PAD.n3714 0.0380882
R44536 PAD.n3823 PAD.n3819 0.0380882
R44537 PAD.n3827 PAD.n3823 0.0380882
R44538 PAD.n3827 PAD.n3712 0.0380882
R44539 PAD.n3831 PAD.n3712 0.0380882
R44540 PAD.n3835 PAD.n3831 0.0380882
R44541 PAD.n3839 PAD.n3835 0.0380882
R44542 PAD.n3839 PAD.n3710 0.0380882
R44543 PAD.n3843 PAD.n3710 0.0380882
R44544 PAD.n3847 PAD.n3843 0.0380882
R44545 PAD.n3851 PAD.n3847 0.0380882
R44546 PAD.n3851 PAD.n3708 0.0380882
R44547 PAD.n3855 PAD.n3708 0.0380882
R44548 PAD.n3859 PAD.n3855 0.0380882
R44549 PAD.n3863 PAD.n3859 0.0380882
R44550 PAD.n3863 PAD.n3706 0.0380882
R44551 PAD.n3867 PAD.n3706 0.0380882
R44552 PAD.n3871 PAD.n3867 0.0380882
R44553 PAD.n3875 PAD.n3871 0.0380882
R44554 PAD.n3875 PAD.n3704 0.0380882
R44555 PAD.n3879 PAD.n3704 0.0380882
R44556 PAD.n3883 PAD.n3879 0.0380882
R44557 PAD.n3887 PAD.n3883 0.0380882
R44558 PAD.n3887 PAD.n3702 0.0380882
R44559 PAD.n3891 PAD.n3702 0.0380882
R44560 PAD.n3895 PAD.n3891 0.0380882
R44561 PAD.n3899 PAD.n3895 0.0380882
R44562 PAD.n3899 PAD.n3700 0.0380882
R44563 PAD.n3903 PAD.n3700 0.0380882
R44564 PAD.n3907 PAD.n3903 0.0380882
R44565 PAD.n3911 PAD.n3907 0.0380882
R44566 PAD.n3911 PAD.n3698 0.0380882
R44567 PAD.n3915 PAD.n3698 0.0380882
R44568 PAD.n3919 PAD.n3915 0.0380882
R44569 PAD.n3923 PAD.n3919 0.0380882
R44570 PAD.n3923 PAD.n3696 0.0380882
R44571 PAD.n3927 PAD.n3696 0.0380882
R44572 PAD.n3931 PAD.n3927 0.0380882
R44573 PAD.n3935 PAD.n3931 0.0380882
R44574 PAD.n3935 PAD.n3694 0.0380882
R44575 PAD.n3939 PAD.n3694 0.0380882
R44576 PAD.n3943 PAD.n3939 0.0380882
R44577 PAD.n3947 PAD.n3943 0.0380882
R44578 PAD.n3947 PAD.n3692 0.0380882
R44579 PAD.n3951 PAD.n3692 0.0380882
R44580 PAD.n3955 PAD.n3951 0.0380882
R44581 PAD.n3959 PAD.n3955 0.0380882
R44582 PAD.n3959 PAD.n3690 0.0380882
R44583 PAD.n3963 PAD.n3690 0.0380882
R44584 PAD.n3967 PAD.n3963 0.0380882
R44585 PAD.n3971 PAD.n3967 0.0380882
R44586 PAD.n3971 PAD.n3688 0.0380882
R44587 PAD.n8464 PAD.n3688 0.0380882
R44588 PAD.n8464 PAD.n3685 0.0380882
R44589 PAD.n3733 PAD.n3732 0.0380882
R44590 PAD.n3734 PAD.n3733 0.0380882
R44591 PAD.n3734 PAD.n3727 0.0380882
R44592 PAD.n3744 PAD.n3727 0.0380882
R44593 PAD.n3745 PAD.n3744 0.0380882
R44594 PAD.n3746 PAD.n3745 0.0380882
R44595 PAD.n3746 PAD.n3725 0.0380882
R44596 PAD.n3756 PAD.n3725 0.0380882
R44597 PAD.n3757 PAD.n3756 0.0380882
R44598 PAD.n3758 PAD.n3757 0.0380882
R44599 PAD.n3758 PAD.n3723 0.0380882
R44600 PAD.n3768 PAD.n3723 0.0380882
R44601 PAD.n3769 PAD.n3768 0.0380882
R44602 PAD.n3770 PAD.n3769 0.0380882
R44603 PAD.n3770 PAD.n3721 0.0380882
R44604 PAD.n3780 PAD.n3721 0.0380882
R44605 PAD.n3781 PAD.n3780 0.0380882
R44606 PAD.n3782 PAD.n3781 0.0380882
R44607 PAD.n3782 PAD.n3719 0.0380882
R44608 PAD.n3792 PAD.n3719 0.0380882
R44609 PAD.n3793 PAD.n3792 0.0380882
R44610 PAD.n3794 PAD.n3793 0.0380882
R44611 PAD.n3794 PAD.n3717 0.0380882
R44612 PAD.n3804 PAD.n3717 0.0380882
R44613 PAD.n3805 PAD.n3804 0.0380882
R44614 PAD.n3806 PAD.n3805 0.0380882
R44615 PAD.n3806 PAD.n3715 0.0380882
R44616 PAD.n3816 PAD.n3715 0.0380882
R44617 PAD.n3817 PAD.n3816 0.0380882
R44618 PAD.n3818 PAD.n3817 0.0380882
R44619 PAD.n3818 PAD.n3713 0.0380882
R44620 PAD.n3828 PAD.n3713 0.0380882
R44621 PAD.n3829 PAD.n3828 0.0380882
R44622 PAD.n3830 PAD.n3829 0.0380882
R44623 PAD.n3830 PAD.n3711 0.0380882
R44624 PAD.n3840 PAD.n3711 0.0380882
R44625 PAD.n3841 PAD.n3840 0.0380882
R44626 PAD.n3842 PAD.n3841 0.0380882
R44627 PAD.n3842 PAD.n3709 0.0380882
R44628 PAD.n3852 PAD.n3709 0.0380882
R44629 PAD.n3853 PAD.n3852 0.0380882
R44630 PAD.n3854 PAD.n3853 0.0380882
R44631 PAD.n3854 PAD.n3707 0.0380882
R44632 PAD.n3864 PAD.n3707 0.0380882
R44633 PAD.n3865 PAD.n3864 0.0380882
R44634 PAD.n3866 PAD.n3865 0.0380882
R44635 PAD.n3866 PAD.n3705 0.0380882
R44636 PAD.n3876 PAD.n3705 0.0380882
R44637 PAD.n3877 PAD.n3876 0.0380882
R44638 PAD.n3878 PAD.n3877 0.0380882
R44639 PAD.n3878 PAD.n3703 0.0380882
R44640 PAD.n3888 PAD.n3703 0.0380882
R44641 PAD.n3889 PAD.n3888 0.0380882
R44642 PAD.n3890 PAD.n3889 0.0380882
R44643 PAD.n3890 PAD.n3701 0.0380882
R44644 PAD.n3900 PAD.n3701 0.0380882
R44645 PAD.n3901 PAD.n3900 0.0380882
R44646 PAD.n3902 PAD.n3901 0.0380882
R44647 PAD.n3902 PAD.n3699 0.0380882
R44648 PAD.n3912 PAD.n3699 0.0380882
R44649 PAD.n3913 PAD.n3912 0.0380882
R44650 PAD.n3914 PAD.n3913 0.0380882
R44651 PAD.n3914 PAD.n3697 0.0380882
R44652 PAD.n3924 PAD.n3697 0.0380882
R44653 PAD.n3925 PAD.n3924 0.0380882
R44654 PAD.n3926 PAD.n3925 0.0380882
R44655 PAD.n3926 PAD.n3695 0.0380882
R44656 PAD.n3936 PAD.n3695 0.0380882
R44657 PAD.n3937 PAD.n3936 0.0380882
R44658 PAD.n3938 PAD.n3937 0.0380882
R44659 PAD.n3938 PAD.n3693 0.0380882
R44660 PAD.n3948 PAD.n3693 0.0380882
R44661 PAD.n3949 PAD.n3948 0.0380882
R44662 PAD.n3950 PAD.n3949 0.0380882
R44663 PAD.n3950 PAD.n3691 0.0380882
R44664 PAD.n3960 PAD.n3691 0.0380882
R44665 PAD.n3961 PAD.n3960 0.0380882
R44666 PAD.n3962 PAD.n3961 0.0380882
R44667 PAD.n3962 PAD.n3689 0.0380882
R44668 PAD.n3972 PAD.n3689 0.0380882
R44669 PAD.n3973 PAD.n3972 0.0380882
R44670 PAD.n8463 PAD.n3973 0.0380882
R44671 PAD.n8463 PAD.n8462 0.0380882
R44672 PAD.n4072 PAD.n4071 0.0380882
R44673 PAD.n4076 PAD.n4071 0.0380882
R44674 PAD.n4080 PAD.n4076 0.0380882
R44675 PAD.n4084 PAD.n4080 0.0380882
R44676 PAD.n4084 PAD.n4067 0.0380882
R44677 PAD.n4088 PAD.n4067 0.0380882
R44678 PAD.n4092 PAD.n4088 0.0380882
R44679 PAD.n4096 PAD.n4092 0.0380882
R44680 PAD.n4096 PAD.n4065 0.0380882
R44681 PAD.n4100 PAD.n4065 0.0380882
R44682 PAD.n4104 PAD.n4100 0.0380882
R44683 PAD.n4108 PAD.n4104 0.0380882
R44684 PAD.n4108 PAD.n4063 0.0380882
R44685 PAD.n4112 PAD.n4063 0.0380882
R44686 PAD.n4116 PAD.n4112 0.0380882
R44687 PAD.n4120 PAD.n4116 0.0380882
R44688 PAD.n4120 PAD.n4061 0.0380882
R44689 PAD.n4124 PAD.n4061 0.0380882
R44690 PAD.n4128 PAD.n4124 0.0380882
R44691 PAD.n4132 PAD.n4128 0.0380882
R44692 PAD.n4132 PAD.n4059 0.0380882
R44693 PAD.n4136 PAD.n4059 0.0380882
R44694 PAD.n4140 PAD.n4136 0.0380882
R44695 PAD.n4144 PAD.n4140 0.0380882
R44696 PAD.n4144 PAD.n4057 0.0380882
R44697 PAD.n4148 PAD.n4057 0.0380882
R44698 PAD.n4152 PAD.n4148 0.0380882
R44699 PAD.n4156 PAD.n4152 0.0380882
R44700 PAD.n4156 PAD.n4055 0.0380882
R44701 PAD.n4160 PAD.n4055 0.0380882
R44702 PAD.n4164 PAD.n4160 0.0380882
R44703 PAD.n4168 PAD.n4164 0.0380882
R44704 PAD.n4168 PAD.n4053 0.0380882
R44705 PAD.n4172 PAD.n4053 0.0380882
R44706 PAD.n4176 PAD.n4172 0.0380882
R44707 PAD.n4180 PAD.n4176 0.0380882
R44708 PAD.n4180 PAD.n4051 0.0380882
R44709 PAD.n4184 PAD.n4051 0.0380882
R44710 PAD.n4188 PAD.n4184 0.0380882
R44711 PAD.n4192 PAD.n4188 0.0380882
R44712 PAD.n4192 PAD.n4049 0.0380882
R44713 PAD.n4196 PAD.n4049 0.0380882
R44714 PAD.n4200 PAD.n4196 0.0380882
R44715 PAD.n4204 PAD.n4200 0.0380882
R44716 PAD.n4204 PAD.n4047 0.0380882
R44717 PAD.n4208 PAD.n4047 0.0380882
R44718 PAD.n4212 PAD.n4208 0.0380882
R44719 PAD.n4216 PAD.n4212 0.0380882
R44720 PAD.n4216 PAD.n4045 0.0380882
R44721 PAD.n4220 PAD.n4045 0.0380882
R44722 PAD.n4224 PAD.n4220 0.0380882
R44723 PAD.n4228 PAD.n4224 0.0380882
R44724 PAD.n4228 PAD.n4043 0.0380882
R44725 PAD.n4232 PAD.n4043 0.0380882
R44726 PAD.n4236 PAD.n4232 0.0380882
R44727 PAD.n4240 PAD.n4236 0.0380882
R44728 PAD.n4240 PAD.n4041 0.0380882
R44729 PAD.n4244 PAD.n4041 0.0380882
R44730 PAD.n4248 PAD.n4244 0.0380882
R44731 PAD.n4252 PAD.n4248 0.0380882
R44732 PAD.n4252 PAD.n4039 0.0380882
R44733 PAD.n4256 PAD.n4039 0.0380882
R44734 PAD.n4260 PAD.n4256 0.0380882
R44735 PAD.n4264 PAD.n4260 0.0380882
R44736 PAD.n4264 PAD.n4037 0.0380882
R44737 PAD.n4268 PAD.n4037 0.0380882
R44738 PAD.n4272 PAD.n4268 0.0380882
R44739 PAD.n4276 PAD.n4272 0.0380882
R44740 PAD.n4276 PAD.n4035 0.0380882
R44741 PAD.n4280 PAD.n4035 0.0380882
R44742 PAD.n4284 PAD.n4280 0.0380882
R44743 PAD.n4288 PAD.n4284 0.0380882
R44744 PAD.n4288 PAD.n4033 0.0380882
R44745 PAD.n4292 PAD.n4033 0.0380882
R44746 PAD.n4296 PAD.n4292 0.0380882
R44747 PAD.n4300 PAD.n4296 0.0380882
R44748 PAD.n4300 PAD.n4031 0.0380882
R44749 PAD.n4304 PAD.n4031 0.0380882
R44750 PAD.n4308 PAD.n4304 0.0380882
R44751 PAD.n4312 PAD.n4308 0.0380882
R44752 PAD.n4312 PAD.n4029 0.0380882
R44753 PAD.n8440 PAD.n4029 0.0380882
R44754 PAD.n8440 PAD.n4026 0.0380882
R44755 PAD.n4074 PAD.n4073 0.0380882
R44756 PAD.n4075 PAD.n4074 0.0380882
R44757 PAD.n4075 PAD.n4068 0.0380882
R44758 PAD.n4085 PAD.n4068 0.0380882
R44759 PAD.n4086 PAD.n4085 0.0380882
R44760 PAD.n4087 PAD.n4086 0.0380882
R44761 PAD.n4087 PAD.n4066 0.0380882
R44762 PAD.n4097 PAD.n4066 0.0380882
R44763 PAD.n4098 PAD.n4097 0.0380882
R44764 PAD.n4099 PAD.n4098 0.0380882
R44765 PAD.n4099 PAD.n4064 0.0380882
R44766 PAD.n4109 PAD.n4064 0.0380882
R44767 PAD.n4110 PAD.n4109 0.0380882
R44768 PAD.n4111 PAD.n4110 0.0380882
R44769 PAD.n4111 PAD.n4062 0.0380882
R44770 PAD.n4121 PAD.n4062 0.0380882
R44771 PAD.n4122 PAD.n4121 0.0380882
R44772 PAD.n4123 PAD.n4122 0.0380882
R44773 PAD.n4123 PAD.n4060 0.0380882
R44774 PAD.n4133 PAD.n4060 0.0380882
R44775 PAD.n4134 PAD.n4133 0.0380882
R44776 PAD.n4135 PAD.n4134 0.0380882
R44777 PAD.n4135 PAD.n4058 0.0380882
R44778 PAD.n4145 PAD.n4058 0.0380882
R44779 PAD.n4146 PAD.n4145 0.0380882
R44780 PAD.n4147 PAD.n4146 0.0380882
R44781 PAD.n4147 PAD.n4056 0.0380882
R44782 PAD.n4157 PAD.n4056 0.0380882
R44783 PAD.n4158 PAD.n4157 0.0380882
R44784 PAD.n4159 PAD.n4158 0.0380882
R44785 PAD.n4159 PAD.n4054 0.0380882
R44786 PAD.n4169 PAD.n4054 0.0380882
R44787 PAD.n4170 PAD.n4169 0.0380882
R44788 PAD.n4171 PAD.n4170 0.0380882
R44789 PAD.n4171 PAD.n4052 0.0380882
R44790 PAD.n4181 PAD.n4052 0.0380882
R44791 PAD.n4182 PAD.n4181 0.0380882
R44792 PAD.n4183 PAD.n4182 0.0380882
R44793 PAD.n4183 PAD.n4050 0.0380882
R44794 PAD.n4193 PAD.n4050 0.0380882
R44795 PAD.n4194 PAD.n4193 0.0380882
R44796 PAD.n4195 PAD.n4194 0.0380882
R44797 PAD.n4195 PAD.n4048 0.0380882
R44798 PAD.n4205 PAD.n4048 0.0380882
R44799 PAD.n4206 PAD.n4205 0.0380882
R44800 PAD.n4207 PAD.n4206 0.0380882
R44801 PAD.n4207 PAD.n4046 0.0380882
R44802 PAD.n4217 PAD.n4046 0.0380882
R44803 PAD.n4218 PAD.n4217 0.0380882
R44804 PAD.n4219 PAD.n4218 0.0380882
R44805 PAD.n4219 PAD.n4044 0.0380882
R44806 PAD.n4229 PAD.n4044 0.0380882
R44807 PAD.n4230 PAD.n4229 0.0380882
R44808 PAD.n4231 PAD.n4230 0.0380882
R44809 PAD.n4231 PAD.n4042 0.0380882
R44810 PAD.n4241 PAD.n4042 0.0380882
R44811 PAD.n4242 PAD.n4241 0.0380882
R44812 PAD.n4243 PAD.n4242 0.0380882
R44813 PAD.n4243 PAD.n4040 0.0380882
R44814 PAD.n4253 PAD.n4040 0.0380882
R44815 PAD.n4254 PAD.n4253 0.0380882
R44816 PAD.n4255 PAD.n4254 0.0380882
R44817 PAD.n4255 PAD.n4038 0.0380882
R44818 PAD.n4265 PAD.n4038 0.0380882
R44819 PAD.n4266 PAD.n4265 0.0380882
R44820 PAD.n4267 PAD.n4266 0.0380882
R44821 PAD.n4267 PAD.n4036 0.0380882
R44822 PAD.n4277 PAD.n4036 0.0380882
R44823 PAD.n4278 PAD.n4277 0.0380882
R44824 PAD.n4279 PAD.n4278 0.0380882
R44825 PAD.n4279 PAD.n4034 0.0380882
R44826 PAD.n4289 PAD.n4034 0.0380882
R44827 PAD.n4290 PAD.n4289 0.0380882
R44828 PAD.n4291 PAD.n4290 0.0380882
R44829 PAD.n4291 PAD.n4032 0.0380882
R44830 PAD.n4301 PAD.n4032 0.0380882
R44831 PAD.n4302 PAD.n4301 0.0380882
R44832 PAD.n4303 PAD.n4302 0.0380882
R44833 PAD.n4303 PAD.n4030 0.0380882
R44834 PAD.n4313 PAD.n4030 0.0380882
R44835 PAD.n4314 PAD.n4313 0.0380882
R44836 PAD.n8439 PAD.n4314 0.0380882
R44837 PAD.n8439 PAD.n8438 0.0380882
R44838 PAD.n4419 PAD.n4418 0.0380882
R44839 PAD.n4427 PAD.n4418 0.0380882
R44840 PAD.n4427 PAD.n4416 0.0380882
R44841 PAD.n4431 PAD.n4416 0.0380882
R44842 PAD.n4431 PAD.n4414 0.0380882
R44843 PAD.n4439 PAD.n4414 0.0380882
R44844 PAD.n4439 PAD.n4412 0.0380882
R44845 PAD.n4443 PAD.n4412 0.0380882
R44846 PAD.n4443 PAD.n4410 0.0380882
R44847 PAD.n4451 PAD.n4410 0.0380882
R44848 PAD.n4451 PAD.n4408 0.0380882
R44849 PAD.n4455 PAD.n4408 0.0380882
R44850 PAD.n4455 PAD.n4406 0.0380882
R44851 PAD.n4463 PAD.n4406 0.0380882
R44852 PAD.n4463 PAD.n4404 0.0380882
R44853 PAD.n4467 PAD.n4404 0.0380882
R44854 PAD.n4467 PAD.n4402 0.0380882
R44855 PAD.n4475 PAD.n4402 0.0380882
R44856 PAD.n4475 PAD.n4400 0.0380882
R44857 PAD.n4479 PAD.n4400 0.0380882
R44858 PAD.n4479 PAD.n4398 0.0380882
R44859 PAD.n4487 PAD.n4398 0.0380882
R44860 PAD.n4487 PAD.n4396 0.0380882
R44861 PAD.n4491 PAD.n4396 0.0380882
R44862 PAD.n4491 PAD.n4394 0.0380882
R44863 PAD.n4499 PAD.n4394 0.0380882
R44864 PAD.n4499 PAD.n4392 0.0380882
R44865 PAD.n4503 PAD.n4392 0.0380882
R44866 PAD.n4503 PAD.n4390 0.0380882
R44867 PAD.n4511 PAD.n4390 0.0380882
R44868 PAD.n4511 PAD.n4388 0.0380882
R44869 PAD.n4515 PAD.n4388 0.0380882
R44870 PAD.n4515 PAD.n4386 0.0380882
R44871 PAD.n4523 PAD.n4386 0.0380882
R44872 PAD.n4523 PAD.n4384 0.0380882
R44873 PAD.n4527 PAD.n4384 0.0380882
R44874 PAD.n4527 PAD.n4382 0.0380882
R44875 PAD.n4535 PAD.n4382 0.0380882
R44876 PAD.n4535 PAD.n4380 0.0380882
R44877 PAD.n4539 PAD.n4380 0.0380882
R44878 PAD.n4539 PAD.n4378 0.0380882
R44879 PAD.n4547 PAD.n4378 0.0380882
R44880 PAD.n4547 PAD.n4376 0.0380882
R44881 PAD.n4551 PAD.n4376 0.0380882
R44882 PAD.n4551 PAD.n4374 0.0380882
R44883 PAD.n4559 PAD.n4374 0.0380882
R44884 PAD.n4559 PAD.n4372 0.0380882
R44885 PAD.n4563 PAD.n4372 0.0380882
R44886 PAD.n4563 PAD.n4370 0.0380882
R44887 PAD.n4571 PAD.n4370 0.0380882
R44888 PAD.n4571 PAD.n4368 0.0380882
R44889 PAD.n4575 PAD.n4368 0.0380882
R44890 PAD.n4575 PAD.n4366 0.0380882
R44891 PAD.n4583 PAD.n4366 0.0380882
R44892 PAD.n4583 PAD.n4364 0.0380882
R44893 PAD.n4587 PAD.n4364 0.0380882
R44894 PAD.n4587 PAD.n4362 0.0380882
R44895 PAD.n4595 PAD.n4362 0.0380882
R44896 PAD.n4595 PAD.n4360 0.0380882
R44897 PAD.n4599 PAD.n4360 0.0380882
R44898 PAD.n4599 PAD.n4358 0.0380882
R44899 PAD.n4607 PAD.n4358 0.0380882
R44900 PAD.n4607 PAD.n4356 0.0380882
R44901 PAD.n4611 PAD.n4356 0.0380882
R44902 PAD.n4611 PAD.n4354 0.0380882
R44903 PAD.n4619 PAD.n4354 0.0380882
R44904 PAD.n4619 PAD.n4352 0.0380882
R44905 PAD.n4623 PAD.n4352 0.0380882
R44906 PAD.n4623 PAD.n4350 0.0380882
R44907 PAD.n4631 PAD.n4350 0.0380882
R44908 PAD.n4631 PAD.n4348 0.0380882
R44909 PAD.n4635 PAD.n4348 0.0380882
R44910 PAD.n4635 PAD.n4346 0.0380882
R44911 PAD.n4643 PAD.n4346 0.0380882
R44912 PAD.n4643 PAD.n4344 0.0380882
R44913 PAD.n4647 PAD.n4344 0.0380882
R44914 PAD.n4647 PAD.n4342 0.0380882
R44915 PAD.n4655 PAD.n4342 0.0380882
R44916 PAD.n4655 PAD.n4340 0.0380882
R44917 PAD.n4660 PAD.n4340 0.0380882
R44918 PAD.n4660 PAD.n4338 0.0380882
R44919 PAD.n4338 PAD.n4337 0.0380882
R44920 PAD.n4668 PAD.n4337 0.0380882
R44921 PAD.n4417 PAD.n4325 0.0380882
R44922 PAD.n4428 PAD.n4417 0.0380882
R44923 PAD.n4429 PAD.n4428 0.0380882
R44924 PAD.n4430 PAD.n4429 0.0380882
R44925 PAD.n4430 PAD.n4413 0.0380882
R44926 PAD.n4440 PAD.n4413 0.0380882
R44927 PAD.n4441 PAD.n4440 0.0380882
R44928 PAD.n4442 PAD.n4441 0.0380882
R44929 PAD.n4442 PAD.n4409 0.0380882
R44930 PAD.n4452 PAD.n4409 0.0380882
R44931 PAD.n4453 PAD.n4452 0.0380882
R44932 PAD.n4454 PAD.n4453 0.0380882
R44933 PAD.n4454 PAD.n4405 0.0380882
R44934 PAD.n4464 PAD.n4405 0.0380882
R44935 PAD.n4465 PAD.n4464 0.0380882
R44936 PAD.n4466 PAD.n4465 0.0380882
R44937 PAD.n4466 PAD.n4401 0.0380882
R44938 PAD.n4476 PAD.n4401 0.0380882
R44939 PAD.n4477 PAD.n4476 0.0380882
R44940 PAD.n4478 PAD.n4477 0.0380882
R44941 PAD.n4478 PAD.n4397 0.0380882
R44942 PAD.n4488 PAD.n4397 0.0380882
R44943 PAD.n4489 PAD.n4488 0.0380882
R44944 PAD.n4490 PAD.n4489 0.0380882
R44945 PAD.n4490 PAD.n4393 0.0380882
R44946 PAD.n4500 PAD.n4393 0.0380882
R44947 PAD.n4501 PAD.n4500 0.0380882
R44948 PAD.n4502 PAD.n4501 0.0380882
R44949 PAD.n4502 PAD.n4389 0.0380882
R44950 PAD.n4512 PAD.n4389 0.0380882
R44951 PAD.n4513 PAD.n4512 0.0380882
R44952 PAD.n4514 PAD.n4513 0.0380882
R44953 PAD.n4514 PAD.n4385 0.0380882
R44954 PAD.n4524 PAD.n4385 0.0380882
R44955 PAD.n4525 PAD.n4524 0.0380882
R44956 PAD.n4526 PAD.n4525 0.0380882
R44957 PAD.n4526 PAD.n4381 0.0380882
R44958 PAD.n4536 PAD.n4381 0.0380882
R44959 PAD.n4537 PAD.n4536 0.0380882
R44960 PAD.n4538 PAD.n4537 0.0380882
R44961 PAD.n4538 PAD.n4377 0.0380882
R44962 PAD.n4548 PAD.n4377 0.0380882
R44963 PAD.n4549 PAD.n4548 0.0380882
R44964 PAD.n4550 PAD.n4549 0.0380882
R44965 PAD.n4550 PAD.n4373 0.0380882
R44966 PAD.n4560 PAD.n4373 0.0380882
R44967 PAD.n4561 PAD.n4560 0.0380882
R44968 PAD.n4562 PAD.n4561 0.0380882
R44969 PAD.n4562 PAD.n4369 0.0380882
R44970 PAD.n4572 PAD.n4369 0.0380882
R44971 PAD.n4573 PAD.n4572 0.0380882
R44972 PAD.n4574 PAD.n4573 0.0380882
R44973 PAD.n4574 PAD.n4365 0.0380882
R44974 PAD.n4584 PAD.n4365 0.0380882
R44975 PAD.n4585 PAD.n4584 0.0380882
R44976 PAD.n4586 PAD.n4585 0.0380882
R44977 PAD.n4586 PAD.n4361 0.0380882
R44978 PAD.n4596 PAD.n4361 0.0380882
R44979 PAD.n4597 PAD.n4596 0.0380882
R44980 PAD.n4598 PAD.n4597 0.0380882
R44981 PAD.n4598 PAD.n4357 0.0380882
R44982 PAD.n4608 PAD.n4357 0.0380882
R44983 PAD.n4609 PAD.n4608 0.0380882
R44984 PAD.n4610 PAD.n4609 0.0380882
R44985 PAD.n4610 PAD.n4353 0.0380882
R44986 PAD.n4620 PAD.n4353 0.0380882
R44987 PAD.n4621 PAD.n4620 0.0380882
R44988 PAD.n4622 PAD.n4621 0.0380882
R44989 PAD.n4622 PAD.n4349 0.0380882
R44990 PAD.n4632 PAD.n4349 0.0380882
R44991 PAD.n4633 PAD.n4632 0.0380882
R44992 PAD.n4634 PAD.n4633 0.0380882
R44993 PAD.n4634 PAD.n4345 0.0380882
R44994 PAD.n4644 PAD.n4345 0.0380882
R44995 PAD.n4645 PAD.n4644 0.0380882
R44996 PAD.n4646 PAD.n4645 0.0380882
R44997 PAD.n4646 PAD.n4341 0.0380882
R44998 PAD.n4656 PAD.n4341 0.0380882
R44999 PAD.n4657 PAD.n4656 0.0380882
R45000 PAD.n4659 PAD.n4657 0.0380882
R45001 PAD.n4659 PAD.n4658 0.0380882
R45002 PAD.n4658 PAD.n4336 0.0380882
R45003 PAD.n4669 PAD.n4336 0.0380882
R45004 PAD.n8394 PAD.n8393 0.0380882
R45005 PAD.n8393 PAD.n4728 0.0380882
R45006 PAD.n8389 PAD.n4728 0.0380882
R45007 PAD.n8389 PAD.n8385 0.0380882
R45008 PAD.n8385 PAD.n8384 0.0380882
R45009 PAD.n8384 PAD.n4730 0.0380882
R45010 PAD.n8380 PAD.n4730 0.0380882
R45011 PAD.n8380 PAD.n8376 0.0380882
R45012 PAD.n8376 PAD.n8375 0.0380882
R45013 PAD.n8375 PAD.n4735 0.0380882
R45014 PAD.n8371 PAD.n4735 0.0380882
R45015 PAD.n8371 PAD.n8367 0.0380882
R45016 PAD.n8367 PAD.n8366 0.0380882
R45017 PAD.n8366 PAD.n4740 0.0380882
R45018 PAD.n8362 PAD.n4740 0.0380882
R45019 PAD.n8362 PAD.n8358 0.0380882
R45020 PAD.n8358 PAD.n8357 0.0380882
R45021 PAD.n8357 PAD.n4745 0.0380882
R45022 PAD.n8353 PAD.n4745 0.0380882
R45023 PAD.n8353 PAD.n8349 0.0380882
R45024 PAD.n8349 PAD.n8348 0.0380882
R45025 PAD.n8348 PAD.n4750 0.0380882
R45026 PAD.n8344 PAD.n4750 0.0380882
R45027 PAD.n8344 PAD.n8340 0.0380882
R45028 PAD.n8340 PAD.n8339 0.0380882
R45029 PAD.n8339 PAD.n4755 0.0380882
R45030 PAD.n8335 PAD.n4755 0.0380882
R45031 PAD.n8335 PAD.n8331 0.0380882
R45032 PAD.n8331 PAD.n8330 0.0380882
R45033 PAD.n8330 PAD.n4760 0.0380882
R45034 PAD.n8326 PAD.n4760 0.0380882
R45035 PAD.n8326 PAD.n8322 0.0380882
R45036 PAD.n8322 PAD.n8321 0.0380882
R45037 PAD.n8321 PAD.n4765 0.0380882
R45038 PAD.n8317 PAD.n4765 0.0380882
R45039 PAD.n8317 PAD.n8313 0.0380882
R45040 PAD.n8313 PAD.n8312 0.0380882
R45041 PAD.n8312 PAD.n4770 0.0380882
R45042 PAD.n8308 PAD.n4770 0.0380882
R45043 PAD.n8308 PAD.n8304 0.0380882
R45044 PAD.n8304 PAD.n8303 0.0380882
R45045 PAD.n8303 PAD.n4775 0.0380882
R45046 PAD.n8299 PAD.n4775 0.0380882
R45047 PAD.n8299 PAD.n8295 0.0380882
R45048 PAD.n8295 PAD.n8294 0.0380882
R45049 PAD.n8294 PAD.n4780 0.0380882
R45050 PAD.n8290 PAD.n4780 0.0380882
R45051 PAD.n8290 PAD.n8286 0.0380882
R45052 PAD.n8286 PAD.n8285 0.0380882
R45053 PAD.n8285 PAD.n4785 0.0380882
R45054 PAD.n8281 PAD.n4785 0.0380882
R45055 PAD.n8281 PAD.n8277 0.0380882
R45056 PAD.n8277 PAD.n8276 0.0380882
R45057 PAD.n8276 PAD.n4790 0.0380882
R45058 PAD.n8272 PAD.n4790 0.0380882
R45059 PAD.n8272 PAD.n8268 0.0380882
R45060 PAD.n8268 PAD.n8267 0.0380882
R45061 PAD.n8267 PAD.n4795 0.0380882
R45062 PAD.n8263 PAD.n4795 0.0380882
R45063 PAD.n8263 PAD.n8259 0.0380882
R45064 PAD.n8259 PAD.n8258 0.0380882
R45065 PAD.n8258 PAD.n4800 0.0380882
R45066 PAD.n8254 PAD.n4800 0.0380882
R45067 PAD.n8254 PAD.n8250 0.0380882
R45068 PAD.n8250 PAD.n8249 0.0380882
R45069 PAD.n8249 PAD.n4805 0.0380882
R45070 PAD.n8245 PAD.n4805 0.0380882
R45071 PAD.n8245 PAD.n8241 0.0380882
R45072 PAD.n8241 PAD.n8240 0.0380882
R45073 PAD.n8240 PAD.n4810 0.0380882
R45074 PAD.n8236 PAD.n4810 0.0380882
R45075 PAD.n8236 PAD.n8232 0.0380882
R45076 PAD.n8232 PAD.n8231 0.0380882
R45077 PAD.n8231 PAD.n4815 0.0380882
R45078 PAD.n8227 PAD.n4815 0.0380882
R45079 PAD.n8227 PAD.n8223 0.0380882
R45080 PAD.n8223 PAD.n8222 0.0380882
R45081 PAD.n8222 PAD.n4820 0.0380882
R45082 PAD.n8218 PAD.n4820 0.0380882
R45083 PAD.n8218 PAD.n8214 0.0380882
R45084 PAD.n8214 PAD.n8213 0.0380882
R45085 PAD.n8213 PAD.n4825 0.0380882
R45086 PAD.n4829 PAD.n4825 0.0380882
R45087 PAD.n8392 PAD.n4676 0.0380882
R45088 PAD.n8392 PAD.n8391 0.0380882
R45089 PAD.n8391 PAD.n8390 0.0380882
R45090 PAD.n8390 PAD.n4729 0.0380882
R45091 PAD.n8383 PAD.n4729 0.0380882
R45092 PAD.n8383 PAD.n8382 0.0380882
R45093 PAD.n8382 PAD.n8381 0.0380882
R45094 PAD.n8381 PAD.n4734 0.0380882
R45095 PAD.n8374 PAD.n4734 0.0380882
R45096 PAD.n8374 PAD.n8373 0.0380882
R45097 PAD.n8373 PAD.n8372 0.0380882
R45098 PAD.n8372 PAD.n4739 0.0380882
R45099 PAD.n8365 PAD.n4739 0.0380882
R45100 PAD.n8365 PAD.n8364 0.0380882
R45101 PAD.n8364 PAD.n8363 0.0380882
R45102 PAD.n8363 PAD.n4744 0.0380882
R45103 PAD.n8356 PAD.n4744 0.0380882
R45104 PAD.n8356 PAD.n8355 0.0380882
R45105 PAD.n8355 PAD.n8354 0.0380882
R45106 PAD.n8354 PAD.n4749 0.0380882
R45107 PAD.n8347 PAD.n4749 0.0380882
R45108 PAD.n8347 PAD.n8346 0.0380882
R45109 PAD.n8346 PAD.n8345 0.0380882
R45110 PAD.n8345 PAD.n4754 0.0380882
R45111 PAD.n8338 PAD.n4754 0.0380882
R45112 PAD.n8338 PAD.n8337 0.0380882
R45113 PAD.n8337 PAD.n8336 0.0380882
R45114 PAD.n8336 PAD.n4759 0.0380882
R45115 PAD.n8329 PAD.n4759 0.0380882
R45116 PAD.n8329 PAD.n8328 0.0380882
R45117 PAD.n8328 PAD.n8327 0.0380882
R45118 PAD.n8327 PAD.n4764 0.0380882
R45119 PAD.n8320 PAD.n4764 0.0380882
R45120 PAD.n8320 PAD.n8319 0.0380882
R45121 PAD.n8319 PAD.n8318 0.0380882
R45122 PAD.n8318 PAD.n4769 0.0380882
R45123 PAD.n8311 PAD.n4769 0.0380882
R45124 PAD.n8311 PAD.n8310 0.0380882
R45125 PAD.n8310 PAD.n8309 0.0380882
R45126 PAD.n8309 PAD.n4774 0.0380882
R45127 PAD.n8302 PAD.n4774 0.0380882
R45128 PAD.n8302 PAD.n8301 0.0380882
R45129 PAD.n8301 PAD.n8300 0.0380882
R45130 PAD.n8300 PAD.n4779 0.0380882
R45131 PAD.n8293 PAD.n4779 0.0380882
R45132 PAD.n8293 PAD.n8292 0.0380882
R45133 PAD.n8292 PAD.n8291 0.0380882
R45134 PAD.n8291 PAD.n4784 0.0380882
R45135 PAD.n8284 PAD.n4784 0.0380882
R45136 PAD.n8284 PAD.n8283 0.0380882
R45137 PAD.n8283 PAD.n8282 0.0380882
R45138 PAD.n8282 PAD.n4789 0.0380882
R45139 PAD.n8275 PAD.n4789 0.0380882
R45140 PAD.n8275 PAD.n8274 0.0380882
R45141 PAD.n8274 PAD.n8273 0.0380882
R45142 PAD.n8273 PAD.n4794 0.0380882
R45143 PAD.n8266 PAD.n4794 0.0380882
R45144 PAD.n8266 PAD.n8265 0.0380882
R45145 PAD.n8265 PAD.n8264 0.0380882
R45146 PAD.n8264 PAD.n4799 0.0380882
R45147 PAD.n8257 PAD.n4799 0.0380882
R45148 PAD.n8257 PAD.n8256 0.0380882
R45149 PAD.n8256 PAD.n8255 0.0380882
R45150 PAD.n8255 PAD.n4804 0.0380882
R45151 PAD.n8248 PAD.n4804 0.0380882
R45152 PAD.n8248 PAD.n8247 0.0380882
R45153 PAD.n8247 PAD.n8246 0.0380882
R45154 PAD.n8246 PAD.n4809 0.0380882
R45155 PAD.n8239 PAD.n4809 0.0380882
R45156 PAD.n8239 PAD.n8238 0.0380882
R45157 PAD.n8238 PAD.n8237 0.0380882
R45158 PAD.n8237 PAD.n4814 0.0380882
R45159 PAD.n8230 PAD.n4814 0.0380882
R45160 PAD.n8230 PAD.n8229 0.0380882
R45161 PAD.n8229 PAD.n8228 0.0380882
R45162 PAD.n8228 PAD.n4819 0.0380882
R45163 PAD.n8221 PAD.n4819 0.0380882
R45164 PAD.n8221 PAD.n8220 0.0380882
R45165 PAD.n8220 PAD.n8219 0.0380882
R45166 PAD.n8219 PAD.n4824 0.0380882
R45167 PAD.n8212 PAD.n4824 0.0380882
R45168 PAD.n8212 PAD.n8211 0.0380882
R45169 PAD.n8211 PAD.n8210 0.0380882
R45170 PAD.n5178 PAD.n5177 0.0380882
R45171 PAD.n5177 PAD.n4848 0.0380882
R45172 PAD.n5171 PAD.n4848 0.0380882
R45173 PAD.n5171 PAD.n4851 0.0380882
R45174 PAD.n5167 PAD.n4851 0.0380882
R45175 PAD.n5167 PAD.n4854 0.0380882
R45176 PAD.n5159 PAD.n4854 0.0380882
R45177 PAD.n5159 PAD.n4856 0.0380882
R45178 PAD.n5155 PAD.n4856 0.0380882
R45179 PAD.n5155 PAD.n4858 0.0380882
R45180 PAD.n5147 PAD.n4858 0.0380882
R45181 PAD.n5147 PAD.n4860 0.0380882
R45182 PAD.n5143 PAD.n4860 0.0380882
R45183 PAD.n5143 PAD.n4862 0.0380882
R45184 PAD.n5135 PAD.n4862 0.0380882
R45185 PAD.n5135 PAD.n4864 0.0380882
R45186 PAD.n5131 PAD.n4864 0.0380882
R45187 PAD.n5131 PAD.n4866 0.0380882
R45188 PAD.n5123 PAD.n4866 0.0380882
R45189 PAD.n5123 PAD.n4868 0.0380882
R45190 PAD.n5119 PAD.n4868 0.0380882
R45191 PAD.n5119 PAD.n4870 0.0380882
R45192 PAD.n5111 PAD.n4870 0.0380882
R45193 PAD.n5111 PAD.n4872 0.0380882
R45194 PAD.n5107 PAD.n4872 0.0380882
R45195 PAD.n5107 PAD.n4874 0.0380882
R45196 PAD.n5099 PAD.n4874 0.0380882
R45197 PAD.n5099 PAD.n4876 0.0380882
R45198 PAD.n5095 PAD.n4876 0.0380882
R45199 PAD.n5095 PAD.n4878 0.0380882
R45200 PAD.n5087 PAD.n4878 0.0380882
R45201 PAD.n5087 PAD.n4880 0.0380882
R45202 PAD.n5083 PAD.n4880 0.0380882
R45203 PAD.n5083 PAD.n4882 0.0380882
R45204 PAD.n5075 PAD.n4882 0.0380882
R45205 PAD.n5075 PAD.n4884 0.0380882
R45206 PAD.n5071 PAD.n4884 0.0380882
R45207 PAD.n5071 PAD.n4886 0.0380882
R45208 PAD.n5063 PAD.n4886 0.0380882
R45209 PAD.n5063 PAD.n4888 0.0380882
R45210 PAD.n5059 PAD.n4888 0.0380882
R45211 PAD.n5059 PAD.n4890 0.0380882
R45212 PAD.n5051 PAD.n4890 0.0380882
R45213 PAD.n5051 PAD.n4892 0.0380882
R45214 PAD.n5047 PAD.n4892 0.0380882
R45215 PAD.n5047 PAD.n4894 0.0380882
R45216 PAD.n5039 PAD.n4894 0.0380882
R45217 PAD.n5039 PAD.n4896 0.0380882
R45218 PAD.n5035 PAD.n4896 0.0380882
R45219 PAD.n5035 PAD.n4898 0.0380882
R45220 PAD.n5027 PAD.n4898 0.0380882
R45221 PAD.n5027 PAD.n4900 0.0380882
R45222 PAD.n5023 PAD.n4900 0.0380882
R45223 PAD.n5023 PAD.n4902 0.0380882
R45224 PAD.n5015 PAD.n4902 0.0380882
R45225 PAD.n5015 PAD.n4904 0.0380882
R45226 PAD.n5011 PAD.n4904 0.0380882
R45227 PAD.n5011 PAD.n4906 0.0380882
R45228 PAD.n5003 PAD.n4906 0.0380882
R45229 PAD.n5003 PAD.n4908 0.0380882
R45230 PAD.n4999 PAD.n4908 0.0380882
R45231 PAD.n4999 PAD.n4910 0.0380882
R45232 PAD.n4991 PAD.n4910 0.0380882
R45233 PAD.n4991 PAD.n4912 0.0380882
R45234 PAD.n4987 PAD.n4912 0.0380882
R45235 PAD.n4987 PAD.n4914 0.0380882
R45236 PAD.n4979 PAD.n4914 0.0380882
R45237 PAD.n4979 PAD.n4916 0.0380882
R45238 PAD.n4975 PAD.n4916 0.0380882
R45239 PAD.n4975 PAD.n4918 0.0380882
R45240 PAD.n4967 PAD.n4918 0.0380882
R45241 PAD.n4967 PAD.n4920 0.0380882
R45242 PAD.n4963 PAD.n4920 0.0380882
R45243 PAD.n4963 PAD.n4922 0.0380882
R45244 PAD.n4955 PAD.n4922 0.0380882
R45245 PAD.n4955 PAD.n4924 0.0380882
R45246 PAD.n4951 PAD.n4924 0.0380882
R45247 PAD.n4951 PAD.n4926 0.0380882
R45248 PAD.n4943 PAD.n4926 0.0380882
R45249 PAD.n4943 PAD.n4928 0.0380882
R45250 PAD.n4939 PAD.n4928 0.0380882
R45251 PAD.n4939 PAD.n4930 0.0380882
R45252 PAD.n4931 PAD.n4930 0.0380882
R45253 PAD.n5179 PAD.n4846 0.0380882
R45254 PAD.n4852 PAD.n4846 0.0380882
R45255 PAD.n5170 PAD.n4852 0.0380882
R45256 PAD.n5170 PAD.n5169 0.0380882
R45257 PAD.n5169 PAD.n5168 0.0380882
R45258 PAD.n5168 PAD.n4853 0.0380882
R45259 PAD.n5158 PAD.n4853 0.0380882
R45260 PAD.n5158 PAD.n5157 0.0380882
R45261 PAD.n5157 PAD.n5156 0.0380882
R45262 PAD.n5156 PAD.n4857 0.0380882
R45263 PAD.n5146 PAD.n4857 0.0380882
R45264 PAD.n5146 PAD.n5145 0.0380882
R45265 PAD.n5145 PAD.n5144 0.0380882
R45266 PAD.n5144 PAD.n4861 0.0380882
R45267 PAD.n5134 PAD.n4861 0.0380882
R45268 PAD.n5134 PAD.n5133 0.0380882
R45269 PAD.n5133 PAD.n5132 0.0380882
R45270 PAD.n5132 PAD.n4865 0.0380882
R45271 PAD.n5122 PAD.n4865 0.0380882
R45272 PAD.n5122 PAD.n5121 0.0380882
R45273 PAD.n5121 PAD.n5120 0.0380882
R45274 PAD.n5120 PAD.n4869 0.0380882
R45275 PAD.n5110 PAD.n4869 0.0380882
R45276 PAD.n5110 PAD.n5109 0.0380882
R45277 PAD.n5109 PAD.n5108 0.0380882
R45278 PAD.n5108 PAD.n4873 0.0380882
R45279 PAD.n5098 PAD.n4873 0.0380882
R45280 PAD.n5098 PAD.n5097 0.0380882
R45281 PAD.n5097 PAD.n5096 0.0380882
R45282 PAD.n5096 PAD.n4877 0.0380882
R45283 PAD.n5086 PAD.n4877 0.0380882
R45284 PAD.n5086 PAD.n5085 0.0380882
R45285 PAD.n5085 PAD.n5084 0.0380882
R45286 PAD.n5084 PAD.n4881 0.0380882
R45287 PAD.n5074 PAD.n4881 0.0380882
R45288 PAD.n5074 PAD.n5073 0.0380882
R45289 PAD.n5073 PAD.n5072 0.0380882
R45290 PAD.n5072 PAD.n4885 0.0380882
R45291 PAD.n5062 PAD.n4885 0.0380882
R45292 PAD.n5062 PAD.n5061 0.0380882
R45293 PAD.n5061 PAD.n5060 0.0380882
R45294 PAD.n5060 PAD.n4889 0.0380882
R45295 PAD.n5050 PAD.n4889 0.0380882
R45296 PAD.n5050 PAD.n5049 0.0380882
R45297 PAD.n5049 PAD.n5048 0.0380882
R45298 PAD.n5048 PAD.n4893 0.0380882
R45299 PAD.n5038 PAD.n4893 0.0380882
R45300 PAD.n5038 PAD.n5037 0.0380882
R45301 PAD.n5037 PAD.n5036 0.0380882
R45302 PAD.n5036 PAD.n4897 0.0380882
R45303 PAD.n5026 PAD.n4897 0.0380882
R45304 PAD.n5026 PAD.n5025 0.0380882
R45305 PAD.n5025 PAD.n5024 0.0380882
R45306 PAD.n5024 PAD.n4901 0.0380882
R45307 PAD.n5014 PAD.n4901 0.0380882
R45308 PAD.n5014 PAD.n5013 0.0380882
R45309 PAD.n5013 PAD.n5012 0.0380882
R45310 PAD.n5012 PAD.n4905 0.0380882
R45311 PAD.n5002 PAD.n4905 0.0380882
R45312 PAD.n5002 PAD.n5001 0.0380882
R45313 PAD.n5001 PAD.n5000 0.0380882
R45314 PAD.n5000 PAD.n4909 0.0380882
R45315 PAD.n4990 PAD.n4909 0.0380882
R45316 PAD.n4990 PAD.n4989 0.0380882
R45317 PAD.n4989 PAD.n4988 0.0380882
R45318 PAD.n4988 PAD.n4913 0.0380882
R45319 PAD.n4978 PAD.n4913 0.0380882
R45320 PAD.n4978 PAD.n4977 0.0380882
R45321 PAD.n4977 PAD.n4976 0.0380882
R45322 PAD.n4976 PAD.n4917 0.0380882
R45323 PAD.n4966 PAD.n4917 0.0380882
R45324 PAD.n4966 PAD.n4965 0.0380882
R45325 PAD.n4965 PAD.n4964 0.0380882
R45326 PAD.n4964 PAD.n4921 0.0380882
R45327 PAD.n4954 PAD.n4921 0.0380882
R45328 PAD.n4954 PAD.n4953 0.0380882
R45329 PAD.n4953 PAD.n4952 0.0380882
R45330 PAD.n4952 PAD.n4925 0.0380882
R45331 PAD.n4942 PAD.n4925 0.0380882
R45332 PAD.n4942 PAD.n4941 0.0380882
R45333 PAD.n4941 PAD.n4940 0.0380882
R45334 PAD.n4940 PAD.n4929 0.0380882
R45335 PAD.n4929 PAD.n4835 0.0380882
R45336 PAD.n8160 PAD.n8159 0.0380882
R45337 PAD.n8159 PAD.n7874 0.0380882
R45338 PAD.n8155 PAD.n7874 0.0380882
R45339 PAD.n8155 PAD.n8151 0.0380882
R45340 PAD.n8151 PAD.n8150 0.0380882
R45341 PAD.n8150 PAD.n7876 0.0380882
R45342 PAD.n8146 PAD.n7876 0.0380882
R45343 PAD.n8146 PAD.n8142 0.0380882
R45344 PAD.n8142 PAD.n8141 0.0380882
R45345 PAD.n8141 PAD.n7881 0.0380882
R45346 PAD.n8137 PAD.n7881 0.0380882
R45347 PAD.n8137 PAD.n8133 0.0380882
R45348 PAD.n8133 PAD.n8132 0.0380882
R45349 PAD.n8132 PAD.n7886 0.0380882
R45350 PAD.n8128 PAD.n7886 0.0380882
R45351 PAD.n8128 PAD.n8124 0.0380882
R45352 PAD.n8124 PAD.n8123 0.0380882
R45353 PAD.n8123 PAD.n7891 0.0380882
R45354 PAD.n8119 PAD.n7891 0.0380882
R45355 PAD.n8119 PAD.n8115 0.0380882
R45356 PAD.n8115 PAD.n8114 0.0380882
R45357 PAD.n8114 PAD.n7896 0.0380882
R45358 PAD.n8110 PAD.n7896 0.0380882
R45359 PAD.n8110 PAD.n8106 0.0380882
R45360 PAD.n8106 PAD.n8105 0.0380882
R45361 PAD.n8105 PAD.n7901 0.0380882
R45362 PAD.n8101 PAD.n7901 0.0380882
R45363 PAD.n8101 PAD.n8097 0.0380882
R45364 PAD.n8097 PAD.n8096 0.0380882
R45365 PAD.n8096 PAD.n7906 0.0380882
R45366 PAD.n8092 PAD.n7906 0.0380882
R45367 PAD.n8092 PAD.n8088 0.0380882
R45368 PAD.n8088 PAD.n8087 0.0380882
R45369 PAD.n8087 PAD.n7911 0.0380882
R45370 PAD.n8083 PAD.n7911 0.0380882
R45371 PAD.n8083 PAD.n8079 0.0380882
R45372 PAD.n8079 PAD.n8078 0.0380882
R45373 PAD.n8078 PAD.n7916 0.0380882
R45374 PAD.n8074 PAD.n7916 0.0380882
R45375 PAD.n8074 PAD.n8070 0.0380882
R45376 PAD.n8070 PAD.n8069 0.0380882
R45377 PAD.n8069 PAD.n7921 0.0380882
R45378 PAD.n8065 PAD.n7921 0.0380882
R45379 PAD.n8065 PAD.n8061 0.0380882
R45380 PAD.n8061 PAD.n8060 0.0380882
R45381 PAD.n8060 PAD.n7926 0.0380882
R45382 PAD.n8056 PAD.n7926 0.0380882
R45383 PAD.n8056 PAD.n8052 0.0380882
R45384 PAD.n8052 PAD.n8051 0.0380882
R45385 PAD.n8051 PAD.n7931 0.0380882
R45386 PAD.n8047 PAD.n7931 0.0380882
R45387 PAD.n8047 PAD.n8043 0.0380882
R45388 PAD.n8043 PAD.n8042 0.0380882
R45389 PAD.n8042 PAD.n7936 0.0380882
R45390 PAD.n8038 PAD.n7936 0.0380882
R45391 PAD.n8038 PAD.n8034 0.0380882
R45392 PAD.n8034 PAD.n8033 0.0380882
R45393 PAD.n8033 PAD.n7941 0.0380882
R45394 PAD.n8029 PAD.n7941 0.0380882
R45395 PAD.n8029 PAD.n8025 0.0380882
R45396 PAD.n8025 PAD.n8024 0.0380882
R45397 PAD.n8024 PAD.n7946 0.0380882
R45398 PAD.n8020 PAD.n7946 0.0380882
R45399 PAD.n8020 PAD.n8016 0.0380882
R45400 PAD.n8016 PAD.n8015 0.0380882
R45401 PAD.n8015 PAD.n7951 0.0380882
R45402 PAD.n8011 PAD.n7951 0.0380882
R45403 PAD.n8011 PAD.n8007 0.0380882
R45404 PAD.n8007 PAD.n8006 0.0380882
R45405 PAD.n8006 PAD.n7956 0.0380882
R45406 PAD.n8002 PAD.n7956 0.0380882
R45407 PAD.n8002 PAD.n7998 0.0380882
R45408 PAD.n7998 PAD.n7997 0.0380882
R45409 PAD.n7997 PAD.n7961 0.0380882
R45410 PAD.n7993 PAD.n7961 0.0380882
R45411 PAD.n7993 PAD.n7989 0.0380882
R45412 PAD.n7989 PAD.n7988 0.0380882
R45413 PAD.n7988 PAD.n7966 0.0380882
R45414 PAD.n7984 PAD.n7966 0.0380882
R45415 PAD.n7984 PAD.n7980 0.0380882
R45416 PAD.n7980 PAD.n7979 0.0380882
R45417 PAD.n7979 PAD.n7973 0.0380882
R45418 PAD.n7973 PAD.n7972 0.0380882
R45419 PAD.n8158 PAD.n5193 0.0380882
R45420 PAD.n8158 PAD.n8157 0.0380882
R45421 PAD.n8157 PAD.n8156 0.0380882
R45422 PAD.n8156 PAD.n7875 0.0380882
R45423 PAD.n8149 PAD.n7875 0.0380882
R45424 PAD.n8149 PAD.n8148 0.0380882
R45425 PAD.n8148 PAD.n8147 0.0380882
R45426 PAD.n8147 PAD.n7880 0.0380882
R45427 PAD.n8140 PAD.n7880 0.0380882
R45428 PAD.n8140 PAD.n8139 0.0380882
R45429 PAD.n8139 PAD.n8138 0.0380882
R45430 PAD.n8138 PAD.n7885 0.0380882
R45431 PAD.n8131 PAD.n7885 0.0380882
R45432 PAD.n8131 PAD.n8130 0.0380882
R45433 PAD.n8130 PAD.n8129 0.0380882
R45434 PAD.n8129 PAD.n7890 0.0380882
R45435 PAD.n8122 PAD.n7890 0.0380882
R45436 PAD.n8122 PAD.n8121 0.0380882
R45437 PAD.n8121 PAD.n8120 0.0380882
R45438 PAD.n8120 PAD.n7895 0.0380882
R45439 PAD.n8113 PAD.n7895 0.0380882
R45440 PAD.n8113 PAD.n8112 0.0380882
R45441 PAD.n8112 PAD.n8111 0.0380882
R45442 PAD.n8111 PAD.n7900 0.0380882
R45443 PAD.n8104 PAD.n7900 0.0380882
R45444 PAD.n8104 PAD.n8103 0.0380882
R45445 PAD.n8103 PAD.n8102 0.0380882
R45446 PAD.n8102 PAD.n7905 0.0380882
R45447 PAD.n8095 PAD.n7905 0.0380882
R45448 PAD.n8095 PAD.n8094 0.0380882
R45449 PAD.n8094 PAD.n8093 0.0380882
R45450 PAD.n8093 PAD.n7910 0.0380882
R45451 PAD.n8086 PAD.n7910 0.0380882
R45452 PAD.n8086 PAD.n8085 0.0380882
R45453 PAD.n8085 PAD.n8084 0.0380882
R45454 PAD.n8084 PAD.n7915 0.0380882
R45455 PAD.n8077 PAD.n7915 0.0380882
R45456 PAD.n8077 PAD.n8076 0.0380882
R45457 PAD.n8076 PAD.n8075 0.0380882
R45458 PAD.n8075 PAD.n7920 0.0380882
R45459 PAD.n8068 PAD.n7920 0.0380882
R45460 PAD.n8068 PAD.n8067 0.0380882
R45461 PAD.n8067 PAD.n8066 0.0380882
R45462 PAD.n8066 PAD.n7925 0.0380882
R45463 PAD.n8059 PAD.n7925 0.0380882
R45464 PAD.n8059 PAD.n8058 0.0380882
R45465 PAD.n8058 PAD.n8057 0.0380882
R45466 PAD.n8057 PAD.n7930 0.0380882
R45467 PAD.n8050 PAD.n7930 0.0380882
R45468 PAD.n8050 PAD.n8049 0.0380882
R45469 PAD.n8049 PAD.n8048 0.0380882
R45470 PAD.n8048 PAD.n7935 0.0380882
R45471 PAD.n8041 PAD.n7935 0.0380882
R45472 PAD.n8041 PAD.n8040 0.0380882
R45473 PAD.n8040 PAD.n8039 0.0380882
R45474 PAD.n8039 PAD.n7940 0.0380882
R45475 PAD.n8032 PAD.n7940 0.0380882
R45476 PAD.n8032 PAD.n8031 0.0380882
R45477 PAD.n8031 PAD.n8030 0.0380882
R45478 PAD.n8030 PAD.n7945 0.0380882
R45479 PAD.n8023 PAD.n7945 0.0380882
R45480 PAD.n8023 PAD.n8022 0.0380882
R45481 PAD.n8022 PAD.n8021 0.0380882
R45482 PAD.n8021 PAD.n7950 0.0380882
R45483 PAD.n8014 PAD.n7950 0.0380882
R45484 PAD.n8014 PAD.n8013 0.0380882
R45485 PAD.n8013 PAD.n8012 0.0380882
R45486 PAD.n8012 PAD.n7955 0.0380882
R45487 PAD.n8005 PAD.n7955 0.0380882
R45488 PAD.n8005 PAD.n8004 0.0380882
R45489 PAD.n8004 PAD.n8003 0.0380882
R45490 PAD.n8003 PAD.n7960 0.0380882
R45491 PAD.n7996 PAD.n7960 0.0380882
R45492 PAD.n7996 PAD.n7995 0.0380882
R45493 PAD.n7995 PAD.n7994 0.0380882
R45494 PAD.n7994 PAD.n7965 0.0380882
R45495 PAD.n7987 PAD.n7965 0.0380882
R45496 PAD.n7987 PAD.n7986 0.0380882
R45497 PAD.n7986 PAD.n7985 0.0380882
R45498 PAD.n7985 PAD.n7970 0.0380882
R45499 PAD.n7978 PAD.n7970 0.0380882
R45500 PAD.n7978 PAD.n7977 0.0380882
R45501 PAD.n7977 PAD.n5186 0.0380882
R45502 PAD.n5542 PAD.n5541 0.0380882
R45503 PAD.n5541 PAD.n5212 0.0380882
R45504 PAD.n5535 PAD.n5212 0.0380882
R45505 PAD.n5535 PAD.n5215 0.0380882
R45506 PAD.n5531 PAD.n5215 0.0380882
R45507 PAD.n5531 PAD.n5218 0.0380882
R45508 PAD.n5523 PAD.n5218 0.0380882
R45509 PAD.n5523 PAD.n5220 0.0380882
R45510 PAD.n5519 PAD.n5220 0.0380882
R45511 PAD.n5519 PAD.n5222 0.0380882
R45512 PAD.n5511 PAD.n5222 0.0380882
R45513 PAD.n5511 PAD.n5224 0.0380882
R45514 PAD.n5507 PAD.n5224 0.0380882
R45515 PAD.n5507 PAD.n5226 0.0380882
R45516 PAD.n5499 PAD.n5226 0.0380882
R45517 PAD.n5499 PAD.n5228 0.0380882
R45518 PAD.n5495 PAD.n5228 0.0380882
R45519 PAD.n5495 PAD.n5230 0.0380882
R45520 PAD.n5487 PAD.n5230 0.0380882
R45521 PAD.n5487 PAD.n5232 0.0380882
R45522 PAD.n5483 PAD.n5232 0.0380882
R45523 PAD.n5483 PAD.n5234 0.0380882
R45524 PAD.n5475 PAD.n5234 0.0380882
R45525 PAD.n5475 PAD.n5236 0.0380882
R45526 PAD.n5471 PAD.n5236 0.0380882
R45527 PAD.n5471 PAD.n5238 0.0380882
R45528 PAD.n5463 PAD.n5238 0.0380882
R45529 PAD.n5463 PAD.n5240 0.0380882
R45530 PAD.n5459 PAD.n5240 0.0380882
R45531 PAD.n5459 PAD.n5242 0.0380882
R45532 PAD.n5451 PAD.n5242 0.0380882
R45533 PAD.n5451 PAD.n5244 0.0380882
R45534 PAD.n5447 PAD.n5244 0.0380882
R45535 PAD.n5447 PAD.n5246 0.0380882
R45536 PAD.n5439 PAD.n5246 0.0380882
R45537 PAD.n5439 PAD.n5248 0.0380882
R45538 PAD.n5435 PAD.n5248 0.0380882
R45539 PAD.n5435 PAD.n5250 0.0380882
R45540 PAD.n5427 PAD.n5250 0.0380882
R45541 PAD.n5427 PAD.n5252 0.0380882
R45542 PAD.n5423 PAD.n5252 0.0380882
R45543 PAD.n5423 PAD.n5254 0.0380882
R45544 PAD.n5415 PAD.n5254 0.0380882
R45545 PAD.n5415 PAD.n5256 0.0380882
R45546 PAD.n5411 PAD.n5256 0.0380882
R45547 PAD.n5411 PAD.n5258 0.0380882
R45548 PAD.n5403 PAD.n5258 0.0380882
R45549 PAD.n5403 PAD.n5260 0.0380882
R45550 PAD.n5399 PAD.n5260 0.0380882
R45551 PAD.n5399 PAD.n5262 0.0380882
R45552 PAD.n5391 PAD.n5262 0.0380882
R45553 PAD.n5391 PAD.n5264 0.0380882
R45554 PAD.n5387 PAD.n5264 0.0380882
R45555 PAD.n5387 PAD.n5266 0.0380882
R45556 PAD.n5379 PAD.n5266 0.0380882
R45557 PAD.n5379 PAD.n5268 0.0380882
R45558 PAD.n5375 PAD.n5268 0.0380882
R45559 PAD.n5375 PAD.n5270 0.0380882
R45560 PAD.n5367 PAD.n5270 0.0380882
R45561 PAD.n5367 PAD.n5272 0.0380882
R45562 PAD.n5363 PAD.n5272 0.0380882
R45563 PAD.n5363 PAD.n5274 0.0380882
R45564 PAD.n5355 PAD.n5274 0.0380882
R45565 PAD.n5355 PAD.n5276 0.0380882
R45566 PAD.n5351 PAD.n5276 0.0380882
R45567 PAD.n5351 PAD.n5278 0.0380882
R45568 PAD.n5343 PAD.n5278 0.0380882
R45569 PAD.n5343 PAD.n5280 0.0380882
R45570 PAD.n5339 PAD.n5280 0.0380882
R45571 PAD.n5339 PAD.n5282 0.0380882
R45572 PAD.n5331 PAD.n5282 0.0380882
R45573 PAD.n5331 PAD.n5284 0.0380882
R45574 PAD.n5327 PAD.n5284 0.0380882
R45575 PAD.n5327 PAD.n5286 0.0380882
R45576 PAD.n5319 PAD.n5286 0.0380882
R45577 PAD.n5319 PAD.n5288 0.0380882
R45578 PAD.n5315 PAD.n5288 0.0380882
R45579 PAD.n5315 PAD.n5290 0.0380882
R45580 PAD.n5307 PAD.n5290 0.0380882
R45581 PAD.n5307 PAD.n5292 0.0380882
R45582 PAD.n5303 PAD.n5292 0.0380882
R45583 PAD.n5303 PAD.n5294 0.0380882
R45584 PAD.n5295 PAD.n5294 0.0380882
R45585 PAD.n5543 PAD.n5210 0.0380882
R45586 PAD.n5216 PAD.n5210 0.0380882
R45587 PAD.n5534 PAD.n5216 0.0380882
R45588 PAD.n5534 PAD.n5533 0.0380882
R45589 PAD.n5533 PAD.n5532 0.0380882
R45590 PAD.n5532 PAD.n5217 0.0380882
R45591 PAD.n5522 PAD.n5217 0.0380882
R45592 PAD.n5522 PAD.n5521 0.0380882
R45593 PAD.n5521 PAD.n5520 0.0380882
R45594 PAD.n5520 PAD.n5221 0.0380882
R45595 PAD.n5510 PAD.n5221 0.0380882
R45596 PAD.n5510 PAD.n5509 0.0380882
R45597 PAD.n5509 PAD.n5508 0.0380882
R45598 PAD.n5508 PAD.n5225 0.0380882
R45599 PAD.n5498 PAD.n5225 0.0380882
R45600 PAD.n5498 PAD.n5497 0.0380882
R45601 PAD.n5497 PAD.n5496 0.0380882
R45602 PAD.n5496 PAD.n5229 0.0380882
R45603 PAD.n5486 PAD.n5229 0.0380882
R45604 PAD.n5486 PAD.n5485 0.0380882
R45605 PAD.n5485 PAD.n5484 0.0380882
R45606 PAD.n5484 PAD.n5233 0.0380882
R45607 PAD.n5474 PAD.n5233 0.0380882
R45608 PAD.n5474 PAD.n5473 0.0380882
R45609 PAD.n5473 PAD.n5472 0.0380882
R45610 PAD.n5472 PAD.n5237 0.0380882
R45611 PAD.n5462 PAD.n5237 0.0380882
R45612 PAD.n5462 PAD.n5461 0.0380882
R45613 PAD.n5461 PAD.n5460 0.0380882
R45614 PAD.n5460 PAD.n5241 0.0380882
R45615 PAD.n5450 PAD.n5241 0.0380882
R45616 PAD.n5450 PAD.n5449 0.0380882
R45617 PAD.n5449 PAD.n5448 0.0380882
R45618 PAD.n5448 PAD.n5245 0.0380882
R45619 PAD.n5438 PAD.n5245 0.0380882
R45620 PAD.n5438 PAD.n5437 0.0380882
R45621 PAD.n5437 PAD.n5436 0.0380882
R45622 PAD.n5436 PAD.n5249 0.0380882
R45623 PAD.n5426 PAD.n5249 0.0380882
R45624 PAD.n5426 PAD.n5425 0.0380882
R45625 PAD.n5425 PAD.n5424 0.0380882
R45626 PAD.n5424 PAD.n5253 0.0380882
R45627 PAD.n5414 PAD.n5253 0.0380882
R45628 PAD.n5414 PAD.n5413 0.0380882
R45629 PAD.n5413 PAD.n5412 0.0380882
R45630 PAD.n5412 PAD.n5257 0.0380882
R45631 PAD.n5402 PAD.n5257 0.0380882
R45632 PAD.n5402 PAD.n5401 0.0380882
R45633 PAD.n5401 PAD.n5400 0.0380882
R45634 PAD.n5400 PAD.n5261 0.0380882
R45635 PAD.n5390 PAD.n5261 0.0380882
R45636 PAD.n5390 PAD.n5389 0.0380882
R45637 PAD.n5389 PAD.n5388 0.0380882
R45638 PAD.n5388 PAD.n5265 0.0380882
R45639 PAD.n5378 PAD.n5265 0.0380882
R45640 PAD.n5378 PAD.n5377 0.0380882
R45641 PAD.n5377 PAD.n5376 0.0380882
R45642 PAD.n5376 PAD.n5269 0.0380882
R45643 PAD.n5366 PAD.n5269 0.0380882
R45644 PAD.n5366 PAD.n5365 0.0380882
R45645 PAD.n5365 PAD.n5364 0.0380882
R45646 PAD.n5364 PAD.n5273 0.0380882
R45647 PAD.n5354 PAD.n5273 0.0380882
R45648 PAD.n5354 PAD.n5353 0.0380882
R45649 PAD.n5353 PAD.n5352 0.0380882
R45650 PAD.n5352 PAD.n5277 0.0380882
R45651 PAD.n5342 PAD.n5277 0.0380882
R45652 PAD.n5342 PAD.n5341 0.0380882
R45653 PAD.n5341 PAD.n5340 0.0380882
R45654 PAD.n5340 PAD.n5281 0.0380882
R45655 PAD.n5330 PAD.n5281 0.0380882
R45656 PAD.n5330 PAD.n5329 0.0380882
R45657 PAD.n5329 PAD.n5328 0.0380882
R45658 PAD.n5328 PAD.n5285 0.0380882
R45659 PAD.n5318 PAD.n5285 0.0380882
R45660 PAD.n5318 PAD.n5317 0.0380882
R45661 PAD.n5317 PAD.n5316 0.0380882
R45662 PAD.n5316 PAD.n5289 0.0380882
R45663 PAD.n5306 PAD.n5289 0.0380882
R45664 PAD.n5306 PAD.n5305 0.0380882
R45665 PAD.n5305 PAD.n5304 0.0380882
R45666 PAD.n5304 PAD.n5293 0.0380882
R45667 PAD.n5293 PAD.n5200 0.0380882
R45668 PAD.n7779 PAD.n7106 0.0380882
R45669 PAD.n7775 PAD.n7106 0.0380882
R45670 PAD.n7775 PAD.n7772 0.0380882
R45671 PAD.n7772 PAD.n7768 0.0380882
R45672 PAD.n7768 PAD.n7108 0.0380882
R45673 PAD.n7764 PAD.n7108 0.0380882
R45674 PAD.n7764 PAD.n7760 0.0380882
R45675 PAD.n7760 PAD.n7756 0.0380882
R45676 PAD.n7756 PAD.n7110 0.0380882
R45677 PAD.n7752 PAD.n7110 0.0380882
R45678 PAD.n7752 PAD.n7748 0.0380882
R45679 PAD.n7748 PAD.n7744 0.0380882
R45680 PAD.n7744 PAD.n7112 0.0380882
R45681 PAD.n7740 PAD.n7112 0.0380882
R45682 PAD.n7740 PAD.n7736 0.0380882
R45683 PAD.n7736 PAD.n7732 0.0380882
R45684 PAD.n7732 PAD.n7114 0.0380882
R45685 PAD.n7728 PAD.n7114 0.0380882
R45686 PAD.n7728 PAD.n7724 0.0380882
R45687 PAD.n7724 PAD.n7720 0.0380882
R45688 PAD.n7720 PAD.n7116 0.0380882
R45689 PAD.n7716 PAD.n7116 0.0380882
R45690 PAD.n7716 PAD.n7712 0.0380882
R45691 PAD.n7712 PAD.n7708 0.0380882
R45692 PAD.n7708 PAD.n7118 0.0380882
R45693 PAD.n7704 PAD.n7118 0.0380882
R45694 PAD.n7704 PAD.n7700 0.0380882
R45695 PAD.n7700 PAD.n7696 0.0380882
R45696 PAD.n7696 PAD.n7120 0.0380882
R45697 PAD.n7692 PAD.n7120 0.0380882
R45698 PAD.n7692 PAD.n7688 0.0380882
R45699 PAD.n7688 PAD.n7684 0.0380882
R45700 PAD.n7684 PAD.n7122 0.0380882
R45701 PAD.n7680 PAD.n7122 0.0380882
R45702 PAD.n7680 PAD.n7676 0.0380882
R45703 PAD.n7676 PAD.n7672 0.0380882
R45704 PAD.n7672 PAD.n7124 0.0380882
R45705 PAD.n7668 PAD.n7124 0.0380882
R45706 PAD.n7668 PAD.n7664 0.0380882
R45707 PAD.n7664 PAD.n7660 0.0380882
R45708 PAD.n7660 PAD.n7126 0.0380882
R45709 PAD.n7656 PAD.n7126 0.0380882
R45710 PAD.n7656 PAD.n7652 0.0380882
R45711 PAD.n7652 PAD.n7648 0.0380882
R45712 PAD.n7648 PAD.n7128 0.0380882
R45713 PAD.n7644 PAD.n7128 0.0380882
R45714 PAD.n7644 PAD.n7640 0.0380882
R45715 PAD.n7640 PAD.n7636 0.0380882
R45716 PAD.n7636 PAD.n7130 0.0380882
R45717 PAD.n7632 PAD.n7130 0.0380882
R45718 PAD.n7632 PAD.n7628 0.0380882
R45719 PAD.n7628 PAD.n7624 0.0380882
R45720 PAD.n7624 PAD.n7132 0.0380882
R45721 PAD.n7620 PAD.n7132 0.0380882
R45722 PAD.n7620 PAD.n7616 0.0380882
R45723 PAD.n7616 PAD.n7612 0.0380882
R45724 PAD.n7612 PAD.n7134 0.0380882
R45725 PAD.n7608 PAD.n7134 0.0380882
R45726 PAD.n7608 PAD.n7604 0.0380882
R45727 PAD.n7604 PAD.n7600 0.0380882
R45728 PAD.n7600 PAD.n7136 0.0380882
R45729 PAD.n7596 PAD.n7136 0.0380882
R45730 PAD.n7596 PAD.n7592 0.0380882
R45731 PAD.n7592 PAD.n7588 0.0380882
R45732 PAD.n7588 PAD.n7138 0.0380882
R45733 PAD.n7584 PAD.n7138 0.0380882
R45734 PAD.n7584 PAD.n7580 0.0380882
R45735 PAD.n7580 PAD.n7576 0.0380882
R45736 PAD.n7576 PAD.n7140 0.0380882
R45737 PAD.n7572 PAD.n7140 0.0380882
R45738 PAD.n7572 PAD.n7568 0.0380882
R45739 PAD.n7568 PAD.n7564 0.0380882
R45740 PAD.n7564 PAD.n7142 0.0380882
R45741 PAD.n7560 PAD.n7142 0.0380882
R45742 PAD.n7560 PAD.n7556 0.0380882
R45743 PAD.n7556 PAD.n7552 0.0380882
R45744 PAD.n7552 PAD.n7144 0.0380882
R45745 PAD.n7548 PAD.n7144 0.0380882
R45746 PAD.n7548 PAD.n7544 0.0380882
R45747 PAD.n7544 PAD.n7540 0.0380882
R45748 PAD.n7540 PAD.n7146 0.0380882
R45749 PAD.n7536 PAD.n7146 0.0380882
R45750 PAD.n7536 PAD.n7532 0.0380882
R45751 PAD.n7778 PAD.n7777 0.0380882
R45752 PAD.n7777 PAD.n7776 0.0380882
R45753 PAD.n7776 PAD.n7107 0.0380882
R45754 PAD.n7767 PAD.n7107 0.0380882
R45755 PAD.n7767 PAD.n7766 0.0380882
R45756 PAD.n7766 PAD.n7765 0.0380882
R45757 PAD.n7765 PAD.n7109 0.0380882
R45758 PAD.n7755 PAD.n7109 0.0380882
R45759 PAD.n7755 PAD.n7754 0.0380882
R45760 PAD.n7754 PAD.n7753 0.0380882
R45761 PAD.n7753 PAD.n7111 0.0380882
R45762 PAD.n7743 PAD.n7111 0.0380882
R45763 PAD.n7743 PAD.n7742 0.0380882
R45764 PAD.n7742 PAD.n7741 0.0380882
R45765 PAD.n7741 PAD.n7113 0.0380882
R45766 PAD.n7731 PAD.n7113 0.0380882
R45767 PAD.n7731 PAD.n7730 0.0380882
R45768 PAD.n7730 PAD.n7729 0.0380882
R45769 PAD.n7729 PAD.n7115 0.0380882
R45770 PAD.n7719 PAD.n7115 0.0380882
R45771 PAD.n7719 PAD.n7718 0.0380882
R45772 PAD.n7718 PAD.n7717 0.0380882
R45773 PAD.n7717 PAD.n7117 0.0380882
R45774 PAD.n7707 PAD.n7117 0.0380882
R45775 PAD.n7707 PAD.n7706 0.0380882
R45776 PAD.n7706 PAD.n7705 0.0380882
R45777 PAD.n7705 PAD.n7119 0.0380882
R45778 PAD.n7695 PAD.n7119 0.0380882
R45779 PAD.n7695 PAD.n7694 0.0380882
R45780 PAD.n7694 PAD.n7693 0.0380882
R45781 PAD.n7693 PAD.n7121 0.0380882
R45782 PAD.n7683 PAD.n7121 0.0380882
R45783 PAD.n7683 PAD.n7682 0.0380882
R45784 PAD.n7682 PAD.n7681 0.0380882
R45785 PAD.n7681 PAD.n7123 0.0380882
R45786 PAD.n7671 PAD.n7123 0.0380882
R45787 PAD.n7671 PAD.n7670 0.0380882
R45788 PAD.n7670 PAD.n7669 0.0380882
R45789 PAD.n7669 PAD.n7125 0.0380882
R45790 PAD.n7659 PAD.n7125 0.0380882
R45791 PAD.n7659 PAD.n7658 0.0380882
R45792 PAD.n7658 PAD.n7657 0.0380882
R45793 PAD.n7657 PAD.n7127 0.0380882
R45794 PAD.n7647 PAD.n7127 0.0380882
R45795 PAD.n7647 PAD.n7646 0.0380882
R45796 PAD.n7646 PAD.n7645 0.0380882
R45797 PAD.n7645 PAD.n7129 0.0380882
R45798 PAD.n7635 PAD.n7129 0.0380882
R45799 PAD.n7635 PAD.n7634 0.0380882
R45800 PAD.n7634 PAD.n7633 0.0380882
R45801 PAD.n7633 PAD.n7131 0.0380882
R45802 PAD.n7623 PAD.n7131 0.0380882
R45803 PAD.n7623 PAD.n7622 0.0380882
R45804 PAD.n7622 PAD.n7621 0.0380882
R45805 PAD.n7621 PAD.n7133 0.0380882
R45806 PAD.n7611 PAD.n7133 0.0380882
R45807 PAD.n7611 PAD.n7610 0.0380882
R45808 PAD.n7610 PAD.n7609 0.0380882
R45809 PAD.n7609 PAD.n7135 0.0380882
R45810 PAD.n7599 PAD.n7135 0.0380882
R45811 PAD.n7599 PAD.n7598 0.0380882
R45812 PAD.n7598 PAD.n7597 0.0380882
R45813 PAD.n7597 PAD.n7137 0.0380882
R45814 PAD.n7587 PAD.n7137 0.0380882
R45815 PAD.n7587 PAD.n7586 0.0380882
R45816 PAD.n7586 PAD.n7585 0.0380882
R45817 PAD.n7585 PAD.n7139 0.0380882
R45818 PAD.n7575 PAD.n7139 0.0380882
R45819 PAD.n7575 PAD.n7574 0.0380882
R45820 PAD.n7574 PAD.n7573 0.0380882
R45821 PAD.n7573 PAD.n7141 0.0380882
R45822 PAD.n7563 PAD.n7141 0.0380882
R45823 PAD.n7563 PAD.n7562 0.0380882
R45824 PAD.n7562 PAD.n7561 0.0380882
R45825 PAD.n7561 PAD.n7143 0.0380882
R45826 PAD.n7551 PAD.n7143 0.0380882
R45827 PAD.n7551 PAD.n7550 0.0380882
R45828 PAD.n7550 PAD.n7549 0.0380882
R45829 PAD.n7549 PAD.n7145 0.0380882
R45830 PAD.n7539 PAD.n7145 0.0380882
R45831 PAD.n7539 PAD.n7538 0.0380882
R45832 PAD.n7538 PAD.n7537 0.0380882
R45833 PAD.n7537 PAD.n7147 0.0380882
R45834 PAD.n7050 PAD.n7049 0.0380882
R45835 PAD.n7049 PAD.n6720 0.0380882
R45836 PAD.n7043 PAD.n6720 0.0380882
R45837 PAD.n7043 PAD.n6723 0.0380882
R45838 PAD.n7039 PAD.n6723 0.0380882
R45839 PAD.n7039 PAD.n6726 0.0380882
R45840 PAD.n7031 PAD.n6726 0.0380882
R45841 PAD.n7031 PAD.n6728 0.0380882
R45842 PAD.n7027 PAD.n6728 0.0380882
R45843 PAD.n7027 PAD.n6730 0.0380882
R45844 PAD.n7019 PAD.n6730 0.0380882
R45845 PAD.n7019 PAD.n6732 0.0380882
R45846 PAD.n7015 PAD.n6732 0.0380882
R45847 PAD.n7015 PAD.n6734 0.0380882
R45848 PAD.n7007 PAD.n6734 0.0380882
R45849 PAD.n7007 PAD.n6736 0.0380882
R45850 PAD.n7003 PAD.n6736 0.0380882
R45851 PAD.n7003 PAD.n6738 0.0380882
R45852 PAD.n6995 PAD.n6738 0.0380882
R45853 PAD.n6995 PAD.n6740 0.0380882
R45854 PAD.n6991 PAD.n6740 0.0380882
R45855 PAD.n6991 PAD.n6742 0.0380882
R45856 PAD.n6983 PAD.n6742 0.0380882
R45857 PAD.n6983 PAD.n6744 0.0380882
R45858 PAD.n6979 PAD.n6744 0.0380882
R45859 PAD.n6979 PAD.n6746 0.0380882
R45860 PAD.n6971 PAD.n6746 0.0380882
R45861 PAD.n6971 PAD.n6748 0.0380882
R45862 PAD.n6967 PAD.n6748 0.0380882
R45863 PAD.n6967 PAD.n6750 0.0380882
R45864 PAD.n6959 PAD.n6750 0.0380882
R45865 PAD.n6959 PAD.n6752 0.0380882
R45866 PAD.n6955 PAD.n6752 0.0380882
R45867 PAD.n6955 PAD.n6754 0.0380882
R45868 PAD.n6947 PAD.n6754 0.0380882
R45869 PAD.n6947 PAD.n6756 0.0380882
R45870 PAD.n6943 PAD.n6756 0.0380882
R45871 PAD.n6943 PAD.n6758 0.0380882
R45872 PAD.n6935 PAD.n6758 0.0380882
R45873 PAD.n6935 PAD.n6760 0.0380882
R45874 PAD.n6931 PAD.n6760 0.0380882
R45875 PAD.n6931 PAD.n6762 0.0380882
R45876 PAD.n6923 PAD.n6762 0.0380882
R45877 PAD.n6923 PAD.n6764 0.0380882
R45878 PAD.n6919 PAD.n6764 0.0380882
R45879 PAD.n6919 PAD.n6766 0.0380882
R45880 PAD.n6911 PAD.n6766 0.0380882
R45881 PAD.n6911 PAD.n6768 0.0380882
R45882 PAD.n6907 PAD.n6768 0.0380882
R45883 PAD.n6907 PAD.n6770 0.0380882
R45884 PAD.n6899 PAD.n6770 0.0380882
R45885 PAD.n6899 PAD.n6772 0.0380882
R45886 PAD.n6895 PAD.n6772 0.0380882
R45887 PAD.n6895 PAD.n6774 0.0380882
R45888 PAD.n6887 PAD.n6774 0.0380882
R45889 PAD.n6887 PAD.n6776 0.0380882
R45890 PAD.n6883 PAD.n6776 0.0380882
R45891 PAD.n6883 PAD.n6778 0.0380882
R45892 PAD.n6875 PAD.n6778 0.0380882
R45893 PAD.n6875 PAD.n6780 0.0380882
R45894 PAD.n6871 PAD.n6780 0.0380882
R45895 PAD.n6871 PAD.n6782 0.0380882
R45896 PAD.n6863 PAD.n6782 0.0380882
R45897 PAD.n6863 PAD.n6784 0.0380882
R45898 PAD.n6859 PAD.n6784 0.0380882
R45899 PAD.n6859 PAD.n6786 0.0380882
R45900 PAD.n6851 PAD.n6786 0.0380882
R45901 PAD.n6851 PAD.n6788 0.0380882
R45902 PAD.n6847 PAD.n6788 0.0380882
R45903 PAD.n6847 PAD.n6790 0.0380882
R45904 PAD.n6839 PAD.n6790 0.0380882
R45905 PAD.n6839 PAD.n6792 0.0380882
R45906 PAD.n6835 PAD.n6792 0.0380882
R45907 PAD.n6835 PAD.n6794 0.0380882
R45908 PAD.n6827 PAD.n6794 0.0380882
R45909 PAD.n6827 PAD.n6796 0.0380882
R45910 PAD.n6823 PAD.n6796 0.0380882
R45911 PAD.n6823 PAD.n6798 0.0380882
R45912 PAD.n6815 PAD.n6798 0.0380882
R45913 PAD.n6815 PAD.n6800 0.0380882
R45914 PAD.n6811 PAD.n6800 0.0380882
R45915 PAD.n6811 PAD.n6802 0.0380882
R45916 PAD.n6803 PAD.n6802 0.0380882
R45917 PAD.n7051 PAD.n6718 0.0380882
R45918 PAD.n6724 PAD.n6718 0.0380882
R45919 PAD.n7042 PAD.n6724 0.0380882
R45920 PAD.n7042 PAD.n7041 0.0380882
R45921 PAD.n7041 PAD.n7040 0.0380882
R45922 PAD.n7040 PAD.n6725 0.0380882
R45923 PAD.n7030 PAD.n6725 0.0380882
R45924 PAD.n7030 PAD.n7029 0.0380882
R45925 PAD.n7029 PAD.n7028 0.0380882
R45926 PAD.n7028 PAD.n6729 0.0380882
R45927 PAD.n7018 PAD.n6729 0.0380882
R45928 PAD.n7018 PAD.n7017 0.0380882
R45929 PAD.n7017 PAD.n7016 0.0380882
R45930 PAD.n7016 PAD.n6733 0.0380882
R45931 PAD.n7006 PAD.n6733 0.0380882
R45932 PAD.n7006 PAD.n7005 0.0380882
R45933 PAD.n7005 PAD.n7004 0.0380882
R45934 PAD.n7004 PAD.n6737 0.0380882
R45935 PAD.n6994 PAD.n6737 0.0380882
R45936 PAD.n6994 PAD.n6993 0.0380882
R45937 PAD.n6993 PAD.n6992 0.0380882
R45938 PAD.n6992 PAD.n6741 0.0380882
R45939 PAD.n6982 PAD.n6741 0.0380882
R45940 PAD.n6982 PAD.n6981 0.0380882
R45941 PAD.n6981 PAD.n6980 0.0380882
R45942 PAD.n6980 PAD.n6745 0.0380882
R45943 PAD.n6970 PAD.n6745 0.0380882
R45944 PAD.n6970 PAD.n6969 0.0380882
R45945 PAD.n6969 PAD.n6968 0.0380882
R45946 PAD.n6968 PAD.n6749 0.0380882
R45947 PAD.n6958 PAD.n6749 0.0380882
R45948 PAD.n6958 PAD.n6957 0.0380882
R45949 PAD.n6957 PAD.n6956 0.0380882
R45950 PAD.n6956 PAD.n6753 0.0380882
R45951 PAD.n6946 PAD.n6753 0.0380882
R45952 PAD.n6946 PAD.n6945 0.0380882
R45953 PAD.n6945 PAD.n6944 0.0380882
R45954 PAD.n6944 PAD.n6757 0.0380882
R45955 PAD.n6934 PAD.n6757 0.0380882
R45956 PAD.n6934 PAD.n6933 0.0380882
R45957 PAD.n6933 PAD.n6932 0.0380882
R45958 PAD.n6932 PAD.n6761 0.0380882
R45959 PAD.n6922 PAD.n6761 0.0380882
R45960 PAD.n6922 PAD.n6921 0.0380882
R45961 PAD.n6921 PAD.n6920 0.0380882
R45962 PAD.n6920 PAD.n6765 0.0380882
R45963 PAD.n6910 PAD.n6765 0.0380882
R45964 PAD.n6910 PAD.n6909 0.0380882
R45965 PAD.n6909 PAD.n6908 0.0380882
R45966 PAD.n6908 PAD.n6769 0.0380882
R45967 PAD.n6898 PAD.n6769 0.0380882
R45968 PAD.n6898 PAD.n6897 0.0380882
R45969 PAD.n6897 PAD.n6896 0.0380882
R45970 PAD.n6896 PAD.n6773 0.0380882
R45971 PAD.n6886 PAD.n6773 0.0380882
R45972 PAD.n6886 PAD.n6885 0.0380882
R45973 PAD.n6885 PAD.n6884 0.0380882
R45974 PAD.n6884 PAD.n6777 0.0380882
R45975 PAD.n6874 PAD.n6777 0.0380882
R45976 PAD.n6874 PAD.n6873 0.0380882
R45977 PAD.n6873 PAD.n6872 0.0380882
R45978 PAD.n6872 PAD.n6781 0.0380882
R45979 PAD.n6862 PAD.n6781 0.0380882
R45980 PAD.n6862 PAD.n6861 0.0380882
R45981 PAD.n6861 PAD.n6860 0.0380882
R45982 PAD.n6860 PAD.n6785 0.0380882
R45983 PAD.n6850 PAD.n6785 0.0380882
R45984 PAD.n6850 PAD.n6849 0.0380882
R45985 PAD.n6849 PAD.n6848 0.0380882
R45986 PAD.n6848 PAD.n6789 0.0380882
R45987 PAD.n6838 PAD.n6789 0.0380882
R45988 PAD.n6838 PAD.n6837 0.0380882
R45989 PAD.n6837 PAD.n6836 0.0380882
R45990 PAD.n6836 PAD.n6793 0.0380882
R45991 PAD.n6826 PAD.n6793 0.0380882
R45992 PAD.n6826 PAD.n6825 0.0380882
R45993 PAD.n6825 PAD.n6824 0.0380882
R45994 PAD.n6824 PAD.n6797 0.0380882
R45995 PAD.n6814 PAD.n6797 0.0380882
R45996 PAD.n6814 PAD.n6813 0.0380882
R45997 PAD.n6813 PAD.n6812 0.0380882
R45998 PAD.n6812 PAD.n6801 0.0380882
R45999 PAD.n6801 PAD.n6705 0.0380882
R46000 PAD.n5891 PAD.n5890 0.0380882
R46001 PAD.n5890 PAD.n5605 0.0380882
R46002 PAD.n5886 PAD.n5605 0.0380882
R46003 PAD.n5886 PAD.n5882 0.0380882
R46004 PAD.n5882 PAD.n5881 0.0380882
R46005 PAD.n5881 PAD.n5607 0.0380882
R46006 PAD.n5877 PAD.n5607 0.0380882
R46007 PAD.n5877 PAD.n5873 0.0380882
R46008 PAD.n5873 PAD.n5872 0.0380882
R46009 PAD.n5872 PAD.n5612 0.0380882
R46010 PAD.n5868 PAD.n5612 0.0380882
R46011 PAD.n5868 PAD.n5864 0.0380882
R46012 PAD.n5864 PAD.n5863 0.0380882
R46013 PAD.n5863 PAD.n5617 0.0380882
R46014 PAD.n5859 PAD.n5617 0.0380882
R46015 PAD.n5859 PAD.n5855 0.0380882
R46016 PAD.n5855 PAD.n5854 0.0380882
R46017 PAD.n5854 PAD.n5622 0.0380882
R46018 PAD.n5850 PAD.n5622 0.0380882
R46019 PAD.n5850 PAD.n5846 0.0380882
R46020 PAD.n5846 PAD.n5845 0.0380882
R46021 PAD.n5845 PAD.n5627 0.0380882
R46022 PAD.n5841 PAD.n5627 0.0380882
R46023 PAD.n5841 PAD.n5837 0.0380882
R46024 PAD.n5837 PAD.n5836 0.0380882
R46025 PAD.n5836 PAD.n5632 0.0380882
R46026 PAD.n5832 PAD.n5632 0.0380882
R46027 PAD.n5832 PAD.n5828 0.0380882
R46028 PAD.n5828 PAD.n5827 0.0380882
R46029 PAD.n5827 PAD.n5637 0.0380882
R46030 PAD.n5823 PAD.n5637 0.0380882
R46031 PAD.n5823 PAD.n5819 0.0380882
R46032 PAD.n5819 PAD.n5818 0.0380882
R46033 PAD.n5818 PAD.n5642 0.0380882
R46034 PAD.n5814 PAD.n5642 0.0380882
R46035 PAD.n5814 PAD.n5810 0.0380882
R46036 PAD.n5810 PAD.n5809 0.0380882
R46037 PAD.n5809 PAD.n5647 0.0380882
R46038 PAD.n5805 PAD.n5647 0.0380882
R46039 PAD.n5805 PAD.n5801 0.0380882
R46040 PAD.n5801 PAD.n5800 0.0380882
R46041 PAD.n5800 PAD.n5652 0.0380882
R46042 PAD.n5796 PAD.n5652 0.0380882
R46043 PAD.n5796 PAD.n5792 0.0380882
R46044 PAD.n5792 PAD.n5791 0.0380882
R46045 PAD.n5791 PAD.n5657 0.0380882
R46046 PAD.n5787 PAD.n5657 0.0380882
R46047 PAD.n5787 PAD.n5783 0.0380882
R46048 PAD.n5783 PAD.n5782 0.0380882
R46049 PAD.n5782 PAD.n5662 0.0380882
R46050 PAD.n5778 PAD.n5662 0.0380882
R46051 PAD.n5778 PAD.n5774 0.0380882
R46052 PAD.n5774 PAD.n5773 0.0380882
R46053 PAD.n5773 PAD.n5667 0.0380882
R46054 PAD.n5769 PAD.n5667 0.0380882
R46055 PAD.n5769 PAD.n5765 0.0380882
R46056 PAD.n5765 PAD.n5764 0.0380882
R46057 PAD.n5764 PAD.n5672 0.0380882
R46058 PAD.n5760 PAD.n5672 0.0380882
R46059 PAD.n5760 PAD.n5756 0.0380882
R46060 PAD.n5756 PAD.n5755 0.0380882
R46061 PAD.n5755 PAD.n5677 0.0380882
R46062 PAD.n5751 PAD.n5677 0.0380882
R46063 PAD.n5751 PAD.n5747 0.0380882
R46064 PAD.n5747 PAD.n5746 0.0380882
R46065 PAD.n5746 PAD.n5682 0.0380882
R46066 PAD.n5742 PAD.n5682 0.0380882
R46067 PAD.n5742 PAD.n5738 0.0380882
R46068 PAD.n5738 PAD.n5737 0.0380882
R46069 PAD.n5737 PAD.n5687 0.0380882
R46070 PAD.n5733 PAD.n5687 0.0380882
R46071 PAD.n5733 PAD.n5729 0.0380882
R46072 PAD.n5729 PAD.n5728 0.0380882
R46073 PAD.n5728 PAD.n5692 0.0380882
R46074 PAD.n5724 PAD.n5692 0.0380882
R46075 PAD.n5724 PAD.n5720 0.0380882
R46076 PAD.n5720 PAD.n5719 0.0380882
R46077 PAD.n5719 PAD.n5697 0.0380882
R46078 PAD.n5715 PAD.n5697 0.0380882
R46079 PAD.n5715 PAD.n5711 0.0380882
R46080 PAD.n5711 PAD.n5710 0.0380882
R46081 PAD.n5710 PAD.n5704 0.0380882
R46082 PAD.n5704 PAD.n5703 0.0380882
R46083 PAD.n5889 PAD.n5545 0.0380882
R46084 PAD.n5889 PAD.n5888 0.0380882
R46085 PAD.n5888 PAD.n5887 0.0380882
R46086 PAD.n5887 PAD.n5606 0.0380882
R46087 PAD.n5880 PAD.n5606 0.0380882
R46088 PAD.n5880 PAD.n5879 0.0380882
R46089 PAD.n5879 PAD.n5878 0.0380882
R46090 PAD.n5878 PAD.n5611 0.0380882
R46091 PAD.n5871 PAD.n5611 0.0380882
R46092 PAD.n5871 PAD.n5870 0.0380882
R46093 PAD.n5870 PAD.n5869 0.0380882
R46094 PAD.n5869 PAD.n5616 0.0380882
R46095 PAD.n5862 PAD.n5616 0.0380882
R46096 PAD.n5862 PAD.n5861 0.0380882
R46097 PAD.n5861 PAD.n5860 0.0380882
R46098 PAD.n5860 PAD.n5621 0.0380882
R46099 PAD.n5853 PAD.n5621 0.0380882
R46100 PAD.n5853 PAD.n5852 0.0380882
R46101 PAD.n5852 PAD.n5851 0.0380882
R46102 PAD.n5851 PAD.n5626 0.0380882
R46103 PAD.n5844 PAD.n5626 0.0380882
R46104 PAD.n5844 PAD.n5843 0.0380882
R46105 PAD.n5843 PAD.n5842 0.0380882
R46106 PAD.n5842 PAD.n5631 0.0380882
R46107 PAD.n5835 PAD.n5631 0.0380882
R46108 PAD.n5835 PAD.n5834 0.0380882
R46109 PAD.n5834 PAD.n5833 0.0380882
R46110 PAD.n5833 PAD.n5636 0.0380882
R46111 PAD.n5826 PAD.n5636 0.0380882
R46112 PAD.n5826 PAD.n5825 0.0380882
R46113 PAD.n5825 PAD.n5824 0.0380882
R46114 PAD.n5824 PAD.n5641 0.0380882
R46115 PAD.n5817 PAD.n5641 0.0380882
R46116 PAD.n5817 PAD.n5816 0.0380882
R46117 PAD.n5816 PAD.n5815 0.0380882
R46118 PAD.n5815 PAD.n5646 0.0380882
R46119 PAD.n5808 PAD.n5646 0.0380882
R46120 PAD.n5808 PAD.n5807 0.0380882
R46121 PAD.n5807 PAD.n5806 0.0380882
R46122 PAD.n5806 PAD.n5651 0.0380882
R46123 PAD.n5799 PAD.n5651 0.0380882
R46124 PAD.n5799 PAD.n5798 0.0380882
R46125 PAD.n5798 PAD.n5797 0.0380882
R46126 PAD.n5797 PAD.n5656 0.0380882
R46127 PAD.n5790 PAD.n5656 0.0380882
R46128 PAD.n5790 PAD.n5789 0.0380882
R46129 PAD.n5789 PAD.n5788 0.0380882
R46130 PAD.n5788 PAD.n5661 0.0380882
R46131 PAD.n5781 PAD.n5661 0.0380882
R46132 PAD.n5781 PAD.n5780 0.0380882
R46133 PAD.n5780 PAD.n5779 0.0380882
R46134 PAD.n5779 PAD.n5666 0.0380882
R46135 PAD.n5772 PAD.n5666 0.0380882
R46136 PAD.n5772 PAD.n5771 0.0380882
R46137 PAD.n5771 PAD.n5770 0.0380882
R46138 PAD.n5770 PAD.n5671 0.0380882
R46139 PAD.n5763 PAD.n5671 0.0380882
R46140 PAD.n5763 PAD.n5762 0.0380882
R46141 PAD.n5762 PAD.n5761 0.0380882
R46142 PAD.n5761 PAD.n5676 0.0380882
R46143 PAD.n5754 PAD.n5676 0.0380882
R46144 PAD.n5754 PAD.n5753 0.0380882
R46145 PAD.n5753 PAD.n5752 0.0380882
R46146 PAD.n5752 PAD.n5681 0.0380882
R46147 PAD.n5745 PAD.n5681 0.0380882
R46148 PAD.n5745 PAD.n5744 0.0380882
R46149 PAD.n5744 PAD.n5743 0.0380882
R46150 PAD.n5743 PAD.n5686 0.0380882
R46151 PAD.n5736 PAD.n5686 0.0380882
R46152 PAD.n5736 PAD.n5735 0.0380882
R46153 PAD.n5735 PAD.n5734 0.0380882
R46154 PAD.n5734 PAD.n5691 0.0380882
R46155 PAD.n5727 PAD.n5691 0.0380882
R46156 PAD.n5727 PAD.n5726 0.0380882
R46157 PAD.n5726 PAD.n5725 0.0380882
R46158 PAD.n5725 PAD.n5696 0.0380882
R46159 PAD.n5718 PAD.n5696 0.0380882
R46160 PAD.n5718 PAD.n5717 0.0380882
R46161 PAD.n5717 PAD.n5716 0.0380882
R46162 PAD.n5716 PAD.n5701 0.0380882
R46163 PAD.n5709 PAD.n5701 0.0380882
R46164 PAD.n5709 PAD.n5708 0.0380882
R46165 PAD.n5708 PAD.n5557 0.0380882
R46166 PAD.n11087 PAD.n10747 0.0380882
R46167 PAD.n11079 PAD.n10747 0.0380882
R46168 PAD.n11079 PAD.n11078 0.0380882
R46169 PAD.n11078 PAD.n11077 0.0380882
R46170 PAD.n11077 PAD.n10758 0.0380882
R46171 PAD.n11067 PAD.n10758 0.0380882
R46172 PAD.n11067 PAD.n11066 0.0380882
R46173 PAD.n11066 PAD.n11065 0.0380882
R46174 PAD.n11065 PAD.n10762 0.0380882
R46175 PAD.n11055 PAD.n10762 0.0380882
R46176 PAD.n11055 PAD.n11054 0.0380882
R46177 PAD.n11054 PAD.n11053 0.0380882
R46178 PAD.n11053 PAD.n10766 0.0380882
R46179 PAD.n11043 PAD.n10766 0.0380882
R46180 PAD.n11043 PAD.n11042 0.0380882
R46181 PAD.n11042 PAD.n11041 0.0380882
R46182 PAD.n11041 PAD.n10770 0.0380882
R46183 PAD.n11031 PAD.n10770 0.0380882
R46184 PAD.n11031 PAD.n11030 0.0380882
R46185 PAD.n11030 PAD.n11029 0.0380882
R46186 PAD.n11029 PAD.n10774 0.0380882
R46187 PAD.n11019 PAD.n10774 0.0380882
R46188 PAD.n11019 PAD.n11018 0.0380882
R46189 PAD.n11018 PAD.n11017 0.0380882
R46190 PAD.n11017 PAD.n10778 0.0380882
R46191 PAD.n11007 PAD.n10778 0.0380882
R46192 PAD.n11007 PAD.n11006 0.0380882
R46193 PAD.n11006 PAD.n11005 0.0380882
R46194 PAD.n11005 PAD.n10782 0.0380882
R46195 PAD.n10995 PAD.n10782 0.0380882
R46196 PAD.n10995 PAD.n10994 0.0380882
R46197 PAD.n10994 PAD.n10993 0.0380882
R46198 PAD.n10993 PAD.n10786 0.0380882
R46199 PAD.n10983 PAD.n10786 0.0380882
R46200 PAD.n10983 PAD.n10982 0.0380882
R46201 PAD.n10982 PAD.n10981 0.0380882
R46202 PAD.n10981 PAD.n10790 0.0380882
R46203 PAD.n10971 PAD.n10790 0.0380882
R46204 PAD.n10971 PAD.n10970 0.0380882
R46205 PAD.n10970 PAD.n10969 0.0380882
R46206 PAD.n10969 PAD.n10794 0.0380882
R46207 PAD.n10959 PAD.n10794 0.0380882
R46208 PAD.n10959 PAD.n10958 0.0380882
R46209 PAD.n10958 PAD.n10957 0.0380882
R46210 PAD.n10957 PAD.n10798 0.0380882
R46211 PAD.n10947 PAD.n10798 0.0380882
R46212 PAD.n10947 PAD.n10946 0.0380882
R46213 PAD.n10946 PAD.n10945 0.0380882
R46214 PAD.n10945 PAD.n10802 0.0380882
R46215 PAD.n10935 PAD.n10802 0.0380882
R46216 PAD.n10935 PAD.n10934 0.0380882
R46217 PAD.n10934 PAD.n10933 0.0380882
R46218 PAD.n10933 PAD.n10806 0.0380882
R46219 PAD.n10923 PAD.n10806 0.0380882
R46220 PAD.n10923 PAD.n10922 0.0380882
R46221 PAD.n10922 PAD.n10921 0.0380882
R46222 PAD.n10921 PAD.n10810 0.0380882
R46223 PAD.n10911 PAD.n10810 0.0380882
R46224 PAD.n10911 PAD.n10910 0.0380882
R46225 PAD.n10910 PAD.n10909 0.0380882
R46226 PAD.n10909 PAD.n10814 0.0380882
R46227 PAD.n10899 PAD.n10814 0.0380882
R46228 PAD.n10899 PAD.n10898 0.0380882
R46229 PAD.n10898 PAD.n10897 0.0380882
R46230 PAD.n10897 PAD.n10818 0.0380882
R46231 PAD.n10887 PAD.n10818 0.0380882
R46232 PAD.n10887 PAD.n10886 0.0380882
R46233 PAD.n10886 PAD.n10885 0.0380882
R46234 PAD.n10885 PAD.n10822 0.0380882
R46235 PAD.n10875 PAD.n10822 0.0380882
R46236 PAD.n10875 PAD.n10874 0.0380882
R46237 PAD.n10874 PAD.n10873 0.0380882
R46238 PAD.n10873 PAD.n10826 0.0380882
R46239 PAD.n10863 PAD.n10826 0.0380882
R46240 PAD.n10863 PAD.n10862 0.0380882
R46241 PAD.n10862 PAD.n10861 0.0380882
R46242 PAD.n10861 PAD.n10830 0.0380882
R46243 PAD.n10851 PAD.n10830 0.0380882
R46244 PAD.n10851 PAD.n10850 0.0380882
R46245 PAD.n10850 PAD.n10849 0.0380882
R46246 PAD.n10849 PAD.n10834 0.0380882
R46247 PAD.n10839 PAD.n10834 0.0380882
R46248 PAD.n10839 PAD.n10734 0.0380882
R46249 PAD.n6692 PAD.n5898 0.0380882
R46250 PAD.n6499 PAD.n5898 0.0380882
R46251 PAD.n6500 PAD.n6499 0.0380882
R46252 PAD.n6501 PAD.n6500 0.0380882
R46253 PAD.n6501 PAD.n6494 0.0380882
R46254 PAD.n6508 PAD.n6494 0.0380882
R46255 PAD.n6509 PAD.n6508 0.0380882
R46256 PAD.n6510 PAD.n6509 0.0380882
R46257 PAD.n6510 PAD.n6491 0.0380882
R46258 PAD.n6517 PAD.n6491 0.0380882
R46259 PAD.n6518 PAD.n6517 0.0380882
R46260 PAD.n6519 PAD.n6518 0.0380882
R46261 PAD.n6519 PAD.n6488 0.0380882
R46262 PAD.n6526 PAD.n6488 0.0380882
R46263 PAD.n6527 PAD.n6526 0.0380882
R46264 PAD.n6528 PAD.n6527 0.0380882
R46265 PAD.n6528 PAD.n6485 0.0380882
R46266 PAD.n6535 PAD.n6485 0.0380882
R46267 PAD.n6536 PAD.n6535 0.0380882
R46268 PAD.n6537 PAD.n6536 0.0380882
R46269 PAD.n6537 PAD.n6482 0.0380882
R46270 PAD.n6544 PAD.n6482 0.0380882
R46271 PAD.n6545 PAD.n6544 0.0380882
R46272 PAD.n6546 PAD.n6545 0.0380882
R46273 PAD.n6546 PAD.n6479 0.0380882
R46274 PAD.n6553 PAD.n6479 0.0380882
R46275 PAD.n6554 PAD.n6553 0.0380882
R46276 PAD.n6555 PAD.n6554 0.0380882
R46277 PAD.n6555 PAD.n6476 0.0380882
R46278 PAD.n6562 PAD.n6476 0.0380882
R46279 PAD.n6563 PAD.n6562 0.0380882
R46280 PAD.n6564 PAD.n6563 0.0380882
R46281 PAD.n6564 PAD.n6473 0.0380882
R46282 PAD.n6571 PAD.n6473 0.0380882
R46283 PAD.n6572 PAD.n6571 0.0380882
R46284 PAD.n6573 PAD.n6572 0.0380882
R46285 PAD.n6573 PAD.n6470 0.0380882
R46286 PAD.n6580 PAD.n6470 0.0380882
R46287 PAD.n6581 PAD.n6580 0.0380882
R46288 PAD.n6582 PAD.n6581 0.0380882
R46289 PAD.n6582 PAD.n6467 0.0380882
R46290 PAD.n6589 PAD.n6467 0.0380882
R46291 PAD.n6590 PAD.n6589 0.0380882
R46292 PAD.n6591 PAD.n6590 0.0380882
R46293 PAD.n6591 PAD.n6464 0.0380882
R46294 PAD.n6598 PAD.n6464 0.0380882
R46295 PAD.n6599 PAD.n6598 0.0380882
R46296 PAD.n6600 PAD.n6599 0.0380882
R46297 PAD.n6600 PAD.n6461 0.0380882
R46298 PAD.n6607 PAD.n6461 0.0380882
R46299 PAD.n6608 PAD.n6607 0.0380882
R46300 PAD.n6609 PAD.n6608 0.0380882
R46301 PAD.n6609 PAD.n6458 0.0380882
R46302 PAD.n6616 PAD.n6458 0.0380882
R46303 PAD.n6617 PAD.n6616 0.0380882
R46304 PAD.n6618 PAD.n6617 0.0380882
R46305 PAD.n6618 PAD.n6455 0.0380882
R46306 PAD.n6625 PAD.n6455 0.0380882
R46307 PAD.n6626 PAD.n6625 0.0380882
R46308 PAD.n6627 PAD.n6626 0.0380882
R46309 PAD.n6627 PAD.n6452 0.0380882
R46310 PAD.n6634 PAD.n6452 0.0380882
R46311 PAD.n6635 PAD.n6634 0.0380882
R46312 PAD.n6636 PAD.n6635 0.0380882
R46313 PAD.n6636 PAD.n6449 0.0380882
R46314 PAD.n6643 PAD.n6449 0.0380882
R46315 PAD.n6644 PAD.n6643 0.0380882
R46316 PAD.n6645 PAD.n6644 0.0380882
R46317 PAD.n6645 PAD.n6446 0.0380882
R46318 PAD.n6652 PAD.n6446 0.0380882
R46319 PAD.n6653 PAD.n6652 0.0380882
R46320 PAD.n6654 PAD.n6653 0.0380882
R46321 PAD.n6654 PAD.n6443 0.0380882
R46322 PAD.n6661 PAD.n6443 0.0380882
R46323 PAD.n6662 PAD.n6661 0.0380882
R46324 PAD.n6663 PAD.n6662 0.0380882
R46325 PAD.n6663 PAD.n6440 0.0380882
R46326 PAD.n6670 PAD.n6440 0.0380882
R46327 PAD.n6671 PAD.n6670 0.0380882
R46328 PAD.n6674 PAD.n6671 0.0380882
R46329 PAD.n6674 PAD.n6673 0.0380882
R46330 PAD.n6673 PAD.n6672 0.0380882
R46331 PAD.n6672 PAD.n5951 0.0380882
R46332 PAD.n6691 PAD.n5900 0.0380882
R46333 PAD.n6498 PAD.n5900 0.0380882
R46334 PAD.n6498 PAD.n6496 0.0380882
R46335 PAD.n6503 PAD.n6496 0.0380882
R46336 PAD.n6505 PAD.n6503 0.0380882
R46337 PAD.n6507 PAD.n6505 0.0380882
R46338 PAD.n6507 PAD.n6493 0.0380882
R46339 PAD.n6512 PAD.n6493 0.0380882
R46340 PAD.n6514 PAD.n6512 0.0380882
R46341 PAD.n6516 PAD.n6514 0.0380882
R46342 PAD.n6516 PAD.n6490 0.0380882
R46343 PAD.n6521 PAD.n6490 0.0380882
R46344 PAD.n6523 PAD.n6521 0.0380882
R46345 PAD.n6525 PAD.n6523 0.0380882
R46346 PAD.n6525 PAD.n6487 0.0380882
R46347 PAD.n6530 PAD.n6487 0.0380882
R46348 PAD.n6532 PAD.n6530 0.0380882
R46349 PAD.n6534 PAD.n6532 0.0380882
R46350 PAD.n6534 PAD.n6484 0.0380882
R46351 PAD.n6539 PAD.n6484 0.0380882
R46352 PAD.n6541 PAD.n6539 0.0380882
R46353 PAD.n6543 PAD.n6541 0.0380882
R46354 PAD.n6543 PAD.n6481 0.0380882
R46355 PAD.n6548 PAD.n6481 0.0380882
R46356 PAD.n6550 PAD.n6548 0.0380882
R46357 PAD.n6552 PAD.n6550 0.0380882
R46358 PAD.n6552 PAD.n6478 0.0380882
R46359 PAD.n6557 PAD.n6478 0.0380882
R46360 PAD.n6559 PAD.n6557 0.0380882
R46361 PAD.n6561 PAD.n6559 0.0380882
R46362 PAD.n6561 PAD.n6475 0.0380882
R46363 PAD.n6566 PAD.n6475 0.0380882
R46364 PAD.n6568 PAD.n6566 0.0380882
R46365 PAD.n6570 PAD.n6568 0.0380882
R46366 PAD.n6570 PAD.n6472 0.0380882
R46367 PAD.n6575 PAD.n6472 0.0380882
R46368 PAD.n6577 PAD.n6575 0.0380882
R46369 PAD.n6579 PAD.n6577 0.0380882
R46370 PAD.n6579 PAD.n6469 0.0380882
R46371 PAD.n6584 PAD.n6469 0.0380882
R46372 PAD.n6586 PAD.n6584 0.0380882
R46373 PAD.n6588 PAD.n6586 0.0380882
R46374 PAD.n6588 PAD.n6466 0.0380882
R46375 PAD.n6593 PAD.n6466 0.0380882
R46376 PAD.n6595 PAD.n6593 0.0380882
R46377 PAD.n6597 PAD.n6595 0.0380882
R46378 PAD.n6597 PAD.n6463 0.0380882
R46379 PAD.n6602 PAD.n6463 0.0380882
R46380 PAD.n6604 PAD.n6602 0.0380882
R46381 PAD.n6606 PAD.n6604 0.0380882
R46382 PAD.n6606 PAD.n6460 0.0380882
R46383 PAD.n6611 PAD.n6460 0.0380882
R46384 PAD.n6613 PAD.n6611 0.0380882
R46385 PAD.n6615 PAD.n6613 0.0380882
R46386 PAD.n6615 PAD.n6457 0.0380882
R46387 PAD.n6620 PAD.n6457 0.0380882
R46388 PAD.n6622 PAD.n6620 0.0380882
R46389 PAD.n6624 PAD.n6622 0.0380882
R46390 PAD.n6624 PAD.n6454 0.0380882
R46391 PAD.n6629 PAD.n6454 0.0380882
R46392 PAD.n6631 PAD.n6629 0.0380882
R46393 PAD.n6633 PAD.n6631 0.0380882
R46394 PAD.n6633 PAD.n6451 0.0380882
R46395 PAD.n6638 PAD.n6451 0.0380882
R46396 PAD.n6640 PAD.n6638 0.0380882
R46397 PAD.n6642 PAD.n6640 0.0380882
R46398 PAD.n6642 PAD.n6448 0.0380882
R46399 PAD.n6647 PAD.n6448 0.0380882
R46400 PAD.n6649 PAD.n6647 0.0380882
R46401 PAD.n6651 PAD.n6649 0.0380882
R46402 PAD.n6651 PAD.n6445 0.0380882
R46403 PAD.n6656 PAD.n6445 0.0380882
R46404 PAD.n6658 PAD.n6656 0.0380882
R46405 PAD.n6660 PAD.n6658 0.0380882
R46406 PAD.n6660 PAD.n6442 0.0380882
R46407 PAD.n6665 PAD.n6442 0.0380882
R46408 PAD.n6667 PAD.n6665 0.0380882
R46409 PAD.n6669 PAD.n6667 0.0380882
R46410 PAD.n6669 PAD.n6438 0.0380882
R46411 PAD.n6675 PAD.n6438 0.0380882
R46412 PAD.n6675 PAD.n6439 0.0380882
R46413 PAD.n6439 PAD.n5950 0.0380882
R46414 PAD.n6687 PAD.n5950 0.0380882
R46415 PAD.n119 PAD.n118 0.0380882
R46416 PAD.n123 PAD.n118 0.0380882
R46417 PAD.n127 PAD.n123 0.0380882
R46418 PAD.n131 PAD.n127 0.0380882
R46419 PAD.n131 PAD.n114 0.0380882
R46420 PAD.n135 PAD.n114 0.0380882
R46421 PAD.n139 PAD.n135 0.0380882
R46422 PAD.n143 PAD.n139 0.0380882
R46423 PAD.n143 PAD.n112 0.0380882
R46424 PAD.n147 PAD.n112 0.0380882
R46425 PAD.n151 PAD.n147 0.0380882
R46426 PAD.n155 PAD.n151 0.0380882
R46427 PAD.n155 PAD.n110 0.0380882
R46428 PAD.n159 PAD.n110 0.0380882
R46429 PAD.n163 PAD.n159 0.0380882
R46430 PAD.n167 PAD.n163 0.0380882
R46431 PAD.n167 PAD.n108 0.0380882
R46432 PAD.n171 PAD.n108 0.0380882
R46433 PAD.n175 PAD.n171 0.0380882
R46434 PAD.n179 PAD.n175 0.0380882
R46435 PAD.n179 PAD.n106 0.0380882
R46436 PAD.n183 PAD.n106 0.0380882
R46437 PAD.n187 PAD.n183 0.0380882
R46438 PAD.n191 PAD.n187 0.0380882
R46439 PAD.n191 PAD.n104 0.0380882
R46440 PAD.n195 PAD.n104 0.0380882
R46441 PAD.n199 PAD.n195 0.0380882
R46442 PAD.n203 PAD.n199 0.0380882
R46443 PAD.n203 PAD.n102 0.0380882
R46444 PAD.n207 PAD.n102 0.0380882
R46445 PAD.n211 PAD.n207 0.0380882
R46446 PAD.n215 PAD.n211 0.0380882
R46447 PAD.n215 PAD.n100 0.0380882
R46448 PAD.n219 PAD.n100 0.0380882
R46449 PAD.n223 PAD.n219 0.0380882
R46450 PAD.n227 PAD.n223 0.0380882
R46451 PAD.n227 PAD.n98 0.0380882
R46452 PAD.n231 PAD.n98 0.0380882
R46453 PAD.n235 PAD.n231 0.0380882
R46454 PAD.n239 PAD.n235 0.0380882
R46455 PAD.n239 PAD.n96 0.0380882
R46456 PAD.n243 PAD.n96 0.0380882
R46457 PAD.n247 PAD.n243 0.0380882
R46458 PAD.n251 PAD.n247 0.0380882
R46459 PAD.n251 PAD.n94 0.0380882
R46460 PAD.n255 PAD.n94 0.0380882
R46461 PAD.n259 PAD.n255 0.0380882
R46462 PAD.n263 PAD.n259 0.0380882
R46463 PAD.n263 PAD.n92 0.0380882
R46464 PAD.n267 PAD.n92 0.0380882
R46465 PAD.n271 PAD.n267 0.0380882
R46466 PAD.n275 PAD.n271 0.0380882
R46467 PAD.n275 PAD.n90 0.0380882
R46468 PAD.n279 PAD.n90 0.0380882
R46469 PAD.n283 PAD.n279 0.0380882
R46470 PAD.n287 PAD.n283 0.0380882
R46471 PAD.n287 PAD.n88 0.0380882
R46472 PAD.n291 PAD.n88 0.0380882
R46473 PAD.n295 PAD.n291 0.0380882
R46474 PAD.n299 PAD.n295 0.0380882
R46475 PAD.n299 PAD.n86 0.0380882
R46476 PAD.n303 PAD.n86 0.0380882
R46477 PAD.n307 PAD.n303 0.0380882
R46478 PAD.n311 PAD.n307 0.0380882
R46479 PAD.n311 PAD.n84 0.0380882
R46480 PAD.n315 PAD.n84 0.0380882
R46481 PAD.n319 PAD.n315 0.0380882
R46482 PAD.n323 PAD.n319 0.0380882
R46483 PAD.n323 PAD.n82 0.0380882
R46484 PAD.n327 PAD.n82 0.0380882
R46485 PAD.n331 PAD.n327 0.0380882
R46486 PAD.n335 PAD.n331 0.0380882
R46487 PAD.n335 PAD.n80 0.0380882
R46488 PAD.n339 PAD.n80 0.0380882
R46489 PAD.n343 PAD.n339 0.0380882
R46490 PAD.n347 PAD.n343 0.0380882
R46491 PAD.n347 PAD.n78 0.0380882
R46492 PAD.n351 PAD.n78 0.0380882
R46493 PAD.n355 PAD.n351 0.0380882
R46494 PAD.n359 PAD.n355 0.0380882
R46495 PAD.n359 PAD.n76 0.0380882
R46496 PAD.n363 PAD.n76 0.0380882
R46497 PAD.n363 PAD.n75 0.0380882
R46498 PAD.n11086 PAD.n10749 0.0380882
R46499 PAD.n11080 PAD.n10749 0.0380882
R46500 PAD.n11080 PAD.n10757 0.0380882
R46501 PAD.n11076 PAD.n10757 0.0380882
R46502 PAD.n11076 PAD.n10759 0.0380882
R46503 PAD.n11068 PAD.n10759 0.0380882
R46504 PAD.n11068 PAD.n10761 0.0380882
R46505 PAD.n11064 PAD.n10761 0.0380882
R46506 PAD.n11064 PAD.n10763 0.0380882
R46507 PAD.n11056 PAD.n10763 0.0380882
R46508 PAD.n11056 PAD.n10765 0.0380882
R46509 PAD.n11052 PAD.n10765 0.0380882
R46510 PAD.n11052 PAD.n10767 0.0380882
R46511 PAD.n11044 PAD.n10767 0.0380882
R46512 PAD.n11044 PAD.n10769 0.0380882
R46513 PAD.n11040 PAD.n10769 0.0380882
R46514 PAD.n11040 PAD.n10771 0.0380882
R46515 PAD.n11032 PAD.n10771 0.0380882
R46516 PAD.n11032 PAD.n10773 0.0380882
R46517 PAD.n11028 PAD.n10773 0.0380882
R46518 PAD.n11028 PAD.n10775 0.0380882
R46519 PAD.n11020 PAD.n10775 0.0380882
R46520 PAD.n11020 PAD.n10777 0.0380882
R46521 PAD.n11016 PAD.n10777 0.0380882
R46522 PAD.n11016 PAD.n10779 0.0380882
R46523 PAD.n11008 PAD.n10779 0.0380882
R46524 PAD.n11008 PAD.n10781 0.0380882
R46525 PAD.n11004 PAD.n10781 0.0380882
R46526 PAD.n11004 PAD.n10783 0.0380882
R46527 PAD.n10996 PAD.n10783 0.0380882
R46528 PAD.n10996 PAD.n10785 0.0380882
R46529 PAD.n10992 PAD.n10785 0.0380882
R46530 PAD.n10992 PAD.n10787 0.0380882
R46531 PAD.n10984 PAD.n10787 0.0380882
R46532 PAD.n10984 PAD.n10789 0.0380882
R46533 PAD.n10980 PAD.n10789 0.0380882
R46534 PAD.n10980 PAD.n10791 0.0380882
R46535 PAD.n10972 PAD.n10791 0.0380882
R46536 PAD.n10972 PAD.n10793 0.0380882
R46537 PAD.n10968 PAD.n10793 0.0380882
R46538 PAD.n10968 PAD.n10795 0.0380882
R46539 PAD.n10960 PAD.n10795 0.0380882
R46540 PAD.n10960 PAD.n10797 0.0380882
R46541 PAD.n10956 PAD.n10797 0.0380882
R46542 PAD.n10956 PAD.n10799 0.0380882
R46543 PAD.n10948 PAD.n10799 0.0380882
R46544 PAD.n10948 PAD.n10801 0.0380882
R46545 PAD.n10944 PAD.n10801 0.0380882
R46546 PAD.n10944 PAD.n10803 0.0380882
R46547 PAD.n10936 PAD.n10803 0.0380882
R46548 PAD.n10936 PAD.n10805 0.0380882
R46549 PAD.n10932 PAD.n10805 0.0380882
R46550 PAD.n10932 PAD.n10807 0.0380882
R46551 PAD.n10924 PAD.n10807 0.0380882
R46552 PAD.n10924 PAD.n10809 0.0380882
R46553 PAD.n10920 PAD.n10809 0.0380882
R46554 PAD.n10920 PAD.n10811 0.0380882
R46555 PAD.n10912 PAD.n10811 0.0380882
R46556 PAD.n10912 PAD.n10813 0.0380882
R46557 PAD.n10908 PAD.n10813 0.0380882
R46558 PAD.n10908 PAD.n10815 0.0380882
R46559 PAD.n10900 PAD.n10815 0.0380882
R46560 PAD.n10900 PAD.n10817 0.0380882
R46561 PAD.n10896 PAD.n10817 0.0380882
R46562 PAD.n10896 PAD.n10819 0.0380882
R46563 PAD.n10888 PAD.n10819 0.0380882
R46564 PAD.n10888 PAD.n10821 0.0380882
R46565 PAD.n10884 PAD.n10821 0.0380882
R46566 PAD.n10884 PAD.n10823 0.0380882
R46567 PAD.n10876 PAD.n10823 0.0380882
R46568 PAD.n10876 PAD.n10825 0.0380882
R46569 PAD.n10872 PAD.n10825 0.0380882
R46570 PAD.n10872 PAD.n10827 0.0380882
R46571 PAD.n10864 PAD.n10827 0.0380882
R46572 PAD.n10864 PAD.n10829 0.0380882
R46573 PAD.n10860 PAD.n10829 0.0380882
R46574 PAD.n10860 PAD.n10831 0.0380882
R46575 PAD.n10852 PAD.n10831 0.0380882
R46576 PAD.n10852 PAD.n10833 0.0380882
R46577 PAD.n10848 PAD.n10833 0.0380882
R46578 PAD.n10848 PAD.n10835 0.0380882
R46579 PAD.n10840 PAD.n10835 0.0380882
R46580 PAD.n10840 PAD.n10838 0.0380882
R46581 PAD.n7810 PAD.n3637 0.0368392
R46582 PAD.n9168 PAD.n12 0.035749
R46583 PAD.n0 PAD 0.0336535
R46584 PAD.n6380 PAD.n6379 0.03245
R46585 PAD.n6379 PAD.n6378 0.03245
R46586 PAD.n5953 PAD.n5558 0.03245
R46587 PAD.n6703 PAD.n5558 0.03245
R46588 PAD.n7798 PAD.n7797 0.03245
R46589 PAD.n7795 PAD.n6706 0.03245
R46590 PAD.n7153 PAD.n6706 0.03245
R46591 PAD.n7526 PAD.n7525 0.03245
R46592 PAD.n7525 PAD.n7524 0.03245
R46593 PAD.n7203 PAD.n5201 0.03245
R46594 PAD.n7823 PAD.n5201 0.03245
R46595 PAD.n7825 PAD.n5187 0.03245
R46596 PAD.n8178 PAD.n5187 0.03245
R46597 PAD.n8180 PAD.n4836 0.03245
R46598 PAD.n8198 PAD.n4836 0.03245
R46599 PAD.n8200 PAD.n4830 0.03245
R46600 PAD.n8208 PAD.n4670 0.03245
R46601 PAD.n8413 PAD.n4670 0.03245
R46602 PAD.n8416 PAD.n8415 0.03245
R46603 PAD.n8415 PAD.n4315 0.03245
R46604 PAD.n8436 PAD.n4316 0.03245
R46605 PAD.n4316 PAD.n3974 0.03245
R46606 PAD.n8460 PAD.n3629 0.03245
R46607 PAD.n8483 PAD.n3629 0.03245
R46608 PAD.n8484 PAD.n3284 0.03245
R46609 PAD.n8509 PAD.n2899 0.03245
R46610 PAD.n8825 PAD.n2899 0.03245
R46611 PAD.n8828 PAD.n8827 0.03245
R46612 PAD.n8828 PAD.n2882 0.03245
R46613 PAD.n9132 PAD.n2491 0.03245
R46614 PAD.n9155 PAD.n2491 0.03245
R46615 PAD.n9157 PAD.n2143 0.03245
R46616 PAD.n9179 PAD.n2143 0.03245
R46617 PAD.n9181 PAD.n2041 0.03245
R46618 PAD.n9449 PAD.n2041 0.03245
R46619 PAD.n9452 PAD.n9451 0.03245
R46620 PAD.n9717 PAD.n9716 0.03245
R46621 PAD.n9718 PAD.n9717 0.03245
R46622 PAD.n9737 PAD.n9736 0.03245
R46623 PAD.n9738 PAD.n9737 0.03245
R46624 PAD.n10003 PAD.n10002 0.03245
R46625 PAD.n10004 PAD.n10003 0.03245
R46626 PAD.n10021 PAD.n10020 0.03245
R46627 PAD.n10358 PAD.n10021 0.03245
R46628 PAD.n10356 PAD.n1115 0.03245
R46629 PAD.n10380 PAD.n773 0.03245
R46630 PAD.n10401 PAD.n773 0.03245
R46631 PAD.n10404 PAD.n10403 0.03245
R46632 PAD.n10403 PAD.n422 0.03245
R46633 PAD.n10708 PAD.n27 0.03245
R46634 PAD.n10731 PAD.n27 0.03245
R46635 PAD.n11529 PAD.n10733 0.03245
R46636 PAD.n11529 PAD.n11528 0.03245
R46637 PAD.n11526 PAD.n10735 0.03245
R46638 PAD.n11504 PAD.n10735 0.03245
R46639 PAD.n7797 PAD.n7796 0.031775
R46640 PAD.n7516 PAD.n7227 0.0317353
R46641 PAD.n120 PAD.n14 0.0317353
R46642 PAD.n10697 PAD.n10696 0.0317353
R46643 PAD.n521 PAD.n430 0.0317353
R46644 PAD.n873 PAD.n779 0.0317353
R46645 PAD.n10367 PAD.n1124 0.0317353
R46646 PAD.n10012 PAD.n1145 0.0317353
R46647 PAD.n9750 PAD.n1580 0.0317353
R46648 PAD.n9726 PAD.n1932 0.0317353
R46649 PAD.n9464 PAD.n2032 0.0317353
R46650 PAD.n9198 PAD.n2135 0.0317353
R46651 PAD.n9167 PAD.n2483 0.0317353
R46652 PAD.n9147 PAD.n2830 0.0317353
R46653 PAD.n9124 PAD.n9120 0.0317353
R46654 PAD.n8817 PAD.n2888 0.0317353
R46655 PAD.n3042 PAD.n2949 0.0317353
R46656 PAD.n3387 PAD.n3293 0.0317353
R46657 PAD.n3732 PAD.n3638 0.0317353
R46658 PAD.n4073 PAD.n3980 0.0317353
R46659 PAD.n8424 PAD.n4325 0.0317353
R46660 PAD.n8402 PAD.n4676 0.0317353
R46661 PAD.n8190 PAD.n5179 0.0317353
R46662 PAD.n8170 PAD.n5193 0.0317353
R46663 PAD.n7815 PAD.n5543 0.0317353
R46664 PAD.n7778 PAD.n7056 0.0317353
R46665 PAD.n7055 PAD.n7051 0.0317353
R46666 PAD.n7806 PAD.n5545 0.0317353
R46667 PAD.n11088 PAD.n11087 0.0317353
R46668 PAD.n6693 PAD.n6692 0.0317353
R46669 PAD.n8510 PAD.n3284 0.031325
R46670 PAD.n9451 PAD.n9450 0.030875
R46671 PAD.n10381 PAD.n1115 0.030875
R46672 PAD.n8200 PAD.n8199 0.030425
R46673 PAD.n8209 PAD.n4830 0.028625
R46674 PAD.n6381 PAD.n5977 0.0284039
R46675 PAD.n5977 PAD.n5952 0.0284039
R46676 PAD.n6685 PAD.n5559 0.0284039
R46677 PAD.n6702 PAD.n5559 0.0284039
R46678 PAD.n7799 PAD.n5556 0.0284039
R46679 PAD.n7794 PAD.n6708 0.0284039
R46680 PAD.n7152 PAD.n6708 0.0284039
R46681 PAD.n7527 PAD.n7151 0.0284039
R46682 PAD.n7523 PAD.n7151 0.0284039
R46683 PAD.n7204 PAD.n5202 0.0284039
R46684 PAD.n7822 PAD.n5202 0.0284039
R46685 PAD.n7826 PAD.n5188 0.0284039
R46686 PAD.n8177 PAD.n5188 0.0284039
R46687 PAD.n8181 PAD.n4837 0.0284039
R46688 PAD.n8197 PAD.n4837 0.0284039
R46689 PAD.n8202 PAD.n8201 0.0284039
R46690 PAD.n8207 PAD.n4671 0.0284039
R46691 PAD.n8412 PAD.n4671 0.0284039
R46692 PAD.n8417 PAD.n4317 0.0284039
R46693 PAD.n8433 PAD.n4317 0.0284039
R46694 PAD.n8435 PAD.n3975 0.0284039
R46695 PAD.n8457 PAD.n3975 0.0284039
R46696 PAD.n8459 PAD.n3630 0.0284039
R46697 PAD.n8482 PAD.n3630 0.0284039
R46698 PAD.n8505 PAD.n3285 0.0284039
R46699 PAD.n8508 PAD.n2900 0.0284039
R46700 PAD.n8824 PAD.n2900 0.0284039
R46701 PAD.n8829 PAD.n2896 0.0284039
R46702 PAD.n8829 PAD.n2897 0.0284039
R46703 PAD.n9131 PAD.n2492 0.0284039
R46704 PAD.n9154 PAD.n2492 0.0284039
R46705 PAD.n9158 PAD.n2144 0.0284039
R46706 PAD.n9178 PAD.n2144 0.0284039
R46707 PAD.n9182 PAD.n2042 0.0284039
R46708 PAD.n9448 PAD.n2042 0.0284039
R46709 PAD.n9453 PAD.n2039 0.0284039
R46710 PAD.n9715 PAD.n1938 0.0284039
R46711 PAD.n9719 PAD.n1938 0.0284039
R46712 PAD.n9735 PAD.n1588 0.0284039
R46713 PAD.n9739 PAD.n1588 0.0284039
R46714 PAD.n10001 PAD.n1485 0.0284039
R46715 PAD.n10005 PAD.n1485 0.0284039
R46716 PAD.n10019 PAD.n1135 0.0284039
R46717 PAD.n10359 PAD.n1135 0.0284039
R46718 PAD.n10376 PAD.n1116 0.0284039
R46719 PAD.n10379 PAD.n774 0.0284039
R46720 PAD.n10400 PAD.n774 0.0284039
R46721 PAD.n10405 PAD.n423 0.0284039
R46722 PAD.n10704 PAD.n423 0.0284039
R46723 PAD.n10707 PAD.n28 0.0284039
R46724 PAD.n10730 PAD.n28 0.0284039
R46725 PAD.n11530 PAD.n24 0.0284039
R46726 PAD.n11530 PAD.n25 0.0284039
R46727 PAD.n11525 PAD.n10737 0.0284039
R46728 PAD.n11503 PAD.n10737 0.0284039
R46729 PAD.n6382 PAD.n5975 0.0284039
R46730 PAD.n5975 PAD.n5973 0.0284039
R46731 PAD.n6684 PAD.n5560 0.0284039
R46732 PAD.n6701 PAD.n5560 0.0284039
R46733 PAD.n7800 PAD.n5554 0.0284039
R46734 PAD.n7793 PAD.n6710 0.0284039
R46735 PAD.n7149 PAD.n6710 0.0284039
R46736 PAD.n7529 PAD.n7150 0.0284039
R46737 PAD.n7522 PAD.n7150 0.0284039
R46738 PAD.n7205 PAD.n5203 0.0284039
R46739 PAD.n7821 PAD.n5203 0.0284039
R46740 PAD.n7827 PAD.n5189 0.0284039
R46741 PAD.n8176 PAD.n5189 0.0284039
R46742 PAD.n8182 PAD.n4838 0.0284039
R46743 PAD.n8196 PAD.n4838 0.0284039
R46744 PAD.n8203 PAD.n4833 0.0284039
R46745 PAD.n8206 PAD.n4672 0.0284039
R46746 PAD.n8411 PAD.n4672 0.0284039
R46747 PAD.n8418 PAD.n4318 0.0284039
R46748 PAD.n8432 PAD.n4318 0.0284039
R46749 PAD.n8455 PAD.n3976 0.0284039
R46750 PAD.n8456 PAD.n8455 0.0284039
R46751 PAD.n8480 PAD.n3632 0.0284039
R46752 PAD.n8481 PAD.n8480 0.0284039
R46753 PAD.n8504 PAD.n3286 0.0284039
R46754 PAD.n8507 PAD.n2902 0.0284039
R46755 PAD.n8823 PAD.n2902 0.0284039
R46756 PAD.n8830 PAD.n2893 0.0284039
R46757 PAD.n8830 PAD.n2895 0.0284039
R46758 PAD.n9130 PAD.n2493 0.0284039
R46759 PAD.n9153 PAD.n2493 0.0284039
R46760 PAD.n9159 PAD.n2145 0.0284039
R46761 PAD.n9177 PAD.n2145 0.0284039
R46762 PAD.n9183 PAD.n2044 0.0284039
R46763 PAD.n9447 PAD.n2044 0.0284039
R46764 PAD.n9454 PAD.n2038 0.0284039
R46765 PAD.n9714 PAD.n1937 0.0284039
R46766 PAD.n9720 PAD.n1937 0.0284039
R46767 PAD.n9734 PAD.n1587 0.0284039
R46768 PAD.n9740 PAD.n1587 0.0284039
R46769 PAD.n10000 PAD.n1484 0.0284039
R46770 PAD.n10006 PAD.n1484 0.0284039
R46771 PAD.n10018 PAD.n1133 0.0284039
R46772 PAD.n10360 PAD.n1133 0.0284039
R46773 PAD.n10375 PAD.n1117 0.0284039
R46774 PAD.n10378 PAD.n775 0.0284039
R46775 PAD.n10399 PAD.n775 0.0284039
R46776 PAD.n10406 PAD.n424 0.0284039
R46777 PAD.n10703 PAD.n424 0.0284039
R46778 PAD.n10706 PAD.n30 0.0284039
R46779 PAD.n10729 PAD.n30 0.0284039
R46780 PAD.n11531 PAD.n22 0.0284039
R46781 PAD.n11531 PAD.n23 0.0284039
R46782 PAD.n11524 PAD.n10739 0.0284039
R46783 PAD.n11502 PAD.n10739 0.0284039
R46784 PAD.n9452 PAD.n1939 0.028175
R46785 PAD.n10357 PAD.n10356 0.028175
R46786 PAD.n6707 PAD.n5556 0.0278144
R46787 PAD.n6709 PAD.n5554 0.0278144
R46788 PAD.n8485 PAD.n8484 0.027725
R46789 PAD.n8506 PAD.n8505 0.0274214
R46790 PAD.n8504 PAD.n2996 0.0274214
R46791 PAD.n7798 PAD.n6704 0.027275
R46792 PAD.n2043 PAD.n2039 0.0270284
R46793 PAD.n10377 PAD.n10376 0.0270284
R46794 PAD.n2045 PAD.n2038 0.0270284
R46795 PAD.n10375 PAD.n827 0.0270284
R46796 PAD.n8201 PAD.n4834 0.0266354
R46797 PAD.n4839 PAD.n4833 0.0266354
R46798 PAD.n7154 PAD.n7153 0.025925
R46799 PAD.n7268 PAD.n7155 0.0259118
R46800 PAD.n10732 PAD.n26 0.0259118
R46801 PAD.n10710 PAD.n10709 0.0259118
R46802 PAD.n10402 PAD.n772 0.0259118
R46803 PAD.n10382 PAD.n10381 0.0259118
R46804 PAD.n10357 PAD.n10355 0.0259118
R46805 PAD.n1296 PAD.n1137 0.0259118
R46806 PAD.n9992 PAD.n1486 0.0259118
R46807 PAD.n1683 PAD.n1589 0.0259118
R46808 PAD.n9706 PAD.n1939 0.0259118
R46809 PAD.n9450 PAD.n2040 0.0259118
R46810 PAD.n9180 PAD.n2142 0.0259118
R46811 PAD.n9156 PAD.n2490 0.0259118
R46812 PAD.n9134 PAD.n9133 0.0259118
R46813 PAD.n8826 PAD.n2898 0.0259118
R46814 PAD.n8511 PAD.n8510 0.0259118
R46815 PAD.n8486 PAD.n8485 0.0259118
R46816 PAD.n8462 PAD.n8461 0.0259118
R46817 PAD.n8438 PAD.n8437 0.0259118
R46818 PAD.n8414 PAD.n4669 0.0259118
R46819 PAD.n8210 PAD.n8209 0.0259118
R46820 PAD.n8199 PAD.n4835 0.0259118
R46821 PAD.n8179 PAD.n5186 0.0259118
R46822 PAD.n7824 PAD.n5200 0.0259118
R46823 PAD.n7154 PAD.n7147 0.0259118
R46824 PAD.n7796 PAD.n6705 0.0259118
R46825 PAD.n6704 PAD.n5557 0.0259118
R46826 PAD.n11527 PAD.n10734 0.0259118
R46827 PAD.n6377 PAD.n5951 0.0259118
R46828 PAD.n8826 PAD.n8825 0.025475
R46829 PAD.n11527 PAD.n11526 0.025475
R46830 PAD.n11106 PAD.n11104 0.0251375
R46831 PAD.n11353 PAD.n11093 0.0251375
R46832 PAD.n11352 PAD.n11091 0.0251375
R46833 PAD.n6226 PAD.n5959 0.0251375
R46834 PAD.n6225 PAD.n5957 0.0251375
R46835 PAD.n6034 PAD.n5969 0.0251375
R46836 PAD.n8202 PAD.n4831 0.0250633
R46837 PAD.n8204 PAD.n8203 0.0250633
R46838 PAD.n9181 PAD.n9180 0.025025
R46839 PAD.n10402 PAD.n10401 0.025025
R46840 PAD.n9453 PAD.n1940 0.0246703
R46841 PAD.n1136 PAD.n1116 0.0246703
R46842 PAD.n9454 PAD.n1941 0.0246703
R46843 PAD.n1134 PAD.n1117 0.0246703
R46844 PAD.n8180 PAD.n8179 0.024575
R46845 PAD.n3631 PAD.n3285 0.0242773
R46846 PAD.n3341 PAD.n3286 0.0242773
R46847 PAD.n7799 PAD.n5555 0.0238843
R46848 PAD.n7800 PAD.n5553 0.0238843
R46849 PAD.n7811 PAD.n7808 0.0228122
R46850 PAD.n8414 PAD.n8413 0.022775
R46851 PAD.n7152 PAD.n7148 0.0227052
R46852 PAD.n7530 PAD.n7149 0.0227052
R46853 PAD.n9718 PAD.n1589 0.022325
R46854 PAD.n10020 PAD.n1137 0.022325
R46855 PAD.n8824 PAD.n2901 0.0223122
R46856 PAD.n11525 PAD.n10736 0.0223122
R46857 PAD.n8823 PAD.n2903 0.0223122
R46858 PAD.n11524 PAD.n10738 0.0223122
R46859 PAD.n13 PAD.n12 0.0221339
R46860 PAD.n9182 PAD.n2141 0.0219192
R46861 PAD.n10400 PAD.n437 0.0219192
R46862 PAD.n9183 PAD.n2140 0.0219192
R46863 PAD.n10399 PAD.n436 0.0219192
R46864 PAD.n8461 PAD.n8460 0.021875
R46865 PAD.n11539 PAD.n13 0.0216978
R46866 PAD.n8181 PAD.n5185 0.0215262
R46867 PAD.n8182 PAD.n5184 0.0215262
R46868 PAD.n6377 PAD.n5953 0.021425
R46869 PAD.n7811 PAD.n7810 0.0210195
R46870 PAD.n7524 PAD.n7155 0.020075
R46871 PAD.n8412 PAD.n4335 0.0199541
R46872 PAD.n8411 PAD.n4334 0.0199541
R46873 PAD.n117 PAD.n116 0.019716
R46874 PAD.n124 PAD.n73 0.019716
R46875 PAD.n125 PAD.n124 0.019716
R46876 PAD.n130 PAD.n72 0.019716
R46877 PAD.n130 PAD.n129 0.019716
R46878 PAD.n136 PAD.n71 0.019716
R46879 PAD.n137 PAD.n136 0.019716
R46880 PAD.n142 PAD.n70 0.019716
R46881 PAD.n142 PAD.n141 0.019716
R46882 PAD.n148 PAD.n69 0.019716
R46883 PAD.n149 PAD.n148 0.019716
R46884 PAD.n154 PAD.n68 0.019716
R46885 PAD.n154 PAD.n153 0.019716
R46886 PAD.n160 PAD.n67 0.019716
R46887 PAD.n161 PAD.n160 0.019716
R46888 PAD.n166 PAD.n66 0.019716
R46889 PAD.n166 PAD.n165 0.019716
R46890 PAD.n172 PAD.n65 0.019716
R46891 PAD.n173 PAD.n172 0.019716
R46892 PAD.n178 PAD.n64 0.019716
R46893 PAD.n178 PAD.n177 0.019716
R46894 PAD.n184 PAD.n63 0.019716
R46895 PAD.n185 PAD.n184 0.019716
R46896 PAD.n190 PAD.n62 0.019716
R46897 PAD.n190 PAD.n189 0.019716
R46898 PAD.n196 PAD.n61 0.019716
R46899 PAD.n197 PAD.n196 0.019716
R46900 PAD.n202 PAD.n60 0.019716
R46901 PAD.n202 PAD.n201 0.019716
R46902 PAD.n208 PAD.n59 0.019716
R46903 PAD.n209 PAD.n208 0.019716
R46904 PAD.n214 PAD.n58 0.019716
R46905 PAD.n214 PAD.n213 0.019716
R46906 PAD.n220 PAD.n57 0.019716
R46907 PAD.n221 PAD.n220 0.019716
R46908 PAD.n226 PAD.n56 0.019716
R46909 PAD.n226 PAD.n225 0.019716
R46910 PAD.n232 PAD.n55 0.019716
R46911 PAD.n233 PAD.n232 0.019716
R46912 PAD.n238 PAD.n54 0.019716
R46913 PAD.n238 PAD.n237 0.019716
R46914 PAD.n244 PAD.n53 0.019716
R46915 PAD.n245 PAD.n244 0.019716
R46916 PAD.n250 PAD.n52 0.019716
R46917 PAD.n250 PAD.n249 0.019716
R46918 PAD.n256 PAD.n51 0.019716
R46919 PAD.n257 PAD.n256 0.019716
R46920 PAD.n262 PAD.n50 0.019716
R46921 PAD.n262 PAD.n261 0.019716
R46922 PAD.n268 PAD.n49 0.019716
R46923 PAD.n269 PAD.n268 0.019716
R46924 PAD.n274 PAD.n48 0.019716
R46925 PAD.n274 PAD.n273 0.019716
R46926 PAD.n280 PAD.n47 0.019716
R46927 PAD.n281 PAD.n280 0.019716
R46928 PAD.n286 PAD.n46 0.019716
R46929 PAD.n286 PAD.n285 0.019716
R46930 PAD.n292 PAD.n45 0.019716
R46931 PAD.n293 PAD.n292 0.019716
R46932 PAD.n298 PAD.n44 0.019716
R46933 PAD.n298 PAD.n297 0.019716
R46934 PAD.n304 PAD.n43 0.019716
R46935 PAD.n305 PAD.n304 0.019716
R46936 PAD.n310 PAD.n42 0.019716
R46937 PAD.n310 PAD.n309 0.019716
R46938 PAD.n316 PAD.n41 0.019716
R46939 PAD.n317 PAD.n316 0.019716
R46940 PAD.n322 PAD.n40 0.019716
R46941 PAD.n322 PAD.n321 0.019716
R46942 PAD.n328 PAD.n39 0.019716
R46943 PAD.n329 PAD.n328 0.019716
R46944 PAD.n334 PAD.n38 0.019716
R46945 PAD.n334 PAD.n333 0.019716
R46946 PAD.n340 PAD.n37 0.019716
R46947 PAD.n341 PAD.n340 0.019716
R46948 PAD.n346 PAD.n36 0.019716
R46949 PAD.n346 PAD.n345 0.019716
R46950 PAD.n352 PAD.n35 0.019716
R46951 PAD.n353 PAD.n352 0.019716
R46952 PAD.n358 PAD.n34 0.019716
R46953 PAD.n358 PAD.n357 0.019716
R46954 PAD.n364 PAD.n33 0.019716
R46955 PAD.n365 PAD.n364 0.019716
R46956 PAD.n7519 PAD.n7201 0.019716
R46957 PAD.n7512 PAD.n7511 0.019716
R46958 PAD.n7512 PAD.n7199 0.019716
R46959 PAD.n7508 PAD.n7507 0.019716
R46960 PAD.n7507 PAD.n7198 0.019716
R46961 PAD.n7501 PAD.n7500 0.019716
R46962 PAD.n7501 PAD.n7197 0.019716
R46963 PAD.n7496 PAD.n7495 0.019716
R46964 PAD.n7495 PAD.n7196 0.019716
R46965 PAD.n7489 PAD.n7488 0.019716
R46966 PAD.n7489 PAD.n7195 0.019716
R46967 PAD.n7484 PAD.n7483 0.019716
R46968 PAD.n7483 PAD.n7194 0.019716
R46969 PAD.n7477 PAD.n7476 0.019716
R46970 PAD.n7477 PAD.n7193 0.019716
R46971 PAD.n7472 PAD.n7471 0.019716
R46972 PAD.n7471 PAD.n7192 0.019716
R46973 PAD.n7465 PAD.n7464 0.019716
R46974 PAD.n7465 PAD.n7191 0.019716
R46975 PAD.n7460 PAD.n7459 0.019716
R46976 PAD.n7459 PAD.n7190 0.019716
R46977 PAD.n7453 PAD.n7452 0.019716
R46978 PAD.n7453 PAD.n7189 0.019716
R46979 PAD.n7448 PAD.n7447 0.019716
R46980 PAD.n7447 PAD.n7188 0.019716
R46981 PAD.n7441 PAD.n7440 0.019716
R46982 PAD.n7441 PAD.n7187 0.019716
R46983 PAD.n7436 PAD.n7435 0.019716
R46984 PAD.n7435 PAD.n7186 0.019716
R46985 PAD.n7429 PAD.n7428 0.019716
R46986 PAD.n7429 PAD.n7185 0.019716
R46987 PAD.n7424 PAD.n7423 0.019716
R46988 PAD.n7423 PAD.n7184 0.019716
R46989 PAD.n7417 PAD.n7416 0.019716
R46990 PAD.n7417 PAD.n7183 0.019716
R46991 PAD.n7412 PAD.n7411 0.019716
R46992 PAD.n7411 PAD.n7182 0.019716
R46993 PAD.n7405 PAD.n7404 0.019716
R46994 PAD.n7405 PAD.n7181 0.019716
R46995 PAD.n7400 PAD.n7399 0.019716
R46996 PAD.n7399 PAD.n7180 0.019716
R46997 PAD.n7393 PAD.n7392 0.019716
R46998 PAD.n7393 PAD.n7179 0.019716
R46999 PAD.n7388 PAD.n7387 0.019716
R47000 PAD.n7387 PAD.n7178 0.019716
R47001 PAD.n7381 PAD.n7380 0.019716
R47002 PAD.n7381 PAD.n7177 0.019716
R47003 PAD.n7376 PAD.n7375 0.019716
R47004 PAD.n7375 PAD.n7176 0.019716
R47005 PAD.n7369 PAD.n7368 0.019716
R47006 PAD.n7369 PAD.n7175 0.019716
R47007 PAD.n7364 PAD.n7363 0.019716
R47008 PAD.n7363 PAD.n7174 0.019716
R47009 PAD.n7357 PAD.n7356 0.019716
R47010 PAD.n7357 PAD.n7173 0.019716
R47011 PAD.n7352 PAD.n7351 0.019716
R47012 PAD.n7351 PAD.n7172 0.019716
R47013 PAD.n7345 PAD.n7344 0.019716
R47014 PAD.n7345 PAD.n7171 0.019716
R47015 PAD.n7340 PAD.n7339 0.019716
R47016 PAD.n7339 PAD.n7170 0.019716
R47017 PAD.n7333 PAD.n7332 0.019716
R47018 PAD.n7333 PAD.n7169 0.019716
R47019 PAD.n7328 PAD.n7327 0.019716
R47020 PAD.n7327 PAD.n7168 0.019716
R47021 PAD.n7321 PAD.n7320 0.019716
R47022 PAD.n7321 PAD.n7167 0.019716
R47023 PAD.n7316 PAD.n7315 0.019716
R47024 PAD.n7315 PAD.n7166 0.019716
R47025 PAD.n7309 PAD.n7308 0.019716
R47026 PAD.n7309 PAD.n7165 0.019716
R47027 PAD.n7304 PAD.n7303 0.019716
R47028 PAD.n7303 PAD.n7164 0.019716
R47029 PAD.n7297 PAD.n7296 0.019716
R47030 PAD.n7297 PAD.n7163 0.019716
R47031 PAD.n7292 PAD.n7291 0.019716
R47032 PAD.n7291 PAD.n7162 0.019716
R47033 PAD.n7285 PAD.n7284 0.019716
R47034 PAD.n7285 PAD.n7161 0.019716
R47035 PAD.n7280 PAD.n7279 0.019716
R47036 PAD.n7279 PAD.n7160 0.019716
R47037 PAD.n7273 PAD.n7272 0.019716
R47038 PAD.n7273 PAD.n7159 0.019716
R47039 PAD.n10693 PAD.n10692 0.019716
R47040 PAD.n10417 PAD.n414 0.019716
R47041 PAD.n10417 PAD.n10416 0.019716
R47042 PAD.n10686 PAD.n413 0.019716
R47043 PAD.n10686 PAD.n10685 0.019716
R47044 PAD.n10422 PAD.n412 0.019716
R47045 PAD.n10422 PAD.n10421 0.019716
R47046 PAD.n10677 PAD.n411 0.019716
R47047 PAD.n10677 PAD.n10676 0.019716
R47048 PAD.n10427 PAD.n410 0.019716
R47049 PAD.n10427 PAD.n10426 0.019716
R47050 PAD.n10668 PAD.n409 0.019716
R47051 PAD.n10668 PAD.n10667 0.019716
R47052 PAD.n10432 PAD.n408 0.019716
R47053 PAD.n10432 PAD.n10431 0.019716
R47054 PAD.n10659 PAD.n407 0.019716
R47055 PAD.n10659 PAD.n10658 0.019716
R47056 PAD.n10437 PAD.n406 0.019716
R47057 PAD.n10437 PAD.n10436 0.019716
R47058 PAD.n10650 PAD.n405 0.019716
R47059 PAD.n10650 PAD.n10649 0.019716
R47060 PAD.n10442 PAD.n404 0.019716
R47061 PAD.n10442 PAD.n10441 0.019716
R47062 PAD.n10641 PAD.n403 0.019716
R47063 PAD.n10641 PAD.n10640 0.019716
R47064 PAD.n10447 PAD.n402 0.019716
R47065 PAD.n10447 PAD.n10446 0.019716
R47066 PAD.n10632 PAD.n401 0.019716
R47067 PAD.n10632 PAD.n10631 0.019716
R47068 PAD.n10452 PAD.n400 0.019716
R47069 PAD.n10452 PAD.n10451 0.019716
R47070 PAD.n10623 PAD.n399 0.019716
R47071 PAD.n10623 PAD.n10622 0.019716
R47072 PAD.n10457 PAD.n398 0.019716
R47073 PAD.n10457 PAD.n10456 0.019716
R47074 PAD.n10614 PAD.n397 0.019716
R47075 PAD.n10614 PAD.n10613 0.019716
R47076 PAD.n10462 PAD.n396 0.019716
R47077 PAD.n10462 PAD.n10461 0.019716
R47078 PAD.n10605 PAD.n395 0.019716
R47079 PAD.n10605 PAD.n10604 0.019716
R47080 PAD.n10467 PAD.n394 0.019716
R47081 PAD.n10467 PAD.n10466 0.019716
R47082 PAD.n10596 PAD.n393 0.019716
R47083 PAD.n10596 PAD.n10595 0.019716
R47084 PAD.n10472 PAD.n392 0.019716
R47085 PAD.n10472 PAD.n10471 0.019716
R47086 PAD.n10587 PAD.n391 0.019716
R47087 PAD.n10587 PAD.n10586 0.019716
R47088 PAD.n10477 PAD.n390 0.019716
R47089 PAD.n10477 PAD.n10476 0.019716
R47090 PAD.n10578 PAD.n389 0.019716
R47091 PAD.n10578 PAD.n10577 0.019716
R47092 PAD.n10482 PAD.n388 0.019716
R47093 PAD.n10482 PAD.n10481 0.019716
R47094 PAD.n10569 PAD.n387 0.019716
R47095 PAD.n10569 PAD.n10568 0.019716
R47096 PAD.n10487 PAD.n386 0.019716
R47097 PAD.n10487 PAD.n10486 0.019716
R47098 PAD.n10560 PAD.n385 0.019716
R47099 PAD.n10560 PAD.n10559 0.019716
R47100 PAD.n10492 PAD.n384 0.019716
R47101 PAD.n10492 PAD.n10491 0.019716
R47102 PAD.n10551 PAD.n383 0.019716
R47103 PAD.n10551 PAD.n10550 0.019716
R47104 PAD.n10497 PAD.n382 0.019716
R47105 PAD.n10497 PAD.n10496 0.019716
R47106 PAD.n10542 PAD.n381 0.019716
R47107 PAD.n10542 PAD.n10541 0.019716
R47108 PAD.n10502 PAD.n380 0.019716
R47109 PAD.n10502 PAD.n10501 0.019716
R47110 PAD.n10533 PAD.n379 0.019716
R47111 PAD.n10533 PAD.n10532 0.019716
R47112 PAD.n10507 PAD.n378 0.019716
R47113 PAD.n10507 PAD.n10506 0.019716
R47114 PAD.n10524 PAD.n377 0.019716
R47115 PAD.n10524 PAD.n10523 0.019716
R47116 PAD.n10512 PAD.n376 0.019716
R47117 PAD.n10512 PAD.n10511 0.019716
R47118 PAD.n10515 PAD.n375 0.019716
R47119 PAD.n10515 PAD.n10514 0.019716
R47120 PAD.n10713 PAD.n374 0.019716
R47121 PAD.n10714 PAD.n10713 0.019716
R47122 PAD.n525 PAD.n524 0.019716
R47123 PAD.n529 PAD.n526 0.019716
R47124 PAD.n529 PAD.n528 0.019716
R47125 PAD.n535 PAD.n517 0.019716
R47126 PAD.n536 PAD.n535 0.019716
R47127 PAD.n541 PAD.n538 0.019716
R47128 PAD.n541 PAD.n540 0.019716
R47129 PAD.n547 PAD.n513 0.019716
R47130 PAD.n548 PAD.n547 0.019716
R47131 PAD.n553 PAD.n550 0.019716
R47132 PAD.n553 PAD.n552 0.019716
R47133 PAD.n559 PAD.n509 0.019716
R47134 PAD.n560 PAD.n559 0.019716
R47135 PAD.n565 PAD.n562 0.019716
R47136 PAD.n565 PAD.n564 0.019716
R47137 PAD.n571 PAD.n505 0.019716
R47138 PAD.n572 PAD.n571 0.019716
R47139 PAD.n577 PAD.n574 0.019716
R47140 PAD.n577 PAD.n576 0.019716
R47141 PAD.n583 PAD.n501 0.019716
R47142 PAD.n584 PAD.n583 0.019716
R47143 PAD.n589 PAD.n586 0.019716
R47144 PAD.n589 PAD.n588 0.019716
R47145 PAD.n595 PAD.n497 0.019716
R47146 PAD.n596 PAD.n595 0.019716
R47147 PAD.n601 PAD.n598 0.019716
R47148 PAD.n601 PAD.n600 0.019716
R47149 PAD.n607 PAD.n493 0.019716
R47150 PAD.n608 PAD.n607 0.019716
R47151 PAD.n613 PAD.n610 0.019716
R47152 PAD.n613 PAD.n612 0.019716
R47153 PAD.n619 PAD.n489 0.019716
R47154 PAD.n620 PAD.n619 0.019716
R47155 PAD.n625 PAD.n622 0.019716
R47156 PAD.n625 PAD.n624 0.019716
R47157 PAD.n631 PAD.n485 0.019716
R47158 PAD.n632 PAD.n631 0.019716
R47159 PAD.n637 PAD.n634 0.019716
R47160 PAD.n637 PAD.n636 0.019716
R47161 PAD.n643 PAD.n481 0.019716
R47162 PAD.n644 PAD.n643 0.019716
R47163 PAD.n649 PAD.n646 0.019716
R47164 PAD.n649 PAD.n648 0.019716
R47165 PAD.n655 PAD.n477 0.019716
R47166 PAD.n656 PAD.n655 0.019716
R47167 PAD.n661 PAD.n658 0.019716
R47168 PAD.n661 PAD.n660 0.019716
R47169 PAD.n667 PAD.n473 0.019716
R47170 PAD.n668 PAD.n667 0.019716
R47171 PAD.n673 PAD.n670 0.019716
R47172 PAD.n673 PAD.n672 0.019716
R47173 PAD.n679 PAD.n469 0.019716
R47174 PAD.n680 PAD.n679 0.019716
R47175 PAD.n685 PAD.n682 0.019716
R47176 PAD.n685 PAD.n684 0.019716
R47177 PAD.n691 PAD.n465 0.019716
R47178 PAD.n692 PAD.n691 0.019716
R47179 PAD.n697 PAD.n694 0.019716
R47180 PAD.n697 PAD.n696 0.019716
R47181 PAD.n703 PAD.n461 0.019716
R47182 PAD.n704 PAD.n703 0.019716
R47183 PAD.n709 PAD.n706 0.019716
R47184 PAD.n709 PAD.n708 0.019716
R47185 PAD.n715 PAD.n457 0.019716
R47186 PAD.n716 PAD.n715 0.019716
R47187 PAD.n721 PAD.n718 0.019716
R47188 PAD.n721 PAD.n720 0.019716
R47189 PAD.n727 PAD.n453 0.019716
R47190 PAD.n728 PAD.n727 0.019716
R47191 PAD.n733 PAD.n730 0.019716
R47192 PAD.n733 PAD.n732 0.019716
R47193 PAD.n739 PAD.n449 0.019716
R47194 PAD.n740 PAD.n739 0.019716
R47195 PAD.n745 PAD.n742 0.019716
R47196 PAD.n745 PAD.n744 0.019716
R47197 PAD.n751 PAD.n445 0.019716
R47198 PAD.n752 PAD.n751 0.019716
R47199 PAD.n757 PAD.n754 0.019716
R47200 PAD.n757 PAD.n756 0.019716
R47201 PAD.n764 PAD.n441 0.019716
R47202 PAD.n765 PAD.n764 0.019716
R47203 PAD.n768 PAD.n767 0.019716
R47204 PAD.n769 PAD.n768 0.019716
R47205 PAD.n870 PAD.n869 0.019716
R47206 PAD.n877 PAD.n823 0.019716
R47207 PAD.n878 PAD.n877 0.019716
R47208 PAD.n883 PAD.n822 0.019716
R47209 PAD.n883 PAD.n882 0.019716
R47210 PAD.n889 PAD.n821 0.019716
R47211 PAD.n890 PAD.n889 0.019716
R47212 PAD.n895 PAD.n820 0.019716
R47213 PAD.n895 PAD.n894 0.019716
R47214 PAD.n901 PAD.n819 0.019716
R47215 PAD.n902 PAD.n901 0.019716
R47216 PAD.n907 PAD.n818 0.019716
R47217 PAD.n907 PAD.n906 0.019716
R47218 PAD.n913 PAD.n817 0.019716
R47219 PAD.n914 PAD.n913 0.019716
R47220 PAD.n919 PAD.n816 0.019716
R47221 PAD.n919 PAD.n918 0.019716
R47222 PAD.n925 PAD.n815 0.019716
R47223 PAD.n926 PAD.n925 0.019716
R47224 PAD.n931 PAD.n814 0.019716
R47225 PAD.n931 PAD.n930 0.019716
R47226 PAD.n937 PAD.n813 0.019716
R47227 PAD.n938 PAD.n937 0.019716
R47228 PAD.n943 PAD.n812 0.019716
R47229 PAD.n943 PAD.n942 0.019716
R47230 PAD.n949 PAD.n811 0.019716
R47231 PAD.n950 PAD.n949 0.019716
R47232 PAD.n955 PAD.n810 0.019716
R47233 PAD.n955 PAD.n954 0.019716
R47234 PAD.n961 PAD.n809 0.019716
R47235 PAD.n962 PAD.n961 0.019716
R47236 PAD.n967 PAD.n808 0.019716
R47237 PAD.n967 PAD.n966 0.019716
R47238 PAD.n973 PAD.n807 0.019716
R47239 PAD.n974 PAD.n973 0.019716
R47240 PAD.n979 PAD.n806 0.019716
R47241 PAD.n979 PAD.n978 0.019716
R47242 PAD.n985 PAD.n805 0.019716
R47243 PAD.n986 PAD.n985 0.019716
R47244 PAD.n991 PAD.n804 0.019716
R47245 PAD.n991 PAD.n990 0.019716
R47246 PAD.n997 PAD.n803 0.019716
R47247 PAD.n998 PAD.n997 0.019716
R47248 PAD.n1003 PAD.n802 0.019716
R47249 PAD.n1003 PAD.n1002 0.019716
R47250 PAD.n1009 PAD.n801 0.019716
R47251 PAD.n1010 PAD.n1009 0.019716
R47252 PAD.n1015 PAD.n800 0.019716
R47253 PAD.n1015 PAD.n1014 0.019716
R47254 PAD.n1021 PAD.n799 0.019716
R47255 PAD.n1022 PAD.n1021 0.019716
R47256 PAD.n1027 PAD.n798 0.019716
R47257 PAD.n1027 PAD.n1026 0.019716
R47258 PAD.n1033 PAD.n797 0.019716
R47259 PAD.n1034 PAD.n1033 0.019716
R47260 PAD.n1039 PAD.n796 0.019716
R47261 PAD.n1039 PAD.n1038 0.019716
R47262 PAD.n1045 PAD.n795 0.019716
R47263 PAD.n1046 PAD.n1045 0.019716
R47264 PAD.n1051 PAD.n794 0.019716
R47265 PAD.n1051 PAD.n1050 0.019716
R47266 PAD.n1057 PAD.n793 0.019716
R47267 PAD.n1058 PAD.n1057 0.019716
R47268 PAD.n1063 PAD.n792 0.019716
R47269 PAD.n1063 PAD.n1062 0.019716
R47270 PAD.n1069 PAD.n791 0.019716
R47271 PAD.n1070 PAD.n1069 0.019716
R47272 PAD.n1075 PAD.n790 0.019716
R47273 PAD.n1075 PAD.n1074 0.019716
R47274 PAD.n1081 PAD.n789 0.019716
R47275 PAD.n1082 PAD.n1081 0.019716
R47276 PAD.n1087 PAD.n788 0.019716
R47277 PAD.n1087 PAD.n1086 0.019716
R47278 PAD.n1093 PAD.n787 0.019716
R47279 PAD.n1094 PAD.n1093 0.019716
R47280 PAD.n1099 PAD.n786 0.019716
R47281 PAD.n1099 PAD.n1098 0.019716
R47282 PAD.n1105 PAD.n785 0.019716
R47283 PAD.n1106 PAD.n1105 0.019716
R47284 PAD.n1111 PAD.n784 0.019716
R47285 PAD.n1111 PAD.n1110 0.019716
R47286 PAD.n10385 PAD.n783 0.019716
R47287 PAD.n10386 PAD.n10385 0.019716
R47288 PAD.n10108 PAD.n10107 0.019716
R47289 PAD.n10112 PAD.n10109 0.019716
R47290 PAD.n10112 PAD.n10111 0.019716
R47291 PAD.n10118 PAD.n10101 0.019716
R47292 PAD.n10119 PAD.n10118 0.019716
R47293 PAD.n10124 PAD.n10121 0.019716
R47294 PAD.n10124 PAD.n10123 0.019716
R47295 PAD.n10130 PAD.n10097 0.019716
R47296 PAD.n10131 PAD.n10130 0.019716
R47297 PAD.n10136 PAD.n10133 0.019716
R47298 PAD.n10136 PAD.n10135 0.019716
R47299 PAD.n10142 PAD.n10093 0.019716
R47300 PAD.n10143 PAD.n10142 0.019716
R47301 PAD.n10148 PAD.n10145 0.019716
R47302 PAD.n10148 PAD.n10147 0.019716
R47303 PAD.n10154 PAD.n10089 0.019716
R47304 PAD.n10155 PAD.n10154 0.019716
R47305 PAD.n10160 PAD.n10157 0.019716
R47306 PAD.n10160 PAD.n10159 0.019716
R47307 PAD.n10166 PAD.n10085 0.019716
R47308 PAD.n10167 PAD.n10166 0.019716
R47309 PAD.n10172 PAD.n10169 0.019716
R47310 PAD.n10172 PAD.n10171 0.019716
R47311 PAD.n10178 PAD.n10081 0.019716
R47312 PAD.n10179 PAD.n10178 0.019716
R47313 PAD.n10184 PAD.n10181 0.019716
R47314 PAD.n10184 PAD.n10183 0.019716
R47315 PAD.n10190 PAD.n10077 0.019716
R47316 PAD.n10191 PAD.n10190 0.019716
R47317 PAD.n10196 PAD.n10193 0.019716
R47318 PAD.n10196 PAD.n10195 0.019716
R47319 PAD.n10202 PAD.n10073 0.019716
R47320 PAD.n10203 PAD.n10202 0.019716
R47321 PAD.n10208 PAD.n10205 0.019716
R47322 PAD.n10208 PAD.n10207 0.019716
R47323 PAD.n10214 PAD.n10069 0.019716
R47324 PAD.n10215 PAD.n10214 0.019716
R47325 PAD.n10220 PAD.n10217 0.019716
R47326 PAD.n10220 PAD.n10219 0.019716
R47327 PAD.n10226 PAD.n10065 0.019716
R47328 PAD.n10227 PAD.n10226 0.019716
R47329 PAD.n10232 PAD.n10229 0.019716
R47330 PAD.n10232 PAD.n10231 0.019716
R47331 PAD.n10238 PAD.n10061 0.019716
R47332 PAD.n10239 PAD.n10238 0.019716
R47333 PAD.n10244 PAD.n10241 0.019716
R47334 PAD.n10244 PAD.n10243 0.019716
R47335 PAD.n10250 PAD.n10057 0.019716
R47336 PAD.n10251 PAD.n10250 0.019716
R47337 PAD.n10256 PAD.n10253 0.019716
R47338 PAD.n10256 PAD.n10255 0.019716
R47339 PAD.n10262 PAD.n10053 0.019716
R47340 PAD.n10263 PAD.n10262 0.019716
R47341 PAD.n10268 PAD.n10265 0.019716
R47342 PAD.n10268 PAD.n10267 0.019716
R47343 PAD.n10274 PAD.n10049 0.019716
R47344 PAD.n10275 PAD.n10274 0.019716
R47345 PAD.n10280 PAD.n10277 0.019716
R47346 PAD.n10280 PAD.n10279 0.019716
R47347 PAD.n10286 PAD.n10045 0.019716
R47348 PAD.n10287 PAD.n10286 0.019716
R47349 PAD.n10292 PAD.n10289 0.019716
R47350 PAD.n10292 PAD.n10291 0.019716
R47351 PAD.n10298 PAD.n10041 0.019716
R47352 PAD.n10299 PAD.n10298 0.019716
R47353 PAD.n10304 PAD.n10301 0.019716
R47354 PAD.n10304 PAD.n10303 0.019716
R47355 PAD.n10310 PAD.n10037 0.019716
R47356 PAD.n10311 PAD.n10310 0.019716
R47357 PAD.n10316 PAD.n10313 0.019716
R47358 PAD.n10316 PAD.n10315 0.019716
R47359 PAD.n10322 PAD.n10033 0.019716
R47360 PAD.n10323 PAD.n10322 0.019716
R47361 PAD.n10328 PAD.n10325 0.019716
R47362 PAD.n10328 PAD.n10327 0.019716
R47363 PAD.n10334 PAD.n10029 0.019716
R47364 PAD.n10335 PAD.n10334 0.019716
R47365 PAD.n10340 PAD.n10337 0.019716
R47366 PAD.n10340 PAD.n10339 0.019716
R47367 PAD.n10347 PAD.n10025 0.019716
R47368 PAD.n10348 PAD.n10347 0.019716
R47369 PAD.n10351 PAD.n10350 0.019716
R47370 PAD.n10352 PAD.n10351 0.019716
R47371 PAD.n1482 PAD.n1190 0.019716
R47372 PAD.n1192 PAD.n1191 0.019716
R47373 PAD.n1192 PAD.n1189 0.019716
R47374 PAD.n1473 PAD.n1472 0.019716
R47375 PAD.n1472 PAD.n1188 0.019716
R47376 PAD.n1197 PAD.n1196 0.019716
R47377 PAD.n1196 PAD.n1187 0.019716
R47378 PAD.n1464 PAD.n1463 0.019716
R47379 PAD.n1463 PAD.n1186 0.019716
R47380 PAD.n1202 PAD.n1201 0.019716
R47381 PAD.n1201 PAD.n1185 0.019716
R47382 PAD.n1455 PAD.n1454 0.019716
R47383 PAD.n1454 PAD.n1184 0.019716
R47384 PAD.n1207 PAD.n1206 0.019716
R47385 PAD.n1206 PAD.n1183 0.019716
R47386 PAD.n1446 PAD.n1445 0.019716
R47387 PAD.n1445 PAD.n1182 0.019716
R47388 PAD.n1212 PAD.n1211 0.019716
R47389 PAD.n1211 PAD.n1181 0.019716
R47390 PAD.n1437 PAD.n1436 0.019716
R47391 PAD.n1436 PAD.n1180 0.019716
R47392 PAD.n1217 PAD.n1216 0.019716
R47393 PAD.n1216 PAD.n1179 0.019716
R47394 PAD.n1428 PAD.n1427 0.019716
R47395 PAD.n1427 PAD.n1178 0.019716
R47396 PAD.n1222 PAD.n1221 0.019716
R47397 PAD.n1221 PAD.n1177 0.019716
R47398 PAD.n1419 PAD.n1418 0.019716
R47399 PAD.n1418 PAD.n1176 0.019716
R47400 PAD.n1227 PAD.n1226 0.019716
R47401 PAD.n1226 PAD.n1175 0.019716
R47402 PAD.n1410 PAD.n1409 0.019716
R47403 PAD.n1409 PAD.n1174 0.019716
R47404 PAD.n1232 PAD.n1231 0.019716
R47405 PAD.n1231 PAD.n1173 0.019716
R47406 PAD.n1401 PAD.n1400 0.019716
R47407 PAD.n1400 PAD.n1172 0.019716
R47408 PAD.n1237 PAD.n1236 0.019716
R47409 PAD.n1236 PAD.n1171 0.019716
R47410 PAD.n1392 PAD.n1391 0.019716
R47411 PAD.n1391 PAD.n1170 0.019716
R47412 PAD.n1242 PAD.n1241 0.019716
R47413 PAD.n1241 PAD.n1169 0.019716
R47414 PAD.n1383 PAD.n1382 0.019716
R47415 PAD.n1382 PAD.n1168 0.019716
R47416 PAD.n1247 PAD.n1246 0.019716
R47417 PAD.n1246 PAD.n1167 0.019716
R47418 PAD.n1374 PAD.n1373 0.019716
R47419 PAD.n1373 PAD.n1166 0.019716
R47420 PAD.n1252 PAD.n1251 0.019716
R47421 PAD.n1251 PAD.n1165 0.019716
R47422 PAD.n1365 PAD.n1364 0.019716
R47423 PAD.n1364 PAD.n1164 0.019716
R47424 PAD.n1257 PAD.n1256 0.019716
R47425 PAD.n1256 PAD.n1163 0.019716
R47426 PAD.n1356 PAD.n1355 0.019716
R47427 PAD.n1355 PAD.n1162 0.019716
R47428 PAD.n1262 PAD.n1261 0.019716
R47429 PAD.n1261 PAD.n1161 0.019716
R47430 PAD.n1347 PAD.n1346 0.019716
R47431 PAD.n1346 PAD.n1160 0.019716
R47432 PAD.n1267 PAD.n1266 0.019716
R47433 PAD.n1266 PAD.n1159 0.019716
R47434 PAD.n1338 PAD.n1337 0.019716
R47435 PAD.n1337 PAD.n1158 0.019716
R47436 PAD.n1272 PAD.n1271 0.019716
R47437 PAD.n1271 PAD.n1157 0.019716
R47438 PAD.n1329 PAD.n1328 0.019716
R47439 PAD.n1328 PAD.n1156 0.019716
R47440 PAD.n1277 PAD.n1276 0.019716
R47441 PAD.n1276 PAD.n1155 0.019716
R47442 PAD.n1320 PAD.n1319 0.019716
R47443 PAD.n1319 PAD.n1154 0.019716
R47444 PAD.n1282 PAD.n1281 0.019716
R47445 PAD.n1281 PAD.n1153 0.019716
R47446 PAD.n1311 PAD.n1310 0.019716
R47447 PAD.n1310 PAD.n1152 0.019716
R47448 PAD.n1287 PAD.n1286 0.019716
R47449 PAD.n1286 PAD.n1151 0.019716
R47450 PAD.n1302 PAD.n1301 0.019716
R47451 PAD.n1301 PAD.n1150 0.019716
R47452 PAD.n1292 PAD.n1291 0.019716
R47453 PAD.n1291 PAD.n1149 0.019716
R47454 PAD.n1578 PAD.n1577 0.019716
R47455 PAD.n9754 PAD.n1530 0.019716
R47456 PAD.n9755 PAD.n9754 0.019716
R47457 PAD.n9760 PAD.n1529 0.019716
R47458 PAD.n9760 PAD.n9759 0.019716
R47459 PAD.n9766 PAD.n1528 0.019716
R47460 PAD.n9767 PAD.n9766 0.019716
R47461 PAD.n9772 PAD.n1527 0.019716
R47462 PAD.n9772 PAD.n9771 0.019716
R47463 PAD.n9778 PAD.n1526 0.019716
R47464 PAD.n9779 PAD.n9778 0.019716
R47465 PAD.n9784 PAD.n1525 0.019716
R47466 PAD.n9784 PAD.n9783 0.019716
R47467 PAD.n9790 PAD.n1524 0.019716
R47468 PAD.n9791 PAD.n9790 0.019716
R47469 PAD.n9796 PAD.n1523 0.019716
R47470 PAD.n9796 PAD.n9795 0.019716
R47471 PAD.n9802 PAD.n1522 0.019716
R47472 PAD.n9803 PAD.n9802 0.019716
R47473 PAD.n9808 PAD.n1521 0.019716
R47474 PAD.n9808 PAD.n9807 0.019716
R47475 PAD.n9814 PAD.n1520 0.019716
R47476 PAD.n9815 PAD.n9814 0.019716
R47477 PAD.n9820 PAD.n1519 0.019716
R47478 PAD.n9820 PAD.n9819 0.019716
R47479 PAD.n9826 PAD.n1518 0.019716
R47480 PAD.n9827 PAD.n9826 0.019716
R47481 PAD.n9832 PAD.n1517 0.019716
R47482 PAD.n9832 PAD.n9831 0.019716
R47483 PAD.n9838 PAD.n1516 0.019716
R47484 PAD.n9839 PAD.n9838 0.019716
R47485 PAD.n9844 PAD.n1515 0.019716
R47486 PAD.n9844 PAD.n9843 0.019716
R47487 PAD.n9850 PAD.n1514 0.019716
R47488 PAD.n9851 PAD.n9850 0.019716
R47489 PAD.n9856 PAD.n1513 0.019716
R47490 PAD.n9856 PAD.n9855 0.019716
R47491 PAD.n9862 PAD.n1512 0.019716
R47492 PAD.n9863 PAD.n9862 0.019716
R47493 PAD.n9868 PAD.n1511 0.019716
R47494 PAD.n9868 PAD.n9867 0.019716
R47495 PAD.n9874 PAD.n1510 0.019716
R47496 PAD.n9875 PAD.n9874 0.019716
R47497 PAD.n9880 PAD.n1509 0.019716
R47498 PAD.n9880 PAD.n9879 0.019716
R47499 PAD.n9886 PAD.n1508 0.019716
R47500 PAD.n9887 PAD.n9886 0.019716
R47501 PAD.n9892 PAD.n1507 0.019716
R47502 PAD.n9892 PAD.n9891 0.019716
R47503 PAD.n9898 PAD.n1506 0.019716
R47504 PAD.n9899 PAD.n9898 0.019716
R47505 PAD.n9904 PAD.n1505 0.019716
R47506 PAD.n9904 PAD.n9903 0.019716
R47507 PAD.n9910 PAD.n1504 0.019716
R47508 PAD.n9911 PAD.n9910 0.019716
R47509 PAD.n9916 PAD.n1503 0.019716
R47510 PAD.n9916 PAD.n9915 0.019716
R47511 PAD.n9922 PAD.n1502 0.019716
R47512 PAD.n9923 PAD.n9922 0.019716
R47513 PAD.n9928 PAD.n1501 0.019716
R47514 PAD.n9928 PAD.n9927 0.019716
R47515 PAD.n9934 PAD.n1500 0.019716
R47516 PAD.n9935 PAD.n9934 0.019716
R47517 PAD.n9940 PAD.n1499 0.019716
R47518 PAD.n9940 PAD.n9939 0.019716
R47519 PAD.n9946 PAD.n1498 0.019716
R47520 PAD.n9947 PAD.n9946 0.019716
R47521 PAD.n9952 PAD.n1497 0.019716
R47522 PAD.n9952 PAD.n9951 0.019716
R47523 PAD.n9958 PAD.n1496 0.019716
R47524 PAD.n9959 PAD.n9958 0.019716
R47525 PAD.n9964 PAD.n1495 0.019716
R47526 PAD.n9964 PAD.n9963 0.019716
R47527 PAD.n9970 PAD.n1494 0.019716
R47528 PAD.n9971 PAD.n9970 0.019716
R47529 PAD.n9976 PAD.n1493 0.019716
R47530 PAD.n9976 PAD.n9975 0.019716
R47531 PAD.n9982 PAD.n1492 0.019716
R47532 PAD.n9983 PAD.n9982 0.019716
R47533 PAD.n9988 PAD.n1491 0.019716
R47534 PAD.n9988 PAD.n9987 0.019716
R47535 PAD.n9995 PAD.n1490 0.019716
R47536 PAD.n9996 PAD.n9995 0.019716
R47537 PAD.n1929 PAD.n1601 0.019716
R47538 PAD.n1928 PAD.n1927 0.019716
R47539 PAD.n1927 PAD.n1926 0.019716
R47540 PAD.n1917 PAD.n1602 0.019716
R47541 PAD.n1918 PAD.n1917 0.019716
R47542 PAD.n1916 PAD.n1915 0.019716
R47543 PAD.n1915 PAD.n1914 0.019716
R47544 PAD.n1905 PAD.n1607 0.019716
R47545 PAD.n1906 PAD.n1905 0.019716
R47546 PAD.n1904 PAD.n1903 0.019716
R47547 PAD.n1903 PAD.n1902 0.019716
R47548 PAD.n1893 PAD.n1611 0.019716
R47549 PAD.n1894 PAD.n1893 0.019716
R47550 PAD.n1892 PAD.n1891 0.019716
R47551 PAD.n1891 PAD.n1890 0.019716
R47552 PAD.n1881 PAD.n1615 0.019716
R47553 PAD.n1882 PAD.n1881 0.019716
R47554 PAD.n1880 PAD.n1879 0.019716
R47555 PAD.n1879 PAD.n1878 0.019716
R47556 PAD.n1869 PAD.n1619 0.019716
R47557 PAD.n1870 PAD.n1869 0.019716
R47558 PAD.n1868 PAD.n1867 0.019716
R47559 PAD.n1867 PAD.n1866 0.019716
R47560 PAD.n1857 PAD.n1623 0.019716
R47561 PAD.n1858 PAD.n1857 0.019716
R47562 PAD.n1856 PAD.n1855 0.019716
R47563 PAD.n1855 PAD.n1854 0.019716
R47564 PAD.n1845 PAD.n1627 0.019716
R47565 PAD.n1846 PAD.n1845 0.019716
R47566 PAD.n1844 PAD.n1843 0.019716
R47567 PAD.n1843 PAD.n1842 0.019716
R47568 PAD.n1833 PAD.n1631 0.019716
R47569 PAD.n1834 PAD.n1833 0.019716
R47570 PAD.n1832 PAD.n1831 0.019716
R47571 PAD.n1831 PAD.n1830 0.019716
R47572 PAD.n1821 PAD.n1635 0.019716
R47573 PAD.n1822 PAD.n1821 0.019716
R47574 PAD.n1820 PAD.n1819 0.019716
R47575 PAD.n1819 PAD.n1818 0.019716
R47576 PAD.n1809 PAD.n1639 0.019716
R47577 PAD.n1810 PAD.n1809 0.019716
R47578 PAD.n1808 PAD.n1807 0.019716
R47579 PAD.n1807 PAD.n1806 0.019716
R47580 PAD.n1797 PAD.n1643 0.019716
R47581 PAD.n1798 PAD.n1797 0.019716
R47582 PAD.n1796 PAD.n1795 0.019716
R47583 PAD.n1795 PAD.n1794 0.019716
R47584 PAD.n1785 PAD.n1647 0.019716
R47585 PAD.n1786 PAD.n1785 0.019716
R47586 PAD.n1784 PAD.n1783 0.019716
R47587 PAD.n1783 PAD.n1782 0.019716
R47588 PAD.n1773 PAD.n1651 0.019716
R47589 PAD.n1774 PAD.n1773 0.019716
R47590 PAD.n1772 PAD.n1771 0.019716
R47591 PAD.n1771 PAD.n1770 0.019716
R47592 PAD.n1761 PAD.n1655 0.019716
R47593 PAD.n1762 PAD.n1761 0.019716
R47594 PAD.n1760 PAD.n1759 0.019716
R47595 PAD.n1759 PAD.n1758 0.019716
R47596 PAD.n1749 PAD.n1659 0.019716
R47597 PAD.n1750 PAD.n1749 0.019716
R47598 PAD.n1748 PAD.n1747 0.019716
R47599 PAD.n1747 PAD.n1746 0.019716
R47600 PAD.n1737 PAD.n1663 0.019716
R47601 PAD.n1738 PAD.n1737 0.019716
R47602 PAD.n1736 PAD.n1735 0.019716
R47603 PAD.n1735 PAD.n1734 0.019716
R47604 PAD.n1725 PAD.n1667 0.019716
R47605 PAD.n1726 PAD.n1725 0.019716
R47606 PAD.n1724 PAD.n1723 0.019716
R47607 PAD.n1723 PAD.n1722 0.019716
R47608 PAD.n1713 PAD.n1671 0.019716
R47609 PAD.n1714 PAD.n1713 0.019716
R47610 PAD.n1712 PAD.n1711 0.019716
R47611 PAD.n1711 PAD.n1710 0.019716
R47612 PAD.n1701 PAD.n1675 0.019716
R47613 PAD.n1702 PAD.n1701 0.019716
R47614 PAD.n1700 PAD.n1699 0.019716
R47615 PAD.n1699 PAD.n1698 0.019716
R47616 PAD.n1689 PAD.n1679 0.019716
R47617 PAD.n1690 PAD.n1689 0.019716
R47618 PAD.n1688 PAD.n1687 0.019716
R47619 PAD.n1687 PAD.n1686 0.019716
R47620 PAD.n2030 PAD.n2029 0.019716
R47621 PAD.n9468 PAD.n1983 0.019716
R47622 PAD.n9469 PAD.n9468 0.019716
R47623 PAD.n9474 PAD.n1982 0.019716
R47624 PAD.n9474 PAD.n9473 0.019716
R47625 PAD.n9480 PAD.n1981 0.019716
R47626 PAD.n9481 PAD.n9480 0.019716
R47627 PAD.n9486 PAD.n1980 0.019716
R47628 PAD.n9486 PAD.n9485 0.019716
R47629 PAD.n9492 PAD.n1979 0.019716
R47630 PAD.n9493 PAD.n9492 0.019716
R47631 PAD.n9498 PAD.n1978 0.019716
R47632 PAD.n9498 PAD.n9497 0.019716
R47633 PAD.n9504 PAD.n1977 0.019716
R47634 PAD.n9505 PAD.n9504 0.019716
R47635 PAD.n9510 PAD.n1976 0.019716
R47636 PAD.n9510 PAD.n9509 0.019716
R47637 PAD.n9516 PAD.n1975 0.019716
R47638 PAD.n9517 PAD.n9516 0.019716
R47639 PAD.n9522 PAD.n1974 0.019716
R47640 PAD.n9522 PAD.n9521 0.019716
R47641 PAD.n9528 PAD.n1973 0.019716
R47642 PAD.n9529 PAD.n9528 0.019716
R47643 PAD.n9534 PAD.n1972 0.019716
R47644 PAD.n9534 PAD.n9533 0.019716
R47645 PAD.n9540 PAD.n1971 0.019716
R47646 PAD.n9541 PAD.n9540 0.019716
R47647 PAD.n9546 PAD.n1970 0.019716
R47648 PAD.n9546 PAD.n9545 0.019716
R47649 PAD.n9552 PAD.n1969 0.019716
R47650 PAD.n9553 PAD.n9552 0.019716
R47651 PAD.n9558 PAD.n1968 0.019716
R47652 PAD.n9558 PAD.n9557 0.019716
R47653 PAD.n9564 PAD.n1967 0.019716
R47654 PAD.n9565 PAD.n9564 0.019716
R47655 PAD.n9570 PAD.n1966 0.019716
R47656 PAD.n9570 PAD.n9569 0.019716
R47657 PAD.n9576 PAD.n1965 0.019716
R47658 PAD.n9577 PAD.n9576 0.019716
R47659 PAD.n9582 PAD.n1964 0.019716
R47660 PAD.n9582 PAD.n9581 0.019716
R47661 PAD.n9588 PAD.n1963 0.019716
R47662 PAD.n9589 PAD.n9588 0.019716
R47663 PAD.n9594 PAD.n1962 0.019716
R47664 PAD.n9594 PAD.n9593 0.019716
R47665 PAD.n9600 PAD.n1961 0.019716
R47666 PAD.n9601 PAD.n9600 0.019716
R47667 PAD.n9606 PAD.n1960 0.019716
R47668 PAD.n9606 PAD.n9605 0.019716
R47669 PAD.n9612 PAD.n1959 0.019716
R47670 PAD.n9613 PAD.n9612 0.019716
R47671 PAD.n9618 PAD.n1958 0.019716
R47672 PAD.n9618 PAD.n9617 0.019716
R47673 PAD.n9624 PAD.n1957 0.019716
R47674 PAD.n9625 PAD.n9624 0.019716
R47675 PAD.n9630 PAD.n1956 0.019716
R47676 PAD.n9630 PAD.n9629 0.019716
R47677 PAD.n9636 PAD.n1955 0.019716
R47678 PAD.n9637 PAD.n9636 0.019716
R47679 PAD.n9642 PAD.n1954 0.019716
R47680 PAD.n9642 PAD.n9641 0.019716
R47681 PAD.n9648 PAD.n1953 0.019716
R47682 PAD.n9649 PAD.n9648 0.019716
R47683 PAD.n9654 PAD.n1952 0.019716
R47684 PAD.n9654 PAD.n9653 0.019716
R47685 PAD.n9660 PAD.n1951 0.019716
R47686 PAD.n9661 PAD.n9660 0.019716
R47687 PAD.n9666 PAD.n1950 0.019716
R47688 PAD.n9666 PAD.n9665 0.019716
R47689 PAD.n9672 PAD.n1949 0.019716
R47690 PAD.n9673 PAD.n9672 0.019716
R47691 PAD.n9678 PAD.n1948 0.019716
R47692 PAD.n9678 PAD.n9677 0.019716
R47693 PAD.n9684 PAD.n1947 0.019716
R47694 PAD.n9685 PAD.n9684 0.019716
R47695 PAD.n9690 PAD.n1946 0.019716
R47696 PAD.n9690 PAD.n9689 0.019716
R47697 PAD.n9696 PAD.n1945 0.019716
R47698 PAD.n9697 PAD.n9696 0.019716
R47699 PAD.n9702 PAD.n1944 0.019716
R47700 PAD.n9702 PAD.n9701 0.019716
R47701 PAD.n9709 PAD.n1943 0.019716
R47702 PAD.n9710 PAD.n9709 0.019716
R47703 PAD.n2133 PAD.n2132 0.019716
R47704 PAD.n9202 PAD.n2087 0.019716
R47705 PAD.n9203 PAD.n9202 0.019716
R47706 PAD.n9208 PAD.n2086 0.019716
R47707 PAD.n9208 PAD.n9207 0.019716
R47708 PAD.n9214 PAD.n2085 0.019716
R47709 PAD.n9215 PAD.n9214 0.019716
R47710 PAD.n9220 PAD.n2084 0.019716
R47711 PAD.n9220 PAD.n9219 0.019716
R47712 PAD.n9226 PAD.n2083 0.019716
R47713 PAD.n9227 PAD.n9226 0.019716
R47714 PAD.n9232 PAD.n2082 0.019716
R47715 PAD.n9232 PAD.n9231 0.019716
R47716 PAD.n9238 PAD.n2081 0.019716
R47717 PAD.n9239 PAD.n9238 0.019716
R47718 PAD.n9244 PAD.n2080 0.019716
R47719 PAD.n9244 PAD.n9243 0.019716
R47720 PAD.n9250 PAD.n2079 0.019716
R47721 PAD.n9251 PAD.n9250 0.019716
R47722 PAD.n9256 PAD.n2078 0.019716
R47723 PAD.n9256 PAD.n9255 0.019716
R47724 PAD.n9262 PAD.n2077 0.019716
R47725 PAD.n9263 PAD.n9262 0.019716
R47726 PAD.n9268 PAD.n2076 0.019716
R47727 PAD.n9268 PAD.n9267 0.019716
R47728 PAD.n9274 PAD.n2075 0.019716
R47729 PAD.n9275 PAD.n9274 0.019716
R47730 PAD.n9280 PAD.n2074 0.019716
R47731 PAD.n9280 PAD.n9279 0.019716
R47732 PAD.n9286 PAD.n2073 0.019716
R47733 PAD.n9287 PAD.n9286 0.019716
R47734 PAD.n9292 PAD.n2072 0.019716
R47735 PAD.n9292 PAD.n9291 0.019716
R47736 PAD.n9298 PAD.n2071 0.019716
R47737 PAD.n9299 PAD.n9298 0.019716
R47738 PAD.n9304 PAD.n2070 0.019716
R47739 PAD.n9304 PAD.n9303 0.019716
R47740 PAD.n9310 PAD.n2069 0.019716
R47741 PAD.n9311 PAD.n9310 0.019716
R47742 PAD.n9316 PAD.n2068 0.019716
R47743 PAD.n9316 PAD.n9315 0.019716
R47744 PAD.n9322 PAD.n2067 0.019716
R47745 PAD.n9323 PAD.n9322 0.019716
R47746 PAD.n9328 PAD.n2066 0.019716
R47747 PAD.n9328 PAD.n9327 0.019716
R47748 PAD.n9334 PAD.n2065 0.019716
R47749 PAD.n9335 PAD.n9334 0.019716
R47750 PAD.n9340 PAD.n2064 0.019716
R47751 PAD.n9340 PAD.n9339 0.019716
R47752 PAD.n9346 PAD.n2063 0.019716
R47753 PAD.n9347 PAD.n9346 0.019716
R47754 PAD.n9352 PAD.n2062 0.019716
R47755 PAD.n9352 PAD.n9351 0.019716
R47756 PAD.n9358 PAD.n2061 0.019716
R47757 PAD.n9359 PAD.n9358 0.019716
R47758 PAD.n9364 PAD.n2060 0.019716
R47759 PAD.n9364 PAD.n9363 0.019716
R47760 PAD.n9370 PAD.n2059 0.019716
R47761 PAD.n9371 PAD.n9370 0.019716
R47762 PAD.n9376 PAD.n2058 0.019716
R47763 PAD.n9376 PAD.n9375 0.019716
R47764 PAD.n9382 PAD.n2057 0.019716
R47765 PAD.n9383 PAD.n9382 0.019716
R47766 PAD.n9388 PAD.n2056 0.019716
R47767 PAD.n9388 PAD.n9387 0.019716
R47768 PAD.n9394 PAD.n2055 0.019716
R47769 PAD.n9395 PAD.n9394 0.019716
R47770 PAD.n9400 PAD.n2054 0.019716
R47771 PAD.n9400 PAD.n9399 0.019716
R47772 PAD.n9406 PAD.n2053 0.019716
R47773 PAD.n9407 PAD.n9406 0.019716
R47774 PAD.n9412 PAD.n2052 0.019716
R47775 PAD.n9412 PAD.n9411 0.019716
R47776 PAD.n9418 PAD.n2051 0.019716
R47777 PAD.n9419 PAD.n9418 0.019716
R47778 PAD.n9424 PAD.n2050 0.019716
R47779 PAD.n9424 PAD.n9423 0.019716
R47780 PAD.n9430 PAD.n2049 0.019716
R47781 PAD.n9431 PAD.n9430 0.019716
R47782 PAD.n9436 PAD.n2048 0.019716
R47783 PAD.n9436 PAD.n9435 0.019716
R47784 PAD.n9442 PAD.n2047 0.019716
R47785 PAD.n9443 PAD.n9442 0.019716
R47786 PAD.n2480 PAD.n2153 0.019716
R47787 PAD.n2479 PAD.n2478 0.019716
R47788 PAD.n2478 PAD.n2477 0.019716
R47789 PAD.n2468 PAD.n2154 0.019716
R47790 PAD.n2469 PAD.n2468 0.019716
R47791 PAD.n2467 PAD.n2466 0.019716
R47792 PAD.n2466 PAD.n2465 0.019716
R47793 PAD.n2456 PAD.n2159 0.019716
R47794 PAD.n2457 PAD.n2456 0.019716
R47795 PAD.n2455 PAD.n2454 0.019716
R47796 PAD.n2454 PAD.n2453 0.019716
R47797 PAD.n2444 PAD.n2163 0.019716
R47798 PAD.n2445 PAD.n2444 0.019716
R47799 PAD.n2443 PAD.n2442 0.019716
R47800 PAD.n2442 PAD.n2441 0.019716
R47801 PAD.n2432 PAD.n2167 0.019716
R47802 PAD.n2433 PAD.n2432 0.019716
R47803 PAD.n2431 PAD.n2430 0.019716
R47804 PAD.n2430 PAD.n2429 0.019716
R47805 PAD.n2420 PAD.n2171 0.019716
R47806 PAD.n2421 PAD.n2420 0.019716
R47807 PAD.n2419 PAD.n2418 0.019716
R47808 PAD.n2418 PAD.n2417 0.019716
R47809 PAD.n2408 PAD.n2175 0.019716
R47810 PAD.n2409 PAD.n2408 0.019716
R47811 PAD.n2407 PAD.n2406 0.019716
R47812 PAD.n2406 PAD.n2405 0.019716
R47813 PAD.n2396 PAD.n2179 0.019716
R47814 PAD.n2397 PAD.n2396 0.019716
R47815 PAD.n2395 PAD.n2394 0.019716
R47816 PAD.n2394 PAD.n2393 0.019716
R47817 PAD.n2384 PAD.n2183 0.019716
R47818 PAD.n2385 PAD.n2384 0.019716
R47819 PAD.n2383 PAD.n2382 0.019716
R47820 PAD.n2382 PAD.n2381 0.019716
R47821 PAD.n2372 PAD.n2187 0.019716
R47822 PAD.n2373 PAD.n2372 0.019716
R47823 PAD.n2371 PAD.n2370 0.019716
R47824 PAD.n2370 PAD.n2369 0.019716
R47825 PAD.n2360 PAD.n2191 0.019716
R47826 PAD.n2361 PAD.n2360 0.019716
R47827 PAD.n2359 PAD.n2358 0.019716
R47828 PAD.n2358 PAD.n2357 0.019716
R47829 PAD.n2348 PAD.n2195 0.019716
R47830 PAD.n2349 PAD.n2348 0.019716
R47831 PAD.n2347 PAD.n2346 0.019716
R47832 PAD.n2346 PAD.n2345 0.019716
R47833 PAD.n2336 PAD.n2199 0.019716
R47834 PAD.n2337 PAD.n2336 0.019716
R47835 PAD.n2335 PAD.n2334 0.019716
R47836 PAD.n2334 PAD.n2333 0.019716
R47837 PAD.n2324 PAD.n2203 0.019716
R47838 PAD.n2325 PAD.n2324 0.019716
R47839 PAD.n2323 PAD.n2322 0.019716
R47840 PAD.n2322 PAD.n2321 0.019716
R47841 PAD.n2312 PAD.n2207 0.019716
R47842 PAD.n2313 PAD.n2312 0.019716
R47843 PAD.n2311 PAD.n2310 0.019716
R47844 PAD.n2310 PAD.n2309 0.019716
R47845 PAD.n2300 PAD.n2211 0.019716
R47846 PAD.n2301 PAD.n2300 0.019716
R47847 PAD.n2299 PAD.n2298 0.019716
R47848 PAD.n2298 PAD.n2297 0.019716
R47849 PAD.n2288 PAD.n2215 0.019716
R47850 PAD.n2289 PAD.n2288 0.019716
R47851 PAD.n2287 PAD.n2286 0.019716
R47852 PAD.n2286 PAD.n2285 0.019716
R47853 PAD.n2276 PAD.n2219 0.019716
R47854 PAD.n2277 PAD.n2276 0.019716
R47855 PAD.n2275 PAD.n2274 0.019716
R47856 PAD.n2274 PAD.n2273 0.019716
R47857 PAD.n2264 PAD.n2223 0.019716
R47858 PAD.n2265 PAD.n2264 0.019716
R47859 PAD.n2263 PAD.n2262 0.019716
R47860 PAD.n2262 PAD.n2261 0.019716
R47861 PAD.n2252 PAD.n2227 0.019716
R47862 PAD.n2253 PAD.n2252 0.019716
R47863 PAD.n2251 PAD.n2250 0.019716
R47864 PAD.n2250 PAD.n2249 0.019716
R47865 PAD.n2240 PAD.n2231 0.019716
R47866 PAD.n2241 PAD.n2240 0.019716
R47867 PAD.n2239 PAD.n2238 0.019716
R47868 PAD.n2238 PAD.n2237 0.019716
R47869 PAD.n2827 PAD.n2500 0.019716
R47870 PAD.n2826 PAD.n2825 0.019716
R47871 PAD.n2825 PAD.n2824 0.019716
R47872 PAD.n2815 PAD.n2501 0.019716
R47873 PAD.n2816 PAD.n2815 0.019716
R47874 PAD.n2814 PAD.n2813 0.019716
R47875 PAD.n2813 PAD.n2812 0.019716
R47876 PAD.n2803 PAD.n2506 0.019716
R47877 PAD.n2804 PAD.n2803 0.019716
R47878 PAD.n2802 PAD.n2801 0.019716
R47879 PAD.n2801 PAD.n2800 0.019716
R47880 PAD.n2791 PAD.n2510 0.019716
R47881 PAD.n2792 PAD.n2791 0.019716
R47882 PAD.n2790 PAD.n2789 0.019716
R47883 PAD.n2789 PAD.n2788 0.019716
R47884 PAD.n2779 PAD.n2514 0.019716
R47885 PAD.n2780 PAD.n2779 0.019716
R47886 PAD.n2778 PAD.n2777 0.019716
R47887 PAD.n2777 PAD.n2776 0.019716
R47888 PAD.n2767 PAD.n2518 0.019716
R47889 PAD.n2768 PAD.n2767 0.019716
R47890 PAD.n2766 PAD.n2765 0.019716
R47891 PAD.n2765 PAD.n2764 0.019716
R47892 PAD.n2755 PAD.n2522 0.019716
R47893 PAD.n2756 PAD.n2755 0.019716
R47894 PAD.n2754 PAD.n2753 0.019716
R47895 PAD.n2753 PAD.n2752 0.019716
R47896 PAD.n2743 PAD.n2526 0.019716
R47897 PAD.n2744 PAD.n2743 0.019716
R47898 PAD.n2742 PAD.n2741 0.019716
R47899 PAD.n2741 PAD.n2740 0.019716
R47900 PAD.n2731 PAD.n2530 0.019716
R47901 PAD.n2732 PAD.n2731 0.019716
R47902 PAD.n2730 PAD.n2729 0.019716
R47903 PAD.n2729 PAD.n2728 0.019716
R47904 PAD.n2719 PAD.n2534 0.019716
R47905 PAD.n2720 PAD.n2719 0.019716
R47906 PAD.n2718 PAD.n2717 0.019716
R47907 PAD.n2717 PAD.n2716 0.019716
R47908 PAD.n2707 PAD.n2538 0.019716
R47909 PAD.n2708 PAD.n2707 0.019716
R47910 PAD.n2706 PAD.n2705 0.019716
R47911 PAD.n2705 PAD.n2704 0.019716
R47912 PAD.n2695 PAD.n2542 0.019716
R47913 PAD.n2696 PAD.n2695 0.019716
R47914 PAD.n2694 PAD.n2693 0.019716
R47915 PAD.n2693 PAD.n2692 0.019716
R47916 PAD.n2683 PAD.n2546 0.019716
R47917 PAD.n2684 PAD.n2683 0.019716
R47918 PAD.n2682 PAD.n2681 0.019716
R47919 PAD.n2681 PAD.n2680 0.019716
R47920 PAD.n2671 PAD.n2550 0.019716
R47921 PAD.n2672 PAD.n2671 0.019716
R47922 PAD.n2670 PAD.n2669 0.019716
R47923 PAD.n2669 PAD.n2668 0.019716
R47924 PAD.n2659 PAD.n2554 0.019716
R47925 PAD.n2660 PAD.n2659 0.019716
R47926 PAD.n2658 PAD.n2657 0.019716
R47927 PAD.n2657 PAD.n2656 0.019716
R47928 PAD.n2647 PAD.n2558 0.019716
R47929 PAD.n2648 PAD.n2647 0.019716
R47930 PAD.n2646 PAD.n2645 0.019716
R47931 PAD.n2645 PAD.n2644 0.019716
R47932 PAD.n2635 PAD.n2562 0.019716
R47933 PAD.n2636 PAD.n2635 0.019716
R47934 PAD.n2634 PAD.n2633 0.019716
R47935 PAD.n2633 PAD.n2632 0.019716
R47936 PAD.n2623 PAD.n2566 0.019716
R47937 PAD.n2624 PAD.n2623 0.019716
R47938 PAD.n2622 PAD.n2621 0.019716
R47939 PAD.n2621 PAD.n2620 0.019716
R47940 PAD.n2611 PAD.n2570 0.019716
R47941 PAD.n2612 PAD.n2611 0.019716
R47942 PAD.n2610 PAD.n2609 0.019716
R47943 PAD.n2609 PAD.n2608 0.019716
R47944 PAD.n2599 PAD.n2574 0.019716
R47945 PAD.n2600 PAD.n2599 0.019716
R47946 PAD.n2598 PAD.n2597 0.019716
R47947 PAD.n2597 PAD.n2596 0.019716
R47948 PAD.n2587 PAD.n2578 0.019716
R47949 PAD.n2588 PAD.n2587 0.019716
R47950 PAD.n2586 PAD.n2585 0.019716
R47951 PAD.n2585 PAD.n2584 0.019716
R47952 PAD.n9117 PAD.n9116 0.019716
R47953 PAD.n8841 PAD.n2875 0.019716
R47954 PAD.n8841 PAD.n8840 0.019716
R47955 PAD.n9110 PAD.n2874 0.019716
R47956 PAD.n9110 PAD.n9109 0.019716
R47957 PAD.n8846 PAD.n2873 0.019716
R47958 PAD.n8846 PAD.n8845 0.019716
R47959 PAD.n9101 PAD.n2872 0.019716
R47960 PAD.n9101 PAD.n9100 0.019716
R47961 PAD.n8851 PAD.n2871 0.019716
R47962 PAD.n8851 PAD.n8850 0.019716
R47963 PAD.n9092 PAD.n2870 0.019716
R47964 PAD.n9092 PAD.n9091 0.019716
R47965 PAD.n8856 PAD.n2869 0.019716
R47966 PAD.n8856 PAD.n8855 0.019716
R47967 PAD.n9083 PAD.n2868 0.019716
R47968 PAD.n9083 PAD.n9082 0.019716
R47969 PAD.n8861 PAD.n2867 0.019716
R47970 PAD.n8861 PAD.n8860 0.019716
R47971 PAD.n9074 PAD.n2866 0.019716
R47972 PAD.n9074 PAD.n9073 0.019716
R47973 PAD.n8866 PAD.n2865 0.019716
R47974 PAD.n8866 PAD.n8865 0.019716
R47975 PAD.n9065 PAD.n2864 0.019716
R47976 PAD.n9065 PAD.n9064 0.019716
R47977 PAD.n8871 PAD.n2863 0.019716
R47978 PAD.n8871 PAD.n8870 0.019716
R47979 PAD.n9056 PAD.n2862 0.019716
R47980 PAD.n9056 PAD.n9055 0.019716
R47981 PAD.n8876 PAD.n2861 0.019716
R47982 PAD.n8876 PAD.n8875 0.019716
R47983 PAD.n9047 PAD.n2860 0.019716
R47984 PAD.n9047 PAD.n9046 0.019716
R47985 PAD.n8881 PAD.n2859 0.019716
R47986 PAD.n8881 PAD.n8880 0.019716
R47987 PAD.n9038 PAD.n2858 0.019716
R47988 PAD.n9038 PAD.n9037 0.019716
R47989 PAD.n8886 PAD.n2857 0.019716
R47990 PAD.n8886 PAD.n8885 0.019716
R47991 PAD.n9029 PAD.n2856 0.019716
R47992 PAD.n9029 PAD.n9028 0.019716
R47993 PAD.n8891 PAD.n2855 0.019716
R47994 PAD.n8891 PAD.n8890 0.019716
R47995 PAD.n9020 PAD.n2854 0.019716
R47996 PAD.n9020 PAD.n9019 0.019716
R47997 PAD.n8896 PAD.n2853 0.019716
R47998 PAD.n8896 PAD.n8895 0.019716
R47999 PAD.n9011 PAD.n2852 0.019716
R48000 PAD.n9011 PAD.n9010 0.019716
R48001 PAD.n8901 PAD.n2851 0.019716
R48002 PAD.n8901 PAD.n8900 0.019716
R48003 PAD.n9002 PAD.n2850 0.019716
R48004 PAD.n9002 PAD.n9001 0.019716
R48005 PAD.n8906 PAD.n2849 0.019716
R48006 PAD.n8906 PAD.n8905 0.019716
R48007 PAD.n8993 PAD.n2848 0.019716
R48008 PAD.n8993 PAD.n8992 0.019716
R48009 PAD.n8911 PAD.n2847 0.019716
R48010 PAD.n8911 PAD.n8910 0.019716
R48011 PAD.n8984 PAD.n2846 0.019716
R48012 PAD.n8984 PAD.n8983 0.019716
R48013 PAD.n8916 PAD.n2845 0.019716
R48014 PAD.n8916 PAD.n8915 0.019716
R48015 PAD.n8975 PAD.n2844 0.019716
R48016 PAD.n8975 PAD.n8974 0.019716
R48017 PAD.n8921 PAD.n2843 0.019716
R48018 PAD.n8921 PAD.n8920 0.019716
R48019 PAD.n8966 PAD.n2842 0.019716
R48020 PAD.n8966 PAD.n8965 0.019716
R48021 PAD.n8926 PAD.n2841 0.019716
R48022 PAD.n8926 PAD.n8925 0.019716
R48023 PAD.n8957 PAD.n2840 0.019716
R48024 PAD.n8957 PAD.n8956 0.019716
R48025 PAD.n8931 PAD.n2839 0.019716
R48026 PAD.n8931 PAD.n8930 0.019716
R48027 PAD.n8948 PAD.n2838 0.019716
R48028 PAD.n8948 PAD.n8947 0.019716
R48029 PAD.n8936 PAD.n2837 0.019716
R48030 PAD.n8936 PAD.n8935 0.019716
R48031 PAD.n8939 PAD.n2836 0.019716
R48032 PAD.n8939 PAD.n8938 0.019716
R48033 PAD.n9137 PAD.n2835 0.019716
R48034 PAD.n9138 PAD.n9137 0.019716
R48035 PAD.n8820 PAD.n8528 0.019716
R48036 PAD.n8813 PAD.n8812 0.019716
R48037 PAD.n8813 PAD.n2945 0.019716
R48038 PAD.n8809 PAD.n8808 0.019716
R48039 PAD.n8808 PAD.n2944 0.019716
R48040 PAD.n8802 PAD.n8801 0.019716
R48041 PAD.n8802 PAD.n2943 0.019716
R48042 PAD.n8797 PAD.n8796 0.019716
R48043 PAD.n8796 PAD.n2942 0.019716
R48044 PAD.n8790 PAD.n8789 0.019716
R48045 PAD.n8790 PAD.n2941 0.019716
R48046 PAD.n8785 PAD.n8784 0.019716
R48047 PAD.n8784 PAD.n2940 0.019716
R48048 PAD.n8778 PAD.n8777 0.019716
R48049 PAD.n8778 PAD.n2939 0.019716
R48050 PAD.n8773 PAD.n8772 0.019716
R48051 PAD.n8772 PAD.n2938 0.019716
R48052 PAD.n8766 PAD.n8765 0.019716
R48053 PAD.n8766 PAD.n2937 0.019716
R48054 PAD.n8761 PAD.n8760 0.019716
R48055 PAD.n8760 PAD.n2936 0.019716
R48056 PAD.n8754 PAD.n8753 0.019716
R48057 PAD.n8754 PAD.n2935 0.019716
R48058 PAD.n8749 PAD.n8748 0.019716
R48059 PAD.n8748 PAD.n2934 0.019716
R48060 PAD.n8742 PAD.n8741 0.019716
R48061 PAD.n8742 PAD.n2933 0.019716
R48062 PAD.n8737 PAD.n8736 0.019716
R48063 PAD.n8736 PAD.n2932 0.019716
R48064 PAD.n8730 PAD.n8729 0.019716
R48065 PAD.n8730 PAD.n2931 0.019716
R48066 PAD.n8725 PAD.n8724 0.019716
R48067 PAD.n8724 PAD.n2930 0.019716
R48068 PAD.n8718 PAD.n8717 0.019716
R48069 PAD.n8718 PAD.n2929 0.019716
R48070 PAD.n8713 PAD.n8712 0.019716
R48071 PAD.n8712 PAD.n2928 0.019716
R48072 PAD.n8706 PAD.n8705 0.019716
R48073 PAD.n8706 PAD.n2927 0.019716
R48074 PAD.n8701 PAD.n8700 0.019716
R48075 PAD.n8700 PAD.n2926 0.019716
R48076 PAD.n8694 PAD.n8693 0.019716
R48077 PAD.n8694 PAD.n2925 0.019716
R48078 PAD.n8689 PAD.n8688 0.019716
R48079 PAD.n8688 PAD.n2924 0.019716
R48080 PAD.n8682 PAD.n8681 0.019716
R48081 PAD.n8682 PAD.n2923 0.019716
R48082 PAD.n8677 PAD.n8676 0.019716
R48083 PAD.n8676 PAD.n2922 0.019716
R48084 PAD.n8670 PAD.n8669 0.019716
R48085 PAD.n8670 PAD.n2921 0.019716
R48086 PAD.n8665 PAD.n8664 0.019716
R48087 PAD.n8664 PAD.n2920 0.019716
R48088 PAD.n8658 PAD.n8657 0.019716
R48089 PAD.n8658 PAD.n2919 0.019716
R48090 PAD.n8653 PAD.n8652 0.019716
R48091 PAD.n8652 PAD.n2918 0.019716
R48092 PAD.n8646 PAD.n8645 0.019716
R48093 PAD.n8646 PAD.n2917 0.019716
R48094 PAD.n8641 PAD.n8640 0.019716
R48095 PAD.n8640 PAD.n2916 0.019716
R48096 PAD.n8634 PAD.n8633 0.019716
R48097 PAD.n8634 PAD.n2915 0.019716
R48098 PAD.n8629 PAD.n8628 0.019716
R48099 PAD.n8628 PAD.n2914 0.019716
R48100 PAD.n8622 PAD.n8621 0.019716
R48101 PAD.n8622 PAD.n2913 0.019716
R48102 PAD.n8617 PAD.n8616 0.019716
R48103 PAD.n8616 PAD.n2912 0.019716
R48104 PAD.n8610 PAD.n8609 0.019716
R48105 PAD.n8610 PAD.n2911 0.019716
R48106 PAD.n8605 PAD.n8604 0.019716
R48107 PAD.n8604 PAD.n2910 0.019716
R48108 PAD.n8598 PAD.n8597 0.019716
R48109 PAD.n8598 PAD.n2909 0.019716
R48110 PAD.n8593 PAD.n8592 0.019716
R48111 PAD.n8592 PAD.n2908 0.019716
R48112 PAD.n8586 PAD.n8585 0.019716
R48113 PAD.n8586 PAD.n2907 0.019716
R48114 PAD.n8581 PAD.n8580 0.019716
R48115 PAD.n8580 PAD.n2906 0.019716
R48116 PAD.n8574 PAD.n8573 0.019716
R48117 PAD.n8574 PAD.n2905 0.019716
R48118 PAD.n3039 PAD.n3038 0.019716
R48119 PAD.n3046 PAD.n2993 0.019716
R48120 PAD.n3047 PAD.n3046 0.019716
R48121 PAD.n3052 PAD.n2992 0.019716
R48122 PAD.n3052 PAD.n3051 0.019716
R48123 PAD.n3058 PAD.n2991 0.019716
R48124 PAD.n3059 PAD.n3058 0.019716
R48125 PAD.n3064 PAD.n2990 0.019716
R48126 PAD.n3064 PAD.n3063 0.019716
R48127 PAD.n3070 PAD.n2989 0.019716
R48128 PAD.n3071 PAD.n3070 0.019716
R48129 PAD.n3076 PAD.n2988 0.019716
R48130 PAD.n3076 PAD.n3075 0.019716
R48131 PAD.n3082 PAD.n2987 0.019716
R48132 PAD.n3083 PAD.n3082 0.019716
R48133 PAD.n3088 PAD.n2986 0.019716
R48134 PAD.n3088 PAD.n3087 0.019716
R48135 PAD.n3094 PAD.n2985 0.019716
R48136 PAD.n3095 PAD.n3094 0.019716
R48137 PAD.n3100 PAD.n2984 0.019716
R48138 PAD.n3100 PAD.n3099 0.019716
R48139 PAD.n3106 PAD.n2983 0.019716
R48140 PAD.n3107 PAD.n3106 0.019716
R48141 PAD.n3112 PAD.n2982 0.019716
R48142 PAD.n3112 PAD.n3111 0.019716
R48143 PAD.n3118 PAD.n2981 0.019716
R48144 PAD.n3119 PAD.n3118 0.019716
R48145 PAD.n3124 PAD.n2980 0.019716
R48146 PAD.n3124 PAD.n3123 0.019716
R48147 PAD.n3130 PAD.n2979 0.019716
R48148 PAD.n3131 PAD.n3130 0.019716
R48149 PAD.n3136 PAD.n2978 0.019716
R48150 PAD.n3136 PAD.n3135 0.019716
R48151 PAD.n3142 PAD.n2977 0.019716
R48152 PAD.n3143 PAD.n3142 0.019716
R48153 PAD.n3148 PAD.n2976 0.019716
R48154 PAD.n3148 PAD.n3147 0.019716
R48155 PAD.n3154 PAD.n2975 0.019716
R48156 PAD.n3155 PAD.n3154 0.019716
R48157 PAD.n3160 PAD.n2974 0.019716
R48158 PAD.n3160 PAD.n3159 0.019716
R48159 PAD.n3166 PAD.n2973 0.019716
R48160 PAD.n3167 PAD.n3166 0.019716
R48161 PAD.n3172 PAD.n2972 0.019716
R48162 PAD.n3172 PAD.n3171 0.019716
R48163 PAD.n3178 PAD.n2971 0.019716
R48164 PAD.n3179 PAD.n3178 0.019716
R48165 PAD.n3184 PAD.n2970 0.019716
R48166 PAD.n3184 PAD.n3183 0.019716
R48167 PAD.n3190 PAD.n2969 0.019716
R48168 PAD.n3191 PAD.n3190 0.019716
R48169 PAD.n3196 PAD.n2968 0.019716
R48170 PAD.n3196 PAD.n3195 0.019716
R48171 PAD.n3202 PAD.n2967 0.019716
R48172 PAD.n3203 PAD.n3202 0.019716
R48173 PAD.n3208 PAD.n2966 0.019716
R48174 PAD.n3208 PAD.n3207 0.019716
R48175 PAD.n3214 PAD.n2965 0.019716
R48176 PAD.n3215 PAD.n3214 0.019716
R48177 PAD.n3220 PAD.n2964 0.019716
R48178 PAD.n3220 PAD.n3219 0.019716
R48179 PAD.n3226 PAD.n2963 0.019716
R48180 PAD.n3227 PAD.n3226 0.019716
R48181 PAD.n3232 PAD.n2962 0.019716
R48182 PAD.n3232 PAD.n3231 0.019716
R48183 PAD.n3238 PAD.n2961 0.019716
R48184 PAD.n3239 PAD.n3238 0.019716
R48185 PAD.n3244 PAD.n2960 0.019716
R48186 PAD.n3244 PAD.n3243 0.019716
R48187 PAD.n3250 PAD.n2959 0.019716
R48188 PAD.n3251 PAD.n3250 0.019716
R48189 PAD.n3256 PAD.n2958 0.019716
R48190 PAD.n3256 PAD.n3255 0.019716
R48191 PAD.n3262 PAD.n2957 0.019716
R48192 PAD.n3263 PAD.n3262 0.019716
R48193 PAD.n3268 PAD.n2956 0.019716
R48194 PAD.n3268 PAD.n3267 0.019716
R48195 PAD.n3274 PAD.n2955 0.019716
R48196 PAD.n3275 PAD.n3274 0.019716
R48197 PAD.n3280 PAD.n2954 0.019716
R48198 PAD.n3280 PAD.n3279 0.019716
R48199 PAD.n8514 PAD.n2953 0.019716
R48200 PAD.n8515 PAD.n8514 0.019716
R48201 PAD.n3384 PAD.n3383 0.019716
R48202 PAD.n3391 PAD.n3337 0.019716
R48203 PAD.n3392 PAD.n3391 0.019716
R48204 PAD.n3397 PAD.n3336 0.019716
R48205 PAD.n3397 PAD.n3396 0.019716
R48206 PAD.n3403 PAD.n3335 0.019716
R48207 PAD.n3404 PAD.n3403 0.019716
R48208 PAD.n3409 PAD.n3334 0.019716
R48209 PAD.n3409 PAD.n3408 0.019716
R48210 PAD.n3415 PAD.n3333 0.019716
R48211 PAD.n3416 PAD.n3415 0.019716
R48212 PAD.n3421 PAD.n3332 0.019716
R48213 PAD.n3421 PAD.n3420 0.019716
R48214 PAD.n3427 PAD.n3331 0.019716
R48215 PAD.n3428 PAD.n3427 0.019716
R48216 PAD.n3433 PAD.n3330 0.019716
R48217 PAD.n3433 PAD.n3432 0.019716
R48218 PAD.n3439 PAD.n3329 0.019716
R48219 PAD.n3440 PAD.n3439 0.019716
R48220 PAD.n3445 PAD.n3328 0.019716
R48221 PAD.n3445 PAD.n3444 0.019716
R48222 PAD.n3451 PAD.n3327 0.019716
R48223 PAD.n3452 PAD.n3451 0.019716
R48224 PAD.n3457 PAD.n3326 0.019716
R48225 PAD.n3457 PAD.n3456 0.019716
R48226 PAD.n3463 PAD.n3325 0.019716
R48227 PAD.n3464 PAD.n3463 0.019716
R48228 PAD.n3469 PAD.n3324 0.019716
R48229 PAD.n3469 PAD.n3468 0.019716
R48230 PAD.n3475 PAD.n3323 0.019716
R48231 PAD.n3476 PAD.n3475 0.019716
R48232 PAD.n3481 PAD.n3322 0.019716
R48233 PAD.n3481 PAD.n3480 0.019716
R48234 PAD.n3487 PAD.n3321 0.019716
R48235 PAD.n3488 PAD.n3487 0.019716
R48236 PAD.n3493 PAD.n3320 0.019716
R48237 PAD.n3493 PAD.n3492 0.019716
R48238 PAD.n3499 PAD.n3319 0.019716
R48239 PAD.n3500 PAD.n3499 0.019716
R48240 PAD.n3505 PAD.n3318 0.019716
R48241 PAD.n3505 PAD.n3504 0.019716
R48242 PAD.n3511 PAD.n3317 0.019716
R48243 PAD.n3512 PAD.n3511 0.019716
R48244 PAD.n3517 PAD.n3316 0.019716
R48245 PAD.n3517 PAD.n3516 0.019716
R48246 PAD.n3523 PAD.n3315 0.019716
R48247 PAD.n3524 PAD.n3523 0.019716
R48248 PAD.n3529 PAD.n3314 0.019716
R48249 PAD.n3529 PAD.n3528 0.019716
R48250 PAD.n3535 PAD.n3313 0.019716
R48251 PAD.n3536 PAD.n3535 0.019716
R48252 PAD.n3541 PAD.n3312 0.019716
R48253 PAD.n3541 PAD.n3540 0.019716
R48254 PAD.n3547 PAD.n3311 0.019716
R48255 PAD.n3548 PAD.n3547 0.019716
R48256 PAD.n3553 PAD.n3310 0.019716
R48257 PAD.n3553 PAD.n3552 0.019716
R48258 PAD.n3559 PAD.n3309 0.019716
R48259 PAD.n3560 PAD.n3559 0.019716
R48260 PAD.n3565 PAD.n3308 0.019716
R48261 PAD.n3565 PAD.n3564 0.019716
R48262 PAD.n3571 PAD.n3307 0.019716
R48263 PAD.n3572 PAD.n3571 0.019716
R48264 PAD.n3577 PAD.n3306 0.019716
R48265 PAD.n3577 PAD.n3576 0.019716
R48266 PAD.n3583 PAD.n3305 0.019716
R48267 PAD.n3584 PAD.n3583 0.019716
R48268 PAD.n3589 PAD.n3304 0.019716
R48269 PAD.n3589 PAD.n3588 0.019716
R48270 PAD.n3595 PAD.n3303 0.019716
R48271 PAD.n3596 PAD.n3595 0.019716
R48272 PAD.n3601 PAD.n3302 0.019716
R48273 PAD.n3601 PAD.n3600 0.019716
R48274 PAD.n3607 PAD.n3301 0.019716
R48275 PAD.n3608 PAD.n3607 0.019716
R48276 PAD.n3613 PAD.n3300 0.019716
R48277 PAD.n3613 PAD.n3612 0.019716
R48278 PAD.n3619 PAD.n3299 0.019716
R48279 PAD.n3620 PAD.n3619 0.019716
R48280 PAD.n3625 PAD.n3298 0.019716
R48281 PAD.n3625 PAD.n3624 0.019716
R48282 PAD.n8489 PAD.n3297 0.019716
R48283 PAD.n8490 PAD.n8489 0.019716
R48284 PAD.n3729 PAD.n3728 0.019716
R48285 PAD.n3736 PAD.n3682 0.019716
R48286 PAD.n3737 PAD.n3736 0.019716
R48287 PAD.n3742 PAD.n3681 0.019716
R48288 PAD.n3742 PAD.n3741 0.019716
R48289 PAD.n3748 PAD.n3680 0.019716
R48290 PAD.n3749 PAD.n3748 0.019716
R48291 PAD.n3754 PAD.n3679 0.019716
R48292 PAD.n3754 PAD.n3753 0.019716
R48293 PAD.n3760 PAD.n3678 0.019716
R48294 PAD.n3761 PAD.n3760 0.019716
R48295 PAD.n3766 PAD.n3677 0.019716
R48296 PAD.n3766 PAD.n3765 0.019716
R48297 PAD.n3772 PAD.n3676 0.019716
R48298 PAD.n3773 PAD.n3772 0.019716
R48299 PAD.n3778 PAD.n3675 0.019716
R48300 PAD.n3778 PAD.n3777 0.019716
R48301 PAD.n3784 PAD.n3674 0.019716
R48302 PAD.n3785 PAD.n3784 0.019716
R48303 PAD.n3790 PAD.n3673 0.019716
R48304 PAD.n3790 PAD.n3789 0.019716
R48305 PAD.n3796 PAD.n3672 0.019716
R48306 PAD.n3797 PAD.n3796 0.019716
R48307 PAD.n3802 PAD.n3671 0.019716
R48308 PAD.n3802 PAD.n3801 0.019716
R48309 PAD.n3808 PAD.n3670 0.019716
R48310 PAD.n3809 PAD.n3808 0.019716
R48311 PAD.n3814 PAD.n3669 0.019716
R48312 PAD.n3814 PAD.n3813 0.019716
R48313 PAD.n3820 PAD.n3668 0.019716
R48314 PAD.n3821 PAD.n3820 0.019716
R48315 PAD.n3826 PAD.n3667 0.019716
R48316 PAD.n3826 PAD.n3825 0.019716
R48317 PAD.n3832 PAD.n3666 0.019716
R48318 PAD.n3833 PAD.n3832 0.019716
R48319 PAD.n3838 PAD.n3665 0.019716
R48320 PAD.n3838 PAD.n3837 0.019716
R48321 PAD.n3844 PAD.n3664 0.019716
R48322 PAD.n3845 PAD.n3844 0.019716
R48323 PAD.n3850 PAD.n3663 0.019716
R48324 PAD.n3850 PAD.n3849 0.019716
R48325 PAD.n3856 PAD.n3662 0.019716
R48326 PAD.n3857 PAD.n3856 0.019716
R48327 PAD.n3862 PAD.n3661 0.019716
R48328 PAD.n3862 PAD.n3861 0.019716
R48329 PAD.n3868 PAD.n3660 0.019716
R48330 PAD.n3869 PAD.n3868 0.019716
R48331 PAD.n3874 PAD.n3659 0.019716
R48332 PAD.n3874 PAD.n3873 0.019716
R48333 PAD.n3880 PAD.n3658 0.019716
R48334 PAD.n3881 PAD.n3880 0.019716
R48335 PAD.n3886 PAD.n3657 0.019716
R48336 PAD.n3886 PAD.n3885 0.019716
R48337 PAD.n3892 PAD.n3656 0.019716
R48338 PAD.n3893 PAD.n3892 0.019716
R48339 PAD.n3898 PAD.n3655 0.019716
R48340 PAD.n3898 PAD.n3897 0.019716
R48341 PAD.n3904 PAD.n3654 0.019716
R48342 PAD.n3905 PAD.n3904 0.019716
R48343 PAD.n3910 PAD.n3653 0.019716
R48344 PAD.n3910 PAD.n3909 0.019716
R48345 PAD.n3916 PAD.n3652 0.019716
R48346 PAD.n3917 PAD.n3916 0.019716
R48347 PAD.n3922 PAD.n3651 0.019716
R48348 PAD.n3922 PAD.n3921 0.019716
R48349 PAD.n3928 PAD.n3650 0.019716
R48350 PAD.n3929 PAD.n3928 0.019716
R48351 PAD.n3934 PAD.n3649 0.019716
R48352 PAD.n3934 PAD.n3933 0.019716
R48353 PAD.n3940 PAD.n3648 0.019716
R48354 PAD.n3941 PAD.n3940 0.019716
R48355 PAD.n3946 PAD.n3647 0.019716
R48356 PAD.n3946 PAD.n3945 0.019716
R48357 PAD.n3952 PAD.n3646 0.019716
R48358 PAD.n3953 PAD.n3952 0.019716
R48359 PAD.n3958 PAD.n3645 0.019716
R48360 PAD.n3958 PAD.n3957 0.019716
R48361 PAD.n3964 PAD.n3644 0.019716
R48362 PAD.n3965 PAD.n3964 0.019716
R48363 PAD.n3970 PAD.n3643 0.019716
R48364 PAD.n3970 PAD.n3969 0.019716
R48365 PAD.n8465 PAD.n3642 0.019716
R48366 PAD.n8466 PAD.n8465 0.019716
R48367 PAD.n4070 PAD.n4069 0.019716
R48368 PAD.n4077 PAD.n4024 0.019716
R48369 PAD.n4078 PAD.n4077 0.019716
R48370 PAD.n4083 PAD.n4023 0.019716
R48371 PAD.n4083 PAD.n4082 0.019716
R48372 PAD.n4089 PAD.n4022 0.019716
R48373 PAD.n4090 PAD.n4089 0.019716
R48374 PAD.n4095 PAD.n4021 0.019716
R48375 PAD.n4095 PAD.n4094 0.019716
R48376 PAD.n4101 PAD.n4020 0.019716
R48377 PAD.n4102 PAD.n4101 0.019716
R48378 PAD.n4107 PAD.n4019 0.019716
R48379 PAD.n4107 PAD.n4106 0.019716
R48380 PAD.n4113 PAD.n4018 0.019716
R48381 PAD.n4114 PAD.n4113 0.019716
R48382 PAD.n4119 PAD.n4017 0.019716
R48383 PAD.n4119 PAD.n4118 0.019716
R48384 PAD.n4125 PAD.n4016 0.019716
R48385 PAD.n4126 PAD.n4125 0.019716
R48386 PAD.n4131 PAD.n4015 0.019716
R48387 PAD.n4131 PAD.n4130 0.019716
R48388 PAD.n4137 PAD.n4014 0.019716
R48389 PAD.n4138 PAD.n4137 0.019716
R48390 PAD.n4143 PAD.n4013 0.019716
R48391 PAD.n4143 PAD.n4142 0.019716
R48392 PAD.n4149 PAD.n4012 0.019716
R48393 PAD.n4150 PAD.n4149 0.019716
R48394 PAD.n4155 PAD.n4011 0.019716
R48395 PAD.n4155 PAD.n4154 0.019716
R48396 PAD.n4161 PAD.n4010 0.019716
R48397 PAD.n4162 PAD.n4161 0.019716
R48398 PAD.n4167 PAD.n4009 0.019716
R48399 PAD.n4167 PAD.n4166 0.019716
R48400 PAD.n4173 PAD.n4008 0.019716
R48401 PAD.n4174 PAD.n4173 0.019716
R48402 PAD.n4179 PAD.n4007 0.019716
R48403 PAD.n4179 PAD.n4178 0.019716
R48404 PAD.n4185 PAD.n4006 0.019716
R48405 PAD.n4186 PAD.n4185 0.019716
R48406 PAD.n4191 PAD.n4005 0.019716
R48407 PAD.n4191 PAD.n4190 0.019716
R48408 PAD.n4197 PAD.n4004 0.019716
R48409 PAD.n4198 PAD.n4197 0.019716
R48410 PAD.n4203 PAD.n4003 0.019716
R48411 PAD.n4203 PAD.n4202 0.019716
R48412 PAD.n4209 PAD.n4002 0.019716
R48413 PAD.n4210 PAD.n4209 0.019716
R48414 PAD.n4215 PAD.n4001 0.019716
R48415 PAD.n4215 PAD.n4214 0.019716
R48416 PAD.n4221 PAD.n4000 0.019716
R48417 PAD.n4222 PAD.n4221 0.019716
R48418 PAD.n4227 PAD.n3999 0.019716
R48419 PAD.n4227 PAD.n4226 0.019716
R48420 PAD.n4233 PAD.n3998 0.019716
R48421 PAD.n4234 PAD.n4233 0.019716
R48422 PAD.n4239 PAD.n3997 0.019716
R48423 PAD.n4239 PAD.n4238 0.019716
R48424 PAD.n4245 PAD.n3996 0.019716
R48425 PAD.n4246 PAD.n4245 0.019716
R48426 PAD.n4251 PAD.n3995 0.019716
R48427 PAD.n4251 PAD.n4250 0.019716
R48428 PAD.n4257 PAD.n3994 0.019716
R48429 PAD.n4258 PAD.n4257 0.019716
R48430 PAD.n4263 PAD.n3993 0.019716
R48431 PAD.n4263 PAD.n4262 0.019716
R48432 PAD.n4269 PAD.n3992 0.019716
R48433 PAD.n4270 PAD.n4269 0.019716
R48434 PAD.n4275 PAD.n3991 0.019716
R48435 PAD.n4275 PAD.n4274 0.019716
R48436 PAD.n4281 PAD.n3990 0.019716
R48437 PAD.n4282 PAD.n4281 0.019716
R48438 PAD.n4287 PAD.n3989 0.019716
R48439 PAD.n4287 PAD.n4286 0.019716
R48440 PAD.n4293 PAD.n3988 0.019716
R48441 PAD.n4294 PAD.n4293 0.019716
R48442 PAD.n4299 PAD.n3987 0.019716
R48443 PAD.n4299 PAD.n4298 0.019716
R48444 PAD.n4305 PAD.n3986 0.019716
R48445 PAD.n4306 PAD.n4305 0.019716
R48446 PAD.n4311 PAD.n3985 0.019716
R48447 PAD.n4311 PAD.n4310 0.019716
R48448 PAD.n8441 PAD.n3984 0.019716
R48449 PAD.n8442 PAD.n8441 0.019716
R48450 PAD.n4422 PAD.n4421 0.019716
R48451 PAD.n4426 PAD.n4423 0.019716
R48452 PAD.n4426 PAD.n4425 0.019716
R48453 PAD.n4432 PAD.n4415 0.019716
R48454 PAD.n4433 PAD.n4432 0.019716
R48455 PAD.n4438 PAD.n4435 0.019716
R48456 PAD.n4438 PAD.n4437 0.019716
R48457 PAD.n4444 PAD.n4411 0.019716
R48458 PAD.n4445 PAD.n4444 0.019716
R48459 PAD.n4450 PAD.n4447 0.019716
R48460 PAD.n4450 PAD.n4449 0.019716
R48461 PAD.n4456 PAD.n4407 0.019716
R48462 PAD.n4457 PAD.n4456 0.019716
R48463 PAD.n4462 PAD.n4459 0.019716
R48464 PAD.n4462 PAD.n4461 0.019716
R48465 PAD.n4468 PAD.n4403 0.019716
R48466 PAD.n4469 PAD.n4468 0.019716
R48467 PAD.n4474 PAD.n4471 0.019716
R48468 PAD.n4474 PAD.n4473 0.019716
R48469 PAD.n4480 PAD.n4399 0.019716
R48470 PAD.n4481 PAD.n4480 0.019716
R48471 PAD.n4486 PAD.n4483 0.019716
R48472 PAD.n4486 PAD.n4485 0.019716
R48473 PAD.n4492 PAD.n4395 0.019716
R48474 PAD.n4493 PAD.n4492 0.019716
R48475 PAD.n4498 PAD.n4495 0.019716
R48476 PAD.n4498 PAD.n4497 0.019716
R48477 PAD.n4504 PAD.n4391 0.019716
R48478 PAD.n4505 PAD.n4504 0.019716
R48479 PAD.n4510 PAD.n4507 0.019716
R48480 PAD.n4510 PAD.n4509 0.019716
R48481 PAD.n4516 PAD.n4387 0.019716
R48482 PAD.n4517 PAD.n4516 0.019716
R48483 PAD.n4522 PAD.n4519 0.019716
R48484 PAD.n4522 PAD.n4521 0.019716
R48485 PAD.n4528 PAD.n4383 0.019716
R48486 PAD.n4529 PAD.n4528 0.019716
R48487 PAD.n4534 PAD.n4531 0.019716
R48488 PAD.n4534 PAD.n4533 0.019716
R48489 PAD.n4540 PAD.n4379 0.019716
R48490 PAD.n4541 PAD.n4540 0.019716
R48491 PAD.n4546 PAD.n4543 0.019716
R48492 PAD.n4546 PAD.n4545 0.019716
R48493 PAD.n4552 PAD.n4375 0.019716
R48494 PAD.n4553 PAD.n4552 0.019716
R48495 PAD.n4558 PAD.n4555 0.019716
R48496 PAD.n4558 PAD.n4557 0.019716
R48497 PAD.n4564 PAD.n4371 0.019716
R48498 PAD.n4565 PAD.n4564 0.019716
R48499 PAD.n4570 PAD.n4567 0.019716
R48500 PAD.n4570 PAD.n4569 0.019716
R48501 PAD.n4576 PAD.n4367 0.019716
R48502 PAD.n4577 PAD.n4576 0.019716
R48503 PAD.n4582 PAD.n4579 0.019716
R48504 PAD.n4582 PAD.n4581 0.019716
R48505 PAD.n4588 PAD.n4363 0.019716
R48506 PAD.n4589 PAD.n4588 0.019716
R48507 PAD.n4594 PAD.n4591 0.019716
R48508 PAD.n4594 PAD.n4593 0.019716
R48509 PAD.n4600 PAD.n4359 0.019716
R48510 PAD.n4601 PAD.n4600 0.019716
R48511 PAD.n4606 PAD.n4603 0.019716
R48512 PAD.n4606 PAD.n4605 0.019716
R48513 PAD.n4612 PAD.n4355 0.019716
R48514 PAD.n4613 PAD.n4612 0.019716
R48515 PAD.n4618 PAD.n4615 0.019716
R48516 PAD.n4618 PAD.n4617 0.019716
R48517 PAD.n4624 PAD.n4351 0.019716
R48518 PAD.n4625 PAD.n4624 0.019716
R48519 PAD.n4630 PAD.n4627 0.019716
R48520 PAD.n4630 PAD.n4629 0.019716
R48521 PAD.n4636 PAD.n4347 0.019716
R48522 PAD.n4637 PAD.n4636 0.019716
R48523 PAD.n4642 PAD.n4639 0.019716
R48524 PAD.n4642 PAD.n4641 0.019716
R48525 PAD.n4648 PAD.n4343 0.019716
R48526 PAD.n4649 PAD.n4648 0.019716
R48527 PAD.n4654 PAD.n4651 0.019716
R48528 PAD.n4654 PAD.n4653 0.019716
R48529 PAD.n4661 PAD.n4339 0.019716
R48530 PAD.n4662 PAD.n4661 0.019716
R48531 PAD.n4665 PAD.n4664 0.019716
R48532 PAD.n4666 PAD.n4665 0.019716
R48533 PAD.n8396 PAD.n4725 0.019716
R48534 PAD.n4727 PAD.n4726 0.019716
R48535 PAD.n4727 PAD.n4723 0.019716
R48536 PAD.n8387 PAD.n8386 0.019716
R48537 PAD.n8386 PAD.n4722 0.019716
R48538 PAD.n4732 PAD.n4731 0.019716
R48539 PAD.n4731 PAD.n4721 0.019716
R48540 PAD.n8378 PAD.n8377 0.019716
R48541 PAD.n8377 PAD.n4720 0.019716
R48542 PAD.n4737 PAD.n4736 0.019716
R48543 PAD.n4736 PAD.n4719 0.019716
R48544 PAD.n8369 PAD.n8368 0.019716
R48545 PAD.n8368 PAD.n4718 0.019716
R48546 PAD.n4742 PAD.n4741 0.019716
R48547 PAD.n4741 PAD.n4717 0.019716
R48548 PAD.n8360 PAD.n8359 0.019716
R48549 PAD.n8359 PAD.n4716 0.019716
R48550 PAD.n4747 PAD.n4746 0.019716
R48551 PAD.n4746 PAD.n4715 0.019716
R48552 PAD.n8351 PAD.n8350 0.019716
R48553 PAD.n8350 PAD.n4714 0.019716
R48554 PAD.n4752 PAD.n4751 0.019716
R48555 PAD.n4751 PAD.n4713 0.019716
R48556 PAD.n8342 PAD.n8341 0.019716
R48557 PAD.n8341 PAD.n4712 0.019716
R48558 PAD.n4757 PAD.n4756 0.019716
R48559 PAD.n4756 PAD.n4711 0.019716
R48560 PAD.n8333 PAD.n8332 0.019716
R48561 PAD.n8332 PAD.n4710 0.019716
R48562 PAD.n4762 PAD.n4761 0.019716
R48563 PAD.n4761 PAD.n4709 0.019716
R48564 PAD.n8324 PAD.n8323 0.019716
R48565 PAD.n8323 PAD.n4708 0.019716
R48566 PAD.n4767 PAD.n4766 0.019716
R48567 PAD.n4766 PAD.n4707 0.019716
R48568 PAD.n8315 PAD.n8314 0.019716
R48569 PAD.n8314 PAD.n4706 0.019716
R48570 PAD.n4772 PAD.n4771 0.019716
R48571 PAD.n4771 PAD.n4705 0.019716
R48572 PAD.n8306 PAD.n8305 0.019716
R48573 PAD.n8305 PAD.n4704 0.019716
R48574 PAD.n4777 PAD.n4776 0.019716
R48575 PAD.n4776 PAD.n4703 0.019716
R48576 PAD.n8297 PAD.n8296 0.019716
R48577 PAD.n8296 PAD.n4702 0.019716
R48578 PAD.n4782 PAD.n4781 0.019716
R48579 PAD.n4781 PAD.n4701 0.019716
R48580 PAD.n8288 PAD.n8287 0.019716
R48581 PAD.n8287 PAD.n4700 0.019716
R48582 PAD.n4787 PAD.n4786 0.019716
R48583 PAD.n4786 PAD.n4699 0.019716
R48584 PAD.n8279 PAD.n8278 0.019716
R48585 PAD.n8278 PAD.n4698 0.019716
R48586 PAD.n4792 PAD.n4791 0.019716
R48587 PAD.n4791 PAD.n4697 0.019716
R48588 PAD.n8270 PAD.n8269 0.019716
R48589 PAD.n8269 PAD.n4696 0.019716
R48590 PAD.n4797 PAD.n4796 0.019716
R48591 PAD.n4796 PAD.n4695 0.019716
R48592 PAD.n8261 PAD.n8260 0.019716
R48593 PAD.n8260 PAD.n4694 0.019716
R48594 PAD.n4802 PAD.n4801 0.019716
R48595 PAD.n4801 PAD.n4693 0.019716
R48596 PAD.n8252 PAD.n8251 0.019716
R48597 PAD.n8251 PAD.n4692 0.019716
R48598 PAD.n4807 PAD.n4806 0.019716
R48599 PAD.n4806 PAD.n4691 0.019716
R48600 PAD.n8243 PAD.n8242 0.019716
R48601 PAD.n8242 PAD.n4690 0.019716
R48602 PAD.n4812 PAD.n4811 0.019716
R48603 PAD.n4811 PAD.n4689 0.019716
R48604 PAD.n8234 PAD.n8233 0.019716
R48605 PAD.n8233 PAD.n4688 0.019716
R48606 PAD.n4817 PAD.n4816 0.019716
R48607 PAD.n4816 PAD.n4687 0.019716
R48608 PAD.n8225 PAD.n8224 0.019716
R48609 PAD.n8224 PAD.n4686 0.019716
R48610 PAD.n4822 PAD.n4821 0.019716
R48611 PAD.n4821 PAD.n4685 0.019716
R48612 PAD.n8216 PAD.n8215 0.019716
R48613 PAD.n8215 PAD.n4684 0.019716
R48614 PAD.n4827 PAD.n4826 0.019716
R48615 PAD.n4826 PAD.n4683 0.019716
R48616 PAD.n5176 PAD.n4849 0.019716
R48617 PAD.n5175 PAD.n5174 0.019716
R48618 PAD.n5174 PAD.n5173 0.019716
R48619 PAD.n5164 PAD.n4850 0.019716
R48620 PAD.n5165 PAD.n5164 0.019716
R48621 PAD.n5163 PAD.n5162 0.019716
R48622 PAD.n5162 PAD.n5161 0.019716
R48623 PAD.n5152 PAD.n4855 0.019716
R48624 PAD.n5153 PAD.n5152 0.019716
R48625 PAD.n5151 PAD.n5150 0.019716
R48626 PAD.n5150 PAD.n5149 0.019716
R48627 PAD.n5140 PAD.n4859 0.019716
R48628 PAD.n5141 PAD.n5140 0.019716
R48629 PAD.n5139 PAD.n5138 0.019716
R48630 PAD.n5138 PAD.n5137 0.019716
R48631 PAD.n5128 PAD.n4863 0.019716
R48632 PAD.n5129 PAD.n5128 0.019716
R48633 PAD.n5127 PAD.n5126 0.019716
R48634 PAD.n5126 PAD.n5125 0.019716
R48635 PAD.n5116 PAD.n4867 0.019716
R48636 PAD.n5117 PAD.n5116 0.019716
R48637 PAD.n5115 PAD.n5114 0.019716
R48638 PAD.n5114 PAD.n5113 0.019716
R48639 PAD.n5104 PAD.n4871 0.019716
R48640 PAD.n5105 PAD.n5104 0.019716
R48641 PAD.n5103 PAD.n5102 0.019716
R48642 PAD.n5102 PAD.n5101 0.019716
R48643 PAD.n5092 PAD.n4875 0.019716
R48644 PAD.n5093 PAD.n5092 0.019716
R48645 PAD.n5091 PAD.n5090 0.019716
R48646 PAD.n5090 PAD.n5089 0.019716
R48647 PAD.n5080 PAD.n4879 0.019716
R48648 PAD.n5081 PAD.n5080 0.019716
R48649 PAD.n5079 PAD.n5078 0.019716
R48650 PAD.n5078 PAD.n5077 0.019716
R48651 PAD.n5068 PAD.n4883 0.019716
R48652 PAD.n5069 PAD.n5068 0.019716
R48653 PAD.n5067 PAD.n5066 0.019716
R48654 PAD.n5066 PAD.n5065 0.019716
R48655 PAD.n5056 PAD.n4887 0.019716
R48656 PAD.n5057 PAD.n5056 0.019716
R48657 PAD.n5055 PAD.n5054 0.019716
R48658 PAD.n5054 PAD.n5053 0.019716
R48659 PAD.n5044 PAD.n4891 0.019716
R48660 PAD.n5045 PAD.n5044 0.019716
R48661 PAD.n5043 PAD.n5042 0.019716
R48662 PAD.n5042 PAD.n5041 0.019716
R48663 PAD.n5032 PAD.n4895 0.019716
R48664 PAD.n5033 PAD.n5032 0.019716
R48665 PAD.n5031 PAD.n5030 0.019716
R48666 PAD.n5030 PAD.n5029 0.019716
R48667 PAD.n5020 PAD.n4899 0.019716
R48668 PAD.n5021 PAD.n5020 0.019716
R48669 PAD.n5019 PAD.n5018 0.019716
R48670 PAD.n5018 PAD.n5017 0.019716
R48671 PAD.n5008 PAD.n4903 0.019716
R48672 PAD.n5009 PAD.n5008 0.019716
R48673 PAD.n5007 PAD.n5006 0.019716
R48674 PAD.n5006 PAD.n5005 0.019716
R48675 PAD.n4996 PAD.n4907 0.019716
R48676 PAD.n4997 PAD.n4996 0.019716
R48677 PAD.n4995 PAD.n4994 0.019716
R48678 PAD.n4994 PAD.n4993 0.019716
R48679 PAD.n4984 PAD.n4911 0.019716
R48680 PAD.n4985 PAD.n4984 0.019716
R48681 PAD.n4983 PAD.n4982 0.019716
R48682 PAD.n4982 PAD.n4981 0.019716
R48683 PAD.n4972 PAD.n4915 0.019716
R48684 PAD.n4973 PAD.n4972 0.019716
R48685 PAD.n4971 PAD.n4970 0.019716
R48686 PAD.n4970 PAD.n4969 0.019716
R48687 PAD.n4960 PAD.n4919 0.019716
R48688 PAD.n4961 PAD.n4960 0.019716
R48689 PAD.n4959 PAD.n4958 0.019716
R48690 PAD.n4958 PAD.n4957 0.019716
R48691 PAD.n4948 PAD.n4923 0.019716
R48692 PAD.n4949 PAD.n4948 0.019716
R48693 PAD.n4947 PAD.n4946 0.019716
R48694 PAD.n4946 PAD.n4945 0.019716
R48695 PAD.n4936 PAD.n4927 0.019716
R48696 PAD.n4937 PAD.n4936 0.019716
R48697 PAD.n4935 PAD.n4934 0.019716
R48698 PAD.n4934 PAD.n4933 0.019716
R48699 PAD.n8162 PAD.n7871 0.019716
R48700 PAD.n7873 PAD.n7872 0.019716
R48701 PAD.n7873 PAD.n7870 0.019716
R48702 PAD.n8153 PAD.n8152 0.019716
R48703 PAD.n8152 PAD.n7869 0.019716
R48704 PAD.n7878 PAD.n7877 0.019716
R48705 PAD.n7877 PAD.n7868 0.019716
R48706 PAD.n8144 PAD.n8143 0.019716
R48707 PAD.n8143 PAD.n7867 0.019716
R48708 PAD.n7883 PAD.n7882 0.019716
R48709 PAD.n7882 PAD.n7866 0.019716
R48710 PAD.n8135 PAD.n8134 0.019716
R48711 PAD.n8134 PAD.n7865 0.019716
R48712 PAD.n7888 PAD.n7887 0.019716
R48713 PAD.n7887 PAD.n7864 0.019716
R48714 PAD.n8126 PAD.n8125 0.019716
R48715 PAD.n8125 PAD.n7863 0.019716
R48716 PAD.n7893 PAD.n7892 0.019716
R48717 PAD.n7892 PAD.n7862 0.019716
R48718 PAD.n8117 PAD.n8116 0.019716
R48719 PAD.n8116 PAD.n7861 0.019716
R48720 PAD.n7898 PAD.n7897 0.019716
R48721 PAD.n7897 PAD.n7860 0.019716
R48722 PAD.n8108 PAD.n8107 0.019716
R48723 PAD.n8107 PAD.n7859 0.019716
R48724 PAD.n7903 PAD.n7902 0.019716
R48725 PAD.n7902 PAD.n7858 0.019716
R48726 PAD.n8099 PAD.n8098 0.019716
R48727 PAD.n8098 PAD.n7857 0.019716
R48728 PAD.n7908 PAD.n7907 0.019716
R48729 PAD.n7907 PAD.n7856 0.019716
R48730 PAD.n8090 PAD.n8089 0.019716
R48731 PAD.n8089 PAD.n7855 0.019716
R48732 PAD.n7913 PAD.n7912 0.019716
R48733 PAD.n7912 PAD.n7854 0.019716
R48734 PAD.n8081 PAD.n8080 0.019716
R48735 PAD.n8080 PAD.n7853 0.019716
R48736 PAD.n7918 PAD.n7917 0.019716
R48737 PAD.n7917 PAD.n7852 0.019716
R48738 PAD.n8072 PAD.n8071 0.019716
R48739 PAD.n8071 PAD.n7851 0.019716
R48740 PAD.n7923 PAD.n7922 0.019716
R48741 PAD.n7922 PAD.n7850 0.019716
R48742 PAD.n8063 PAD.n8062 0.019716
R48743 PAD.n8062 PAD.n7849 0.019716
R48744 PAD.n7928 PAD.n7927 0.019716
R48745 PAD.n7927 PAD.n7848 0.019716
R48746 PAD.n8054 PAD.n8053 0.019716
R48747 PAD.n8053 PAD.n7847 0.019716
R48748 PAD.n7933 PAD.n7932 0.019716
R48749 PAD.n7932 PAD.n7846 0.019716
R48750 PAD.n8045 PAD.n8044 0.019716
R48751 PAD.n8044 PAD.n7845 0.019716
R48752 PAD.n7938 PAD.n7937 0.019716
R48753 PAD.n7937 PAD.n7844 0.019716
R48754 PAD.n8036 PAD.n8035 0.019716
R48755 PAD.n8035 PAD.n7843 0.019716
R48756 PAD.n7943 PAD.n7942 0.019716
R48757 PAD.n7942 PAD.n7842 0.019716
R48758 PAD.n8027 PAD.n8026 0.019716
R48759 PAD.n8026 PAD.n7841 0.019716
R48760 PAD.n7948 PAD.n7947 0.019716
R48761 PAD.n7947 PAD.n7840 0.019716
R48762 PAD.n8018 PAD.n8017 0.019716
R48763 PAD.n8017 PAD.n7839 0.019716
R48764 PAD.n7953 PAD.n7952 0.019716
R48765 PAD.n7952 PAD.n7838 0.019716
R48766 PAD.n8009 PAD.n8008 0.019716
R48767 PAD.n8008 PAD.n7837 0.019716
R48768 PAD.n7958 PAD.n7957 0.019716
R48769 PAD.n7957 PAD.n7836 0.019716
R48770 PAD.n8000 PAD.n7999 0.019716
R48771 PAD.n7999 PAD.n7835 0.019716
R48772 PAD.n7963 PAD.n7962 0.019716
R48773 PAD.n7962 PAD.n7834 0.019716
R48774 PAD.n7991 PAD.n7990 0.019716
R48775 PAD.n7990 PAD.n7833 0.019716
R48776 PAD.n7968 PAD.n7967 0.019716
R48777 PAD.n7967 PAD.n7832 0.019716
R48778 PAD.n7982 PAD.n7981 0.019716
R48779 PAD.n7981 PAD.n7831 0.019716
R48780 PAD.n7975 PAD.n7974 0.019716
R48781 PAD.n7974 PAD.n7830 0.019716
R48782 PAD.n5540 PAD.n5213 0.019716
R48783 PAD.n5539 PAD.n5538 0.019716
R48784 PAD.n5538 PAD.n5537 0.019716
R48785 PAD.n5528 PAD.n5214 0.019716
R48786 PAD.n5529 PAD.n5528 0.019716
R48787 PAD.n5527 PAD.n5526 0.019716
R48788 PAD.n5526 PAD.n5525 0.019716
R48789 PAD.n5516 PAD.n5219 0.019716
R48790 PAD.n5517 PAD.n5516 0.019716
R48791 PAD.n5515 PAD.n5514 0.019716
R48792 PAD.n5514 PAD.n5513 0.019716
R48793 PAD.n5504 PAD.n5223 0.019716
R48794 PAD.n5505 PAD.n5504 0.019716
R48795 PAD.n5503 PAD.n5502 0.019716
R48796 PAD.n5502 PAD.n5501 0.019716
R48797 PAD.n5492 PAD.n5227 0.019716
R48798 PAD.n5493 PAD.n5492 0.019716
R48799 PAD.n5491 PAD.n5490 0.019716
R48800 PAD.n5490 PAD.n5489 0.019716
R48801 PAD.n5480 PAD.n5231 0.019716
R48802 PAD.n5481 PAD.n5480 0.019716
R48803 PAD.n5479 PAD.n5478 0.019716
R48804 PAD.n5478 PAD.n5477 0.019716
R48805 PAD.n5468 PAD.n5235 0.019716
R48806 PAD.n5469 PAD.n5468 0.019716
R48807 PAD.n5467 PAD.n5466 0.019716
R48808 PAD.n5466 PAD.n5465 0.019716
R48809 PAD.n5456 PAD.n5239 0.019716
R48810 PAD.n5457 PAD.n5456 0.019716
R48811 PAD.n5455 PAD.n5454 0.019716
R48812 PAD.n5454 PAD.n5453 0.019716
R48813 PAD.n5444 PAD.n5243 0.019716
R48814 PAD.n5445 PAD.n5444 0.019716
R48815 PAD.n5443 PAD.n5442 0.019716
R48816 PAD.n5442 PAD.n5441 0.019716
R48817 PAD.n5432 PAD.n5247 0.019716
R48818 PAD.n5433 PAD.n5432 0.019716
R48819 PAD.n5431 PAD.n5430 0.019716
R48820 PAD.n5430 PAD.n5429 0.019716
R48821 PAD.n5420 PAD.n5251 0.019716
R48822 PAD.n5421 PAD.n5420 0.019716
R48823 PAD.n5419 PAD.n5418 0.019716
R48824 PAD.n5418 PAD.n5417 0.019716
R48825 PAD.n5408 PAD.n5255 0.019716
R48826 PAD.n5409 PAD.n5408 0.019716
R48827 PAD.n5407 PAD.n5406 0.019716
R48828 PAD.n5406 PAD.n5405 0.019716
R48829 PAD.n5396 PAD.n5259 0.019716
R48830 PAD.n5397 PAD.n5396 0.019716
R48831 PAD.n5395 PAD.n5394 0.019716
R48832 PAD.n5394 PAD.n5393 0.019716
R48833 PAD.n5384 PAD.n5263 0.019716
R48834 PAD.n5385 PAD.n5384 0.019716
R48835 PAD.n5383 PAD.n5382 0.019716
R48836 PAD.n5382 PAD.n5381 0.019716
R48837 PAD.n5372 PAD.n5267 0.019716
R48838 PAD.n5373 PAD.n5372 0.019716
R48839 PAD.n5371 PAD.n5370 0.019716
R48840 PAD.n5370 PAD.n5369 0.019716
R48841 PAD.n5360 PAD.n5271 0.019716
R48842 PAD.n5361 PAD.n5360 0.019716
R48843 PAD.n5359 PAD.n5358 0.019716
R48844 PAD.n5358 PAD.n5357 0.019716
R48845 PAD.n5348 PAD.n5275 0.019716
R48846 PAD.n5349 PAD.n5348 0.019716
R48847 PAD.n5347 PAD.n5346 0.019716
R48848 PAD.n5346 PAD.n5345 0.019716
R48849 PAD.n5336 PAD.n5279 0.019716
R48850 PAD.n5337 PAD.n5336 0.019716
R48851 PAD.n5335 PAD.n5334 0.019716
R48852 PAD.n5334 PAD.n5333 0.019716
R48853 PAD.n5324 PAD.n5283 0.019716
R48854 PAD.n5325 PAD.n5324 0.019716
R48855 PAD.n5323 PAD.n5322 0.019716
R48856 PAD.n5322 PAD.n5321 0.019716
R48857 PAD.n5312 PAD.n5287 0.019716
R48858 PAD.n5313 PAD.n5312 0.019716
R48859 PAD.n5311 PAD.n5310 0.019716
R48860 PAD.n5310 PAD.n5309 0.019716
R48861 PAD.n5300 PAD.n5291 0.019716
R48862 PAD.n5301 PAD.n5300 0.019716
R48863 PAD.n5299 PAD.n5298 0.019716
R48864 PAD.n5298 PAD.n5297 0.019716
R48865 PAD.n7781 PAD.n7104 0.019716
R48866 PAD.n7774 PAD.n7773 0.019716
R48867 PAD.n7774 PAD.n7102 0.019716
R48868 PAD.n7770 PAD.n7769 0.019716
R48869 PAD.n7769 PAD.n7101 0.019716
R48870 PAD.n7763 PAD.n7762 0.019716
R48871 PAD.n7763 PAD.n7100 0.019716
R48872 PAD.n7758 PAD.n7757 0.019716
R48873 PAD.n7757 PAD.n7099 0.019716
R48874 PAD.n7751 PAD.n7750 0.019716
R48875 PAD.n7751 PAD.n7098 0.019716
R48876 PAD.n7746 PAD.n7745 0.019716
R48877 PAD.n7745 PAD.n7097 0.019716
R48878 PAD.n7739 PAD.n7738 0.019716
R48879 PAD.n7739 PAD.n7096 0.019716
R48880 PAD.n7734 PAD.n7733 0.019716
R48881 PAD.n7733 PAD.n7095 0.019716
R48882 PAD.n7727 PAD.n7726 0.019716
R48883 PAD.n7727 PAD.n7094 0.019716
R48884 PAD.n7722 PAD.n7721 0.019716
R48885 PAD.n7721 PAD.n7093 0.019716
R48886 PAD.n7715 PAD.n7714 0.019716
R48887 PAD.n7715 PAD.n7092 0.019716
R48888 PAD.n7710 PAD.n7709 0.019716
R48889 PAD.n7709 PAD.n7091 0.019716
R48890 PAD.n7703 PAD.n7702 0.019716
R48891 PAD.n7703 PAD.n7090 0.019716
R48892 PAD.n7698 PAD.n7697 0.019716
R48893 PAD.n7697 PAD.n7089 0.019716
R48894 PAD.n7691 PAD.n7690 0.019716
R48895 PAD.n7691 PAD.n7088 0.019716
R48896 PAD.n7686 PAD.n7685 0.019716
R48897 PAD.n7685 PAD.n7087 0.019716
R48898 PAD.n7679 PAD.n7678 0.019716
R48899 PAD.n7679 PAD.n7086 0.019716
R48900 PAD.n7674 PAD.n7673 0.019716
R48901 PAD.n7673 PAD.n7085 0.019716
R48902 PAD.n7667 PAD.n7666 0.019716
R48903 PAD.n7667 PAD.n7084 0.019716
R48904 PAD.n7662 PAD.n7661 0.019716
R48905 PAD.n7661 PAD.n7083 0.019716
R48906 PAD.n7655 PAD.n7654 0.019716
R48907 PAD.n7655 PAD.n7082 0.019716
R48908 PAD.n7650 PAD.n7649 0.019716
R48909 PAD.n7649 PAD.n7081 0.019716
R48910 PAD.n7643 PAD.n7642 0.019716
R48911 PAD.n7643 PAD.n7080 0.019716
R48912 PAD.n7638 PAD.n7637 0.019716
R48913 PAD.n7637 PAD.n7079 0.019716
R48914 PAD.n7631 PAD.n7630 0.019716
R48915 PAD.n7631 PAD.n7078 0.019716
R48916 PAD.n7626 PAD.n7625 0.019716
R48917 PAD.n7625 PAD.n7077 0.019716
R48918 PAD.n7619 PAD.n7618 0.019716
R48919 PAD.n7619 PAD.n7076 0.019716
R48920 PAD.n7614 PAD.n7613 0.019716
R48921 PAD.n7613 PAD.n7075 0.019716
R48922 PAD.n7607 PAD.n7606 0.019716
R48923 PAD.n7607 PAD.n7074 0.019716
R48924 PAD.n7602 PAD.n7601 0.019716
R48925 PAD.n7601 PAD.n7073 0.019716
R48926 PAD.n7595 PAD.n7594 0.019716
R48927 PAD.n7595 PAD.n7072 0.019716
R48928 PAD.n7590 PAD.n7589 0.019716
R48929 PAD.n7589 PAD.n7071 0.019716
R48930 PAD.n7583 PAD.n7582 0.019716
R48931 PAD.n7583 PAD.n7070 0.019716
R48932 PAD.n7578 PAD.n7577 0.019716
R48933 PAD.n7577 PAD.n7069 0.019716
R48934 PAD.n7571 PAD.n7570 0.019716
R48935 PAD.n7571 PAD.n7068 0.019716
R48936 PAD.n7566 PAD.n7565 0.019716
R48937 PAD.n7565 PAD.n7067 0.019716
R48938 PAD.n7559 PAD.n7558 0.019716
R48939 PAD.n7559 PAD.n7066 0.019716
R48940 PAD.n7554 PAD.n7553 0.019716
R48941 PAD.n7553 PAD.n7065 0.019716
R48942 PAD.n7547 PAD.n7546 0.019716
R48943 PAD.n7547 PAD.n7064 0.019716
R48944 PAD.n7542 PAD.n7541 0.019716
R48945 PAD.n7541 PAD.n7063 0.019716
R48946 PAD.n7535 PAD.n7534 0.019716
R48947 PAD.n7535 PAD.n7062 0.019716
R48948 PAD.n7048 PAD.n6721 0.019716
R48949 PAD.n7047 PAD.n7046 0.019716
R48950 PAD.n7046 PAD.n7045 0.019716
R48951 PAD.n7036 PAD.n6722 0.019716
R48952 PAD.n7037 PAD.n7036 0.019716
R48953 PAD.n7035 PAD.n7034 0.019716
R48954 PAD.n7034 PAD.n7033 0.019716
R48955 PAD.n7024 PAD.n6727 0.019716
R48956 PAD.n7025 PAD.n7024 0.019716
R48957 PAD.n7023 PAD.n7022 0.019716
R48958 PAD.n7022 PAD.n7021 0.019716
R48959 PAD.n7012 PAD.n6731 0.019716
R48960 PAD.n7013 PAD.n7012 0.019716
R48961 PAD.n7011 PAD.n7010 0.019716
R48962 PAD.n7010 PAD.n7009 0.019716
R48963 PAD.n7000 PAD.n6735 0.019716
R48964 PAD.n7001 PAD.n7000 0.019716
R48965 PAD.n6999 PAD.n6998 0.019716
R48966 PAD.n6998 PAD.n6997 0.019716
R48967 PAD.n6988 PAD.n6739 0.019716
R48968 PAD.n6989 PAD.n6988 0.019716
R48969 PAD.n6987 PAD.n6986 0.019716
R48970 PAD.n6986 PAD.n6985 0.019716
R48971 PAD.n6976 PAD.n6743 0.019716
R48972 PAD.n6977 PAD.n6976 0.019716
R48973 PAD.n6975 PAD.n6974 0.019716
R48974 PAD.n6974 PAD.n6973 0.019716
R48975 PAD.n6964 PAD.n6747 0.019716
R48976 PAD.n6965 PAD.n6964 0.019716
R48977 PAD.n6963 PAD.n6962 0.019716
R48978 PAD.n6962 PAD.n6961 0.019716
R48979 PAD.n6952 PAD.n6751 0.019716
R48980 PAD.n6953 PAD.n6952 0.019716
R48981 PAD.n6951 PAD.n6950 0.019716
R48982 PAD.n6950 PAD.n6949 0.019716
R48983 PAD.n6940 PAD.n6755 0.019716
R48984 PAD.n6941 PAD.n6940 0.019716
R48985 PAD.n6939 PAD.n6938 0.019716
R48986 PAD.n6938 PAD.n6937 0.019716
R48987 PAD.n6928 PAD.n6759 0.019716
R48988 PAD.n6929 PAD.n6928 0.019716
R48989 PAD.n6927 PAD.n6926 0.019716
R48990 PAD.n6926 PAD.n6925 0.019716
R48991 PAD.n6916 PAD.n6763 0.019716
R48992 PAD.n6917 PAD.n6916 0.019716
R48993 PAD.n6915 PAD.n6914 0.019716
R48994 PAD.n6914 PAD.n6913 0.019716
R48995 PAD.n6904 PAD.n6767 0.019716
R48996 PAD.n6905 PAD.n6904 0.019716
R48997 PAD.n6903 PAD.n6902 0.019716
R48998 PAD.n6902 PAD.n6901 0.019716
R48999 PAD.n6892 PAD.n6771 0.019716
R49000 PAD.n6893 PAD.n6892 0.019716
R49001 PAD.n6891 PAD.n6890 0.019716
R49002 PAD.n6890 PAD.n6889 0.019716
R49003 PAD.n6880 PAD.n6775 0.019716
R49004 PAD.n6881 PAD.n6880 0.019716
R49005 PAD.n6879 PAD.n6878 0.019716
R49006 PAD.n6878 PAD.n6877 0.019716
R49007 PAD.n6868 PAD.n6779 0.019716
R49008 PAD.n6869 PAD.n6868 0.019716
R49009 PAD.n6867 PAD.n6866 0.019716
R49010 PAD.n6866 PAD.n6865 0.019716
R49011 PAD.n6856 PAD.n6783 0.019716
R49012 PAD.n6857 PAD.n6856 0.019716
R49013 PAD.n6855 PAD.n6854 0.019716
R49014 PAD.n6854 PAD.n6853 0.019716
R49015 PAD.n6844 PAD.n6787 0.019716
R49016 PAD.n6845 PAD.n6844 0.019716
R49017 PAD.n6843 PAD.n6842 0.019716
R49018 PAD.n6842 PAD.n6841 0.019716
R49019 PAD.n6832 PAD.n6791 0.019716
R49020 PAD.n6833 PAD.n6832 0.019716
R49021 PAD.n6831 PAD.n6830 0.019716
R49022 PAD.n6830 PAD.n6829 0.019716
R49023 PAD.n6820 PAD.n6795 0.019716
R49024 PAD.n6821 PAD.n6820 0.019716
R49025 PAD.n6819 PAD.n6818 0.019716
R49026 PAD.n6818 PAD.n6817 0.019716
R49027 PAD.n6808 PAD.n6799 0.019716
R49028 PAD.n6809 PAD.n6808 0.019716
R49029 PAD.n6807 PAD.n6806 0.019716
R49030 PAD.n6806 PAD.n6805 0.019716
R49031 PAD.n5893 PAD.n5602 0.019716
R49032 PAD.n5604 PAD.n5603 0.019716
R49033 PAD.n5604 PAD.n5601 0.019716
R49034 PAD.n5884 PAD.n5883 0.019716
R49035 PAD.n5883 PAD.n5600 0.019716
R49036 PAD.n5609 PAD.n5608 0.019716
R49037 PAD.n5608 PAD.n5599 0.019716
R49038 PAD.n5875 PAD.n5874 0.019716
R49039 PAD.n5874 PAD.n5598 0.019716
R49040 PAD.n5614 PAD.n5613 0.019716
R49041 PAD.n5613 PAD.n5597 0.019716
R49042 PAD.n5866 PAD.n5865 0.019716
R49043 PAD.n5865 PAD.n5596 0.019716
R49044 PAD.n5619 PAD.n5618 0.019716
R49045 PAD.n5618 PAD.n5595 0.019716
R49046 PAD.n5857 PAD.n5856 0.019716
R49047 PAD.n5856 PAD.n5594 0.019716
R49048 PAD.n5624 PAD.n5623 0.019716
R49049 PAD.n5623 PAD.n5593 0.019716
R49050 PAD.n5848 PAD.n5847 0.019716
R49051 PAD.n5847 PAD.n5592 0.019716
R49052 PAD.n5629 PAD.n5628 0.019716
R49053 PAD.n5628 PAD.n5591 0.019716
R49054 PAD.n5839 PAD.n5838 0.019716
R49055 PAD.n5838 PAD.n5590 0.019716
R49056 PAD.n5634 PAD.n5633 0.019716
R49057 PAD.n5633 PAD.n5589 0.019716
R49058 PAD.n5830 PAD.n5829 0.019716
R49059 PAD.n5829 PAD.n5588 0.019716
R49060 PAD.n5639 PAD.n5638 0.019716
R49061 PAD.n5638 PAD.n5587 0.019716
R49062 PAD.n5821 PAD.n5820 0.019716
R49063 PAD.n5820 PAD.n5586 0.019716
R49064 PAD.n5644 PAD.n5643 0.019716
R49065 PAD.n5643 PAD.n5585 0.019716
R49066 PAD.n5812 PAD.n5811 0.019716
R49067 PAD.n5811 PAD.n5584 0.019716
R49068 PAD.n5649 PAD.n5648 0.019716
R49069 PAD.n5648 PAD.n5583 0.019716
R49070 PAD.n5803 PAD.n5802 0.019716
R49071 PAD.n5802 PAD.n5582 0.019716
R49072 PAD.n5654 PAD.n5653 0.019716
R49073 PAD.n5653 PAD.n5581 0.019716
R49074 PAD.n5794 PAD.n5793 0.019716
R49075 PAD.n5793 PAD.n5580 0.019716
R49076 PAD.n5659 PAD.n5658 0.019716
R49077 PAD.n5658 PAD.n5579 0.019716
R49078 PAD.n5785 PAD.n5784 0.019716
R49079 PAD.n5784 PAD.n5578 0.019716
R49080 PAD.n5664 PAD.n5663 0.019716
R49081 PAD.n5663 PAD.n5577 0.019716
R49082 PAD.n5776 PAD.n5775 0.019716
R49083 PAD.n5775 PAD.n5576 0.019716
R49084 PAD.n5669 PAD.n5668 0.019716
R49085 PAD.n5668 PAD.n5575 0.019716
R49086 PAD.n5767 PAD.n5766 0.019716
R49087 PAD.n5766 PAD.n5574 0.019716
R49088 PAD.n5674 PAD.n5673 0.019716
R49089 PAD.n5673 PAD.n5573 0.019716
R49090 PAD.n5758 PAD.n5757 0.019716
R49091 PAD.n5757 PAD.n5572 0.019716
R49092 PAD.n5679 PAD.n5678 0.019716
R49093 PAD.n5678 PAD.n5571 0.019716
R49094 PAD.n5749 PAD.n5748 0.019716
R49095 PAD.n5748 PAD.n5570 0.019716
R49096 PAD.n5684 PAD.n5683 0.019716
R49097 PAD.n5683 PAD.n5569 0.019716
R49098 PAD.n5740 PAD.n5739 0.019716
R49099 PAD.n5739 PAD.n5568 0.019716
R49100 PAD.n5689 PAD.n5688 0.019716
R49101 PAD.n5688 PAD.n5567 0.019716
R49102 PAD.n5731 PAD.n5730 0.019716
R49103 PAD.n5730 PAD.n5566 0.019716
R49104 PAD.n5694 PAD.n5693 0.019716
R49105 PAD.n5693 PAD.n5565 0.019716
R49106 PAD.n5722 PAD.n5721 0.019716
R49107 PAD.n5721 PAD.n5564 0.019716
R49108 PAD.n5699 PAD.n5698 0.019716
R49109 PAD.n5698 PAD.n5563 0.019716
R49110 PAD.n5713 PAD.n5712 0.019716
R49111 PAD.n5712 PAD.n5562 0.019716
R49112 PAD.n5706 PAD.n5705 0.019716
R49113 PAD.n5705 PAD.n5561 0.019716
R49114 PAD.n11084 PAD.n11083 0.019716
R49115 PAD.n11083 PAD.n11082 0.019716
R49116 PAD.n11073 PAD.n10756 0.019716
R49117 PAD.n11074 PAD.n11073 0.019716
R49118 PAD.n11072 PAD.n11071 0.019716
R49119 PAD.n11071 PAD.n11070 0.019716
R49120 PAD.n11061 PAD.n10760 0.019716
R49121 PAD.n11062 PAD.n11061 0.019716
R49122 PAD.n11060 PAD.n11059 0.019716
R49123 PAD.n11059 PAD.n11058 0.019716
R49124 PAD.n11049 PAD.n10764 0.019716
R49125 PAD.n11050 PAD.n11049 0.019716
R49126 PAD.n11048 PAD.n11047 0.019716
R49127 PAD.n11047 PAD.n11046 0.019716
R49128 PAD.n11037 PAD.n10768 0.019716
R49129 PAD.n11038 PAD.n11037 0.019716
R49130 PAD.n11036 PAD.n11035 0.019716
R49131 PAD.n11035 PAD.n11034 0.019716
R49132 PAD.n11025 PAD.n10772 0.019716
R49133 PAD.n11026 PAD.n11025 0.019716
R49134 PAD.n11024 PAD.n11023 0.019716
R49135 PAD.n11023 PAD.n11022 0.019716
R49136 PAD.n11013 PAD.n10776 0.019716
R49137 PAD.n11014 PAD.n11013 0.019716
R49138 PAD.n11012 PAD.n11011 0.019716
R49139 PAD.n11011 PAD.n11010 0.019716
R49140 PAD.n11001 PAD.n10780 0.019716
R49141 PAD.n11002 PAD.n11001 0.019716
R49142 PAD.n11000 PAD.n10999 0.019716
R49143 PAD.n10999 PAD.n10998 0.019716
R49144 PAD.n10989 PAD.n10784 0.019716
R49145 PAD.n10990 PAD.n10989 0.019716
R49146 PAD.n10988 PAD.n10987 0.019716
R49147 PAD.n10987 PAD.n10986 0.019716
R49148 PAD.n10977 PAD.n10788 0.019716
R49149 PAD.n10978 PAD.n10977 0.019716
R49150 PAD.n10976 PAD.n10975 0.019716
R49151 PAD.n10975 PAD.n10974 0.019716
R49152 PAD.n10965 PAD.n10792 0.019716
R49153 PAD.n10966 PAD.n10965 0.019716
R49154 PAD.n10964 PAD.n10963 0.019716
R49155 PAD.n10963 PAD.n10962 0.019716
R49156 PAD.n10953 PAD.n10796 0.019716
R49157 PAD.n10954 PAD.n10953 0.019716
R49158 PAD.n10952 PAD.n10951 0.019716
R49159 PAD.n10951 PAD.n10950 0.019716
R49160 PAD.n10941 PAD.n10800 0.019716
R49161 PAD.n10942 PAD.n10941 0.019716
R49162 PAD.n10940 PAD.n10939 0.019716
R49163 PAD.n10939 PAD.n10938 0.019716
R49164 PAD.n10929 PAD.n10804 0.019716
R49165 PAD.n10930 PAD.n10929 0.019716
R49166 PAD.n10928 PAD.n10927 0.019716
R49167 PAD.n10927 PAD.n10926 0.019716
R49168 PAD.n10917 PAD.n10808 0.019716
R49169 PAD.n10918 PAD.n10917 0.019716
R49170 PAD.n10916 PAD.n10915 0.019716
R49171 PAD.n10915 PAD.n10914 0.019716
R49172 PAD.n10905 PAD.n10812 0.019716
R49173 PAD.n10906 PAD.n10905 0.019716
R49174 PAD.n10904 PAD.n10903 0.019716
R49175 PAD.n10903 PAD.n10902 0.019716
R49176 PAD.n10893 PAD.n10816 0.019716
R49177 PAD.n10894 PAD.n10893 0.019716
R49178 PAD.n10892 PAD.n10891 0.019716
R49179 PAD.n10891 PAD.n10890 0.019716
R49180 PAD.n10881 PAD.n10820 0.019716
R49181 PAD.n10882 PAD.n10881 0.019716
R49182 PAD.n10880 PAD.n10879 0.019716
R49183 PAD.n10879 PAD.n10878 0.019716
R49184 PAD.n10869 PAD.n10824 0.019716
R49185 PAD.n10870 PAD.n10869 0.019716
R49186 PAD.n10868 PAD.n10867 0.019716
R49187 PAD.n10867 PAD.n10866 0.019716
R49188 PAD.n10857 PAD.n10828 0.019716
R49189 PAD.n10858 PAD.n10857 0.019716
R49190 PAD.n10856 PAD.n10855 0.019716
R49191 PAD.n10855 PAD.n10854 0.019716
R49192 PAD.n10845 PAD.n10832 0.019716
R49193 PAD.n10846 PAD.n10845 0.019716
R49194 PAD.n10844 PAD.n10843 0.019716
R49195 PAD.n10843 PAD.n10842 0.019716
R49196 PAD.n10837 PAD.n10836 0.019716
R49197 PAD.n5905 PAD.n5902 0.019716
R49198 PAD.n5906 PAD.n5905 0.019716
R49199 PAD.n6495 PAD.n6397 0.019716
R49200 PAD.n6495 PAD.n5907 0.019716
R49201 PAD.n6504 PAD.n6398 0.019716
R49202 PAD.n6504 PAD.n5908 0.019716
R49203 PAD.n6492 PAD.n6399 0.019716
R49204 PAD.n6492 PAD.n5909 0.019716
R49205 PAD.n6513 PAD.n6400 0.019716
R49206 PAD.n6513 PAD.n5910 0.019716
R49207 PAD.n6489 PAD.n6401 0.019716
R49208 PAD.n6489 PAD.n5911 0.019716
R49209 PAD.n6522 PAD.n6402 0.019716
R49210 PAD.n6522 PAD.n5912 0.019716
R49211 PAD.n6486 PAD.n6403 0.019716
R49212 PAD.n6486 PAD.n5913 0.019716
R49213 PAD.n6531 PAD.n6404 0.019716
R49214 PAD.n6531 PAD.n5914 0.019716
R49215 PAD.n6483 PAD.n6405 0.019716
R49216 PAD.n6483 PAD.n5915 0.019716
R49217 PAD.n6540 PAD.n6406 0.019716
R49218 PAD.n6540 PAD.n5916 0.019716
R49219 PAD.n6480 PAD.n6407 0.019716
R49220 PAD.n6480 PAD.n5917 0.019716
R49221 PAD.n6549 PAD.n6408 0.019716
R49222 PAD.n6549 PAD.n5918 0.019716
R49223 PAD.n6477 PAD.n6409 0.019716
R49224 PAD.n6477 PAD.n5919 0.019716
R49225 PAD.n6558 PAD.n6410 0.019716
R49226 PAD.n6558 PAD.n5920 0.019716
R49227 PAD.n6474 PAD.n6411 0.019716
R49228 PAD.n6474 PAD.n5921 0.019716
R49229 PAD.n6567 PAD.n6412 0.019716
R49230 PAD.n6567 PAD.n5922 0.019716
R49231 PAD.n6471 PAD.n6413 0.019716
R49232 PAD.n6471 PAD.n5923 0.019716
R49233 PAD.n6576 PAD.n6414 0.019716
R49234 PAD.n6576 PAD.n5924 0.019716
R49235 PAD.n6468 PAD.n6415 0.019716
R49236 PAD.n6468 PAD.n5925 0.019716
R49237 PAD.n6585 PAD.n6416 0.019716
R49238 PAD.n6585 PAD.n5926 0.019716
R49239 PAD.n6465 PAD.n6417 0.019716
R49240 PAD.n6465 PAD.n5927 0.019716
R49241 PAD.n6594 PAD.n6418 0.019716
R49242 PAD.n6594 PAD.n5928 0.019716
R49243 PAD.n6462 PAD.n6419 0.019716
R49244 PAD.n6462 PAD.n5929 0.019716
R49245 PAD.n6603 PAD.n6420 0.019716
R49246 PAD.n6603 PAD.n5930 0.019716
R49247 PAD.n6459 PAD.n6421 0.019716
R49248 PAD.n6459 PAD.n5931 0.019716
R49249 PAD.n6612 PAD.n6422 0.019716
R49250 PAD.n6612 PAD.n5932 0.019716
R49251 PAD.n6456 PAD.n6423 0.019716
R49252 PAD.n6456 PAD.n5933 0.019716
R49253 PAD.n6621 PAD.n6424 0.019716
R49254 PAD.n6621 PAD.n5934 0.019716
R49255 PAD.n6453 PAD.n6425 0.019716
R49256 PAD.n6453 PAD.n5935 0.019716
R49257 PAD.n6630 PAD.n6426 0.019716
R49258 PAD.n6630 PAD.n5936 0.019716
R49259 PAD.n6450 PAD.n6427 0.019716
R49260 PAD.n6450 PAD.n5937 0.019716
R49261 PAD.n6639 PAD.n6428 0.019716
R49262 PAD.n6639 PAD.n5938 0.019716
R49263 PAD.n6447 PAD.n6429 0.019716
R49264 PAD.n6447 PAD.n5939 0.019716
R49265 PAD.n6648 PAD.n6430 0.019716
R49266 PAD.n6648 PAD.n5940 0.019716
R49267 PAD.n6444 PAD.n6431 0.019716
R49268 PAD.n6444 PAD.n5941 0.019716
R49269 PAD.n6657 PAD.n6432 0.019716
R49270 PAD.n6657 PAD.n5942 0.019716
R49271 PAD.n6441 PAD.n6433 0.019716
R49272 PAD.n6441 PAD.n5943 0.019716
R49273 PAD.n6666 PAD.n6434 0.019716
R49274 PAD.n6666 PAD.n5944 0.019716
R49275 PAD.n6437 PAD.n6435 0.019716
R49276 PAD.n6437 PAD.n5945 0.019716
R49277 PAD.n6677 PAD.n6436 0.019716
R49278 PAD.n6436 PAD.n5946 0.019716
R49279 PAD.n6688 PAD.n5947 0.019716
R49280 PAD.n11085 PAD.n11084 0.019716
R49281 PAD.n11081 PAD.n10756 0.019716
R49282 PAD.n11082 PAD.n11081 0.019716
R49283 PAD.n11075 PAD.n11072 0.019716
R49284 PAD.n11075 PAD.n11074 0.019716
R49285 PAD.n11069 PAD.n10760 0.019716
R49286 PAD.n11070 PAD.n11069 0.019716
R49287 PAD.n11063 PAD.n11060 0.019716
R49288 PAD.n11063 PAD.n11062 0.019716
R49289 PAD.n11057 PAD.n10764 0.019716
R49290 PAD.n11058 PAD.n11057 0.019716
R49291 PAD.n11051 PAD.n11048 0.019716
R49292 PAD.n11051 PAD.n11050 0.019716
R49293 PAD.n11045 PAD.n10768 0.019716
R49294 PAD.n11046 PAD.n11045 0.019716
R49295 PAD.n11039 PAD.n11036 0.019716
R49296 PAD.n11039 PAD.n11038 0.019716
R49297 PAD.n11033 PAD.n10772 0.019716
R49298 PAD.n11034 PAD.n11033 0.019716
R49299 PAD.n11027 PAD.n11024 0.019716
R49300 PAD.n11027 PAD.n11026 0.019716
R49301 PAD.n11021 PAD.n10776 0.019716
R49302 PAD.n11022 PAD.n11021 0.019716
R49303 PAD.n11015 PAD.n11012 0.019716
R49304 PAD.n11015 PAD.n11014 0.019716
R49305 PAD.n11009 PAD.n10780 0.019716
R49306 PAD.n11010 PAD.n11009 0.019716
R49307 PAD.n11003 PAD.n11000 0.019716
R49308 PAD.n11003 PAD.n11002 0.019716
R49309 PAD.n10997 PAD.n10784 0.019716
R49310 PAD.n10998 PAD.n10997 0.019716
R49311 PAD.n10991 PAD.n10988 0.019716
R49312 PAD.n10991 PAD.n10990 0.019716
R49313 PAD.n10985 PAD.n10788 0.019716
R49314 PAD.n10986 PAD.n10985 0.019716
R49315 PAD.n10979 PAD.n10976 0.019716
R49316 PAD.n10979 PAD.n10978 0.019716
R49317 PAD.n10973 PAD.n10792 0.019716
R49318 PAD.n10974 PAD.n10973 0.019716
R49319 PAD.n10967 PAD.n10964 0.019716
R49320 PAD.n10967 PAD.n10966 0.019716
R49321 PAD.n10961 PAD.n10796 0.019716
R49322 PAD.n10962 PAD.n10961 0.019716
R49323 PAD.n10955 PAD.n10952 0.019716
R49324 PAD.n10955 PAD.n10954 0.019716
R49325 PAD.n10949 PAD.n10800 0.019716
R49326 PAD.n10950 PAD.n10949 0.019716
R49327 PAD.n10943 PAD.n10940 0.019716
R49328 PAD.n10943 PAD.n10942 0.019716
R49329 PAD.n10937 PAD.n10804 0.019716
R49330 PAD.n10938 PAD.n10937 0.019716
R49331 PAD.n10931 PAD.n10928 0.019716
R49332 PAD.n10931 PAD.n10930 0.019716
R49333 PAD.n10925 PAD.n10808 0.019716
R49334 PAD.n10926 PAD.n10925 0.019716
R49335 PAD.n10919 PAD.n10916 0.019716
R49336 PAD.n10919 PAD.n10918 0.019716
R49337 PAD.n10913 PAD.n10812 0.019716
R49338 PAD.n10914 PAD.n10913 0.019716
R49339 PAD.n10907 PAD.n10904 0.019716
R49340 PAD.n10907 PAD.n10906 0.019716
R49341 PAD.n10901 PAD.n10816 0.019716
R49342 PAD.n10902 PAD.n10901 0.019716
R49343 PAD.n10895 PAD.n10892 0.019716
R49344 PAD.n10895 PAD.n10894 0.019716
R49345 PAD.n10889 PAD.n10820 0.019716
R49346 PAD.n10890 PAD.n10889 0.019716
R49347 PAD.n10883 PAD.n10880 0.019716
R49348 PAD.n10883 PAD.n10882 0.019716
R49349 PAD.n10877 PAD.n10824 0.019716
R49350 PAD.n10878 PAD.n10877 0.019716
R49351 PAD.n10871 PAD.n10868 0.019716
R49352 PAD.n10871 PAD.n10870 0.019716
R49353 PAD.n10865 PAD.n10828 0.019716
R49354 PAD.n10866 PAD.n10865 0.019716
R49355 PAD.n10859 PAD.n10856 0.019716
R49356 PAD.n10859 PAD.n10858 0.019716
R49357 PAD.n10853 PAD.n10832 0.019716
R49358 PAD.n10854 PAD.n10853 0.019716
R49359 PAD.n10847 PAD.n10844 0.019716
R49360 PAD.n10847 PAD.n10846 0.019716
R49361 PAD.n10841 PAD.n10836 0.019716
R49362 PAD.n10842 PAD.n10841 0.019716
R49363 PAD.n116 PAD.n74 0.019716
R49364 PAD.n117 PAD.n73 0.019716
R49365 PAD.n126 PAD.n72 0.019716
R49366 PAD.n126 PAD.n125 0.019716
R49367 PAD.n128 PAD.n71 0.019716
R49368 PAD.n129 PAD.n128 0.019716
R49369 PAD.n138 PAD.n70 0.019716
R49370 PAD.n138 PAD.n137 0.019716
R49371 PAD.n140 PAD.n69 0.019716
R49372 PAD.n141 PAD.n140 0.019716
R49373 PAD.n150 PAD.n68 0.019716
R49374 PAD.n150 PAD.n149 0.019716
R49375 PAD.n152 PAD.n67 0.019716
R49376 PAD.n153 PAD.n152 0.019716
R49377 PAD.n162 PAD.n66 0.019716
R49378 PAD.n162 PAD.n161 0.019716
R49379 PAD.n164 PAD.n65 0.019716
R49380 PAD.n165 PAD.n164 0.019716
R49381 PAD.n174 PAD.n64 0.019716
R49382 PAD.n174 PAD.n173 0.019716
R49383 PAD.n176 PAD.n63 0.019716
R49384 PAD.n177 PAD.n176 0.019716
R49385 PAD.n186 PAD.n62 0.019716
R49386 PAD.n186 PAD.n185 0.019716
R49387 PAD.n188 PAD.n61 0.019716
R49388 PAD.n189 PAD.n188 0.019716
R49389 PAD.n198 PAD.n60 0.019716
R49390 PAD.n198 PAD.n197 0.019716
R49391 PAD.n200 PAD.n59 0.019716
R49392 PAD.n201 PAD.n200 0.019716
R49393 PAD.n210 PAD.n58 0.019716
R49394 PAD.n210 PAD.n209 0.019716
R49395 PAD.n212 PAD.n57 0.019716
R49396 PAD.n213 PAD.n212 0.019716
R49397 PAD.n222 PAD.n56 0.019716
R49398 PAD.n222 PAD.n221 0.019716
R49399 PAD.n224 PAD.n55 0.019716
R49400 PAD.n225 PAD.n224 0.019716
R49401 PAD.n234 PAD.n54 0.019716
R49402 PAD.n234 PAD.n233 0.019716
R49403 PAD.n236 PAD.n53 0.019716
R49404 PAD.n237 PAD.n236 0.019716
R49405 PAD.n246 PAD.n52 0.019716
R49406 PAD.n246 PAD.n245 0.019716
R49407 PAD.n248 PAD.n51 0.019716
R49408 PAD.n249 PAD.n248 0.019716
R49409 PAD.n258 PAD.n50 0.019716
R49410 PAD.n258 PAD.n257 0.019716
R49411 PAD.n260 PAD.n49 0.019716
R49412 PAD.n261 PAD.n260 0.019716
R49413 PAD.n270 PAD.n48 0.019716
R49414 PAD.n270 PAD.n269 0.019716
R49415 PAD.n272 PAD.n47 0.019716
R49416 PAD.n273 PAD.n272 0.019716
R49417 PAD.n282 PAD.n46 0.019716
R49418 PAD.n282 PAD.n281 0.019716
R49419 PAD.n284 PAD.n45 0.019716
R49420 PAD.n285 PAD.n284 0.019716
R49421 PAD.n294 PAD.n44 0.019716
R49422 PAD.n294 PAD.n293 0.019716
R49423 PAD.n296 PAD.n43 0.019716
R49424 PAD.n297 PAD.n296 0.019716
R49425 PAD.n306 PAD.n42 0.019716
R49426 PAD.n306 PAD.n305 0.019716
R49427 PAD.n308 PAD.n41 0.019716
R49428 PAD.n309 PAD.n308 0.019716
R49429 PAD.n318 PAD.n40 0.019716
R49430 PAD.n318 PAD.n317 0.019716
R49431 PAD.n320 PAD.n39 0.019716
R49432 PAD.n321 PAD.n320 0.019716
R49433 PAD.n330 PAD.n38 0.019716
R49434 PAD.n330 PAD.n329 0.019716
R49435 PAD.n332 PAD.n37 0.019716
R49436 PAD.n333 PAD.n332 0.019716
R49437 PAD.n342 PAD.n36 0.019716
R49438 PAD.n342 PAD.n341 0.019716
R49439 PAD.n344 PAD.n35 0.019716
R49440 PAD.n345 PAD.n344 0.019716
R49441 PAD.n354 PAD.n34 0.019716
R49442 PAD.n354 PAD.n353 0.019716
R49443 PAD.n356 PAD.n33 0.019716
R49444 PAD.n357 PAD.n356 0.019716
R49445 PAD.n366 PAD.n365 0.019716
R49446 PAD.n10692 PAD.n415 0.019716
R49447 PAD.n10693 PAD.n414 0.019716
R49448 PAD.n10415 PAD.n413 0.019716
R49449 PAD.n10416 PAD.n10415 0.019716
R49450 PAD.n10684 PAD.n412 0.019716
R49451 PAD.n10685 PAD.n10684 0.019716
R49452 PAD.n10420 PAD.n411 0.019716
R49453 PAD.n10421 PAD.n10420 0.019716
R49454 PAD.n10675 PAD.n410 0.019716
R49455 PAD.n10676 PAD.n10675 0.019716
R49456 PAD.n10425 PAD.n409 0.019716
R49457 PAD.n10426 PAD.n10425 0.019716
R49458 PAD.n10666 PAD.n408 0.019716
R49459 PAD.n10667 PAD.n10666 0.019716
R49460 PAD.n10430 PAD.n407 0.019716
R49461 PAD.n10431 PAD.n10430 0.019716
R49462 PAD.n10657 PAD.n406 0.019716
R49463 PAD.n10658 PAD.n10657 0.019716
R49464 PAD.n10435 PAD.n405 0.019716
R49465 PAD.n10436 PAD.n10435 0.019716
R49466 PAD.n10648 PAD.n404 0.019716
R49467 PAD.n10649 PAD.n10648 0.019716
R49468 PAD.n10440 PAD.n403 0.019716
R49469 PAD.n10441 PAD.n10440 0.019716
R49470 PAD.n10639 PAD.n402 0.019716
R49471 PAD.n10640 PAD.n10639 0.019716
R49472 PAD.n10445 PAD.n401 0.019716
R49473 PAD.n10446 PAD.n10445 0.019716
R49474 PAD.n10630 PAD.n400 0.019716
R49475 PAD.n10631 PAD.n10630 0.019716
R49476 PAD.n10450 PAD.n399 0.019716
R49477 PAD.n10451 PAD.n10450 0.019716
R49478 PAD.n10621 PAD.n398 0.019716
R49479 PAD.n10622 PAD.n10621 0.019716
R49480 PAD.n10455 PAD.n397 0.019716
R49481 PAD.n10456 PAD.n10455 0.019716
R49482 PAD.n10612 PAD.n396 0.019716
R49483 PAD.n10613 PAD.n10612 0.019716
R49484 PAD.n10460 PAD.n395 0.019716
R49485 PAD.n10461 PAD.n10460 0.019716
R49486 PAD.n10603 PAD.n394 0.019716
R49487 PAD.n10604 PAD.n10603 0.019716
R49488 PAD.n10465 PAD.n393 0.019716
R49489 PAD.n10466 PAD.n10465 0.019716
R49490 PAD.n10594 PAD.n392 0.019716
R49491 PAD.n10595 PAD.n10594 0.019716
R49492 PAD.n10470 PAD.n391 0.019716
R49493 PAD.n10471 PAD.n10470 0.019716
R49494 PAD.n10585 PAD.n390 0.019716
R49495 PAD.n10586 PAD.n10585 0.019716
R49496 PAD.n10475 PAD.n389 0.019716
R49497 PAD.n10476 PAD.n10475 0.019716
R49498 PAD.n10576 PAD.n388 0.019716
R49499 PAD.n10577 PAD.n10576 0.019716
R49500 PAD.n10480 PAD.n387 0.019716
R49501 PAD.n10481 PAD.n10480 0.019716
R49502 PAD.n10567 PAD.n386 0.019716
R49503 PAD.n10568 PAD.n10567 0.019716
R49504 PAD.n10485 PAD.n385 0.019716
R49505 PAD.n10486 PAD.n10485 0.019716
R49506 PAD.n10558 PAD.n384 0.019716
R49507 PAD.n10559 PAD.n10558 0.019716
R49508 PAD.n10490 PAD.n383 0.019716
R49509 PAD.n10491 PAD.n10490 0.019716
R49510 PAD.n10549 PAD.n382 0.019716
R49511 PAD.n10550 PAD.n10549 0.019716
R49512 PAD.n10495 PAD.n381 0.019716
R49513 PAD.n10496 PAD.n10495 0.019716
R49514 PAD.n10540 PAD.n380 0.019716
R49515 PAD.n10541 PAD.n10540 0.019716
R49516 PAD.n10500 PAD.n379 0.019716
R49517 PAD.n10501 PAD.n10500 0.019716
R49518 PAD.n10531 PAD.n378 0.019716
R49519 PAD.n10532 PAD.n10531 0.019716
R49520 PAD.n10505 PAD.n377 0.019716
R49521 PAD.n10506 PAD.n10505 0.019716
R49522 PAD.n10522 PAD.n376 0.019716
R49523 PAD.n10523 PAD.n10522 0.019716
R49524 PAD.n10510 PAD.n375 0.019716
R49525 PAD.n10511 PAD.n10510 0.019716
R49526 PAD.n10513 PAD.n374 0.019716
R49527 PAD.n10514 PAD.n10513 0.019716
R49528 PAD.n10715 PAD.n10714 0.019716
R49529 PAD.n524 PAD.n523 0.019716
R49530 PAD.n526 PAD.n525 0.019716
R49531 PAD.n527 PAD.n517 0.019716
R49532 PAD.n528 PAD.n527 0.019716
R49533 PAD.n538 PAD.n537 0.019716
R49534 PAD.n537 PAD.n536 0.019716
R49535 PAD.n539 PAD.n513 0.019716
R49536 PAD.n540 PAD.n539 0.019716
R49537 PAD.n550 PAD.n549 0.019716
R49538 PAD.n549 PAD.n548 0.019716
R49539 PAD.n551 PAD.n509 0.019716
R49540 PAD.n552 PAD.n551 0.019716
R49541 PAD.n562 PAD.n561 0.019716
R49542 PAD.n561 PAD.n560 0.019716
R49543 PAD.n563 PAD.n505 0.019716
R49544 PAD.n564 PAD.n563 0.019716
R49545 PAD.n574 PAD.n573 0.019716
R49546 PAD.n573 PAD.n572 0.019716
R49547 PAD.n575 PAD.n501 0.019716
R49548 PAD.n576 PAD.n575 0.019716
R49549 PAD.n586 PAD.n585 0.019716
R49550 PAD.n585 PAD.n584 0.019716
R49551 PAD.n587 PAD.n497 0.019716
R49552 PAD.n588 PAD.n587 0.019716
R49553 PAD.n598 PAD.n597 0.019716
R49554 PAD.n597 PAD.n596 0.019716
R49555 PAD.n599 PAD.n493 0.019716
R49556 PAD.n600 PAD.n599 0.019716
R49557 PAD.n610 PAD.n609 0.019716
R49558 PAD.n609 PAD.n608 0.019716
R49559 PAD.n611 PAD.n489 0.019716
R49560 PAD.n612 PAD.n611 0.019716
R49561 PAD.n622 PAD.n621 0.019716
R49562 PAD.n621 PAD.n620 0.019716
R49563 PAD.n623 PAD.n485 0.019716
R49564 PAD.n624 PAD.n623 0.019716
R49565 PAD.n634 PAD.n633 0.019716
R49566 PAD.n633 PAD.n632 0.019716
R49567 PAD.n635 PAD.n481 0.019716
R49568 PAD.n636 PAD.n635 0.019716
R49569 PAD.n646 PAD.n645 0.019716
R49570 PAD.n645 PAD.n644 0.019716
R49571 PAD.n647 PAD.n477 0.019716
R49572 PAD.n648 PAD.n647 0.019716
R49573 PAD.n658 PAD.n657 0.019716
R49574 PAD.n657 PAD.n656 0.019716
R49575 PAD.n659 PAD.n473 0.019716
R49576 PAD.n660 PAD.n659 0.019716
R49577 PAD.n670 PAD.n669 0.019716
R49578 PAD.n669 PAD.n668 0.019716
R49579 PAD.n671 PAD.n469 0.019716
R49580 PAD.n672 PAD.n671 0.019716
R49581 PAD.n682 PAD.n681 0.019716
R49582 PAD.n681 PAD.n680 0.019716
R49583 PAD.n683 PAD.n465 0.019716
R49584 PAD.n684 PAD.n683 0.019716
R49585 PAD.n694 PAD.n693 0.019716
R49586 PAD.n693 PAD.n692 0.019716
R49587 PAD.n695 PAD.n461 0.019716
R49588 PAD.n696 PAD.n695 0.019716
R49589 PAD.n706 PAD.n705 0.019716
R49590 PAD.n705 PAD.n704 0.019716
R49591 PAD.n707 PAD.n457 0.019716
R49592 PAD.n708 PAD.n707 0.019716
R49593 PAD.n718 PAD.n717 0.019716
R49594 PAD.n717 PAD.n716 0.019716
R49595 PAD.n719 PAD.n453 0.019716
R49596 PAD.n720 PAD.n719 0.019716
R49597 PAD.n730 PAD.n729 0.019716
R49598 PAD.n729 PAD.n728 0.019716
R49599 PAD.n731 PAD.n449 0.019716
R49600 PAD.n732 PAD.n731 0.019716
R49601 PAD.n742 PAD.n741 0.019716
R49602 PAD.n741 PAD.n740 0.019716
R49603 PAD.n743 PAD.n445 0.019716
R49604 PAD.n744 PAD.n743 0.019716
R49605 PAD.n754 PAD.n753 0.019716
R49606 PAD.n753 PAD.n752 0.019716
R49607 PAD.n755 PAD.n441 0.019716
R49608 PAD.n756 PAD.n755 0.019716
R49609 PAD.n767 PAD.n766 0.019716
R49610 PAD.n766 PAD.n765 0.019716
R49611 PAD.n770 PAD.n769 0.019716
R49612 PAD.n869 PAD.n824 0.019716
R49613 PAD.n870 PAD.n823 0.019716
R49614 PAD.n879 PAD.n822 0.019716
R49615 PAD.n879 PAD.n878 0.019716
R49616 PAD.n881 PAD.n821 0.019716
R49617 PAD.n882 PAD.n881 0.019716
R49618 PAD.n891 PAD.n820 0.019716
R49619 PAD.n891 PAD.n890 0.019716
R49620 PAD.n893 PAD.n819 0.019716
R49621 PAD.n894 PAD.n893 0.019716
R49622 PAD.n903 PAD.n818 0.019716
R49623 PAD.n903 PAD.n902 0.019716
R49624 PAD.n905 PAD.n817 0.019716
R49625 PAD.n906 PAD.n905 0.019716
R49626 PAD.n915 PAD.n816 0.019716
R49627 PAD.n915 PAD.n914 0.019716
R49628 PAD.n917 PAD.n815 0.019716
R49629 PAD.n918 PAD.n917 0.019716
R49630 PAD.n927 PAD.n814 0.019716
R49631 PAD.n927 PAD.n926 0.019716
R49632 PAD.n929 PAD.n813 0.019716
R49633 PAD.n930 PAD.n929 0.019716
R49634 PAD.n939 PAD.n812 0.019716
R49635 PAD.n939 PAD.n938 0.019716
R49636 PAD.n941 PAD.n811 0.019716
R49637 PAD.n942 PAD.n941 0.019716
R49638 PAD.n951 PAD.n810 0.019716
R49639 PAD.n951 PAD.n950 0.019716
R49640 PAD.n953 PAD.n809 0.019716
R49641 PAD.n954 PAD.n953 0.019716
R49642 PAD.n963 PAD.n808 0.019716
R49643 PAD.n963 PAD.n962 0.019716
R49644 PAD.n965 PAD.n807 0.019716
R49645 PAD.n966 PAD.n965 0.019716
R49646 PAD.n975 PAD.n806 0.019716
R49647 PAD.n975 PAD.n974 0.019716
R49648 PAD.n977 PAD.n805 0.019716
R49649 PAD.n978 PAD.n977 0.019716
R49650 PAD.n987 PAD.n804 0.019716
R49651 PAD.n987 PAD.n986 0.019716
R49652 PAD.n989 PAD.n803 0.019716
R49653 PAD.n990 PAD.n989 0.019716
R49654 PAD.n999 PAD.n802 0.019716
R49655 PAD.n999 PAD.n998 0.019716
R49656 PAD.n1001 PAD.n801 0.019716
R49657 PAD.n1002 PAD.n1001 0.019716
R49658 PAD.n1011 PAD.n800 0.019716
R49659 PAD.n1011 PAD.n1010 0.019716
R49660 PAD.n1013 PAD.n799 0.019716
R49661 PAD.n1014 PAD.n1013 0.019716
R49662 PAD.n1023 PAD.n798 0.019716
R49663 PAD.n1023 PAD.n1022 0.019716
R49664 PAD.n1025 PAD.n797 0.019716
R49665 PAD.n1026 PAD.n1025 0.019716
R49666 PAD.n1035 PAD.n796 0.019716
R49667 PAD.n1035 PAD.n1034 0.019716
R49668 PAD.n1037 PAD.n795 0.019716
R49669 PAD.n1038 PAD.n1037 0.019716
R49670 PAD.n1047 PAD.n794 0.019716
R49671 PAD.n1047 PAD.n1046 0.019716
R49672 PAD.n1049 PAD.n793 0.019716
R49673 PAD.n1050 PAD.n1049 0.019716
R49674 PAD.n1059 PAD.n792 0.019716
R49675 PAD.n1059 PAD.n1058 0.019716
R49676 PAD.n1061 PAD.n791 0.019716
R49677 PAD.n1062 PAD.n1061 0.019716
R49678 PAD.n1071 PAD.n790 0.019716
R49679 PAD.n1071 PAD.n1070 0.019716
R49680 PAD.n1073 PAD.n789 0.019716
R49681 PAD.n1074 PAD.n1073 0.019716
R49682 PAD.n1083 PAD.n788 0.019716
R49683 PAD.n1083 PAD.n1082 0.019716
R49684 PAD.n1085 PAD.n787 0.019716
R49685 PAD.n1086 PAD.n1085 0.019716
R49686 PAD.n1095 PAD.n786 0.019716
R49687 PAD.n1095 PAD.n1094 0.019716
R49688 PAD.n1097 PAD.n785 0.019716
R49689 PAD.n1098 PAD.n1097 0.019716
R49690 PAD.n1107 PAD.n784 0.019716
R49691 PAD.n1107 PAD.n1106 0.019716
R49692 PAD.n1109 PAD.n783 0.019716
R49693 PAD.n1110 PAD.n1109 0.019716
R49694 PAD.n10387 PAD.n10386 0.019716
R49695 PAD.n10107 PAD.n10106 0.019716
R49696 PAD.n10109 PAD.n10108 0.019716
R49697 PAD.n10110 PAD.n10101 0.019716
R49698 PAD.n10111 PAD.n10110 0.019716
R49699 PAD.n10121 PAD.n10120 0.019716
R49700 PAD.n10120 PAD.n10119 0.019716
R49701 PAD.n10122 PAD.n10097 0.019716
R49702 PAD.n10123 PAD.n10122 0.019716
R49703 PAD.n10133 PAD.n10132 0.019716
R49704 PAD.n10132 PAD.n10131 0.019716
R49705 PAD.n10134 PAD.n10093 0.019716
R49706 PAD.n10135 PAD.n10134 0.019716
R49707 PAD.n10145 PAD.n10144 0.019716
R49708 PAD.n10144 PAD.n10143 0.019716
R49709 PAD.n10146 PAD.n10089 0.019716
R49710 PAD.n10147 PAD.n10146 0.019716
R49711 PAD.n10157 PAD.n10156 0.019716
R49712 PAD.n10156 PAD.n10155 0.019716
R49713 PAD.n10158 PAD.n10085 0.019716
R49714 PAD.n10159 PAD.n10158 0.019716
R49715 PAD.n10169 PAD.n10168 0.019716
R49716 PAD.n10168 PAD.n10167 0.019716
R49717 PAD.n10170 PAD.n10081 0.019716
R49718 PAD.n10171 PAD.n10170 0.019716
R49719 PAD.n10181 PAD.n10180 0.019716
R49720 PAD.n10180 PAD.n10179 0.019716
R49721 PAD.n10182 PAD.n10077 0.019716
R49722 PAD.n10183 PAD.n10182 0.019716
R49723 PAD.n10193 PAD.n10192 0.019716
R49724 PAD.n10192 PAD.n10191 0.019716
R49725 PAD.n10194 PAD.n10073 0.019716
R49726 PAD.n10195 PAD.n10194 0.019716
R49727 PAD.n10205 PAD.n10204 0.019716
R49728 PAD.n10204 PAD.n10203 0.019716
R49729 PAD.n10206 PAD.n10069 0.019716
R49730 PAD.n10207 PAD.n10206 0.019716
R49731 PAD.n10217 PAD.n10216 0.019716
R49732 PAD.n10216 PAD.n10215 0.019716
R49733 PAD.n10218 PAD.n10065 0.019716
R49734 PAD.n10219 PAD.n10218 0.019716
R49735 PAD.n10229 PAD.n10228 0.019716
R49736 PAD.n10228 PAD.n10227 0.019716
R49737 PAD.n10230 PAD.n10061 0.019716
R49738 PAD.n10231 PAD.n10230 0.019716
R49739 PAD.n10241 PAD.n10240 0.019716
R49740 PAD.n10240 PAD.n10239 0.019716
R49741 PAD.n10242 PAD.n10057 0.019716
R49742 PAD.n10243 PAD.n10242 0.019716
R49743 PAD.n10253 PAD.n10252 0.019716
R49744 PAD.n10252 PAD.n10251 0.019716
R49745 PAD.n10254 PAD.n10053 0.019716
R49746 PAD.n10255 PAD.n10254 0.019716
R49747 PAD.n10265 PAD.n10264 0.019716
R49748 PAD.n10264 PAD.n10263 0.019716
R49749 PAD.n10266 PAD.n10049 0.019716
R49750 PAD.n10267 PAD.n10266 0.019716
R49751 PAD.n10277 PAD.n10276 0.019716
R49752 PAD.n10276 PAD.n10275 0.019716
R49753 PAD.n10278 PAD.n10045 0.019716
R49754 PAD.n10279 PAD.n10278 0.019716
R49755 PAD.n10289 PAD.n10288 0.019716
R49756 PAD.n10288 PAD.n10287 0.019716
R49757 PAD.n10290 PAD.n10041 0.019716
R49758 PAD.n10291 PAD.n10290 0.019716
R49759 PAD.n10301 PAD.n10300 0.019716
R49760 PAD.n10300 PAD.n10299 0.019716
R49761 PAD.n10302 PAD.n10037 0.019716
R49762 PAD.n10303 PAD.n10302 0.019716
R49763 PAD.n10313 PAD.n10312 0.019716
R49764 PAD.n10312 PAD.n10311 0.019716
R49765 PAD.n10314 PAD.n10033 0.019716
R49766 PAD.n10315 PAD.n10314 0.019716
R49767 PAD.n10325 PAD.n10324 0.019716
R49768 PAD.n10324 PAD.n10323 0.019716
R49769 PAD.n10326 PAD.n10029 0.019716
R49770 PAD.n10327 PAD.n10326 0.019716
R49771 PAD.n10337 PAD.n10336 0.019716
R49772 PAD.n10336 PAD.n10335 0.019716
R49773 PAD.n10338 PAD.n10025 0.019716
R49774 PAD.n10339 PAD.n10338 0.019716
R49775 PAD.n10350 PAD.n10349 0.019716
R49776 PAD.n10349 PAD.n10348 0.019716
R49777 PAD.n10353 PAD.n10352 0.019716
R49778 PAD.n1482 PAD.n1481 0.019716
R49779 PAD.n1191 PAD.n1190 0.019716
R49780 PAD.n1474 PAD.n1473 0.019716
R49781 PAD.n1474 PAD.n1189 0.019716
R49782 PAD.n1198 PAD.n1197 0.019716
R49783 PAD.n1198 PAD.n1188 0.019716
R49784 PAD.n1465 PAD.n1464 0.019716
R49785 PAD.n1465 PAD.n1187 0.019716
R49786 PAD.n1203 PAD.n1202 0.019716
R49787 PAD.n1203 PAD.n1186 0.019716
R49788 PAD.n1456 PAD.n1455 0.019716
R49789 PAD.n1456 PAD.n1185 0.019716
R49790 PAD.n1208 PAD.n1207 0.019716
R49791 PAD.n1208 PAD.n1184 0.019716
R49792 PAD.n1447 PAD.n1446 0.019716
R49793 PAD.n1447 PAD.n1183 0.019716
R49794 PAD.n1213 PAD.n1212 0.019716
R49795 PAD.n1213 PAD.n1182 0.019716
R49796 PAD.n1438 PAD.n1437 0.019716
R49797 PAD.n1438 PAD.n1181 0.019716
R49798 PAD.n1218 PAD.n1217 0.019716
R49799 PAD.n1218 PAD.n1180 0.019716
R49800 PAD.n1429 PAD.n1428 0.019716
R49801 PAD.n1429 PAD.n1179 0.019716
R49802 PAD.n1223 PAD.n1222 0.019716
R49803 PAD.n1223 PAD.n1178 0.019716
R49804 PAD.n1420 PAD.n1419 0.019716
R49805 PAD.n1420 PAD.n1177 0.019716
R49806 PAD.n1228 PAD.n1227 0.019716
R49807 PAD.n1228 PAD.n1176 0.019716
R49808 PAD.n1411 PAD.n1410 0.019716
R49809 PAD.n1411 PAD.n1175 0.019716
R49810 PAD.n1233 PAD.n1232 0.019716
R49811 PAD.n1233 PAD.n1174 0.019716
R49812 PAD.n1402 PAD.n1401 0.019716
R49813 PAD.n1402 PAD.n1173 0.019716
R49814 PAD.n1238 PAD.n1237 0.019716
R49815 PAD.n1238 PAD.n1172 0.019716
R49816 PAD.n1393 PAD.n1392 0.019716
R49817 PAD.n1393 PAD.n1171 0.019716
R49818 PAD.n1243 PAD.n1242 0.019716
R49819 PAD.n1243 PAD.n1170 0.019716
R49820 PAD.n1384 PAD.n1383 0.019716
R49821 PAD.n1384 PAD.n1169 0.019716
R49822 PAD.n1248 PAD.n1247 0.019716
R49823 PAD.n1248 PAD.n1168 0.019716
R49824 PAD.n1375 PAD.n1374 0.019716
R49825 PAD.n1375 PAD.n1167 0.019716
R49826 PAD.n1253 PAD.n1252 0.019716
R49827 PAD.n1253 PAD.n1166 0.019716
R49828 PAD.n1366 PAD.n1365 0.019716
R49829 PAD.n1366 PAD.n1165 0.019716
R49830 PAD.n1258 PAD.n1257 0.019716
R49831 PAD.n1258 PAD.n1164 0.019716
R49832 PAD.n1357 PAD.n1356 0.019716
R49833 PAD.n1357 PAD.n1163 0.019716
R49834 PAD.n1263 PAD.n1262 0.019716
R49835 PAD.n1263 PAD.n1162 0.019716
R49836 PAD.n1348 PAD.n1347 0.019716
R49837 PAD.n1348 PAD.n1161 0.019716
R49838 PAD.n1268 PAD.n1267 0.019716
R49839 PAD.n1268 PAD.n1160 0.019716
R49840 PAD.n1339 PAD.n1338 0.019716
R49841 PAD.n1339 PAD.n1159 0.019716
R49842 PAD.n1273 PAD.n1272 0.019716
R49843 PAD.n1273 PAD.n1158 0.019716
R49844 PAD.n1330 PAD.n1329 0.019716
R49845 PAD.n1330 PAD.n1157 0.019716
R49846 PAD.n1278 PAD.n1277 0.019716
R49847 PAD.n1278 PAD.n1156 0.019716
R49848 PAD.n1321 PAD.n1320 0.019716
R49849 PAD.n1321 PAD.n1155 0.019716
R49850 PAD.n1283 PAD.n1282 0.019716
R49851 PAD.n1283 PAD.n1154 0.019716
R49852 PAD.n1312 PAD.n1311 0.019716
R49853 PAD.n1312 PAD.n1153 0.019716
R49854 PAD.n1288 PAD.n1287 0.019716
R49855 PAD.n1288 PAD.n1152 0.019716
R49856 PAD.n1303 PAD.n1302 0.019716
R49857 PAD.n1303 PAD.n1151 0.019716
R49858 PAD.n1293 PAD.n1292 0.019716
R49859 PAD.n1293 PAD.n1150 0.019716
R49860 PAD.n1294 PAD.n1149 0.019716
R49861 PAD.n1577 PAD.n1531 0.019716
R49862 PAD.n1578 PAD.n1530 0.019716
R49863 PAD.n9756 PAD.n1529 0.019716
R49864 PAD.n9756 PAD.n9755 0.019716
R49865 PAD.n9758 PAD.n1528 0.019716
R49866 PAD.n9759 PAD.n9758 0.019716
R49867 PAD.n9768 PAD.n1527 0.019716
R49868 PAD.n9768 PAD.n9767 0.019716
R49869 PAD.n9770 PAD.n1526 0.019716
R49870 PAD.n9771 PAD.n9770 0.019716
R49871 PAD.n9780 PAD.n1525 0.019716
R49872 PAD.n9780 PAD.n9779 0.019716
R49873 PAD.n9782 PAD.n1524 0.019716
R49874 PAD.n9783 PAD.n9782 0.019716
R49875 PAD.n9792 PAD.n1523 0.019716
R49876 PAD.n9792 PAD.n9791 0.019716
R49877 PAD.n9794 PAD.n1522 0.019716
R49878 PAD.n9795 PAD.n9794 0.019716
R49879 PAD.n9804 PAD.n1521 0.019716
R49880 PAD.n9804 PAD.n9803 0.019716
R49881 PAD.n9806 PAD.n1520 0.019716
R49882 PAD.n9807 PAD.n9806 0.019716
R49883 PAD.n9816 PAD.n1519 0.019716
R49884 PAD.n9816 PAD.n9815 0.019716
R49885 PAD.n9818 PAD.n1518 0.019716
R49886 PAD.n9819 PAD.n9818 0.019716
R49887 PAD.n9828 PAD.n1517 0.019716
R49888 PAD.n9828 PAD.n9827 0.019716
R49889 PAD.n9830 PAD.n1516 0.019716
R49890 PAD.n9831 PAD.n9830 0.019716
R49891 PAD.n9840 PAD.n1515 0.019716
R49892 PAD.n9840 PAD.n9839 0.019716
R49893 PAD.n9842 PAD.n1514 0.019716
R49894 PAD.n9843 PAD.n9842 0.019716
R49895 PAD.n9852 PAD.n1513 0.019716
R49896 PAD.n9852 PAD.n9851 0.019716
R49897 PAD.n9854 PAD.n1512 0.019716
R49898 PAD.n9855 PAD.n9854 0.019716
R49899 PAD.n9864 PAD.n1511 0.019716
R49900 PAD.n9864 PAD.n9863 0.019716
R49901 PAD.n9866 PAD.n1510 0.019716
R49902 PAD.n9867 PAD.n9866 0.019716
R49903 PAD.n9876 PAD.n1509 0.019716
R49904 PAD.n9876 PAD.n9875 0.019716
R49905 PAD.n9878 PAD.n1508 0.019716
R49906 PAD.n9879 PAD.n9878 0.019716
R49907 PAD.n9888 PAD.n1507 0.019716
R49908 PAD.n9888 PAD.n9887 0.019716
R49909 PAD.n9890 PAD.n1506 0.019716
R49910 PAD.n9891 PAD.n9890 0.019716
R49911 PAD.n9900 PAD.n1505 0.019716
R49912 PAD.n9900 PAD.n9899 0.019716
R49913 PAD.n9902 PAD.n1504 0.019716
R49914 PAD.n9903 PAD.n9902 0.019716
R49915 PAD.n9912 PAD.n1503 0.019716
R49916 PAD.n9912 PAD.n9911 0.019716
R49917 PAD.n9914 PAD.n1502 0.019716
R49918 PAD.n9915 PAD.n9914 0.019716
R49919 PAD.n9924 PAD.n1501 0.019716
R49920 PAD.n9924 PAD.n9923 0.019716
R49921 PAD.n9926 PAD.n1500 0.019716
R49922 PAD.n9927 PAD.n9926 0.019716
R49923 PAD.n9936 PAD.n1499 0.019716
R49924 PAD.n9936 PAD.n9935 0.019716
R49925 PAD.n9938 PAD.n1498 0.019716
R49926 PAD.n9939 PAD.n9938 0.019716
R49927 PAD.n9948 PAD.n1497 0.019716
R49928 PAD.n9948 PAD.n9947 0.019716
R49929 PAD.n9950 PAD.n1496 0.019716
R49930 PAD.n9951 PAD.n9950 0.019716
R49931 PAD.n9960 PAD.n1495 0.019716
R49932 PAD.n9960 PAD.n9959 0.019716
R49933 PAD.n9962 PAD.n1494 0.019716
R49934 PAD.n9963 PAD.n9962 0.019716
R49935 PAD.n9972 PAD.n1493 0.019716
R49936 PAD.n9972 PAD.n9971 0.019716
R49937 PAD.n9974 PAD.n1492 0.019716
R49938 PAD.n9975 PAD.n9974 0.019716
R49939 PAD.n9984 PAD.n1491 0.019716
R49940 PAD.n9984 PAD.n9983 0.019716
R49941 PAD.n9986 PAD.n1490 0.019716
R49942 PAD.n9987 PAD.n9986 0.019716
R49943 PAD.n9997 PAD.n9996 0.019716
R49944 PAD.n1601 PAD.n1599 0.019716
R49945 PAD.n1929 PAD.n1928 0.019716
R49946 PAD.n1925 PAD.n1602 0.019716
R49947 PAD.n1926 PAD.n1925 0.019716
R49948 PAD.n1919 PAD.n1916 0.019716
R49949 PAD.n1919 PAD.n1918 0.019716
R49950 PAD.n1913 PAD.n1607 0.019716
R49951 PAD.n1914 PAD.n1913 0.019716
R49952 PAD.n1907 PAD.n1904 0.019716
R49953 PAD.n1907 PAD.n1906 0.019716
R49954 PAD.n1901 PAD.n1611 0.019716
R49955 PAD.n1902 PAD.n1901 0.019716
R49956 PAD.n1895 PAD.n1892 0.019716
R49957 PAD.n1895 PAD.n1894 0.019716
R49958 PAD.n1889 PAD.n1615 0.019716
R49959 PAD.n1890 PAD.n1889 0.019716
R49960 PAD.n1883 PAD.n1880 0.019716
R49961 PAD.n1883 PAD.n1882 0.019716
R49962 PAD.n1877 PAD.n1619 0.019716
R49963 PAD.n1878 PAD.n1877 0.019716
R49964 PAD.n1871 PAD.n1868 0.019716
R49965 PAD.n1871 PAD.n1870 0.019716
R49966 PAD.n1865 PAD.n1623 0.019716
R49967 PAD.n1866 PAD.n1865 0.019716
R49968 PAD.n1859 PAD.n1856 0.019716
R49969 PAD.n1859 PAD.n1858 0.019716
R49970 PAD.n1853 PAD.n1627 0.019716
R49971 PAD.n1854 PAD.n1853 0.019716
R49972 PAD.n1847 PAD.n1844 0.019716
R49973 PAD.n1847 PAD.n1846 0.019716
R49974 PAD.n1841 PAD.n1631 0.019716
R49975 PAD.n1842 PAD.n1841 0.019716
R49976 PAD.n1835 PAD.n1832 0.019716
R49977 PAD.n1835 PAD.n1834 0.019716
R49978 PAD.n1829 PAD.n1635 0.019716
R49979 PAD.n1830 PAD.n1829 0.019716
R49980 PAD.n1823 PAD.n1820 0.019716
R49981 PAD.n1823 PAD.n1822 0.019716
R49982 PAD.n1817 PAD.n1639 0.019716
R49983 PAD.n1818 PAD.n1817 0.019716
R49984 PAD.n1811 PAD.n1808 0.019716
R49985 PAD.n1811 PAD.n1810 0.019716
R49986 PAD.n1805 PAD.n1643 0.019716
R49987 PAD.n1806 PAD.n1805 0.019716
R49988 PAD.n1799 PAD.n1796 0.019716
R49989 PAD.n1799 PAD.n1798 0.019716
R49990 PAD.n1793 PAD.n1647 0.019716
R49991 PAD.n1794 PAD.n1793 0.019716
R49992 PAD.n1787 PAD.n1784 0.019716
R49993 PAD.n1787 PAD.n1786 0.019716
R49994 PAD.n1781 PAD.n1651 0.019716
R49995 PAD.n1782 PAD.n1781 0.019716
R49996 PAD.n1775 PAD.n1772 0.019716
R49997 PAD.n1775 PAD.n1774 0.019716
R49998 PAD.n1769 PAD.n1655 0.019716
R49999 PAD.n1770 PAD.n1769 0.019716
R50000 PAD.n1763 PAD.n1760 0.019716
R50001 PAD.n1763 PAD.n1762 0.019716
R50002 PAD.n1757 PAD.n1659 0.019716
R50003 PAD.n1758 PAD.n1757 0.019716
R50004 PAD.n1751 PAD.n1748 0.019716
R50005 PAD.n1751 PAD.n1750 0.019716
R50006 PAD.n1745 PAD.n1663 0.019716
R50007 PAD.n1746 PAD.n1745 0.019716
R50008 PAD.n1739 PAD.n1736 0.019716
R50009 PAD.n1739 PAD.n1738 0.019716
R50010 PAD.n1733 PAD.n1667 0.019716
R50011 PAD.n1734 PAD.n1733 0.019716
R50012 PAD.n1727 PAD.n1724 0.019716
R50013 PAD.n1727 PAD.n1726 0.019716
R50014 PAD.n1721 PAD.n1671 0.019716
R50015 PAD.n1722 PAD.n1721 0.019716
R50016 PAD.n1715 PAD.n1712 0.019716
R50017 PAD.n1715 PAD.n1714 0.019716
R50018 PAD.n1709 PAD.n1675 0.019716
R50019 PAD.n1710 PAD.n1709 0.019716
R50020 PAD.n1703 PAD.n1700 0.019716
R50021 PAD.n1703 PAD.n1702 0.019716
R50022 PAD.n1697 PAD.n1679 0.019716
R50023 PAD.n1698 PAD.n1697 0.019716
R50024 PAD.n1691 PAD.n1688 0.019716
R50025 PAD.n1691 PAD.n1690 0.019716
R50026 PAD.n1686 PAD.n1685 0.019716
R50027 PAD.n2029 PAD.n1984 0.019716
R50028 PAD.n2030 PAD.n1983 0.019716
R50029 PAD.n9470 PAD.n1982 0.019716
R50030 PAD.n9470 PAD.n9469 0.019716
R50031 PAD.n9472 PAD.n1981 0.019716
R50032 PAD.n9473 PAD.n9472 0.019716
R50033 PAD.n9482 PAD.n1980 0.019716
R50034 PAD.n9482 PAD.n9481 0.019716
R50035 PAD.n9484 PAD.n1979 0.019716
R50036 PAD.n9485 PAD.n9484 0.019716
R50037 PAD.n9494 PAD.n1978 0.019716
R50038 PAD.n9494 PAD.n9493 0.019716
R50039 PAD.n9496 PAD.n1977 0.019716
R50040 PAD.n9497 PAD.n9496 0.019716
R50041 PAD.n9506 PAD.n1976 0.019716
R50042 PAD.n9506 PAD.n9505 0.019716
R50043 PAD.n9508 PAD.n1975 0.019716
R50044 PAD.n9509 PAD.n9508 0.019716
R50045 PAD.n9518 PAD.n1974 0.019716
R50046 PAD.n9518 PAD.n9517 0.019716
R50047 PAD.n9520 PAD.n1973 0.019716
R50048 PAD.n9521 PAD.n9520 0.019716
R50049 PAD.n9530 PAD.n1972 0.019716
R50050 PAD.n9530 PAD.n9529 0.019716
R50051 PAD.n9532 PAD.n1971 0.019716
R50052 PAD.n9533 PAD.n9532 0.019716
R50053 PAD.n9542 PAD.n1970 0.019716
R50054 PAD.n9542 PAD.n9541 0.019716
R50055 PAD.n9544 PAD.n1969 0.019716
R50056 PAD.n9545 PAD.n9544 0.019716
R50057 PAD.n9554 PAD.n1968 0.019716
R50058 PAD.n9554 PAD.n9553 0.019716
R50059 PAD.n9556 PAD.n1967 0.019716
R50060 PAD.n9557 PAD.n9556 0.019716
R50061 PAD.n9566 PAD.n1966 0.019716
R50062 PAD.n9566 PAD.n9565 0.019716
R50063 PAD.n9568 PAD.n1965 0.019716
R50064 PAD.n9569 PAD.n9568 0.019716
R50065 PAD.n9578 PAD.n1964 0.019716
R50066 PAD.n9578 PAD.n9577 0.019716
R50067 PAD.n9580 PAD.n1963 0.019716
R50068 PAD.n9581 PAD.n9580 0.019716
R50069 PAD.n9590 PAD.n1962 0.019716
R50070 PAD.n9590 PAD.n9589 0.019716
R50071 PAD.n9592 PAD.n1961 0.019716
R50072 PAD.n9593 PAD.n9592 0.019716
R50073 PAD.n9602 PAD.n1960 0.019716
R50074 PAD.n9602 PAD.n9601 0.019716
R50075 PAD.n9604 PAD.n1959 0.019716
R50076 PAD.n9605 PAD.n9604 0.019716
R50077 PAD.n9614 PAD.n1958 0.019716
R50078 PAD.n9614 PAD.n9613 0.019716
R50079 PAD.n9616 PAD.n1957 0.019716
R50080 PAD.n9617 PAD.n9616 0.019716
R50081 PAD.n9626 PAD.n1956 0.019716
R50082 PAD.n9626 PAD.n9625 0.019716
R50083 PAD.n9628 PAD.n1955 0.019716
R50084 PAD.n9629 PAD.n9628 0.019716
R50085 PAD.n9638 PAD.n1954 0.019716
R50086 PAD.n9638 PAD.n9637 0.019716
R50087 PAD.n9640 PAD.n1953 0.019716
R50088 PAD.n9641 PAD.n9640 0.019716
R50089 PAD.n9650 PAD.n1952 0.019716
R50090 PAD.n9650 PAD.n9649 0.019716
R50091 PAD.n9652 PAD.n1951 0.019716
R50092 PAD.n9653 PAD.n9652 0.019716
R50093 PAD.n9662 PAD.n1950 0.019716
R50094 PAD.n9662 PAD.n9661 0.019716
R50095 PAD.n9664 PAD.n1949 0.019716
R50096 PAD.n9665 PAD.n9664 0.019716
R50097 PAD.n9674 PAD.n1948 0.019716
R50098 PAD.n9674 PAD.n9673 0.019716
R50099 PAD.n9676 PAD.n1947 0.019716
R50100 PAD.n9677 PAD.n9676 0.019716
R50101 PAD.n9686 PAD.n1946 0.019716
R50102 PAD.n9686 PAD.n9685 0.019716
R50103 PAD.n9688 PAD.n1945 0.019716
R50104 PAD.n9689 PAD.n9688 0.019716
R50105 PAD.n9698 PAD.n1944 0.019716
R50106 PAD.n9698 PAD.n9697 0.019716
R50107 PAD.n9700 PAD.n1943 0.019716
R50108 PAD.n9701 PAD.n9700 0.019716
R50109 PAD.n9711 PAD.n9710 0.019716
R50110 PAD.n2132 PAD.n2088 0.019716
R50111 PAD.n2133 PAD.n2087 0.019716
R50112 PAD.n9204 PAD.n2086 0.019716
R50113 PAD.n9204 PAD.n9203 0.019716
R50114 PAD.n9206 PAD.n2085 0.019716
R50115 PAD.n9207 PAD.n9206 0.019716
R50116 PAD.n9216 PAD.n2084 0.019716
R50117 PAD.n9216 PAD.n9215 0.019716
R50118 PAD.n9218 PAD.n2083 0.019716
R50119 PAD.n9219 PAD.n9218 0.019716
R50120 PAD.n9228 PAD.n2082 0.019716
R50121 PAD.n9228 PAD.n9227 0.019716
R50122 PAD.n9230 PAD.n2081 0.019716
R50123 PAD.n9231 PAD.n9230 0.019716
R50124 PAD.n9240 PAD.n2080 0.019716
R50125 PAD.n9240 PAD.n9239 0.019716
R50126 PAD.n9242 PAD.n2079 0.019716
R50127 PAD.n9243 PAD.n9242 0.019716
R50128 PAD.n9252 PAD.n2078 0.019716
R50129 PAD.n9252 PAD.n9251 0.019716
R50130 PAD.n9254 PAD.n2077 0.019716
R50131 PAD.n9255 PAD.n9254 0.019716
R50132 PAD.n9264 PAD.n2076 0.019716
R50133 PAD.n9264 PAD.n9263 0.019716
R50134 PAD.n9266 PAD.n2075 0.019716
R50135 PAD.n9267 PAD.n9266 0.019716
R50136 PAD.n9276 PAD.n2074 0.019716
R50137 PAD.n9276 PAD.n9275 0.019716
R50138 PAD.n9278 PAD.n2073 0.019716
R50139 PAD.n9279 PAD.n9278 0.019716
R50140 PAD.n9288 PAD.n2072 0.019716
R50141 PAD.n9288 PAD.n9287 0.019716
R50142 PAD.n9290 PAD.n2071 0.019716
R50143 PAD.n9291 PAD.n9290 0.019716
R50144 PAD.n9300 PAD.n2070 0.019716
R50145 PAD.n9300 PAD.n9299 0.019716
R50146 PAD.n9302 PAD.n2069 0.019716
R50147 PAD.n9303 PAD.n9302 0.019716
R50148 PAD.n9312 PAD.n2068 0.019716
R50149 PAD.n9312 PAD.n9311 0.019716
R50150 PAD.n9314 PAD.n2067 0.019716
R50151 PAD.n9315 PAD.n9314 0.019716
R50152 PAD.n9324 PAD.n2066 0.019716
R50153 PAD.n9324 PAD.n9323 0.019716
R50154 PAD.n9326 PAD.n2065 0.019716
R50155 PAD.n9327 PAD.n9326 0.019716
R50156 PAD.n9336 PAD.n2064 0.019716
R50157 PAD.n9336 PAD.n9335 0.019716
R50158 PAD.n9338 PAD.n2063 0.019716
R50159 PAD.n9339 PAD.n9338 0.019716
R50160 PAD.n9348 PAD.n2062 0.019716
R50161 PAD.n9348 PAD.n9347 0.019716
R50162 PAD.n9350 PAD.n2061 0.019716
R50163 PAD.n9351 PAD.n9350 0.019716
R50164 PAD.n9360 PAD.n2060 0.019716
R50165 PAD.n9360 PAD.n9359 0.019716
R50166 PAD.n9362 PAD.n2059 0.019716
R50167 PAD.n9363 PAD.n9362 0.019716
R50168 PAD.n9372 PAD.n2058 0.019716
R50169 PAD.n9372 PAD.n9371 0.019716
R50170 PAD.n9374 PAD.n2057 0.019716
R50171 PAD.n9375 PAD.n9374 0.019716
R50172 PAD.n9384 PAD.n2056 0.019716
R50173 PAD.n9384 PAD.n9383 0.019716
R50174 PAD.n9386 PAD.n2055 0.019716
R50175 PAD.n9387 PAD.n9386 0.019716
R50176 PAD.n9396 PAD.n2054 0.019716
R50177 PAD.n9396 PAD.n9395 0.019716
R50178 PAD.n9398 PAD.n2053 0.019716
R50179 PAD.n9399 PAD.n9398 0.019716
R50180 PAD.n9408 PAD.n2052 0.019716
R50181 PAD.n9408 PAD.n9407 0.019716
R50182 PAD.n9410 PAD.n2051 0.019716
R50183 PAD.n9411 PAD.n9410 0.019716
R50184 PAD.n9420 PAD.n2050 0.019716
R50185 PAD.n9420 PAD.n9419 0.019716
R50186 PAD.n9422 PAD.n2049 0.019716
R50187 PAD.n9423 PAD.n9422 0.019716
R50188 PAD.n9432 PAD.n2048 0.019716
R50189 PAD.n9432 PAD.n9431 0.019716
R50190 PAD.n9434 PAD.n2047 0.019716
R50191 PAD.n9435 PAD.n9434 0.019716
R50192 PAD.n9444 PAD.n9443 0.019716
R50193 PAD.n2153 PAD.n2151 0.019716
R50194 PAD.n2480 PAD.n2479 0.019716
R50195 PAD.n2476 PAD.n2154 0.019716
R50196 PAD.n2477 PAD.n2476 0.019716
R50197 PAD.n2470 PAD.n2467 0.019716
R50198 PAD.n2470 PAD.n2469 0.019716
R50199 PAD.n2464 PAD.n2159 0.019716
R50200 PAD.n2465 PAD.n2464 0.019716
R50201 PAD.n2458 PAD.n2455 0.019716
R50202 PAD.n2458 PAD.n2457 0.019716
R50203 PAD.n2452 PAD.n2163 0.019716
R50204 PAD.n2453 PAD.n2452 0.019716
R50205 PAD.n2446 PAD.n2443 0.019716
R50206 PAD.n2446 PAD.n2445 0.019716
R50207 PAD.n2440 PAD.n2167 0.019716
R50208 PAD.n2441 PAD.n2440 0.019716
R50209 PAD.n2434 PAD.n2431 0.019716
R50210 PAD.n2434 PAD.n2433 0.019716
R50211 PAD.n2428 PAD.n2171 0.019716
R50212 PAD.n2429 PAD.n2428 0.019716
R50213 PAD.n2422 PAD.n2419 0.019716
R50214 PAD.n2422 PAD.n2421 0.019716
R50215 PAD.n2416 PAD.n2175 0.019716
R50216 PAD.n2417 PAD.n2416 0.019716
R50217 PAD.n2410 PAD.n2407 0.019716
R50218 PAD.n2410 PAD.n2409 0.019716
R50219 PAD.n2404 PAD.n2179 0.019716
R50220 PAD.n2405 PAD.n2404 0.019716
R50221 PAD.n2398 PAD.n2395 0.019716
R50222 PAD.n2398 PAD.n2397 0.019716
R50223 PAD.n2392 PAD.n2183 0.019716
R50224 PAD.n2393 PAD.n2392 0.019716
R50225 PAD.n2386 PAD.n2383 0.019716
R50226 PAD.n2386 PAD.n2385 0.019716
R50227 PAD.n2380 PAD.n2187 0.019716
R50228 PAD.n2381 PAD.n2380 0.019716
R50229 PAD.n2374 PAD.n2371 0.019716
R50230 PAD.n2374 PAD.n2373 0.019716
R50231 PAD.n2368 PAD.n2191 0.019716
R50232 PAD.n2369 PAD.n2368 0.019716
R50233 PAD.n2362 PAD.n2359 0.019716
R50234 PAD.n2362 PAD.n2361 0.019716
R50235 PAD.n2356 PAD.n2195 0.019716
R50236 PAD.n2357 PAD.n2356 0.019716
R50237 PAD.n2350 PAD.n2347 0.019716
R50238 PAD.n2350 PAD.n2349 0.019716
R50239 PAD.n2344 PAD.n2199 0.019716
R50240 PAD.n2345 PAD.n2344 0.019716
R50241 PAD.n2338 PAD.n2335 0.019716
R50242 PAD.n2338 PAD.n2337 0.019716
R50243 PAD.n2332 PAD.n2203 0.019716
R50244 PAD.n2333 PAD.n2332 0.019716
R50245 PAD.n2326 PAD.n2323 0.019716
R50246 PAD.n2326 PAD.n2325 0.019716
R50247 PAD.n2320 PAD.n2207 0.019716
R50248 PAD.n2321 PAD.n2320 0.019716
R50249 PAD.n2314 PAD.n2311 0.019716
R50250 PAD.n2314 PAD.n2313 0.019716
R50251 PAD.n2308 PAD.n2211 0.019716
R50252 PAD.n2309 PAD.n2308 0.019716
R50253 PAD.n2302 PAD.n2299 0.019716
R50254 PAD.n2302 PAD.n2301 0.019716
R50255 PAD.n2296 PAD.n2215 0.019716
R50256 PAD.n2297 PAD.n2296 0.019716
R50257 PAD.n2290 PAD.n2287 0.019716
R50258 PAD.n2290 PAD.n2289 0.019716
R50259 PAD.n2284 PAD.n2219 0.019716
R50260 PAD.n2285 PAD.n2284 0.019716
R50261 PAD.n2278 PAD.n2275 0.019716
R50262 PAD.n2278 PAD.n2277 0.019716
R50263 PAD.n2272 PAD.n2223 0.019716
R50264 PAD.n2273 PAD.n2272 0.019716
R50265 PAD.n2266 PAD.n2263 0.019716
R50266 PAD.n2266 PAD.n2265 0.019716
R50267 PAD.n2260 PAD.n2227 0.019716
R50268 PAD.n2261 PAD.n2260 0.019716
R50269 PAD.n2254 PAD.n2251 0.019716
R50270 PAD.n2254 PAD.n2253 0.019716
R50271 PAD.n2248 PAD.n2231 0.019716
R50272 PAD.n2249 PAD.n2248 0.019716
R50273 PAD.n2242 PAD.n2239 0.019716
R50274 PAD.n2242 PAD.n2241 0.019716
R50275 PAD.n2237 PAD.n2236 0.019716
R50276 PAD.n2500 PAD.n2498 0.019716
R50277 PAD.n2827 PAD.n2826 0.019716
R50278 PAD.n2823 PAD.n2501 0.019716
R50279 PAD.n2824 PAD.n2823 0.019716
R50280 PAD.n2817 PAD.n2814 0.019716
R50281 PAD.n2817 PAD.n2816 0.019716
R50282 PAD.n2811 PAD.n2506 0.019716
R50283 PAD.n2812 PAD.n2811 0.019716
R50284 PAD.n2805 PAD.n2802 0.019716
R50285 PAD.n2805 PAD.n2804 0.019716
R50286 PAD.n2799 PAD.n2510 0.019716
R50287 PAD.n2800 PAD.n2799 0.019716
R50288 PAD.n2793 PAD.n2790 0.019716
R50289 PAD.n2793 PAD.n2792 0.019716
R50290 PAD.n2787 PAD.n2514 0.019716
R50291 PAD.n2788 PAD.n2787 0.019716
R50292 PAD.n2781 PAD.n2778 0.019716
R50293 PAD.n2781 PAD.n2780 0.019716
R50294 PAD.n2775 PAD.n2518 0.019716
R50295 PAD.n2776 PAD.n2775 0.019716
R50296 PAD.n2769 PAD.n2766 0.019716
R50297 PAD.n2769 PAD.n2768 0.019716
R50298 PAD.n2763 PAD.n2522 0.019716
R50299 PAD.n2764 PAD.n2763 0.019716
R50300 PAD.n2757 PAD.n2754 0.019716
R50301 PAD.n2757 PAD.n2756 0.019716
R50302 PAD.n2751 PAD.n2526 0.019716
R50303 PAD.n2752 PAD.n2751 0.019716
R50304 PAD.n2745 PAD.n2742 0.019716
R50305 PAD.n2745 PAD.n2744 0.019716
R50306 PAD.n2739 PAD.n2530 0.019716
R50307 PAD.n2740 PAD.n2739 0.019716
R50308 PAD.n2733 PAD.n2730 0.019716
R50309 PAD.n2733 PAD.n2732 0.019716
R50310 PAD.n2727 PAD.n2534 0.019716
R50311 PAD.n2728 PAD.n2727 0.019716
R50312 PAD.n2721 PAD.n2718 0.019716
R50313 PAD.n2721 PAD.n2720 0.019716
R50314 PAD.n2715 PAD.n2538 0.019716
R50315 PAD.n2716 PAD.n2715 0.019716
R50316 PAD.n2709 PAD.n2706 0.019716
R50317 PAD.n2709 PAD.n2708 0.019716
R50318 PAD.n2703 PAD.n2542 0.019716
R50319 PAD.n2704 PAD.n2703 0.019716
R50320 PAD.n2697 PAD.n2694 0.019716
R50321 PAD.n2697 PAD.n2696 0.019716
R50322 PAD.n2691 PAD.n2546 0.019716
R50323 PAD.n2692 PAD.n2691 0.019716
R50324 PAD.n2685 PAD.n2682 0.019716
R50325 PAD.n2685 PAD.n2684 0.019716
R50326 PAD.n2679 PAD.n2550 0.019716
R50327 PAD.n2680 PAD.n2679 0.019716
R50328 PAD.n2673 PAD.n2670 0.019716
R50329 PAD.n2673 PAD.n2672 0.019716
R50330 PAD.n2667 PAD.n2554 0.019716
R50331 PAD.n2668 PAD.n2667 0.019716
R50332 PAD.n2661 PAD.n2658 0.019716
R50333 PAD.n2661 PAD.n2660 0.019716
R50334 PAD.n2655 PAD.n2558 0.019716
R50335 PAD.n2656 PAD.n2655 0.019716
R50336 PAD.n2649 PAD.n2646 0.019716
R50337 PAD.n2649 PAD.n2648 0.019716
R50338 PAD.n2643 PAD.n2562 0.019716
R50339 PAD.n2644 PAD.n2643 0.019716
R50340 PAD.n2637 PAD.n2634 0.019716
R50341 PAD.n2637 PAD.n2636 0.019716
R50342 PAD.n2631 PAD.n2566 0.019716
R50343 PAD.n2632 PAD.n2631 0.019716
R50344 PAD.n2625 PAD.n2622 0.019716
R50345 PAD.n2625 PAD.n2624 0.019716
R50346 PAD.n2619 PAD.n2570 0.019716
R50347 PAD.n2620 PAD.n2619 0.019716
R50348 PAD.n2613 PAD.n2610 0.019716
R50349 PAD.n2613 PAD.n2612 0.019716
R50350 PAD.n2607 PAD.n2574 0.019716
R50351 PAD.n2608 PAD.n2607 0.019716
R50352 PAD.n2601 PAD.n2598 0.019716
R50353 PAD.n2601 PAD.n2600 0.019716
R50354 PAD.n2595 PAD.n2578 0.019716
R50355 PAD.n2596 PAD.n2595 0.019716
R50356 PAD.n2589 PAD.n2586 0.019716
R50357 PAD.n2589 PAD.n2588 0.019716
R50358 PAD.n2584 PAD.n2583 0.019716
R50359 PAD.n9116 PAD.n2876 0.019716
R50360 PAD.n9117 PAD.n2875 0.019716
R50361 PAD.n8839 PAD.n2874 0.019716
R50362 PAD.n8840 PAD.n8839 0.019716
R50363 PAD.n9108 PAD.n2873 0.019716
R50364 PAD.n9109 PAD.n9108 0.019716
R50365 PAD.n8844 PAD.n2872 0.019716
R50366 PAD.n8845 PAD.n8844 0.019716
R50367 PAD.n9099 PAD.n2871 0.019716
R50368 PAD.n9100 PAD.n9099 0.019716
R50369 PAD.n8849 PAD.n2870 0.019716
R50370 PAD.n8850 PAD.n8849 0.019716
R50371 PAD.n9090 PAD.n2869 0.019716
R50372 PAD.n9091 PAD.n9090 0.019716
R50373 PAD.n8854 PAD.n2868 0.019716
R50374 PAD.n8855 PAD.n8854 0.019716
R50375 PAD.n9081 PAD.n2867 0.019716
R50376 PAD.n9082 PAD.n9081 0.019716
R50377 PAD.n8859 PAD.n2866 0.019716
R50378 PAD.n8860 PAD.n8859 0.019716
R50379 PAD.n9072 PAD.n2865 0.019716
R50380 PAD.n9073 PAD.n9072 0.019716
R50381 PAD.n8864 PAD.n2864 0.019716
R50382 PAD.n8865 PAD.n8864 0.019716
R50383 PAD.n9063 PAD.n2863 0.019716
R50384 PAD.n9064 PAD.n9063 0.019716
R50385 PAD.n8869 PAD.n2862 0.019716
R50386 PAD.n8870 PAD.n8869 0.019716
R50387 PAD.n9054 PAD.n2861 0.019716
R50388 PAD.n9055 PAD.n9054 0.019716
R50389 PAD.n8874 PAD.n2860 0.019716
R50390 PAD.n8875 PAD.n8874 0.019716
R50391 PAD.n9045 PAD.n2859 0.019716
R50392 PAD.n9046 PAD.n9045 0.019716
R50393 PAD.n8879 PAD.n2858 0.019716
R50394 PAD.n8880 PAD.n8879 0.019716
R50395 PAD.n9036 PAD.n2857 0.019716
R50396 PAD.n9037 PAD.n9036 0.019716
R50397 PAD.n8884 PAD.n2856 0.019716
R50398 PAD.n8885 PAD.n8884 0.019716
R50399 PAD.n9027 PAD.n2855 0.019716
R50400 PAD.n9028 PAD.n9027 0.019716
R50401 PAD.n8889 PAD.n2854 0.019716
R50402 PAD.n8890 PAD.n8889 0.019716
R50403 PAD.n9018 PAD.n2853 0.019716
R50404 PAD.n9019 PAD.n9018 0.019716
R50405 PAD.n8894 PAD.n2852 0.019716
R50406 PAD.n8895 PAD.n8894 0.019716
R50407 PAD.n9009 PAD.n2851 0.019716
R50408 PAD.n9010 PAD.n9009 0.019716
R50409 PAD.n8899 PAD.n2850 0.019716
R50410 PAD.n8900 PAD.n8899 0.019716
R50411 PAD.n9000 PAD.n2849 0.019716
R50412 PAD.n9001 PAD.n9000 0.019716
R50413 PAD.n8904 PAD.n2848 0.019716
R50414 PAD.n8905 PAD.n8904 0.019716
R50415 PAD.n8991 PAD.n2847 0.019716
R50416 PAD.n8992 PAD.n8991 0.019716
R50417 PAD.n8909 PAD.n2846 0.019716
R50418 PAD.n8910 PAD.n8909 0.019716
R50419 PAD.n8982 PAD.n2845 0.019716
R50420 PAD.n8983 PAD.n8982 0.019716
R50421 PAD.n8914 PAD.n2844 0.019716
R50422 PAD.n8915 PAD.n8914 0.019716
R50423 PAD.n8973 PAD.n2843 0.019716
R50424 PAD.n8974 PAD.n8973 0.019716
R50425 PAD.n8919 PAD.n2842 0.019716
R50426 PAD.n8920 PAD.n8919 0.019716
R50427 PAD.n8964 PAD.n2841 0.019716
R50428 PAD.n8965 PAD.n8964 0.019716
R50429 PAD.n8924 PAD.n2840 0.019716
R50430 PAD.n8925 PAD.n8924 0.019716
R50431 PAD.n8955 PAD.n2839 0.019716
R50432 PAD.n8956 PAD.n8955 0.019716
R50433 PAD.n8929 PAD.n2838 0.019716
R50434 PAD.n8930 PAD.n8929 0.019716
R50435 PAD.n8946 PAD.n2837 0.019716
R50436 PAD.n8947 PAD.n8946 0.019716
R50437 PAD.n8934 PAD.n2836 0.019716
R50438 PAD.n8935 PAD.n8934 0.019716
R50439 PAD.n8937 PAD.n2835 0.019716
R50440 PAD.n8938 PAD.n8937 0.019716
R50441 PAD.n9139 PAD.n9138 0.019716
R50442 PAD.n8820 PAD.n8819 0.019716
R50443 PAD.n8812 PAD.n8528 0.019716
R50444 PAD.n8810 PAD.n8809 0.019716
R50445 PAD.n8810 PAD.n2945 0.019716
R50446 PAD.n8801 PAD.n8800 0.019716
R50447 PAD.n8800 PAD.n2944 0.019716
R50448 PAD.n8798 PAD.n8797 0.019716
R50449 PAD.n8798 PAD.n2943 0.019716
R50450 PAD.n8789 PAD.n8788 0.019716
R50451 PAD.n8788 PAD.n2942 0.019716
R50452 PAD.n8786 PAD.n8785 0.019716
R50453 PAD.n8786 PAD.n2941 0.019716
R50454 PAD.n8777 PAD.n8776 0.019716
R50455 PAD.n8776 PAD.n2940 0.019716
R50456 PAD.n8774 PAD.n8773 0.019716
R50457 PAD.n8774 PAD.n2939 0.019716
R50458 PAD.n8765 PAD.n8764 0.019716
R50459 PAD.n8764 PAD.n2938 0.019716
R50460 PAD.n8762 PAD.n8761 0.019716
R50461 PAD.n8762 PAD.n2937 0.019716
R50462 PAD.n8753 PAD.n8752 0.019716
R50463 PAD.n8752 PAD.n2936 0.019716
R50464 PAD.n8750 PAD.n8749 0.019716
R50465 PAD.n8750 PAD.n2935 0.019716
R50466 PAD.n8741 PAD.n8740 0.019716
R50467 PAD.n8740 PAD.n2934 0.019716
R50468 PAD.n8738 PAD.n8737 0.019716
R50469 PAD.n8738 PAD.n2933 0.019716
R50470 PAD.n8729 PAD.n8728 0.019716
R50471 PAD.n8728 PAD.n2932 0.019716
R50472 PAD.n8726 PAD.n8725 0.019716
R50473 PAD.n8726 PAD.n2931 0.019716
R50474 PAD.n8717 PAD.n8716 0.019716
R50475 PAD.n8716 PAD.n2930 0.019716
R50476 PAD.n8714 PAD.n8713 0.019716
R50477 PAD.n8714 PAD.n2929 0.019716
R50478 PAD.n8705 PAD.n8704 0.019716
R50479 PAD.n8704 PAD.n2928 0.019716
R50480 PAD.n8702 PAD.n8701 0.019716
R50481 PAD.n8702 PAD.n2927 0.019716
R50482 PAD.n8693 PAD.n8692 0.019716
R50483 PAD.n8692 PAD.n2926 0.019716
R50484 PAD.n8690 PAD.n8689 0.019716
R50485 PAD.n8690 PAD.n2925 0.019716
R50486 PAD.n8681 PAD.n8680 0.019716
R50487 PAD.n8680 PAD.n2924 0.019716
R50488 PAD.n8678 PAD.n8677 0.019716
R50489 PAD.n8678 PAD.n2923 0.019716
R50490 PAD.n8669 PAD.n8668 0.019716
R50491 PAD.n8668 PAD.n2922 0.019716
R50492 PAD.n8666 PAD.n8665 0.019716
R50493 PAD.n8666 PAD.n2921 0.019716
R50494 PAD.n8657 PAD.n8656 0.019716
R50495 PAD.n8656 PAD.n2920 0.019716
R50496 PAD.n8654 PAD.n8653 0.019716
R50497 PAD.n8654 PAD.n2919 0.019716
R50498 PAD.n8645 PAD.n8644 0.019716
R50499 PAD.n8644 PAD.n2918 0.019716
R50500 PAD.n8642 PAD.n8641 0.019716
R50501 PAD.n8642 PAD.n2917 0.019716
R50502 PAD.n8633 PAD.n8632 0.019716
R50503 PAD.n8632 PAD.n2916 0.019716
R50504 PAD.n8630 PAD.n8629 0.019716
R50505 PAD.n8630 PAD.n2915 0.019716
R50506 PAD.n8621 PAD.n8620 0.019716
R50507 PAD.n8620 PAD.n2914 0.019716
R50508 PAD.n8618 PAD.n8617 0.019716
R50509 PAD.n8618 PAD.n2913 0.019716
R50510 PAD.n8609 PAD.n8608 0.019716
R50511 PAD.n8608 PAD.n2912 0.019716
R50512 PAD.n8606 PAD.n8605 0.019716
R50513 PAD.n8606 PAD.n2911 0.019716
R50514 PAD.n8597 PAD.n8596 0.019716
R50515 PAD.n8596 PAD.n2910 0.019716
R50516 PAD.n8594 PAD.n8593 0.019716
R50517 PAD.n8594 PAD.n2909 0.019716
R50518 PAD.n8585 PAD.n8584 0.019716
R50519 PAD.n8584 PAD.n2908 0.019716
R50520 PAD.n8582 PAD.n8581 0.019716
R50521 PAD.n8582 PAD.n2907 0.019716
R50522 PAD.n8573 PAD.n8572 0.019716
R50523 PAD.n8572 PAD.n2906 0.019716
R50524 PAD.n8570 PAD.n2905 0.019716
R50525 PAD.n3038 PAD.n2994 0.019716
R50526 PAD.n3039 PAD.n2993 0.019716
R50527 PAD.n3048 PAD.n2992 0.019716
R50528 PAD.n3048 PAD.n3047 0.019716
R50529 PAD.n3050 PAD.n2991 0.019716
R50530 PAD.n3051 PAD.n3050 0.019716
R50531 PAD.n3060 PAD.n2990 0.019716
R50532 PAD.n3060 PAD.n3059 0.019716
R50533 PAD.n3062 PAD.n2989 0.019716
R50534 PAD.n3063 PAD.n3062 0.019716
R50535 PAD.n3072 PAD.n2988 0.019716
R50536 PAD.n3072 PAD.n3071 0.019716
R50537 PAD.n3074 PAD.n2987 0.019716
R50538 PAD.n3075 PAD.n3074 0.019716
R50539 PAD.n3084 PAD.n2986 0.019716
R50540 PAD.n3084 PAD.n3083 0.019716
R50541 PAD.n3086 PAD.n2985 0.019716
R50542 PAD.n3087 PAD.n3086 0.019716
R50543 PAD.n3096 PAD.n2984 0.019716
R50544 PAD.n3096 PAD.n3095 0.019716
R50545 PAD.n3098 PAD.n2983 0.019716
R50546 PAD.n3099 PAD.n3098 0.019716
R50547 PAD.n3108 PAD.n2982 0.019716
R50548 PAD.n3108 PAD.n3107 0.019716
R50549 PAD.n3110 PAD.n2981 0.019716
R50550 PAD.n3111 PAD.n3110 0.019716
R50551 PAD.n3120 PAD.n2980 0.019716
R50552 PAD.n3120 PAD.n3119 0.019716
R50553 PAD.n3122 PAD.n2979 0.019716
R50554 PAD.n3123 PAD.n3122 0.019716
R50555 PAD.n3132 PAD.n2978 0.019716
R50556 PAD.n3132 PAD.n3131 0.019716
R50557 PAD.n3134 PAD.n2977 0.019716
R50558 PAD.n3135 PAD.n3134 0.019716
R50559 PAD.n3144 PAD.n2976 0.019716
R50560 PAD.n3144 PAD.n3143 0.019716
R50561 PAD.n3146 PAD.n2975 0.019716
R50562 PAD.n3147 PAD.n3146 0.019716
R50563 PAD.n3156 PAD.n2974 0.019716
R50564 PAD.n3156 PAD.n3155 0.019716
R50565 PAD.n3158 PAD.n2973 0.019716
R50566 PAD.n3159 PAD.n3158 0.019716
R50567 PAD.n3168 PAD.n2972 0.019716
R50568 PAD.n3168 PAD.n3167 0.019716
R50569 PAD.n3170 PAD.n2971 0.019716
R50570 PAD.n3171 PAD.n3170 0.019716
R50571 PAD.n3180 PAD.n2970 0.019716
R50572 PAD.n3180 PAD.n3179 0.019716
R50573 PAD.n3182 PAD.n2969 0.019716
R50574 PAD.n3183 PAD.n3182 0.019716
R50575 PAD.n3192 PAD.n2968 0.019716
R50576 PAD.n3192 PAD.n3191 0.019716
R50577 PAD.n3194 PAD.n2967 0.019716
R50578 PAD.n3195 PAD.n3194 0.019716
R50579 PAD.n3204 PAD.n2966 0.019716
R50580 PAD.n3204 PAD.n3203 0.019716
R50581 PAD.n3206 PAD.n2965 0.019716
R50582 PAD.n3207 PAD.n3206 0.019716
R50583 PAD.n3216 PAD.n2964 0.019716
R50584 PAD.n3216 PAD.n3215 0.019716
R50585 PAD.n3218 PAD.n2963 0.019716
R50586 PAD.n3219 PAD.n3218 0.019716
R50587 PAD.n3228 PAD.n2962 0.019716
R50588 PAD.n3228 PAD.n3227 0.019716
R50589 PAD.n3230 PAD.n2961 0.019716
R50590 PAD.n3231 PAD.n3230 0.019716
R50591 PAD.n3240 PAD.n2960 0.019716
R50592 PAD.n3240 PAD.n3239 0.019716
R50593 PAD.n3242 PAD.n2959 0.019716
R50594 PAD.n3243 PAD.n3242 0.019716
R50595 PAD.n3252 PAD.n2958 0.019716
R50596 PAD.n3252 PAD.n3251 0.019716
R50597 PAD.n3254 PAD.n2957 0.019716
R50598 PAD.n3255 PAD.n3254 0.019716
R50599 PAD.n3264 PAD.n2956 0.019716
R50600 PAD.n3264 PAD.n3263 0.019716
R50601 PAD.n3266 PAD.n2955 0.019716
R50602 PAD.n3267 PAD.n3266 0.019716
R50603 PAD.n3276 PAD.n2954 0.019716
R50604 PAD.n3276 PAD.n3275 0.019716
R50605 PAD.n3278 PAD.n2953 0.019716
R50606 PAD.n3279 PAD.n3278 0.019716
R50607 PAD.n8516 PAD.n8515 0.019716
R50608 PAD.n3383 PAD.n3338 0.019716
R50609 PAD.n3384 PAD.n3337 0.019716
R50610 PAD.n3393 PAD.n3336 0.019716
R50611 PAD.n3393 PAD.n3392 0.019716
R50612 PAD.n3395 PAD.n3335 0.019716
R50613 PAD.n3396 PAD.n3395 0.019716
R50614 PAD.n3405 PAD.n3334 0.019716
R50615 PAD.n3405 PAD.n3404 0.019716
R50616 PAD.n3407 PAD.n3333 0.019716
R50617 PAD.n3408 PAD.n3407 0.019716
R50618 PAD.n3417 PAD.n3332 0.019716
R50619 PAD.n3417 PAD.n3416 0.019716
R50620 PAD.n3419 PAD.n3331 0.019716
R50621 PAD.n3420 PAD.n3419 0.019716
R50622 PAD.n3429 PAD.n3330 0.019716
R50623 PAD.n3429 PAD.n3428 0.019716
R50624 PAD.n3431 PAD.n3329 0.019716
R50625 PAD.n3432 PAD.n3431 0.019716
R50626 PAD.n3441 PAD.n3328 0.019716
R50627 PAD.n3441 PAD.n3440 0.019716
R50628 PAD.n3443 PAD.n3327 0.019716
R50629 PAD.n3444 PAD.n3443 0.019716
R50630 PAD.n3453 PAD.n3326 0.019716
R50631 PAD.n3453 PAD.n3452 0.019716
R50632 PAD.n3455 PAD.n3325 0.019716
R50633 PAD.n3456 PAD.n3455 0.019716
R50634 PAD.n3465 PAD.n3324 0.019716
R50635 PAD.n3465 PAD.n3464 0.019716
R50636 PAD.n3467 PAD.n3323 0.019716
R50637 PAD.n3468 PAD.n3467 0.019716
R50638 PAD.n3477 PAD.n3322 0.019716
R50639 PAD.n3477 PAD.n3476 0.019716
R50640 PAD.n3479 PAD.n3321 0.019716
R50641 PAD.n3480 PAD.n3479 0.019716
R50642 PAD.n3489 PAD.n3320 0.019716
R50643 PAD.n3489 PAD.n3488 0.019716
R50644 PAD.n3491 PAD.n3319 0.019716
R50645 PAD.n3492 PAD.n3491 0.019716
R50646 PAD.n3501 PAD.n3318 0.019716
R50647 PAD.n3501 PAD.n3500 0.019716
R50648 PAD.n3503 PAD.n3317 0.019716
R50649 PAD.n3504 PAD.n3503 0.019716
R50650 PAD.n3513 PAD.n3316 0.019716
R50651 PAD.n3513 PAD.n3512 0.019716
R50652 PAD.n3515 PAD.n3315 0.019716
R50653 PAD.n3516 PAD.n3515 0.019716
R50654 PAD.n3525 PAD.n3314 0.019716
R50655 PAD.n3525 PAD.n3524 0.019716
R50656 PAD.n3527 PAD.n3313 0.019716
R50657 PAD.n3528 PAD.n3527 0.019716
R50658 PAD.n3537 PAD.n3312 0.019716
R50659 PAD.n3537 PAD.n3536 0.019716
R50660 PAD.n3539 PAD.n3311 0.019716
R50661 PAD.n3540 PAD.n3539 0.019716
R50662 PAD.n3549 PAD.n3310 0.019716
R50663 PAD.n3549 PAD.n3548 0.019716
R50664 PAD.n3551 PAD.n3309 0.019716
R50665 PAD.n3552 PAD.n3551 0.019716
R50666 PAD.n3561 PAD.n3308 0.019716
R50667 PAD.n3561 PAD.n3560 0.019716
R50668 PAD.n3563 PAD.n3307 0.019716
R50669 PAD.n3564 PAD.n3563 0.019716
R50670 PAD.n3573 PAD.n3306 0.019716
R50671 PAD.n3573 PAD.n3572 0.019716
R50672 PAD.n3575 PAD.n3305 0.019716
R50673 PAD.n3576 PAD.n3575 0.019716
R50674 PAD.n3585 PAD.n3304 0.019716
R50675 PAD.n3585 PAD.n3584 0.019716
R50676 PAD.n3587 PAD.n3303 0.019716
R50677 PAD.n3588 PAD.n3587 0.019716
R50678 PAD.n3597 PAD.n3302 0.019716
R50679 PAD.n3597 PAD.n3596 0.019716
R50680 PAD.n3599 PAD.n3301 0.019716
R50681 PAD.n3600 PAD.n3599 0.019716
R50682 PAD.n3609 PAD.n3300 0.019716
R50683 PAD.n3609 PAD.n3608 0.019716
R50684 PAD.n3611 PAD.n3299 0.019716
R50685 PAD.n3612 PAD.n3611 0.019716
R50686 PAD.n3621 PAD.n3298 0.019716
R50687 PAD.n3621 PAD.n3620 0.019716
R50688 PAD.n3623 PAD.n3297 0.019716
R50689 PAD.n3624 PAD.n3623 0.019716
R50690 PAD.n8491 PAD.n8490 0.019716
R50691 PAD.n3728 PAD.n3683 0.019716
R50692 PAD.n3729 PAD.n3682 0.019716
R50693 PAD.n3738 PAD.n3681 0.019716
R50694 PAD.n3738 PAD.n3737 0.019716
R50695 PAD.n3740 PAD.n3680 0.019716
R50696 PAD.n3741 PAD.n3740 0.019716
R50697 PAD.n3750 PAD.n3679 0.019716
R50698 PAD.n3750 PAD.n3749 0.019716
R50699 PAD.n3752 PAD.n3678 0.019716
R50700 PAD.n3753 PAD.n3752 0.019716
R50701 PAD.n3762 PAD.n3677 0.019716
R50702 PAD.n3762 PAD.n3761 0.019716
R50703 PAD.n3764 PAD.n3676 0.019716
R50704 PAD.n3765 PAD.n3764 0.019716
R50705 PAD.n3774 PAD.n3675 0.019716
R50706 PAD.n3774 PAD.n3773 0.019716
R50707 PAD.n3776 PAD.n3674 0.019716
R50708 PAD.n3777 PAD.n3776 0.019716
R50709 PAD.n3786 PAD.n3673 0.019716
R50710 PAD.n3786 PAD.n3785 0.019716
R50711 PAD.n3788 PAD.n3672 0.019716
R50712 PAD.n3789 PAD.n3788 0.019716
R50713 PAD.n3798 PAD.n3671 0.019716
R50714 PAD.n3798 PAD.n3797 0.019716
R50715 PAD.n3800 PAD.n3670 0.019716
R50716 PAD.n3801 PAD.n3800 0.019716
R50717 PAD.n3810 PAD.n3669 0.019716
R50718 PAD.n3810 PAD.n3809 0.019716
R50719 PAD.n3812 PAD.n3668 0.019716
R50720 PAD.n3813 PAD.n3812 0.019716
R50721 PAD.n3822 PAD.n3667 0.019716
R50722 PAD.n3822 PAD.n3821 0.019716
R50723 PAD.n3824 PAD.n3666 0.019716
R50724 PAD.n3825 PAD.n3824 0.019716
R50725 PAD.n3834 PAD.n3665 0.019716
R50726 PAD.n3834 PAD.n3833 0.019716
R50727 PAD.n3836 PAD.n3664 0.019716
R50728 PAD.n3837 PAD.n3836 0.019716
R50729 PAD.n3846 PAD.n3663 0.019716
R50730 PAD.n3846 PAD.n3845 0.019716
R50731 PAD.n3848 PAD.n3662 0.019716
R50732 PAD.n3849 PAD.n3848 0.019716
R50733 PAD.n3858 PAD.n3661 0.019716
R50734 PAD.n3858 PAD.n3857 0.019716
R50735 PAD.n3860 PAD.n3660 0.019716
R50736 PAD.n3861 PAD.n3860 0.019716
R50737 PAD.n3870 PAD.n3659 0.019716
R50738 PAD.n3870 PAD.n3869 0.019716
R50739 PAD.n3872 PAD.n3658 0.019716
R50740 PAD.n3873 PAD.n3872 0.019716
R50741 PAD.n3882 PAD.n3657 0.019716
R50742 PAD.n3882 PAD.n3881 0.019716
R50743 PAD.n3884 PAD.n3656 0.019716
R50744 PAD.n3885 PAD.n3884 0.019716
R50745 PAD.n3894 PAD.n3655 0.019716
R50746 PAD.n3894 PAD.n3893 0.019716
R50747 PAD.n3896 PAD.n3654 0.019716
R50748 PAD.n3897 PAD.n3896 0.019716
R50749 PAD.n3906 PAD.n3653 0.019716
R50750 PAD.n3906 PAD.n3905 0.019716
R50751 PAD.n3908 PAD.n3652 0.019716
R50752 PAD.n3909 PAD.n3908 0.019716
R50753 PAD.n3918 PAD.n3651 0.019716
R50754 PAD.n3918 PAD.n3917 0.019716
R50755 PAD.n3920 PAD.n3650 0.019716
R50756 PAD.n3921 PAD.n3920 0.019716
R50757 PAD.n3930 PAD.n3649 0.019716
R50758 PAD.n3930 PAD.n3929 0.019716
R50759 PAD.n3932 PAD.n3648 0.019716
R50760 PAD.n3933 PAD.n3932 0.019716
R50761 PAD.n3942 PAD.n3647 0.019716
R50762 PAD.n3942 PAD.n3941 0.019716
R50763 PAD.n3944 PAD.n3646 0.019716
R50764 PAD.n3945 PAD.n3944 0.019716
R50765 PAD.n3954 PAD.n3645 0.019716
R50766 PAD.n3954 PAD.n3953 0.019716
R50767 PAD.n3956 PAD.n3644 0.019716
R50768 PAD.n3957 PAD.n3956 0.019716
R50769 PAD.n3966 PAD.n3643 0.019716
R50770 PAD.n3966 PAD.n3965 0.019716
R50771 PAD.n3968 PAD.n3642 0.019716
R50772 PAD.n3969 PAD.n3968 0.019716
R50773 PAD.n8467 PAD.n8466 0.019716
R50774 PAD.n4069 PAD.n4025 0.019716
R50775 PAD.n4070 PAD.n4024 0.019716
R50776 PAD.n4079 PAD.n4023 0.019716
R50777 PAD.n4079 PAD.n4078 0.019716
R50778 PAD.n4081 PAD.n4022 0.019716
R50779 PAD.n4082 PAD.n4081 0.019716
R50780 PAD.n4091 PAD.n4021 0.019716
R50781 PAD.n4091 PAD.n4090 0.019716
R50782 PAD.n4093 PAD.n4020 0.019716
R50783 PAD.n4094 PAD.n4093 0.019716
R50784 PAD.n4103 PAD.n4019 0.019716
R50785 PAD.n4103 PAD.n4102 0.019716
R50786 PAD.n4105 PAD.n4018 0.019716
R50787 PAD.n4106 PAD.n4105 0.019716
R50788 PAD.n4115 PAD.n4017 0.019716
R50789 PAD.n4115 PAD.n4114 0.019716
R50790 PAD.n4117 PAD.n4016 0.019716
R50791 PAD.n4118 PAD.n4117 0.019716
R50792 PAD.n4127 PAD.n4015 0.019716
R50793 PAD.n4127 PAD.n4126 0.019716
R50794 PAD.n4129 PAD.n4014 0.019716
R50795 PAD.n4130 PAD.n4129 0.019716
R50796 PAD.n4139 PAD.n4013 0.019716
R50797 PAD.n4139 PAD.n4138 0.019716
R50798 PAD.n4141 PAD.n4012 0.019716
R50799 PAD.n4142 PAD.n4141 0.019716
R50800 PAD.n4151 PAD.n4011 0.019716
R50801 PAD.n4151 PAD.n4150 0.019716
R50802 PAD.n4153 PAD.n4010 0.019716
R50803 PAD.n4154 PAD.n4153 0.019716
R50804 PAD.n4163 PAD.n4009 0.019716
R50805 PAD.n4163 PAD.n4162 0.019716
R50806 PAD.n4165 PAD.n4008 0.019716
R50807 PAD.n4166 PAD.n4165 0.019716
R50808 PAD.n4175 PAD.n4007 0.019716
R50809 PAD.n4175 PAD.n4174 0.019716
R50810 PAD.n4177 PAD.n4006 0.019716
R50811 PAD.n4178 PAD.n4177 0.019716
R50812 PAD.n4187 PAD.n4005 0.019716
R50813 PAD.n4187 PAD.n4186 0.019716
R50814 PAD.n4189 PAD.n4004 0.019716
R50815 PAD.n4190 PAD.n4189 0.019716
R50816 PAD.n4199 PAD.n4003 0.019716
R50817 PAD.n4199 PAD.n4198 0.019716
R50818 PAD.n4201 PAD.n4002 0.019716
R50819 PAD.n4202 PAD.n4201 0.019716
R50820 PAD.n4211 PAD.n4001 0.019716
R50821 PAD.n4211 PAD.n4210 0.019716
R50822 PAD.n4213 PAD.n4000 0.019716
R50823 PAD.n4214 PAD.n4213 0.019716
R50824 PAD.n4223 PAD.n3999 0.019716
R50825 PAD.n4223 PAD.n4222 0.019716
R50826 PAD.n4225 PAD.n3998 0.019716
R50827 PAD.n4226 PAD.n4225 0.019716
R50828 PAD.n4235 PAD.n3997 0.019716
R50829 PAD.n4235 PAD.n4234 0.019716
R50830 PAD.n4237 PAD.n3996 0.019716
R50831 PAD.n4238 PAD.n4237 0.019716
R50832 PAD.n4247 PAD.n3995 0.019716
R50833 PAD.n4247 PAD.n4246 0.019716
R50834 PAD.n4249 PAD.n3994 0.019716
R50835 PAD.n4250 PAD.n4249 0.019716
R50836 PAD.n4259 PAD.n3993 0.019716
R50837 PAD.n4259 PAD.n4258 0.019716
R50838 PAD.n4261 PAD.n3992 0.019716
R50839 PAD.n4262 PAD.n4261 0.019716
R50840 PAD.n4271 PAD.n3991 0.019716
R50841 PAD.n4271 PAD.n4270 0.019716
R50842 PAD.n4273 PAD.n3990 0.019716
R50843 PAD.n4274 PAD.n4273 0.019716
R50844 PAD.n4283 PAD.n3989 0.019716
R50845 PAD.n4283 PAD.n4282 0.019716
R50846 PAD.n4285 PAD.n3988 0.019716
R50847 PAD.n4286 PAD.n4285 0.019716
R50848 PAD.n4295 PAD.n3987 0.019716
R50849 PAD.n4295 PAD.n4294 0.019716
R50850 PAD.n4297 PAD.n3986 0.019716
R50851 PAD.n4298 PAD.n4297 0.019716
R50852 PAD.n4307 PAD.n3985 0.019716
R50853 PAD.n4307 PAD.n4306 0.019716
R50854 PAD.n4309 PAD.n3984 0.019716
R50855 PAD.n4310 PAD.n4309 0.019716
R50856 PAD.n8443 PAD.n8442 0.019716
R50857 PAD.n4421 PAD.n4420 0.019716
R50858 PAD.n4423 PAD.n4422 0.019716
R50859 PAD.n4424 PAD.n4415 0.019716
R50860 PAD.n4425 PAD.n4424 0.019716
R50861 PAD.n4435 PAD.n4434 0.019716
R50862 PAD.n4434 PAD.n4433 0.019716
R50863 PAD.n4436 PAD.n4411 0.019716
R50864 PAD.n4437 PAD.n4436 0.019716
R50865 PAD.n4447 PAD.n4446 0.019716
R50866 PAD.n4446 PAD.n4445 0.019716
R50867 PAD.n4448 PAD.n4407 0.019716
R50868 PAD.n4449 PAD.n4448 0.019716
R50869 PAD.n4459 PAD.n4458 0.019716
R50870 PAD.n4458 PAD.n4457 0.019716
R50871 PAD.n4460 PAD.n4403 0.019716
R50872 PAD.n4461 PAD.n4460 0.019716
R50873 PAD.n4471 PAD.n4470 0.019716
R50874 PAD.n4470 PAD.n4469 0.019716
R50875 PAD.n4472 PAD.n4399 0.019716
R50876 PAD.n4473 PAD.n4472 0.019716
R50877 PAD.n4483 PAD.n4482 0.019716
R50878 PAD.n4482 PAD.n4481 0.019716
R50879 PAD.n4484 PAD.n4395 0.019716
R50880 PAD.n4485 PAD.n4484 0.019716
R50881 PAD.n4495 PAD.n4494 0.019716
R50882 PAD.n4494 PAD.n4493 0.019716
R50883 PAD.n4496 PAD.n4391 0.019716
R50884 PAD.n4497 PAD.n4496 0.019716
R50885 PAD.n4507 PAD.n4506 0.019716
R50886 PAD.n4506 PAD.n4505 0.019716
R50887 PAD.n4508 PAD.n4387 0.019716
R50888 PAD.n4509 PAD.n4508 0.019716
R50889 PAD.n4519 PAD.n4518 0.019716
R50890 PAD.n4518 PAD.n4517 0.019716
R50891 PAD.n4520 PAD.n4383 0.019716
R50892 PAD.n4521 PAD.n4520 0.019716
R50893 PAD.n4531 PAD.n4530 0.019716
R50894 PAD.n4530 PAD.n4529 0.019716
R50895 PAD.n4532 PAD.n4379 0.019716
R50896 PAD.n4533 PAD.n4532 0.019716
R50897 PAD.n4543 PAD.n4542 0.019716
R50898 PAD.n4542 PAD.n4541 0.019716
R50899 PAD.n4544 PAD.n4375 0.019716
R50900 PAD.n4545 PAD.n4544 0.019716
R50901 PAD.n4555 PAD.n4554 0.019716
R50902 PAD.n4554 PAD.n4553 0.019716
R50903 PAD.n4556 PAD.n4371 0.019716
R50904 PAD.n4557 PAD.n4556 0.019716
R50905 PAD.n4567 PAD.n4566 0.019716
R50906 PAD.n4566 PAD.n4565 0.019716
R50907 PAD.n4568 PAD.n4367 0.019716
R50908 PAD.n4569 PAD.n4568 0.019716
R50909 PAD.n4579 PAD.n4578 0.019716
R50910 PAD.n4578 PAD.n4577 0.019716
R50911 PAD.n4580 PAD.n4363 0.019716
R50912 PAD.n4581 PAD.n4580 0.019716
R50913 PAD.n4591 PAD.n4590 0.019716
R50914 PAD.n4590 PAD.n4589 0.019716
R50915 PAD.n4592 PAD.n4359 0.019716
R50916 PAD.n4593 PAD.n4592 0.019716
R50917 PAD.n4603 PAD.n4602 0.019716
R50918 PAD.n4602 PAD.n4601 0.019716
R50919 PAD.n4604 PAD.n4355 0.019716
R50920 PAD.n4605 PAD.n4604 0.019716
R50921 PAD.n4615 PAD.n4614 0.019716
R50922 PAD.n4614 PAD.n4613 0.019716
R50923 PAD.n4616 PAD.n4351 0.019716
R50924 PAD.n4617 PAD.n4616 0.019716
R50925 PAD.n4627 PAD.n4626 0.019716
R50926 PAD.n4626 PAD.n4625 0.019716
R50927 PAD.n4628 PAD.n4347 0.019716
R50928 PAD.n4629 PAD.n4628 0.019716
R50929 PAD.n4639 PAD.n4638 0.019716
R50930 PAD.n4638 PAD.n4637 0.019716
R50931 PAD.n4640 PAD.n4343 0.019716
R50932 PAD.n4641 PAD.n4640 0.019716
R50933 PAD.n4651 PAD.n4650 0.019716
R50934 PAD.n4650 PAD.n4649 0.019716
R50935 PAD.n4652 PAD.n4339 0.019716
R50936 PAD.n4653 PAD.n4652 0.019716
R50937 PAD.n4664 PAD.n4663 0.019716
R50938 PAD.n4663 PAD.n4662 0.019716
R50939 PAD.n4667 PAD.n4666 0.019716
R50940 PAD.n8396 PAD.n8395 0.019716
R50941 PAD.n4726 PAD.n4725 0.019716
R50942 PAD.n8388 PAD.n8387 0.019716
R50943 PAD.n8388 PAD.n4723 0.019716
R50944 PAD.n4733 PAD.n4732 0.019716
R50945 PAD.n4733 PAD.n4722 0.019716
R50946 PAD.n8379 PAD.n8378 0.019716
R50947 PAD.n8379 PAD.n4721 0.019716
R50948 PAD.n4738 PAD.n4737 0.019716
R50949 PAD.n4738 PAD.n4720 0.019716
R50950 PAD.n8370 PAD.n8369 0.019716
R50951 PAD.n8370 PAD.n4719 0.019716
R50952 PAD.n4743 PAD.n4742 0.019716
R50953 PAD.n4743 PAD.n4718 0.019716
R50954 PAD.n8361 PAD.n8360 0.019716
R50955 PAD.n8361 PAD.n4717 0.019716
R50956 PAD.n4748 PAD.n4747 0.019716
R50957 PAD.n4748 PAD.n4716 0.019716
R50958 PAD.n8352 PAD.n8351 0.019716
R50959 PAD.n8352 PAD.n4715 0.019716
R50960 PAD.n4753 PAD.n4752 0.019716
R50961 PAD.n4753 PAD.n4714 0.019716
R50962 PAD.n8343 PAD.n8342 0.019716
R50963 PAD.n8343 PAD.n4713 0.019716
R50964 PAD.n4758 PAD.n4757 0.019716
R50965 PAD.n4758 PAD.n4712 0.019716
R50966 PAD.n8334 PAD.n8333 0.019716
R50967 PAD.n8334 PAD.n4711 0.019716
R50968 PAD.n4763 PAD.n4762 0.019716
R50969 PAD.n4763 PAD.n4710 0.019716
R50970 PAD.n8325 PAD.n8324 0.019716
R50971 PAD.n8325 PAD.n4709 0.019716
R50972 PAD.n4768 PAD.n4767 0.019716
R50973 PAD.n4768 PAD.n4708 0.019716
R50974 PAD.n8316 PAD.n8315 0.019716
R50975 PAD.n8316 PAD.n4707 0.019716
R50976 PAD.n4773 PAD.n4772 0.019716
R50977 PAD.n4773 PAD.n4706 0.019716
R50978 PAD.n8307 PAD.n8306 0.019716
R50979 PAD.n8307 PAD.n4705 0.019716
R50980 PAD.n4778 PAD.n4777 0.019716
R50981 PAD.n4778 PAD.n4704 0.019716
R50982 PAD.n8298 PAD.n8297 0.019716
R50983 PAD.n8298 PAD.n4703 0.019716
R50984 PAD.n4783 PAD.n4782 0.019716
R50985 PAD.n4783 PAD.n4702 0.019716
R50986 PAD.n8289 PAD.n8288 0.019716
R50987 PAD.n8289 PAD.n4701 0.019716
R50988 PAD.n4788 PAD.n4787 0.019716
R50989 PAD.n4788 PAD.n4700 0.019716
R50990 PAD.n8280 PAD.n8279 0.019716
R50991 PAD.n8280 PAD.n4699 0.019716
R50992 PAD.n4793 PAD.n4792 0.019716
R50993 PAD.n4793 PAD.n4698 0.019716
R50994 PAD.n8271 PAD.n8270 0.019716
R50995 PAD.n8271 PAD.n4697 0.019716
R50996 PAD.n4798 PAD.n4797 0.019716
R50997 PAD.n4798 PAD.n4696 0.019716
R50998 PAD.n8262 PAD.n8261 0.019716
R50999 PAD.n8262 PAD.n4695 0.019716
R51000 PAD.n4803 PAD.n4802 0.019716
R51001 PAD.n4803 PAD.n4694 0.019716
R51002 PAD.n8253 PAD.n8252 0.019716
R51003 PAD.n8253 PAD.n4693 0.019716
R51004 PAD.n4808 PAD.n4807 0.019716
R51005 PAD.n4808 PAD.n4692 0.019716
R51006 PAD.n8244 PAD.n8243 0.019716
R51007 PAD.n8244 PAD.n4691 0.019716
R51008 PAD.n4813 PAD.n4812 0.019716
R51009 PAD.n4813 PAD.n4690 0.019716
R51010 PAD.n8235 PAD.n8234 0.019716
R51011 PAD.n8235 PAD.n4689 0.019716
R51012 PAD.n4818 PAD.n4817 0.019716
R51013 PAD.n4818 PAD.n4688 0.019716
R51014 PAD.n8226 PAD.n8225 0.019716
R51015 PAD.n8226 PAD.n4687 0.019716
R51016 PAD.n4823 PAD.n4822 0.019716
R51017 PAD.n4823 PAD.n4686 0.019716
R51018 PAD.n8217 PAD.n8216 0.019716
R51019 PAD.n8217 PAD.n4685 0.019716
R51020 PAD.n4828 PAD.n4827 0.019716
R51021 PAD.n4828 PAD.n4684 0.019716
R51022 PAD.n4832 PAD.n4683 0.019716
R51023 PAD.n4849 PAD.n4847 0.019716
R51024 PAD.n5176 PAD.n5175 0.019716
R51025 PAD.n5172 PAD.n4850 0.019716
R51026 PAD.n5173 PAD.n5172 0.019716
R51027 PAD.n5166 PAD.n5163 0.019716
R51028 PAD.n5166 PAD.n5165 0.019716
R51029 PAD.n5160 PAD.n4855 0.019716
R51030 PAD.n5161 PAD.n5160 0.019716
R51031 PAD.n5154 PAD.n5151 0.019716
R51032 PAD.n5154 PAD.n5153 0.019716
R51033 PAD.n5148 PAD.n4859 0.019716
R51034 PAD.n5149 PAD.n5148 0.019716
R51035 PAD.n5142 PAD.n5139 0.019716
R51036 PAD.n5142 PAD.n5141 0.019716
R51037 PAD.n5136 PAD.n4863 0.019716
R51038 PAD.n5137 PAD.n5136 0.019716
R51039 PAD.n5130 PAD.n5127 0.019716
R51040 PAD.n5130 PAD.n5129 0.019716
R51041 PAD.n5124 PAD.n4867 0.019716
R51042 PAD.n5125 PAD.n5124 0.019716
R51043 PAD.n5118 PAD.n5115 0.019716
R51044 PAD.n5118 PAD.n5117 0.019716
R51045 PAD.n5112 PAD.n4871 0.019716
R51046 PAD.n5113 PAD.n5112 0.019716
R51047 PAD.n5106 PAD.n5103 0.019716
R51048 PAD.n5106 PAD.n5105 0.019716
R51049 PAD.n5100 PAD.n4875 0.019716
R51050 PAD.n5101 PAD.n5100 0.019716
R51051 PAD.n5094 PAD.n5091 0.019716
R51052 PAD.n5094 PAD.n5093 0.019716
R51053 PAD.n5088 PAD.n4879 0.019716
R51054 PAD.n5089 PAD.n5088 0.019716
R51055 PAD.n5082 PAD.n5079 0.019716
R51056 PAD.n5082 PAD.n5081 0.019716
R51057 PAD.n5076 PAD.n4883 0.019716
R51058 PAD.n5077 PAD.n5076 0.019716
R51059 PAD.n5070 PAD.n5067 0.019716
R51060 PAD.n5070 PAD.n5069 0.019716
R51061 PAD.n5064 PAD.n4887 0.019716
R51062 PAD.n5065 PAD.n5064 0.019716
R51063 PAD.n5058 PAD.n5055 0.019716
R51064 PAD.n5058 PAD.n5057 0.019716
R51065 PAD.n5052 PAD.n4891 0.019716
R51066 PAD.n5053 PAD.n5052 0.019716
R51067 PAD.n5046 PAD.n5043 0.019716
R51068 PAD.n5046 PAD.n5045 0.019716
R51069 PAD.n5040 PAD.n4895 0.019716
R51070 PAD.n5041 PAD.n5040 0.019716
R51071 PAD.n5034 PAD.n5031 0.019716
R51072 PAD.n5034 PAD.n5033 0.019716
R51073 PAD.n5028 PAD.n4899 0.019716
R51074 PAD.n5029 PAD.n5028 0.019716
R51075 PAD.n5022 PAD.n5019 0.019716
R51076 PAD.n5022 PAD.n5021 0.019716
R51077 PAD.n5016 PAD.n4903 0.019716
R51078 PAD.n5017 PAD.n5016 0.019716
R51079 PAD.n5010 PAD.n5007 0.019716
R51080 PAD.n5010 PAD.n5009 0.019716
R51081 PAD.n5004 PAD.n4907 0.019716
R51082 PAD.n5005 PAD.n5004 0.019716
R51083 PAD.n4998 PAD.n4995 0.019716
R51084 PAD.n4998 PAD.n4997 0.019716
R51085 PAD.n4992 PAD.n4911 0.019716
R51086 PAD.n4993 PAD.n4992 0.019716
R51087 PAD.n4986 PAD.n4983 0.019716
R51088 PAD.n4986 PAD.n4985 0.019716
R51089 PAD.n4980 PAD.n4915 0.019716
R51090 PAD.n4981 PAD.n4980 0.019716
R51091 PAD.n4974 PAD.n4971 0.019716
R51092 PAD.n4974 PAD.n4973 0.019716
R51093 PAD.n4968 PAD.n4919 0.019716
R51094 PAD.n4969 PAD.n4968 0.019716
R51095 PAD.n4962 PAD.n4959 0.019716
R51096 PAD.n4962 PAD.n4961 0.019716
R51097 PAD.n4956 PAD.n4923 0.019716
R51098 PAD.n4957 PAD.n4956 0.019716
R51099 PAD.n4950 PAD.n4947 0.019716
R51100 PAD.n4950 PAD.n4949 0.019716
R51101 PAD.n4944 PAD.n4927 0.019716
R51102 PAD.n4945 PAD.n4944 0.019716
R51103 PAD.n4938 PAD.n4935 0.019716
R51104 PAD.n4938 PAD.n4937 0.019716
R51105 PAD.n4933 PAD.n4932 0.019716
R51106 PAD.n8162 PAD.n8161 0.019716
R51107 PAD.n7872 PAD.n7871 0.019716
R51108 PAD.n8154 PAD.n8153 0.019716
R51109 PAD.n8154 PAD.n7870 0.019716
R51110 PAD.n7879 PAD.n7878 0.019716
R51111 PAD.n7879 PAD.n7869 0.019716
R51112 PAD.n8145 PAD.n8144 0.019716
R51113 PAD.n8145 PAD.n7868 0.019716
R51114 PAD.n7884 PAD.n7883 0.019716
R51115 PAD.n7884 PAD.n7867 0.019716
R51116 PAD.n8136 PAD.n8135 0.019716
R51117 PAD.n8136 PAD.n7866 0.019716
R51118 PAD.n7889 PAD.n7888 0.019716
R51119 PAD.n7889 PAD.n7865 0.019716
R51120 PAD.n8127 PAD.n8126 0.019716
R51121 PAD.n8127 PAD.n7864 0.019716
R51122 PAD.n7894 PAD.n7893 0.019716
R51123 PAD.n7894 PAD.n7863 0.019716
R51124 PAD.n8118 PAD.n8117 0.019716
R51125 PAD.n8118 PAD.n7862 0.019716
R51126 PAD.n7899 PAD.n7898 0.019716
R51127 PAD.n7899 PAD.n7861 0.019716
R51128 PAD.n8109 PAD.n8108 0.019716
R51129 PAD.n8109 PAD.n7860 0.019716
R51130 PAD.n7904 PAD.n7903 0.019716
R51131 PAD.n7904 PAD.n7859 0.019716
R51132 PAD.n8100 PAD.n8099 0.019716
R51133 PAD.n8100 PAD.n7858 0.019716
R51134 PAD.n7909 PAD.n7908 0.019716
R51135 PAD.n7909 PAD.n7857 0.019716
R51136 PAD.n8091 PAD.n8090 0.019716
R51137 PAD.n8091 PAD.n7856 0.019716
R51138 PAD.n7914 PAD.n7913 0.019716
R51139 PAD.n7914 PAD.n7855 0.019716
R51140 PAD.n8082 PAD.n8081 0.019716
R51141 PAD.n8082 PAD.n7854 0.019716
R51142 PAD.n7919 PAD.n7918 0.019716
R51143 PAD.n7919 PAD.n7853 0.019716
R51144 PAD.n8073 PAD.n8072 0.019716
R51145 PAD.n8073 PAD.n7852 0.019716
R51146 PAD.n7924 PAD.n7923 0.019716
R51147 PAD.n7924 PAD.n7851 0.019716
R51148 PAD.n8064 PAD.n8063 0.019716
R51149 PAD.n8064 PAD.n7850 0.019716
R51150 PAD.n7929 PAD.n7928 0.019716
R51151 PAD.n7929 PAD.n7849 0.019716
R51152 PAD.n8055 PAD.n8054 0.019716
R51153 PAD.n8055 PAD.n7848 0.019716
R51154 PAD.n7934 PAD.n7933 0.019716
R51155 PAD.n7934 PAD.n7847 0.019716
R51156 PAD.n8046 PAD.n8045 0.019716
R51157 PAD.n8046 PAD.n7846 0.019716
R51158 PAD.n7939 PAD.n7938 0.019716
R51159 PAD.n7939 PAD.n7845 0.019716
R51160 PAD.n8037 PAD.n8036 0.019716
R51161 PAD.n8037 PAD.n7844 0.019716
R51162 PAD.n7944 PAD.n7943 0.019716
R51163 PAD.n7944 PAD.n7843 0.019716
R51164 PAD.n8028 PAD.n8027 0.019716
R51165 PAD.n8028 PAD.n7842 0.019716
R51166 PAD.n7949 PAD.n7948 0.019716
R51167 PAD.n7949 PAD.n7841 0.019716
R51168 PAD.n8019 PAD.n8018 0.019716
R51169 PAD.n8019 PAD.n7840 0.019716
R51170 PAD.n7954 PAD.n7953 0.019716
R51171 PAD.n7954 PAD.n7839 0.019716
R51172 PAD.n8010 PAD.n8009 0.019716
R51173 PAD.n8010 PAD.n7838 0.019716
R51174 PAD.n7959 PAD.n7958 0.019716
R51175 PAD.n7959 PAD.n7837 0.019716
R51176 PAD.n8001 PAD.n8000 0.019716
R51177 PAD.n8001 PAD.n7836 0.019716
R51178 PAD.n7964 PAD.n7963 0.019716
R51179 PAD.n7964 PAD.n7835 0.019716
R51180 PAD.n7992 PAD.n7991 0.019716
R51181 PAD.n7992 PAD.n7834 0.019716
R51182 PAD.n7969 PAD.n7968 0.019716
R51183 PAD.n7969 PAD.n7833 0.019716
R51184 PAD.n7983 PAD.n7982 0.019716
R51185 PAD.n7983 PAD.n7832 0.019716
R51186 PAD.n7976 PAD.n7975 0.019716
R51187 PAD.n7976 PAD.n7831 0.019716
R51188 PAD.n7971 PAD.n7830 0.019716
R51189 PAD.n5213 PAD.n5211 0.019716
R51190 PAD.n5540 PAD.n5539 0.019716
R51191 PAD.n5536 PAD.n5214 0.019716
R51192 PAD.n5537 PAD.n5536 0.019716
R51193 PAD.n5530 PAD.n5527 0.019716
R51194 PAD.n5530 PAD.n5529 0.019716
R51195 PAD.n5524 PAD.n5219 0.019716
R51196 PAD.n5525 PAD.n5524 0.019716
R51197 PAD.n5518 PAD.n5515 0.019716
R51198 PAD.n5518 PAD.n5517 0.019716
R51199 PAD.n5512 PAD.n5223 0.019716
R51200 PAD.n5513 PAD.n5512 0.019716
R51201 PAD.n5506 PAD.n5503 0.019716
R51202 PAD.n5506 PAD.n5505 0.019716
R51203 PAD.n5500 PAD.n5227 0.019716
R51204 PAD.n5501 PAD.n5500 0.019716
R51205 PAD.n5494 PAD.n5491 0.019716
R51206 PAD.n5494 PAD.n5493 0.019716
R51207 PAD.n5488 PAD.n5231 0.019716
R51208 PAD.n5489 PAD.n5488 0.019716
R51209 PAD.n5482 PAD.n5479 0.019716
R51210 PAD.n5482 PAD.n5481 0.019716
R51211 PAD.n5476 PAD.n5235 0.019716
R51212 PAD.n5477 PAD.n5476 0.019716
R51213 PAD.n5470 PAD.n5467 0.019716
R51214 PAD.n5470 PAD.n5469 0.019716
R51215 PAD.n5464 PAD.n5239 0.019716
R51216 PAD.n5465 PAD.n5464 0.019716
R51217 PAD.n5458 PAD.n5455 0.019716
R51218 PAD.n5458 PAD.n5457 0.019716
R51219 PAD.n5452 PAD.n5243 0.019716
R51220 PAD.n5453 PAD.n5452 0.019716
R51221 PAD.n5446 PAD.n5443 0.019716
R51222 PAD.n5446 PAD.n5445 0.019716
R51223 PAD.n5440 PAD.n5247 0.019716
R51224 PAD.n5441 PAD.n5440 0.019716
R51225 PAD.n5434 PAD.n5431 0.019716
R51226 PAD.n5434 PAD.n5433 0.019716
R51227 PAD.n5428 PAD.n5251 0.019716
R51228 PAD.n5429 PAD.n5428 0.019716
R51229 PAD.n5422 PAD.n5419 0.019716
R51230 PAD.n5422 PAD.n5421 0.019716
R51231 PAD.n5416 PAD.n5255 0.019716
R51232 PAD.n5417 PAD.n5416 0.019716
R51233 PAD.n5410 PAD.n5407 0.019716
R51234 PAD.n5410 PAD.n5409 0.019716
R51235 PAD.n5404 PAD.n5259 0.019716
R51236 PAD.n5405 PAD.n5404 0.019716
R51237 PAD.n5398 PAD.n5395 0.019716
R51238 PAD.n5398 PAD.n5397 0.019716
R51239 PAD.n5392 PAD.n5263 0.019716
R51240 PAD.n5393 PAD.n5392 0.019716
R51241 PAD.n5386 PAD.n5383 0.019716
R51242 PAD.n5386 PAD.n5385 0.019716
R51243 PAD.n5380 PAD.n5267 0.019716
R51244 PAD.n5381 PAD.n5380 0.019716
R51245 PAD.n5374 PAD.n5371 0.019716
R51246 PAD.n5374 PAD.n5373 0.019716
R51247 PAD.n5368 PAD.n5271 0.019716
R51248 PAD.n5369 PAD.n5368 0.019716
R51249 PAD.n5362 PAD.n5359 0.019716
R51250 PAD.n5362 PAD.n5361 0.019716
R51251 PAD.n5356 PAD.n5275 0.019716
R51252 PAD.n5357 PAD.n5356 0.019716
R51253 PAD.n5350 PAD.n5347 0.019716
R51254 PAD.n5350 PAD.n5349 0.019716
R51255 PAD.n5344 PAD.n5279 0.019716
R51256 PAD.n5345 PAD.n5344 0.019716
R51257 PAD.n5338 PAD.n5335 0.019716
R51258 PAD.n5338 PAD.n5337 0.019716
R51259 PAD.n5332 PAD.n5283 0.019716
R51260 PAD.n5333 PAD.n5332 0.019716
R51261 PAD.n5326 PAD.n5323 0.019716
R51262 PAD.n5326 PAD.n5325 0.019716
R51263 PAD.n5320 PAD.n5287 0.019716
R51264 PAD.n5321 PAD.n5320 0.019716
R51265 PAD.n5314 PAD.n5311 0.019716
R51266 PAD.n5314 PAD.n5313 0.019716
R51267 PAD.n5308 PAD.n5291 0.019716
R51268 PAD.n5309 PAD.n5308 0.019716
R51269 PAD.n5302 PAD.n5299 0.019716
R51270 PAD.n5302 PAD.n5301 0.019716
R51271 PAD.n5297 PAD.n5296 0.019716
R51272 PAD.n7519 PAD.n7518 0.019716
R51273 PAD.n7511 PAD.n7201 0.019716
R51274 PAD.n7509 PAD.n7508 0.019716
R51275 PAD.n7509 PAD.n7199 0.019716
R51276 PAD.n7500 PAD.n7499 0.019716
R51277 PAD.n7499 PAD.n7198 0.019716
R51278 PAD.n7497 PAD.n7496 0.019716
R51279 PAD.n7497 PAD.n7197 0.019716
R51280 PAD.n7488 PAD.n7487 0.019716
R51281 PAD.n7487 PAD.n7196 0.019716
R51282 PAD.n7485 PAD.n7484 0.019716
R51283 PAD.n7485 PAD.n7195 0.019716
R51284 PAD.n7476 PAD.n7475 0.019716
R51285 PAD.n7475 PAD.n7194 0.019716
R51286 PAD.n7473 PAD.n7472 0.019716
R51287 PAD.n7473 PAD.n7193 0.019716
R51288 PAD.n7464 PAD.n7463 0.019716
R51289 PAD.n7463 PAD.n7192 0.019716
R51290 PAD.n7461 PAD.n7460 0.019716
R51291 PAD.n7461 PAD.n7191 0.019716
R51292 PAD.n7452 PAD.n7451 0.019716
R51293 PAD.n7451 PAD.n7190 0.019716
R51294 PAD.n7449 PAD.n7448 0.019716
R51295 PAD.n7449 PAD.n7189 0.019716
R51296 PAD.n7440 PAD.n7439 0.019716
R51297 PAD.n7439 PAD.n7188 0.019716
R51298 PAD.n7437 PAD.n7436 0.019716
R51299 PAD.n7437 PAD.n7187 0.019716
R51300 PAD.n7428 PAD.n7427 0.019716
R51301 PAD.n7427 PAD.n7186 0.019716
R51302 PAD.n7425 PAD.n7424 0.019716
R51303 PAD.n7425 PAD.n7185 0.019716
R51304 PAD.n7416 PAD.n7415 0.019716
R51305 PAD.n7415 PAD.n7184 0.019716
R51306 PAD.n7413 PAD.n7412 0.019716
R51307 PAD.n7413 PAD.n7183 0.019716
R51308 PAD.n7404 PAD.n7403 0.019716
R51309 PAD.n7403 PAD.n7182 0.019716
R51310 PAD.n7401 PAD.n7400 0.019716
R51311 PAD.n7401 PAD.n7181 0.019716
R51312 PAD.n7392 PAD.n7391 0.019716
R51313 PAD.n7391 PAD.n7180 0.019716
R51314 PAD.n7389 PAD.n7388 0.019716
R51315 PAD.n7389 PAD.n7179 0.019716
R51316 PAD.n7380 PAD.n7379 0.019716
R51317 PAD.n7379 PAD.n7178 0.019716
R51318 PAD.n7377 PAD.n7376 0.019716
R51319 PAD.n7377 PAD.n7177 0.019716
R51320 PAD.n7368 PAD.n7367 0.019716
R51321 PAD.n7367 PAD.n7176 0.019716
R51322 PAD.n7365 PAD.n7364 0.019716
R51323 PAD.n7365 PAD.n7175 0.019716
R51324 PAD.n7356 PAD.n7355 0.019716
R51325 PAD.n7355 PAD.n7174 0.019716
R51326 PAD.n7353 PAD.n7352 0.019716
R51327 PAD.n7353 PAD.n7173 0.019716
R51328 PAD.n7344 PAD.n7343 0.019716
R51329 PAD.n7343 PAD.n7172 0.019716
R51330 PAD.n7341 PAD.n7340 0.019716
R51331 PAD.n7341 PAD.n7171 0.019716
R51332 PAD.n7332 PAD.n7331 0.019716
R51333 PAD.n7331 PAD.n7170 0.019716
R51334 PAD.n7329 PAD.n7328 0.019716
R51335 PAD.n7329 PAD.n7169 0.019716
R51336 PAD.n7320 PAD.n7319 0.019716
R51337 PAD.n7319 PAD.n7168 0.019716
R51338 PAD.n7317 PAD.n7316 0.019716
R51339 PAD.n7317 PAD.n7167 0.019716
R51340 PAD.n7308 PAD.n7307 0.019716
R51341 PAD.n7307 PAD.n7166 0.019716
R51342 PAD.n7305 PAD.n7304 0.019716
R51343 PAD.n7305 PAD.n7165 0.019716
R51344 PAD.n7296 PAD.n7295 0.019716
R51345 PAD.n7295 PAD.n7164 0.019716
R51346 PAD.n7293 PAD.n7292 0.019716
R51347 PAD.n7293 PAD.n7163 0.019716
R51348 PAD.n7284 PAD.n7283 0.019716
R51349 PAD.n7283 PAD.n7162 0.019716
R51350 PAD.n7281 PAD.n7280 0.019716
R51351 PAD.n7281 PAD.n7161 0.019716
R51352 PAD.n7272 PAD.n7271 0.019716
R51353 PAD.n7271 PAD.n7160 0.019716
R51354 PAD.n7269 PAD.n7159 0.019716
R51355 PAD.n7781 PAD.n7780 0.019716
R51356 PAD.n7773 PAD.n7104 0.019716
R51357 PAD.n7771 PAD.n7770 0.019716
R51358 PAD.n7771 PAD.n7102 0.019716
R51359 PAD.n7762 PAD.n7761 0.019716
R51360 PAD.n7761 PAD.n7101 0.019716
R51361 PAD.n7759 PAD.n7758 0.019716
R51362 PAD.n7759 PAD.n7100 0.019716
R51363 PAD.n7750 PAD.n7749 0.019716
R51364 PAD.n7749 PAD.n7099 0.019716
R51365 PAD.n7747 PAD.n7746 0.019716
R51366 PAD.n7747 PAD.n7098 0.019716
R51367 PAD.n7738 PAD.n7737 0.019716
R51368 PAD.n7737 PAD.n7097 0.019716
R51369 PAD.n7735 PAD.n7734 0.019716
R51370 PAD.n7735 PAD.n7096 0.019716
R51371 PAD.n7726 PAD.n7725 0.019716
R51372 PAD.n7725 PAD.n7095 0.019716
R51373 PAD.n7723 PAD.n7722 0.019716
R51374 PAD.n7723 PAD.n7094 0.019716
R51375 PAD.n7714 PAD.n7713 0.019716
R51376 PAD.n7713 PAD.n7093 0.019716
R51377 PAD.n7711 PAD.n7710 0.019716
R51378 PAD.n7711 PAD.n7092 0.019716
R51379 PAD.n7702 PAD.n7701 0.019716
R51380 PAD.n7701 PAD.n7091 0.019716
R51381 PAD.n7699 PAD.n7698 0.019716
R51382 PAD.n7699 PAD.n7090 0.019716
R51383 PAD.n7690 PAD.n7689 0.019716
R51384 PAD.n7689 PAD.n7089 0.019716
R51385 PAD.n7687 PAD.n7686 0.019716
R51386 PAD.n7687 PAD.n7088 0.019716
R51387 PAD.n7678 PAD.n7677 0.019716
R51388 PAD.n7677 PAD.n7087 0.019716
R51389 PAD.n7675 PAD.n7674 0.019716
R51390 PAD.n7675 PAD.n7086 0.019716
R51391 PAD.n7666 PAD.n7665 0.019716
R51392 PAD.n7665 PAD.n7085 0.019716
R51393 PAD.n7663 PAD.n7662 0.019716
R51394 PAD.n7663 PAD.n7084 0.019716
R51395 PAD.n7654 PAD.n7653 0.019716
R51396 PAD.n7653 PAD.n7083 0.019716
R51397 PAD.n7651 PAD.n7650 0.019716
R51398 PAD.n7651 PAD.n7082 0.019716
R51399 PAD.n7642 PAD.n7641 0.019716
R51400 PAD.n7641 PAD.n7081 0.019716
R51401 PAD.n7639 PAD.n7638 0.019716
R51402 PAD.n7639 PAD.n7080 0.019716
R51403 PAD.n7630 PAD.n7629 0.019716
R51404 PAD.n7629 PAD.n7079 0.019716
R51405 PAD.n7627 PAD.n7626 0.019716
R51406 PAD.n7627 PAD.n7078 0.019716
R51407 PAD.n7618 PAD.n7617 0.019716
R51408 PAD.n7617 PAD.n7077 0.019716
R51409 PAD.n7615 PAD.n7614 0.019716
R51410 PAD.n7615 PAD.n7076 0.019716
R51411 PAD.n7606 PAD.n7605 0.019716
R51412 PAD.n7605 PAD.n7075 0.019716
R51413 PAD.n7603 PAD.n7602 0.019716
R51414 PAD.n7603 PAD.n7074 0.019716
R51415 PAD.n7594 PAD.n7593 0.019716
R51416 PAD.n7593 PAD.n7073 0.019716
R51417 PAD.n7591 PAD.n7590 0.019716
R51418 PAD.n7591 PAD.n7072 0.019716
R51419 PAD.n7582 PAD.n7581 0.019716
R51420 PAD.n7581 PAD.n7071 0.019716
R51421 PAD.n7579 PAD.n7578 0.019716
R51422 PAD.n7579 PAD.n7070 0.019716
R51423 PAD.n7570 PAD.n7569 0.019716
R51424 PAD.n7569 PAD.n7069 0.019716
R51425 PAD.n7567 PAD.n7566 0.019716
R51426 PAD.n7567 PAD.n7068 0.019716
R51427 PAD.n7558 PAD.n7557 0.019716
R51428 PAD.n7557 PAD.n7067 0.019716
R51429 PAD.n7555 PAD.n7554 0.019716
R51430 PAD.n7555 PAD.n7066 0.019716
R51431 PAD.n7546 PAD.n7545 0.019716
R51432 PAD.n7545 PAD.n7065 0.019716
R51433 PAD.n7543 PAD.n7542 0.019716
R51434 PAD.n7543 PAD.n7064 0.019716
R51435 PAD.n7534 PAD.n7533 0.019716
R51436 PAD.n7533 PAD.n7063 0.019716
R51437 PAD.n7531 PAD.n7062 0.019716
R51438 PAD.n6721 PAD.n6719 0.019716
R51439 PAD.n7048 PAD.n7047 0.019716
R51440 PAD.n7044 PAD.n6722 0.019716
R51441 PAD.n7045 PAD.n7044 0.019716
R51442 PAD.n7038 PAD.n7035 0.019716
R51443 PAD.n7038 PAD.n7037 0.019716
R51444 PAD.n7032 PAD.n6727 0.019716
R51445 PAD.n7033 PAD.n7032 0.019716
R51446 PAD.n7026 PAD.n7023 0.019716
R51447 PAD.n7026 PAD.n7025 0.019716
R51448 PAD.n7020 PAD.n6731 0.019716
R51449 PAD.n7021 PAD.n7020 0.019716
R51450 PAD.n7014 PAD.n7011 0.019716
R51451 PAD.n7014 PAD.n7013 0.019716
R51452 PAD.n7008 PAD.n6735 0.019716
R51453 PAD.n7009 PAD.n7008 0.019716
R51454 PAD.n7002 PAD.n6999 0.019716
R51455 PAD.n7002 PAD.n7001 0.019716
R51456 PAD.n6996 PAD.n6739 0.019716
R51457 PAD.n6997 PAD.n6996 0.019716
R51458 PAD.n6990 PAD.n6987 0.019716
R51459 PAD.n6990 PAD.n6989 0.019716
R51460 PAD.n6984 PAD.n6743 0.019716
R51461 PAD.n6985 PAD.n6984 0.019716
R51462 PAD.n6978 PAD.n6975 0.019716
R51463 PAD.n6978 PAD.n6977 0.019716
R51464 PAD.n6972 PAD.n6747 0.019716
R51465 PAD.n6973 PAD.n6972 0.019716
R51466 PAD.n6966 PAD.n6963 0.019716
R51467 PAD.n6966 PAD.n6965 0.019716
R51468 PAD.n6960 PAD.n6751 0.019716
R51469 PAD.n6961 PAD.n6960 0.019716
R51470 PAD.n6954 PAD.n6951 0.019716
R51471 PAD.n6954 PAD.n6953 0.019716
R51472 PAD.n6948 PAD.n6755 0.019716
R51473 PAD.n6949 PAD.n6948 0.019716
R51474 PAD.n6942 PAD.n6939 0.019716
R51475 PAD.n6942 PAD.n6941 0.019716
R51476 PAD.n6936 PAD.n6759 0.019716
R51477 PAD.n6937 PAD.n6936 0.019716
R51478 PAD.n6930 PAD.n6927 0.019716
R51479 PAD.n6930 PAD.n6929 0.019716
R51480 PAD.n6924 PAD.n6763 0.019716
R51481 PAD.n6925 PAD.n6924 0.019716
R51482 PAD.n6918 PAD.n6915 0.019716
R51483 PAD.n6918 PAD.n6917 0.019716
R51484 PAD.n6912 PAD.n6767 0.019716
R51485 PAD.n6913 PAD.n6912 0.019716
R51486 PAD.n6906 PAD.n6903 0.019716
R51487 PAD.n6906 PAD.n6905 0.019716
R51488 PAD.n6900 PAD.n6771 0.019716
R51489 PAD.n6901 PAD.n6900 0.019716
R51490 PAD.n6894 PAD.n6891 0.019716
R51491 PAD.n6894 PAD.n6893 0.019716
R51492 PAD.n6888 PAD.n6775 0.019716
R51493 PAD.n6889 PAD.n6888 0.019716
R51494 PAD.n6882 PAD.n6879 0.019716
R51495 PAD.n6882 PAD.n6881 0.019716
R51496 PAD.n6876 PAD.n6779 0.019716
R51497 PAD.n6877 PAD.n6876 0.019716
R51498 PAD.n6870 PAD.n6867 0.019716
R51499 PAD.n6870 PAD.n6869 0.019716
R51500 PAD.n6864 PAD.n6783 0.019716
R51501 PAD.n6865 PAD.n6864 0.019716
R51502 PAD.n6858 PAD.n6855 0.019716
R51503 PAD.n6858 PAD.n6857 0.019716
R51504 PAD.n6852 PAD.n6787 0.019716
R51505 PAD.n6853 PAD.n6852 0.019716
R51506 PAD.n6846 PAD.n6843 0.019716
R51507 PAD.n6846 PAD.n6845 0.019716
R51508 PAD.n6840 PAD.n6791 0.019716
R51509 PAD.n6841 PAD.n6840 0.019716
R51510 PAD.n6834 PAD.n6831 0.019716
R51511 PAD.n6834 PAD.n6833 0.019716
R51512 PAD.n6828 PAD.n6795 0.019716
R51513 PAD.n6829 PAD.n6828 0.019716
R51514 PAD.n6822 PAD.n6819 0.019716
R51515 PAD.n6822 PAD.n6821 0.019716
R51516 PAD.n6816 PAD.n6799 0.019716
R51517 PAD.n6817 PAD.n6816 0.019716
R51518 PAD.n6810 PAD.n6807 0.019716
R51519 PAD.n6810 PAD.n6809 0.019716
R51520 PAD.n6805 PAD.n6804 0.019716
R51521 PAD.n5893 PAD.n5892 0.019716
R51522 PAD.n5603 PAD.n5602 0.019716
R51523 PAD.n5885 PAD.n5884 0.019716
R51524 PAD.n5885 PAD.n5601 0.019716
R51525 PAD.n5610 PAD.n5609 0.019716
R51526 PAD.n5610 PAD.n5600 0.019716
R51527 PAD.n5876 PAD.n5875 0.019716
R51528 PAD.n5876 PAD.n5599 0.019716
R51529 PAD.n5615 PAD.n5614 0.019716
R51530 PAD.n5615 PAD.n5598 0.019716
R51531 PAD.n5867 PAD.n5866 0.019716
R51532 PAD.n5867 PAD.n5597 0.019716
R51533 PAD.n5620 PAD.n5619 0.019716
R51534 PAD.n5620 PAD.n5596 0.019716
R51535 PAD.n5858 PAD.n5857 0.019716
R51536 PAD.n5858 PAD.n5595 0.019716
R51537 PAD.n5625 PAD.n5624 0.019716
R51538 PAD.n5625 PAD.n5594 0.019716
R51539 PAD.n5849 PAD.n5848 0.019716
R51540 PAD.n5849 PAD.n5593 0.019716
R51541 PAD.n5630 PAD.n5629 0.019716
R51542 PAD.n5630 PAD.n5592 0.019716
R51543 PAD.n5840 PAD.n5839 0.019716
R51544 PAD.n5840 PAD.n5591 0.019716
R51545 PAD.n5635 PAD.n5634 0.019716
R51546 PAD.n5635 PAD.n5590 0.019716
R51547 PAD.n5831 PAD.n5830 0.019716
R51548 PAD.n5831 PAD.n5589 0.019716
R51549 PAD.n5640 PAD.n5639 0.019716
R51550 PAD.n5640 PAD.n5588 0.019716
R51551 PAD.n5822 PAD.n5821 0.019716
R51552 PAD.n5822 PAD.n5587 0.019716
R51553 PAD.n5645 PAD.n5644 0.019716
R51554 PAD.n5645 PAD.n5586 0.019716
R51555 PAD.n5813 PAD.n5812 0.019716
R51556 PAD.n5813 PAD.n5585 0.019716
R51557 PAD.n5650 PAD.n5649 0.019716
R51558 PAD.n5650 PAD.n5584 0.019716
R51559 PAD.n5804 PAD.n5803 0.019716
R51560 PAD.n5804 PAD.n5583 0.019716
R51561 PAD.n5655 PAD.n5654 0.019716
R51562 PAD.n5655 PAD.n5582 0.019716
R51563 PAD.n5795 PAD.n5794 0.019716
R51564 PAD.n5795 PAD.n5581 0.019716
R51565 PAD.n5660 PAD.n5659 0.019716
R51566 PAD.n5660 PAD.n5580 0.019716
R51567 PAD.n5786 PAD.n5785 0.019716
R51568 PAD.n5786 PAD.n5579 0.019716
R51569 PAD.n5665 PAD.n5664 0.019716
R51570 PAD.n5665 PAD.n5578 0.019716
R51571 PAD.n5777 PAD.n5776 0.019716
R51572 PAD.n5777 PAD.n5577 0.019716
R51573 PAD.n5670 PAD.n5669 0.019716
R51574 PAD.n5670 PAD.n5576 0.019716
R51575 PAD.n5768 PAD.n5767 0.019716
R51576 PAD.n5768 PAD.n5575 0.019716
R51577 PAD.n5675 PAD.n5674 0.019716
R51578 PAD.n5675 PAD.n5574 0.019716
R51579 PAD.n5759 PAD.n5758 0.019716
R51580 PAD.n5759 PAD.n5573 0.019716
R51581 PAD.n5680 PAD.n5679 0.019716
R51582 PAD.n5680 PAD.n5572 0.019716
R51583 PAD.n5750 PAD.n5749 0.019716
R51584 PAD.n5750 PAD.n5571 0.019716
R51585 PAD.n5685 PAD.n5684 0.019716
R51586 PAD.n5685 PAD.n5570 0.019716
R51587 PAD.n5741 PAD.n5740 0.019716
R51588 PAD.n5741 PAD.n5569 0.019716
R51589 PAD.n5690 PAD.n5689 0.019716
R51590 PAD.n5690 PAD.n5568 0.019716
R51591 PAD.n5732 PAD.n5731 0.019716
R51592 PAD.n5732 PAD.n5567 0.019716
R51593 PAD.n5695 PAD.n5694 0.019716
R51594 PAD.n5695 PAD.n5566 0.019716
R51595 PAD.n5723 PAD.n5722 0.019716
R51596 PAD.n5723 PAD.n5565 0.019716
R51597 PAD.n5700 PAD.n5699 0.019716
R51598 PAD.n5700 PAD.n5564 0.019716
R51599 PAD.n5714 PAD.n5713 0.019716
R51600 PAD.n5714 PAD.n5563 0.019716
R51601 PAD.n5707 PAD.n5706 0.019716
R51602 PAD.n5707 PAD.n5562 0.019716
R51603 PAD.n5702 PAD.n5561 0.019716
R51604 PAD.n6690 PAD.n5902 0.019716
R51605 PAD.n6497 PAD.n6397 0.019716
R51606 PAD.n6497 PAD.n5906 0.019716
R51607 PAD.n6502 PAD.n6398 0.019716
R51608 PAD.n6502 PAD.n5907 0.019716
R51609 PAD.n6506 PAD.n6399 0.019716
R51610 PAD.n6506 PAD.n5908 0.019716
R51611 PAD.n6511 PAD.n6400 0.019716
R51612 PAD.n6511 PAD.n5909 0.019716
R51613 PAD.n6515 PAD.n6401 0.019716
R51614 PAD.n6515 PAD.n5910 0.019716
R51615 PAD.n6520 PAD.n6402 0.019716
R51616 PAD.n6520 PAD.n5911 0.019716
R51617 PAD.n6524 PAD.n6403 0.019716
R51618 PAD.n6524 PAD.n5912 0.019716
R51619 PAD.n6529 PAD.n6404 0.019716
R51620 PAD.n6529 PAD.n5913 0.019716
R51621 PAD.n6533 PAD.n6405 0.019716
R51622 PAD.n6533 PAD.n5914 0.019716
R51623 PAD.n6538 PAD.n6406 0.019716
R51624 PAD.n6538 PAD.n5915 0.019716
R51625 PAD.n6542 PAD.n6407 0.019716
R51626 PAD.n6542 PAD.n5916 0.019716
R51627 PAD.n6547 PAD.n6408 0.019716
R51628 PAD.n6547 PAD.n5917 0.019716
R51629 PAD.n6551 PAD.n6409 0.019716
R51630 PAD.n6551 PAD.n5918 0.019716
R51631 PAD.n6556 PAD.n6410 0.019716
R51632 PAD.n6556 PAD.n5919 0.019716
R51633 PAD.n6560 PAD.n6411 0.019716
R51634 PAD.n6560 PAD.n5920 0.019716
R51635 PAD.n6565 PAD.n6412 0.019716
R51636 PAD.n6565 PAD.n5921 0.019716
R51637 PAD.n6569 PAD.n6413 0.019716
R51638 PAD.n6569 PAD.n5922 0.019716
R51639 PAD.n6574 PAD.n6414 0.019716
R51640 PAD.n6574 PAD.n5923 0.019716
R51641 PAD.n6578 PAD.n6415 0.019716
R51642 PAD.n6578 PAD.n5924 0.019716
R51643 PAD.n6583 PAD.n6416 0.019716
R51644 PAD.n6583 PAD.n5925 0.019716
R51645 PAD.n6587 PAD.n6417 0.019716
R51646 PAD.n6587 PAD.n5926 0.019716
R51647 PAD.n6592 PAD.n6418 0.019716
R51648 PAD.n6592 PAD.n5927 0.019716
R51649 PAD.n6596 PAD.n6419 0.019716
R51650 PAD.n6596 PAD.n5928 0.019716
R51651 PAD.n6601 PAD.n6420 0.019716
R51652 PAD.n6601 PAD.n5929 0.019716
R51653 PAD.n6605 PAD.n6421 0.019716
R51654 PAD.n6605 PAD.n5930 0.019716
R51655 PAD.n6610 PAD.n6422 0.019716
R51656 PAD.n6610 PAD.n5931 0.019716
R51657 PAD.n6614 PAD.n6423 0.019716
R51658 PAD.n6614 PAD.n5932 0.019716
R51659 PAD.n6619 PAD.n6424 0.019716
R51660 PAD.n6619 PAD.n5933 0.019716
R51661 PAD.n6623 PAD.n6425 0.019716
R51662 PAD.n6623 PAD.n5934 0.019716
R51663 PAD.n6628 PAD.n6426 0.019716
R51664 PAD.n6628 PAD.n5935 0.019716
R51665 PAD.n6632 PAD.n6427 0.019716
R51666 PAD.n6632 PAD.n5936 0.019716
R51667 PAD.n6637 PAD.n6428 0.019716
R51668 PAD.n6637 PAD.n5937 0.019716
R51669 PAD.n6641 PAD.n6429 0.019716
R51670 PAD.n6641 PAD.n5938 0.019716
R51671 PAD.n6646 PAD.n6430 0.019716
R51672 PAD.n6646 PAD.n5939 0.019716
R51673 PAD.n6650 PAD.n6431 0.019716
R51674 PAD.n6650 PAD.n5940 0.019716
R51675 PAD.n6655 PAD.n6432 0.019716
R51676 PAD.n6655 PAD.n5941 0.019716
R51677 PAD.n6659 PAD.n6433 0.019716
R51678 PAD.n6659 PAD.n5942 0.019716
R51679 PAD.n6664 PAD.n6434 0.019716
R51680 PAD.n6664 PAD.n5943 0.019716
R51681 PAD.n6668 PAD.n6435 0.019716
R51682 PAD.n6668 PAD.n5944 0.019716
R51683 PAD.n6677 PAD.n6676 0.019716
R51684 PAD.n6676 PAD.n5945 0.019716
R51685 PAD.n5949 PAD.n5947 0.019716
R51686 PAD.n5949 PAD.n5946 0.019716
R51687 PAD.n9133 PAD.n2882 0.019625
R51688 PAD.n10733 PAD.n10732 0.019625
R51689 PAD.n9719 PAD.n1590 0.0195611
R51690 PAD.n10019 PAD.n1138 0.0195611
R51691 PAD.n9720 PAD.n1591 0.0195611
R51692 PAD.n10018 PAD.n1139 0.0195611
R51693 PAD.n9157 PAD.n9156 0.019175
R51694 PAD.n10709 PAD.n422 0.019175
R51695 PAD.n8459 PAD.n8458 0.0191681
R51696 PAD.n3686 PAD.n3632 0.0191681
R51697 PAD.n6686 PAD.n6685 0.0187751
R51698 PAD.n6684 PAD.n5948 0.0187751
R51699 PAD.n7825 PAD.n7824 0.018725
R51700 PAD.n7523 PAD.n7156 0.0175961
R51701 PAD.n7522 PAD.n7157 0.0175961
R51702 PAD.n6392 PAD.n6391 0.017282
R51703 PAD.n6392 PAD.n5897 0.017282
R51704 PAD.n6695 PAD.n6694 0.017282
R51705 PAD.n6695 PAD.n5544 0.017282
R51706 PAD.n7805 PAD.n5546 0.017282
R51707 PAD.n7054 PAD.n5546 0.017282
R51708 PAD.n7788 PAD.n7787 0.017282
R51709 PAD.n7787 PAD.n7786 0.017282
R51710 PAD.n7212 PAD.n7210 0.017282
R51711 PAD.n7220 PAD.n7210 0.017282
R51712 PAD.n7227 PAD.n7220 0.017282
R51713 PAD.n7227 PAD.n7226 0.017282
R51714 PAD.n7226 PAD.n5209 0.017282
R51715 PAD.n7816 PAD.n5209 0.017282
R51716 PAD.n8169 PAD.n5194 0.017282
R51717 PAD.n8171 PAD.n5180 0.017282
R51718 PAD.n8189 PAD.n5180 0.017282
R51719 PAD.n8191 PAD.n4677 0.017282
R51720 PAD.n8401 PAD.n4677 0.017282
R51721 PAD.n8404 PAD.n8403 0.017282
R51722 PAD.n8404 PAD.n4326 0.017282
R51723 PAD.n8423 PAD.n4326 0.017282
R51724 PAD.n8427 PAD.n8425 0.017282
R51725 PAD.n8427 PAD.n8426 0.017282
R51726 PAD.n8449 PAD.n8448 0.017282
R51727 PAD.n8450 PAD.n8449 0.017282
R51728 PAD.n8475 PAD.n8474 0.017282
R51729 PAD.n8497 PAD.n8496 0.017282
R51730 PAD.n8499 PAD.n8497 0.017282
R51731 PAD.n8499 PAD.n8498 0.017282
R51732 PAD.n8523 PAD.n8522 0.017282
R51733 PAD.n8524 PAD.n8523 0.017282
R51734 PAD.n8836 PAD.n8835 0.017282
R51735 PAD.n9125 PAD.n8836 0.017282
R51736 PAD.n9123 PAD.n2831 0.017282
R51737 PAD.n9146 PAD.n2831 0.017282
R51738 PAD.n9148 PAD.n2484 0.017282
R51739 PAD.n9166 PAD.n2484 0.017282
R51740 PAD.n9170 PAD.n9169 0.017282
R51741 PAD.n9169 PAD.n2137 0.017282
R51742 PAD.n9194 PAD.n9193 0.017282
R51743 PAD.n9193 PAD.n9192 0.017282
R51744 PAD.n2034 PAD.n1933 0.017282
R51745 PAD.n9725 PAD.n1933 0.017282
R51746 PAD.n9729 PAD.n9728 0.017282
R51747 PAD.n9728 PAD.n9727 0.017282
R51748 PAD.n1584 PAD.n1583 0.017282
R51749 PAD.n1583 PAD.n1146 0.017282
R51750 PAD.n10011 PAD.n1146 0.017282
R51751 PAD.n10013 PAD.n1125 0.017282
R51752 PAD.n10365 PAD.n1125 0.017282
R51753 PAD.n10370 PAD.n10368 0.017282
R51754 PAD.n10370 PAD.n10369 0.017282
R51755 PAD.n10393 PAD.n10392 0.017282
R51756 PAD.n10394 PAD.n10393 0.017282
R51757 PAD.n10412 PAD.n10411 0.017282
R51758 PAD.n10698 PAD.n10412 0.017282
R51759 PAD.n10722 PAD.n370 0.017282
R51760 PAD.n10723 PAD.n10722 0.017282
R51761 PAD.n10724 PAD.n10723 0.017282
R51762 PAD.n11537 PAD.n15 0.017282
R51763 PAD.n10746 PAD.n15 0.017282
R51764 PAD.n11519 PAD.n11089 0.017282
R51765 PAD.n11519 PAD.n11518 0.017282
R51766 PAD.n2897 PAD.n2883 0.0172031
R51767 PAD.n29 PAD.n24 0.0172031
R51768 PAD.n2895 PAD.n2878 0.0172031
R51769 PAD.n31 PAD.n22 0.0172031
R51770 PAD.n8437 PAD.n4315 0.016925
R51771 PAD.n9158 PAD.n2489 0.01681
R51772 PAD.n10705 PAD.n10704 0.01681
R51773 PAD.n9159 PAD.n2488 0.01681
R51774 PAD.n10703 PAD.n417 0.01681
R51775 PAD.n8522 PAD.n2949 0.0167406
R51776 PAD.n10698 PAD.n10697 0.0167406
R51777 PAD.n9738 PAD.n1486 0.016475
R51778 PAD.n10002 PAD.n1486 0.016475
R51779 PAD.n11518 PAD.n11517 0.0164699
R51780 PAD.n7826 PAD.n5199 0.016417
R51781 PAD.n7827 PAD.n5198 0.016417
R51782 PAD.n9167 PAD.n9166 0.0161992
R51783 PAD.n10013 PAD.n10012 0.0161992
R51784 PAD.n8437 PAD.n8436 0.016025
R51785 PAD.n6694 PAD.n6693 0.0156579
R51786 PAD.n8402 PAD.n8401 0.0156579
R51787 PAD.n6393 PAD.n5955 0.0154799
R51788 PAD.n6394 PAD.n6393 0.0154799
R51789 PAD.n6696 PAD.n5896 0.0154799
R51790 PAD.n6697 PAD.n6696 0.0154799
R51791 PAD.n7804 PAD.n5548 0.0154799
R51792 PAD.n7053 PAD.n5548 0.0154799
R51793 PAD.n7789 PAD.n6717 0.0154799
R51794 PAD.n7785 PAD.n6717 0.0154799
R51795 PAD.n7213 PAD.n7211 0.0154799
R51796 PAD.n7219 PAD.n7211 0.0154799
R51797 PAD.n7219 PAD.n7208 0.0154799
R51798 PAD.n7225 PAD.n7208 0.0154799
R51799 PAD.n7225 PAD.n5207 0.0154799
R51800 PAD.n7817 PAD.n5207 0.0154799
R51801 PAD.n7813 PAD.n5195 0.0154799
R51802 PAD.n8168 PAD.n5195 0.0154799
R51803 PAD.n8172 PAD.n5181 0.0154799
R51804 PAD.n8188 PAD.n5181 0.0154799
R51805 PAD.n8192 PAD.n4678 0.0154799
R51806 PAD.n8400 PAD.n4678 0.0154799
R51807 PAD.n8405 PAD.n4675 0.0154799
R51808 PAD.n8405 PAD.n4327 0.0154799
R51809 PAD.n8422 PAD.n4327 0.0154799
R51810 PAD.n8428 PAD.n4323 0.0154799
R51811 PAD.n8428 PAD.n4324 0.0154799
R51812 PAD.n8447 PAD.n3979 0.0154799
R51813 PAD.n8451 PAD.n3979 0.0154799
R51814 PAD.n8471 PAD.n3635 0.0154799
R51815 PAD.n8476 PAD.n3635 0.0154799
R51816 PAD.n8495 PAD.n3291 0.0154799
R51817 PAD.n8500 PAD.n3291 0.0154799
R51818 PAD.n8500 PAD.n3292 0.0154799
R51819 PAD.n8521 PAD.n2948 0.0154799
R51820 PAD.n8525 PAD.n2948 0.0154799
R51821 PAD.n8834 PAD.n2886 0.0154799
R51822 PAD.n9126 PAD.n2886 0.0154799
R51823 PAD.n9122 PAD.n2832 0.0154799
R51824 PAD.n9145 PAD.n2832 0.0154799
R51825 PAD.n9149 PAD.n2485 0.0154799
R51826 PAD.n9165 PAD.n2485 0.0154799
R51827 PAD.n9173 PAD.n2149 0.0154799
R51828 PAD.n2149 PAD.n2136 0.0154799
R51829 PAD.n9191 PAD.n2136 0.0154799
R51830 PAD.n9195 PAD.n2036 0.0154799
R51831 PAD.n2036 PAD.n2033 0.0154799
R51832 PAD.n9461 PAD.n1934 0.0154799
R51833 PAD.n9724 PAD.n1934 0.0154799
R51834 PAD.n9730 PAD.n1597 0.0154799
R51835 PAD.n1597 PAD.n1581 0.0154799
R51836 PAD.n9747 PAD.n1582 0.0154799
R51837 PAD.n1582 PAD.n1147 0.0154799
R51838 PAD.n10010 PAD.n1147 0.0154799
R51839 PAD.n10014 PAD.n1126 0.0154799
R51840 PAD.n10364 PAD.n1126 0.0154799
R51841 PAD.n10371 PAD.n1122 0.0154799
R51842 PAD.n10371 PAD.n1123 0.0154799
R51843 PAD.n10391 PAD.n778 0.0154799
R51844 PAD.n10395 PAD.n778 0.0154799
R51845 PAD.n10410 PAD.n428 0.0154799
R51846 PAD.n10699 PAD.n428 0.0154799
R51847 PAD.n10721 PAD.n371 0.0154799
R51848 PAD.n10721 PAD.n369 0.0154799
R51849 PAD.n10725 PAD.n369 0.0154799
R51850 PAD.n11536 PAD.n17 0.0154799
R51851 PAD.n10751 PAD.n17 0.0154799
R51852 PAD.n11520 PAD.n10744 0.0154799
R51853 PAD.n11520 PAD.n10745 0.0154799
R51854 PAD.n5970 PAD.n5954 0.0154799
R51855 PAD.n6395 PAD.n5954 0.0154799
R51856 PAD.n6681 PAD.n5895 0.0154799
R51857 PAD.n6698 PAD.n5895 0.0154799
R51858 PAD.n7803 PAD.n5550 0.0154799
R51859 PAD.n7052 PAD.n5550 0.0154799
R51860 PAD.n7790 PAD.n6715 0.0154799
R51861 PAD.n7784 PAD.n6715 0.0154799
R51862 PAD.n7217 PAD.n7214 0.0154799
R51863 PAD.n7218 PAD.n7217 0.0154799
R51864 PAD.n7218 PAD.n7202 0.0154799
R51865 PAD.n7224 PAD.n7202 0.0154799
R51866 PAD.n7224 PAD.n5205 0.0154799
R51867 PAD.n7818 PAD.n5205 0.0154799
R51868 PAD.n8166 PAD.n5196 0.0154799
R51869 PAD.n8167 PAD.n8166 0.0154799
R51870 PAD.n8173 PAD.n5182 0.0154799
R51871 PAD.n8187 PAD.n5182 0.0154799
R51872 PAD.n8193 PAD.n4680 0.0154799
R51873 PAD.n8399 PAD.n4680 0.0154799
R51874 PAD.n8406 PAD.n4674 0.0154799
R51875 PAD.n8406 PAD.n4329 0.0154799
R51876 PAD.n8421 PAD.n4329 0.0154799
R51877 PAD.n8429 PAD.n4320 0.0154799
R51878 PAD.n8429 PAD.n4322 0.0154799
R51879 PAD.n8446 PAD.n3978 0.0154799
R51880 PAD.n8452 PAD.n3978 0.0154799
R51881 PAD.n8470 PAD.n3634 0.0154799
R51882 PAD.n8477 PAD.n3634 0.0154799
R51883 PAD.n8494 PAD.n3288 0.0154799
R51884 PAD.n8501 PAD.n3288 0.0154799
R51885 PAD.n8501 PAD.n3290 0.0154799
R51886 PAD.n8520 PAD.n2947 0.0154799
R51887 PAD.n8526 PAD.n2947 0.0154799
R51888 PAD.n8833 PAD.n2884 0.0154799
R51889 PAD.n9127 PAD.n2884 0.0154799
R51890 PAD.n9121 PAD.n2833 0.0154799
R51891 PAD.n9144 PAD.n2833 0.0154799
R51892 PAD.n9150 PAD.n2486 0.0154799
R51893 PAD.n9164 PAD.n2486 0.0154799
R51894 PAD.n9174 PAD.n2138 0.0154799
R51895 PAD.n9188 PAD.n2138 0.0154799
R51896 PAD.n9190 PAD.n9188 0.0154799
R51897 PAD.n9457 PAD.n2035 0.0154799
R51898 PAD.n9458 PAD.n9457 0.0154799
R51899 PAD.n9460 PAD.n1935 0.0154799
R51900 PAD.n9723 PAD.n1935 0.0154799
R51901 PAD.n9731 PAD.n1585 0.0154799
R51902 PAD.n9743 PAD.n1585 0.0154799
R51903 PAD.n9746 PAD.n9745 0.0154799
R51904 PAD.n9745 PAD.n1148 0.0154799
R51905 PAD.n10009 PAD.n1148 0.0154799
R51906 PAD.n10015 PAD.n1128 0.0154799
R51907 PAD.n10363 PAD.n1128 0.0154799
R51908 PAD.n10372 PAD.n1119 0.0154799
R51909 PAD.n10372 PAD.n1121 0.0154799
R51910 PAD.n10390 PAD.n777 0.0154799
R51911 PAD.n10396 PAD.n777 0.0154799
R51912 PAD.n10409 PAD.n426 0.0154799
R51913 PAD.n10700 PAD.n426 0.0154799
R51914 PAD.n10720 PAD.n372 0.0154799
R51915 PAD.n10720 PAD.n368 0.0154799
R51916 PAD.n10726 PAD.n368 0.0154799
R51917 PAD.n11535 PAD.n19 0.0154799
R51918 PAD.n10752 PAD.n19 0.0154799
R51919 PAD.n11521 PAD.n10742 0.0154799
R51920 PAD.n11521 PAD.n10743 0.0154799
R51921 PAD.n8425 PAD.n8424 0.0151165
R51922 PAD.n8521 PAD.n2950 0.0149966
R51923 PAD.n10699 PAD.n429 0.0149966
R51924 PAD.n8520 PAD.n2951 0.0149966
R51925 PAD.n10700 PAD.n427 0.0149966
R51926 PAD.n8434 PAD.n8433 0.014845
R51927 PAD.n8432 PAD.n4027 0.014845
R51928 PAD.n11092 PAD.n10745 0.014755
R51929 PAD.n11094 PAD.n10743 0.014755
R51930 PAD.n9194 PAD.n2135 0.0145752
R51931 PAD.n9727 PAD.n1580 0.0145752
R51932 PAD.n9165 PAD.n2148 0.0145134
R51933 PAD.n10014 PAD.n1144 0.0145134
R51934 PAD.n9164 PAD.n2147 0.0145134
R51935 PAD.n10015 PAD.n1143 0.0145134
R51936 PAD.n9739 PAD.n1487 0.014452
R51937 PAD.n10001 PAD.n1487 0.014452
R51938 PAD.n9740 PAD.n1488 0.014452
R51939 PAD.n10000 PAD.n1488 0.014452
R51940 PAD.n11515 PAD.n11093 0.01445
R51941 PAD.n11354 PAD.n11353 0.01445
R51942 PAD.n11354 PAD.n11351 0.01445
R51943 PAD.n11358 PAD.n11351 0.01445
R51944 PAD.n11359 PAD.n11358 0.01445
R51945 PAD.n11360 PAD.n11359 0.01445
R51946 PAD.n11360 PAD.n11349 0.01445
R51947 PAD.n11364 PAD.n11349 0.01445
R51948 PAD.n11365 PAD.n11364 0.01445
R51949 PAD.n11366 PAD.n11365 0.01445
R51950 PAD.n11366 PAD.n11347 0.01445
R51951 PAD.n11370 PAD.n11347 0.01445
R51952 PAD.n11371 PAD.n11370 0.01445
R51953 PAD.n11372 PAD.n11371 0.01445
R51954 PAD.n11372 PAD.n11345 0.01445
R51955 PAD.n11376 PAD.n11345 0.01445
R51956 PAD.n11377 PAD.n11376 0.01445
R51957 PAD.n11378 PAD.n11377 0.01445
R51958 PAD.n11378 PAD.n11343 0.01445
R51959 PAD.n11382 PAD.n11343 0.01445
R51960 PAD.n11383 PAD.n11382 0.01445
R51961 PAD.n11384 PAD.n11383 0.01445
R51962 PAD.n11384 PAD.n11341 0.01445
R51963 PAD.n11388 PAD.n11341 0.01445
R51964 PAD.n11389 PAD.n11388 0.01445
R51965 PAD.n11390 PAD.n11389 0.01445
R51966 PAD.n11390 PAD.n11339 0.01445
R51967 PAD.n11394 PAD.n11339 0.01445
R51968 PAD.n11395 PAD.n11394 0.01445
R51969 PAD.n11396 PAD.n11395 0.01445
R51970 PAD.n11396 PAD.n11337 0.01445
R51971 PAD.n11400 PAD.n11337 0.01445
R51972 PAD.n11401 PAD.n11400 0.01445
R51973 PAD.n11402 PAD.n11401 0.01445
R51974 PAD.n11402 PAD.n11335 0.01445
R51975 PAD.n11406 PAD.n11335 0.01445
R51976 PAD.n11407 PAD.n11406 0.01445
R51977 PAD.n11408 PAD.n11407 0.01445
R51978 PAD.n11408 PAD.n11333 0.01445
R51979 PAD.n11412 PAD.n11333 0.01445
R51980 PAD.n11413 PAD.n11412 0.01445
R51981 PAD.n11414 PAD.n11413 0.01445
R51982 PAD.n11414 PAD.n11331 0.01445
R51983 PAD.n11418 PAD.n11331 0.01445
R51984 PAD.n11419 PAD.n11418 0.01445
R51985 PAD.n11420 PAD.n11419 0.01445
R51986 PAD.n11420 PAD.n11329 0.01445
R51987 PAD.n11424 PAD.n11329 0.01445
R51988 PAD.n11425 PAD.n11424 0.01445
R51989 PAD.n11426 PAD.n11425 0.01445
R51990 PAD.n11426 PAD.n11327 0.01445
R51991 PAD.n11430 PAD.n11327 0.01445
R51992 PAD.n11431 PAD.n11430 0.01445
R51993 PAD.n11432 PAD.n11431 0.01445
R51994 PAD.n11432 PAD.n11325 0.01445
R51995 PAD.n11436 PAD.n11325 0.01445
R51996 PAD.n11437 PAD.n11436 0.01445
R51997 PAD.n11438 PAD.n11437 0.01445
R51998 PAD.n11438 PAD.n11323 0.01445
R51999 PAD.n11442 PAD.n11323 0.01445
R52000 PAD.n11443 PAD.n11442 0.01445
R52001 PAD.n11444 PAD.n11443 0.01445
R52002 PAD.n11444 PAD.n11321 0.01445
R52003 PAD.n11448 PAD.n11321 0.01445
R52004 PAD.n11449 PAD.n11448 0.01445
R52005 PAD.n11450 PAD.n11449 0.01445
R52006 PAD.n11450 PAD.n11319 0.01445
R52007 PAD.n11454 PAD.n11319 0.01445
R52008 PAD.n11455 PAD.n11454 0.01445
R52009 PAD.n11456 PAD.n11455 0.01445
R52010 PAD.n11456 PAD.n11317 0.01445
R52011 PAD.n11460 PAD.n11317 0.01445
R52012 PAD.n11461 PAD.n11460 0.01445
R52013 PAD.n11462 PAD.n11461 0.01445
R52014 PAD.n11462 PAD.n11315 0.01445
R52015 PAD.n11466 PAD.n11315 0.01445
R52016 PAD.n11467 PAD.n11466 0.01445
R52017 PAD.n11468 PAD.n11467 0.01445
R52018 PAD.n11468 PAD.n11313 0.01445
R52019 PAD.n11472 PAD.n11313 0.01445
R52020 PAD.n11473 PAD.n11472 0.01445
R52021 PAD.n11474 PAD.n11473 0.01445
R52022 PAD.n11474 PAD.n11311 0.01445
R52023 PAD.n11478 PAD.n11311 0.01445
R52024 PAD.n11479 PAD.n11478 0.01445
R52025 PAD.n11480 PAD.n11479 0.01445
R52026 PAD.n11480 PAD.n11309 0.01445
R52027 PAD.n11484 PAD.n11309 0.01445
R52028 PAD.n11485 PAD.n11484 0.01445
R52029 PAD.n11486 PAD.n11485 0.01445
R52030 PAD.n11486 PAD.n11307 0.01445
R52031 PAD.n11490 PAD.n11307 0.01445
R52032 PAD.n11491 PAD.n11490 0.01445
R52033 PAD.n11492 PAD.n11491 0.01445
R52034 PAD.n11492 PAD.n11305 0.01445
R52035 PAD.n11496 PAD.n11305 0.01445
R52036 PAD.n11497 PAD.n11496 0.01445
R52037 PAD.n11498 PAD.n11497 0.01445
R52038 PAD.n11516 PAD.n11091 0.01445
R52039 PAD.n11355 PAD.n11352 0.01445
R52040 PAD.n11356 PAD.n11355 0.01445
R52041 PAD.n11357 PAD.n11356 0.01445
R52042 PAD.n11357 PAD.n11350 0.01445
R52043 PAD.n11361 PAD.n11350 0.01445
R52044 PAD.n11362 PAD.n11361 0.01445
R52045 PAD.n11363 PAD.n11362 0.01445
R52046 PAD.n11363 PAD.n11348 0.01445
R52047 PAD.n11367 PAD.n11348 0.01445
R52048 PAD.n11368 PAD.n11367 0.01445
R52049 PAD.n11369 PAD.n11368 0.01445
R52050 PAD.n11369 PAD.n11346 0.01445
R52051 PAD.n11373 PAD.n11346 0.01445
R52052 PAD.n11374 PAD.n11373 0.01445
R52053 PAD.n11375 PAD.n11374 0.01445
R52054 PAD.n11375 PAD.n11344 0.01445
R52055 PAD.n11379 PAD.n11344 0.01445
R52056 PAD.n11380 PAD.n11379 0.01445
R52057 PAD.n11381 PAD.n11380 0.01445
R52058 PAD.n11381 PAD.n11342 0.01445
R52059 PAD.n11385 PAD.n11342 0.01445
R52060 PAD.n11386 PAD.n11385 0.01445
R52061 PAD.n11387 PAD.n11386 0.01445
R52062 PAD.n11387 PAD.n11340 0.01445
R52063 PAD.n11391 PAD.n11340 0.01445
R52064 PAD.n11392 PAD.n11391 0.01445
R52065 PAD.n11393 PAD.n11392 0.01445
R52066 PAD.n11393 PAD.n11338 0.01445
R52067 PAD.n11397 PAD.n11338 0.01445
R52068 PAD.n11398 PAD.n11397 0.01445
R52069 PAD.n11399 PAD.n11398 0.01445
R52070 PAD.n11399 PAD.n11336 0.01445
R52071 PAD.n11403 PAD.n11336 0.01445
R52072 PAD.n11404 PAD.n11403 0.01445
R52073 PAD.n11405 PAD.n11404 0.01445
R52074 PAD.n11405 PAD.n11334 0.01445
R52075 PAD.n11409 PAD.n11334 0.01445
R52076 PAD.n11410 PAD.n11409 0.01445
R52077 PAD.n11411 PAD.n11410 0.01445
R52078 PAD.n11411 PAD.n11332 0.01445
R52079 PAD.n11415 PAD.n11332 0.01445
R52080 PAD.n11416 PAD.n11415 0.01445
R52081 PAD.n11417 PAD.n11416 0.01445
R52082 PAD.n11417 PAD.n11330 0.01445
R52083 PAD.n11421 PAD.n11330 0.01445
R52084 PAD.n11422 PAD.n11421 0.01445
R52085 PAD.n11423 PAD.n11422 0.01445
R52086 PAD.n11423 PAD.n11328 0.01445
R52087 PAD.n11427 PAD.n11328 0.01445
R52088 PAD.n11428 PAD.n11427 0.01445
R52089 PAD.n11429 PAD.n11428 0.01445
R52090 PAD.n11429 PAD.n11326 0.01445
R52091 PAD.n11433 PAD.n11326 0.01445
R52092 PAD.n11434 PAD.n11433 0.01445
R52093 PAD.n11435 PAD.n11434 0.01445
R52094 PAD.n11435 PAD.n11324 0.01445
R52095 PAD.n11439 PAD.n11324 0.01445
R52096 PAD.n11440 PAD.n11439 0.01445
R52097 PAD.n11441 PAD.n11440 0.01445
R52098 PAD.n11441 PAD.n11322 0.01445
R52099 PAD.n11445 PAD.n11322 0.01445
R52100 PAD.n11446 PAD.n11445 0.01445
R52101 PAD.n11447 PAD.n11446 0.01445
R52102 PAD.n11447 PAD.n11320 0.01445
R52103 PAD.n11451 PAD.n11320 0.01445
R52104 PAD.n11452 PAD.n11451 0.01445
R52105 PAD.n11453 PAD.n11452 0.01445
R52106 PAD.n11453 PAD.n11318 0.01445
R52107 PAD.n11457 PAD.n11318 0.01445
R52108 PAD.n11458 PAD.n11457 0.01445
R52109 PAD.n11459 PAD.n11458 0.01445
R52110 PAD.n11459 PAD.n11316 0.01445
R52111 PAD.n11463 PAD.n11316 0.01445
R52112 PAD.n11464 PAD.n11463 0.01445
R52113 PAD.n11465 PAD.n11464 0.01445
R52114 PAD.n11465 PAD.n11314 0.01445
R52115 PAD.n11469 PAD.n11314 0.01445
R52116 PAD.n11470 PAD.n11469 0.01445
R52117 PAD.n11471 PAD.n11470 0.01445
R52118 PAD.n11471 PAD.n11312 0.01445
R52119 PAD.n11475 PAD.n11312 0.01445
R52120 PAD.n11476 PAD.n11475 0.01445
R52121 PAD.n11477 PAD.n11476 0.01445
R52122 PAD.n11477 PAD.n11310 0.01445
R52123 PAD.n11481 PAD.n11310 0.01445
R52124 PAD.n11482 PAD.n11481 0.01445
R52125 PAD.n11483 PAD.n11482 0.01445
R52126 PAD.n11483 PAD.n11308 0.01445
R52127 PAD.n11487 PAD.n11308 0.01445
R52128 PAD.n11488 PAD.n11487 0.01445
R52129 PAD.n11489 PAD.n11488 0.01445
R52130 PAD.n11489 PAD.n11306 0.01445
R52131 PAD.n11493 PAD.n11306 0.01445
R52132 PAD.n11494 PAD.n11493 0.01445
R52133 PAD.n11495 PAD.n11494 0.01445
R52134 PAD.n11495 PAD.n11304 0.01445
R52135 PAD.n11499 PAD.n11304 0.01445
R52136 PAD.n6388 PAD.n5959 0.01445
R52137 PAD.n6227 PAD.n6226 0.01445
R52138 PAD.n6228 PAD.n6227 0.01445
R52139 PAD.n6228 PAD.n6223 0.01445
R52140 PAD.n6232 PAD.n6223 0.01445
R52141 PAD.n6233 PAD.n6232 0.01445
R52142 PAD.n6234 PAD.n6233 0.01445
R52143 PAD.n6234 PAD.n6221 0.01445
R52144 PAD.n6238 PAD.n6221 0.01445
R52145 PAD.n6239 PAD.n6238 0.01445
R52146 PAD.n6240 PAD.n6239 0.01445
R52147 PAD.n6240 PAD.n6219 0.01445
R52148 PAD.n6244 PAD.n6219 0.01445
R52149 PAD.n6245 PAD.n6244 0.01445
R52150 PAD.n6246 PAD.n6245 0.01445
R52151 PAD.n6246 PAD.n6217 0.01445
R52152 PAD.n6250 PAD.n6217 0.01445
R52153 PAD.n6251 PAD.n6250 0.01445
R52154 PAD.n6252 PAD.n6251 0.01445
R52155 PAD.n6252 PAD.n6215 0.01445
R52156 PAD.n6256 PAD.n6215 0.01445
R52157 PAD.n6257 PAD.n6256 0.01445
R52158 PAD.n6258 PAD.n6257 0.01445
R52159 PAD.n6258 PAD.n6213 0.01445
R52160 PAD.n6262 PAD.n6213 0.01445
R52161 PAD.n6263 PAD.n6262 0.01445
R52162 PAD.n6264 PAD.n6263 0.01445
R52163 PAD.n6264 PAD.n6211 0.01445
R52164 PAD.n6268 PAD.n6211 0.01445
R52165 PAD.n6269 PAD.n6268 0.01445
R52166 PAD.n6270 PAD.n6269 0.01445
R52167 PAD.n6270 PAD.n6209 0.01445
R52168 PAD.n6274 PAD.n6209 0.01445
R52169 PAD.n6275 PAD.n6274 0.01445
R52170 PAD.n6276 PAD.n6275 0.01445
R52171 PAD.n6276 PAD.n6207 0.01445
R52172 PAD.n6280 PAD.n6207 0.01445
R52173 PAD.n6281 PAD.n6280 0.01445
R52174 PAD.n6282 PAD.n6281 0.01445
R52175 PAD.n6282 PAD.n6205 0.01445
R52176 PAD.n6286 PAD.n6205 0.01445
R52177 PAD.n6287 PAD.n6286 0.01445
R52178 PAD.n6288 PAD.n6287 0.01445
R52179 PAD.n6288 PAD.n6203 0.01445
R52180 PAD.n6292 PAD.n6203 0.01445
R52181 PAD.n6293 PAD.n6292 0.01445
R52182 PAD.n6294 PAD.n6293 0.01445
R52183 PAD.n6294 PAD.n6201 0.01445
R52184 PAD.n6298 PAD.n6201 0.01445
R52185 PAD.n6299 PAD.n6298 0.01445
R52186 PAD.n6300 PAD.n6299 0.01445
R52187 PAD.n6300 PAD.n6199 0.01445
R52188 PAD.n6304 PAD.n6199 0.01445
R52189 PAD.n6305 PAD.n6304 0.01445
R52190 PAD.n6306 PAD.n6305 0.01445
R52191 PAD.n6306 PAD.n6197 0.01445
R52192 PAD.n6310 PAD.n6197 0.01445
R52193 PAD.n6311 PAD.n6310 0.01445
R52194 PAD.n6312 PAD.n6311 0.01445
R52195 PAD.n6312 PAD.n6195 0.01445
R52196 PAD.n6316 PAD.n6195 0.01445
R52197 PAD.n6317 PAD.n6316 0.01445
R52198 PAD.n6318 PAD.n6317 0.01445
R52199 PAD.n6318 PAD.n6193 0.01445
R52200 PAD.n6322 PAD.n6193 0.01445
R52201 PAD.n6323 PAD.n6322 0.01445
R52202 PAD.n6324 PAD.n6323 0.01445
R52203 PAD.n6324 PAD.n6191 0.01445
R52204 PAD.n6328 PAD.n6191 0.01445
R52205 PAD.n6329 PAD.n6328 0.01445
R52206 PAD.n6330 PAD.n6329 0.01445
R52207 PAD.n6330 PAD.n6189 0.01445
R52208 PAD.n6334 PAD.n6189 0.01445
R52209 PAD.n6335 PAD.n6334 0.01445
R52210 PAD.n6336 PAD.n6335 0.01445
R52211 PAD.n6336 PAD.n6187 0.01445
R52212 PAD.n6340 PAD.n6187 0.01445
R52213 PAD.n6341 PAD.n6340 0.01445
R52214 PAD.n6342 PAD.n6341 0.01445
R52215 PAD.n6342 PAD.n6185 0.01445
R52216 PAD.n6346 PAD.n6185 0.01445
R52217 PAD.n6347 PAD.n6346 0.01445
R52218 PAD.n6348 PAD.n6347 0.01445
R52219 PAD.n6348 PAD.n6183 0.01445
R52220 PAD.n6352 PAD.n6183 0.01445
R52221 PAD.n6353 PAD.n6352 0.01445
R52222 PAD.n6354 PAD.n6353 0.01445
R52223 PAD.n6354 PAD.n6181 0.01445
R52224 PAD.n6358 PAD.n6181 0.01445
R52225 PAD.n6359 PAD.n6358 0.01445
R52226 PAD.n6360 PAD.n6359 0.01445
R52227 PAD.n6360 PAD.n6179 0.01445
R52228 PAD.n6364 PAD.n6179 0.01445
R52229 PAD.n6365 PAD.n6364 0.01445
R52230 PAD.n6366 PAD.n6365 0.01445
R52231 PAD.n6366 PAD.n6177 0.01445
R52232 PAD.n6370 PAD.n6177 0.01445
R52233 PAD.n6371 PAD.n6370 0.01445
R52234 PAD.n6389 PAD.n5957 0.01445
R52235 PAD.n6225 PAD.n6224 0.01445
R52236 PAD.n6229 PAD.n6224 0.01445
R52237 PAD.n6230 PAD.n6229 0.01445
R52238 PAD.n6231 PAD.n6230 0.01445
R52239 PAD.n6231 PAD.n6222 0.01445
R52240 PAD.n6235 PAD.n6222 0.01445
R52241 PAD.n6236 PAD.n6235 0.01445
R52242 PAD.n6237 PAD.n6236 0.01445
R52243 PAD.n6237 PAD.n6220 0.01445
R52244 PAD.n6241 PAD.n6220 0.01445
R52245 PAD.n6242 PAD.n6241 0.01445
R52246 PAD.n6243 PAD.n6242 0.01445
R52247 PAD.n6243 PAD.n6218 0.01445
R52248 PAD.n6247 PAD.n6218 0.01445
R52249 PAD.n6248 PAD.n6247 0.01445
R52250 PAD.n6249 PAD.n6248 0.01445
R52251 PAD.n6249 PAD.n6216 0.01445
R52252 PAD.n6253 PAD.n6216 0.01445
R52253 PAD.n6254 PAD.n6253 0.01445
R52254 PAD.n6255 PAD.n6254 0.01445
R52255 PAD.n6255 PAD.n6214 0.01445
R52256 PAD.n6259 PAD.n6214 0.01445
R52257 PAD.n6260 PAD.n6259 0.01445
R52258 PAD.n6261 PAD.n6260 0.01445
R52259 PAD.n6261 PAD.n6212 0.01445
R52260 PAD.n6265 PAD.n6212 0.01445
R52261 PAD.n6266 PAD.n6265 0.01445
R52262 PAD.n6267 PAD.n6266 0.01445
R52263 PAD.n6267 PAD.n6210 0.01445
R52264 PAD.n6271 PAD.n6210 0.01445
R52265 PAD.n6272 PAD.n6271 0.01445
R52266 PAD.n6273 PAD.n6272 0.01445
R52267 PAD.n6273 PAD.n6208 0.01445
R52268 PAD.n6277 PAD.n6208 0.01445
R52269 PAD.n6278 PAD.n6277 0.01445
R52270 PAD.n6279 PAD.n6278 0.01445
R52271 PAD.n6279 PAD.n6206 0.01445
R52272 PAD.n6283 PAD.n6206 0.01445
R52273 PAD.n6284 PAD.n6283 0.01445
R52274 PAD.n6285 PAD.n6284 0.01445
R52275 PAD.n6285 PAD.n6204 0.01445
R52276 PAD.n6289 PAD.n6204 0.01445
R52277 PAD.n6290 PAD.n6289 0.01445
R52278 PAD.n6291 PAD.n6290 0.01445
R52279 PAD.n6291 PAD.n6202 0.01445
R52280 PAD.n6295 PAD.n6202 0.01445
R52281 PAD.n6296 PAD.n6295 0.01445
R52282 PAD.n6297 PAD.n6296 0.01445
R52283 PAD.n6297 PAD.n6200 0.01445
R52284 PAD.n6301 PAD.n6200 0.01445
R52285 PAD.n6302 PAD.n6301 0.01445
R52286 PAD.n6303 PAD.n6302 0.01445
R52287 PAD.n6303 PAD.n6198 0.01445
R52288 PAD.n6307 PAD.n6198 0.01445
R52289 PAD.n6308 PAD.n6307 0.01445
R52290 PAD.n6309 PAD.n6308 0.01445
R52291 PAD.n6309 PAD.n6196 0.01445
R52292 PAD.n6313 PAD.n6196 0.01445
R52293 PAD.n6314 PAD.n6313 0.01445
R52294 PAD.n6315 PAD.n6314 0.01445
R52295 PAD.n6315 PAD.n6194 0.01445
R52296 PAD.n6319 PAD.n6194 0.01445
R52297 PAD.n6320 PAD.n6319 0.01445
R52298 PAD.n6321 PAD.n6320 0.01445
R52299 PAD.n6321 PAD.n6192 0.01445
R52300 PAD.n6325 PAD.n6192 0.01445
R52301 PAD.n6326 PAD.n6325 0.01445
R52302 PAD.n6327 PAD.n6326 0.01445
R52303 PAD.n6327 PAD.n6190 0.01445
R52304 PAD.n6331 PAD.n6190 0.01445
R52305 PAD.n6332 PAD.n6331 0.01445
R52306 PAD.n6333 PAD.n6332 0.01445
R52307 PAD.n6333 PAD.n6188 0.01445
R52308 PAD.n6337 PAD.n6188 0.01445
R52309 PAD.n6338 PAD.n6337 0.01445
R52310 PAD.n6339 PAD.n6338 0.01445
R52311 PAD.n6339 PAD.n6186 0.01445
R52312 PAD.n6343 PAD.n6186 0.01445
R52313 PAD.n6344 PAD.n6343 0.01445
R52314 PAD.n6345 PAD.n6344 0.01445
R52315 PAD.n6345 PAD.n6184 0.01445
R52316 PAD.n6349 PAD.n6184 0.01445
R52317 PAD.n6350 PAD.n6349 0.01445
R52318 PAD.n6351 PAD.n6350 0.01445
R52319 PAD.n6351 PAD.n6182 0.01445
R52320 PAD.n6355 PAD.n6182 0.01445
R52321 PAD.n6356 PAD.n6355 0.01445
R52322 PAD.n6357 PAD.n6356 0.01445
R52323 PAD.n6357 PAD.n6180 0.01445
R52324 PAD.n6361 PAD.n6180 0.01445
R52325 PAD.n6362 PAD.n6361 0.01445
R52326 PAD.n6363 PAD.n6362 0.01445
R52327 PAD.n6363 PAD.n6178 0.01445
R52328 PAD.n6367 PAD.n6178 0.01445
R52329 PAD.n6368 PAD.n6367 0.01445
R52330 PAD.n6369 PAD.n6368 0.01445
R52331 PAD.n6369 PAD.n5978 0.01445
R52332 PAD.n6391 PAD.n6390 0.0143045
R52333 PAD.n7824 PAD.n7823 0.014225
R52334 PAD.n8435 PAD.n8434 0.014059
R52335 PAD.n4027 PAD.n3976 0.014059
R52336 PAD.n8475 PAD.n3293 0.0140338
R52337 PAD.n5899 PAD.n5896 0.0140302
R52338 PAD.n8400 PAD.n4679 0.0140302
R52339 PAD.n6681 PAD.n5901 0.0140302
R52340 PAD.n8399 PAD.n4681 0.0140302
R52341 PAD.n9156 PAD.n9155 0.013775
R52342 PAD.n10709 PAD.n10708 0.013775
R52343 PAD.n9171 PAD.n9170 0.0137632
R52344 PAD.n4328 PAD.n4323 0.013547
R52345 PAD.n4330 PAD.n4320 0.013547
R52346 PAD.n7786 PAD.n7056 0.0134925
R52347 PAD.n7815 PAD.n7814 0.0134925
R52348 PAD.n9133 PAD.n9132 0.013325
R52349 PAD.n10732 PAD.n10731 0.013325
R52350 PAD.n9196 PAD.n9195 0.0130638
R52351 PAD.n9748 PAD.n1581 0.0130638
R52352 PAD.n9189 PAD.n2035 0.0130638
R52353 PAD.n9744 PAD.n9743 0.0130638
R52354 PAD.n8835 PAD.n2888 0.0129511
R52355 PAD.n10394 PAD.n430 0.0129511
R52356 PAD.n7203 PAD.n7155 0.012875
R52357 PAD.n5958 PAD.n5955 0.0128221
R52358 PAD.n5970 PAD.n5960 0.0128221
R52359 PAD.n8474 PAD.n8473 0.0128158
R52360 PAD.n8476 PAD.n3294 0.0125805
R52361 PAD.n11536 PAD.n16 0.0125805
R52362 PAD.n8477 PAD.n3295 0.0125805
R52363 PAD.n11535 PAD.n18 0.0125805
R52364 PAD.n7822 PAD.n5199 0.0124869
R52365 PAD.n7821 PAD.n5198 0.0124869
R52366 PAD.n9147 PAD.n9146 0.0124098
R52367 PAD.n10368 PAD.n10367 0.0124098
R52368 PAD.n11538 PAD.n14 0.0124098
R52369 PAD.n11102 PAD.n11094 0.0123125
R52370 PAD.n11101 PAD.n11092 0.0123125
R52371 PAD.n5967 PAD.n5958 0.0123125
R52372 PAD.n5968 PAD.n5960 0.0123125
R52373 PAD.n7785 PAD.n7057 0.0120973
R52374 PAD.n7813 PAD.n5208 0.0120973
R52375 PAD.n7784 PAD.n7058 0.0120973
R52376 PAD.n5206 PAD.n5196 0.0120973
R52377 PAD.n9154 PAD.n2489 0.0120939
R52378 PAD.n10707 PAD.n10705 0.0120939
R52379 PAD.n9153 PAD.n2488 0.0120939
R52380 PAD.n10706 PAD.n417 0.0120939
R52381 PAD.n11505 PAD.n11499 0.011975
R52382 PAD.n6376 PAD.n5978 0.011975
R52383 PAD.n7806 PAD.n7805 0.0118684
R52384 PAD.n8190 PAD.n8189 0.0118684
R52385 PAD.n9131 PAD.n2883 0.0117009
R52386 PAD.n10730 PAD.n29 0.0117009
R52387 PAD.n9130 PAD.n2878 0.0117009
R52388 PAD.n10729 PAD.n31 0.0117009
R52389 PAD.n8834 PAD.n2889 0.0116141
R52390 PAD.n10395 PAD.n431 0.0116141
R52391 PAD.n8833 PAD.n2890 0.0116141
R52392 PAD.n10396 PAD.n432 0.0116141
R52393 PAD.n7812 PAD.n5194 0.0115977
R52394 PAD.n6378 PAD.n6377 0.011525
R52395 PAD.n8448 PAD.n3980 0.0113271
R52396 PAD.n7204 PAD.n7156 0.0113079
R52397 PAD.n7205 PAD.n7157 0.0113079
R52398 PAD.n9145 PAD.n2496 0.0111309
R52399 PAD.n1127 PAD.n1122 0.0111309
R52400 PAD.n9144 PAD.n2495 0.0111309
R52401 PAD.n1129 PAD.n1119 0.0111309
R52402 PAD.n8461 PAD.n3974 0.011075
R52403 PAD.n2034 PAD.n2032 0.0107857
R52404 PAD.n9726 PAD.n9725 0.0107857
R52405 PAD.n7804 PAD.n5547 0.0106477
R52406 PAD.n8188 PAD.n4845 0.0106477
R52407 PAD.n7803 PAD.n5549 0.0106477
R52408 PAD.n8187 PAD.n4844 0.0106477
R52409 PAD.n9736 PAD.n1589 0.010625
R52410 PAD.n10004 PAD.n1137 0.010625
R52411 PAD.n74 PAD.n18 0.0105588
R52412 PAD.n366 PAD.n31 0.0105588
R52413 PAD.n7518 PAD.n7202 0.0105588
R52414 PAD.n7269 PAD.n7157 0.0105588
R52415 PAD.n7517 PAD.n7208 0.0105588
R52416 PAD.n7270 PAD.n7156 0.0105588
R52417 PAD.n427 PAD.n415 0.0105588
R52418 PAD.n10715 PAD.n417 0.0105588
R52419 PAD.n10695 PAD.n429 0.0105588
R52420 PAD.n10705 PAD.n416 0.0105588
R52421 PAD.n523 PAD.n432 0.0105588
R52422 PAD.n770 PAD.n436 0.0105588
R52423 PAD.n522 PAD.n431 0.0105588
R52424 PAD.n771 PAD.n437 0.0105588
R52425 PAD.n824 PAD.n781 0.0105588
R52426 PAD.n10387 PAD.n827 0.0105588
R52427 PAD.n872 PAD.n780 0.0105588
R52428 PAD.n10377 PAD.n826 0.0105588
R52429 PAD.n10106 PAD.n1129 0.0105588
R52430 PAD.n10353 PAD.n1134 0.0105588
R52431 PAD.n10105 PAD.n1127 0.0105588
R52432 PAD.n10354 PAD.n1136 0.0105588
R52433 PAD.n1481 PAD.n1143 0.0105588
R52434 PAD.n1294 PAD.n1139 0.0105588
R52435 PAD.n1480 PAD.n1144 0.0105588
R52436 PAD.n1295 PAD.n1138 0.0105588
R52437 PAD.n9744 PAD.n1531 0.0105588
R52438 PAD.n9997 PAD.n1488 0.0105588
R52439 PAD.n9749 PAD.n9748 0.0105588
R52440 PAD.n1535 PAD.n1487 0.0105588
R52441 PAD.n1599 PAD.n1595 0.0105588
R52442 PAD.n1685 PAD.n1591 0.0105588
R52443 PAD.n1931 PAD.n1596 0.0105588
R52444 PAD.n1684 PAD.n1590 0.0105588
R52445 PAD.n9459 PAD.n1984 0.0105588
R52446 PAD.n9711 PAD.n1941 0.0105588
R52447 PAD.n9463 PAD.n9462 0.0105588
R52448 PAD.n1987 PAD.n1940 0.0105588
R52449 PAD.n9189 PAD.n2088 0.0105588
R52450 PAD.n9444 PAD.n2045 0.0105588
R52451 PAD.n9197 PAD.n9196 0.0105588
R52452 PAD.n2090 PAD.n2043 0.0105588
R52453 PAD.n2151 PAD.n2147 0.0105588
R52454 PAD.n2236 PAD.n2140 0.0105588
R52455 PAD.n2482 PAD.n2148 0.0105588
R52456 PAD.n2235 PAD.n2141 0.0105588
R52457 PAD.n2498 PAD.n2495 0.0105588
R52458 PAD.n2583 PAD.n2488 0.0105588
R52459 PAD.n2829 PAD.n2496 0.0105588
R52460 PAD.n2582 PAD.n2489 0.0105588
R52461 PAD.n2885 PAD.n2876 0.0105588
R52462 PAD.n9139 PAD.n2878 0.0105588
R52463 PAD.n9119 PAD.n2887 0.0105588
R52464 PAD.n2883 PAD.n2877 0.0105588
R52465 PAD.n8819 PAD.n2890 0.0105588
R52466 PAD.n8570 PAD.n2903 0.0105588
R52467 PAD.n8818 PAD.n2889 0.0105588
R52468 PAD.n8571 PAD.n2901 0.0105588
R52469 PAD.n2994 PAD.n2951 0.0105588
R52470 PAD.n8516 PAD.n2996 0.0105588
R52471 PAD.n3041 PAD.n2950 0.0105588
R52472 PAD.n8506 PAD.n2995 0.0105588
R52473 PAD.n3338 PAD.n3295 0.0105588
R52474 PAD.n8491 PAD.n3341 0.0105588
R52475 PAD.n3386 PAD.n3294 0.0105588
R52476 PAD.n3631 PAD.n3340 0.0105588
R52477 PAD.n3683 PAD.n3640 0.0105588
R52478 PAD.n8467 PAD.n3686 0.0105588
R52479 PAD.n3731 PAD.n3639 0.0105588
R52480 PAD.n8458 PAD.n3685 0.0105588
R52481 PAD.n4025 PAD.n3982 0.0105588
R52482 PAD.n8443 PAD.n4027 0.0105588
R52483 PAD.n4072 PAD.n3981 0.0105588
R52484 PAD.n8434 PAD.n4026 0.0105588
R52485 PAD.n4420 PAD.n4330 0.0105588
R52486 PAD.n4667 PAD.n4334 0.0105588
R52487 PAD.n4419 PAD.n4328 0.0105588
R52488 PAD.n4668 PAD.n4335 0.0105588
R52489 PAD.n8395 PAD.n4681 0.0105588
R52490 PAD.n8204 PAD.n4832 0.0105588
R52491 PAD.n8394 PAD.n4679 0.0105588
R52492 PAD.n4831 PAD.n4829 0.0105588
R52493 PAD.n4847 PAD.n4844 0.0105588
R52494 PAD.n4932 PAD.n4839 0.0105588
R52495 PAD.n5178 PAD.n4845 0.0105588
R52496 PAD.n4931 PAD.n4834 0.0105588
R52497 PAD.n8161 PAD.n5191 0.0105588
R52498 PAD.n7971 PAD.n5184 0.0105588
R52499 PAD.n8160 PAD.n5192 0.0105588
R52500 PAD.n7972 PAD.n5185 0.0105588
R52501 PAD.n5211 PAD.n5206 0.0105588
R52502 PAD.n5296 PAD.n5198 0.0105588
R52503 PAD.n5542 PAD.n5208 0.0105588
R52504 PAD.n5295 PAD.n5199 0.0105588
R52505 PAD.n7780 PAD.n7058 0.0105588
R52506 PAD.n7531 PAD.n7530 0.0105588
R52507 PAD.n7779 PAD.n7057 0.0105588
R52508 PAD.n7532 PAD.n7148 0.0105588
R52509 PAD.n6719 PAD.n6714 0.0105588
R52510 PAD.n6804 PAD.n6709 0.0105588
R52511 PAD.n7050 PAD.n6716 0.0105588
R52512 PAD.n6803 PAD.n6707 0.0105588
R52513 PAD.n5892 PAD.n5549 0.0105588
R52514 PAD.n5702 PAD.n5553 0.0105588
R52515 PAD.n5891 PAD.n5547 0.0105588
R52516 PAD.n5703 PAD.n5555 0.0105588
R52517 PAD.n6691 PAD.n5899 0.0105588
R52518 PAD.n6687 PAD.n6686 0.0105588
R52519 PAD.n119 PAD.n16 0.0105588
R52520 PAD.n75 PAD.n29 0.0105588
R52521 PAD.n11086 PAD.n10748 0.0105588
R52522 PAD.n10838 PAD.n10736 0.0105588
R52523 PAD.n11085 PAD.n10750 0.0105588
R52524 PAD.n10837 PAD.n10738 0.0105588
R52525 PAD.n6690 PAD.n5901 0.0105588
R52526 PAD.n6688 PAD.n5948 0.0105588
R52527 PAD.n8450 PAD.n3638 0.0102444
R52528 PAD.n11089 PAD.n11088 0.0102444
R52529 PAD.n8416 PAD.n8414 0.010175
R52530 PAD.n11505 PAD.n11504 0.010175
R52531 PAD.n8447 PAD.n3981 0.0101644
R52532 PAD.n8446 PAD.n3982 0.0101644
R52533 PAD.n6686 PAD.n5952 0.0101288
R52534 PAD.n5973 PAD.n5948 0.0101288
R52535 PAD.n8458 PAD.n8457 0.00973581
R52536 PAD.n8456 PAD.n3686 0.00973581
R52537 PAD.n7055 PAD.n7054 0.00970301
R52538 PAD.n8171 PAD.n8170 0.00970301
R52539 PAD.n11101 PAD.n11090 0.00969267
R52540 PAD.n9462 PAD.n9461 0.00968121
R52541 PAD.n9724 PAD.n1596 0.00968121
R52542 PAD.n9460 PAD.n9459 0.00968121
R52543 PAD.n9723 PAD.n1595 0.00968121
R52544 PAD.n9735 PAD.n1590 0.00934279
R52545 PAD.n10005 PAD.n1138 0.00934279
R52546 PAD.n9734 PAD.n1591 0.00934279
R52547 PAD.n10006 PAD.n1139 0.00934279
R52548 PAD.n8451 PAD.n3639 0.00919799
R52549 PAD.n10748 PAD.n10744 0.00919799
R52550 PAD.n8452 PAD.n3640 0.00919799
R52551 PAD.n10750 PAD.n10742 0.00919799
R52552 PAD.n9124 PAD.n9123 0.00916165
R52553 PAD.n10369 PAD.n779 0.00916165
R52554 PAD.n8417 PAD.n4335 0.00894978
R52555 PAD.n11503 PAD.n11303 0.00894978
R52556 PAD.n8418 PAD.n4334 0.00894978
R52557 PAD.n11502 PAD.n11253 0.00894978
R52558 PAD.n7053 PAD.n6716 0.00871477
R52559 PAD.n8172 PAD.n5192 0.00871477
R52560 PAD.n7052 PAD.n6714 0.00871477
R52561 PAD.n8173 PAD.n5191 0.00871477
R52562 PAD.n11253 PAD.n11156 0.0087125
R52563 PAD.n11498 PAD.n11303 0.0087125
R52564 PAD.n6371 PAD.n5976 0.0087125
R52565 PAD.n6372 PAD.n5972 0.0087125
R52566 PAD.n9125 PAD.n9124 0.0086203
R52567 PAD.n10392 PAD.n779 0.0086203
R52568 PAD.n8179 PAD.n8178 0.008375
R52569 PAD.n9122 PAD.n2887 0.00823154
R52570 PAD.n1123 PAD.n780 0.00823154
R52571 PAD.n9121 PAD.n2885 0.00823154
R52572 PAD.n1121 PAD.n781 0.00823154
R52573 PAD.n5967 PAD.n5956 0.00813094
R52574 PAD.n9168 PAD.n11 0.00808277
R52575 PAD.n7788 PAD.n7055 0.00807895
R52576 PAD.n8170 PAD.n8169 0.00807895
R52577 PAD.n11511 PAD.n11102 0.00796421
R52578 PAD.n11104 PAD.n11095 0.00796421
R52579 PAD.n11301 PAD.n11252 0.00796421
R52580 PAD.n11251 PAD.n11107 0.00796421
R52581 PAD.n11300 PAD.n11250 0.00796421
R52582 PAD.n11249 PAD.n11108 0.00796421
R52583 PAD.n11299 PAD.n11248 0.00796421
R52584 PAD.n11247 PAD.n11109 0.00796421
R52585 PAD.n11298 PAD.n11246 0.00796421
R52586 PAD.n11245 PAD.n11110 0.00796421
R52587 PAD.n11297 PAD.n11244 0.00796421
R52588 PAD.n11243 PAD.n11111 0.00796421
R52589 PAD.n11296 PAD.n11242 0.00796421
R52590 PAD.n11241 PAD.n11112 0.00796421
R52591 PAD.n11295 PAD.n11240 0.00796421
R52592 PAD.n11239 PAD.n11113 0.00796421
R52593 PAD.n11294 PAD.n11238 0.00796421
R52594 PAD.n11237 PAD.n11114 0.00796421
R52595 PAD.n11293 PAD.n11236 0.00796421
R52596 PAD.n11235 PAD.n11115 0.00796421
R52597 PAD.n11292 PAD.n11234 0.00796421
R52598 PAD.n11233 PAD.n11116 0.00796421
R52599 PAD.n11291 PAD.n11232 0.00796421
R52600 PAD.n11231 PAD.n11117 0.00796421
R52601 PAD.n11290 PAD.n11230 0.00796421
R52602 PAD.n11229 PAD.n11118 0.00796421
R52603 PAD.n11289 PAD.n11228 0.00796421
R52604 PAD.n11227 PAD.n11119 0.00796421
R52605 PAD.n11288 PAD.n11226 0.00796421
R52606 PAD.n11225 PAD.n11120 0.00796421
R52607 PAD.n11287 PAD.n11224 0.00796421
R52608 PAD.n11223 PAD.n11121 0.00796421
R52609 PAD.n11286 PAD.n11222 0.00796421
R52610 PAD.n11221 PAD.n11122 0.00796421
R52611 PAD.n11285 PAD.n11220 0.00796421
R52612 PAD.n11219 PAD.n11123 0.00796421
R52613 PAD.n11284 PAD.n11218 0.00796421
R52614 PAD.n11217 PAD.n11124 0.00796421
R52615 PAD.n11283 PAD.n11216 0.00796421
R52616 PAD.n11215 PAD.n11125 0.00796421
R52617 PAD.n11282 PAD.n11214 0.00796421
R52618 PAD.n11213 PAD.n11126 0.00796421
R52619 PAD.n11281 PAD.n11212 0.00796421
R52620 PAD.n11211 PAD.n11127 0.00796421
R52621 PAD.n11280 PAD.n11210 0.00796421
R52622 PAD.n11209 PAD.n11128 0.00796421
R52623 PAD.n11279 PAD.n11208 0.00796421
R52624 PAD.n11207 PAD.n11129 0.00796421
R52625 PAD.n11278 PAD.n11206 0.00796421
R52626 PAD.n11205 PAD.n11130 0.00796421
R52627 PAD.n11277 PAD.n11204 0.00796421
R52628 PAD.n11203 PAD.n11131 0.00796421
R52629 PAD.n11276 PAD.n11202 0.00796421
R52630 PAD.n11201 PAD.n11132 0.00796421
R52631 PAD.n11275 PAD.n11200 0.00796421
R52632 PAD.n11199 PAD.n11133 0.00796421
R52633 PAD.n11274 PAD.n11198 0.00796421
R52634 PAD.n11197 PAD.n11134 0.00796421
R52635 PAD.n11273 PAD.n11196 0.00796421
R52636 PAD.n11195 PAD.n11135 0.00796421
R52637 PAD.n11272 PAD.n11194 0.00796421
R52638 PAD.n11193 PAD.n11136 0.00796421
R52639 PAD.n11271 PAD.n11192 0.00796421
R52640 PAD.n11191 PAD.n11137 0.00796421
R52641 PAD.n11270 PAD.n11190 0.00796421
R52642 PAD.n11189 PAD.n11138 0.00796421
R52643 PAD.n11269 PAD.n11188 0.00796421
R52644 PAD.n11187 PAD.n11139 0.00796421
R52645 PAD.n11268 PAD.n11186 0.00796421
R52646 PAD.n11185 PAD.n11140 0.00796421
R52647 PAD.n11267 PAD.n11184 0.00796421
R52648 PAD.n11183 PAD.n11141 0.00796421
R52649 PAD.n11266 PAD.n11182 0.00796421
R52650 PAD.n11181 PAD.n11142 0.00796421
R52651 PAD.n11265 PAD.n11180 0.00796421
R52652 PAD.n11179 PAD.n11143 0.00796421
R52653 PAD.n11264 PAD.n11178 0.00796421
R52654 PAD.n11177 PAD.n11144 0.00796421
R52655 PAD.n11263 PAD.n11176 0.00796421
R52656 PAD.n11175 PAD.n11145 0.00796421
R52657 PAD.n11262 PAD.n11174 0.00796421
R52658 PAD.n11173 PAD.n11146 0.00796421
R52659 PAD.n11261 PAD.n11172 0.00796421
R52660 PAD.n11171 PAD.n11147 0.00796421
R52661 PAD.n11260 PAD.n11170 0.00796421
R52662 PAD.n11169 PAD.n11148 0.00796421
R52663 PAD.n11259 PAD.n11168 0.00796421
R52664 PAD.n11167 PAD.n11149 0.00796421
R52665 PAD.n11258 PAD.n11166 0.00796421
R52666 PAD.n11165 PAD.n11150 0.00796421
R52667 PAD.n11257 PAD.n11164 0.00796421
R52668 PAD.n11163 PAD.n11151 0.00796421
R52669 PAD.n11256 PAD.n11162 0.00796421
R52670 PAD.n11161 PAD.n11152 0.00796421
R52671 PAD.n11255 PAD.n11160 0.00796421
R52672 PAD.n11159 PAD.n11153 0.00796421
R52673 PAD.n11254 PAD.n11158 0.00796421
R52674 PAD.n11157 PAD.n11154 0.00796421
R52675 PAD.n11156 PAD.n11155 0.00796421
R52676 PAD.n6384 PAD.n5968 0.00796421
R52677 PAD.n5969 PAD.n5961 0.00796421
R52678 PAD.n6033 PAD.n6030 0.00796421
R52679 PAD.n6037 PAD.n6035 0.00796421
R52680 PAD.n6036 PAD.n6029 0.00796421
R52681 PAD.n6040 PAD.n6038 0.00796421
R52682 PAD.n6039 PAD.n6028 0.00796421
R52683 PAD.n6043 PAD.n6041 0.00796421
R52684 PAD.n6042 PAD.n6027 0.00796421
R52685 PAD.n6046 PAD.n6044 0.00796421
R52686 PAD.n6045 PAD.n6026 0.00796421
R52687 PAD.n6049 PAD.n6047 0.00796421
R52688 PAD.n6048 PAD.n6025 0.00796421
R52689 PAD.n6052 PAD.n6050 0.00796421
R52690 PAD.n6051 PAD.n6024 0.00796421
R52691 PAD.n6055 PAD.n6053 0.00796421
R52692 PAD.n6054 PAD.n6023 0.00796421
R52693 PAD.n6058 PAD.n6056 0.00796421
R52694 PAD.n6057 PAD.n6022 0.00796421
R52695 PAD.n6061 PAD.n6059 0.00796421
R52696 PAD.n6060 PAD.n6021 0.00796421
R52697 PAD.n6064 PAD.n6062 0.00796421
R52698 PAD.n6063 PAD.n6020 0.00796421
R52699 PAD.n6067 PAD.n6065 0.00796421
R52700 PAD.n6066 PAD.n6019 0.00796421
R52701 PAD.n6070 PAD.n6068 0.00796421
R52702 PAD.n6069 PAD.n6018 0.00796421
R52703 PAD.n6073 PAD.n6071 0.00796421
R52704 PAD.n6072 PAD.n6017 0.00796421
R52705 PAD.n6076 PAD.n6074 0.00796421
R52706 PAD.n6075 PAD.n6016 0.00796421
R52707 PAD.n6079 PAD.n6077 0.00796421
R52708 PAD.n6078 PAD.n6015 0.00796421
R52709 PAD.n6082 PAD.n6080 0.00796421
R52710 PAD.n6081 PAD.n6014 0.00796421
R52711 PAD.n6085 PAD.n6083 0.00796421
R52712 PAD.n6084 PAD.n6013 0.00796421
R52713 PAD.n6088 PAD.n6086 0.00796421
R52714 PAD.n6087 PAD.n6012 0.00796421
R52715 PAD.n6091 PAD.n6089 0.00796421
R52716 PAD.n6090 PAD.n6011 0.00796421
R52717 PAD.n6094 PAD.n6092 0.00796421
R52718 PAD.n6093 PAD.n6010 0.00796421
R52719 PAD.n6097 PAD.n6095 0.00796421
R52720 PAD.n6096 PAD.n6009 0.00796421
R52721 PAD.n6100 PAD.n6098 0.00796421
R52722 PAD.n6099 PAD.n6008 0.00796421
R52723 PAD.n6103 PAD.n6101 0.00796421
R52724 PAD.n6102 PAD.n6007 0.00796421
R52725 PAD.n6106 PAD.n6104 0.00796421
R52726 PAD.n6105 PAD.n6006 0.00796421
R52727 PAD.n6109 PAD.n6107 0.00796421
R52728 PAD.n6108 PAD.n6005 0.00796421
R52729 PAD.n6112 PAD.n6110 0.00796421
R52730 PAD.n6111 PAD.n6004 0.00796421
R52731 PAD.n6115 PAD.n6113 0.00796421
R52732 PAD.n6114 PAD.n6003 0.00796421
R52733 PAD.n6118 PAD.n6116 0.00796421
R52734 PAD.n6117 PAD.n6002 0.00796421
R52735 PAD.n6121 PAD.n6119 0.00796421
R52736 PAD.n6120 PAD.n6001 0.00796421
R52737 PAD.n6124 PAD.n6122 0.00796421
R52738 PAD.n6123 PAD.n6000 0.00796421
R52739 PAD.n6127 PAD.n6125 0.00796421
R52740 PAD.n6126 PAD.n5999 0.00796421
R52741 PAD.n6130 PAD.n6128 0.00796421
R52742 PAD.n6129 PAD.n5998 0.00796421
R52743 PAD.n6133 PAD.n6131 0.00796421
R52744 PAD.n6132 PAD.n5997 0.00796421
R52745 PAD.n6136 PAD.n6134 0.00796421
R52746 PAD.n6135 PAD.n5996 0.00796421
R52747 PAD.n6139 PAD.n6137 0.00796421
R52748 PAD.n6138 PAD.n5995 0.00796421
R52749 PAD.n6142 PAD.n6140 0.00796421
R52750 PAD.n6141 PAD.n5994 0.00796421
R52751 PAD.n6145 PAD.n6143 0.00796421
R52752 PAD.n6144 PAD.n5993 0.00796421
R52753 PAD.n6148 PAD.n6146 0.00796421
R52754 PAD.n6147 PAD.n5992 0.00796421
R52755 PAD.n6151 PAD.n6149 0.00796421
R52756 PAD.n6150 PAD.n5991 0.00796421
R52757 PAD.n6154 PAD.n6152 0.00796421
R52758 PAD.n6153 PAD.n5990 0.00796421
R52759 PAD.n6157 PAD.n6155 0.00796421
R52760 PAD.n6156 PAD.n5989 0.00796421
R52761 PAD.n6160 PAD.n6158 0.00796421
R52762 PAD.n6159 PAD.n5988 0.00796421
R52763 PAD.n6163 PAD.n6161 0.00796421
R52764 PAD.n6162 PAD.n5987 0.00796421
R52765 PAD.n6166 PAD.n6164 0.00796421
R52766 PAD.n6165 PAD.n5986 0.00796421
R52767 PAD.n6169 PAD.n6167 0.00796421
R52768 PAD.n6168 PAD.n5985 0.00796421
R52769 PAD.n6172 PAD.n6170 0.00796421
R52770 PAD.n6171 PAD.n5984 0.00796421
R52771 PAD.n6175 PAD.n6173 0.00796421
R52772 PAD.n6174 PAD.n5983 0.00796421
R52773 PAD.n6032 PAD.n6031 0.00796421
R52774 PAD.n6372 PAD.n6176 0.00796421
R52775 PAD.n6176 PAD.n6032 0.00796421
R52776 PAD.n11155 PAD.n11154 0.00796421
R52777 PAD.n11158 PAD.n11157 0.00796421
R52778 PAD.n11254 PAD.n11153 0.00796421
R52779 PAD.n11160 PAD.n11159 0.00796421
R52780 PAD.n11255 PAD.n11152 0.00796421
R52781 PAD.n11162 PAD.n11161 0.00796421
R52782 PAD.n11256 PAD.n11151 0.00796421
R52783 PAD.n11164 PAD.n11163 0.00796421
R52784 PAD.n11257 PAD.n11150 0.00796421
R52785 PAD.n11166 PAD.n11165 0.00796421
R52786 PAD.n11258 PAD.n11149 0.00796421
R52787 PAD.n11168 PAD.n11167 0.00796421
R52788 PAD.n11259 PAD.n11148 0.00796421
R52789 PAD.n11170 PAD.n11169 0.00796421
R52790 PAD.n11260 PAD.n11147 0.00796421
R52791 PAD.n11172 PAD.n11171 0.00796421
R52792 PAD.n11261 PAD.n11146 0.00796421
R52793 PAD.n11174 PAD.n11173 0.00796421
R52794 PAD.n11262 PAD.n11145 0.00796421
R52795 PAD.n11176 PAD.n11175 0.00796421
R52796 PAD.n11263 PAD.n11144 0.00796421
R52797 PAD.n11178 PAD.n11177 0.00796421
R52798 PAD.n11264 PAD.n11143 0.00796421
R52799 PAD.n11180 PAD.n11179 0.00796421
R52800 PAD.n11265 PAD.n11142 0.00796421
R52801 PAD.n11182 PAD.n11181 0.00796421
R52802 PAD.n11266 PAD.n11141 0.00796421
R52803 PAD.n11184 PAD.n11183 0.00796421
R52804 PAD.n11267 PAD.n11140 0.00796421
R52805 PAD.n11186 PAD.n11185 0.00796421
R52806 PAD.n11268 PAD.n11139 0.00796421
R52807 PAD.n11188 PAD.n11187 0.00796421
R52808 PAD.n11269 PAD.n11138 0.00796421
R52809 PAD.n11190 PAD.n11189 0.00796421
R52810 PAD.n11270 PAD.n11137 0.00796421
R52811 PAD.n11192 PAD.n11191 0.00796421
R52812 PAD.n11271 PAD.n11136 0.00796421
R52813 PAD.n11194 PAD.n11193 0.00796421
R52814 PAD.n11272 PAD.n11135 0.00796421
R52815 PAD.n11196 PAD.n11195 0.00796421
R52816 PAD.n11273 PAD.n11134 0.00796421
R52817 PAD.n11198 PAD.n11197 0.00796421
R52818 PAD.n11274 PAD.n11133 0.00796421
R52819 PAD.n11200 PAD.n11199 0.00796421
R52820 PAD.n11275 PAD.n11132 0.00796421
R52821 PAD.n11202 PAD.n11201 0.00796421
R52822 PAD.n11276 PAD.n11131 0.00796421
R52823 PAD.n11204 PAD.n11203 0.00796421
R52824 PAD.n11277 PAD.n11130 0.00796421
R52825 PAD.n11206 PAD.n11205 0.00796421
R52826 PAD.n11278 PAD.n11129 0.00796421
R52827 PAD.n11208 PAD.n11207 0.00796421
R52828 PAD.n11279 PAD.n11128 0.00796421
R52829 PAD.n11210 PAD.n11209 0.00796421
R52830 PAD.n11280 PAD.n11127 0.00796421
R52831 PAD.n11212 PAD.n11211 0.00796421
R52832 PAD.n11281 PAD.n11126 0.00796421
R52833 PAD.n11214 PAD.n11213 0.00796421
R52834 PAD.n11282 PAD.n11125 0.00796421
R52835 PAD.n11216 PAD.n11215 0.00796421
R52836 PAD.n11283 PAD.n11124 0.00796421
R52837 PAD.n11218 PAD.n11217 0.00796421
R52838 PAD.n11284 PAD.n11123 0.00796421
R52839 PAD.n11220 PAD.n11219 0.00796421
R52840 PAD.n11285 PAD.n11122 0.00796421
R52841 PAD.n11222 PAD.n11221 0.00796421
R52842 PAD.n11286 PAD.n11121 0.00796421
R52843 PAD.n11224 PAD.n11223 0.00796421
R52844 PAD.n11287 PAD.n11120 0.00796421
R52845 PAD.n11226 PAD.n11225 0.00796421
R52846 PAD.n11288 PAD.n11119 0.00796421
R52847 PAD.n11228 PAD.n11227 0.00796421
R52848 PAD.n11289 PAD.n11118 0.00796421
R52849 PAD.n11230 PAD.n11229 0.00796421
R52850 PAD.n11290 PAD.n11117 0.00796421
R52851 PAD.n11232 PAD.n11231 0.00796421
R52852 PAD.n11291 PAD.n11116 0.00796421
R52853 PAD.n11234 PAD.n11233 0.00796421
R52854 PAD.n11292 PAD.n11115 0.00796421
R52855 PAD.n11236 PAD.n11235 0.00796421
R52856 PAD.n11293 PAD.n11114 0.00796421
R52857 PAD.n11238 PAD.n11237 0.00796421
R52858 PAD.n11294 PAD.n11113 0.00796421
R52859 PAD.n11240 PAD.n11239 0.00796421
R52860 PAD.n11295 PAD.n11112 0.00796421
R52861 PAD.n11242 PAD.n11241 0.00796421
R52862 PAD.n11296 PAD.n11111 0.00796421
R52863 PAD.n11244 PAD.n11243 0.00796421
R52864 PAD.n11297 PAD.n11110 0.00796421
R52865 PAD.n11246 PAD.n11245 0.00796421
R52866 PAD.n11298 PAD.n11109 0.00796421
R52867 PAD.n11248 PAD.n11247 0.00796421
R52868 PAD.n11299 PAD.n11108 0.00796421
R52869 PAD.n11250 PAD.n11249 0.00796421
R52870 PAD.n11300 PAD.n11107 0.00796421
R52871 PAD.n11252 PAD.n11251 0.00796421
R52872 PAD.n11301 PAD.n11106 0.00796421
R52873 PAD.n6387 PAD.n5961 0.00796421
R52874 PAD.n11514 PAD.n11095 0.00796421
R52875 PAD.n6385 PAD.n6384 0.00796421
R52876 PAD.n11512 PAD.n11511 0.00796421
R52877 PAD.n6034 PAD.n6033 0.00796421
R52878 PAD.n6035 PAD.n6030 0.00796421
R52879 PAD.n6037 PAD.n6036 0.00796421
R52880 PAD.n6038 PAD.n6029 0.00796421
R52881 PAD.n6040 PAD.n6039 0.00796421
R52882 PAD.n6041 PAD.n6028 0.00796421
R52883 PAD.n6043 PAD.n6042 0.00796421
R52884 PAD.n6044 PAD.n6027 0.00796421
R52885 PAD.n6046 PAD.n6045 0.00796421
R52886 PAD.n6047 PAD.n6026 0.00796421
R52887 PAD.n6049 PAD.n6048 0.00796421
R52888 PAD.n6050 PAD.n6025 0.00796421
R52889 PAD.n6052 PAD.n6051 0.00796421
R52890 PAD.n6053 PAD.n6024 0.00796421
R52891 PAD.n6055 PAD.n6054 0.00796421
R52892 PAD.n6056 PAD.n6023 0.00796421
R52893 PAD.n6058 PAD.n6057 0.00796421
R52894 PAD.n6059 PAD.n6022 0.00796421
R52895 PAD.n6061 PAD.n6060 0.00796421
R52896 PAD.n6062 PAD.n6021 0.00796421
R52897 PAD.n6064 PAD.n6063 0.00796421
R52898 PAD.n6065 PAD.n6020 0.00796421
R52899 PAD.n6067 PAD.n6066 0.00796421
R52900 PAD.n6068 PAD.n6019 0.00796421
R52901 PAD.n6070 PAD.n6069 0.00796421
R52902 PAD.n6071 PAD.n6018 0.00796421
R52903 PAD.n6073 PAD.n6072 0.00796421
R52904 PAD.n6074 PAD.n6017 0.00796421
R52905 PAD.n6076 PAD.n6075 0.00796421
R52906 PAD.n6077 PAD.n6016 0.00796421
R52907 PAD.n6079 PAD.n6078 0.00796421
R52908 PAD.n6080 PAD.n6015 0.00796421
R52909 PAD.n6082 PAD.n6081 0.00796421
R52910 PAD.n6083 PAD.n6014 0.00796421
R52911 PAD.n6085 PAD.n6084 0.00796421
R52912 PAD.n6086 PAD.n6013 0.00796421
R52913 PAD.n6088 PAD.n6087 0.00796421
R52914 PAD.n6089 PAD.n6012 0.00796421
R52915 PAD.n6091 PAD.n6090 0.00796421
R52916 PAD.n6092 PAD.n6011 0.00796421
R52917 PAD.n6094 PAD.n6093 0.00796421
R52918 PAD.n6095 PAD.n6010 0.00796421
R52919 PAD.n6097 PAD.n6096 0.00796421
R52920 PAD.n6098 PAD.n6009 0.00796421
R52921 PAD.n6100 PAD.n6099 0.00796421
R52922 PAD.n6101 PAD.n6008 0.00796421
R52923 PAD.n6103 PAD.n6102 0.00796421
R52924 PAD.n6104 PAD.n6007 0.00796421
R52925 PAD.n6106 PAD.n6105 0.00796421
R52926 PAD.n6107 PAD.n6006 0.00796421
R52927 PAD.n6109 PAD.n6108 0.00796421
R52928 PAD.n6110 PAD.n6005 0.00796421
R52929 PAD.n6112 PAD.n6111 0.00796421
R52930 PAD.n6113 PAD.n6004 0.00796421
R52931 PAD.n6115 PAD.n6114 0.00796421
R52932 PAD.n6116 PAD.n6003 0.00796421
R52933 PAD.n6118 PAD.n6117 0.00796421
R52934 PAD.n6119 PAD.n6002 0.00796421
R52935 PAD.n6121 PAD.n6120 0.00796421
R52936 PAD.n6122 PAD.n6001 0.00796421
R52937 PAD.n6124 PAD.n6123 0.00796421
R52938 PAD.n6125 PAD.n6000 0.00796421
R52939 PAD.n6127 PAD.n6126 0.00796421
R52940 PAD.n6128 PAD.n5999 0.00796421
R52941 PAD.n6130 PAD.n6129 0.00796421
R52942 PAD.n6131 PAD.n5998 0.00796421
R52943 PAD.n6133 PAD.n6132 0.00796421
R52944 PAD.n6134 PAD.n5997 0.00796421
R52945 PAD.n6136 PAD.n6135 0.00796421
R52946 PAD.n6137 PAD.n5996 0.00796421
R52947 PAD.n6139 PAD.n6138 0.00796421
R52948 PAD.n6140 PAD.n5995 0.00796421
R52949 PAD.n6142 PAD.n6141 0.00796421
R52950 PAD.n6143 PAD.n5994 0.00796421
R52951 PAD.n6145 PAD.n6144 0.00796421
R52952 PAD.n6146 PAD.n5993 0.00796421
R52953 PAD.n6148 PAD.n6147 0.00796421
R52954 PAD.n6149 PAD.n5992 0.00796421
R52955 PAD.n6151 PAD.n6150 0.00796421
R52956 PAD.n6152 PAD.n5991 0.00796421
R52957 PAD.n6154 PAD.n6153 0.00796421
R52958 PAD.n6155 PAD.n5990 0.00796421
R52959 PAD.n6157 PAD.n6156 0.00796421
R52960 PAD.n6158 PAD.n5989 0.00796421
R52961 PAD.n6160 PAD.n6159 0.00796421
R52962 PAD.n6161 PAD.n5988 0.00796421
R52963 PAD.n6163 PAD.n6162 0.00796421
R52964 PAD.n6164 PAD.n5987 0.00796421
R52965 PAD.n6166 PAD.n6165 0.00796421
R52966 PAD.n6167 PAD.n5986 0.00796421
R52967 PAD.n6169 PAD.n6168 0.00796421
R52968 PAD.n6170 PAD.n5985 0.00796421
R52969 PAD.n6172 PAD.n6171 0.00796421
R52970 PAD.n6173 PAD.n5984 0.00796421
R52971 PAD.n6175 PAD.n6174 0.00796421
R52972 PAD.n6031 PAD.n5983 0.00796421
R52973 PAD.n9180 PAD.n9179 0.007925
R52974 PAD.n10404 PAD.n10402 0.007925
R52975 PAD.n9126 PAD.n2887 0.00774832
R52976 PAD.n10391 PAD.n780 0.00774832
R52977 PAD.n9127 PAD.n2885 0.00774832
R52978 PAD.n10390 PAD.n781 0.00774832
R52979 PAD.n8472 PAD.n3638 0.00753759
R52980 PAD.n11088 PAD.n10746 0.00753759
R52981 PAD.n8827 PAD.n8826 0.007475
R52982 PAD.n11528 PAD.n11527 0.007475
R52983 PAD.n8177 PAD.n5185 0.00737773
R52984 PAD.n8176 PAD.n5184 0.00737773
R52985 PAD.n7789 PAD.n6716 0.0072651
R52986 PAD.n8168 PAD.n5192 0.0072651
R52987 PAD.n7790 PAD.n6714 0.0072651
R52988 PAD.n8167 PAD.n5191 0.0072651
R52989 PAD.n11517 PAD.n11516 0.0071375
R52990 PAD.n6390 PAD.n6389 0.0071375
R52991 PAD.n6380 PAD.n6376 0.007025
R52992 PAD.n7526 PAD.n7154 0.007025
R52993 PAD.n9192 PAD.n2032 0.00699624
R52994 PAD.n9729 PAD.n9726 0.00699624
R52995 PAD.n3637 PAD.n3636 0.0069926
R52996 PAD.n9178 PAD.n2141 0.00698472
R52997 PAD.n10405 PAD.n437 0.00698472
R52998 PAD.n9177 PAD.n2140 0.00698472
R52999 PAD.n10406 PAD.n436 0.00698472
R53000 PAD.n8471 PAD.n3639 0.00678188
R53001 PAD.n10751 PAD.n10748 0.00678188
R53002 PAD.n8470 PAD.n3640 0.00678188
R53003 PAD.n10752 PAD.n10750 0.00678188
R53004 PAD.n2901 PAD.n2896 0.0065917
R53005 PAD.n10736 PAD.n25 0.0065917
R53006 PAD.n2903 PAD.n2893 0.0065917
R53007 PAD.n10738 PAD.n23 0.0065917
R53008 PAD.n8426 PAD.n3980 0.00645489
R53009 PAD.n9462 PAD.n2033 0.00629866
R53010 PAD.n9730 PAD.n1596 0.00629866
R53011 PAD.n9459 PAD.n9458 0.00629866
R53012 PAD.n9731 PAD.n1595 0.00629866
R53013 PAD.n11508 PAD.n11253 0.0062375
R53014 PAD.n11506 PAD.n11303 0.0062375
R53015 PAD.n6375 PAD.n5976 0.0062375
R53016 PAD.n6374 PAD.n5972 0.0062375
R53017 PAD.n6381 PAD.n5976 0.00619869
R53018 PAD.n7527 PAD.n7148 0.00619869
R53019 PAD.n6382 PAD.n5972 0.00619869
R53020 PAD.n7530 PAD.n7529 0.00619869
R53021 PAD.n7814 PAD.n7812 0.00618421
R53022 PAD.n8191 PAD.n8190 0.00591353
R53023 PAD.n4324 PAD.n3981 0.00581544
R53024 PAD.n4322 PAD.n3982 0.00581544
R53025 PAD.n6704 PAD.n6703 0.005675
R53026 PAD.n9148 PAD.n9147 0.00537218
R53027 PAD.n6697 PAD.n5547 0.00533221
R53028 PAD.n8192 PAD.n4845 0.00533221
R53029 PAD.n6698 PAD.n5549 0.00533221
R53030 PAD.n8193 PAD.n4844 0.00533221
R53031 PAD.n8485 PAD.n8483 0.005225
R53032 PAD.n6702 PAD.n5555 0.00501965
R53033 PAD.n6701 PAD.n5553 0.00501965
R53034 PAD.n8473 PAD.n8472 0.00496617
R53035 PAD.n9149 PAD.n2496 0.00484899
R53036 PAD.n10364 PAD.n1127 0.00484899
R53037 PAD.n9150 PAD.n2495 0.00484899
R53038 PAD.n10363 PAD.n1129 0.00484899
R53039 PAD.n8524 PAD.n2888 0.00483083
R53040 PAD.n10411 PAD.n430 0.00483083
R53041 PAD.n9716 PAD.n1939 0.004775
R53042 PAD.n10358 PAD.n10357 0.004775
R53043 PAD.n8482 PAD.n3631 0.00462664
R53044 PAD.n8481 PAD.n3341 0.00462664
R53045 PAD.n8525 PAD.n2889 0.00436577
R53046 PAD.n10410 PAD.n431 0.00436577
R53047 PAD.n8526 PAD.n2890 0.00436577
R53048 PAD.n10409 PAD.n432 0.00436577
R53049 PAD.n8209 PAD.n8208 0.004325
R53050 PAD.n7212 PAD.n7056 0.00428947
R53051 PAD.n7816 PAD.n7815 0.00428947
R53052 PAD.n9715 PAD.n1940 0.00423362
R53053 PAD.n10359 PAD.n1136 0.00423362
R53054 PAD.n9714 PAD.n1941 0.00423362
R53055 PAD.n10360 PAD.n1134 0.00423362
R53056 PAD.n9172 PAD.n9171 0.0040188
R53057 PAD.n7213 PAD.n7057 0.00388255
R53058 PAD.n7817 PAD.n5208 0.00388255
R53059 PAD.n7214 PAD.n7058 0.00388255
R53060 PAD.n7818 PAD.n5206 0.00388255
R53061 PAD.n8207 PAD.n4831 0.00384061
R53062 PAD.n8206 PAD.n8204 0.00384061
R53063 PAD.n8496 PAD.n3293 0.00374812
R53064 PAD.n10724 PAD.n14 0.00374812
R53065 PAD.n7807 PAD.n7806 0.00347744
R53066 PAD.n8495 PAD.n3294 0.00339933
R53067 PAD.n10725 PAD.n16 0.00339933
R53068 PAD.n8494 PAD.n3295 0.00339933
R53069 PAD.n10726 PAD.n18 0.00339933
R53070 PAD.n2137 PAD.n2135 0.00320677
R53071 PAD.n1584 PAD.n1580 0.00320677
R53072 PAD.n7807 PAD.n5544 0.00293609
R53073 PAD.n10366 PAD.n10365 0.00293609
R53074 PAD.n10367 PAD.n10366 0.00293609
R53075 PAD.n9196 PAD.n9191 0.00291611
R53076 PAD.n9748 PAD.n9747 0.00291611
R53077 PAD.n9190 PAD.n9189 0.00291611
R53078 PAD.n9746 PAD.n9744 0.00291611
R53079 PAD.n8424 PAD.n8423 0.00266541
R53080 PAD.n11514 PAD.n11094 0.0026375
R53081 PAD.n11515 PAD.n11092 0.0026375
R53082 PAD.n6388 PAD.n5958 0.0026375
R53083 PAD.n6387 PAD.n5960 0.0026375
R53084 PAD.n8199 PAD.n8198 0.002525
R53085 PAD.n8422 PAD.n4328 0.00243289
R53086 PAD.n8421 PAD.n4330 0.00243289
R53087 PAD.n8197 PAD.n4834 0.00226856
R53088 PAD.n8196 PAD.n4839 0.00226856
R53089 PAD.n6693 PAD.n5897 0.00212406
R53090 PAD.n8403 PAD.n8402 0.00212406
R53091 PAD.n11538 PAD.n11537 0.00212406
R53092 PAD.n9450 PAD.n9449 0.002075
R53093 PAD.n10381 PAD.n10380 0.002075
R53094 PAD.n6394 PAD.n5899 0.00194966
R53095 PAD.n4679 PAD.n4675 0.00194966
R53096 PAD.n6395 PAD.n5901 0.00194966
R53097 PAD.n4681 PAD.n4674 0.00194966
R53098 PAD.n9448 PAD.n2043 0.00187555
R53099 PAD.n10379 PAD.n10377 0.00187555
R53100 PAD.n9447 PAD.n2045 0.00187555
R53101 PAD.n10378 PAD.n827 0.00187555
R53102 PAD.n8510 PAD.n8509 0.001625
R53103 PAD.n9172 PAD.n9167 0.00158271
R53104 PAD.n10012 PAD.n10011 0.00158271
R53105 PAD.n8508 PAD.n8506 0.00148253
R53106 PAD.n8507 PAD.n2996 0.00148253
R53107 PAD.n9173 PAD.n2148 0.00146644
R53108 PAD.n10010 PAD.n1144 0.00146644
R53109 PAD.n9174 PAD.n2147 0.00146644
R53110 PAD.n10009 PAD.n1143 0.00146644
R53111 PAD.n11103 PAD.n11097 0.00128471
R53112 PAD.n11103 PAD.n11098 0.00128471
R53113 PAD.n7796 PAD.n7795 0.001175
R53114 PAD.n7794 PAD.n6707 0.00108952
R53115 PAD.n7793 PAD.n6709 0.00108952
R53116 PAD.n6386 PAD.n5966 0.00106946
R53117 PAD.n8165 PAD.n7829 0.00106946
R53118 PAD.n8445 PAD.n3977 0.00106946
R53119 PAD.n11534 PAD.n11533 0.00106946
R53120 PAD.n6682 PAD.n6680 0.00106487
R53121 PAD.n10016 PAD.n1142 0.00106487
R53122 PAD.n9186 PAD.n9185 0.0010465
R53123 PAD.n8498 PAD.n2949 0.00104135
R53124 PAD.n10697 PAD.n370 0.00104135
R53125 PAD.n8454 PAD.n8453 0.00103731
R53126 PAD.n9129 PAD.n9128 0.00103731
R53127 PAD.n5982 PAD.n5963 0.00103272
R53128 PAD.n5981 PAD.n5964 0.00103272
R53129 PAD.n5980 PAD.n5962 0.00103272
R53130 PAD.n5979 PAD.n5965 0.00103272
R53131 PAD.n8503 PAD.n3287 0.00102813
R53132 PAD.n9141 PAD.n9140 0.00102813
R53133 PAD.n4321 PAD.n3983 0.00101894
R53134 PAD.n9143 PAD.n9142 0.00101894
R53135 PAD.n4841 PAD.n4682 0.00100976
R53136 PAD.n9733 PAD.n1592 0.00100517
R53137 PAD.n9742 PAD.n1586 0.00100057
R53138 PAD.n7061 PAD.n7060 0.000991389
R53139 PAD.n8164 PAD.n8163 0.000991389
R53140 PAD.n10398 PAD.n776 0.000991389
R53141 PAD.n3292 PAD.n2950 0.000983221
R53142 PAD.n429 PAD.n371 0.000983221
R53143 PAD.n3290 PAD.n2951 0.000983221
R53144 PAD.n427 PAD.n372 0.000983221
R53145 PAD.n7215 PAD.n7158 0.000982204
R53146 PAD.n10701 PAD.n425 0.000982204
R53147 PAD.n7819 PAD.n5197 0.000977612
R53148 PAD.n8175 PAD.n8174 0.00097302
R53149 PAD.n9721 PAD.n1936 0.00097302
R53150 PAD.n10408 PAD.n433 0.00097302
R53151 PAD.n8409 PAD.n8408 0.000963835
R53152 PAD.n11532 PAD.n21 0.000959242
R53153 PAD.n10755 PAD.n10754 0.000959242
R53154 PAD.n8469 PAD.n3641 0.00095465
R53155 PAD.n2894 PAD.n2892 0.00095465
R53156 PAD.n6700 PAD.n5551 0.000945465
R53157 PAD.n8518 PAD.n2904 0.000945465
R53158 PAD.n6679 PAD.n5894 0.000940873
R53159 PAD.n8431 PAD.n8430 0.00093628
R53160 PAD.n9152 PAD.n9151 0.00093628
R53161 PAD.n1594 PAD.n1593 0.00093628
R53162 PAD.n9456 PAD.n2037 0.000927095
R53163 PAD.n10727 PAD.n367 0.000922503
R53164 PAD.n11507 PAD.n11096 0.000922503
R53165 PAD.n11302 PAD.n11099 0.000922503
R53166 PAD.n11510 PAD.n11509 0.000922503
R53167 PAD.n11513 PAD.n11100 0.000922503
R53168 PAD.n7782 PAD.n7103 0.00091791
R53169 PAD.n7801 PAD.n5552 0.000908726
R53170 PAD.n10361 PAD.n1132 0.000908726
R53171 PAD.n10373 PAD.n1118 0.000908726
R53172 PAD.n1536 PAD.n1489 0.000904133
R53173 PAD.n1141 PAD.n1130 0.000904133
R53174 PAD.n7221 PAD.n5204 0.000894948
R53175 PAD.n8184 PAD.n8183 0.000890356
R53176 PAD.n1986 PAD.n1985 0.000890356
R53177 PAD.n435 PAD.n434 0.000890356
R53178 PAD.n11523 PAD.n11522 0.000890356
R53179 PAD.n10008 PAD.n1140 0.000876579
R53180 PAD.n6678 PAD.n6396 0.000871986
R53181 PAD.n8397 PAD.n4724 0.000871986
R53182 PAD.n3684 PAD.n3633 0.000871986
R53183 PAD.n8832 PAD.n8831 0.000871986
R53184 PAD.n9446 PAD.n9445 0.000862801
R53185 PAD.n419 PAD.n418 0.000858209
R53186 PAD.n4332 PAD.n4319 0.000853617
R53187 PAD.n9161 PAD.n9160 0.000853617
R53188 PAD.n10388 PAD.n825 0.000844432
R53189 PAD.n11501 PAD.n11500 0.000844432
R53190 PAD.n9187 PAD.n2091 0.000839839
R53191 PAD.n10717 PAD.n32 0.000839839
R53192 PAD.n6383 PAD.n5971 0.000835247
R53193 PAD.n7216 PAD.n7105 0.000835247
R53194 PAD.n7223 PAD.n7222 0.000835247
R53195 PAD.n10719 PAD.n10718 0.000835247
R53196 PAD.n6712 PAD.n6711 0.000826062
R53197 PAD.n7792 PAD.n6712 0.000826062
R53198 PAD.n7059 PAD.n6713 0.000826062
R53199 PAD.n1120 PAD.n782 0.000826062
R53200 PAD.n3289 PAD.n2997 0.00082147
R53201 PAD.n9998 PAD.n1534 0.00082147
R53202 PAD.n5974 PAD.n5971 0.000816877
R53203 PAD.n1534 PAD.n1533 0.000816877
R53204 PAD.n8186 PAD.n8185 0.000807692
R53205 PAD.n9713 PAD.n1942 0.000807692
R53206 PAD.n10374 PAD.n828 0.000807692
R53207 PAD.n11500 PAD.n10741 0.000807692
R53208 PAD.n7520 PAD.n7200 0.0008031
R53209 PAD.n9162 PAD.n9161 0.000798507
R53210 PAD.n1532 PAD.n1483 0.000793915
R53211 PAD.n6689 PAD.n5903 0.000789323
R53212 PAD.n8407 PAD.n4673 0.000789323
R53213 PAD.n8479 PAD.n8478 0.000789323
R53214 PAD.n8517 PAD.n2952 0.000789323
R53215 PAD.n8479 PAD.n3633 0.000780138
R53216 PAD.n10719 PAD.n10716 0.000775545
R53217 PAD.n8420 PAD.n8419 0.000770953
R53218 PAD.n9163 PAD.n9162 0.000770953
R53219 PAD.n9175 PAD.n2139 0.000770953
R53220 PAD.n8185 PAD.n8184 0.000761768
R53221 PAD.n8195 PAD.n4840 0.000761768
R53222 PAD.n4843 PAD.n4842 0.000761768
R53223 PAD.n11522 PAD.n10741 0.000761768
R53224 PAD.n8205 PAD.n4673 0.000757176
R53225 PAD.n8420 PAD.n4331 0.000757176
R53226 PAD.n3342 PAD.n3296 0.000757176
R53227 PAD.n8492 PAD.n3339 0.000757176
R53228 PAD.n5974 PAD.n5903 0.000752583
R53229 PAD.n7206 PAD.n7200 0.000752583
R53230 PAD.n1533 PAD.n1532 0.000752583
R53231 PAD.n418 PAD.n373 0.000752583
R53232 PAD.n8502 PAD.n2997 0.000747991
R53233 PAD.n6711 PAD.n5552 0.000743398
R53234 PAD.n7792 PAD.n7791 0.000743398
R53235 PAD.n9455 PAD.n1988 0.000743398
R53236 PAD.n9713 PAD.n9712 0.000743398
R53237 PAD.n10374 PAD.n10373 0.000743398
R53238 PAD.n10389 PAD.n782 0.000743398
R53239 PAD.n8519 PAD.n8517 0.000738806
R53240 PAD.n6386 PAD.n6383 0.000734214
R53241 PAD.n7222 PAD.n7221 0.000734214
R53242 PAD.n9999 PAD.n1489 0.000734214
R53243 PAD.n10718 PAD.n10717 0.000734214
R53244 PAD.n7528 PAD.n7105 0.000729621
R53245 PAD.n2091 PAD.n2046 0.000729621
R53246 PAD.n8195 PAD.n8194 0.000725029
R53247 PAD.n9456 PAD.n9455 0.000725029
R53248 PAD.n11501 PAD.n11097 0.000725029
R53249 PAD.n7223 PAD.n7207 0.000720436
R53250 PAD.n8430 PAD.n4319 0.000715844
R53251 PAD.n8493 PAD.n3296 0.000706659
R53252 PAD.n8822 PAD.n2904 0.000706659
R53253 PAD.n8398 PAD.n8397 0.000697474
R53254 PAD.n8831 PAD.n2892 0.000697474
R53255 PAD.n9176 PAD.n2146 0.000692882
R53256 PAD.n9184 PAD.n2139 0.000692882
R53257 PAD.n8410 PAD.n8409 0.000688289
R53258 PAD.n8493 PAD.n8492 0.000688289
R53259 PAD.n9163 PAD.n2146 0.000688289
R53260 PAD.n9176 PAD.n9175 0.000688289
R53261 PAD.n8821 PAD.n8527 0.000683697
R53262 PAD.n8822 PAD.n8821 0.000679104
R53263 PAD.n2946 PAD.n2891 0.000679104
R53264 PAD.n1985 PAD.n1936 0.000679104
R53265 PAD.n11523 PAD.n10740 0.000679104
R53266 PAD.n4333 PAD.n4332 0.000674512
R53267 PAD.n8527 PAD 0.000674512
R53268 PAD.n10407 PAD.n435 0.000674512
R53269 PAD.n6396 PAD.n5904 0.00066992
R53270 PAD.n7521 PAD.n7158 0.00066992
R53271 PAD.n10008 PAD.n10007 0.00066992
R53272 PAD.n10702 PAD.n10701 0.00066992
R53273 PAD.n8194 PAD.n4843 0.000665327
R53274 PAD.n10362 PAD.n1130 0.000665327
R53275 PAD.n7802 PAD.n7801 0.000660735
R53276 PAD.n7060 PAD.n7059 0.000660735
R53277 PAD.n8183 PAD.n5183 0.000660735
R53278 PAD.n1131 PAD.n1118 0.000660735
R53279 PAD.n825 PAD.n776 0.000660735
R53280 PAD.n9151 PAD.n2487 0.000656142
R53281 PAD.n7783 PAD.n7782 0.00065155
R53282 PAD.n7820 PAD.n7819 0.00065155
R53283 PAD.n9742 PAD.n9741 0.00065155
R53284 PAD.n10728 PAD.n10727 0.00065155
R53285 PAD.n9445 PAD.n2089 0.000646958
R53286 PAD.n11507 PAD.n11098 0.000646958
R53287 PAD.n11302 PAD.n11096 0.000646958
R53288 PAD.n11509 PAD.n11099 0.000646958
R53289 PAD.n11510 PAD.n11100 0.000646958
R53290 PAD.n11513 PAD.n11105 0.000646958
R53291 PAD.n4842 PAD.n4841 0.000642365
R53292 PAD.n2089 PAD.n2037 0.000642365
R53293 PAD.n9732 PAD.n1594 0.00063318
R53294 PAD.n6699 PAD.n5894 0.000628588
R53295 PAD.n4321 PAD.n4028 0.000628588
R53296 PAD.n8410 PAD.n4331 0.000623995
R53297 PAD.n8419 PAD.n4333 0.000623995
R53298 PAD.n3339 PAD.n3287 0.000623995
R53299 PAD.n8519 PAD.n8518 0.000623995
R53300 PAD PAD.n2946 0.000614811
R53301 PAD.n6689 PAD.n5904 0.000610218
R53302 PAD.n6683 PAD.n6678 0.000610218
R53303 PAD.n3687 PAD.n3641 0.000610218
R53304 PAD.n8468 PAD.n3684 0.000610218
R53305 PAD.n8408 PAD.n8407 0.000605626
R53306 PAD.n8478 PAD.n3342 0.000605626
R53307 PAD.n9185 PAD.n9184 0.000605626
R53308 PAD.n10007 PAD.n1483 0.000605626
R53309 PAD.n10017 PAD.n1140 0.000605626
R53310 PAD.n8832 PAD.n2891 0.000601033
R53311 PAD.n1988 PAD.n1942 0.000601033
R53312 PAD.n7521 PAD.n7520 0.000596441
R53313 PAD.n7207 PAD.n7206 0.000596441
R53314 PAD.n8175 PAD.n5190 0.000596441
R53315 PAD.n9722 PAD.n9721 0.000596441
R53316 PAD.n10397 PAD.n433 0.000596441
R53317 PAD.n10753 PAD.n21 0.000596441
R53318 PAD.n10754 PAD.n10753 0.000596441
R53319 PAD.n6683 PAD.n6682 0.000587256
R53320 PAD.n7216 PAD.n7215 0.000587256
R53321 PAD.n8469 PAD.n8468 0.000587256
R53322 PAD.n10017 PAD.n10016 0.000587256
R53323 PAD.n434 PAD.n425 0.000587256
R53324 PAD.n7791 PAD.n6713 0.000582664
R53325 PAD.n8186 PAD.n4840 0.000582664
R53326 PAD.n1132 PAD.n1131 0.000582664
R53327 PAD.n6700 PAD.n6699 0.000578071
R53328 PAD.n7783 PAD.n7061 0.000578071
R53329 PAD.n10362 PAD.n10361 0.000578071
R53330 PAD.n10398 PAD.n10397 0.000578071
R53331 PAD.n10728 PAD.n32 0.000578071
R53332 PAD.n367 PAD.n20 0.000578071
R53333 PAD.n2894 PAD.n2879 0.000573479
R53334 PAD.n9143 PAD.n2494 0.000573479
R53335 PAD.n7829 PAD.n7828 0.000568886
R53336 PAD.n1593 PAD.n1586 0.000568886
R53337 PAD.n11534 PAD.n20 0.000568886
R53338 PAD.n8163 PAD.n5190 0.000564294
R53339 PAD.n10389 PAD.n10388 0.000564294
R53340 PAD.n8398 PAD.n4682 0.000559702
R53341 PAD.n9152 PAD.n2494 0.000559702
R53342 PAD.n9160 PAD.n2487 0.000559702
R53343 PAD.n9446 PAD.n2046 0.000559702
R53344 PAD.n9142 PAD.n9141 0.000550517
R53345 PAD.n9722 PAD.n1592 0.000550517
R53346 PAD.n7802 PAD.n5551 0.000545924
R53347 PAD.n8445 PAD.n8444 0.000545924
R53348 PAD.n8503 PAD.n8502 0.000541332
R53349 PAD.n3289 PAD.n2952 0.000541332
R53350 PAD.n9128 PAD.n2879 0.000541332
R53351 PAD.n9140 PAD.n2834 0.000541332
R53352 PAD.n10702 PAD.n419 0.000541332
R53353 PAD.n10716 PAD.n373 0.000541332
R53354 PAD.n6373 PAD.n5963 0.000536739
R53355 PAD.n5982 PAD.n5964 0.000536739
R53356 PAD.n5981 PAD.n5962 0.000536739
R53357 PAD.n5980 PAD.n5965 0.000536739
R53358 PAD.n5979 PAD.n5966 0.000536739
R53359 PAD.n8454 PAD.n3977 0.000532147
R53360 PAD.n9129 PAD.n2834 0.000532147
R53361 PAD.n7820 PAD.n5204 0.000522962
R53362 PAD.n7828 PAD.n5197 0.000522962
R53363 PAD.n8205 PAD.n4724 0.000522962
R53364 PAD.n9187 PAD.n9186 0.000522962
R53365 PAD.n8174 PAD.n5183 0.00051837
R53366 PAD.n9712 PAD.n1986 0.00051837
R53367 PAD.n1120 PAD.n828 0.00051837
R53368 PAD.n8165 PAD.n8164 0.000513777
R53369 PAD.n9733 PAD.n9732 0.000513777
R53370 PAD.n9741 PAD.n1536 0.000513777
R53371 PAD.n9999 PAD.n9998 0.000513777
R53372 PAD.n11533 PAD.n11532 0.000513777
R53373 PAD.n10755 PAD.n10740 0.000513777
R53374 PAD.n6680 PAD.n6679 0.000504592
R53375 PAD.n7528 PAD.n7103 0.000504592
R53376 PAD.n8431 PAD.n4028 0.000504592
R53377 PAD.n8444 PAD.n3983 0.000504592
R53378 PAD.n8453 PAD.n3687 0.000504592
R53379 PAD.n1142 PAD.n1141 0.000504592
R53380 PAD.n10408 PAD.n10407 0.000504592
R53381 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.pdrive_y_<0>.t4 115.13
R53382 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t0 GF_NI_BI_T_BASE_0.pdrive_y_<0>.n0 6.10848
R53383 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t1 GF_NI_BI_T_BASE_0.pdrive_y_<0>.n0 2.68197
R53384 GF_NI_BI_T_BASE_0.pdrive_y_<0>.n0 GF_NI_BI_T_BASE_0.pdrive_y_<0> 1.59856
R53385 GF_NI_BI_T_BASE_0.pdrive_y_<0>.n0 GF_NI_BI_T_BASE_0.pdrive_y_<0> 1.11644
R53386 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t3 GF_NI_BI_T_BASE_0.pdrive_y_<0> 0.773893
R53387 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.pdrive_y_<0>.t2 0.767197
R53388 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.pdrive_y_<0>.t1 0.7304
R53389 GF_NI_BI_T_BASE_0.pdrive_x_<1>.n1 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t4 113.415
R53390 GF_NI_BI_T_BASE_0.pdrive_x_<1>.n1 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t5 112.626
R53391 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t0 GF_NI_BI_T_BASE_0.pdrive_x_<1>.n0 6.12025
R53392 GF_NI_BI_T_BASE_0.pdrive_x_<1> GF_NI_BI_T_BASE_0.pdrive_x_<1>.n1 2.40503
R53393 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t3 GF_NI_BI_T_BASE_0.pdrive_x_<1>.n0 2.26404
R53394 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t2 GF_NI_BI_T_BASE_0.pdrive_x_<1> 1.43572
R53395 GF_NI_BI_T_BASE_0.pdrive_x_<1>.n0 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t2 1.0357
R53396 GF_NI_BI_T_BASE_0.pdrive_x_<1> GF_NI_BI_T_BASE_0.pdrive_x_<1>.t1 0.779435
R53397 GF_NI_BI_T_BASE_0.pdrive_x_<1> GF_NI_BI_T_BASE_0.pdrive_x_<1>.t3 0.7439
R53398 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.pdrive_y_<1>.t4 115.45
R53399 GF_NI_BI_T_BASE_0.pdrive_y_<1>.t0 GF_NI_BI_T_BASE_0.pdrive_y_<1>.n0 6.10848
R53400 GF_NI_BI_T_BASE_0.pdrive_y_<1>.t3 GF_NI_BI_T_BASE_0.pdrive_y_<1>.n0 2.68197
R53401 GF_NI_BI_T_BASE_0.pdrive_y_<1>.n0 GF_NI_BI_T_BASE_0.pdrive_y_<1> 1.59857
R53402 GF_NI_BI_T_BASE_0.pdrive_y_<1>.n0 GF_NI_BI_T_BASE_0.pdrive_y_<1> 1.11715
R53403 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.pdrive_y_<1>.t2 0.773875
R53404 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.pdrive_y_<1>.t1 0.766858
R53405 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.pdrive_y_<1>.t3 0.7304
R53406 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t2 4.05318
R53407 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n1 1.23426
R53408 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n0 1.23426
R53409 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D 1.10335
R53410 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t1 1.02238
R53411 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t0 1.0223
R53412 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n2 0.943559
R53413 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t6 0.618613
R53414 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t3 0.618613
R53415 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t4 0.618613
R53416 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t5 0.618613
R53417 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t6 6.51577
R53418 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t5 3.11732
R53419 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S 2.17664
R53420 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t4 1.85326
R53421 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t0 1.57786
R53422 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t2 1.56968
R53423 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t3 1.23492
R53424 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t1 1.02385
R53425 GF_NI_BI_T_BASE_0.ndrive_x_<1> GF_NI_BI_T_BASE_0.ndrive_x_<1>.t3 90.8824
R53426 GF_NI_BI_T_BASE_0.ndrive_x_<1>.t1 GF_NI_BI_T_BASE_0.ndrive_x_<1>.n0 7.28458
R53427 GF_NI_BI_T_BASE_0.ndrive_x_<1>.n0 GF_NI_BI_T_BASE_0.ndrive_x_<1>.t2 6.03391
R53428 GF_NI_BI_T_BASE_0.ndrive_x_<1>.n0 GF_NI_BI_T_BASE_0.ndrive_x_<1> 1.45646
R53429 GF_NI_BI_T_BASE_0.ndrive_x_<1> GF_NI_BI_T_BASE_0.ndrive_x_<1>.t1 0.951421
R53430 GF_NI_BI_T_BASE_0.ndrive_x_<1>.t0 GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.773893
R53431 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB.t3 82.1164
R53432 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB.t2 42.2319
R53433 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB.t1 2.04837
R53434 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB.t0 1.49421
R53435 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t5 80.4772
R53436 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t7 80.4772
R53437 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t4 62.5719
R53438 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t8 62.5719
R53439 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t6 45.4098
R53440 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t3 34.4148
R53441 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n1 8.06816
R53442 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n0 8.06816
R53443 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n2 6.31953
R53444 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n4 6.08116
R53445 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n3 4.80357
R53446 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t1 4.54043
R53447 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t0 1.1409
R53448 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 0.702557
R53449 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t4 45.4098
R53450 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t6 45.4098
R53451 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t9 45.4098
R53452 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t2 45.4098
R53453 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t3 34.4148
R53454 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t8 34.4148
R53455 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t7 34.4148
R53456 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t5 34.4148
R53457 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n6 9.02147
R53458 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n2 6.99208
R53459 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n5 6.273
R53460 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n3 6.273
R53461 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n1 6.273
R53462 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n0 6.273
R53463 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 5.57458
R53464 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n6 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 4.26721
R53465 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 4.26721
R53466 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 4.26721
R53467 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 2.39238
R53468 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t1 2.0632
R53469 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n6 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n4 1.30787
R53470 GF_NI_BI_T_BASE_0.pdrive_x_<0>.n2 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t5 113.251
R53471 GF_NI_BI_T_BASE_0.pdrive_x_<0>.n2 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t4 112.769
R53472 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t0 GF_NI_BI_T_BASE_0.pdrive_x_<0>.n1 6.12025
R53473 GF_NI_BI_T_BASE_0.pdrive_x_<0> GF_NI_BI_T_BASE_0.pdrive_x_<0>.n2 2.39
R53474 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t1 GF_NI_BI_T_BASE_0.pdrive_x_<0>.n1 2.26404
R53475 GF_NI_BI_T_BASE_0.pdrive_x_<0> GF_NI_BI_T_BASE_0.pdrive_x_<0>.n0 1.4357
R53476 GF_NI_BI_T_BASE_0.pdrive_x_<0>.n1 GF_NI_BI_T_BASE_0.pdrive_x_<0>.n0 1.03582
R53477 GF_NI_BI_T_BASE_0.pdrive_x_<0> GF_NI_BI_T_BASE_0.pdrive_x_<0>.t2 0.779294
R53478 GF_NI_BI_T_BASE_0.pdrive_x_<0> GF_NI_BI_T_BASE_0.pdrive_x_<0>.t1 0.7466
R53479 GF_NI_BI_T_BASE_0.pdrive_x_<0>.n0 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t3 0.66992
R53480 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t14 39.4055
R53481 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t13 35.4055
R53482 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t15 34.8841
R53483 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t11 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n0 4.05527
R53484 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t12 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n0 4.06684
R53485 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n12 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n8 6.3635
R53486 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n1 1.35467
R53487 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n14 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n13 5.38559
R53488 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n11 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n10 4.06578
R53489 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n3 4.0005
R53490 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n8 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t2 3.98107
R53491 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n11 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n9 3.16412
R53492 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n1 3.19389
R53493 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n8 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n7 2.94036
R53494 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n6 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n5 2.2505
R53495 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n12 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n11 2.2505
R53496 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n4 1.19063
R53497 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t4 3.19366
R53498 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n9 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t6 1.03341
R53499 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n14 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n2 1.03297
R53500 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n7 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t1 0.9105
R53501 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n7 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t0 0.9105
R53502 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n13 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n6 0.888086
R53503 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n10 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t10 0.847012
R53504 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n10 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t9 0.847012
R53505 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t6 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t5 0.5465
R53506 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t8 0.5465
R53507 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t7 0.5465
R53508 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n13 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n12 0.397741
R53509 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.291816
R53510 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n6 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.1355
R53511 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n14 0.122942
R53512 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n9 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.122187
R53513 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n5 1.38073
R53514 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t2 33.2287
R53515 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t1 25.193
R53516 PU.n3 PU.t2 40.5155
R53517 PU.n8 PU.n6 37.3205
R53518 PU.n0 PU.t3 35.5619
R53519 PU.n0 PU.t4 34.9362
R53520 PU.n3 PU.t5 26.3326
R53521 PU.n6 PU.n5 7.47146
R53522 PU.n1 PU.n0 4.00141
R53523 PU PU.n3 4.00106
R53524 PU.n2 PU.t1 3.17811
R53525 PU.n8 PU.n7 2.25122
R53526 PU PU.n8 1.98787
R53527 PU.n5 PU.t0 1.36552
R53528 PU.n7 PU.t6 1.31518
R53529 PU.n5 PU.n4 0.80237
R53530 PU.n4 PU.n2 0.45653
R53531 PU.n4 PU 0.163278
R53532 PU.n6 PU.n1 0.127056
R53533 PU.n2 PU 0.0456808
R53534 PU.n1 PU 0.00756793
R53535 PU.n7 PU 0.001225
R53536 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t3 82.1164
R53537 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t1 44.3219
R53538 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t2 42.2319
R53539 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t4 28.0534
R53540 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.n0 4.00859
R53541 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t0 1.33388
R53542 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D 6.03467
R53543 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t1 4.66477
R53544 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t3 3.2416
R53545 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t2 3.17822
R53546 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t3 37.5434
R53547 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t5 37.5434
R53548 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t2 25.3941
R53549 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t4 25.3941
R53550 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.n0 8.44221
R53551 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.n1 4.90922
R53552 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t0 2.6373
R53553 GF_NI_BI_T_BASE_0.pdrive_x_<2>.n3 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t4 113.415
R53554 GF_NI_BI_T_BASE_0.pdrive_x_<2>.n3 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t5 112.603
R53555 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t1 GF_NI_BI_T_BASE_0.pdrive_x_<2>.n2 6.12025
R53556 GF_NI_BI_T_BASE_0.pdrive_x_<2> GF_NI_BI_T_BASE_0.pdrive_x_<2>.n3 2.40448
R53557 GF_NI_BI_T_BASE_0.pdrive_x_<2>.n0 GF_NI_BI_T_BASE_0.pdrive_x_<2>.n2 2.26404
R53558 GF_NI_BI_T_BASE_0.pdrive_x_<2> GF_NI_BI_T_BASE_0.pdrive_x_<2>.n1 1.4357
R53559 GF_NI_BI_T_BASE_0.pdrive_x_<2>.n2 GF_NI_BI_T_BASE_0.pdrive_x_<2>.n1 1.03582
R53560 GF_NI_BI_T_BASE_0.pdrive_x_<2> GF_NI_BI_T_BASE_0.pdrive_x_<2>.t2 0.779294
R53561 GF_NI_BI_T_BASE_0.pdrive_x_<2> GF_NI_BI_T_BASE_0.pdrive_x_<2>.n0 0.7439
R53562 GF_NI_BI_T_BASE_0.pdrive_x_<2>.n1 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t3 0.66992
R53563 GF_NI_BI_T_BASE_0.pdrive_x_<2>.n0 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t0 0.360167
R53564 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t7 79.0838
R53565 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t4 78.041
R53566 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t6 34.4148
R53567 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t5 34.4148
R53568 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t2 34.4148
R53569 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t3 34.4148
R53570 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n2 10.9956
R53571 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n3 10.9956
R53572 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n4 10.9956
R53573 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n5 9.95826
R53574 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n1 8.49628
R53575 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t0 2.12938
R53576 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t1 1.97771
R53577 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n0 1.32326
R53578 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n6 1.25751
R53579 GF_NI_BI_T_BASE_0.ndrive_x_<3> GF_NI_BI_T_BASE_0.ndrive_x_<3>.t3 90.7152
R53580 GF_NI_BI_T_BASE_0.ndrive_x_<3>.t1 GF_NI_BI_T_BASE_0.ndrive_x_<3>.n0 7.28458
R53581 GF_NI_BI_T_BASE_0.ndrive_x_<3>.n0 GF_NI_BI_T_BASE_0.ndrive_x_<3>.t2 6.03391
R53582 GF_NI_BI_T_BASE_0.ndrive_x_<3>.n0 GF_NI_BI_T_BASE_0.ndrive_x_<3> 1.45646
R53583 GF_NI_BI_T_BASE_0.ndrive_x_<3> GF_NI_BI_T_BASE_0.ndrive_x_<3>.t1 0.951421
R53584 GF_NI_BI_T_BASE_0.ndrive_x_<3>.t0 GF_NI_BI_T_BASE_0.ndrive_x_<3> 0.773893
R53585 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t2 79.0838
R53586 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t6 78.041
R53587 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t3 34.4148
R53588 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t7 34.4148
R53589 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t4 34.4148
R53590 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t5 34.4148
R53591 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n2 10.9956
R53592 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n3 10.9956
R53593 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n4 10.9956
R53594 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n5 9.95826
R53595 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n1 8.49628
R53596 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t1 2.12938
R53597 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t0 1.97771
R53598 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n0 1.32326
R53599 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n6 1.25751
R53600 GF_NI_BI_T_BASE_0.ndrive_Y_<1> GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t5 90.7338
R53601 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n0 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t4 5.90425
R53602 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n2 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t2 2.41832
R53603 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n1 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t1 1.84043
R53604 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n0 GF_NI_BI_T_BASE_0.ndrive_Y_<1> 1.5749
R53605 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n3 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n2 1.48076
R53606 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n1 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n0 1.09118
R53607 GF_NI_BI_T_BASE_0.ndrive_Y_<1> GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n3 0.9455
R53608 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n2 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n1 0.578395
R53609 GF_NI_BI_T_BASE_0.ndrive_Y_<1> GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t3 0.500893
R53610 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n3 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t0 0.360167
R53611 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t7 40.4112
R53612 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t6 40.4112
R53613 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t13 40.4112
R53614 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t10 40.4112
R53615 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t2 40.4112
R53616 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t11 40.4112
R53617 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t4 35.3012
R53618 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t3 35.3012
R53619 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t9 35.3012
R53620 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t5 35.3012
R53621 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t12 35.3012
R53622 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t8 35.3012
R53623 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D 4.78544
R53624 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n0 4.13606
R53625 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n1 4.0005
R53626 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n5 4.0005
R53627 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n4 4.0005
R53628 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n3 4.0005
R53629 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n2 4.0005
R53630 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t0 3.91697
R53631 Y.n9 Y 9.72218
R53632 Y.n13 Y.n12 6.3005
R53633 Y Y.n13 3.18489
R53634 Y.n3 Y.n2 2.08611
R53635 Y.n1 Y.n0 2.08611
R53636 Y.n7 Y.n6 1.67295
R53637 Y.n7 Y.n5 1.09506
R53638 Y.n8 Y.n4 1.09506
R53639 Y.n2 Y.t7 1.0925
R53640 Y.n2 Y.t11 1.0925
R53641 Y.n0 Y.t8 1.0925
R53642 Y.n0 Y.t6 1.0925
R53643 Y.n13 Y.t10 1.0925
R53644 Y.n13 Y.t9 1.0925
R53645 Y.n12 Y.n11 0.825895
R53646 Y.n10 Y.n9 0.770237
R53647 Y.n8 Y.n7 0.578395
R53648 Y.n11 Y.n10 0.578395
R53649 Y.n6 Y.t5 0.5205
R53650 Y.n6 Y.t4 0.5205
R53651 Y.n5 Y.t3 0.5205
R53652 Y.n5 Y.t1 0.5205
R53653 Y.n4 Y.t2 0.5205
R53654 Y.n4 Y.t0 0.5205
R53655 Y.n9 Y.n8 0.457605
R53656 Y.n10 Y.n3 0.336924
R53657 Y.n11 Y.n1 0.336924
R53658 Y Y.n12 0.1355
R53659 Y.n3 Y 0.0456808
R53660 Y.n1 Y 0.0456808
R53661 PDRV0.n21 PDRV0.n20 227.274
R53662 PDRV0.n30 PDRV0.n29 227.274
R53663 PDRV0.n21 PDRV0.t0 113.636
R53664 PDRV0.n30 PDRV0.t0 113.636
R53665 PDRV0.n1 PDRV0.t2 46.7726
R53666 PDRV0.n1 PDRV0.t1 41.2455
R53667 PDRV0.n3 PDRV0 21.925
R53668 PDRV0.n22 PDRV0.n11 10.5005
R53669 PDRV0.n22 PDRV0.n7 10.5005
R53670 PDRV0.n8 PDRV0.n7 10.5005
R53671 PDRV0.n18 PDRV0.n13 10.5005
R53672 PDRV0.n14 PDRV0.n5 10.5005
R53673 PDRV0.n31 PDRV0.n5 10.5005
R53674 PDRV0.n31 PDRV0.n6 10.5005
R53675 PDRV0.n27 PDRV0.n8 7.3505
R53676 PDRV0.n16 PDRV0.n13 6.3005
R53677 PDRV0.n18 PDRV0.n17 6.3005
R53678 PDRV0.n27 PDRV0.n26 6.3005
R53679 PDRV0.n25 PDRV0.n8 6.3005
R53680 PDRV0.n29 PDRV0.n8 6.3005
R53681 PDRV0.n24 PDRV0.n7 6.3005
R53682 PDRV0.n30 PDRV0.n7 6.3005
R53683 PDRV0.n23 PDRV0.n22 6.3005
R53684 PDRV0.n22 PDRV0.n21 6.3005
R53685 PDRV0.n11 PDRV0.n10 6.3005
R53686 PDRV0.n32 PDRV0.n31 6.3005
R53687 PDRV0.n31 PDRV0.n30 6.3005
R53688 PDRV0.n5 PDRV0.n0 6.3005
R53689 PDRV0.n21 PDRV0.n5 6.3005
R53690 PDRV0.n15 PDRV0.n14 6.3005
R53691 PDRV0.n29 PDRV0.n6 6.3005
R53692 PDRV0.n28 PDRV0.n9 5.18619
R53693 PDRV0.n4 PDRV0.n3 4.53118
R53694 PDRV0.n2 PDRV0.n1 4.0005
R53695 PDRV0.n28 PDRV0.n27 2.86464
R53696 PDRV0.n9 PDRV0.n6 2.32205
R53697 PDRV0.n13 PDRV0.n12 2.32205
R53698 PDRV0.n19 PDRV0.n18 2.32205
R53699 PDRV0.n19 PDRV0.n11 2.32205
R53700 PDRV0.n14 PDRV0.n12 2.32205
R53701 PDRV0.n3 PDRV0.n2 2.2505
R53702 PDRV0.n20 PDRV0.n12 1.99047
R53703 PDRV0.n20 PDRV0.n19 1.99047
R53704 PDRV0.n9 PDRV0.n4 1.99047
R53705 PDRV0.n29 PDRV0.n28 1.71918
R53706 PDRV0.n23 PDRV0.n10 0.1505
R53707 PDRV0.n25 PDRV0.n24 0.1505
R53708 PDRV0.n15 PDRV0.n0 0.1505
R53709 PDRV0.n32 PDRV0.n4 0.1235
R53710 PDRV0.n26 PDRV0.n25 0.1055
R53711 PDRV0.n16 PDRV0.n15 0.1055
R53712 PDRV0.n17 PDRV0.n10 0.1055
R53713 PDRV0.n26 PDRV0 0.0755
R53714 PDRV0 PDRV0.n23 0.0755
R53715 PDRV0.n24 PDRV0 0.0755
R53716 PDRV0 PDRV0.n16 0.0755
R53717 PDRV0.n17 PDRV0 0.0755
R53718 PDRV0 PDRV0.n0 0.0755
R53719 PDRV0 PDRV0.n32 0.0755
R53720 PDRV0 PDRV0.n4 0.0455
R53721 PDRV0.n2 PDRV0 0.002
R53722 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t3 38.8469
R53723 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t2 22.5262
R53724 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.n0 12.9666
R53725 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t1 2.79762
R53726 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t7 79.0838
R53727 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t5 78.041
R53728 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t2 34.4148
R53729 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t6 34.4148
R53730 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t3 34.4148
R53731 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t4 34.4148
R53732 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n4 10.9956
R53733 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n3 10.9956
R53734 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n2 10.9956
R53735 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n5 9.95826
R53736 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n1 8.49628
R53737 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t1 2.12938
R53738 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t0 1.97771
R53739 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n0 1.32326
R53740 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n6 1.25751
R53741 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.pdrive_y_<3>.t4 115.088
R53742 GF_NI_BI_T_BASE_0.pdrive_y_<3>.t0 GF_NI_BI_T_BASE_0.pdrive_y_<3>.n1 6.10848
R53743 GF_NI_BI_T_BASE_0.pdrive_y_<3>.n0 GF_NI_BI_T_BASE_0.pdrive_y_<3>.n1 2.68197
R53744 GF_NI_BI_T_BASE_0.pdrive_y_<3>.n2 GF_NI_BI_T_BASE_0.pdrive_y_<3> 1.59857
R53745 GF_NI_BI_T_BASE_0.pdrive_y_<3>.n2 GF_NI_BI_T_BASE_0.pdrive_y_<3> 0.781133
R53746 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.pdrive_y_<3>.n0 0.7304
R53747 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.pdrive_y_<3>.t2 0.500875
R53748 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.pdrive_y_<3>.t3 0.493858
R53749 GF_NI_BI_T_BASE_0.pdrive_y_<3>.n0 GF_NI_BI_T_BASE_0.pdrive_y_<3>.t1 0.360167
R53750 GF_NI_BI_T_BASE_0.pdrive_y_<3>.n1 GF_NI_BI_T_BASE_0.pdrive_y_<3>.n2 0.336519
R53751 a_5575_63014.t0 a_5575_63014.n2 4.28715
R53752 a_5575_63014.n3 a_5575_63014.t5 5.32188
R53753 a_5575_63014.t1 a_5575_63014.n0 4.29256
R53754 a_5575_63014.n3 a_5575_63014.n1 2.84024
R53755 a_5575_63014.t4 a_5575_63014.n0 1.30198
R53756 a_5575_63014.n1 a_5575_63014.n2 0.00322045
R53757 a_5575_63014.n1 a_5575_63014.t3 2.34839
R53758 a_5575_63014.n0 a_5575_63014.n3 2.28727
R53759 a_5575_63014.n2 a_5575_63014.t2 8.1298
R53760 GF_NI_BI_T_BASE_0.ndrive_Y_<3> GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t5 89.3064
R53761 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n1 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t4 5.90425
R53762 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n3 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t0 2.41832
R53763 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n2 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t3 1.84043
R53764 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n1 GF_NI_BI_T_BASE_0.ndrive_Y_<3> 1.5749
R53765 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n0 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n3 1.48076
R53766 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n2 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n1 1.09118
R53767 GF_NI_BI_T_BASE_0.ndrive_Y_<3> GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n0 0.9455
R53768 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n3 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n2 0.578395
R53769 GF_NI_BI_T_BASE_0.ndrive_Y_<3> GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t2 0.500893
R53770 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n0 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t1 0.360167
R53771 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t0 35.9269
R53772 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t1 30.9212
R53773 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A 25.1335
R53774 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.n0 4.0005
R53775 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t2 37.5434
R53776 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t4 37.5434
R53777 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t5 25.3941
R53778 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t3 25.3941
R53779 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.n0 8.44221
R53780 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.n1 4.90922
R53781 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t1 2.6373
R53782 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS.t1 22.3936
R53783 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t2 82.1164
R53784 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t3 82.1164
R53785 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.n1 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t6 44.3219
R53786 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t5 42.2319
R53787 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t7 42.2319
R53788 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.n1 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t4 28.0534
R53789 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN 11.0504
R53790 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.n0 7.90454
R53791 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN 7.30826
R53792 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.n1 4.09808
R53793 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t0 1.53534
R53794 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t1 1.33388
R53795 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t4 37.5434
R53796 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t2 37.5434
R53797 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t3 25.3941
R53798 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t5 25.3941
R53799 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.n0 8.44221
R53800 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.n1 4.90922
R53801 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t1 2.6373
R53802 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t4 37.5434
R53803 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t2 37.5434
R53804 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t3 25.3941
R53805 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t5 25.3941
R53806 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.n0 8.44221
R53807 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314531_1.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.n1 4.40816
R53808 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314531_1.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t0 2.2762
R53809 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314531_1.D 2.08654
R53810 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t2 24.9619
R53811 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t0 2.39238
R53812 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t1 2.0632
R53813 GF_NI_BI_T_BASE_0.ndrive_y_<2> GF_NI_BI_T_BASE_0.ndrive_y_<2>.t5 90.9292
R53814 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n1 GF_NI_BI_T_BASE_0.ndrive_y_<2> 12.0008
R53815 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n0 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t4 5.90425
R53816 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n3 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t2 2.41832
R53817 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n0 GF_NI_BI_T_BASE_0.ndrive_y_<2> 1.5749
R53818 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n4 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n3 1.48076
R53819 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n2 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n1 1.48076
R53820 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n2 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n0 1.09118
R53821 GF_NI_BI_T_BASE_0.ndrive_y_<2> GF_NI_BI_T_BASE_0.ndrive_y_<2>.n4 0.9455
R53822 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n3 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n2 0.578395
R53823 GF_NI_BI_T_BASE_0.ndrive_y_<2> GF_NI_BI_T_BASE_0.ndrive_y_<2>.t3 0.500893
R53824 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n4 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t0 0.360167
R53825 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n1 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t1 0.360167
R53826 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314531_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB.t0 2.36868
R53827 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314531_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB.t1 2.08654
R53828 GF_NI_BI_T_BASE_0.pdrive_x_<3>.n3 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t5 113.317
R53829 GF_NI_BI_T_BASE_0.pdrive_x_<3>.n3 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t4 112.746
R53830 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t0 GF_NI_BI_T_BASE_0.pdrive_x_<3>.n1 6.12025
R53831 GF_NI_BI_T_BASE_0.pdrive_x_<3> GF_NI_BI_T_BASE_0.pdrive_x_<3>.n3 2.39
R53832 GF_NI_BI_T_BASE_0.pdrive_x_<3>.n0 GF_NI_BI_T_BASE_0.pdrive_x_<3>.n1 2.26404
R53833 GF_NI_BI_T_BASE_0.pdrive_x_<3>.n2 GF_NI_BI_T_BASE_0.pdrive_x_<3> 1.43572
R53834 GF_NI_BI_T_BASE_0.pdrive_x_<3>.n1 GF_NI_BI_T_BASE_0.pdrive_x_<3>.n2 1.0357
R53835 GF_NI_BI_T_BASE_0.pdrive_x_<3> GF_NI_BI_T_BASE_0.pdrive_x_<3>.t3 0.779435
R53836 GF_NI_BI_T_BASE_0.pdrive_x_<3> GF_NI_BI_T_BASE_0.pdrive_x_<3>.n0 0.7466
R53837 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t2 GF_NI_BI_T_BASE_0.pdrive_x_<3>.n2 0.396936
R53838 GF_NI_BI_T_BASE_0.pdrive_x_<3>.n0 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t1 0.360167
R53839 IE.n0 IE.t2 35.9269
R53840 IE.n0 IE.t0 30.9212
R53841 IE IE.n0 4.0005
R53842 IE.n2 IE 3.56853
R53843 IE.n2 IE.n1 2.25122
R53844 IE.n1 IE.t1 1.31518
R53845 IE IE.n2 0.63879
R53846 IE.n1 IE 0.001225
R53847 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t4 37.5434
R53848 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t5 37.5434
R53849 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t2 25.3941
R53850 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t3 25.3941
R53851 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.n0 8.44221
R53852 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.n1 4.90922
R53853 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t1 2.6373
R53854 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t3 37.5434
R53855 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t4 37.5434
R53856 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t2 26.1617
R53857 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t5 25.3941
R53858 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t6 25.3941
R53859 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n0 8.44221
R53860 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n1 4.40816
R53861 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t0 2.2999
R53862 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t1 2.0632
R53863 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t8 80.4772
R53864 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t4 80.4772
R53865 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t7 62.5719
R53866 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t5 62.5719
R53867 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t3 45.4098
R53868 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t6 34.4148
R53869 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n1 8.06816
R53870 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n0 8.06816
R53871 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n2 6.31953
R53872 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n4 6.08116
R53873 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n3 4.80357
R53874 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t1 4.54043
R53875 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t2 1.1409
R53876 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 0.702557
R53877 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t6 80.4772
R53878 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t3 80.4772
R53879 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t8 62.5719
R53880 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t7 62.5719
R53881 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t4 45.4098
R53882 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t5 34.4148
R53883 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n1 8.06816
R53884 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n0 8.06816
R53885 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n2 6.31953
R53886 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n4 6.08116
R53887 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n3 4.80357
R53888 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t2 4.54043
R53889 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t1 1.1409
R53890 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 0.702585
R53891 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n1 3.11956
R53892 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n0 2.91689
R53893 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n0 0.0638785
R53894 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n2 0.055602
R53895 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n1 6.35009
R53896 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n2 11.9543
R53897 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 11.0117
R53898 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t0 1.0925
R53899 GF_NI_BI_T_BASE_0.pdrive_y_<2> GF_NI_BI_T_BASE_0.pdrive_y_<2>.t4 115.388
R53900 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t2 GF_NI_BI_T_BASE_0.pdrive_y_<2>.n1 6.10848
R53901 GF_NI_BI_T_BASE_0.pdrive_y_<2>.n0 GF_NI_BI_T_BASE_0.pdrive_y_<2>.n1 2.68197
R53902 GF_NI_BI_T_BASE_0.pdrive_y_<2>.n2 GF_NI_BI_T_BASE_0.pdrive_y_<2> 1.59856
R53903 GF_NI_BI_T_BASE_0.pdrive_y_<2>.n2 GF_NI_BI_T_BASE_0.pdrive_y_<2> 0.780424
R53904 GF_NI_BI_T_BASE_0.pdrive_y_<2> GF_NI_BI_T_BASE_0.pdrive_y_<2>.n0 0.7304
R53905 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t1 GF_NI_BI_T_BASE_0.pdrive_y_<2> 0.500893
R53906 GF_NI_BI_T_BASE_0.pdrive_y_<2> GF_NI_BI_T_BASE_0.pdrive_y_<2>.t3 0.494197
R53907 GF_NI_BI_T_BASE_0.pdrive_y_<2>.n0 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t0 0.360167
R53908 GF_NI_BI_T_BASE_0.pdrive_y_<2>.n1 GF_NI_BI_T_BASE_0.pdrive_y_<2>.n2 0.336519
R53909 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t3 22.8162
R53910 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t4 22.3026
R53911 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t2 20.1892
R53912 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n1 11.9677
R53913 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t1 1.55917
R53914 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t0 1.45173
R53915 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n0 1.38831
R53916 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t2 19.4535
R53917 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t1 13.1326
R53918 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t0 8.30501
R53919 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t0 8.14999
R53920 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.n0 5.61641
R53921 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t3 44.3219
R53922 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t2 28.0534
R53923 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.n0 4.18151
R53924 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t1 1.76195
R53925 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t0 1.56963
R53926 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314531_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB.t0 2.36868
R53927 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314531_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB.t1 2.08654
R53928 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS 11.0117
R53929 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS.t1 11.0117
R53930 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.MINUS.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.MINUS.t1 22.3936
R53931 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t5 82.1164
R53932 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t4 44.3219
R53933 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t2 42.2319
R53934 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t3 28.0534
R53935 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.n0 4.09808
R53936 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t1 1.53534
R53937 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t0 1.33388
R53938 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t5 79.0838
R53939 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t3 78.041
R53940 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t6 34.4148
R53941 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t4 34.4148
R53942 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t7 34.4148
R53943 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t2 34.4148
R53944 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n4 10.9956
R53945 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n3 10.9956
R53946 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n2 10.9956
R53947 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n5 9.95826
R53948 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n1 8.49628
R53949 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t1 2.12938
R53950 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t0 1.97771
R53951 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n0 1.32326
R53952 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n6 1.25751
R53953 OE.n22 OE.n8 227.274
R53954 OE.n23 OE.n4 227.274
R53955 OE.n44 OE.n39 227.274
R53956 OE.n55 OE.n45 227.274
R53957 OE.n92 OE.n78 227.274
R53958 OE.n93 OE.n74 227.274
R53959 OE.t2 OE.n22 113.636
R53960 OE.n23 OE.t2 113.636
R53961 OE.t1 OE.n44 113.636
R53962 OE.n55 OE.t1 113.636
R53963 OE.t0 OE.n92 113.636
R53964 OE.n93 OE.t0 113.636
R53965 OE.n33 OE.t6 46.7726
R53966 OE.n67 OE.t9 46.7726
R53967 OE.n103 OE.t3 46.7726
R53968 OE.n0 OE.t10 46.7726
R53969 OE.n33 OE.t8 41.2455
R53970 OE.n67 OE.t4 41.2455
R53971 OE.n103 OE.t7 41.2455
R53972 OE.n0 OE.t5 41.2455
R53973 OE.n107 OE 25.7369
R53974 OE.n17 OE.n16 10.5005
R53975 OE.n21 OE.n9 10.5005
R53976 OE.n21 OE.n3 10.5005
R53977 OE.n31 OE.n3 10.5005
R53978 OE.n29 OE.n28 10.5005
R53979 OE.n13 OE.n7 10.5005
R53980 OE.n24 OE.n7 10.5005
R53981 OE.n25 OE.n24 10.5005
R53982 OE.n63 OE.n62 10.5005
R53983 OE.n60 OE.n41 10.5005
R53984 OE.n56 OE.n41 10.5005
R53985 OE.n56 OE.n43 10.5005
R53986 OE.n65 OE.n38 10.5005
R53987 OE.n54 OE.n38 10.5005
R53988 OE.n54 OE.n46 10.5005
R53989 OE.n87 OE.n86 10.5005
R53990 OE.n91 OE.n79 10.5005
R53991 OE.n91 OE.n73 10.5005
R53992 OE.n101 OE.n73 10.5005
R53993 OE.n99 OE.n98 10.5005
R53994 OE.n83 OE.n77 10.5005
R53995 OE.n94 OE.n77 10.5005
R53996 OE.n95 OE.n94 10.5005
R53997 OE.n70 OE.n35 7.68484
R53998 OE.n50 OE.n46 7.3505
R53999 OE.n48 OE.n43 7.3505
R54000 OE.n108 OE.n107 6.57761
R54001 OE.n18 OE.n17 6.3005
R54002 OE.n16 OE.n15 6.3005
R54003 OE.n3 OE.n1 6.3005
R54004 OE.n23 OE.n3 6.3005
R54005 OE.n21 OE.n20 6.3005
R54006 OE.n22 OE.n21 6.3005
R54007 OE.n19 OE.n9 6.3005
R54008 OE.n26 OE.n25 6.3005
R54009 OE.n24 OE.n6 6.3005
R54010 OE.n24 OE.n23 6.3005
R54011 OE.n12 OE.n7 6.3005
R54012 OE.n22 OE.n7 6.3005
R54013 OE.n14 OE.n13 6.3005
R54014 OE.n28 OE.n27 6.3005
R54015 OE.n29 OE.n2 6.3005
R54016 OE.n32 OE.n31 6.3005
R54017 OE.n52 OE.n46 6.3005
R54018 OE.n46 OE.n45 6.3005
R54019 OE.n54 OE.n53 6.3005
R54020 OE.n55 OE.n54 6.3005
R54021 OE.n38 OE.n36 6.3005
R54022 OE.n44 OE.n38 6.3005
R54023 OE.n48 OE.n47 6.3005
R54024 OE.n51 OE.n50 6.3005
R54025 OE.n43 OE.n42 6.3005
R54026 OE.n45 OE.n43 6.3005
R54027 OE.n57 OE.n56 6.3005
R54028 OE.n56 OE.n55 6.3005
R54029 OE.n58 OE.n41 6.3005
R54030 OE.n44 OE.n41 6.3005
R54031 OE.n60 OE.n59 6.3005
R54032 OE.n63 OE.n37 6.3005
R54033 OE.n62 OE.n40 6.3005
R54034 OE.n66 OE.n65 6.3005
R54035 OE.n88 OE.n87 6.3005
R54036 OE.n86 OE.n85 6.3005
R54037 OE.n73 OE.n71 6.3005
R54038 OE.n93 OE.n73 6.3005
R54039 OE.n91 OE.n90 6.3005
R54040 OE.n92 OE.n91 6.3005
R54041 OE.n89 OE.n79 6.3005
R54042 OE.n96 OE.n95 6.3005
R54043 OE.n94 OE.n76 6.3005
R54044 OE.n94 OE.n93 6.3005
R54045 OE.n82 OE.n77 6.3005
R54046 OE.n92 OE.n77 6.3005
R54047 OE.n84 OE.n83 6.3005
R54048 OE.n98 OE.n97 6.3005
R54049 OE.n99 OE.n72 6.3005
R54050 OE.n102 OE.n101 6.3005
R54051 OE.n35 OE.n32 4.67458
R54052 OE.n69 OE.n66 4.67458
R54053 OE.n105 OE.n102 4.67458
R54054 OE.n107 OE.n106 4.54195
R54055 OE.n70 OE.n69 4.22221
R54056 OE.n106 OE.n105 4.22221
R54057 OE.n34 OE.n33 4.0005
R54058 OE.n68 OE.n67 4.0005
R54059 OE.n104 OE.n103 4.0005
R54060 OE.n108 OE.n0 4.0005
R54061 OE.n50 OE.n49 2.86464
R54062 OE.n49 OE.n48 2.86464
R54063 OE.n106 OE.n70 2.62471
R54064 OE.n35 OE.n34 2.49418
R54065 OE.n69 OE.n68 2.49418
R54066 OE.n105 OE.n104 2.49418
R54067 OE.n17 OE.n10 2.32205
R54068 OE.n16 OE.n11 2.32205
R54069 OE.n10 OE.n9 2.32205
R54070 OE.n30 OE.n29 2.32205
R54071 OE.n28 OE.n5 2.32205
R54072 OE.n25 OE.n5 2.32205
R54073 OE.n13 OE.n11 2.32205
R54074 OE.n31 OE.n30 2.32205
R54075 OE.n64 OE.n63 2.32205
R54076 OE.n61 OE.n60 2.32205
R54077 OE.n62 OE.n61 2.32205
R54078 OE.n65 OE.n64 2.32205
R54079 OE.n87 OE.n80 2.32205
R54080 OE.n86 OE.n81 2.32205
R54081 OE.n80 OE.n79 2.32205
R54082 OE.n100 OE.n99 2.32205
R54083 OE.n98 OE.n75 2.32205
R54084 OE.n95 OE.n75 2.32205
R54085 OE.n83 OE.n81 2.32205
R54086 OE.n101 OE.n100 2.32205
R54087 OE.n10 OE.n8 1.99047
R54088 OE.n11 OE.n8 1.99047
R54089 OE.n5 OE.n4 1.99047
R54090 OE.n30 OE.n4 1.99047
R54091 OE.n61 OE.n39 1.99047
R54092 OE.n64 OE.n39 1.99047
R54093 OE.n80 OE.n78 1.99047
R54094 OE.n81 OE.n78 1.99047
R54095 OE.n75 OE.n74 1.99047
R54096 OE.n100 OE.n74 1.99047
R54097 OE.n49 OE.n45 1.71918
R54098 OE.n20 OE.n19 0.1505
R54099 OE.n14 OE.n12 0.1505
R54100 OE.n26 OE.n6 0.1505
R54101 OE.n53 OE.n52 0.1505
R54102 OE.n59 OE.n58 0.1505
R54103 OE.n57 OE.n42 0.1505
R54104 OE.n90 OE.n89 0.1505
R54105 OE.n84 OE.n82 0.1505
R54106 OE.n96 OE.n76 0.1505
R54107 OE.n32 OE.n2 0.148132
R54108 OE.n66 OE.n37 0.148132
R54109 OE.n102 OE.n72 0.148132
R54110 OE.n19 OE.n18 0.1055
R54111 OE.n15 OE.n14 0.1055
R54112 OE.n27 OE.n26 0.1055
R54113 OE.n52 OE.n51 0.1055
R54114 OE.n47 OE.n42 0.1055
R54115 OE.n59 OE.n40 0.1055
R54116 OE.n89 OE.n88 0.1055
R54117 OE.n85 OE.n84 0.1055
R54118 OE.n97 OE.n96 0.1055
R54119 OE.n32 OE.n1 0.1005
R54120 OE.n66 OE.n36 0.1005
R54121 OE.n102 OE.n71 0.1005
R54122 OE.n18 OE 0.0755
R54123 OE.n15 OE 0.0755
R54124 OE.n20 OE 0.0755
R54125 OE OE.n1 0.0755
R54126 OE.n12 OE 0.0755
R54127 OE OE.n6 0.0755
R54128 OE OE.n2 0.0755
R54129 OE.n27 OE 0.0755
R54130 OE OE.n36 0.0755
R54131 OE.n53 OE 0.0755
R54132 OE.n51 OE 0.0755
R54133 OE.n47 OE 0.0755
R54134 OE.n58 OE 0.0755
R54135 OE OE.n57 0.0755
R54136 OE OE.n37 0.0755
R54137 OE.n40 OE 0.0755
R54138 OE.n88 OE 0.0755
R54139 OE.n85 OE 0.0755
R54140 OE.n90 OE 0.0755
R54141 OE OE.n71 0.0755
R54142 OE.n82 OE 0.0755
R54143 OE OE.n76 0.0755
R54144 OE OE.n72 0.0755
R54145 OE.n97 OE 0.0755
R54146 OE OE.n108 0.004
R54147 OE.n34 OE 0.00168421
R54148 OE.n68 OE 0.00168421
R54149 OE.n104 OE 0.00168421
R54150 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.D GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S.n0 1.15854
R54151 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S.t1 0.5465
R54152 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S.t0 0.5465
R54153 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t3 38.8469
R54154 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t2 22.5262
R54155 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.n0 12.9666
R54156 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t1 2.79762
R54157 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.ndrive_x_<2>.t3 90.7537
R54158 GF_NI_BI_T_BASE_0.ndrive_x_<2>.n0 GF_NI_BI_T_BASE_0.ndrive_x_<2>.n1 7.28458
R54159 GF_NI_BI_T_BASE_0.ndrive_x_<2>.n1 GF_NI_BI_T_BASE_0.ndrive_x_<2>.t2 6.03391
R54160 GF_NI_BI_T_BASE_0.ndrive_x_<2>.n1 GF_NI_BI_T_BASE_0.ndrive_x_<2> 1.45646
R54161 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.ndrive_x_<2>.n0 0.951421
R54162 GF_NI_BI_T_BASE_0.ndrive_x_<2>.t1 GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.500893
R54163 GF_NI_BI_T_BASE_0.ndrive_x_<2>.n0 GF_NI_BI_T_BASE_0.ndrive_x_<2>.t0 0.360167
R54164 PDRV1.n19 PDRV1.n18 227.274
R54165 PDRV1.n30 PDRV1.n29 227.274
R54166 PDRV1.n19 PDRV1.t0 113.636
R54167 PDRV1.n30 PDRV1.t0 113.636
R54168 PDRV1.n12 PDRV1.t2 46.7726
R54169 PDRV1.n12 PDRV1.t1 41.2455
R54170 PDRV1.n14 PDRV1 30.9297
R54171 PDRV1.n17 PDRV1.n2 10.5005
R54172 PDRV1.n31 PDRV1.n2 10.5005
R54173 PDRV1.n31 PDRV1.n3 10.5005
R54174 PDRV1.n23 PDRV1.n6 10.5005
R54175 PDRV1.n20 PDRV1.n8 10.5005
R54176 PDRV1.n20 PDRV1.n4 10.5005
R54177 PDRV1.n27 PDRV1.n4 10.5005
R54178 PDRV1.n10 PDRV1.n8 7.3505
R54179 PDRV1.n11 PDRV1.n10 6.3005
R54180 PDRV1.n27 PDRV1.n26 6.3005
R54181 PDRV1.n22 PDRV1.n4 6.3005
R54182 PDRV1.n30 PDRV1.n4 6.3005
R54183 PDRV1.n21 PDRV1.n20 6.3005
R54184 PDRV1.n20 PDRV1.n19 6.3005
R54185 PDRV1.n8 PDRV1.n7 6.3005
R54186 PDRV1.n18 PDRV1.n8 6.3005
R54187 PDRV1.n25 PDRV1.n6 6.3005
R54188 PDRV1.n24 PDRV1.n23 6.3005
R54189 PDRV1.n3 PDRV1.n1 6.3005
R54190 PDRV1.n32 PDRV1.n31 6.3005
R54191 PDRV1.n31 PDRV1.n30 6.3005
R54192 PDRV1.n2 PDRV1.n0 6.3005
R54193 PDRV1.n19 PDRV1.n2 6.3005
R54194 PDRV1.n18 PDRV1.n17 6.3005
R54195 PDRV1.n16 PDRV1.n9 5.18619
R54196 PDRV1.n15 PDRV1.n14 4.53118
R54197 PDRV1.n13 PDRV1.n12 4.0005
R54198 PDRV1.n10 PDRV1.n9 2.86464
R54199 PDRV1.n17 PDRV1.n16 2.32205
R54200 PDRV1.n5 PDRV1.n3 2.32205
R54201 PDRV1.n28 PDRV1.n6 2.32205
R54202 PDRV1.n28 PDRV1.n27 2.32205
R54203 PDRV1.n23 PDRV1.n5 2.32205
R54204 PDRV1.n14 PDRV1.n13 2.2505
R54205 PDRV1.n29 PDRV1.n28 1.99047
R54206 PDRV1.n29 PDRV1.n5 1.99047
R54207 PDRV1.n16 PDRV1.n15 1.99047
R54208 PDRV1.n18 PDRV1.n9 1.71918
R54209 PDRV1.n21 PDRV1.n7 0.1505
R54210 PDRV1.n26 PDRV1.n22 0.1505
R54211 PDRV1.n32 PDRV1.n1 0.1505
R54212 PDRV1.n15 PDRV1.n0 0.1235
R54213 PDRV1.n11 PDRV1.n7 0.1055
R54214 PDRV1.n24 PDRV1.n1 0.1055
R54215 PDRV1.n26 PDRV1.n25 0.1055
R54216 PDRV1 PDRV1.n11 0.0755
R54217 PDRV1 PDRV1.n21 0.0755
R54218 PDRV1.n22 PDRV1 0.0755
R54219 PDRV1 PDRV1.n24 0.0755
R54220 PDRV1.n25 PDRV1 0.0755
R54221 PDRV1 PDRV1.n0 0.0755
R54222 PDRV1 PDRV1.n32 0.0755
R54223 PDRV1.n15 PDRV1 0.0455
R54224 PDRV1.n13 PDRV1 0.002
R54225 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t3 38.8469
R54226 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t2 22.5262
R54227 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t1 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.n0 12.9666
R54228 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t1 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t0 2.79762
R54229 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t4 82.1164
R54230 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t5 82.1164
R54231 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t3 42.2319
R54232 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t2 42.2319
R54233 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB 10.4346
R54234 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB 9.25386
R54235 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.n0 7.14721
R54236 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t0 2.04837
R54237 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t1 1.49421
R54238 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t3 38.8469
R54239 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t2 22.5262
R54240 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t1 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.n0 12.9564
R54241 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t1 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t0 2.79762
R54242 A.n0 A.t2 46.7726
R54243 A.n0 A.t0 41.2455
R54244 A.n2 A 24.6463
R54245 A.n3 A.n2 7.84234
R54246 A.n2 A.n1 5.59634
R54247 A.n3 A.n0 4.0005
R54248 A A.t1 2.6293
R54249 A.n1 A.t1 2.60635
R54250 A.n1 A 0.02345
R54251 A A.n3 0.0025
R54252 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t8 41.7148
R54253 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t7 41.7148
R54254 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t4 34.2225
R54255 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t3 34.0869
R54256 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t6 30.0869
R54257 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t5 30.0869
R54258 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t0 4.67357
R54259 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n2 4.0005
R54260 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n3 4.0005
R54261 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S 2.87207
R54262 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t2 1.81789
R54263 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t1 1.22475
R54264 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n0 1.14881
R54265 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.D GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S.n0 1.15854
R54266 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S.t1 0.5465
R54267 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S.t0 0.5465
R54268 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t2 82.1164
R54269 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t3 42.2319
R54270 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t0 2.04837
R54271 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t1 1.49421
R54272 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_2.PLUS.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_2.PLUS.t1 22.3936
R54273 PD.n5 PD.t3 35.5619
R54274 PD PD.t2 35.4693
R54275 PD.n5 PD.t4 34.9362
R54276 PD.n2 PD.t1 33.3819
R54277 PD.n3 PD.t0 28.9398
R54278 PD PD.n7 23.3129
R54279 PD.n2 PD.t5 16.3212
R54280 PD.n3 PD.n2 12.3062
R54281 PD.n1 PD 4.84629
R54282 PD.n7 PD.n4 4.73379
R54283 PD.n7 PD.n6 4.00668
R54284 PD PD.n3 4.00168
R54285 PD.n6 PD.n5 4.0005
R54286 PD.n4 PD 2.3055
R54287 PD.n1 PD.n0 2.25122
R54288 PD.n0 PD.t6 1.31518
R54289 PD PD.n1 0.4505
R54290 PD.n6 PD 0.00642105
R54291 PD.n4 PD 0.00405263
R54292 PD.n0 PD 0.001225
R54293 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_4.PLUS.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_4.PLUS.t1 22.3936
R54294 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_1.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D.n0 1.15854
R54295 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D.t0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D.n0 0.5465
R54296 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D.n0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D.t1 0.5465
R54297 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.D GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S.n0 1.15854
R54298 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S.t1 0.5465
R54299 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S.t0 0.5465
R54300 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_2.D GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S.n0 1.15854
R54301 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S.t0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S.n0 0.5465
R54302 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S.t1 0.5465
C0 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.894376f
C1 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A PD 0.055616f
C2 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.012707f
C3 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVSS 9.648331f
C4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D 0.66544f
C5 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.003886f
C6 GF_NI_BI_T_BASE_0.ndrive_y_<0> GF_NI_BI_T_BASE_0.ndrive_Y_<1> 0.031279f
C7 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.035148f
C8 GF_NI_BI_T_BASE_0.ndrive_Y_<3> GF_NI_BI_T_BASE_0.ndrive_x_<3> 10.302f
C9 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S 2.30509f
C10 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B 2.46651f
C11 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_y_<0> 0.737025f
C12 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS VDD 8.9e-19
C13 IE CS 0.002438f
C14 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB PAD 0.10231f
C15 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVDD 6.99663f
C16 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB VDD 0.135207f
C17 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.007263f
C18 GF_NI_BI_T_BASE_0.pdrive_x_<2> GF_NI_BI_T_BASE_0.pdrive_x_<3> 0.048189f
C19 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 0.002385f
C20 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.ndrive_x_<3> 0.001965f
C21 Y A 0.06578f
C22 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS DVSS 0.053427f
C23 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S 0.060445f
C24 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.ndrive_y_<2> 6.12e-19
C25 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.658049f
C26 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.pdrive_y_<3> 1.53e-19
C27 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 0.01198f
C28 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 0.001011f
C29 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 2.42536f
C30 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB DVSS 17.3344f
C31 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.ndrive_y_<2> 7.22e-19
C32 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.pdrive_x_<3> 0.981343f
C33 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.523505f
C34 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 0.09891f
C35 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.ndrive_Y_<1> 3.42e-19
C36 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS DVDD 0.352022f
C37 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 4.94e-20
C38 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL PDRV0 0.025119f
C39 PAD OE 1.52682f
C40 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z VDD 0.171557f
C41 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 0.324691f
C42 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.504632f
C43 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB DVDD 0.478421f
C44 VDD OE 9.91496f
C45 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.pdrive_x_<1> 5.58e-20
C46 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.pdrive_x_<0> 0.718068f
C47 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.ndrive_y_<0> 0.00714f
C48 GF_NI_BI_T_BASE_0.pdrive_x_<1> GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.925558f
C49 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z CS 0.045524f
C50 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D VDD 0.17922f
C51 GF_NI_BI_T_BASE_0.pdrive_y_<2> PAD 10.1896f
C52 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.00192f
C53 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S 0.08422f
C54 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVSS 5.60287f
C55 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.pdrive_y_<1> 1.53e-19
C56 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 0.01198f
C57 DVSS OE 3.49109f
C58 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z PU 0.05345f
C59 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_y_<3> 0.737025f
C60 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 0.026278f
C61 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.035199f
C62 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.ndrive_x_<0> 0.033783f
C63 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D DVSS 0.663936f
C64 OE PU 1.84835f
C65 GF_NI_BI_T_BASE_0.ndrive_Y_<1> GF_NI_BI_T_BASE_0.ndrive_x_<1> 14.8135f
C66 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS PDRV0 0.017469f
C67 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D PU 2.31e-19
C68 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.039646f
C69 GF_NI_BI_T_BASE_0.pdrive_y_<2> DVSS 2.5147f
C70 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVDD 3.53635f
C71 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL A 5.38e-19
C72 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S 0.328757f
C73 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS VDD 1.56815f
C74 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S 0.329817f
C75 DVDD OE 7.68857f
C76 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 0.003533f
C77 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.007532f
C78 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D DVDD 1.95425f
C79 GF_NI_BI_T_BASE_0.pdrive_x_<0> GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.048189f
C80 GF_NI_BI_T_BASE_0.pdrive_y_<0> PAD 10.1953f
C81 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S 0.001012f
C82 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z PD 0.046863f
C83 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 0.505117f
C84 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS DVSS 1.07738f
C85 GF_NI_BI_T_BASE_0.pdrive_y_<2> DVDD 16.7894f
C86 PAD VDD 1.40781f
C87 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB 1.47047f
C88 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_y_<1> 0.737025f
C89 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 0.026278f
C90 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.035214f
C91 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D PD 1.33e-19
C92 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.pdrive_x_<0> 0.003333f
C93 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN 0.001515f
C94 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.pdrive_x_<0> 4.33e-19
C95 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN OE 0.032111f
C96 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.ndrive_x_<3> 0.01433f
C97 GF_NI_BI_T_BASE_0.pdrive_y_<0> DVSS 2.40379f
C98 GF_NI_BI_T_BASE_0.pdrive_x_<3> GF_NI_BI_T_BASE_0.ndrive_Y_<3> 4.4e-19
C99 GF_NI_BI_T_BASE_0.pdrive_y_<2> GF_NI_BI_T_BASE_0.pdrive_y_<3> 0.124712f
C100 PAD DVSS 0.239006p
C101 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS DVDD 5.16559f
C102 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S OE 2.94e-19
C103 PDRV0 OE 0.526899f
C104 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S OE 0.001031f
C105 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D 3.11e-20
C106 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S 0.329551f
C107 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D PDRV0 9.62e-20
C108 DVSS VDD 31.77f
C109 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D 0.575641f
C110 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S 0.014194f
C111 VDD PU 3.27456f
C112 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS PD 0.106114f
C113 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B SL 1.61e-19
C114 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.ndrive_Y_<3> 0.003293f
C115 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D 1.21e-19
C116 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 0.505117f
C117 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.ndrive_x_<1> 6.12e-19
C118 PDRV1 CS 0.039881f
C119 GF_NI_BI_T_BASE_0.pdrive_y_<0> DVDD 18.047901f
C120 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.pdrive_y_<2> 0.026792f
C121 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.pdrive_x_<3> 0.00224f
C122 DVDD PAD 0.310183p
C123 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.051146f
C124 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.003589f
C125 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_y_<2> 1.11498f
C126 DVDD VDD 49.6715f
C127 DVSS PU 6.93148f
C128 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.ndrive_Y_<1> 0.001369f
C129 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS PDRV0 0.195056f
C130 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D 0.316661f
C131 GF_NI_BI_T_BASE_0.pdrive_y_<3> PAD 10.1904f
C132 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.00138f
C133 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D 3.68e-20
C134 OE A 7.46897f
C135 VDD PD 4.66088f
C136 DVDD DVSS 0.360357p
C137 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S 0.003533f
C138 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D 0.217321f
C139 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN PAD 0.227696f
C140 DVDD PU 3.58093f
C141 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S PAD 0.005824f
C142 GF_NI_BI_T_BASE_0.ndrive_Y_<1> GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.13555f
C143 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN VDD 0.415098f
C144 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S PAD 0.289643f
C145 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S DVSS 0.758941f
C146 DVSS PD 6.47201f
C147 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.051146f
C148 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.pdrive_x_<0> 0.002263f
C149 GF_NI_BI_T_BASE_0.pdrive_y_<3> DVSS 2.51644f
C150 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S VDD 0.290069f
C151 VDD PDRV0 2.40295f
C152 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D DVSS 4.62523f
C153 PU PD 0.774032f
C154 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 2.21763f
C155 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_y_<0> 1.12772f
C156 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN DVSS 2.65347f
C157 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 4.43546f
C158 GF_NI_BI_T_BASE_0.pdrive_x_<1> GF_NI_BI_T_BASE_0.ndrive_Y_<1> 0.668765f
C159 GF_NI_BI_T_BASE_0.pdrive_x_<0> GF_NI_BI_T_BASE_0.ndrive_Y_<1> 0.981139f
C160 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 0.02501f
C161 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.pdrive_y_<1> 0.124934f
C162 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 1.8e-19
C163 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 5.42e-20
C164 GF_NI_BI_T_BASE_0.pdrive_y_<1> PAD 10.1967f
C165 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S DVSS 0.733838f
C166 DVSS PDRV0 2.24294f
C167 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.ndrive_x_<0> 7.02e-19
C168 DVDD PD 2.85463f
C169 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S DVDD 0.355101f
C170 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S DVSS 2.82117f
C171 GF_NI_BI_T_BASE_0.pdrive_y_<3> DVDD 17.9191f
C172 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D DVDD 4.00081f
C173 PDRV0 PU 1.1538f
C174 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.ndrive_Y_<1> 0.360786f
C175 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D DVSS 1.72154f
C176 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S 6.92e-19
C177 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN DVDD 1.7492f
C178 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.ndrive_Y_<1> 0.002206f
C179 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.pdrive_y_<0> 0.020536f
C180 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 2.21936f
C181 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S DVDD 1.06223f
C182 DVDD PDRV0 3.29565f
C183 GF_NI_BI_T_BASE_0.pdrive_y_<1> DVSS 2.57525f
C184 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D DVSS 4.60927f
C185 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.pdrive_y_<3> 2.92427f
C186 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S DVDD 5.23952f
C187 VDD A 3.8089f
C188 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D VDD 0.074173f
C189 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.055041f
C190 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D DVDD 6.16e-19
C191 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<3> 0.864692f
C192 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 2.21816f
C193 PDRV0 PD 7.52e-20
C194 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 0.407297f
C195 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.pdrive_x_<3> 6.39e-19
C196 DVSS A 2.11336f
C197 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D DVSS 2.04024f
C198 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S DVSS 2.85457f
C199 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D DVDD 3.93821f
C200 GF_NI_BI_T_BASE_0.ndrive_y_<2> GF_NI_BI_T_BASE_0.pdrive_y_<2> 0.06919f
C201 GF_NI_BI_T_BASE_0.pdrive_y_<1> DVDD 16.784801f
C202 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S DVSS 2.75596f
C203 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S 1.03718f
C204 PU A 0.097708f
C205 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D PU 0.029892f
C206 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.003319f
C207 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S 0.014957f
C208 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 6.5e-19
C209 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.ndrive_x_<2> 3.42e-19
C210 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S PAD 0.289643f
C211 DVDD A 4.11342f
C212 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.pdrive_x_<0> 9.2e-19
C213 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D DVDD 0.09529f
C214 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S DVDD 5.45873f
C215 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S DVDD 5.61526f
C216 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S VDD 0.002554f
C217 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.05515f
C218 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.858187f
C219 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB 0.001515f
C220 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D PD 0.011323f
C221 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S 0.395973f
C222 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.ndrive_x_<0> 0.002977f
C223 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 4.24e-20
C224 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB 5.44729f
C225 GF_NI_BI_T_BASE_0.ndrive_y_<2> PAD 6.37203f
C226 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.ndrive_Y_<1> 6.85e-19
C227 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S DVSS 2.75548f
C228 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S 1.90189f
C229 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.pdrive_y_<3> 0.020536f
C230 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A SL 5.29e-20
C231 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN A 1.16e-19
C232 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.001819f
C233 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z IE 1.4e-19
C234 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB 0.002247f
C235 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S 2.30331f
C236 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S A 0.001505f
C237 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S PDRV0 0.0011f
C238 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D SL 0.397451f
C239 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.pdrive_y_<1> 2.80754f
C240 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S DVDD 5.23942f
C241 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z CS 0.05398f
C242 GF_NI_BI_T_BASE_0.ndrive_y_<2> DVSS 9.63284f
C243 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D 0.178647f
C244 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 0.01198f
C245 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D CS 9.64e-20
C246 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB PDRV1 4.26e-19
C247 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB OE 0.040755f
C248 GF_NI_BI_T_BASE_0.ndrive_y_<0> GF_NI_BI_T_BASE_0.pdrive_y_<0> 2.38e-19
C249 GF_NI_BI_T_BASE_0.ndrive_y_<0> PAD 5.88153f
C250 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S Y 0.002641f
C251 GF_NI_BI_T_BASE_0.ndrive_y_<2> DVDD 11.7338f
C252 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 9.98e-19
C253 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 0.032032f
C254 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.ndrive_Y_<3> 0.360444f
C255 GF_NI_BI_T_BASE_0.ndrive_y_<0> DVSS 12.183001f
C256 GF_NI_BI_T_BASE_0.ndrive_y_<2> GF_NI_BI_T_BASE_0.pdrive_y_<3> 0.069955f
C257 GF_NI_BI_T_BASE_0.ndrive_y_<2> GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 0.00245f
C258 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.328973f
C259 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S 0.520068f
C260 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 0.01198f
C261 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.80907f
C262 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.005985f
C263 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 0.026278f
C264 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.ndrive_y_<2> 6.12e-19
C265 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S 1.90189f
C266 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.pdrive_y_<1> 0.026792f
C267 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.ndrive_Y_<1> 3.42e-19
C268 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.091634f
C269 GF_NI_BI_T_BASE_0.ndrive_y_<0> DVDD 8.54006f
C270 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.ndrive_y_<2> 1.8828f
C271 GF_NI_BI_T_BASE_0.ndrive_x_<3> PAD 6.09734f
C272 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.ndrive_Y_<1> 3.42e-19
C273 VDD CS 2.82934f
C274 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<2> 0.861977f
C275 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB VDD 0.136728f
C276 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB SL 1.29e-19
C277 DVSS CS 4.28108f
C278 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A PDRV1 0.00363f
C279 GF_NI_BI_T_BASE_0.ndrive_x_<3> DVSS 12.039901f
C280 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.013839f
C281 CS PU 0.371306f
C282 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 0.024516f
C283 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB DVSS 2.65303f
C284 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.544964f
C285 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<3> 0.544964f
C286 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.069442f
C287 GF_NI_BI_T_BASE_0.ndrive_x_<1> PAD 5.87598f
C288 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.pdrive_y_<2> 2.80754f
C289 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 0.34223f
C290 DVDD CS 1.35642f
C291 GF_NI_BI_T_BASE_0.ndrive_x_<3> DVDD 5.83927f
C292 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<0> 0.869906f
C293 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB DVDD 1.30327f
C294 CS PD 4.7968f
C295 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z PDRV1 0.047826f
C296 GF_NI_BI_T_BASE_0.ndrive_x_<1> DVSS 9.78378f
C297 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.ndrive_x_<3> 3.33e-19
C298 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.ndrive_x_<3> 0.039995f
C299 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D OE 9.09e-19
C300 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN 0.011456f
C301 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.544964f
C302 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<0> 0.544964f
C303 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.ndrive_x_<3> 0.007481f
C304 Y SL 0.121675f
C305 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS PDRV1 9.81e-19
C306 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.ndrive_y_<0> 1.8897f
C307 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 0.426986f
C308 PDRV0 CS 0.037684f
C309 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.ndrive_y_<2> 3.7e-19
C310 GF_NI_BI_T_BASE_0.ndrive_x_<1> DVDD 9.370099f
C311 GF_NI_BI_T_BASE_0.pdrive_y_<2> GF_NI_BI_T_BASE_0.pdrive_x_<2> 2.31053f
C312 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.077321f
C313 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB PDRV0 0.006824f
C314 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB 0.005324f
C315 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_Y_<3> 1.11322f
C316 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.pdrive_y_<2> 0.465424f
C317 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B VDD 0.529523f
C318 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN PDRV1 5.15e-19
C319 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D DVSS 4.60821f
C320 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S 7.55e-19
C321 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN PDRV1 0.086411f
C322 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 1.10297f
C323 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 8.486509f
C324 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 3.36825f
C325 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.pdrive_y_<0> 2.92427f
C326 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D CS 0.016805f
C327 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B DVSS 4.77406f
C328 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB OE 0.037408f
C329 GF_NI_BI_T_BASE_0.pdrive_x_<2> PAD 20.8838f
C330 GF_NI_BI_T_BASE_0.pdrive_x_<3> PAD 20.2053f
C331 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.ndrive_x_<3> 1.76852f
C332 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D DVDD 3.93443f
C333 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B PU 0.200243f
C334 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S 0.561221f
C335 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_Y_<1> 1.11846f
C336 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 0.016985f
C337 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL SL 3.57e-19
C338 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD VDD 0.600426f
C339 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.041607f
C340 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.069353f
C341 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B DVDD 2.29153f
C342 GF_NI_BI_T_BASE_0.ndrive_x_<2> PAD 7.42368f
C343 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D DVSS 4.60532f
C344 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 0.00366f
C345 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.pdrive_y_<3> 0.02501f
C346 GF_NI_BI_T_BASE_0.pdrive_x_<3> DVSS 5.56575f
C347 GF_NI_BI_T_BASE_0.pdrive_x_<2> DVSS 4.80498f
C348 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 2.31e-19
C349 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B PD 1.53932f
C350 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.215003f
C351 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD DVSS 1.9996f
C352 w_4468_53342# PDRV1 0.003048f
C353 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.071453f
C354 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.pdrive_x_<0> 2.34844f
C355 GF_NI_BI_T_BASE_0.pdrive_x_<1> PAD 20.890501f
C356 GF_NI_BI_T_BASE_0.pdrive_x_<0> PAD 20.2173f
C357 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD PU 0.052014f
C358 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S VDD 1.4802f
C359 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 1.90189f
C360 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D DVDD 4.00037f
C361 GF_NI_BI_T_BASE_0.ndrive_x_<2> DVSS 11.047901f
C362 GF_NI_BI_T_BASE_0.pdrive_x_<2> DVDD 30.158598f
C363 GF_NI_BI_T_BASE_0.pdrive_x_<3> DVDD 29.843302f
C364 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB PAD 0.1164f
C365 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z IE 0.001596f
C366 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD DVDD 0.606126f
C367 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.pdrive_y_<0> 1.64e-19
C368 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S DVSS 1.23577f
C369 GF_NI_BI_T_BASE_0.ndrive_x_<0> PAD 5.05035f
C370 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB VDD 0.137153f
C371 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S PU 0.021163f
C372 GF_NI_BI_T_BASE_0.pdrive_x_<1> DVSS 4.80913f
C373 GF_NI_BI_T_BASE_0.pdrive_x_<0> DVSS 5.52466f
C374 GF_NI_BI_T_BASE_0.pdrive_x_<3> GF_NI_BI_T_BASE_0.pdrive_y_<3> 2.34446f
C375 GF_NI_BI_T_BASE_0.ndrive_y_<2> GF_NI_BI_T_BASE_0.ndrive_x_<3> 9.95829f
C376 GF_NI_BI_T_BASE_0.ndrive_x_<2> DVDD 15.306601f
C377 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.pdrive_x_<3> 0.718047f
C378 GF_NI_BI_T_BASE_0.pdrive_x_<2> GF_NI_BI_T_BASE_0.pdrive_y_<3> 0.071453f
C379 GF_NI_BI_T_BASE_0.pdrive_x_<2> GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 5.58e-20
C380 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A OE 0.006481f
C381 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD PD 0.013731f
C382 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 0.051023f
C383 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.pdrive_x_<3> 9.56e-19
C384 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S DVDD 0.415966f
C385 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB DVSS 4.8944f
C386 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.ndrive_x_<1> 1.76505f
C387 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 0.08661f
C388 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS PDRV1 0.009499f
C389 GF_NI_BI_T_BASE_0.ndrive_x_<0> DVSS 17.7526f
C390 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.pdrive_y_<3> 0.158648f
C391 GF_NI_BI_T_BASE_0.pdrive_x_<1> DVDD 30.213099f
C392 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 0.001369f
C393 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.184422f
C394 GF_NI_BI_T_BASE_0.pdrive_x_<0> DVDD 29.688698f
C395 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.pdrive_y_<2> 0.06401f
C396 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL 0.247434f
C397 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.ndrive_x_<2> 3.42e-19
C398 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S PD 0.223029f
C399 OE SL 2.07268f
C400 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B A 9.24e-21
C401 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB DVDD 1.73731f
C402 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 0.00366f
C403 GF_NI_BI_T_BASE_0.ndrive_x_<0> DVDD 7.91147f
C404 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.ndrive_x_<2> 1.77749f
C405 GF_NI_BI_T_BASE_0.ndrive_Y_<3> PAD 5.0955f
C406 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z 1.53428f
C407 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.ndrive_y_<0> 0.371612f
C408 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL PDRV1 2.27e-19
C409 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 5.97e-20
C410 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D 1.98091f
C411 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 1.90189f
C412 VDD IE 1.31152f
C413 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.088175f
C414 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.pdrive_x_<3> 8.77e-19
C415 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.pdrive_y_<0> 0.055976f
C416 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A PAD 0.107351f
C417 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN 0.007733f
C418 GF_NI_BI_T_BASE_0.ndrive_Y_<3> DVSS 16.0696f
C419 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 0.211601f
C420 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S 1.29e-20
C421 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A VDD 0.156744f
C422 DVSS IE 1.19482f
C423 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 0.519126f
C424 GF_NI_BI_T_BASE_0.ndrive_y_<0> GF_NI_BI_T_BASE_0.ndrive_x_<1> 10.0071f
C425 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.86434f
C426 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.ndrive_Y_<1> 0.158279f
C427 GF_NI_BI_T_BASE_0.pdrive_x_<1> GF_NI_BI_T_BASE_0.pdrive_y_<1> 2.29406f
C428 GF_NI_BI_T_BASE_0.pdrive_x_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 5.58e-20
C429 GF_NI_BI_T_BASE_0.ndrive_Y_<1> PAD 7.99617f
C430 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D VDD 0.740129f
C431 IE PU 1.65e-19
C432 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 0.002397f
C433 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.ndrive_y_<2> 1.2931f
C434 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS PDRV1 0.047903f
C435 GF_NI_BI_T_BASE_0.ndrive_Y_<3> DVDD 12.3656f
C436 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVSS 11.0223f
C437 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN OE 0.206275f
C438 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S 6.63e-20
C439 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB PDRV1 1.35e-19
C440 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 2.42579f
C441 VDD SL 3.37013f
C442 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS 4.05e-19
C443 DVDD IE 1.1774f
C444 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN OE 0.226999f
C445 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D DVSS 0.378193f
C446 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.pdrive_x_<0> 8.77e-19
C447 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D PU 0.840559f
C448 GF_NI_BI_T_BASE_0.ndrive_Y_<1> DVSS 10.754701f
C449 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.ndrive_Y_<3> 1.27008f
C450 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB OE 0.023843f
C451 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVDD 3.81385f
C452 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z VDD 0.180657f
C453 DVSS SL 3.47057f
C454 IE PD 0.814654f
C455 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.pdrive_y_<2> 0.004504f
C456 PU SL 1.23934f
C457 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.ndrive_x_<0> 1.79768f
C458 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D DVDD 0.162547f
C459 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS VDD 0.001344f
C460 GF_NI_BI_T_BASE_0.ndrive_y_<2> GF_NI_BI_T_BASE_0.pdrive_x_<3> 0.074402f
C461 GF_NI_BI_T_BASE_0.ndrive_Y_<1> DVDD 17.7908f
C462 GF_NI_BI_T_BASE_0.ndrive_y_<2> GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.217482f
C463 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVSS 4.88418f
C464 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.pdrive_y_<3> 0.055976f
C465 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 0.491713f
C466 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.ndrive_x_<1> 6.12e-19
C467 OE PDRV1 2.66488f
C468 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z PU 2.62886f
C469 DVDD SL 3.75991f
C470 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D PD 0.100418f
C471 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D PDRV1 0.002909f
C472 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.835267f
C473 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.pdrive_x_<1> 0.184422f
C474 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS DVSS 0.073995f
C475 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.ndrive_y_<2> 14.653599f
C476 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A 0.5167f
C477 w_4468_53342# OE 0.158111f
C478 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVDD 3.13259f
C479 PD SL 0.002085f
C480 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 1.67859f
C481 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN PAD 0.109854f
C482 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN VDD 0.29195f
C483 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S 0.562071f
C484 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN VDD 0.36641f
C485 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.ndrive_y_<0> 1.29246f
C486 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS DVDD 0.373441f
C487 OE Y 2.47359f
C488 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN SL 9.91e-20
C489 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z PD 2.63281f
C490 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB PAD 0.005919f
C491 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S 0.050642f
C492 GF_NI_BI_T_BASE_0.ndrive_Y_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 3.7e-19
C493 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS PDRV1 0.092117f
C494 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.pdrive_y_<1> 0.064015f
C495 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.ndrive_Y_<3> 1.92044f
C496 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 0.505117f
C497 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN DVSS 2.2585f
C498 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB VDD 0.136965f
C499 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D IE 5.96e-20
C500 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN DVSS 3.77203f
C501 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.ndrive_y_<2> 0.34647f
C502 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.290394f
C503 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.ndrive_Y_<1> 0.463637f
C504 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z PDRV0 1.79e-19
C505 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.ndrive_Y_<1> 1.27145f
C506 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A A 0.001333f
C507 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB 9.573371f
C508 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S 1.67734f
C509 PAD PDRV1 7.17e-21
C510 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB DVSS 2.56716f
C511 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S 1.67734f
C512 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN DVDD 1.75818f
C513 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS OE 5.33e-19
C514 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 3.40047f
C515 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D 0.079431f
C516 VDD PDRV1 3.11946f
C517 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN DVDD 2.35832f
C518 w_4468_53342# PAD 1.7719f
C519 GF_NI_BI_T_BASE_0.ndrive_y_<0> GF_NI_BI_T_BASE_0.pdrive_x_<0> 7.63e-19
C520 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB DVDD 1.30605f
C521 w_4468_53342# VDD 0.007089f
C522 SL A 8.864361f
C523 GF_NI_BI_T_BASE_0.pdrive_x_<3> GF_NI_BI_T_BASE_0.ndrive_x_<3> 7.34e-19
C524 DVSS PDRV1 3.24858f
C525 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 2.42579f
C526 PDRV1 PU 0.034849f
C527 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 0.001033f
C528 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.ndrive_y_<0> 10.427401f
C529 VDD Y 1.78812f
C530 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL OE 0.001094f
C531 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D 0.303391f
C532 w_4468_53342# DVSS 0.22053f
C533 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN 0.712898f
C534 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN PDRV0 0.011436f
C535 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 2.42388f
C536 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.ndrive_x_<3> 0.003209f
C537 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S 1.67859f
C538 GF_NI_BI_T_BASE_0.ndrive_y_<2> GF_NI_BI_T_BASE_0.ndrive_Y_<3> 0.003823f
C539 DVDD PDRV1 4.97419f
C540 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S 4.38e-19
C541 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 2.30393f
C542 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB 5.39405f
C543 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.pdrive_y_<2> 1.53e-19
C544 DVSS Y 0.978702f
C545 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S 0.001643f
C546 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S GF_NI_BI_T_BASE_0.ndrive_Y_<1> 1.90029f
C547 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.00245f
C548 w_4468_53342# DVDD 3.9053f
C549 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 1.28e-19
C550 PU Y 0.228424f
C551 PDRV1 PD 0.032008f
C552 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A VDD 0.606688f
C553 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.ndrive_y_<2> 0.001225f
C554 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS VDD 0.001064f
C555 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.pdrive_y_<1> 0.005045f
C556 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 2.2174f
C557 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.pdrive_x_<0> 6.39e-19
C558 DVDD Y 2.10223f
C559 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVSS 1.44042f
C560 PDRV0 PDRV1 6.88206f
C561 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB OE 0.001064f
C562 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S 2.30471f
C563 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB 0.042012f
C564 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A PU 0.001361f
C565 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.ndrive_x_<0> 0.00719f
C566 w_4468_53342# GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN 0.001159f
C567 PD Y 1.13e-19
C568 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.pdrive_y_<0> 1.53e-19
C569 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL PAD 0.598535f
C570 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_y_<2> 0.737025f
C571 w_4468_53342# GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S 0.001239f
C572 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB A 1.54e-19
C573 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVDD 2.37178f
C574 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL VDD 0.671373f
C575 GF_NI_BI_T_BASE_0.pdrive_x_<1> GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.156934f
C576 GF_NI_BI_T_BASE_0.pdrive_x_<0> GF_NI_BI_T_BASE_0.ndrive_x_<1> 0.074382f
C577 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S 0.561221f
C578 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D PDRV1 0.001902f
C579 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS DVDD 0.43338f
C580 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.pdrive_x_<3> 5.58e-20
C581 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.ndrive_y_<0> 0.001918f
C582 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D GF_NI_BI_T_BASE_0.pdrive_x_<2> 0.86434f
C583 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS 0.035159f
C584 A VSS 12.077827f
C585 SL VSS 12.379984f
C586 Y VSS 4.675856f
C587 PD VSS 14.765371f
C588 PU VSS 11.35394f
C589 CS VSS 9.431071f
C590 IE VSS 1.56335f
C591 PDRV1 VSS 13.508398f
C592 OE VSS 19.974787f
C593 PDRV0 VSS 11.475904f
C594 VDD VSS 0.150513p
C595 DVSS VSS 0.207472p
C596 PAD VSS 96.8862f
C597 DVDD VSS 1.073375p
C598 GF_NI_BI_T_BASE_0.ndrive_x_<3> VSS 26.985743f
C599 GF_NI_BI_T_BASE_0.ndrive_Y_<3> VSS 22.96035f
C600 GF_NI_BI_T_BASE_0.pdrive_y_<3> VSS 21.603668f
C601 GF_NI_BI_T_BASE_0.pdrive_x_<3> VSS 5.376266f
C602 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S VSS 1.797274f
C603 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D VSS 1.300121f
C604 GF_NI_BI_T_BASE_0.pdrive_x_<2> VSS 7.15483f
C605 GF_NI_BI_T_BASE_0.pdrive_y_<2> VSS 20.644226f
C606 GF_NI_BI_T_BASE_0.ndrive_y_<2> VSS 28.465302f
C607 GF_NI_BI_T_BASE_0.ndrive_x_<2> VSS 32.64671f
C608 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D VSS 1.297077f
C609 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S VSS 1.730447f
C610 GF_NI_BI_T_BASE_0.ndrive_x_<1> VSS 32.776463f
C611 GF_NI_BI_T_BASE_0.ndrive_Y_<1> VSS 31.33064f
C612 GF_NI_BI_T_BASE_0.pdrive_y_<1> VSS 21.372349f
C613 GF_NI_BI_T_BASE_0.pdrive_x_<1> VSS 7.13999f
C614 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S VSS 1.731697f
C615 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D VSS 1.297201f
C616 GF_NI_BI_T_BASE_0.pdrive_x_<0> VSS 5.363458f
C617 GF_NI_BI_T_BASE_0.pdrive_y_<0> VSS 22.27423f
C618 GF_NI_BI_T_BASE_0.ndrive_y_<0> VSS 25.177105f
C619 GF_NI_BI_T_BASE_0.ndrive_x_<0> VSS 25.017963f
C620 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D VSS 1.300839f
C621 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S VSS 1.800334f
C622 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB VSS 8.662611f
C623 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL VSS 10.852985f
C624 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A VSS 15.26673f
C625 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S VSS 0.327138f
C626 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB VSS 9.65207f
C627 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN VSS 10.13205f
C628 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB VSS 10.53255f
C629 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN VSS 12.82096f
C630 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB VSS 4.70695f
C631 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN VSS 5.64779f
C632 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D VSS 0.810347f
C633 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS VSS 0.15084f
C634 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS VSS 0.151523f
C635 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS VSS 0.148863f
C636 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS VSS 6.718945f
C637 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S VSS 4.01574f
C638 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A VSS 2.984452f
C639 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S VSS 2.342603f
C640 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D VSS 0.629369f
C641 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D VSS 4.25674f
C642 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D VSS 1.299001f
C643 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B VSS 7.37456f
C644 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD VSS 3.170621f
C645 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z VSS 10.767779f
C646 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z VSS 4.74982f
C647 w_4468_53342# VSS 39.222f
C648 PD.t6 VSS 0.330098f
C649 PD.n0 VSS 0.161778f
C650 PD.n1 VSS 1.42326f
C651 PD.t5 VSS 0.301061f
C652 PD.t1 VSS 0.599977f
C653 PD.n2 VSS 1.00615f
C654 PD.t0 VSS 0.61187f
C655 PD.n3 VSS 0.453604f
C656 PD.t2 VSS 0.700879f
C657 PD.n4 VSS 0.945303f
C658 PD.t4 VSS 0.677816f
C659 PD.t3 VSS 0.684698f
C660 PD.n5 VSS 0.775303f
C661 PD.n6 VSS 0.285615f
C662 PD.n7 VSS 6.7579f
C663 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t1 VSS 0.138169f
C664 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t0 VSS 0.478686f
C665 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t3 VSS 0.476171f
C666 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t2 VSS 0.963705f
C667 A.t0 VSS 1.06886f
C668 A.t2 VSS 1.15581f
C669 A.n0 VSS 1.38467f
C670 A.t1 VSS 0.470715f
C671 A.n1 VSS 1.14038f
C672 A.n2 VSS 10.5601f
C673 A.n3 VSS 1.12803f
C674 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t3 VSS 1.00379f
C675 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t4 VSS 2.03153f
C676 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t1 VSS 0.291265f
C677 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t0 VSS 1.00909f
C678 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.n0 VSS 3.98221f
C679 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t2 VSS 1.00379f
C680 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t5 VSS 2.03153f
C681 PDRV1.n0 VSS 0.046183f
C682 PDRV1.n1 VSS 0.075216f
C683 PDRV1.n2 VSS 0.065406f
C684 PDRV1.n3 VSS 0.075216f
C685 PDRV1.t0 VSS 0.23982f
C686 PDRV1.n4 VSS 0.065406f
C687 PDRV1.n6 VSS 0.055595f
C688 PDRV1.n7 VSS 0.075216f
C689 PDRV1.n8 VSS 0.075216f
C690 PDRV1.n9 VSS 0.024889f
C691 PDRV1.n10 VSS 0.055595f
C692 PDRV1.n11 VSS 0.039243f
C693 PDRV1.t1 VSS 0.690467f
C694 PDRV1.t2 VSS 0.746637f
C695 PDRV1.n12 VSS 0.894481f
C696 PDRV1.n13 VSS 0.053823f
C697 PDRV1.n14 VSS 6.80904f
C698 PDRV1.n15 VSS 0.829167f
C699 PDRV1.n16 VSS 0.030706f
C700 PDRV1.n17 VSS 0.075216f
C701 PDRV1.n18 VSS 0.575569f
C702 PDRV1.n19 VSS 0.35973f
C703 PDRV1.n20 VSS 0.065406f
C704 PDRV1.n21 VSS 0.049054f
C705 PDRV1.n22 VSS 0.049054f
C706 PDRV1.n23 VSS 0.055595f
C707 PDRV1.n24 VSS 0.039243f
C708 PDRV1.n25 VSS 0.039243f
C709 PDRV1.n26 VSS 0.075216f
C710 PDRV1.n27 VSS 0.075216f
C711 PDRV1.n29 VSS 0.575569f
C712 PDRV1.n30 VSS 0.35973f
C713 PDRV1.n31 VSS 0.065406f
C714 PDRV1.n32 VSS 0.049054f
C715 GF_NI_BI_T_BASE_0.ndrive_x_<2>.t1 VSS 0.993106f
C716 GF_NI_BI_T_BASE_0.ndrive_x_<2>.t0 VSS 1.27447f
C717 GF_NI_BI_T_BASE_0.ndrive_x_<2>.n0 VSS 1.65686f
C718 GF_NI_BI_T_BASE_0.ndrive_x_<2>.t2 VSS 0.104886f
C719 GF_NI_BI_T_BASE_0.ndrive_x_<2>.n1 VSS 1.69595f
C720 GF_NI_BI_T_BASE_0.ndrive_x_<2>.t3 VSS 12.2133f
C721 OE.t5 VSS 0.516087f
C722 OE.t10 VSS 0.558071f
C723 OE.n0 VSS 0.668576f
C724 OE.n1 VSS 0.028517f
C725 OE.n2 VSS 0.036509f
C726 OE.n3 VSS 0.048887f
C727 OE.n4 VSS 0.430206f
C728 OE.n6 VSS 0.036665f
C729 OE.n7 VSS 0.048887f
C730 OE.n8 VSS 0.430206f
C731 OE.n9 VSS 0.05622f
C732 OE.n12 VSS 0.036665f
C733 OE.n13 VSS 0.05622f
C734 OE.n14 VSS 0.05622f
C735 OE.n15 VSS 0.029332f
C736 OE.n16 VSS 0.041554f
C737 OE.n17 VSS 0.041554f
C738 OE.n18 VSS 0.029332f
C739 OE.n19 VSS 0.05622f
C740 OE.n20 VSS 0.036665f
C741 OE.n21 VSS 0.048887f
C742 OE.n22 VSS 0.268879f
C743 OE.t2 VSS 0.179253f
C744 OE.n23 VSS 0.268879f
C745 OE.n24 VSS 0.048887f
C746 OE.n25 VSS 0.05622f
C747 OE.n26 VSS 0.05622f
C748 OE.n27 VSS 0.029332f
C749 OE.n28 VSS 0.041554f
C750 OE.n29 VSS 0.041554f
C751 OE.n31 VSS 0.05622f
C752 OE.n32 VSS 0.503198f
C753 OE.t8 VSS 0.516087f
C754 OE.t6 VSS 0.558071f
C755 OE.n33 VSS 0.668576f
C756 OE.n34 VSS 0.06711f
C757 OE.n35 VSS 2.03839f
C758 OE.n36 VSS 0.028517f
C759 OE.n37 VSS 0.036509f
C760 OE.n38 VSS 0.048887f
C761 OE.n39 VSS 0.430206f
C762 OE.n40 VSS 0.029332f
C763 OE.n41 VSS 0.048887f
C764 OE.n42 VSS 0.05622f
C765 OE.n43 VSS 0.05622f
C766 OE.n44 VSS 0.268879f
C767 OE.t1 VSS 0.179253f
C768 OE.n45 VSS 0.430206f
C769 OE.n46 VSS 0.05622f
C770 OE.n47 VSS 0.029332f
C771 OE.n48 VSS 0.041554f
C772 OE.n50 VSS 0.041554f
C773 OE.n51 VSS 0.029332f
C774 OE.n52 VSS 0.05622f
C775 OE.n53 VSS 0.036665f
C776 OE.n54 VSS 0.048887f
C777 OE.n55 VSS 0.268879f
C778 OE.n56 VSS 0.048887f
C779 OE.n57 VSS 0.036665f
C780 OE.n58 VSS 0.036665f
C781 OE.n59 VSS 0.05622f
C782 OE.n60 VSS 0.05622f
C783 OE.n62 VSS 0.041554f
C784 OE.n63 VSS 0.041554f
C785 OE.n65 VSS 0.05622f
C786 OE.n66 VSS 0.503198f
C787 OE.t4 VSS 0.516087f
C788 OE.t9 VSS 0.558071f
C789 OE.n67 VSS 0.668576f
C790 OE.n68 VSS 0.06711f
C791 OE.n69 VSS 1.65083f
C792 OE.n70 VSS 1.77035f
C793 OE.n71 VSS 0.028517f
C794 OE.n72 VSS 0.036509f
C795 OE.n73 VSS 0.048887f
C796 OE.n74 VSS 0.430206f
C797 OE.n76 VSS 0.036665f
C798 OE.n77 VSS 0.048887f
C799 OE.n78 VSS 0.430206f
C800 OE.n79 VSS 0.05622f
C801 OE.n82 VSS 0.036665f
C802 OE.n83 VSS 0.05622f
C803 OE.n84 VSS 0.05622f
C804 OE.n85 VSS 0.029332f
C805 OE.n86 VSS 0.041554f
C806 OE.n87 VSS 0.041554f
C807 OE.n88 VSS 0.029332f
C808 OE.n89 VSS 0.05622f
C809 OE.n90 VSS 0.036665f
C810 OE.n91 VSS 0.048887f
C811 OE.n92 VSS 0.268879f
C812 OE.t0 VSS 0.179253f
C813 OE.n93 VSS 0.268879f
C814 OE.n94 VSS 0.048887f
C815 OE.n95 VSS 0.05622f
C816 OE.n96 VSS 0.05622f
C817 OE.n97 VSS 0.029332f
C818 OE.n98 VSS 0.041554f
C819 OE.n99 VSS 0.041554f
C820 OE.n101 VSS 0.05622f
C821 OE.n102 VSS 0.503198f
C822 OE.t7 VSS 0.516087f
C823 OE.t3 VSS 0.558071f
C824 OE.n103 VSS 0.668576f
C825 OE.n104 VSS 0.06711f
C826 OE.n105 VSS 1.65083f
C827 OE.n106 VSS 1.49371f
C828 OE.n107 VSS 5.33715f
C829 OE.n108 VSS 0.463845f
C830 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t0 VSS 1.34784f
C831 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t1 VSS 1.14179f
C832 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n0 VSS 0.748383f
C833 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t6 VSS 0.437171f
C834 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t7 VSS 0.437171f
C835 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t2 VSS 0.437171f
C836 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t4 VSS 0.437171f
C837 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t3 VSS 0.940081f
C838 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t5 VSS 0.944921f
C839 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n1 VSS 1.00241f
C840 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n2 VSS 0.469225f
C841 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n3 VSS 0.302143f
C842 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n4 VSS 0.302143f
C843 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n5 VSS 0.446667f
C844 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n6 VSS 0.582197f
C845 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t4 VSS 0.536852f
C846 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t3 VSS 0.287306f
C847 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.n0 VSS 0.382086f
C848 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t1 VSS 0.206579f
C849 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t2 VSS 0.528517f
C850 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t5 VSS 1.06955f
C851 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN.t0 VSS 0.505447f
C852 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.n0 VSS 0.131232f
C853 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t2 VSS 0.097441f
C854 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t1 VSS 0.418367f
C855 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t0 VSS 0.035864f
C856 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t1 VSS 0.159919f
C857 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t0 VSS 0.463729f
C858 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n0 VSS 1.04783f
C859 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t3 VSS 0.198371f
C860 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t4 VSS 0.195341f
C861 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n1 VSS 0.973754f
C862 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t2 VSS 0.157997f
C863 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t3 VSS 1.24183f
C864 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t1 VSS 1.23656f
C865 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t0 VSS 1.58691f
C866 GF_NI_BI_T_BASE_0.pdrive_y_<2>.n0 VSS 2.47086f
C867 GF_NI_BI_T_BASE_0.pdrive_y_<2>.n1 VSS 1.25671f
C868 GF_NI_BI_T_BASE_0.pdrive_y_<2>.n2 VSS 0.898858f
C869 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t2 VSS 0.134046f
C870 GF_NI_BI_T_BASE_0.pdrive_y_<2>.t4 VSS 6.27852f
C871 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t1 VSS 0.210383f
C872 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n0 VSS 0.232277f
C873 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n1 VSS 0.046696f
C874 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t0 VSS 0.019531f
C875 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n2 VSS 1.35751f
C876 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t2 VSS 0.033306f
C877 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t1 VSS 1.57587f
C878 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t0 VSS 1.51789f
C879 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t7 VSS 1.25234f
C880 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t3 VSS 1.37161f
C881 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n0 VSS 0.981389f
C882 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t8 VSS 1.25234f
C883 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t6 VSS 1.37161f
C884 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n1 VSS 0.981389f
C885 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n2 VSS 0.25845f
C886 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t2 VSS 1.89864f
C887 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n3 VSS 1.19395f
C888 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t5 VSS 0.631878f
C889 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t4 VSS 0.727229f
C890 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n4 VSS 0.820403f
C891 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t2 VSS 1.55639f
C892 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t0 VSS 1.49904f
C893 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t1 VSS 1.87506f
C894 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t5 VSS 1.23679f
C895 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t4 VSS 1.35457f
C896 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n0 VSS 0.969197f
C897 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t7 VSS 1.23679f
C898 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t8 VSS 1.35457f
C899 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n1 VSS 0.969197f
C900 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n2 VSS 0.255239f
C901 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n3 VSS 1.17912f
C902 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t6 VSS 0.624028f
C903 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t3 VSS 0.718195f
C904 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n4 VSS 0.810212f
C905 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t0 VSS 0.51572f
C906 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t1 VSS 0.181706f
C907 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t2 VSS 0.418935f
C908 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t3 VSS 0.50148f
C909 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t5 VSS 0.284525f
C910 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t4 VSS 0.50148f
C911 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t6 VSS 0.284525f
C912 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n0 VSS 0.726879f
C913 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n1 VSS 0.721995f
C914 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t1 VSS 1.61065f
C915 GF_NI_BI_T_BASE_0.pdrive_x_<3>.n0 VSS 2.36388f
C916 GF_NI_BI_T_BASE_0.pdrive_x_<3>.n1 VSS 1.88831f
C917 GF_NI_BI_T_BASE_0.pdrive_x_<3>.n2 VSS 1.37203f
C918 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t2 VSS 0.99663f
C919 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t3 VSS 0.803601f
C920 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t0 VSS 0.136052f
C921 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t5 VSS 6.08062f
C922 GF_NI_BI_T_BASE_0.pdrive_x_<3>.t4 VSS 6.00179f
C923 GF_NI_BI_T_BASE_0.pdrive_x_<3>.n3 VSS 33.0065f
C924 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t3 VSS 1.01484f
C925 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t4 VSS 0.10226f
C926 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n0 VSS 0.746002f
C927 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t5 VSS 12.126599f
C928 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t1 VSS 1.13289f
C929 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n1 VSS 3.49749f
C930 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n2 VSS 0.805369f
C931 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t2 VSS 2.56725f
C932 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n3 VSS 1.27451f
C933 GF_NI_BI_T_BASE_0.ndrive_y_<2>.t0 VSS 1.30236f
C934 GF_NI_BI_T_BASE_0.ndrive_y_<2>.n4 VSS 1.19632f
C935 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t1 VSS 0.090077f
C936 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t0 VSS 0.265454f
C937 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t2 VSS 0.142651f
C938 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t5 VSS 0.923628f
C939 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t2 VSS 1.86913f
C940 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t7 VSS 0.923628f
C941 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t3 VSS 1.86913f
C942 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.n0 VSS 3.58291f
C943 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t0 VSS 0.361015f
C944 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t1 VSS 0.88331f
C945 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t6 VSS 0.938193f
C946 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.t4 VSS 0.502091f
C947 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN.n1 VSS 0.667727f
C948 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.Z VSS 4.43443f
C949 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A VSS 2.41435f
C950 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t0 VSS 0.457031f
C951 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t1 VSS 0.306336f
C952 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.n0 VSS 0.487855f
C953 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t2 VSS 0.94601f
C954 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t1 VSS 1.21403f
C955 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n0 VSS 1.11518f
C956 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t0 VSS 2.39313f
C957 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t4 VSS 0.095324f
C958 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n1 VSS 0.695405f
C959 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t3 VSS 2.20897f
C960 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n2 VSS 1.03087f
C961 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.n3 VSS 1.18807f
C962 GF_NI_BI_T_BASE_0.ndrive_Y_<3>.t5 VSS 10.826099f
C963 GF_NI_BI_T_BASE_0.pdrive_y_<3>.t3 VSS 1.26189f
C964 GF_NI_BI_T_BASE_0.pdrive_y_<3>.t2 VSS 1.25662f
C965 GF_NI_BI_T_BASE_0.pdrive_y_<3>.t1 VSS 1.61254f
C966 GF_NI_BI_T_BASE_0.pdrive_y_<3>.n0 VSS 2.51077f
C967 GF_NI_BI_T_BASE_0.pdrive_y_<3>.n1 VSS 1.27701f
C968 GF_NI_BI_T_BASE_0.pdrive_y_<3>.n2 VSS 0.913487f
C969 GF_NI_BI_T_BASE_0.pdrive_y_<3>.t0 VSS 0.13621f
C970 GF_NI_BI_T_BASE_0.pdrive_y_<3>.t4 VSS 6.32474f
C971 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t0 VSS 1.29746f
C972 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t1 VSS 1.09911f
C973 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n0 VSS 0.720406f
C974 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t2 VSS 0.420829f
C975 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t3 VSS 0.420829f
C976 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t4 VSS 0.420829f
C977 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t6 VSS 0.420829f
C978 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t5 VSS 0.904937f
C979 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t7 VSS 0.909597f
C980 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n1 VSS 0.964934f
C981 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n2 VSS 0.451683f
C982 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n3 VSS 0.290848f
C983 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n4 VSS 0.290848f
C984 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n5 VSS 0.429969f
C985 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n6 VSS 0.560433f
C986 PDRV0.n0 VSS 0.039234f
C987 PDRV0.t1 VSS 0.552244f
C988 PDRV0.t2 VSS 0.59717f
C989 PDRV0.n1 VSS 0.715417f
C990 PDRV0.n2 VSS 0.043049f
C991 PDRV0.n3 VSS 4.95179f
C992 PDRV0.n4 VSS 0.663178f
C993 PDRV0.n5 VSS 0.052312f
C994 PDRV0.n6 VSS 0.060159f
C995 PDRV0.t0 VSS 0.191811f
C996 PDRV0.n7 VSS 0.052312f
C997 PDRV0.n8 VSS 0.060159f
C998 PDRV0.n9 VSS 0.024559f
C999 PDRV0.n10 VSS 0.060159f
C1000 PDRV0.n11 VSS 0.060159f
C1001 PDRV0.n13 VSS 0.044465f
C1002 PDRV0.n14 VSS 0.060159f
C1003 PDRV0.n15 VSS 0.060159f
C1004 PDRV0.n16 VSS 0.031387f
C1005 PDRV0.n17 VSS 0.031387f
C1006 PDRV0.n18 VSS 0.044465f
C1007 PDRV0.n20 VSS 0.460347f
C1008 PDRV0.n21 VSS 0.287717f
C1009 PDRV0.n22 VSS 0.052312f
C1010 PDRV0.n23 VSS 0.039234f
C1011 PDRV0.n24 VSS 0.039234f
C1012 PDRV0.n25 VSS 0.060159f
C1013 PDRV0.n26 VSS 0.031387f
C1014 PDRV0.n27 VSS 0.044465f
C1015 PDRV0.n28 VSS 0.019906f
C1016 PDRV0.n29 VSS 0.460347f
C1017 PDRV0.n30 VSS 0.287717f
C1018 PDRV0.n31 VSS 0.052312f
C1019 PDRV0.n32 VSS 0.036937f
C1020 Y.t8 VSS 0.039999f
C1021 Y.t6 VSS 0.039999f
C1022 Y.n0 VSS 0.080758f
C1023 Y.n1 VSS 0.046305f
C1024 Y.t7 VSS 0.039999f
C1025 Y.t11 VSS 0.039999f
C1026 Y.n2 VSS 0.080758f
C1027 Y.n3 VSS 0.046305f
C1028 Y.t2 VSS 0.09333f
C1029 Y.t0 VSS 0.09333f
C1030 Y.n4 VSS 0.275451f
C1031 Y.t3 VSS 0.09333f
C1032 Y.t1 VSS 0.09333f
C1033 Y.n5 VSS 0.275451f
C1034 Y.t5 VSS 0.09333f
C1035 Y.t4 VSS 0.09333f
C1036 Y.n6 VSS 0.387786f
C1037 Y.n7 VSS 0.618155f
C1038 Y.n8 VSS 0.388772f
C1039 Y.n9 VSS 1.39079f
C1040 Y.n10 VSS 0.287072f
C1041 Y.n11 VSS 0.29272f
C1042 Y.n12 VSS 0.168405f
C1043 Y.t10 VSS 0.039999f
C1044 Y.t9 VSS 0.039999f
C1045 Y.n13 VSS 0.080763f
C1046 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D VSS 1.19647f
C1047 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t1 VSS 0.063962f
C1048 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t0 VSS 0.300506f
C1049 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t11 VSS 0.169311f
C1050 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t8 VSS 0.221117f
C1051 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n0 VSS 0.251108f
C1052 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t2 VSS 0.169311f
C1053 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t12 VSS 0.221117f
C1054 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n1 VSS 0.249078f
C1055 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t7 VSS 0.169311f
C1056 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t4 VSS 0.221117f
C1057 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n2 VSS 0.249078f
C1058 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t6 VSS 0.169311f
C1059 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t3 VSS 0.221117f
C1060 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n3 VSS 0.249078f
C1061 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t13 VSS 0.169311f
C1062 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t9 VSS 0.221117f
C1063 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n4 VSS 0.249078f
C1064 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t10 VSS 0.169311f
C1065 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t5 VSS 0.221117f
C1066 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n5 VSS 0.249078f
C1067 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t3 VSS 0.93914f
C1068 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t2 VSS 2.37575f
C1069 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t4 VSS 0.094632f
C1070 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n0 VSS 0.690355f
C1071 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t1 VSS 2.19293f
C1072 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n1 VSS 1.02339f
C1073 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n2 VSS 1.17944f
C1074 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t0 VSS 1.20522f
C1075 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.n3 VSS 1.10708f
C1076 GF_NI_BI_T_BASE_0.ndrive_Y_<1>.t5 VSS 11.5531f
C1077 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t0 VSS 1.29746f
C1078 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t1 VSS 1.09911f
C1079 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n0 VSS 0.720406f
C1080 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t3 VSS 0.420829f
C1081 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t5 VSS 0.420829f
C1082 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t4 VSS 0.420829f
C1083 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t7 VSS 0.420829f
C1084 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t2 VSS 0.909597f
C1085 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t6 VSS 0.904937f
C1086 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n1 VSS 0.964934f
C1087 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n2 VSS 0.451683f
C1088 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n3 VSS 0.290848f
C1089 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n4 VSS 0.290848f
C1090 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n5 VSS 0.429969f
C1091 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n6 VSS 0.560433f
C1092 GF_NI_BI_T_BASE_0.ndrive_x_<3>.t1 VSS 3.10443f
C1093 GF_NI_BI_T_BASE_0.ndrive_x_<3>.t0 VSS 0.767595f
C1094 GF_NI_BI_T_BASE_0.ndrive_x_<3>.t2 VSS 0.111079f
C1095 GF_NI_BI_T_BASE_0.ndrive_x_<3>.n0 VSS 1.79609f
C1096 GF_NI_BI_T_BASE_0.ndrive_x_<3>.t3 VSS 12.4708f
C1097 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t1 VSS 1.34784f
C1098 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t0 VSS 1.14179f
C1099 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n0 VSS 0.748383f
C1100 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t6 VSS 0.437171f
C1101 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t3 VSS 0.437171f
C1102 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t2 VSS 0.437171f
C1103 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t5 VSS 0.437171f
C1104 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t7 VSS 0.944921f
C1105 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t4 VSS 0.940081f
C1106 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n1 VSS 1.00241f
C1107 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n2 VSS 0.469225f
C1108 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n3 VSS 0.302143f
C1109 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n4 VSS 0.302143f
C1110 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n5 VSS 0.446667f
C1111 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n6 VSS 0.582197f
C1112 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t0 VSS 1.56917f
C1113 GF_NI_BI_T_BASE_0.pdrive_x_<2>.n0 VSS 2.30162f
C1114 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t2 VSS 0.782832f
C1115 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t3 VSS 0.691979f
C1116 GF_NI_BI_T_BASE_0.pdrive_x_<2>.n1 VSS 1.61579f
C1117 GF_NI_BI_T_BASE_0.pdrive_x_<2>.n2 VSS 1.83962f
C1118 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t1 VSS 0.132547f
C1119 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t5 VSS 5.82992f
C1120 GF_NI_BI_T_BASE_0.pdrive_x_<2>.t4 VSS 5.94087f
C1121 GF_NI_BI_T_BASE_0.pdrive_x_<2>.n3 VSS 32.157803f
C1122 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t1 VSS 0.811404f
C1123 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t4 VSS 0.434237f
C1124 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.n0 VSS 0.574127f
C1125 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t2 VSS 0.798807f
C1126 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t3 VSS 1.61653f
C1127 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN.t0 VSS 0.763937f
C1128 PU.t4 VSS 0.431002f
C1129 PU.t3 VSS 0.435378f
C1130 PU.n0 VSS 0.492992f
C1131 PU.n1 VSS 0.036137f
C1132 PU.t1 VSS 0.104731f
C1133 PU.n2 VSS 0.101125f
C1134 PU.t5 VSS 0.261445f
C1135 PU.t2 VSS 0.470018f
C1136 PU.n3 VSS 0.46747f
C1137 PU.n4 VSS 0.376861f
C1138 PU.t0 VSS 0.188953f
C1139 PU.n5 VSS 0.844412f
C1140 PU.n6 VSS 5.01223f
C1141 PU.t6 VSS 0.209899f
C1142 PU.n7 VSS 0.10287f
C1143 PU.n8 VSS 5.28119f
C1144 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n0 VSS 0.560838f
C1145 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n1 VSS 0.34898f
C1146 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t8 VSS 0.071338f
C1147 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t7 VSS 0.071338f
C1148 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n2 VSS 0.14835f
C1149 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t13 VSS 0.445267f
C1150 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t15 VSS 0.314023f
C1151 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n3 VSS 0.431502f
C1152 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n4 VSS 0.441196f
C1153 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t14 VSS 0.473114f
C1154 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t4 VSS 0.0925f
C1155 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t3 VSS 0.092507f
C1156 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t11 VSS 0.066482f
C1157 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t12 VSS 0.067162f
C1158 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n5 VSS 0.738258f
C1159 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n6 VSS 0.349573f
C1160 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t2 VSS 0.065232f
C1161 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t1 VSS 0.047558f
C1162 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t0 VSS 0.047558f
C1163 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n7 VSS 0.215887f
C1164 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n8 VSS 0.625782f
C1165 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t6 VSS 0.219696f
C1166 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t5 VSS 0.071338f
C1167 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n9 VSS 0.097229f
C1168 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t10 VSS 0.051125f
C1169 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t9 VSS 0.051125f
C1170 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n10 VSS 0.199205f
C1171 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n11 VSS 0.577838f
C1172 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n12 VSS 0.977898f
C1173 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n13 VSS 0.58506f
C1174 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n14 VSS 0.199987f
C1175 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t1 VSS 3.96081f
C1176 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t2 VSS 0.800753f
C1177 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t3 VSS 0.70782f
C1178 GF_NI_BI_T_BASE_0.pdrive_x_<0>.n0 VSS 1.65277f
C1179 GF_NI_BI_T_BASE_0.pdrive_x_<0>.n1 VSS 1.88173f
C1180 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t0 VSS 0.135582f
C1181 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t4 VSS 5.98219f
C1182 GF_NI_BI_T_BASE_0.pdrive_x_<0>.t5 VSS 6.05673f
C1183 GF_NI_BI_T_BASE_0.pdrive_x_<0>.n2 VSS 32.894302f
C1184 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t1 VSS 0.245849f
C1185 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t5 VSS 0.975903f
C1186 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t2 VSS 1.12317f
C1187 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n0 VSS 1.10814f
C1188 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t7 VSS 0.975903f
C1189 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t9 VSS 1.12317f
C1190 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n1 VSS 1.10814f
C1191 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n2 VSS 2.87718f
C1192 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t8 VSS 0.975903f
C1193 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t6 VSS 1.12317f
C1194 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n3 VSS 1.10814f
C1195 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n4 VSS 2.37169f
C1196 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t3 VSS 0.975903f
C1197 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t4 VSS 1.12317f
C1198 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n5 VSS 1.10814f
C1199 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.n6 VSS 2.10472f
C1200 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB.t0 VSS 0.72451f
C1201 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t0 VSS 1.57596f
C1202 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t2 VSS 1.51789f
C1203 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t1 VSS 1.89864f
C1204 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t8 VSS 1.25234f
C1205 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t7 VSS 1.37161f
C1206 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n0 VSS 0.981389f
C1207 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t4 VSS 1.25234f
C1208 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t5 VSS 1.37161f
C1209 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n1 VSS 0.981389f
C1210 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n2 VSS 0.25845f
C1211 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n3 VSS 1.19395f
C1212 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t3 VSS 0.631878f
C1213 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t6 VSS 0.727229f
C1214 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n4 VSS 0.820403f
C1215 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB.t0 VSS 0.239584f
C1216 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB.t1 VSS 0.830038f
C1217 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB.t2 VSS 0.825677f
C1218 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB.t3 VSS 1.67106f
C1219 GF_NI_BI_T_BASE_0.ndrive_x_<1>.t1 VSS 3.19703f
C1220 GF_NI_BI_T_BASE_0.ndrive_x_<1>.t0 VSS 0.790491f
C1221 GF_NI_BI_T_BASE_0.ndrive_x_<1>.t2 VSS 0.114393f
C1222 GF_NI_BI_T_BASE_0.ndrive_x_<1>.n0 VSS 1.84967f
C1223 GF_NI_BI_T_BASE_0.ndrive_x_<1>.t3 VSS 12.944799f
C1224 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t3 VSS 0.133905f
C1225 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t1 VSS 0.152948f
C1226 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t2 VSS 0.097738f
C1227 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t6 VSS 0.036976f
C1228 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t0 VSS 0.097639f
C1229 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t5 VSS 0.113596f
C1230 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t4 VSS 0.086707f
C1231 GF_NI_BI_T_BASE_0.pdrive_y_<1>.t3 VSS 4.07002f
C1232 GF_NI_BI_T_BASE_0.pdrive_y_<1>.n0 VSS 2.16219f
C1233 GF_NI_BI_T_BASE_0.pdrive_y_<1>.t1 VSS 0.90553f
C1234 GF_NI_BI_T_BASE_0.pdrive_y_<1>.t2 VSS 0.905248f
C1235 GF_NI_BI_T_BASE_0.pdrive_y_<1>.t0 VSS 0.134451f
C1236 GF_NI_BI_T_BASE_0.pdrive_y_<1>.t4 VSS 6.29957f
C1237 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t2 VSS 2.30771f
C1238 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t3 VSS 3.87089f
C1239 GF_NI_BI_T_BASE_0.pdrive_x_<1>.n0 VSS 1.83972f
C1240 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t1 VSS 0.782923f
C1241 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t0 VSS 0.132551f
C1242 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t5 VSS 5.83096f
C1243 GF_NI_BI_T_BASE_0.pdrive_x_<1>.t4 VSS 5.94093f
C1244 GF_NI_BI_T_BASE_0.pdrive_x_<1>.n1 VSS 32.1564f
C1245 GF_NI_BI_T_BASE_0.pdrive_y_<0>.n0 VSS 2.19038f
C1246 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t1 VSS 4.1233f
C1247 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t2 VSS 0.917535f
C1248 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t3 VSS 0.917053f
C1249 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t0 VSS 0.136211f
C1250 GF_NI_BI_T_BASE_0.pdrive_y_<0>.t4 VSS 6.32639f
C1251 PAD.t21 VSS 0.012461f
C1252 PAD.t4 VSS 0.028954f
C1253 PAD.n0 VSS 0.03269f
C1254 PAD.n1 VSS 0.037321f
C1255 PAD.n2 VSS 0.026054f
C1256 PAD.n3 VSS 0.013705f
C1257 PAD.t3 VSS 0.012461f
C1258 PAD.t5 VSS 0.012461f
C1259 PAD.n4 VSS 0.026495f
C1260 PAD.n5 VSS 0.030045f
C1261 PAD.n6 VSS 0.030045f
C1262 PAD.n7 VSS 0.026054f
C1263 PAD.n8 VSS 0.018382f
C1264 PAD.n9 VSS 0.024675f
C1265 PAD.n10 VSS 10.1417f
C1266 PAD.n11 VSS 12.772201f
C1267 PAD.n12 VSS 13.1467f
C1268 PAD.n13 VSS 14.5427f
C1269 PAD.n14 VSS 0.043273f
C1270 PAD.n15 VSS 0.062274f
C1271 PAD.n16 VSS 0.039761f
C1272 PAD.n17 VSS 0.069765f
C1273 PAD.n18 VSS 0.039761f
C1274 PAD.n19 VSS 0.069765f
C1275 PAD.n20 VSS 0.157866f
C1276 PAD.n21 VSS 0.596934f
C1277 PAD.n22 VSS 0.039258f
C1278 PAD.n23 VSS 0.029919f
C1279 PAD.n24 VSS 0.039258f
C1280 PAD.n25 VSS 0.029919f
C1281 PAD.n26 VSS 0.030555f
C1282 PAD.n27 VSS 0.042895f
C1283 PAD.n28 VSS 0.049115f
C1284 PAD.n29 VSS 0.029436f
C1285 PAD.n30 VSS 0.049115f
C1286 PAD.n31 VSS 0.029436f
C1287 PAD.n32 VSS 0.448934f
C1288 PAD.n74 VSS 0.023109f
C1289 PAD.n75 VSS 0.023109f
C1290 PAD.n76 VSS 0.036461f
C1291 PAD.n77 VSS 0.036461f
C1292 PAD.n78 VSS 0.036461f
C1293 PAD.n79 VSS 0.036461f
C1294 PAD.n80 VSS 0.036461f
C1295 PAD.n81 VSS 0.036461f
C1296 PAD.n82 VSS 0.036461f
C1297 PAD.n83 VSS 0.036461f
C1298 PAD.n84 VSS 0.036461f
C1299 PAD.n85 VSS 0.036461f
C1300 PAD.n86 VSS 0.036461f
C1301 PAD.n87 VSS 0.036461f
C1302 PAD.n88 VSS 0.036461f
C1303 PAD.n89 VSS 0.036461f
C1304 PAD.n90 VSS 0.036461f
C1305 PAD.n91 VSS 0.036461f
C1306 PAD.n92 VSS 0.036461f
C1307 PAD.n93 VSS 0.036461f
C1308 PAD.n94 VSS 0.036461f
C1309 PAD.n95 VSS 0.036461f
C1310 PAD.n96 VSS 0.036461f
C1311 PAD.n97 VSS 0.036461f
C1312 PAD.n98 VSS 0.036461f
C1313 PAD.n99 VSS 0.036461f
C1314 PAD.n100 VSS 0.036461f
C1315 PAD.n101 VSS 0.036461f
C1316 PAD.n102 VSS 0.036461f
C1317 PAD.n103 VSS 0.036461f
C1318 PAD.n104 VSS 0.036461f
C1319 PAD.n105 VSS 0.036461f
C1320 PAD.n106 VSS 0.036461f
C1321 PAD.n107 VSS 0.036461f
C1322 PAD.n108 VSS 0.036461f
C1323 PAD.n109 VSS 0.036461f
C1324 PAD.n110 VSS 0.036461f
C1325 PAD.n111 VSS 0.036461f
C1326 PAD.n112 VSS 0.036461f
C1327 PAD.n113 VSS 0.036461f
C1328 PAD.n114 VSS 0.036461f
C1329 PAD.n115 VSS 0.036461f
C1330 PAD.n117 VSS 0.036461f
C1331 PAD.n118 VSS 0.036461f
C1332 PAD.n119 VSS 0.023109f
C1333 PAD.n120 VSS 0.03338f
C1334 PAD.n121 VSS 0.036461f
C1335 PAD.n122 VSS 0.036461f
C1336 PAD.n123 VSS 0.036461f
C1337 PAD.n124 VSS 0.036461f
C1338 PAD.n126 VSS 0.036461f
C1339 PAD.n127 VSS 0.036461f
C1340 PAD.n128 VSS 0.036461f
C1341 PAD.n130 VSS 0.036461f
C1342 PAD.n131 VSS 0.036461f
C1343 PAD.n132 VSS 0.036461f
C1344 PAD.n133 VSS 0.036461f
C1345 PAD.n134 VSS 0.036461f
C1346 PAD.n135 VSS 0.036461f
C1347 PAD.n136 VSS 0.036461f
C1348 PAD.n138 VSS 0.036461f
C1349 PAD.n139 VSS 0.036461f
C1350 PAD.n140 VSS 0.036461f
C1351 PAD.n142 VSS 0.036461f
C1352 PAD.n143 VSS 0.036461f
C1353 PAD.n144 VSS 0.036461f
C1354 PAD.n145 VSS 0.036461f
C1355 PAD.n146 VSS 0.036461f
C1356 PAD.n147 VSS 0.036461f
C1357 PAD.n148 VSS 0.036461f
C1358 PAD.n150 VSS 0.036461f
C1359 PAD.n151 VSS 0.036461f
C1360 PAD.n152 VSS 0.036461f
C1361 PAD.n154 VSS 0.036461f
C1362 PAD.n155 VSS 0.036461f
C1363 PAD.n156 VSS 0.036461f
C1364 PAD.n157 VSS 0.036461f
C1365 PAD.n158 VSS 0.036461f
C1366 PAD.n159 VSS 0.036461f
C1367 PAD.n160 VSS 0.036461f
C1368 PAD.n162 VSS 0.036461f
C1369 PAD.n163 VSS 0.036461f
C1370 PAD.n164 VSS 0.036461f
C1371 PAD.n166 VSS 0.036461f
C1372 PAD.n167 VSS 0.036461f
C1373 PAD.n168 VSS 0.036461f
C1374 PAD.n169 VSS 0.036461f
C1375 PAD.n170 VSS 0.036461f
C1376 PAD.n171 VSS 0.036461f
C1377 PAD.n172 VSS 0.036461f
C1378 PAD.n174 VSS 0.036461f
C1379 PAD.n175 VSS 0.036461f
C1380 PAD.n176 VSS 0.036461f
C1381 PAD.n178 VSS 0.036461f
C1382 PAD.n179 VSS 0.036461f
C1383 PAD.n180 VSS 0.036461f
C1384 PAD.n181 VSS 0.036461f
C1385 PAD.n182 VSS 0.036461f
C1386 PAD.n183 VSS 0.036461f
C1387 PAD.n184 VSS 0.036461f
C1388 PAD.n186 VSS 0.036461f
C1389 PAD.n187 VSS 0.036461f
C1390 PAD.n188 VSS 0.036461f
C1391 PAD.n190 VSS 0.036461f
C1392 PAD.n191 VSS 0.036461f
C1393 PAD.n192 VSS 0.036461f
C1394 PAD.n193 VSS 0.036461f
C1395 PAD.n194 VSS 0.036461f
C1396 PAD.n195 VSS 0.036461f
C1397 PAD.n196 VSS 0.036461f
C1398 PAD.n198 VSS 0.036461f
C1399 PAD.n199 VSS 0.036461f
C1400 PAD.n200 VSS 0.036461f
C1401 PAD.n202 VSS 0.036461f
C1402 PAD.n203 VSS 0.036461f
C1403 PAD.n204 VSS 0.036461f
C1404 PAD.n205 VSS 0.036461f
C1405 PAD.n206 VSS 0.036461f
C1406 PAD.n207 VSS 0.036461f
C1407 PAD.n208 VSS 0.036461f
C1408 PAD.n210 VSS 0.036461f
C1409 PAD.n211 VSS 0.036461f
C1410 PAD.n212 VSS 0.036461f
C1411 PAD.n214 VSS 0.036461f
C1412 PAD.n215 VSS 0.036461f
C1413 PAD.n216 VSS 0.036461f
C1414 PAD.n217 VSS 0.036461f
C1415 PAD.n218 VSS 0.036461f
C1416 PAD.n219 VSS 0.036461f
C1417 PAD.n220 VSS 0.036461f
C1418 PAD.n222 VSS 0.036461f
C1419 PAD.n223 VSS 0.036461f
C1420 PAD.n224 VSS 0.036461f
C1421 PAD.n226 VSS 0.036461f
C1422 PAD.n227 VSS 0.036461f
C1423 PAD.n228 VSS 0.036461f
C1424 PAD.n229 VSS 0.036461f
C1425 PAD.n230 VSS 0.036461f
C1426 PAD.n231 VSS 0.036461f
C1427 PAD.n232 VSS 0.036461f
C1428 PAD.n234 VSS 0.036461f
C1429 PAD.n235 VSS 0.036461f
C1430 PAD.n236 VSS 0.036461f
C1431 PAD.n238 VSS 0.036461f
C1432 PAD.n239 VSS 0.036461f
C1433 PAD.n240 VSS 0.036461f
C1434 PAD.n241 VSS 0.036461f
C1435 PAD.n242 VSS 0.036461f
C1436 PAD.n243 VSS 0.036461f
C1437 PAD.n244 VSS 0.036461f
C1438 PAD.n246 VSS 0.036461f
C1439 PAD.n247 VSS 0.036461f
C1440 PAD.n248 VSS 0.036461f
C1441 PAD.n250 VSS 0.036461f
C1442 PAD.n251 VSS 0.036461f
C1443 PAD.n252 VSS 0.036461f
C1444 PAD.n253 VSS 0.036461f
C1445 PAD.n254 VSS 0.036461f
C1446 PAD.n255 VSS 0.036461f
C1447 PAD.n256 VSS 0.036461f
C1448 PAD.n258 VSS 0.036461f
C1449 PAD.n259 VSS 0.036461f
C1450 PAD.n260 VSS 0.036461f
C1451 PAD.n262 VSS 0.036461f
C1452 PAD.n263 VSS 0.036461f
C1453 PAD.n264 VSS 0.036461f
C1454 PAD.n265 VSS 0.036461f
C1455 PAD.n266 VSS 0.036461f
C1456 PAD.n267 VSS 0.036461f
C1457 PAD.n268 VSS 0.036461f
C1458 PAD.n270 VSS 0.036461f
C1459 PAD.n271 VSS 0.036461f
C1460 PAD.n272 VSS 0.036461f
C1461 PAD.n274 VSS 0.036461f
C1462 PAD.n275 VSS 0.036461f
C1463 PAD.n276 VSS 0.036461f
C1464 PAD.n277 VSS 0.036461f
C1465 PAD.n278 VSS 0.036461f
C1466 PAD.n279 VSS 0.036461f
C1467 PAD.n280 VSS 0.036461f
C1468 PAD.n282 VSS 0.036461f
C1469 PAD.n283 VSS 0.036461f
C1470 PAD.n284 VSS 0.036461f
C1471 PAD.n286 VSS 0.036461f
C1472 PAD.n287 VSS 0.036461f
C1473 PAD.n288 VSS 0.036461f
C1474 PAD.n289 VSS 0.036461f
C1475 PAD.n290 VSS 0.036461f
C1476 PAD.n291 VSS 0.036461f
C1477 PAD.n292 VSS 0.036461f
C1478 PAD.n294 VSS 0.036461f
C1479 PAD.n295 VSS 0.036461f
C1480 PAD.n296 VSS 0.036461f
C1481 PAD.n298 VSS 0.036461f
C1482 PAD.n299 VSS 0.036461f
C1483 PAD.n300 VSS 0.036461f
C1484 PAD.n301 VSS 0.036461f
C1485 PAD.n302 VSS 0.036461f
C1486 PAD.n303 VSS 0.036461f
C1487 PAD.n304 VSS 0.036461f
C1488 PAD.n306 VSS 0.036461f
C1489 PAD.n307 VSS 0.036461f
C1490 PAD.n308 VSS 0.036461f
C1491 PAD.n310 VSS 0.036461f
C1492 PAD.n311 VSS 0.036461f
C1493 PAD.n312 VSS 0.036461f
C1494 PAD.n313 VSS 0.036461f
C1495 PAD.n314 VSS 0.036461f
C1496 PAD.n315 VSS 0.036461f
C1497 PAD.n316 VSS 0.036461f
C1498 PAD.n318 VSS 0.036461f
C1499 PAD.n319 VSS 0.036461f
C1500 PAD.n320 VSS 0.036461f
C1501 PAD.n322 VSS 0.036461f
C1502 PAD.n323 VSS 0.036461f
C1503 PAD.n324 VSS 0.036461f
C1504 PAD.n325 VSS 0.036461f
C1505 PAD.n326 VSS 0.036461f
C1506 PAD.n327 VSS 0.036461f
C1507 PAD.n328 VSS 0.036461f
C1508 PAD.n330 VSS 0.036461f
C1509 PAD.n331 VSS 0.036461f
C1510 PAD.n332 VSS 0.036461f
C1511 PAD.n334 VSS 0.036461f
C1512 PAD.n335 VSS 0.036461f
C1513 PAD.n336 VSS 0.036461f
C1514 PAD.n337 VSS 0.036461f
C1515 PAD.n338 VSS 0.036461f
C1516 PAD.n339 VSS 0.036461f
C1517 PAD.n340 VSS 0.036461f
C1518 PAD.n342 VSS 0.036461f
C1519 PAD.n343 VSS 0.036461f
C1520 PAD.n344 VSS 0.036461f
C1521 PAD.n346 VSS 0.036461f
C1522 PAD.n347 VSS 0.036461f
C1523 PAD.n348 VSS 0.036461f
C1524 PAD.n349 VSS 0.036461f
C1525 PAD.n350 VSS 0.036461f
C1526 PAD.n351 VSS 0.036461f
C1527 PAD.n352 VSS 0.036461f
C1528 PAD.n354 VSS 0.036461f
C1529 PAD.n355 VSS 0.036461f
C1530 PAD.n356 VSS 0.036461f
C1531 PAD.n358 VSS 0.036461f
C1532 PAD.n359 VSS 0.036461f
C1533 PAD.n360 VSS 0.036461f
C1534 PAD.n361 VSS 0.036461f
C1535 PAD.n362 VSS 0.036461f
C1536 PAD.n363 VSS 0.036461f
C1537 PAD.n364 VSS 0.036461f
C1538 PAD.n366 VSS 0.023109f
C1539 PAD.n367 VSS 0.537734f
C1540 PAD.n368 VSS 0.069765f
C1541 PAD.n369 VSS 0.069765f
C1542 PAD.n370 VSS 0.032141f
C1543 PAD.n371 VSS 0.036008f
C1544 PAD.n372 VSS 0.036008f
C1545 PAD.n373 VSS 0.315733f
C1546 PAD.n415 VSS 0.023109f
C1547 PAD.n416 VSS 0.023109f
C1548 PAD.n417 VSS 0.029436f
C1549 PAD.n418 VSS 0.656134f
C1550 PAD.n419 VSS 0.429201f
C1551 PAD.n420 VSS 0.036461f
C1552 PAD.n421 VSS 0.036461f
C1553 PAD.n422 VSS 0.033984f
C1554 PAD.n423 VSS 0.049115f
C1555 PAD.n424 VSS 0.049115f
C1556 PAD.n425 VSS 0.611734f
C1557 PAD.n426 VSS 0.069765f
C1558 PAD.n427 VSS 0.039761f
C1559 PAD.n428 VSS 0.069765f
C1560 PAD.n429 VSS 0.039761f
C1561 PAD.n430 VSS 0.046286f
C1562 PAD.n431 VSS 0.039761f
C1563 PAD.n432 VSS 0.039761f
C1564 PAD.n433 VSS 0.611734f
C1565 PAD.n434 VSS 0.513067f
C1566 PAD.n435 VSS 0.606801f
C1567 PAD.n436 VSS 0.029436f
C1568 PAD.n437 VSS 0.029436f
C1569 PAD.n438 VSS 0.036461f
C1570 PAD.n439 VSS 0.036461f
C1571 PAD.n440 VSS 0.036461f
C1572 PAD.n442 VSS 0.036461f
C1573 PAD.n443 VSS 0.036461f
C1574 PAD.n444 VSS 0.036461f
C1575 PAD.n446 VSS 0.036461f
C1576 PAD.n447 VSS 0.036461f
C1577 PAD.n448 VSS 0.036461f
C1578 PAD.n450 VSS 0.036461f
C1579 PAD.n451 VSS 0.036461f
C1580 PAD.n452 VSS 0.036461f
C1581 PAD.n454 VSS 0.036461f
C1582 PAD.n455 VSS 0.036461f
C1583 PAD.n456 VSS 0.036461f
C1584 PAD.n458 VSS 0.036461f
C1585 PAD.n459 VSS 0.036461f
C1586 PAD.n460 VSS 0.036461f
C1587 PAD.n462 VSS 0.036461f
C1588 PAD.n463 VSS 0.036461f
C1589 PAD.n464 VSS 0.036461f
C1590 PAD.n466 VSS 0.036461f
C1591 PAD.n467 VSS 0.036461f
C1592 PAD.n468 VSS 0.036461f
C1593 PAD.n470 VSS 0.036461f
C1594 PAD.n471 VSS 0.036461f
C1595 PAD.n472 VSS 0.036461f
C1596 PAD.n474 VSS 0.036461f
C1597 PAD.n475 VSS 0.036461f
C1598 PAD.n476 VSS 0.036461f
C1599 PAD.n478 VSS 0.036461f
C1600 PAD.n479 VSS 0.036461f
C1601 PAD.n480 VSS 0.036461f
C1602 PAD.n482 VSS 0.036461f
C1603 PAD.n483 VSS 0.036461f
C1604 PAD.n484 VSS 0.036461f
C1605 PAD.n486 VSS 0.036461f
C1606 PAD.n487 VSS 0.036461f
C1607 PAD.n488 VSS 0.036461f
C1608 PAD.n490 VSS 0.036461f
C1609 PAD.n491 VSS 0.036461f
C1610 PAD.n492 VSS 0.036461f
C1611 PAD.n494 VSS 0.036461f
C1612 PAD.n495 VSS 0.036461f
C1613 PAD.n496 VSS 0.036461f
C1614 PAD.n498 VSS 0.036461f
C1615 PAD.n499 VSS 0.036461f
C1616 PAD.n500 VSS 0.036461f
C1617 PAD.n502 VSS 0.036461f
C1618 PAD.n503 VSS 0.036461f
C1619 PAD.n504 VSS 0.036461f
C1620 PAD.n506 VSS 0.036461f
C1621 PAD.n507 VSS 0.036461f
C1622 PAD.n508 VSS 0.036461f
C1623 PAD.n510 VSS 0.036461f
C1624 PAD.n511 VSS 0.036461f
C1625 PAD.n512 VSS 0.036461f
C1626 PAD.n514 VSS 0.036461f
C1627 PAD.n515 VSS 0.036461f
C1628 PAD.n516 VSS 0.036461f
C1629 PAD.n518 VSS 0.036461f
C1630 PAD.n519 VSS 0.036461f
C1631 PAD.n520 VSS 0.036461f
C1632 PAD.n521 VSS 0.03338f
C1633 PAD.n522 VSS 0.023109f
C1634 PAD.n523 VSS 0.023109f
C1635 PAD.n525 VSS 0.036461f
C1636 PAD.n527 VSS 0.036461f
C1637 PAD.n529 VSS 0.036461f
C1638 PAD.n530 VSS 0.036461f
C1639 PAD.n531 VSS 0.036461f
C1640 PAD.n532 VSS 0.036461f
C1641 PAD.n533 VSS 0.036461f
C1642 PAD.n534 VSS 0.036461f
C1643 PAD.n535 VSS 0.036461f
C1644 PAD.n537 VSS 0.036461f
C1645 PAD.n539 VSS 0.036461f
C1646 PAD.n541 VSS 0.036461f
C1647 PAD.n542 VSS 0.036461f
C1648 PAD.n543 VSS 0.036461f
C1649 PAD.n544 VSS 0.036461f
C1650 PAD.n545 VSS 0.036461f
C1651 PAD.n546 VSS 0.036461f
C1652 PAD.n547 VSS 0.036461f
C1653 PAD.n549 VSS 0.036461f
C1654 PAD.n551 VSS 0.036461f
C1655 PAD.n553 VSS 0.036461f
C1656 PAD.n554 VSS 0.036461f
C1657 PAD.n555 VSS 0.036461f
C1658 PAD.n556 VSS 0.036461f
C1659 PAD.n557 VSS 0.036461f
C1660 PAD.n558 VSS 0.036461f
C1661 PAD.n559 VSS 0.036461f
C1662 PAD.n561 VSS 0.036461f
C1663 PAD.n563 VSS 0.036461f
C1664 PAD.n565 VSS 0.036461f
C1665 PAD.n566 VSS 0.036461f
C1666 PAD.n567 VSS 0.036461f
C1667 PAD.n568 VSS 0.036461f
C1668 PAD.n569 VSS 0.036461f
C1669 PAD.n570 VSS 0.036461f
C1670 PAD.n571 VSS 0.036461f
C1671 PAD.n573 VSS 0.036461f
C1672 PAD.n575 VSS 0.036461f
C1673 PAD.n577 VSS 0.036461f
C1674 PAD.n578 VSS 0.036461f
C1675 PAD.n579 VSS 0.036461f
C1676 PAD.n580 VSS 0.036461f
C1677 PAD.n581 VSS 0.036461f
C1678 PAD.n582 VSS 0.036461f
C1679 PAD.n583 VSS 0.036461f
C1680 PAD.n585 VSS 0.036461f
C1681 PAD.n587 VSS 0.036461f
C1682 PAD.n589 VSS 0.036461f
C1683 PAD.n590 VSS 0.036461f
C1684 PAD.n591 VSS 0.036461f
C1685 PAD.n592 VSS 0.036461f
C1686 PAD.n593 VSS 0.036461f
C1687 PAD.n594 VSS 0.036461f
C1688 PAD.n595 VSS 0.036461f
C1689 PAD.n597 VSS 0.036461f
C1690 PAD.n599 VSS 0.036461f
C1691 PAD.n601 VSS 0.036461f
C1692 PAD.n602 VSS 0.036461f
C1693 PAD.n603 VSS 0.036461f
C1694 PAD.n604 VSS 0.036461f
C1695 PAD.n605 VSS 0.036461f
C1696 PAD.n606 VSS 0.036461f
C1697 PAD.n607 VSS 0.036461f
C1698 PAD.n609 VSS 0.036461f
C1699 PAD.n611 VSS 0.036461f
C1700 PAD.n613 VSS 0.036461f
C1701 PAD.n614 VSS 0.036461f
C1702 PAD.n615 VSS 0.036461f
C1703 PAD.n616 VSS 0.036461f
C1704 PAD.n617 VSS 0.036461f
C1705 PAD.n618 VSS 0.036461f
C1706 PAD.n619 VSS 0.036461f
C1707 PAD.n621 VSS 0.036461f
C1708 PAD.n623 VSS 0.036461f
C1709 PAD.n625 VSS 0.036461f
C1710 PAD.n626 VSS 0.036461f
C1711 PAD.n627 VSS 0.036461f
C1712 PAD.n628 VSS 0.036461f
C1713 PAD.n629 VSS 0.036461f
C1714 PAD.n630 VSS 0.036461f
C1715 PAD.n631 VSS 0.036461f
C1716 PAD.n633 VSS 0.036461f
C1717 PAD.n635 VSS 0.036461f
C1718 PAD.n637 VSS 0.036461f
C1719 PAD.n638 VSS 0.036461f
C1720 PAD.n639 VSS 0.036461f
C1721 PAD.n640 VSS 0.036461f
C1722 PAD.n641 VSS 0.036461f
C1723 PAD.n642 VSS 0.036461f
C1724 PAD.n643 VSS 0.036461f
C1725 PAD.n645 VSS 0.036461f
C1726 PAD.n647 VSS 0.036461f
C1727 PAD.n649 VSS 0.036461f
C1728 PAD.n650 VSS 0.036461f
C1729 PAD.n651 VSS 0.036461f
C1730 PAD.n652 VSS 0.036461f
C1731 PAD.n653 VSS 0.036461f
C1732 PAD.n654 VSS 0.036461f
C1733 PAD.n655 VSS 0.036461f
C1734 PAD.n657 VSS 0.036461f
C1735 PAD.n659 VSS 0.036461f
C1736 PAD.n661 VSS 0.036461f
C1737 PAD.n662 VSS 0.036461f
C1738 PAD.n663 VSS 0.036461f
C1739 PAD.n664 VSS 0.036461f
C1740 PAD.n665 VSS 0.036461f
C1741 PAD.n666 VSS 0.036461f
C1742 PAD.n667 VSS 0.036461f
C1743 PAD.n669 VSS 0.036461f
C1744 PAD.n671 VSS 0.036461f
C1745 PAD.n673 VSS 0.036461f
C1746 PAD.n674 VSS 0.036461f
C1747 PAD.n675 VSS 0.036461f
C1748 PAD.n676 VSS 0.036461f
C1749 PAD.n677 VSS 0.036461f
C1750 PAD.n678 VSS 0.036461f
C1751 PAD.n679 VSS 0.036461f
C1752 PAD.n681 VSS 0.036461f
C1753 PAD.n683 VSS 0.036461f
C1754 PAD.n685 VSS 0.036461f
C1755 PAD.n686 VSS 0.036461f
C1756 PAD.n687 VSS 0.036461f
C1757 PAD.n688 VSS 0.036461f
C1758 PAD.n689 VSS 0.036461f
C1759 PAD.n690 VSS 0.036461f
C1760 PAD.n691 VSS 0.036461f
C1761 PAD.n693 VSS 0.036461f
C1762 PAD.n695 VSS 0.036461f
C1763 PAD.n697 VSS 0.036461f
C1764 PAD.n698 VSS 0.036461f
C1765 PAD.n699 VSS 0.036461f
C1766 PAD.n700 VSS 0.036461f
C1767 PAD.n701 VSS 0.036461f
C1768 PAD.n702 VSS 0.036461f
C1769 PAD.n703 VSS 0.036461f
C1770 PAD.n705 VSS 0.036461f
C1771 PAD.n707 VSS 0.036461f
C1772 PAD.n709 VSS 0.036461f
C1773 PAD.n710 VSS 0.036461f
C1774 PAD.n711 VSS 0.036461f
C1775 PAD.n712 VSS 0.036461f
C1776 PAD.n713 VSS 0.036461f
C1777 PAD.n714 VSS 0.036461f
C1778 PAD.n715 VSS 0.036461f
C1779 PAD.n717 VSS 0.036461f
C1780 PAD.n719 VSS 0.036461f
C1781 PAD.n721 VSS 0.036461f
C1782 PAD.n722 VSS 0.036461f
C1783 PAD.n723 VSS 0.036461f
C1784 PAD.n724 VSS 0.036461f
C1785 PAD.n725 VSS 0.036461f
C1786 PAD.n726 VSS 0.036461f
C1787 PAD.n727 VSS 0.036461f
C1788 PAD.n729 VSS 0.036461f
C1789 PAD.n731 VSS 0.036461f
C1790 PAD.n733 VSS 0.036461f
C1791 PAD.n734 VSS 0.036461f
C1792 PAD.n735 VSS 0.036461f
C1793 PAD.n736 VSS 0.036461f
C1794 PAD.n737 VSS 0.036461f
C1795 PAD.n738 VSS 0.036461f
C1796 PAD.n739 VSS 0.036461f
C1797 PAD.n741 VSS 0.036461f
C1798 PAD.n743 VSS 0.036461f
C1799 PAD.n745 VSS 0.036461f
C1800 PAD.n746 VSS 0.036461f
C1801 PAD.n747 VSS 0.036461f
C1802 PAD.n748 VSS 0.036461f
C1803 PAD.n749 VSS 0.036461f
C1804 PAD.n750 VSS 0.036461f
C1805 PAD.n751 VSS 0.036461f
C1806 PAD.n753 VSS 0.036461f
C1807 PAD.n755 VSS 0.036461f
C1808 PAD.n757 VSS 0.036461f
C1809 PAD.n758 VSS 0.036461f
C1810 PAD.n759 VSS 0.036461f
C1811 PAD.n760 VSS 0.036461f
C1812 PAD.n761 VSS 0.036461f
C1813 PAD.n762 VSS 0.036461f
C1814 PAD.n763 VSS 0.036461f
C1815 PAD.n764 VSS 0.036461f
C1816 PAD.n766 VSS 0.036461f
C1817 PAD.n768 VSS 0.036461f
C1818 PAD.n770 VSS 0.023109f
C1819 PAD.n771 VSS 0.023109f
C1820 PAD.n772 VSS 0.030555f
C1821 PAD.n773 VSS 0.042895f
C1822 PAD.n774 VSS 0.049115f
C1823 PAD.n775 VSS 0.049115f
C1824 PAD.n776 VSS 0.700534f
C1825 PAD.n777 VSS 0.069765f
C1826 PAD.n778 VSS 0.069765f
C1827 PAD.n779 VSS 0.046286f
C1828 PAD.n780 VSS 0.039761f
C1829 PAD.n781 VSS 0.039761f
C1830 PAD.n782 VSS 0.611734f
C1831 PAD.n824 VSS 0.023109f
C1832 PAD.n825 VSS 0.542667f
C1833 PAD.n826 VSS 0.023109f
C1834 PAD.n827 VSS 0.029436f
C1835 PAD.n828 VSS 0.350267f
C1836 PAD.n829 VSS 0.036461f
C1837 PAD.n830 VSS 0.036461f
C1838 PAD.n831 VSS 0.036461f
C1839 PAD.n832 VSS 0.036461f
C1840 PAD.n833 VSS 0.036461f
C1841 PAD.n834 VSS 0.036461f
C1842 PAD.n835 VSS 0.036461f
C1843 PAD.n836 VSS 0.036461f
C1844 PAD.n837 VSS 0.036461f
C1845 PAD.n838 VSS 0.036461f
C1846 PAD.n839 VSS 0.036461f
C1847 PAD.n840 VSS 0.036461f
C1848 PAD.n841 VSS 0.036461f
C1849 PAD.n842 VSS 0.036461f
C1850 PAD.n843 VSS 0.036461f
C1851 PAD.n844 VSS 0.036461f
C1852 PAD.n845 VSS 0.036461f
C1853 PAD.n846 VSS 0.036461f
C1854 PAD.n847 VSS 0.036461f
C1855 PAD.n848 VSS 0.036461f
C1856 PAD.n849 VSS 0.036461f
C1857 PAD.n850 VSS 0.036461f
C1858 PAD.n851 VSS 0.036461f
C1859 PAD.n852 VSS 0.036461f
C1860 PAD.n853 VSS 0.036461f
C1861 PAD.n854 VSS 0.036461f
C1862 PAD.n855 VSS 0.036461f
C1863 PAD.n856 VSS 0.036461f
C1864 PAD.n857 VSS 0.036461f
C1865 PAD.n858 VSS 0.036461f
C1866 PAD.n859 VSS 0.036461f
C1867 PAD.n860 VSS 0.036461f
C1868 PAD.n861 VSS 0.036461f
C1869 PAD.n862 VSS 0.036461f
C1870 PAD.n863 VSS 0.036461f
C1871 PAD.n864 VSS 0.036461f
C1872 PAD.n865 VSS 0.036461f
C1873 PAD.n866 VSS 0.036461f
C1874 PAD.n867 VSS 0.036461f
C1875 PAD.n868 VSS 0.036461f
C1876 PAD.n870 VSS 0.036461f
C1877 PAD.n871 VSS 0.036461f
C1878 PAD.n872 VSS 0.023109f
C1879 PAD.n873 VSS 0.03338f
C1880 PAD.n874 VSS 0.036461f
C1881 PAD.n875 VSS 0.036461f
C1882 PAD.n876 VSS 0.036461f
C1883 PAD.n877 VSS 0.036461f
C1884 PAD.n879 VSS 0.036461f
C1885 PAD.n880 VSS 0.036461f
C1886 PAD.n881 VSS 0.036461f
C1887 PAD.n883 VSS 0.036461f
C1888 PAD.n884 VSS 0.036461f
C1889 PAD.n885 VSS 0.036461f
C1890 PAD.n886 VSS 0.036461f
C1891 PAD.n887 VSS 0.036461f
C1892 PAD.n888 VSS 0.036461f
C1893 PAD.n889 VSS 0.036461f
C1894 PAD.n891 VSS 0.036461f
C1895 PAD.n892 VSS 0.036461f
C1896 PAD.n893 VSS 0.036461f
C1897 PAD.n895 VSS 0.036461f
C1898 PAD.n896 VSS 0.036461f
C1899 PAD.n897 VSS 0.036461f
C1900 PAD.n898 VSS 0.036461f
C1901 PAD.n899 VSS 0.036461f
C1902 PAD.n900 VSS 0.036461f
C1903 PAD.n901 VSS 0.036461f
C1904 PAD.n903 VSS 0.036461f
C1905 PAD.n904 VSS 0.036461f
C1906 PAD.n905 VSS 0.036461f
C1907 PAD.n907 VSS 0.036461f
C1908 PAD.n908 VSS 0.036461f
C1909 PAD.n909 VSS 0.036461f
C1910 PAD.n910 VSS 0.036461f
C1911 PAD.n911 VSS 0.036461f
C1912 PAD.n912 VSS 0.036461f
C1913 PAD.n913 VSS 0.036461f
C1914 PAD.n915 VSS 0.036461f
C1915 PAD.n916 VSS 0.036461f
C1916 PAD.n917 VSS 0.036461f
C1917 PAD.n919 VSS 0.036461f
C1918 PAD.n920 VSS 0.036461f
C1919 PAD.n921 VSS 0.036461f
C1920 PAD.n922 VSS 0.036461f
C1921 PAD.n923 VSS 0.036461f
C1922 PAD.n924 VSS 0.036461f
C1923 PAD.n925 VSS 0.036461f
C1924 PAD.n927 VSS 0.036461f
C1925 PAD.n928 VSS 0.036461f
C1926 PAD.n929 VSS 0.036461f
C1927 PAD.n931 VSS 0.036461f
C1928 PAD.n932 VSS 0.036461f
C1929 PAD.n933 VSS 0.036461f
C1930 PAD.n934 VSS 0.036461f
C1931 PAD.n935 VSS 0.036461f
C1932 PAD.n936 VSS 0.036461f
C1933 PAD.n937 VSS 0.036461f
C1934 PAD.n939 VSS 0.036461f
C1935 PAD.n940 VSS 0.036461f
C1936 PAD.n941 VSS 0.036461f
C1937 PAD.n943 VSS 0.036461f
C1938 PAD.n944 VSS 0.036461f
C1939 PAD.n945 VSS 0.036461f
C1940 PAD.n946 VSS 0.036461f
C1941 PAD.n947 VSS 0.036461f
C1942 PAD.n948 VSS 0.036461f
C1943 PAD.n949 VSS 0.036461f
C1944 PAD.n951 VSS 0.036461f
C1945 PAD.n952 VSS 0.036461f
C1946 PAD.n953 VSS 0.036461f
C1947 PAD.n955 VSS 0.036461f
C1948 PAD.n956 VSS 0.036461f
C1949 PAD.n957 VSS 0.036461f
C1950 PAD.n958 VSS 0.036461f
C1951 PAD.n959 VSS 0.036461f
C1952 PAD.n960 VSS 0.036461f
C1953 PAD.n961 VSS 0.036461f
C1954 PAD.n963 VSS 0.036461f
C1955 PAD.n964 VSS 0.036461f
C1956 PAD.n965 VSS 0.036461f
C1957 PAD.n967 VSS 0.036461f
C1958 PAD.n968 VSS 0.036461f
C1959 PAD.n969 VSS 0.036461f
C1960 PAD.n970 VSS 0.036461f
C1961 PAD.n971 VSS 0.036461f
C1962 PAD.n972 VSS 0.036461f
C1963 PAD.n973 VSS 0.036461f
C1964 PAD.n975 VSS 0.036461f
C1965 PAD.n976 VSS 0.036461f
C1966 PAD.n977 VSS 0.036461f
C1967 PAD.n979 VSS 0.036461f
C1968 PAD.n980 VSS 0.036461f
C1969 PAD.n981 VSS 0.036461f
C1970 PAD.n982 VSS 0.036461f
C1971 PAD.n983 VSS 0.036461f
C1972 PAD.n984 VSS 0.036461f
C1973 PAD.n985 VSS 0.036461f
C1974 PAD.n987 VSS 0.036461f
C1975 PAD.n988 VSS 0.036461f
C1976 PAD.n989 VSS 0.036461f
C1977 PAD.n991 VSS 0.036461f
C1978 PAD.n992 VSS 0.036461f
C1979 PAD.n993 VSS 0.036461f
C1980 PAD.n994 VSS 0.036461f
C1981 PAD.n995 VSS 0.036461f
C1982 PAD.n996 VSS 0.036461f
C1983 PAD.n997 VSS 0.036461f
C1984 PAD.n999 VSS 0.036461f
C1985 PAD.n1000 VSS 0.036461f
C1986 PAD.n1001 VSS 0.036461f
C1987 PAD.n1003 VSS 0.036461f
C1988 PAD.n1004 VSS 0.036461f
C1989 PAD.n1005 VSS 0.036461f
C1990 PAD.n1006 VSS 0.036461f
C1991 PAD.n1007 VSS 0.036461f
C1992 PAD.n1008 VSS 0.036461f
C1993 PAD.n1009 VSS 0.036461f
C1994 PAD.n1011 VSS 0.036461f
C1995 PAD.n1012 VSS 0.036461f
C1996 PAD.n1013 VSS 0.036461f
C1997 PAD.n1015 VSS 0.036461f
C1998 PAD.n1016 VSS 0.036461f
C1999 PAD.n1017 VSS 0.036461f
C2000 PAD.n1018 VSS 0.036461f
C2001 PAD.n1019 VSS 0.036461f
C2002 PAD.n1020 VSS 0.036461f
C2003 PAD.n1021 VSS 0.036461f
C2004 PAD.n1023 VSS 0.036461f
C2005 PAD.n1024 VSS 0.036461f
C2006 PAD.n1025 VSS 0.036461f
C2007 PAD.n1027 VSS 0.036461f
C2008 PAD.n1028 VSS 0.036461f
C2009 PAD.n1029 VSS 0.036461f
C2010 PAD.n1030 VSS 0.036461f
C2011 PAD.n1031 VSS 0.036461f
C2012 PAD.n1032 VSS 0.036461f
C2013 PAD.n1033 VSS 0.036461f
C2014 PAD.n1035 VSS 0.036461f
C2015 PAD.n1036 VSS 0.036461f
C2016 PAD.n1037 VSS 0.036461f
C2017 PAD.n1039 VSS 0.036461f
C2018 PAD.n1040 VSS 0.036461f
C2019 PAD.n1041 VSS 0.036461f
C2020 PAD.n1042 VSS 0.036461f
C2021 PAD.n1043 VSS 0.036461f
C2022 PAD.n1044 VSS 0.036461f
C2023 PAD.n1045 VSS 0.036461f
C2024 PAD.n1047 VSS 0.036461f
C2025 PAD.n1048 VSS 0.036461f
C2026 PAD.n1049 VSS 0.036461f
C2027 PAD.n1051 VSS 0.036461f
C2028 PAD.n1052 VSS 0.036461f
C2029 PAD.n1053 VSS 0.036461f
C2030 PAD.n1054 VSS 0.036461f
C2031 PAD.n1055 VSS 0.036461f
C2032 PAD.n1056 VSS 0.036461f
C2033 PAD.n1057 VSS 0.036461f
C2034 PAD.n1059 VSS 0.036461f
C2035 PAD.n1060 VSS 0.036461f
C2036 PAD.n1061 VSS 0.036461f
C2037 PAD.n1063 VSS 0.036461f
C2038 PAD.n1064 VSS 0.036461f
C2039 PAD.n1065 VSS 0.036461f
C2040 PAD.n1066 VSS 0.036461f
C2041 PAD.n1067 VSS 0.036461f
C2042 PAD.n1068 VSS 0.036461f
C2043 PAD.n1069 VSS 0.036461f
C2044 PAD.n1071 VSS 0.036461f
C2045 PAD.n1072 VSS 0.036461f
C2046 PAD.n1073 VSS 0.036461f
C2047 PAD.n1075 VSS 0.036461f
C2048 PAD.n1076 VSS 0.036461f
C2049 PAD.n1077 VSS 0.036461f
C2050 PAD.n1078 VSS 0.036461f
C2051 PAD.n1079 VSS 0.036461f
C2052 PAD.n1080 VSS 0.036461f
C2053 PAD.n1081 VSS 0.036461f
C2054 PAD.n1083 VSS 0.036461f
C2055 PAD.n1084 VSS 0.036461f
C2056 PAD.n1085 VSS 0.036461f
C2057 PAD.n1087 VSS 0.036461f
C2058 PAD.n1088 VSS 0.036461f
C2059 PAD.n1089 VSS 0.036461f
C2060 PAD.n1090 VSS 0.036461f
C2061 PAD.n1091 VSS 0.036461f
C2062 PAD.n1092 VSS 0.036461f
C2063 PAD.n1093 VSS 0.036461f
C2064 PAD.n1095 VSS 0.036461f
C2065 PAD.n1096 VSS 0.036461f
C2066 PAD.n1097 VSS 0.036461f
C2067 PAD.n1099 VSS 0.036461f
C2068 PAD.n1100 VSS 0.036461f
C2069 PAD.n1101 VSS 0.036461f
C2070 PAD.n1102 VSS 0.036461f
C2071 PAD.n1103 VSS 0.036461f
C2072 PAD.n1104 VSS 0.036461f
C2073 PAD.n1105 VSS 0.036461f
C2074 PAD.n1107 VSS 0.036461f
C2075 PAD.n1108 VSS 0.036461f
C2076 PAD.n1109 VSS 0.036461f
C2077 PAD.n1111 VSS 0.036461f
C2078 PAD.n1112 VSS 0.036461f
C2079 PAD.n1113 VSS 0.036461f
C2080 PAD.n1114 VSS 0.036461f
C2081 PAD.n1115 VSS 0.041838f
C2082 PAD.n1116 VSS 0.045829f
C2083 PAD.n1117 VSS 0.045829f
C2084 PAD.n1118 VSS 0.611734f
C2085 PAD.n1119 VSS 0.059638f
C2086 PAD.n1120 VSS 0.37f
C2087 PAD.n1121 VSS 0.052887f
C2088 PAD.n1122 VSS 0.059638f
C2089 PAD.n1123 VSS 0.052887f
C2090 PAD.n1124 VSS 0.03338f
C2091 PAD.n1125 VSS 0.062274f
C2092 PAD.n1126 VSS 0.069765f
C2093 PAD.n1127 VSS 0.039761f
C2094 PAD.n1128 VSS 0.069765f
C2095 PAD.n1129 VSS 0.039761f
C2096 PAD.n1130 VSS 0.611735f
C2097 PAD.n1131 VSS 0.261467f
C2098 PAD.n1132 VSS 0.527867f
C2099 PAD.n1133 VSS 0.049115f
C2100 PAD.n1134 VSS 0.029436f
C2101 PAD.n1135 VSS 0.049115f
C2102 PAD.n1136 VSS 0.029436f
C2103 PAD.n1137 VSS 0.033773f
C2104 PAD.n1138 VSS 0.029436f
C2105 PAD.n1139 VSS 0.029436f
C2106 PAD.n1140 VSS 0.518001f
C2107 PAD.n1141 VSS 0.439067f
C2108 PAD.n1142 VSS 0.611734f
C2109 PAD.n1143 VSS 0.039761f
C2110 PAD.n1144 VSS 0.039761f
C2111 PAD.n1145 VSS 0.03338f
C2112 PAD.n1146 VSS 0.062274f
C2113 PAD.n1147 VSS 0.069765f
C2114 PAD.n1148 VSS 0.069765f
C2115 PAD.n1190 VSS 0.036461f
C2116 PAD.n1192 VSS 0.036461f
C2117 PAD.n1193 VSS 0.036461f
C2118 PAD.n1194 VSS 0.036461f
C2119 PAD.n1195 VSS 0.036461f
C2120 PAD.n1196 VSS 0.036461f
C2121 PAD.n1198 VSS 0.036461f
C2122 PAD.n1199 VSS 0.036461f
C2123 PAD.n1200 VSS 0.036461f
C2124 PAD.n1201 VSS 0.036461f
C2125 PAD.n1203 VSS 0.036461f
C2126 PAD.n1204 VSS 0.036461f
C2127 PAD.n1205 VSS 0.036461f
C2128 PAD.n1206 VSS 0.036461f
C2129 PAD.n1208 VSS 0.036461f
C2130 PAD.n1209 VSS 0.036461f
C2131 PAD.n1210 VSS 0.036461f
C2132 PAD.n1211 VSS 0.036461f
C2133 PAD.n1213 VSS 0.036461f
C2134 PAD.n1214 VSS 0.036461f
C2135 PAD.n1215 VSS 0.036461f
C2136 PAD.n1216 VSS 0.036461f
C2137 PAD.n1218 VSS 0.036461f
C2138 PAD.n1219 VSS 0.036461f
C2139 PAD.n1220 VSS 0.036461f
C2140 PAD.n1221 VSS 0.036461f
C2141 PAD.n1223 VSS 0.036461f
C2142 PAD.n1224 VSS 0.036461f
C2143 PAD.n1225 VSS 0.036461f
C2144 PAD.n1226 VSS 0.036461f
C2145 PAD.n1228 VSS 0.036461f
C2146 PAD.n1229 VSS 0.036461f
C2147 PAD.n1230 VSS 0.036461f
C2148 PAD.n1231 VSS 0.036461f
C2149 PAD.n1233 VSS 0.036461f
C2150 PAD.n1234 VSS 0.036461f
C2151 PAD.n1235 VSS 0.036461f
C2152 PAD.n1236 VSS 0.036461f
C2153 PAD.n1238 VSS 0.036461f
C2154 PAD.n1239 VSS 0.036461f
C2155 PAD.n1240 VSS 0.036461f
C2156 PAD.n1241 VSS 0.036461f
C2157 PAD.n1243 VSS 0.036461f
C2158 PAD.n1244 VSS 0.036461f
C2159 PAD.n1245 VSS 0.036461f
C2160 PAD.n1246 VSS 0.036461f
C2161 PAD.n1248 VSS 0.036461f
C2162 PAD.n1249 VSS 0.036461f
C2163 PAD.n1250 VSS 0.036461f
C2164 PAD.n1251 VSS 0.036461f
C2165 PAD.n1253 VSS 0.036461f
C2166 PAD.n1254 VSS 0.036461f
C2167 PAD.n1255 VSS 0.036461f
C2168 PAD.n1256 VSS 0.036461f
C2169 PAD.n1258 VSS 0.036461f
C2170 PAD.n1259 VSS 0.036461f
C2171 PAD.n1260 VSS 0.036461f
C2172 PAD.n1261 VSS 0.036461f
C2173 PAD.n1263 VSS 0.036461f
C2174 PAD.n1264 VSS 0.036461f
C2175 PAD.n1265 VSS 0.036461f
C2176 PAD.n1266 VSS 0.036461f
C2177 PAD.n1268 VSS 0.036461f
C2178 PAD.n1269 VSS 0.036461f
C2179 PAD.n1270 VSS 0.036461f
C2180 PAD.n1271 VSS 0.036461f
C2181 PAD.n1273 VSS 0.036461f
C2182 PAD.n1274 VSS 0.036461f
C2183 PAD.n1275 VSS 0.036461f
C2184 PAD.n1276 VSS 0.036461f
C2185 PAD.n1278 VSS 0.036461f
C2186 PAD.n1279 VSS 0.036461f
C2187 PAD.n1280 VSS 0.036461f
C2188 PAD.n1281 VSS 0.036461f
C2189 PAD.n1283 VSS 0.036461f
C2190 PAD.n1284 VSS 0.036461f
C2191 PAD.n1285 VSS 0.036461f
C2192 PAD.n1286 VSS 0.036461f
C2193 PAD.n1288 VSS 0.036461f
C2194 PAD.n1289 VSS 0.036461f
C2195 PAD.n1290 VSS 0.036461f
C2196 PAD.n1291 VSS 0.036461f
C2197 PAD.n1293 VSS 0.036461f
C2198 PAD.n1294 VSS 0.023109f
C2199 PAD.n1295 VSS 0.023109f
C2200 PAD.n1296 VSS 0.030555f
C2201 PAD.n1297 VSS 0.036461f
C2202 PAD.n1298 VSS 0.036461f
C2203 PAD.n1299 VSS 0.036461f
C2204 PAD.n1300 VSS 0.036461f
C2205 PAD.n1301 VSS 0.036461f
C2206 PAD.n1303 VSS 0.036461f
C2207 PAD.n1304 VSS 0.036461f
C2208 PAD.n1305 VSS 0.036461f
C2209 PAD.n1306 VSS 0.036461f
C2210 PAD.n1307 VSS 0.036461f
C2211 PAD.n1308 VSS 0.036461f
C2212 PAD.n1309 VSS 0.036461f
C2213 PAD.n1310 VSS 0.036461f
C2214 PAD.n1312 VSS 0.036461f
C2215 PAD.n1313 VSS 0.036461f
C2216 PAD.n1314 VSS 0.036461f
C2217 PAD.n1315 VSS 0.036461f
C2218 PAD.n1316 VSS 0.036461f
C2219 PAD.n1317 VSS 0.036461f
C2220 PAD.n1318 VSS 0.036461f
C2221 PAD.n1319 VSS 0.036461f
C2222 PAD.n1321 VSS 0.036461f
C2223 PAD.n1322 VSS 0.036461f
C2224 PAD.n1323 VSS 0.036461f
C2225 PAD.n1324 VSS 0.036461f
C2226 PAD.n1325 VSS 0.036461f
C2227 PAD.n1326 VSS 0.036461f
C2228 PAD.n1327 VSS 0.036461f
C2229 PAD.n1328 VSS 0.036461f
C2230 PAD.n1330 VSS 0.036461f
C2231 PAD.n1331 VSS 0.036461f
C2232 PAD.n1332 VSS 0.036461f
C2233 PAD.n1333 VSS 0.036461f
C2234 PAD.n1334 VSS 0.036461f
C2235 PAD.n1335 VSS 0.036461f
C2236 PAD.n1336 VSS 0.036461f
C2237 PAD.n1337 VSS 0.036461f
C2238 PAD.n1339 VSS 0.036461f
C2239 PAD.n1340 VSS 0.036461f
C2240 PAD.n1341 VSS 0.036461f
C2241 PAD.n1342 VSS 0.036461f
C2242 PAD.n1343 VSS 0.036461f
C2243 PAD.n1344 VSS 0.036461f
C2244 PAD.n1345 VSS 0.036461f
C2245 PAD.n1346 VSS 0.036461f
C2246 PAD.n1348 VSS 0.036461f
C2247 PAD.n1349 VSS 0.036461f
C2248 PAD.n1350 VSS 0.036461f
C2249 PAD.n1351 VSS 0.036461f
C2250 PAD.n1352 VSS 0.036461f
C2251 PAD.n1353 VSS 0.036461f
C2252 PAD.n1354 VSS 0.036461f
C2253 PAD.n1355 VSS 0.036461f
C2254 PAD.n1357 VSS 0.036461f
C2255 PAD.n1358 VSS 0.036461f
C2256 PAD.n1359 VSS 0.036461f
C2257 PAD.n1360 VSS 0.036461f
C2258 PAD.n1361 VSS 0.036461f
C2259 PAD.n1362 VSS 0.036461f
C2260 PAD.n1363 VSS 0.036461f
C2261 PAD.n1364 VSS 0.036461f
C2262 PAD.n1366 VSS 0.036461f
C2263 PAD.n1367 VSS 0.036461f
C2264 PAD.n1368 VSS 0.036461f
C2265 PAD.n1369 VSS 0.036461f
C2266 PAD.n1370 VSS 0.036461f
C2267 PAD.n1371 VSS 0.036461f
C2268 PAD.n1372 VSS 0.036461f
C2269 PAD.n1373 VSS 0.036461f
C2270 PAD.n1375 VSS 0.036461f
C2271 PAD.n1376 VSS 0.036461f
C2272 PAD.n1377 VSS 0.036461f
C2273 PAD.n1378 VSS 0.036461f
C2274 PAD.n1379 VSS 0.036461f
C2275 PAD.n1380 VSS 0.036461f
C2276 PAD.n1381 VSS 0.036461f
C2277 PAD.n1382 VSS 0.036461f
C2278 PAD.n1384 VSS 0.036461f
C2279 PAD.n1385 VSS 0.036461f
C2280 PAD.n1386 VSS 0.036461f
C2281 PAD.n1387 VSS 0.036461f
C2282 PAD.n1388 VSS 0.036461f
C2283 PAD.n1389 VSS 0.036461f
C2284 PAD.n1390 VSS 0.036461f
C2285 PAD.n1391 VSS 0.036461f
C2286 PAD.n1393 VSS 0.036461f
C2287 PAD.n1394 VSS 0.036461f
C2288 PAD.n1395 VSS 0.036461f
C2289 PAD.n1396 VSS 0.036461f
C2290 PAD.n1397 VSS 0.036461f
C2291 PAD.n1398 VSS 0.036461f
C2292 PAD.n1399 VSS 0.036461f
C2293 PAD.n1400 VSS 0.036461f
C2294 PAD.n1402 VSS 0.036461f
C2295 PAD.n1403 VSS 0.036461f
C2296 PAD.n1404 VSS 0.036461f
C2297 PAD.n1405 VSS 0.036461f
C2298 PAD.n1406 VSS 0.036461f
C2299 PAD.n1407 VSS 0.036461f
C2300 PAD.n1408 VSS 0.036461f
C2301 PAD.n1409 VSS 0.036461f
C2302 PAD.n1411 VSS 0.036461f
C2303 PAD.n1412 VSS 0.036461f
C2304 PAD.n1413 VSS 0.036461f
C2305 PAD.n1414 VSS 0.036461f
C2306 PAD.n1415 VSS 0.036461f
C2307 PAD.n1416 VSS 0.036461f
C2308 PAD.n1417 VSS 0.036461f
C2309 PAD.n1418 VSS 0.036461f
C2310 PAD.n1420 VSS 0.036461f
C2311 PAD.n1421 VSS 0.036461f
C2312 PAD.n1422 VSS 0.036461f
C2313 PAD.n1423 VSS 0.036461f
C2314 PAD.n1424 VSS 0.036461f
C2315 PAD.n1425 VSS 0.036461f
C2316 PAD.n1426 VSS 0.036461f
C2317 PAD.n1427 VSS 0.036461f
C2318 PAD.n1429 VSS 0.036461f
C2319 PAD.n1430 VSS 0.036461f
C2320 PAD.n1431 VSS 0.036461f
C2321 PAD.n1432 VSS 0.036461f
C2322 PAD.n1433 VSS 0.036461f
C2323 PAD.n1434 VSS 0.036461f
C2324 PAD.n1435 VSS 0.036461f
C2325 PAD.n1436 VSS 0.036461f
C2326 PAD.n1438 VSS 0.036461f
C2327 PAD.n1439 VSS 0.036461f
C2328 PAD.n1440 VSS 0.036461f
C2329 PAD.n1441 VSS 0.036461f
C2330 PAD.n1442 VSS 0.036461f
C2331 PAD.n1443 VSS 0.036461f
C2332 PAD.n1444 VSS 0.036461f
C2333 PAD.n1445 VSS 0.036461f
C2334 PAD.n1447 VSS 0.036461f
C2335 PAD.n1448 VSS 0.036461f
C2336 PAD.n1449 VSS 0.036461f
C2337 PAD.n1450 VSS 0.036461f
C2338 PAD.n1451 VSS 0.036461f
C2339 PAD.n1452 VSS 0.036461f
C2340 PAD.n1453 VSS 0.036461f
C2341 PAD.n1454 VSS 0.036461f
C2342 PAD.n1456 VSS 0.036461f
C2343 PAD.n1457 VSS 0.036461f
C2344 PAD.n1458 VSS 0.036461f
C2345 PAD.n1459 VSS 0.036461f
C2346 PAD.n1460 VSS 0.036461f
C2347 PAD.n1461 VSS 0.036461f
C2348 PAD.n1462 VSS 0.036461f
C2349 PAD.n1463 VSS 0.036461f
C2350 PAD.n1465 VSS 0.036461f
C2351 PAD.n1466 VSS 0.036461f
C2352 PAD.n1467 VSS 0.036461f
C2353 PAD.n1468 VSS 0.036461f
C2354 PAD.n1469 VSS 0.036461f
C2355 PAD.n1470 VSS 0.036461f
C2356 PAD.n1471 VSS 0.036461f
C2357 PAD.n1472 VSS 0.036461f
C2358 PAD.n1474 VSS 0.036461f
C2359 PAD.n1475 VSS 0.036461f
C2360 PAD.n1476 VSS 0.036461f
C2361 PAD.n1477 VSS 0.036461f
C2362 PAD.n1478 VSS 0.036461f
C2363 PAD.n1479 VSS 0.036461f
C2364 PAD.n1480 VSS 0.023109f
C2365 PAD.n1481 VSS 0.023109f
C2366 PAD.n1483 VSS 0.429201f
C2367 PAD.n1484 VSS 0.049115f
C2368 PAD.n1485 VSS 0.049115f
C2369 PAD.n1486 VSS 0.033773f
C2370 PAD.n1487 VSS 0.029436f
C2371 PAD.n1488 VSS 0.029436f
C2372 PAD.n1489 VSS 0.685734f
C2373 PAD.n1531 VSS 0.023109f
C2374 PAD.n1532 VSS 0.587068f
C2375 PAD.n1533 VSS 0.611734f
C2376 PAD.n1534 VSS 0.685734f
C2377 PAD.n1535 VSS 0.023109f
C2378 PAD.n1536 VSS 0.448934f
C2379 PAD.n1537 VSS 0.036461f
C2380 PAD.n1538 VSS 0.036461f
C2381 PAD.n1539 VSS 0.036461f
C2382 PAD.n1540 VSS 0.036461f
C2383 PAD.n1541 VSS 0.036461f
C2384 PAD.n1542 VSS 0.036461f
C2385 PAD.n1543 VSS 0.036461f
C2386 PAD.n1544 VSS 0.036461f
C2387 PAD.n1545 VSS 0.036461f
C2388 PAD.n1546 VSS 0.036461f
C2389 PAD.n1547 VSS 0.036461f
C2390 PAD.n1548 VSS 0.036461f
C2391 PAD.n1549 VSS 0.036461f
C2392 PAD.n1550 VSS 0.036461f
C2393 PAD.n1551 VSS 0.036461f
C2394 PAD.n1552 VSS 0.036461f
C2395 PAD.n1553 VSS 0.036461f
C2396 PAD.n1554 VSS 0.036461f
C2397 PAD.n1555 VSS 0.036461f
C2398 PAD.n1556 VSS 0.036461f
C2399 PAD.n1557 VSS 0.036461f
C2400 PAD.n1558 VSS 0.036461f
C2401 PAD.n1559 VSS 0.036461f
C2402 PAD.n1560 VSS 0.036461f
C2403 PAD.n1561 VSS 0.036461f
C2404 PAD.n1562 VSS 0.036461f
C2405 PAD.n1563 VSS 0.036461f
C2406 PAD.n1564 VSS 0.036461f
C2407 PAD.n1565 VSS 0.036461f
C2408 PAD.n1566 VSS 0.036461f
C2409 PAD.n1567 VSS 0.036461f
C2410 PAD.n1568 VSS 0.036461f
C2411 PAD.n1569 VSS 0.036461f
C2412 PAD.n1570 VSS 0.036461f
C2413 PAD.n1571 VSS 0.036461f
C2414 PAD.n1572 VSS 0.036461f
C2415 PAD.n1573 VSS 0.036461f
C2416 PAD.n1574 VSS 0.036461f
C2417 PAD.n1575 VSS 0.036461f
C2418 PAD.n1576 VSS 0.036461f
C2419 PAD.n1578 VSS 0.036461f
C2420 PAD.n1579 VSS 0.036461f
C2421 PAD.n1580 VSS 0.046286f
C2422 PAD.n1581 VSS 0.064139f
C2423 PAD.n1582 VSS 0.069765f
C2424 PAD.n1583 VSS 0.062274f
C2425 PAD.n1584 VSS 0.036159f
C2426 PAD.n1585 VSS 0.069765f
C2427 PAD.n1586 VSS 0.611734f
C2428 PAD.n1587 VSS 0.049115f
C2429 PAD.n1588 VSS 0.049115f
C2430 PAD.n1589 VSS 0.033773f
C2431 PAD.n1590 VSS 0.029436f
C2432 PAD.n1591 VSS 0.029436f
C2433 PAD.n1592 VSS 0.596934f
C2434 PAD.n1593 VSS 0.542667f
C2435 PAD.n1594 VSS 0.611734f
C2436 PAD.n1595 VSS 0.039761f
C2437 PAD.n1596 VSS 0.039761f
C2438 PAD.n1597 VSS 0.069765f
C2439 PAD.n1598 VSS 0.036461f
C2440 PAD.n1599 VSS 0.023109f
C2441 PAD.n1600 VSS 0.036461f
C2442 PAD.n1603 VSS 0.036461f
C2443 PAD.n1604 VSS 0.036461f
C2444 PAD.n1605 VSS 0.036461f
C2445 PAD.n1606 VSS 0.036461f
C2446 PAD.n1608 VSS 0.036461f
C2447 PAD.n1609 VSS 0.036461f
C2448 PAD.n1610 VSS 0.036461f
C2449 PAD.n1612 VSS 0.036461f
C2450 PAD.n1613 VSS 0.036461f
C2451 PAD.n1614 VSS 0.036461f
C2452 PAD.n1616 VSS 0.036461f
C2453 PAD.n1617 VSS 0.036461f
C2454 PAD.n1618 VSS 0.036461f
C2455 PAD.n1620 VSS 0.036461f
C2456 PAD.n1621 VSS 0.036461f
C2457 PAD.n1622 VSS 0.036461f
C2458 PAD.n1624 VSS 0.036461f
C2459 PAD.n1625 VSS 0.036461f
C2460 PAD.n1626 VSS 0.036461f
C2461 PAD.n1628 VSS 0.036461f
C2462 PAD.n1629 VSS 0.036461f
C2463 PAD.n1630 VSS 0.036461f
C2464 PAD.n1632 VSS 0.036461f
C2465 PAD.n1633 VSS 0.036461f
C2466 PAD.n1634 VSS 0.036461f
C2467 PAD.n1636 VSS 0.036461f
C2468 PAD.n1637 VSS 0.036461f
C2469 PAD.n1638 VSS 0.036461f
C2470 PAD.n1640 VSS 0.036461f
C2471 PAD.n1641 VSS 0.036461f
C2472 PAD.n1642 VSS 0.036461f
C2473 PAD.n1644 VSS 0.036461f
C2474 PAD.n1645 VSS 0.036461f
C2475 PAD.n1646 VSS 0.036461f
C2476 PAD.n1648 VSS 0.036461f
C2477 PAD.n1649 VSS 0.036461f
C2478 PAD.n1650 VSS 0.036461f
C2479 PAD.n1652 VSS 0.036461f
C2480 PAD.n1653 VSS 0.036461f
C2481 PAD.n1654 VSS 0.036461f
C2482 PAD.n1656 VSS 0.036461f
C2483 PAD.n1657 VSS 0.036461f
C2484 PAD.n1658 VSS 0.036461f
C2485 PAD.n1660 VSS 0.036461f
C2486 PAD.n1661 VSS 0.036461f
C2487 PAD.n1662 VSS 0.036461f
C2488 PAD.n1664 VSS 0.036461f
C2489 PAD.n1665 VSS 0.036461f
C2490 PAD.n1666 VSS 0.036461f
C2491 PAD.n1668 VSS 0.036461f
C2492 PAD.n1669 VSS 0.036461f
C2493 PAD.n1670 VSS 0.036461f
C2494 PAD.n1672 VSS 0.036461f
C2495 PAD.n1673 VSS 0.036461f
C2496 PAD.n1674 VSS 0.036461f
C2497 PAD.n1676 VSS 0.036461f
C2498 PAD.n1677 VSS 0.036461f
C2499 PAD.n1678 VSS 0.036461f
C2500 PAD.n1680 VSS 0.036461f
C2501 PAD.n1681 VSS 0.036461f
C2502 PAD.n1682 VSS 0.036461f
C2503 PAD.n1683 VSS 0.030555f
C2504 PAD.n1684 VSS 0.023109f
C2505 PAD.n1685 VSS 0.023109f
C2506 PAD.n1687 VSS 0.036461f
C2507 PAD.n1689 VSS 0.036461f
C2508 PAD.n1691 VSS 0.036461f
C2509 PAD.n1692 VSS 0.036461f
C2510 PAD.n1693 VSS 0.036461f
C2511 PAD.n1694 VSS 0.036461f
C2512 PAD.n1695 VSS 0.036461f
C2513 PAD.n1696 VSS 0.036461f
C2514 PAD.n1697 VSS 0.036461f
C2515 PAD.n1699 VSS 0.036461f
C2516 PAD.n1701 VSS 0.036461f
C2517 PAD.n1703 VSS 0.036461f
C2518 PAD.n1704 VSS 0.036461f
C2519 PAD.n1705 VSS 0.036461f
C2520 PAD.n1706 VSS 0.036461f
C2521 PAD.n1707 VSS 0.036461f
C2522 PAD.n1708 VSS 0.036461f
C2523 PAD.n1709 VSS 0.036461f
C2524 PAD.n1711 VSS 0.036461f
C2525 PAD.n1713 VSS 0.036461f
C2526 PAD.n1715 VSS 0.036461f
C2527 PAD.n1716 VSS 0.036461f
C2528 PAD.n1717 VSS 0.036461f
C2529 PAD.n1718 VSS 0.036461f
C2530 PAD.n1719 VSS 0.036461f
C2531 PAD.n1720 VSS 0.036461f
C2532 PAD.n1721 VSS 0.036461f
C2533 PAD.n1723 VSS 0.036461f
C2534 PAD.n1725 VSS 0.036461f
C2535 PAD.n1727 VSS 0.036461f
C2536 PAD.n1728 VSS 0.036461f
C2537 PAD.n1729 VSS 0.036461f
C2538 PAD.n1730 VSS 0.036461f
C2539 PAD.n1731 VSS 0.036461f
C2540 PAD.n1732 VSS 0.036461f
C2541 PAD.n1733 VSS 0.036461f
C2542 PAD.n1735 VSS 0.036461f
C2543 PAD.n1737 VSS 0.036461f
C2544 PAD.n1739 VSS 0.036461f
C2545 PAD.n1740 VSS 0.036461f
C2546 PAD.n1741 VSS 0.036461f
C2547 PAD.n1742 VSS 0.036461f
C2548 PAD.n1743 VSS 0.036461f
C2549 PAD.n1744 VSS 0.036461f
C2550 PAD.n1745 VSS 0.036461f
C2551 PAD.n1747 VSS 0.036461f
C2552 PAD.n1749 VSS 0.036461f
C2553 PAD.n1751 VSS 0.036461f
C2554 PAD.n1752 VSS 0.036461f
C2555 PAD.n1753 VSS 0.036461f
C2556 PAD.n1754 VSS 0.036461f
C2557 PAD.n1755 VSS 0.036461f
C2558 PAD.n1756 VSS 0.036461f
C2559 PAD.n1757 VSS 0.036461f
C2560 PAD.n1759 VSS 0.036461f
C2561 PAD.n1761 VSS 0.036461f
C2562 PAD.n1763 VSS 0.036461f
C2563 PAD.n1764 VSS 0.036461f
C2564 PAD.n1765 VSS 0.036461f
C2565 PAD.n1766 VSS 0.036461f
C2566 PAD.n1767 VSS 0.036461f
C2567 PAD.n1768 VSS 0.036461f
C2568 PAD.n1769 VSS 0.036461f
C2569 PAD.n1771 VSS 0.036461f
C2570 PAD.n1773 VSS 0.036461f
C2571 PAD.n1775 VSS 0.036461f
C2572 PAD.n1776 VSS 0.036461f
C2573 PAD.n1777 VSS 0.036461f
C2574 PAD.n1778 VSS 0.036461f
C2575 PAD.n1779 VSS 0.036461f
C2576 PAD.n1780 VSS 0.036461f
C2577 PAD.n1781 VSS 0.036461f
C2578 PAD.n1783 VSS 0.036461f
C2579 PAD.n1785 VSS 0.036461f
C2580 PAD.n1787 VSS 0.036461f
C2581 PAD.n1788 VSS 0.036461f
C2582 PAD.n1789 VSS 0.036461f
C2583 PAD.n1790 VSS 0.036461f
C2584 PAD.n1791 VSS 0.036461f
C2585 PAD.n1792 VSS 0.036461f
C2586 PAD.n1793 VSS 0.036461f
C2587 PAD.n1795 VSS 0.036461f
C2588 PAD.n1797 VSS 0.036461f
C2589 PAD.n1799 VSS 0.036461f
C2590 PAD.n1800 VSS 0.036461f
C2591 PAD.n1801 VSS 0.036461f
C2592 PAD.n1802 VSS 0.036461f
C2593 PAD.n1803 VSS 0.036461f
C2594 PAD.n1804 VSS 0.036461f
C2595 PAD.n1805 VSS 0.036461f
C2596 PAD.n1807 VSS 0.036461f
C2597 PAD.n1809 VSS 0.036461f
C2598 PAD.n1811 VSS 0.036461f
C2599 PAD.n1812 VSS 0.036461f
C2600 PAD.n1813 VSS 0.036461f
C2601 PAD.n1814 VSS 0.036461f
C2602 PAD.n1815 VSS 0.036461f
C2603 PAD.n1816 VSS 0.036461f
C2604 PAD.n1817 VSS 0.036461f
C2605 PAD.n1819 VSS 0.036461f
C2606 PAD.n1821 VSS 0.036461f
C2607 PAD.n1823 VSS 0.036461f
C2608 PAD.n1824 VSS 0.036461f
C2609 PAD.n1825 VSS 0.036461f
C2610 PAD.n1826 VSS 0.036461f
C2611 PAD.n1827 VSS 0.036461f
C2612 PAD.n1828 VSS 0.036461f
C2613 PAD.n1829 VSS 0.036461f
C2614 PAD.n1831 VSS 0.036461f
C2615 PAD.n1833 VSS 0.036461f
C2616 PAD.n1835 VSS 0.036461f
C2617 PAD.n1836 VSS 0.036461f
C2618 PAD.n1837 VSS 0.036461f
C2619 PAD.n1838 VSS 0.036461f
C2620 PAD.n1839 VSS 0.036461f
C2621 PAD.n1840 VSS 0.036461f
C2622 PAD.n1841 VSS 0.036461f
C2623 PAD.n1843 VSS 0.036461f
C2624 PAD.n1845 VSS 0.036461f
C2625 PAD.n1847 VSS 0.036461f
C2626 PAD.n1848 VSS 0.036461f
C2627 PAD.n1849 VSS 0.036461f
C2628 PAD.n1850 VSS 0.036461f
C2629 PAD.n1851 VSS 0.036461f
C2630 PAD.n1852 VSS 0.036461f
C2631 PAD.n1853 VSS 0.036461f
C2632 PAD.n1855 VSS 0.036461f
C2633 PAD.n1857 VSS 0.036461f
C2634 PAD.n1859 VSS 0.036461f
C2635 PAD.n1860 VSS 0.036461f
C2636 PAD.n1861 VSS 0.036461f
C2637 PAD.n1862 VSS 0.036461f
C2638 PAD.n1863 VSS 0.036461f
C2639 PAD.n1864 VSS 0.036461f
C2640 PAD.n1865 VSS 0.036461f
C2641 PAD.n1867 VSS 0.036461f
C2642 PAD.n1869 VSS 0.036461f
C2643 PAD.n1871 VSS 0.036461f
C2644 PAD.n1872 VSS 0.036461f
C2645 PAD.n1873 VSS 0.036461f
C2646 PAD.n1874 VSS 0.036461f
C2647 PAD.n1875 VSS 0.036461f
C2648 PAD.n1876 VSS 0.036461f
C2649 PAD.n1877 VSS 0.036461f
C2650 PAD.n1879 VSS 0.036461f
C2651 PAD.n1881 VSS 0.036461f
C2652 PAD.n1883 VSS 0.036461f
C2653 PAD.n1884 VSS 0.036461f
C2654 PAD.n1885 VSS 0.036461f
C2655 PAD.n1886 VSS 0.036461f
C2656 PAD.n1887 VSS 0.036461f
C2657 PAD.n1888 VSS 0.036461f
C2658 PAD.n1889 VSS 0.036461f
C2659 PAD.n1891 VSS 0.036461f
C2660 PAD.n1893 VSS 0.036461f
C2661 PAD.n1895 VSS 0.036461f
C2662 PAD.n1896 VSS 0.036461f
C2663 PAD.n1897 VSS 0.036461f
C2664 PAD.n1898 VSS 0.036461f
C2665 PAD.n1899 VSS 0.036461f
C2666 PAD.n1900 VSS 0.036461f
C2667 PAD.n1901 VSS 0.036461f
C2668 PAD.n1903 VSS 0.036461f
C2669 PAD.n1905 VSS 0.036461f
C2670 PAD.n1907 VSS 0.036461f
C2671 PAD.n1908 VSS 0.036461f
C2672 PAD.n1909 VSS 0.036461f
C2673 PAD.n1910 VSS 0.036461f
C2674 PAD.n1911 VSS 0.036461f
C2675 PAD.n1912 VSS 0.036461f
C2676 PAD.n1913 VSS 0.036461f
C2677 PAD.n1915 VSS 0.036461f
C2678 PAD.n1917 VSS 0.036461f
C2679 PAD.n1919 VSS 0.036461f
C2680 PAD.n1920 VSS 0.036461f
C2681 PAD.n1921 VSS 0.036461f
C2682 PAD.n1922 VSS 0.036461f
C2683 PAD.n1923 VSS 0.036461f
C2684 PAD.n1924 VSS 0.036461f
C2685 PAD.n1925 VSS 0.036461f
C2686 PAD.n1927 VSS 0.036461f
C2687 PAD.n1929 VSS 0.036461f
C2688 PAD.n1930 VSS 0.036461f
C2689 PAD.n1931 VSS 0.023109f
C2690 PAD.n1932 VSS 0.03338f
C2691 PAD.n1933 VSS 0.062274f
C2692 PAD.n1934 VSS 0.069765f
C2693 PAD.n1935 VSS 0.069765f
C2694 PAD.n1936 VSS 0.700534f
C2695 PAD.n1937 VSS 0.049115f
C2696 PAD.n1938 VSS 0.049115f
C2697 PAD.n1939 VSS 0.033773f
C2698 PAD.n1940 VSS 0.029436f
C2699 PAD.n1941 VSS 0.029436f
C2700 PAD.n1942 VSS 0.439067f
C2701 PAD.n1984 VSS 0.023109f
C2702 PAD.n1985 VSS 0.611734f
C2703 PAD.n1986 VSS 0.439067f
C2704 PAD.n1987 VSS 0.023109f
C2705 PAD.n1988 VSS 0.37f
C2706 PAD.n1989 VSS 0.036461f
C2707 PAD.n1990 VSS 0.036461f
C2708 PAD.n1991 VSS 0.036461f
C2709 PAD.n1992 VSS 0.036461f
C2710 PAD.n1993 VSS 0.036461f
C2711 PAD.n1994 VSS 0.036461f
C2712 PAD.n1995 VSS 0.036461f
C2713 PAD.n1996 VSS 0.036461f
C2714 PAD.n1997 VSS 0.036461f
C2715 PAD.n1998 VSS 0.036461f
C2716 PAD.n1999 VSS 0.036461f
C2717 PAD.n2000 VSS 0.036461f
C2718 PAD.n2001 VSS 0.036461f
C2719 PAD.n2002 VSS 0.036461f
C2720 PAD.n2003 VSS 0.036461f
C2721 PAD.n2004 VSS 0.036461f
C2722 PAD.n2005 VSS 0.036461f
C2723 PAD.n2006 VSS 0.036461f
C2724 PAD.n2007 VSS 0.036461f
C2725 PAD.n2008 VSS 0.036461f
C2726 PAD.n2009 VSS 0.036461f
C2727 PAD.n2010 VSS 0.036461f
C2728 PAD.n2011 VSS 0.036461f
C2729 PAD.n2012 VSS 0.036461f
C2730 PAD.n2013 VSS 0.036461f
C2731 PAD.n2014 VSS 0.036461f
C2732 PAD.n2015 VSS 0.036461f
C2733 PAD.n2016 VSS 0.036461f
C2734 PAD.n2017 VSS 0.036461f
C2735 PAD.n2018 VSS 0.036461f
C2736 PAD.n2019 VSS 0.036461f
C2737 PAD.n2020 VSS 0.036461f
C2738 PAD.n2021 VSS 0.036461f
C2739 PAD.n2022 VSS 0.036461f
C2740 PAD.n2023 VSS 0.036461f
C2741 PAD.n2024 VSS 0.036461f
C2742 PAD.n2025 VSS 0.036461f
C2743 PAD.n2026 VSS 0.036461f
C2744 PAD.n2027 VSS 0.036461f
C2745 PAD.n2028 VSS 0.036461f
C2746 PAD.n2030 VSS 0.036461f
C2747 PAD.n2031 VSS 0.036461f
C2748 PAD.n2032 VSS 0.046286f
C2749 PAD.n2033 VSS 0.048386f
C2750 PAD.n2034 VSS 0.050221f
C2751 PAD.n2035 VSS 0.064139f
C2752 PAD.n2036 VSS 0.069765f
C2753 PAD.n2037 VSS 0.611734f
C2754 PAD.n2038 VSS 0.047905f
C2755 PAD.n2039 VSS 0.047905f
C2756 PAD.n2040 VSS 0.030555f
C2757 PAD.n2041 VSS 0.042895f
C2758 PAD.n2042 VSS 0.049115f
C2759 PAD.n2043 VSS 0.029436f
C2760 PAD.n2044 VSS 0.049115f
C2761 PAD.n2045 VSS 0.029436f
C2762 PAD.n2046 VSS 0.3108f
C2763 PAD.n2088 VSS 0.023109f
C2764 PAD.n2089 VSS 0.3108f
C2765 PAD.n2090 VSS 0.023109f
C2766 PAD.n2091 VSS 0.611735f
C2767 PAD.n2092 VSS 0.036461f
C2768 PAD.n2093 VSS 0.036461f
C2769 PAD.n2094 VSS 0.036461f
C2770 PAD.n2095 VSS 0.036461f
C2771 PAD.n2096 VSS 0.036461f
C2772 PAD.n2097 VSS 0.036461f
C2773 PAD.n2098 VSS 0.036461f
C2774 PAD.n2099 VSS 0.036461f
C2775 PAD.n2100 VSS 0.036461f
C2776 PAD.n2101 VSS 0.036461f
C2777 PAD.n2102 VSS 0.036461f
C2778 PAD.n2103 VSS 0.036461f
C2779 PAD.n2104 VSS 0.036461f
C2780 PAD.n2105 VSS 0.036461f
C2781 PAD.n2106 VSS 0.036461f
C2782 PAD.n2107 VSS 0.036461f
C2783 PAD.n2108 VSS 0.036461f
C2784 PAD.n2109 VSS 0.036461f
C2785 PAD.n2110 VSS 0.036461f
C2786 PAD.n2111 VSS 0.036461f
C2787 PAD.n2112 VSS 0.036461f
C2788 PAD.n2113 VSS 0.036461f
C2789 PAD.n2114 VSS 0.036461f
C2790 PAD.n2115 VSS 0.036461f
C2791 PAD.n2116 VSS 0.036461f
C2792 PAD.n2117 VSS 0.036461f
C2793 PAD.n2118 VSS 0.036461f
C2794 PAD.n2119 VSS 0.036461f
C2795 PAD.n2120 VSS 0.036461f
C2796 PAD.n2121 VSS 0.036461f
C2797 PAD.n2122 VSS 0.036461f
C2798 PAD.n2123 VSS 0.036461f
C2799 PAD.n2124 VSS 0.036461f
C2800 PAD.n2125 VSS 0.036461f
C2801 PAD.n2126 VSS 0.036461f
C2802 PAD.n2127 VSS 0.036461f
C2803 PAD.n2128 VSS 0.036461f
C2804 PAD.n2129 VSS 0.036461f
C2805 PAD.n2130 VSS 0.036461f
C2806 PAD.n2131 VSS 0.036461f
C2807 PAD.n2133 VSS 0.036461f
C2808 PAD.n2134 VSS 0.036461f
C2809 PAD.n2135 VSS 0.046286f
C2810 PAD.n2136 VSS 0.069765f
C2811 PAD.n2137 VSS 0.036159f
C2812 PAD.n2138 VSS 0.069765f
C2813 PAD.n2139 VSS 0.498267f
C2814 PAD.n2140 VSS 0.029436f
C2815 PAD.n2141 VSS 0.029436f
C2816 PAD.n2142 VSS 0.030555f
C2817 PAD.n2143 VSS 0.042895f
C2818 PAD.n2144 VSS 0.049115f
C2819 PAD.n2145 VSS 0.049115f
C2820 PAD.n2146 VSS 0.409467f
C2821 PAD.n2147 VSS 0.039761f
C2822 PAD.n2148 VSS 0.039761f
C2823 PAD.n2149 VSS 0.069765f
C2824 PAD.n2150 VSS 0.036461f
C2825 PAD.n2151 VSS 0.023109f
C2826 PAD.n2152 VSS 0.036461f
C2827 PAD.n2155 VSS 0.036461f
C2828 PAD.n2156 VSS 0.036461f
C2829 PAD.n2157 VSS 0.036461f
C2830 PAD.n2158 VSS 0.036461f
C2831 PAD.n2160 VSS 0.036461f
C2832 PAD.n2161 VSS 0.036461f
C2833 PAD.n2162 VSS 0.036461f
C2834 PAD.n2164 VSS 0.036461f
C2835 PAD.n2165 VSS 0.036461f
C2836 PAD.n2166 VSS 0.036461f
C2837 PAD.n2168 VSS 0.036461f
C2838 PAD.n2169 VSS 0.036461f
C2839 PAD.n2170 VSS 0.036461f
C2840 PAD.n2172 VSS 0.036461f
C2841 PAD.n2173 VSS 0.036461f
C2842 PAD.n2174 VSS 0.036461f
C2843 PAD.n2176 VSS 0.036461f
C2844 PAD.n2177 VSS 0.036461f
C2845 PAD.n2178 VSS 0.036461f
C2846 PAD.n2180 VSS 0.036461f
C2847 PAD.n2181 VSS 0.036461f
C2848 PAD.n2182 VSS 0.036461f
C2849 PAD.n2184 VSS 0.036461f
C2850 PAD.n2185 VSS 0.036461f
C2851 PAD.n2186 VSS 0.036461f
C2852 PAD.n2188 VSS 0.036461f
C2853 PAD.n2189 VSS 0.036461f
C2854 PAD.n2190 VSS 0.036461f
C2855 PAD.n2192 VSS 0.036461f
C2856 PAD.n2193 VSS 0.036461f
C2857 PAD.n2194 VSS 0.036461f
C2858 PAD.n2196 VSS 0.036461f
C2859 PAD.n2197 VSS 0.036461f
C2860 PAD.n2198 VSS 0.036461f
C2861 PAD.n2200 VSS 0.036461f
C2862 PAD.n2201 VSS 0.036461f
C2863 PAD.n2202 VSS 0.036461f
C2864 PAD.n2204 VSS 0.036461f
C2865 PAD.n2205 VSS 0.036461f
C2866 PAD.n2206 VSS 0.036461f
C2867 PAD.n2208 VSS 0.036461f
C2868 PAD.n2209 VSS 0.036461f
C2869 PAD.n2210 VSS 0.036461f
C2870 PAD.n2212 VSS 0.036461f
C2871 PAD.n2213 VSS 0.036461f
C2872 PAD.n2214 VSS 0.036461f
C2873 PAD.n2216 VSS 0.036461f
C2874 PAD.n2217 VSS 0.036461f
C2875 PAD.n2218 VSS 0.036461f
C2876 PAD.n2220 VSS 0.036461f
C2877 PAD.n2221 VSS 0.036461f
C2878 PAD.n2222 VSS 0.036461f
C2879 PAD.n2224 VSS 0.036461f
C2880 PAD.n2225 VSS 0.036461f
C2881 PAD.n2226 VSS 0.036461f
C2882 PAD.n2228 VSS 0.036461f
C2883 PAD.n2229 VSS 0.036461f
C2884 PAD.n2230 VSS 0.036461f
C2885 PAD.n2232 VSS 0.036461f
C2886 PAD.n2233 VSS 0.036461f
C2887 PAD.n2234 VSS 0.036461f
C2888 PAD.n2235 VSS 0.023109f
C2889 PAD.n2236 VSS 0.023109f
C2890 PAD.n2238 VSS 0.036461f
C2891 PAD.n2240 VSS 0.036461f
C2892 PAD.n2242 VSS 0.036461f
C2893 PAD.n2243 VSS 0.036461f
C2894 PAD.n2244 VSS 0.036461f
C2895 PAD.n2245 VSS 0.036461f
C2896 PAD.n2246 VSS 0.036461f
C2897 PAD.n2247 VSS 0.036461f
C2898 PAD.n2248 VSS 0.036461f
C2899 PAD.n2250 VSS 0.036461f
C2900 PAD.n2252 VSS 0.036461f
C2901 PAD.n2254 VSS 0.036461f
C2902 PAD.n2255 VSS 0.036461f
C2903 PAD.n2256 VSS 0.036461f
C2904 PAD.n2257 VSS 0.036461f
C2905 PAD.n2258 VSS 0.036461f
C2906 PAD.n2259 VSS 0.036461f
C2907 PAD.n2260 VSS 0.036461f
C2908 PAD.n2262 VSS 0.036461f
C2909 PAD.n2264 VSS 0.036461f
C2910 PAD.n2266 VSS 0.036461f
C2911 PAD.n2267 VSS 0.036461f
C2912 PAD.n2268 VSS 0.036461f
C2913 PAD.n2269 VSS 0.036461f
C2914 PAD.n2270 VSS 0.036461f
C2915 PAD.n2271 VSS 0.036461f
C2916 PAD.n2272 VSS 0.036461f
C2917 PAD.n2274 VSS 0.036461f
C2918 PAD.n2276 VSS 0.036461f
C2919 PAD.n2278 VSS 0.036461f
C2920 PAD.n2279 VSS 0.036461f
C2921 PAD.n2280 VSS 0.036461f
C2922 PAD.n2281 VSS 0.036461f
C2923 PAD.n2282 VSS 0.036461f
C2924 PAD.n2283 VSS 0.036461f
C2925 PAD.n2284 VSS 0.036461f
C2926 PAD.n2286 VSS 0.036461f
C2927 PAD.n2288 VSS 0.036461f
C2928 PAD.n2290 VSS 0.036461f
C2929 PAD.n2291 VSS 0.036461f
C2930 PAD.n2292 VSS 0.036461f
C2931 PAD.n2293 VSS 0.036461f
C2932 PAD.n2294 VSS 0.036461f
C2933 PAD.n2295 VSS 0.036461f
C2934 PAD.n2296 VSS 0.036461f
C2935 PAD.n2298 VSS 0.036461f
C2936 PAD.n2300 VSS 0.036461f
C2937 PAD.n2302 VSS 0.036461f
C2938 PAD.n2303 VSS 0.036461f
C2939 PAD.n2304 VSS 0.036461f
C2940 PAD.n2305 VSS 0.036461f
C2941 PAD.n2306 VSS 0.036461f
C2942 PAD.n2307 VSS 0.036461f
C2943 PAD.n2308 VSS 0.036461f
C2944 PAD.n2310 VSS 0.036461f
C2945 PAD.n2312 VSS 0.036461f
C2946 PAD.n2314 VSS 0.036461f
C2947 PAD.n2315 VSS 0.036461f
C2948 PAD.n2316 VSS 0.036461f
C2949 PAD.n2317 VSS 0.036461f
C2950 PAD.n2318 VSS 0.036461f
C2951 PAD.n2319 VSS 0.036461f
C2952 PAD.n2320 VSS 0.036461f
C2953 PAD.n2322 VSS 0.036461f
C2954 PAD.n2324 VSS 0.036461f
C2955 PAD.n2326 VSS 0.036461f
C2956 PAD.n2327 VSS 0.036461f
C2957 PAD.n2328 VSS 0.036461f
C2958 PAD.n2329 VSS 0.036461f
C2959 PAD.n2330 VSS 0.036461f
C2960 PAD.n2331 VSS 0.036461f
C2961 PAD.n2332 VSS 0.036461f
C2962 PAD.n2334 VSS 0.036461f
C2963 PAD.n2336 VSS 0.036461f
C2964 PAD.n2338 VSS 0.036461f
C2965 PAD.n2339 VSS 0.036461f
C2966 PAD.n2340 VSS 0.036461f
C2967 PAD.n2341 VSS 0.036461f
C2968 PAD.n2342 VSS 0.036461f
C2969 PAD.n2343 VSS 0.036461f
C2970 PAD.n2344 VSS 0.036461f
C2971 PAD.n2346 VSS 0.036461f
C2972 PAD.n2348 VSS 0.036461f
C2973 PAD.n2350 VSS 0.036461f
C2974 PAD.n2351 VSS 0.036461f
C2975 PAD.n2352 VSS 0.036461f
C2976 PAD.n2353 VSS 0.036461f
C2977 PAD.n2354 VSS 0.036461f
C2978 PAD.n2355 VSS 0.036461f
C2979 PAD.n2356 VSS 0.036461f
C2980 PAD.n2358 VSS 0.036461f
C2981 PAD.n2360 VSS 0.036461f
C2982 PAD.n2362 VSS 0.036461f
C2983 PAD.n2363 VSS 0.036461f
C2984 PAD.n2364 VSS 0.036461f
C2985 PAD.n2365 VSS 0.036461f
C2986 PAD.n2366 VSS 0.036461f
C2987 PAD.n2367 VSS 0.036461f
C2988 PAD.n2368 VSS 0.036461f
C2989 PAD.n2370 VSS 0.036461f
C2990 PAD.n2372 VSS 0.036461f
C2991 PAD.n2374 VSS 0.036461f
C2992 PAD.n2375 VSS 0.036461f
C2993 PAD.n2376 VSS 0.036461f
C2994 PAD.n2377 VSS 0.036461f
C2995 PAD.n2378 VSS 0.036461f
C2996 PAD.n2379 VSS 0.036461f
C2997 PAD.n2380 VSS 0.036461f
C2998 PAD.n2382 VSS 0.036461f
C2999 PAD.n2384 VSS 0.036461f
C3000 PAD.n2386 VSS 0.036461f
C3001 PAD.n2387 VSS 0.036461f
C3002 PAD.n2388 VSS 0.036461f
C3003 PAD.n2389 VSS 0.036461f
C3004 PAD.n2390 VSS 0.036461f
C3005 PAD.n2391 VSS 0.036461f
C3006 PAD.n2392 VSS 0.036461f
C3007 PAD.n2394 VSS 0.036461f
C3008 PAD.n2396 VSS 0.036461f
C3009 PAD.n2398 VSS 0.036461f
C3010 PAD.n2399 VSS 0.036461f
C3011 PAD.n2400 VSS 0.036461f
C3012 PAD.n2401 VSS 0.036461f
C3013 PAD.n2402 VSS 0.036461f
C3014 PAD.n2403 VSS 0.036461f
C3015 PAD.n2404 VSS 0.036461f
C3016 PAD.n2406 VSS 0.036461f
C3017 PAD.n2408 VSS 0.036461f
C3018 PAD.n2410 VSS 0.036461f
C3019 PAD.n2411 VSS 0.036461f
C3020 PAD.n2412 VSS 0.036461f
C3021 PAD.n2413 VSS 0.036461f
C3022 PAD.n2414 VSS 0.036461f
C3023 PAD.n2415 VSS 0.036461f
C3024 PAD.n2416 VSS 0.036461f
C3025 PAD.n2418 VSS 0.036461f
C3026 PAD.n2420 VSS 0.036461f
C3027 PAD.n2422 VSS 0.036461f
C3028 PAD.n2423 VSS 0.036461f
C3029 PAD.n2424 VSS 0.036461f
C3030 PAD.n2425 VSS 0.036461f
C3031 PAD.n2426 VSS 0.036461f
C3032 PAD.n2427 VSS 0.036461f
C3033 PAD.n2428 VSS 0.036461f
C3034 PAD.n2430 VSS 0.036461f
C3035 PAD.n2432 VSS 0.036461f
C3036 PAD.n2434 VSS 0.036461f
C3037 PAD.n2435 VSS 0.036461f
C3038 PAD.n2436 VSS 0.036461f
C3039 PAD.n2437 VSS 0.036461f
C3040 PAD.n2438 VSS 0.036461f
C3041 PAD.n2439 VSS 0.036461f
C3042 PAD.n2440 VSS 0.036461f
C3043 PAD.n2442 VSS 0.036461f
C3044 PAD.n2444 VSS 0.036461f
C3045 PAD.n2446 VSS 0.036461f
C3046 PAD.n2447 VSS 0.036461f
C3047 PAD.n2448 VSS 0.036461f
C3048 PAD.n2449 VSS 0.036461f
C3049 PAD.n2450 VSS 0.036461f
C3050 PAD.n2451 VSS 0.036461f
C3051 PAD.n2452 VSS 0.036461f
C3052 PAD.n2454 VSS 0.036461f
C3053 PAD.n2456 VSS 0.036461f
C3054 PAD.n2458 VSS 0.036461f
C3055 PAD.n2459 VSS 0.036461f
C3056 PAD.n2460 VSS 0.036461f
C3057 PAD.n2461 VSS 0.036461f
C3058 PAD.n2462 VSS 0.036461f
C3059 PAD.n2463 VSS 0.036461f
C3060 PAD.n2464 VSS 0.036461f
C3061 PAD.n2466 VSS 0.036461f
C3062 PAD.n2468 VSS 0.036461f
C3063 PAD.n2470 VSS 0.036461f
C3064 PAD.n2471 VSS 0.036461f
C3065 PAD.n2472 VSS 0.036461f
C3066 PAD.n2473 VSS 0.036461f
C3067 PAD.n2474 VSS 0.036461f
C3068 PAD.n2475 VSS 0.036461f
C3069 PAD.n2476 VSS 0.036461f
C3070 PAD.n2478 VSS 0.036461f
C3071 PAD.n2480 VSS 0.036461f
C3072 PAD.n2481 VSS 0.036461f
C3073 PAD.n2482 VSS 0.023109f
C3074 PAD.n2483 VSS 0.03338f
C3075 PAD.n2484 VSS 0.062274f
C3076 PAD.n2485 VSS 0.069765f
C3077 PAD.n2486 VSS 0.069765f
C3078 PAD.n2487 VSS 0.231867f
C3079 PAD.n2488 VSS 0.029436f
C3080 PAD.n2489 VSS 0.029436f
C3081 PAD.n2490 VSS 0.030555f
C3082 PAD.n2491 VSS 0.042895f
C3083 PAD.n2492 VSS 0.049115f
C3084 PAD.n2493 VSS 0.049115f
C3085 PAD.n2494 VSS 0.143067f
C3086 PAD.n2495 VSS 0.039761f
C3087 PAD.n2496 VSS 0.039761f
C3088 PAD.n2497 VSS 0.036461f
C3089 PAD.n2498 VSS 0.023109f
C3090 PAD.n2499 VSS 0.036461f
C3091 PAD.n2502 VSS 0.036461f
C3092 PAD.n2503 VSS 0.036461f
C3093 PAD.n2504 VSS 0.036461f
C3094 PAD.n2505 VSS 0.036461f
C3095 PAD.n2507 VSS 0.036461f
C3096 PAD.n2508 VSS 0.036461f
C3097 PAD.n2509 VSS 0.036461f
C3098 PAD.n2511 VSS 0.036461f
C3099 PAD.n2512 VSS 0.036461f
C3100 PAD.n2513 VSS 0.036461f
C3101 PAD.n2515 VSS 0.036461f
C3102 PAD.n2516 VSS 0.036461f
C3103 PAD.n2517 VSS 0.036461f
C3104 PAD.n2519 VSS 0.036461f
C3105 PAD.n2520 VSS 0.036461f
C3106 PAD.n2521 VSS 0.036461f
C3107 PAD.n2523 VSS 0.036461f
C3108 PAD.n2524 VSS 0.036461f
C3109 PAD.n2525 VSS 0.036461f
C3110 PAD.n2527 VSS 0.036461f
C3111 PAD.n2528 VSS 0.036461f
C3112 PAD.n2529 VSS 0.036461f
C3113 PAD.n2531 VSS 0.036461f
C3114 PAD.n2532 VSS 0.036461f
C3115 PAD.n2533 VSS 0.036461f
C3116 PAD.n2535 VSS 0.036461f
C3117 PAD.n2536 VSS 0.036461f
C3118 PAD.n2537 VSS 0.036461f
C3119 PAD.n2539 VSS 0.036461f
C3120 PAD.n2540 VSS 0.036461f
C3121 PAD.n2541 VSS 0.036461f
C3122 PAD.n2543 VSS 0.036461f
C3123 PAD.n2544 VSS 0.036461f
C3124 PAD.n2545 VSS 0.036461f
C3125 PAD.n2547 VSS 0.036461f
C3126 PAD.n2548 VSS 0.036461f
C3127 PAD.n2549 VSS 0.036461f
C3128 PAD.n2551 VSS 0.036461f
C3129 PAD.n2552 VSS 0.036461f
C3130 PAD.n2553 VSS 0.036461f
C3131 PAD.n2555 VSS 0.036461f
C3132 PAD.n2556 VSS 0.036461f
C3133 PAD.n2557 VSS 0.036461f
C3134 PAD.n2559 VSS 0.036461f
C3135 PAD.n2560 VSS 0.036461f
C3136 PAD.n2561 VSS 0.036461f
C3137 PAD.n2563 VSS 0.036461f
C3138 PAD.n2564 VSS 0.036461f
C3139 PAD.n2565 VSS 0.036461f
C3140 PAD.n2567 VSS 0.036461f
C3141 PAD.n2568 VSS 0.036461f
C3142 PAD.n2569 VSS 0.036461f
C3143 PAD.n2571 VSS 0.036461f
C3144 PAD.n2572 VSS 0.036461f
C3145 PAD.n2573 VSS 0.036461f
C3146 PAD.n2575 VSS 0.036461f
C3147 PAD.n2576 VSS 0.036461f
C3148 PAD.n2577 VSS 0.036461f
C3149 PAD.n2579 VSS 0.036461f
C3150 PAD.n2580 VSS 0.036461f
C3151 PAD.n2581 VSS 0.036461f
C3152 PAD.n2582 VSS 0.023109f
C3153 PAD.n2583 VSS 0.023109f
C3154 PAD.n2585 VSS 0.036461f
C3155 PAD.n2587 VSS 0.036461f
C3156 PAD.n2589 VSS 0.036461f
C3157 PAD.n2590 VSS 0.036461f
C3158 PAD.n2591 VSS 0.036461f
C3159 PAD.n2592 VSS 0.036461f
C3160 PAD.n2593 VSS 0.036461f
C3161 PAD.n2594 VSS 0.036461f
C3162 PAD.n2595 VSS 0.036461f
C3163 PAD.n2597 VSS 0.036461f
C3164 PAD.n2599 VSS 0.036461f
C3165 PAD.n2601 VSS 0.036461f
C3166 PAD.n2602 VSS 0.036461f
C3167 PAD.n2603 VSS 0.036461f
C3168 PAD.n2604 VSS 0.036461f
C3169 PAD.n2605 VSS 0.036461f
C3170 PAD.n2606 VSS 0.036461f
C3171 PAD.n2607 VSS 0.036461f
C3172 PAD.n2609 VSS 0.036461f
C3173 PAD.n2611 VSS 0.036461f
C3174 PAD.n2613 VSS 0.036461f
C3175 PAD.n2614 VSS 0.036461f
C3176 PAD.n2615 VSS 0.036461f
C3177 PAD.n2616 VSS 0.036461f
C3178 PAD.n2617 VSS 0.036461f
C3179 PAD.n2618 VSS 0.036461f
C3180 PAD.n2619 VSS 0.036461f
C3181 PAD.n2621 VSS 0.036461f
C3182 PAD.n2623 VSS 0.036461f
C3183 PAD.n2625 VSS 0.036461f
C3184 PAD.n2626 VSS 0.036461f
C3185 PAD.n2627 VSS 0.036461f
C3186 PAD.n2628 VSS 0.036461f
C3187 PAD.n2629 VSS 0.036461f
C3188 PAD.n2630 VSS 0.036461f
C3189 PAD.n2631 VSS 0.036461f
C3190 PAD.n2633 VSS 0.036461f
C3191 PAD.n2635 VSS 0.036461f
C3192 PAD.n2637 VSS 0.036461f
C3193 PAD.n2638 VSS 0.036461f
C3194 PAD.n2639 VSS 0.036461f
C3195 PAD.n2640 VSS 0.036461f
C3196 PAD.n2641 VSS 0.036461f
C3197 PAD.n2642 VSS 0.036461f
C3198 PAD.n2643 VSS 0.036461f
C3199 PAD.n2645 VSS 0.036461f
C3200 PAD.n2647 VSS 0.036461f
C3201 PAD.n2649 VSS 0.036461f
C3202 PAD.n2650 VSS 0.036461f
C3203 PAD.n2651 VSS 0.036461f
C3204 PAD.n2652 VSS 0.036461f
C3205 PAD.n2653 VSS 0.036461f
C3206 PAD.n2654 VSS 0.036461f
C3207 PAD.n2655 VSS 0.036461f
C3208 PAD.n2657 VSS 0.036461f
C3209 PAD.n2659 VSS 0.036461f
C3210 PAD.n2661 VSS 0.036461f
C3211 PAD.n2662 VSS 0.036461f
C3212 PAD.n2663 VSS 0.036461f
C3213 PAD.n2664 VSS 0.036461f
C3214 PAD.n2665 VSS 0.036461f
C3215 PAD.n2666 VSS 0.036461f
C3216 PAD.n2667 VSS 0.036461f
C3217 PAD.n2669 VSS 0.036461f
C3218 PAD.n2671 VSS 0.036461f
C3219 PAD.n2673 VSS 0.036461f
C3220 PAD.n2674 VSS 0.036461f
C3221 PAD.n2675 VSS 0.036461f
C3222 PAD.n2676 VSS 0.036461f
C3223 PAD.n2677 VSS 0.036461f
C3224 PAD.n2678 VSS 0.036461f
C3225 PAD.n2679 VSS 0.036461f
C3226 PAD.n2681 VSS 0.036461f
C3227 PAD.n2683 VSS 0.036461f
C3228 PAD.n2685 VSS 0.036461f
C3229 PAD.n2686 VSS 0.036461f
C3230 PAD.n2687 VSS 0.036461f
C3231 PAD.n2688 VSS 0.036461f
C3232 PAD.n2689 VSS 0.036461f
C3233 PAD.n2690 VSS 0.036461f
C3234 PAD.n2691 VSS 0.036461f
C3235 PAD.n2693 VSS 0.036461f
C3236 PAD.n2695 VSS 0.036461f
C3237 PAD.n2697 VSS 0.036461f
C3238 PAD.n2698 VSS 0.036461f
C3239 PAD.n2699 VSS 0.036461f
C3240 PAD.n2700 VSS 0.036461f
C3241 PAD.n2701 VSS 0.036461f
C3242 PAD.n2702 VSS 0.036461f
C3243 PAD.n2703 VSS 0.036461f
C3244 PAD.n2705 VSS 0.036461f
C3245 PAD.n2707 VSS 0.036461f
C3246 PAD.n2709 VSS 0.036461f
C3247 PAD.n2710 VSS 0.036461f
C3248 PAD.n2711 VSS 0.036461f
C3249 PAD.n2712 VSS 0.036461f
C3250 PAD.n2713 VSS 0.036461f
C3251 PAD.n2714 VSS 0.036461f
C3252 PAD.n2715 VSS 0.036461f
C3253 PAD.n2717 VSS 0.036461f
C3254 PAD.n2719 VSS 0.036461f
C3255 PAD.n2721 VSS 0.036461f
C3256 PAD.n2722 VSS 0.036461f
C3257 PAD.n2723 VSS 0.036461f
C3258 PAD.n2724 VSS 0.036461f
C3259 PAD.n2725 VSS 0.036461f
C3260 PAD.n2726 VSS 0.036461f
C3261 PAD.n2727 VSS 0.036461f
C3262 PAD.n2729 VSS 0.036461f
C3263 PAD.n2731 VSS 0.036461f
C3264 PAD.n2733 VSS 0.036461f
C3265 PAD.n2734 VSS 0.036461f
C3266 PAD.n2735 VSS 0.036461f
C3267 PAD.n2736 VSS 0.036461f
C3268 PAD.n2737 VSS 0.036461f
C3269 PAD.n2738 VSS 0.036461f
C3270 PAD.n2739 VSS 0.036461f
C3271 PAD.n2741 VSS 0.036461f
C3272 PAD.n2743 VSS 0.036461f
C3273 PAD.n2745 VSS 0.036461f
C3274 PAD.n2746 VSS 0.036461f
C3275 PAD.n2747 VSS 0.036461f
C3276 PAD.n2748 VSS 0.036461f
C3277 PAD.n2749 VSS 0.036461f
C3278 PAD.n2750 VSS 0.036461f
C3279 PAD.n2751 VSS 0.036461f
C3280 PAD.n2753 VSS 0.036461f
C3281 PAD.n2755 VSS 0.036461f
C3282 PAD.n2757 VSS 0.036461f
C3283 PAD.n2758 VSS 0.036461f
C3284 PAD.n2759 VSS 0.036461f
C3285 PAD.n2760 VSS 0.036461f
C3286 PAD.n2761 VSS 0.036461f
C3287 PAD.n2762 VSS 0.036461f
C3288 PAD.n2763 VSS 0.036461f
C3289 PAD.n2765 VSS 0.036461f
C3290 PAD.n2767 VSS 0.036461f
C3291 PAD.n2769 VSS 0.036461f
C3292 PAD.n2770 VSS 0.036461f
C3293 PAD.n2771 VSS 0.036461f
C3294 PAD.n2772 VSS 0.036461f
C3295 PAD.n2773 VSS 0.036461f
C3296 PAD.n2774 VSS 0.036461f
C3297 PAD.n2775 VSS 0.036461f
C3298 PAD.n2777 VSS 0.036461f
C3299 PAD.n2779 VSS 0.036461f
C3300 PAD.n2781 VSS 0.036461f
C3301 PAD.n2782 VSS 0.036461f
C3302 PAD.n2783 VSS 0.036461f
C3303 PAD.n2784 VSS 0.036461f
C3304 PAD.n2785 VSS 0.036461f
C3305 PAD.n2786 VSS 0.036461f
C3306 PAD.n2787 VSS 0.036461f
C3307 PAD.n2789 VSS 0.036461f
C3308 PAD.n2791 VSS 0.036461f
C3309 PAD.n2793 VSS 0.036461f
C3310 PAD.n2794 VSS 0.036461f
C3311 PAD.n2795 VSS 0.036461f
C3312 PAD.n2796 VSS 0.036461f
C3313 PAD.n2797 VSS 0.036461f
C3314 PAD.n2798 VSS 0.036461f
C3315 PAD.n2799 VSS 0.036461f
C3316 PAD.n2801 VSS 0.036461f
C3317 PAD.n2803 VSS 0.036461f
C3318 PAD.n2805 VSS 0.036461f
C3319 PAD.n2806 VSS 0.036461f
C3320 PAD.n2807 VSS 0.036461f
C3321 PAD.n2808 VSS 0.036461f
C3322 PAD.n2809 VSS 0.036461f
C3323 PAD.n2810 VSS 0.036461f
C3324 PAD.n2811 VSS 0.036461f
C3325 PAD.n2813 VSS 0.036461f
C3326 PAD.n2815 VSS 0.036461f
C3327 PAD.n2817 VSS 0.036461f
C3328 PAD.n2818 VSS 0.036461f
C3329 PAD.n2819 VSS 0.036461f
C3330 PAD.n2820 VSS 0.036461f
C3331 PAD.n2821 VSS 0.036461f
C3332 PAD.n2822 VSS 0.036461f
C3333 PAD.n2823 VSS 0.036461f
C3334 PAD.n2825 VSS 0.036461f
C3335 PAD.n2827 VSS 0.036461f
C3336 PAD.n2828 VSS 0.036461f
C3337 PAD.n2829 VSS 0.023109f
C3338 PAD.n2830 VSS 0.03338f
C3339 PAD.n2831 VSS 0.062274f
C3340 PAD.n2832 VSS 0.069765f
C3341 PAD.n2833 VSS 0.069765f
C3342 PAD.n2834 VSS 0.078933f
C3343 PAD.n2876 VSS 0.023109f
C3344 PAD.n2877 VSS 0.023109f
C3345 PAD.n2878 VSS 0.029436f
C3346 PAD.n2879 VSS 0.123333f
C3347 PAD.n2880 VSS 0.036461f
C3348 PAD.n2881 VSS 0.036461f
C3349 PAD.n2882 VSS 0.034286f
C3350 PAD.n2883 VSS 0.029436f
C3351 PAD.n2884 VSS 0.069765f
C3352 PAD.n2885 VSS 0.039761f
C3353 PAD.n2886 VSS 0.069765f
C3354 PAD.n2887 VSS 0.039761f
C3355 PAD.n2888 VSS 0.046286f
C3356 PAD.n2889 VSS 0.039761f
C3357 PAD.n2890 VSS 0.039761f
C3358 PAD.n2891 VSS 0.300934f
C3359 PAD.n2892 VSS 0.700534f
C3360 PAD.n2893 VSS 0.029919f
C3361 PAD.n2894 VSS 0.567334f
C3362 PAD.n2895 VSS 0.039258f
C3363 PAD.n2896 VSS 0.029919f
C3364 PAD.n2897 VSS 0.039258f
C3365 PAD.n2898 VSS 0.030555f
C3366 PAD.n2899 VSS 0.042895f
C3367 PAD.n2900 VSS 0.049115f
C3368 PAD.n2901 VSS 0.029436f
C3369 PAD.n2902 VSS 0.049115f
C3370 PAD.n2903 VSS 0.029436f
C3371 PAD.n2904 VSS 0.700534f
C3372 PAD.n2946 VSS 0.315733f
C3373 PAD.n2947 VSS 0.069765f
C3374 PAD.n2948 VSS 0.069765f
C3375 PAD.n2949 VSS 0.046286f
C3376 PAD.n2950 VSS 0.039761f
C3377 PAD.n2951 VSS 0.039761f
C3378 PAD.n2952 VSS 0.3552f
C3379 PAD.n2994 VSS 0.023109f
C3380 PAD.n2995 VSS 0.023109f
C3381 PAD.n2996 VSS 0.029436f
C3382 PAD.n2997 VSS 0.611735f
C3383 PAD.n2998 VSS 0.036461f
C3384 PAD.n2999 VSS 0.036461f
C3385 PAD.n3000 VSS 0.036461f
C3386 PAD.n3001 VSS 0.036461f
C3387 PAD.n3002 VSS 0.036461f
C3388 PAD.n3003 VSS 0.036461f
C3389 PAD.n3004 VSS 0.036461f
C3390 PAD.n3005 VSS 0.036461f
C3391 PAD.n3006 VSS 0.036461f
C3392 PAD.n3007 VSS 0.036461f
C3393 PAD.n3008 VSS 0.036461f
C3394 PAD.n3009 VSS 0.036461f
C3395 PAD.n3010 VSS 0.036461f
C3396 PAD.n3011 VSS 0.036461f
C3397 PAD.n3012 VSS 0.036461f
C3398 PAD.n3013 VSS 0.036461f
C3399 PAD.n3014 VSS 0.036461f
C3400 PAD.n3015 VSS 0.036461f
C3401 PAD.n3016 VSS 0.036461f
C3402 PAD.n3017 VSS 0.036461f
C3403 PAD.n3018 VSS 0.036461f
C3404 PAD.n3019 VSS 0.036461f
C3405 PAD.n3020 VSS 0.036461f
C3406 PAD.n3021 VSS 0.036461f
C3407 PAD.n3022 VSS 0.036461f
C3408 PAD.n3023 VSS 0.036461f
C3409 PAD.n3024 VSS 0.036461f
C3410 PAD.n3025 VSS 0.036461f
C3411 PAD.n3026 VSS 0.036461f
C3412 PAD.n3027 VSS 0.036461f
C3413 PAD.n3028 VSS 0.036461f
C3414 PAD.n3029 VSS 0.036461f
C3415 PAD.n3030 VSS 0.036461f
C3416 PAD.n3031 VSS 0.036461f
C3417 PAD.n3032 VSS 0.036461f
C3418 PAD.n3033 VSS 0.036461f
C3419 PAD.n3034 VSS 0.036461f
C3420 PAD.n3035 VSS 0.036461f
C3421 PAD.n3036 VSS 0.036461f
C3422 PAD.n3037 VSS 0.036461f
C3423 PAD.n3039 VSS 0.036461f
C3424 PAD.n3040 VSS 0.036461f
C3425 PAD.n3041 VSS 0.023109f
C3426 PAD.n3042 VSS 0.03338f
C3427 PAD.n3043 VSS 0.036461f
C3428 PAD.n3044 VSS 0.036461f
C3429 PAD.n3045 VSS 0.036461f
C3430 PAD.n3046 VSS 0.036461f
C3431 PAD.n3048 VSS 0.036461f
C3432 PAD.n3049 VSS 0.036461f
C3433 PAD.n3050 VSS 0.036461f
C3434 PAD.n3052 VSS 0.036461f
C3435 PAD.n3053 VSS 0.036461f
C3436 PAD.n3054 VSS 0.036461f
C3437 PAD.n3055 VSS 0.036461f
C3438 PAD.n3056 VSS 0.036461f
C3439 PAD.n3057 VSS 0.036461f
C3440 PAD.n3058 VSS 0.036461f
C3441 PAD.n3060 VSS 0.036461f
C3442 PAD.n3061 VSS 0.036461f
C3443 PAD.n3062 VSS 0.036461f
C3444 PAD.n3064 VSS 0.036461f
C3445 PAD.n3065 VSS 0.036461f
C3446 PAD.n3066 VSS 0.036461f
C3447 PAD.n3067 VSS 0.036461f
C3448 PAD.n3068 VSS 0.036461f
C3449 PAD.n3069 VSS 0.036461f
C3450 PAD.n3070 VSS 0.036461f
C3451 PAD.n3072 VSS 0.036461f
C3452 PAD.n3073 VSS 0.036461f
C3453 PAD.n3074 VSS 0.036461f
C3454 PAD.n3076 VSS 0.036461f
C3455 PAD.n3077 VSS 0.036461f
C3456 PAD.n3078 VSS 0.036461f
C3457 PAD.n3079 VSS 0.036461f
C3458 PAD.n3080 VSS 0.036461f
C3459 PAD.n3081 VSS 0.036461f
C3460 PAD.n3082 VSS 0.036461f
C3461 PAD.n3084 VSS 0.036461f
C3462 PAD.n3085 VSS 0.036461f
C3463 PAD.n3086 VSS 0.036461f
C3464 PAD.n3088 VSS 0.036461f
C3465 PAD.n3089 VSS 0.036461f
C3466 PAD.n3090 VSS 0.036461f
C3467 PAD.n3091 VSS 0.036461f
C3468 PAD.n3092 VSS 0.036461f
C3469 PAD.n3093 VSS 0.036461f
C3470 PAD.n3094 VSS 0.036461f
C3471 PAD.n3096 VSS 0.036461f
C3472 PAD.n3097 VSS 0.036461f
C3473 PAD.n3098 VSS 0.036461f
C3474 PAD.n3100 VSS 0.036461f
C3475 PAD.n3101 VSS 0.036461f
C3476 PAD.n3102 VSS 0.036461f
C3477 PAD.n3103 VSS 0.036461f
C3478 PAD.n3104 VSS 0.036461f
C3479 PAD.n3105 VSS 0.036461f
C3480 PAD.n3106 VSS 0.036461f
C3481 PAD.n3108 VSS 0.036461f
C3482 PAD.n3109 VSS 0.036461f
C3483 PAD.n3110 VSS 0.036461f
C3484 PAD.n3112 VSS 0.036461f
C3485 PAD.n3113 VSS 0.036461f
C3486 PAD.n3114 VSS 0.036461f
C3487 PAD.n3115 VSS 0.036461f
C3488 PAD.n3116 VSS 0.036461f
C3489 PAD.n3117 VSS 0.036461f
C3490 PAD.n3118 VSS 0.036461f
C3491 PAD.n3120 VSS 0.036461f
C3492 PAD.n3121 VSS 0.036461f
C3493 PAD.n3122 VSS 0.036461f
C3494 PAD.n3124 VSS 0.036461f
C3495 PAD.n3125 VSS 0.036461f
C3496 PAD.n3126 VSS 0.036461f
C3497 PAD.n3127 VSS 0.036461f
C3498 PAD.n3128 VSS 0.036461f
C3499 PAD.n3129 VSS 0.036461f
C3500 PAD.n3130 VSS 0.036461f
C3501 PAD.n3132 VSS 0.036461f
C3502 PAD.n3133 VSS 0.036461f
C3503 PAD.n3134 VSS 0.036461f
C3504 PAD.n3136 VSS 0.036461f
C3505 PAD.n3137 VSS 0.036461f
C3506 PAD.n3138 VSS 0.036461f
C3507 PAD.n3139 VSS 0.036461f
C3508 PAD.n3140 VSS 0.036461f
C3509 PAD.n3141 VSS 0.036461f
C3510 PAD.n3142 VSS 0.036461f
C3511 PAD.n3144 VSS 0.036461f
C3512 PAD.n3145 VSS 0.036461f
C3513 PAD.n3146 VSS 0.036461f
C3514 PAD.n3148 VSS 0.036461f
C3515 PAD.n3149 VSS 0.036461f
C3516 PAD.n3150 VSS 0.036461f
C3517 PAD.n3151 VSS 0.036461f
C3518 PAD.n3152 VSS 0.036461f
C3519 PAD.n3153 VSS 0.036461f
C3520 PAD.n3154 VSS 0.036461f
C3521 PAD.n3156 VSS 0.036461f
C3522 PAD.n3157 VSS 0.036461f
C3523 PAD.n3158 VSS 0.036461f
C3524 PAD.n3160 VSS 0.036461f
C3525 PAD.n3161 VSS 0.036461f
C3526 PAD.n3162 VSS 0.036461f
C3527 PAD.n3163 VSS 0.036461f
C3528 PAD.n3164 VSS 0.036461f
C3529 PAD.n3165 VSS 0.036461f
C3530 PAD.n3166 VSS 0.036461f
C3531 PAD.n3168 VSS 0.036461f
C3532 PAD.n3169 VSS 0.036461f
C3533 PAD.n3170 VSS 0.036461f
C3534 PAD.n3172 VSS 0.036461f
C3535 PAD.n3173 VSS 0.036461f
C3536 PAD.n3174 VSS 0.036461f
C3537 PAD.n3175 VSS 0.036461f
C3538 PAD.n3176 VSS 0.036461f
C3539 PAD.n3177 VSS 0.036461f
C3540 PAD.n3178 VSS 0.036461f
C3541 PAD.n3180 VSS 0.036461f
C3542 PAD.n3181 VSS 0.036461f
C3543 PAD.n3182 VSS 0.036461f
C3544 PAD.n3184 VSS 0.036461f
C3545 PAD.n3185 VSS 0.036461f
C3546 PAD.n3186 VSS 0.036461f
C3547 PAD.n3187 VSS 0.036461f
C3548 PAD.n3188 VSS 0.036461f
C3549 PAD.n3189 VSS 0.036461f
C3550 PAD.n3190 VSS 0.036461f
C3551 PAD.n3192 VSS 0.036461f
C3552 PAD.n3193 VSS 0.036461f
C3553 PAD.n3194 VSS 0.036461f
C3554 PAD.n3196 VSS 0.036461f
C3555 PAD.n3197 VSS 0.036461f
C3556 PAD.n3198 VSS 0.036461f
C3557 PAD.n3199 VSS 0.036461f
C3558 PAD.n3200 VSS 0.036461f
C3559 PAD.n3201 VSS 0.036461f
C3560 PAD.n3202 VSS 0.036461f
C3561 PAD.n3204 VSS 0.036461f
C3562 PAD.n3205 VSS 0.036461f
C3563 PAD.n3206 VSS 0.036461f
C3564 PAD.n3208 VSS 0.036461f
C3565 PAD.n3209 VSS 0.036461f
C3566 PAD.n3210 VSS 0.036461f
C3567 PAD.n3211 VSS 0.036461f
C3568 PAD.n3212 VSS 0.036461f
C3569 PAD.n3213 VSS 0.036461f
C3570 PAD.n3214 VSS 0.036461f
C3571 PAD.n3216 VSS 0.036461f
C3572 PAD.n3217 VSS 0.036461f
C3573 PAD.n3218 VSS 0.036461f
C3574 PAD.n3220 VSS 0.036461f
C3575 PAD.n3221 VSS 0.036461f
C3576 PAD.n3222 VSS 0.036461f
C3577 PAD.n3223 VSS 0.036461f
C3578 PAD.n3224 VSS 0.036461f
C3579 PAD.n3225 VSS 0.036461f
C3580 PAD.n3226 VSS 0.036461f
C3581 PAD.n3228 VSS 0.036461f
C3582 PAD.n3229 VSS 0.036461f
C3583 PAD.n3230 VSS 0.036461f
C3584 PAD.n3232 VSS 0.036461f
C3585 PAD.n3233 VSS 0.036461f
C3586 PAD.n3234 VSS 0.036461f
C3587 PAD.n3235 VSS 0.036461f
C3588 PAD.n3236 VSS 0.036461f
C3589 PAD.n3237 VSS 0.036461f
C3590 PAD.n3238 VSS 0.036461f
C3591 PAD.n3240 VSS 0.036461f
C3592 PAD.n3241 VSS 0.036461f
C3593 PAD.n3242 VSS 0.036461f
C3594 PAD.n3244 VSS 0.036461f
C3595 PAD.n3245 VSS 0.036461f
C3596 PAD.n3246 VSS 0.036461f
C3597 PAD.n3247 VSS 0.036461f
C3598 PAD.n3248 VSS 0.036461f
C3599 PAD.n3249 VSS 0.036461f
C3600 PAD.n3250 VSS 0.036461f
C3601 PAD.n3252 VSS 0.036461f
C3602 PAD.n3253 VSS 0.036461f
C3603 PAD.n3254 VSS 0.036461f
C3604 PAD.n3256 VSS 0.036461f
C3605 PAD.n3257 VSS 0.036461f
C3606 PAD.n3258 VSS 0.036461f
C3607 PAD.n3259 VSS 0.036461f
C3608 PAD.n3260 VSS 0.036461f
C3609 PAD.n3261 VSS 0.036461f
C3610 PAD.n3262 VSS 0.036461f
C3611 PAD.n3264 VSS 0.036461f
C3612 PAD.n3265 VSS 0.036461f
C3613 PAD.n3266 VSS 0.036461f
C3614 PAD.n3268 VSS 0.036461f
C3615 PAD.n3269 VSS 0.036461f
C3616 PAD.n3270 VSS 0.036461f
C3617 PAD.n3271 VSS 0.036461f
C3618 PAD.n3272 VSS 0.036461f
C3619 PAD.n3273 VSS 0.036461f
C3620 PAD.n3274 VSS 0.036461f
C3621 PAD.n3276 VSS 0.036461f
C3622 PAD.n3277 VSS 0.036461f
C3623 PAD.n3278 VSS 0.036461f
C3624 PAD.n3280 VSS 0.036461f
C3625 PAD.n3281 VSS 0.036461f
C3626 PAD.n3282 VSS 0.036461f
C3627 PAD.n3283 VSS 0.036461f
C3628 PAD.n3284 VSS 0.04214f
C3629 PAD.n3285 VSS 0.045483f
C3630 PAD.n3286 VSS 0.045483f
C3631 PAD.n3287 VSS 0.700534f
C3632 PAD.n3288 VSS 0.069765f
C3633 PAD.n3289 VSS 0.389734f
C3634 PAD.n3290 VSS 0.036008f
C3635 PAD.n3291 VSS 0.069765f
C3636 PAD.n3292 VSS 0.036008f
C3637 PAD.n3293 VSS 0.046286f
C3638 PAD.n3294 VSS 0.039761f
C3639 PAD.n3295 VSS 0.039761f
C3640 PAD.n3296 VSS 0.498267f
C3641 PAD.n3338 VSS 0.023109f
C3642 PAD.n3339 VSS 0.409467f
C3643 PAD.n3340 VSS 0.023109f
C3644 PAD.n3341 VSS 0.029436f
C3645 PAD.n3342 VSS 0.389734f
C3646 PAD.n3343 VSS 0.036461f
C3647 PAD.n3344 VSS 0.036461f
C3648 PAD.n3345 VSS 0.036461f
C3649 PAD.n3346 VSS 0.036461f
C3650 PAD.n3347 VSS 0.036461f
C3651 PAD.n3348 VSS 0.036461f
C3652 PAD.n3349 VSS 0.036461f
C3653 PAD.n3350 VSS 0.036461f
C3654 PAD.n3351 VSS 0.036461f
C3655 PAD.n3352 VSS 0.036461f
C3656 PAD.n3353 VSS 0.036461f
C3657 PAD.n3354 VSS 0.036461f
C3658 PAD.n3355 VSS 0.036461f
C3659 PAD.n3356 VSS 0.036461f
C3660 PAD.n3357 VSS 0.036461f
C3661 PAD.n3358 VSS 0.036461f
C3662 PAD.n3359 VSS 0.036461f
C3663 PAD.n3360 VSS 0.036461f
C3664 PAD.n3361 VSS 0.036461f
C3665 PAD.n3362 VSS 0.036461f
C3666 PAD.n3363 VSS 0.036461f
C3667 PAD.n3364 VSS 0.036461f
C3668 PAD.n3365 VSS 0.036461f
C3669 PAD.n3366 VSS 0.036461f
C3670 PAD.n3367 VSS 0.036461f
C3671 PAD.n3368 VSS 0.036461f
C3672 PAD.n3369 VSS 0.036461f
C3673 PAD.n3370 VSS 0.036461f
C3674 PAD.n3371 VSS 0.036461f
C3675 PAD.n3372 VSS 0.036461f
C3676 PAD.n3373 VSS 0.036461f
C3677 PAD.n3374 VSS 0.036461f
C3678 PAD.n3375 VSS 0.036461f
C3679 PAD.n3376 VSS 0.036461f
C3680 PAD.n3377 VSS 0.036461f
C3681 PAD.n3378 VSS 0.036461f
C3682 PAD.n3379 VSS 0.036461f
C3683 PAD.n3380 VSS 0.036461f
C3684 PAD.n3381 VSS 0.036461f
C3685 PAD.n3382 VSS 0.036461f
C3686 PAD.n3384 VSS 0.036461f
C3687 PAD.n3385 VSS 0.036461f
C3688 PAD.n3386 VSS 0.023109f
C3689 PAD.n3387 VSS 0.03338f
C3690 PAD.n3388 VSS 0.036461f
C3691 PAD.n3389 VSS 0.036461f
C3692 PAD.n3390 VSS 0.036461f
C3693 PAD.n3391 VSS 0.036461f
C3694 PAD.n3393 VSS 0.036461f
C3695 PAD.n3394 VSS 0.036461f
C3696 PAD.n3395 VSS 0.036461f
C3697 PAD.n3397 VSS 0.036461f
C3698 PAD.n3398 VSS 0.036461f
C3699 PAD.n3399 VSS 0.036461f
C3700 PAD.n3400 VSS 0.036461f
C3701 PAD.n3401 VSS 0.036461f
C3702 PAD.n3402 VSS 0.036461f
C3703 PAD.n3403 VSS 0.036461f
C3704 PAD.n3405 VSS 0.036461f
C3705 PAD.n3406 VSS 0.036461f
C3706 PAD.n3407 VSS 0.036461f
C3707 PAD.n3409 VSS 0.036461f
C3708 PAD.n3410 VSS 0.036461f
C3709 PAD.n3411 VSS 0.036461f
C3710 PAD.n3412 VSS 0.036461f
C3711 PAD.n3413 VSS 0.036461f
C3712 PAD.n3414 VSS 0.036461f
C3713 PAD.n3415 VSS 0.036461f
C3714 PAD.n3417 VSS 0.036461f
C3715 PAD.n3418 VSS 0.036461f
C3716 PAD.n3419 VSS 0.036461f
C3717 PAD.n3421 VSS 0.036461f
C3718 PAD.n3422 VSS 0.036461f
C3719 PAD.n3423 VSS 0.036461f
C3720 PAD.n3424 VSS 0.036461f
C3721 PAD.n3425 VSS 0.036461f
C3722 PAD.n3426 VSS 0.036461f
C3723 PAD.n3427 VSS 0.036461f
C3724 PAD.n3429 VSS 0.036461f
C3725 PAD.n3430 VSS 0.036461f
C3726 PAD.n3431 VSS 0.036461f
C3727 PAD.n3433 VSS 0.036461f
C3728 PAD.n3434 VSS 0.036461f
C3729 PAD.n3435 VSS 0.036461f
C3730 PAD.n3436 VSS 0.036461f
C3731 PAD.n3437 VSS 0.036461f
C3732 PAD.n3438 VSS 0.036461f
C3733 PAD.n3439 VSS 0.036461f
C3734 PAD.n3441 VSS 0.036461f
C3735 PAD.n3442 VSS 0.036461f
C3736 PAD.n3443 VSS 0.036461f
C3737 PAD.n3445 VSS 0.036461f
C3738 PAD.n3446 VSS 0.036461f
C3739 PAD.n3447 VSS 0.036461f
C3740 PAD.n3448 VSS 0.036461f
C3741 PAD.n3449 VSS 0.036461f
C3742 PAD.n3450 VSS 0.036461f
C3743 PAD.n3451 VSS 0.036461f
C3744 PAD.n3453 VSS 0.036461f
C3745 PAD.n3454 VSS 0.036461f
C3746 PAD.n3455 VSS 0.036461f
C3747 PAD.n3457 VSS 0.036461f
C3748 PAD.n3458 VSS 0.036461f
C3749 PAD.n3459 VSS 0.036461f
C3750 PAD.n3460 VSS 0.036461f
C3751 PAD.n3461 VSS 0.036461f
C3752 PAD.n3462 VSS 0.036461f
C3753 PAD.n3463 VSS 0.036461f
C3754 PAD.n3465 VSS 0.036461f
C3755 PAD.n3466 VSS 0.036461f
C3756 PAD.n3467 VSS 0.036461f
C3757 PAD.n3469 VSS 0.036461f
C3758 PAD.n3470 VSS 0.036461f
C3759 PAD.n3471 VSS 0.036461f
C3760 PAD.n3472 VSS 0.036461f
C3761 PAD.n3473 VSS 0.036461f
C3762 PAD.n3474 VSS 0.036461f
C3763 PAD.n3475 VSS 0.036461f
C3764 PAD.n3477 VSS 0.036461f
C3765 PAD.n3478 VSS 0.036461f
C3766 PAD.n3479 VSS 0.036461f
C3767 PAD.n3481 VSS 0.036461f
C3768 PAD.n3482 VSS 0.036461f
C3769 PAD.n3483 VSS 0.036461f
C3770 PAD.n3484 VSS 0.036461f
C3771 PAD.n3485 VSS 0.036461f
C3772 PAD.n3486 VSS 0.036461f
C3773 PAD.n3487 VSS 0.036461f
C3774 PAD.n3489 VSS 0.036461f
C3775 PAD.n3490 VSS 0.036461f
C3776 PAD.n3491 VSS 0.036461f
C3777 PAD.n3493 VSS 0.036461f
C3778 PAD.n3494 VSS 0.036461f
C3779 PAD.n3495 VSS 0.036461f
C3780 PAD.n3496 VSS 0.036461f
C3781 PAD.n3497 VSS 0.036461f
C3782 PAD.n3498 VSS 0.036461f
C3783 PAD.n3499 VSS 0.036461f
C3784 PAD.n3501 VSS 0.036461f
C3785 PAD.n3502 VSS 0.036461f
C3786 PAD.n3503 VSS 0.036461f
C3787 PAD.n3505 VSS 0.036461f
C3788 PAD.n3506 VSS 0.036461f
C3789 PAD.n3507 VSS 0.036461f
C3790 PAD.n3508 VSS 0.036461f
C3791 PAD.n3509 VSS 0.036461f
C3792 PAD.n3510 VSS 0.036461f
C3793 PAD.n3511 VSS 0.036461f
C3794 PAD.n3513 VSS 0.036461f
C3795 PAD.n3514 VSS 0.036461f
C3796 PAD.n3515 VSS 0.036461f
C3797 PAD.n3517 VSS 0.036461f
C3798 PAD.n3518 VSS 0.036461f
C3799 PAD.n3519 VSS 0.036461f
C3800 PAD.n3520 VSS 0.036461f
C3801 PAD.n3521 VSS 0.036461f
C3802 PAD.n3522 VSS 0.036461f
C3803 PAD.n3523 VSS 0.036461f
C3804 PAD.n3525 VSS 0.036461f
C3805 PAD.n3526 VSS 0.036461f
C3806 PAD.n3527 VSS 0.036461f
C3807 PAD.n3529 VSS 0.036461f
C3808 PAD.n3530 VSS 0.036461f
C3809 PAD.n3531 VSS 0.036461f
C3810 PAD.n3532 VSS 0.036461f
C3811 PAD.n3533 VSS 0.036461f
C3812 PAD.n3534 VSS 0.036461f
C3813 PAD.n3535 VSS 0.036461f
C3814 PAD.n3537 VSS 0.036461f
C3815 PAD.n3538 VSS 0.036461f
C3816 PAD.n3539 VSS 0.036461f
C3817 PAD.n3541 VSS 0.036461f
C3818 PAD.n3542 VSS 0.036461f
C3819 PAD.n3543 VSS 0.036461f
C3820 PAD.n3544 VSS 0.036461f
C3821 PAD.n3545 VSS 0.036461f
C3822 PAD.n3546 VSS 0.036461f
C3823 PAD.n3547 VSS 0.036461f
C3824 PAD.n3549 VSS 0.036461f
C3825 PAD.n3550 VSS 0.036461f
C3826 PAD.n3551 VSS 0.036461f
C3827 PAD.n3553 VSS 0.036461f
C3828 PAD.n3554 VSS 0.036461f
C3829 PAD.n3555 VSS 0.036461f
C3830 PAD.n3556 VSS 0.036461f
C3831 PAD.n3557 VSS 0.036461f
C3832 PAD.n3558 VSS 0.036461f
C3833 PAD.n3559 VSS 0.036461f
C3834 PAD.n3561 VSS 0.036461f
C3835 PAD.n3562 VSS 0.036461f
C3836 PAD.n3563 VSS 0.036461f
C3837 PAD.n3565 VSS 0.036461f
C3838 PAD.n3566 VSS 0.036461f
C3839 PAD.n3567 VSS 0.036461f
C3840 PAD.n3568 VSS 0.036461f
C3841 PAD.n3569 VSS 0.036461f
C3842 PAD.n3570 VSS 0.036461f
C3843 PAD.n3571 VSS 0.036461f
C3844 PAD.n3573 VSS 0.036461f
C3845 PAD.n3574 VSS 0.036461f
C3846 PAD.n3575 VSS 0.036461f
C3847 PAD.n3577 VSS 0.036461f
C3848 PAD.n3578 VSS 0.036461f
C3849 PAD.n3579 VSS 0.036461f
C3850 PAD.n3580 VSS 0.036461f
C3851 PAD.n3581 VSS 0.036461f
C3852 PAD.n3582 VSS 0.036461f
C3853 PAD.n3583 VSS 0.036461f
C3854 PAD.n3585 VSS 0.036461f
C3855 PAD.n3586 VSS 0.036461f
C3856 PAD.n3587 VSS 0.036461f
C3857 PAD.n3589 VSS 0.036461f
C3858 PAD.n3590 VSS 0.036461f
C3859 PAD.n3591 VSS 0.036461f
C3860 PAD.n3592 VSS 0.036461f
C3861 PAD.n3593 VSS 0.036461f
C3862 PAD.n3594 VSS 0.036461f
C3863 PAD.n3595 VSS 0.036461f
C3864 PAD.n3597 VSS 0.036461f
C3865 PAD.n3598 VSS 0.036461f
C3866 PAD.n3599 VSS 0.036461f
C3867 PAD.n3601 VSS 0.036461f
C3868 PAD.n3602 VSS 0.036461f
C3869 PAD.n3603 VSS 0.036461f
C3870 PAD.n3604 VSS 0.036461f
C3871 PAD.n3605 VSS 0.036461f
C3872 PAD.n3606 VSS 0.036461f
C3873 PAD.n3607 VSS 0.036461f
C3874 PAD.n3609 VSS 0.036461f
C3875 PAD.n3610 VSS 0.036461f
C3876 PAD.n3611 VSS 0.036461f
C3877 PAD.n3613 VSS 0.036461f
C3878 PAD.n3614 VSS 0.036461f
C3879 PAD.n3615 VSS 0.036461f
C3880 PAD.n3616 VSS 0.036461f
C3881 PAD.n3617 VSS 0.036461f
C3882 PAD.n3618 VSS 0.036461f
C3883 PAD.n3619 VSS 0.036461f
C3884 PAD.n3621 VSS 0.036461f
C3885 PAD.n3622 VSS 0.036461f
C3886 PAD.n3623 VSS 0.036461f
C3887 PAD.n3625 VSS 0.036461f
C3888 PAD.n3626 VSS 0.036461f
C3889 PAD.n3627 VSS 0.036461f
C3890 PAD.n3628 VSS 0.036461f
C3891 PAD.n3629 VSS 0.042895f
C3892 PAD.n3630 VSS 0.049115f
C3893 PAD.n3631 VSS 0.029436f
C3894 PAD.n3632 VSS 0.040987f
C3895 PAD.n3633 VSS 0.700534f
C3896 PAD.n3634 VSS 0.069765f
C3897 PAD.n3635 VSS 0.069765f
C3898 PAD.n3636 VSS 12.709f
C3899 PAD.n3637 VSS 14.5471f
C3900 PAD.n3638 VSS 0.046286f
C3901 PAD.n3639 VSS 0.039761f
C3902 PAD.n3640 VSS 0.039761f
C3903 PAD.n3641 VSS 0.606801f
C3904 PAD.n3683 VSS 0.023109f
C3905 PAD.n3684 VSS 0.518001f
C3906 PAD.n3685 VSS 0.023109f
C3907 PAD.n3686 VSS 0.029436f
C3908 PAD.n3687 VSS 0.123333f
C3909 PAD.n3688 VSS 0.036461f
C3910 PAD.n3689 VSS 0.036461f
C3911 PAD.n3690 VSS 0.036461f
C3912 PAD.n3691 VSS 0.036461f
C3913 PAD.n3692 VSS 0.036461f
C3914 PAD.n3693 VSS 0.036461f
C3915 PAD.n3694 VSS 0.036461f
C3916 PAD.n3695 VSS 0.036461f
C3917 PAD.n3696 VSS 0.036461f
C3918 PAD.n3697 VSS 0.036461f
C3919 PAD.n3698 VSS 0.036461f
C3920 PAD.n3699 VSS 0.036461f
C3921 PAD.n3700 VSS 0.036461f
C3922 PAD.n3701 VSS 0.036461f
C3923 PAD.n3702 VSS 0.036461f
C3924 PAD.n3703 VSS 0.036461f
C3925 PAD.n3704 VSS 0.036461f
C3926 PAD.n3705 VSS 0.036461f
C3927 PAD.n3706 VSS 0.036461f
C3928 PAD.n3707 VSS 0.036461f
C3929 PAD.n3708 VSS 0.036461f
C3930 PAD.n3709 VSS 0.036461f
C3931 PAD.n3710 VSS 0.036461f
C3932 PAD.n3711 VSS 0.036461f
C3933 PAD.n3712 VSS 0.036461f
C3934 PAD.n3713 VSS 0.036461f
C3935 PAD.n3714 VSS 0.036461f
C3936 PAD.n3715 VSS 0.036461f
C3937 PAD.n3716 VSS 0.036461f
C3938 PAD.n3717 VSS 0.036461f
C3939 PAD.n3718 VSS 0.036461f
C3940 PAD.n3719 VSS 0.036461f
C3941 PAD.n3720 VSS 0.036461f
C3942 PAD.n3721 VSS 0.036461f
C3943 PAD.n3722 VSS 0.036461f
C3944 PAD.n3723 VSS 0.036461f
C3945 PAD.n3724 VSS 0.036461f
C3946 PAD.n3725 VSS 0.036461f
C3947 PAD.n3726 VSS 0.036461f
C3948 PAD.n3727 VSS 0.036461f
C3949 PAD.n3729 VSS 0.036461f
C3950 PAD.n3730 VSS 0.036461f
C3951 PAD.n3731 VSS 0.023109f
C3952 PAD.n3732 VSS 0.03338f
C3953 PAD.n3733 VSS 0.036461f
C3954 PAD.n3734 VSS 0.036461f
C3955 PAD.n3735 VSS 0.036461f
C3956 PAD.n3736 VSS 0.036461f
C3957 PAD.n3738 VSS 0.036461f
C3958 PAD.n3739 VSS 0.036461f
C3959 PAD.n3740 VSS 0.036461f
C3960 PAD.n3742 VSS 0.036461f
C3961 PAD.n3743 VSS 0.036461f
C3962 PAD.n3744 VSS 0.036461f
C3963 PAD.n3745 VSS 0.036461f
C3964 PAD.n3746 VSS 0.036461f
C3965 PAD.n3747 VSS 0.036461f
C3966 PAD.n3748 VSS 0.036461f
C3967 PAD.n3750 VSS 0.036461f
C3968 PAD.n3751 VSS 0.036461f
C3969 PAD.n3752 VSS 0.036461f
C3970 PAD.n3754 VSS 0.036461f
C3971 PAD.n3755 VSS 0.036461f
C3972 PAD.n3756 VSS 0.036461f
C3973 PAD.n3757 VSS 0.036461f
C3974 PAD.n3758 VSS 0.036461f
C3975 PAD.n3759 VSS 0.036461f
C3976 PAD.n3760 VSS 0.036461f
C3977 PAD.n3762 VSS 0.036461f
C3978 PAD.n3763 VSS 0.036461f
C3979 PAD.n3764 VSS 0.036461f
C3980 PAD.n3766 VSS 0.036461f
C3981 PAD.n3767 VSS 0.036461f
C3982 PAD.n3768 VSS 0.036461f
C3983 PAD.n3769 VSS 0.036461f
C3984 PAD.n3770 VSS 0.036461f
C3985 PAD.n3771 VSS 0.036461f
C3986 PAD.n3772 VSS 0.036461f
C3987 PAD.n3774 VSS 0.036461f
C3988 PAD.n3775 VSS 0.036461f
C3989 PAD.n3776 VSS 0.036461f
C3990 PAD.n3778 VSS 0.036461f
C3991 PAD.n3779 VSS 0.036461f
C3992 PAD.n3780 VSS 0.036461f
C3993 PAD.n3781 VSS 0.036461f
C3994 PAD.n3782 VSS 0.036461f
C3995 PAD.n3783 VSS 0.036461f
C3996 PAD.n3784 VSS 0.036461f
C3997 PAD.n3786 VSS 0.036461f
C3998 PAD.n3787 VSS 0.036461f
C3999 PAD.n3788 VSS 0.036461f
C4000 PAD.n3790 VSS 0.036461f
C4001 PAD.n3791 VSS 0.036461f
C4002 PAD.n3792 VSS 0.036461f
C4003 PAD.n3793 VSS 0.036461f
C4004 PAD.n3794 VSS 0.036461f
C4005 PAD.n3795 VSS 0.036461f
C4006 PAD.n3796 VSS 0.036461f
C4007 PAD.n3798 VSS 0.036461f
C4008 PAD.n3799 VSS 0.036461f
C4009 PAD.n3800 VSS 0.036461f
C4010 PAD.n3802 VSS 0.036461f
C4011 PAD.n3803 VSS 0.036461f
C4012 PAD.n3804 VSS 0.036461f
C4013 PAD.n3805 VSS 0.036461f
C4014 PAD.n3806 VSS 0.036461f
C4015 PAD.n3807 VSS 0.036461f
C4016 PAD.n3808 VSS 0.036461f
C4017 PAD.n3810 VSS 0.036461f
C4018 PAD.n3811 VSS 0.036461f
C4019 PAD.n3812 VSS 0.036461f
C4020 PAD.n3814 VSS 0.036461f
C4021 PAD.n3815 VSS 0.036461f
C4022 PAD.n3816 VSS 0.036461f
C4023 PAD.n3817 VSS 0.036461f
C4024 PAD.n3818 VSS 0.036461f
C4025 PAD.n3819 VSS 0.036461f
C4026 PAD.n3820 VSS 0.036461f
C4027 PAD.n3822 VSS 0.036461f
C4028 PAD.n3823 VSS 0.036461f
C4029 PAD.n3824 VSS 0.036461f
C4030 PAD.n3826 VSS 0.036461f
C4031 PAD.n3827 VSS 0.036461f
C4032 PAD.n3828 VSS 0.036461f
C4033 PAD.n3829 VSS 0.036461f
C4034 PAD.n3830 VSS 0.036461f
C4035 PAD.n3831 VSS 0.036461f
C4036 PAD.n3832 VSS 0.036461f
C4037 PAD.n3834 VSS 0.036461f
C4038 PAD.n3835 VSS 0.036461f
C4039 PAD.n3836 VSS 0.036461f
C4040 PAD.n3838 VSS 0.036461f
C4041 PAD.n3839 VSS 0.036461f
C4042 PAD.n3840 VSS 0.036461f
C4043 PAD.n3841 VSS 0.036461f
C4044 PAD.n3842 VSS 0.036461f
C4045 PAD.n3843 VSS 0.036461f
C4046 PAD.n3844 VSS 0.036461f
C4047 PAD.n3846 VSS 0.036461f
C4048 PAD.n3847 VSS 0.036461f
C4049 PAD.n3848 VSS 0.036461f
C4050 PAD.n3850 VSS 0.036461f
C4051 PAD.n3851 VSS 0.036461f
C4052 PAD.n3852 VSS 0.036461f
C4053 PAD.n3853 VSS 0.036461f
C4054 PAD.n3854 VSS 0.036461f
C4055 PAD.n3855 VSS 0.036461f
C4056 PAD.n3856 VSS 0.036461f
C4057 PAD.n3858 VSS 0.036461f
C4058 PAD.n3859 VSS 0.036461f
C4059 PAD.n3860 VSS 0.036461f
C4060 PAD.n3862 VSS 0.036461f
C4061 PAD.n3863 VSS 0.036461f
C4062 PAD.n3864 VSS 0.036461f
C4063 PAD.n3865 VSS 0.036461f
C4064 PAD.n3866 VSS 0.036461f
C4065 PAD.n3867 VSS 0.036461f
C4066 PAD.n3868 VSS 0.036461f
C4067 PAD.n3870 VSS 0.036461f
C4068 PAD.n3871 VSS 0.036461f
C4069 PAD.n3872 VSS 0.036461f
C4070 PAD.n3874 VSS 0.036461f
C4071 PAD.n3875 VSS 0.036461f
C4072 PAD.n3876 VSS 0.036461f
C4073 PAD.n3877 VSS 0.036461f
C4074 PAD.n3878 VSS 0.036461f
C4075 PAD.n3879 VSS 0.036461f
C4076 PAD.n3880 VSS 0.036461f
C4077 PAD.n3882 VSS 0.036461f
C4078 PAD.n3883 VSS 0.036461f
C4079 PAD.n3884 VSS 0.036461f
C4080 PAD.n3886 VSS 0.036461f
C4081 PAD.n3887 VSS 0.036461f
C4082 PAD.n3888 VSS 0.036461f
C4083 PAD.n3889 VSS 0.036461f
C4084 PAD.n3890 VSS 0.036461f
C4085 PAD.n3891 VSS 0.036461f
C4086 PAD.n3892 VSS 0.036461f
C4087 PAD.n3894 VSS 0.036461f
C4088 PAD.n3895 VSS 0.036461f
C4089 PAD.n3896 VSS 0.036461f
C4090 PAD.n3898 VSS 0.036461f
C4091 PAD.n3899 VSS 0.036461f
C4092 PAD.n3900 VSS 0.036461f
C4093 PAD.n3901 VSS 0.036461f
C4094 PAD.n3902 VSS 0.036461f
C4095 PAD.n3903 VSS 0.036461f
C4096 PAD.n3904 VSS 0.036461f
C4097 PAD.n3906 VSS 0.036461f
C4098 PAD.n3907 VSS 0.036461f
C4099 PAD.n3908 VSS 0.036461f
C4100 PAD.n3910 VSS 0.036461f
C4101 PAD.n3911 VSS 0.036461f
C4102 PAD.n3912 VSS 0.036461f
C4103 PAD.n3913 VSS 0.036461f
C4104 PAD.n3914 VSS 0.036461f
C4105 PAD.n3915 VSS 0.036461f
C4106 PAD.n3916 VSS 0.036461f
C4107 PAD.n3918 VSS 0.036461f
C4108 PAD.n3919 VSS 0.036461f
C4109 PAD.n3920 VSS 0.036461f
C4110 PAD.n3922 VSS 0.036461f
C4111 PAD.n3923 VSS 0.036461f
C4112 PAD.n3924 VSS 0.036461f
C4113 PAD.n3925 VSS 0.036461f
C4114 PAD.n3926 VSS 0.036461f
C4115 PAD.n3927 VSS 0.036461f
C4116 PAD.n3928 VSS 0.036461f
C4117 PAD.n3930 VSS 0.036461f
C4118 PAD.n3931 VSS 0.036461f
C4119 PAD.n3932 VSS 0.036461f
C4120 PAD.n3934 VSS 0.036461f
C4121 PAD.n3935 VSS 0.036461f
C4122 PAD.n3936 VSS 0.036461f
C4123 PAD.n3937 VSS 0.036461f
C4124 PAD.n3938 VSS 0.036461f
C4125 PAD.n3939 VSS 0.036461f
C4126 PAD.n3940 VSS 0.036461f
C4127 PAD.n3942 VSS 0.036461f
C4128 PAD.n3943 VSS 0.036461f
C4129 PAD.n3944 VSS 0.036461f
C4130 PAD.n3946 VSS 0.036461f
C4131 PAD.n3947 VSS 0.036461f
C4132 PAD.n3948 VSS 0.036461f
C4133 PAD.n3949 VSS 0.036461f
C4134 PAD.n3950 VSS 0.036461f
C4135 PAD.n3951 VSS 0.036461f
C4136 PAD.n3952 VSS 0.036461f
C4137 PAD.n3954 VSS 0.036461f
C4138 PAD.n3955 VSS 0.036461f
C4139 PAD.n3956 VSS 0.036461f
C4140 PAD.n3958 VSS 0.036461f
C4141 PAD.n3959 VSS 0.036461f
C4142 PAD.n3960 VSS 0.036461f
C4143 PAD.n3961 VSS 0.036461f
C4144 PAD.n3962 VSS 0.036461f
C4145 PAD.n3963 VSS 0.036461f
C4146 PAD.n3964 VSS 0.036461f
C4147 PAD.n3966 VSS 0.036461f
C4148 PAD.n3967 VSS 0.036461f
C4149 PAD.n3968 VSS 0.036461f
C4150 PAD.n3970 VSS 0.036461f
C4151 PAD.n3971 VSS 0.036461f
C4152 PAD.n3972 VSS 0.036461f
C4153 PAD.n3973 VSS 0.036461f
C4154 PAD.n3974 VSS 0.028547f
C4155 PAD.n3975 VSS 0.049115f
C4156 PAD.n3976 VSS 0.03649f
C4157 PAD.n3977 VSS 0.646268f
C4158 PAD.n3978 VSS 0.069765f
C4159 PAD.n3979 VSS 0.069765f
C4160 PAD.n3980 VSS 0.046286f
C4161 PAD.n3981 VSS 0.039761f
C4162 PAD.n3982 VSS 0.039761f
C4163 PAD.n3983 VSS 0.562401f
C4164 PAD.n4025 VSS 0.023109f
C4165 PAD.n4026 VSS 0.023109f
C4166 PAD.n4027 VSS 0.029436f
C4167 PAD.n4028 VSS 0.143067f
C4168 PAD.n4029 VSS 0.036461f
C4169 PAD.n4030 VSS 0.036461f
C4170 PAD.n4031 VSS 0.036461f
C4171 PAD.n4032 VSS 0.036461f
C4172 PAD.n4033 VSS 0.036461f
C4173 PAD.n4034 VSS 0.036461f
C4174 PAD.n4035 VSS 0.036461f
C4175 PAD.n4036 VSS 0.036461f
C4176 PAD.n4037 VSS 0.036461f
C4177 PAD.n4038 VSS 0.036461f
C4178 PAD.n4039 VSS 0.036461f
C4179 PAD.n4040 VSS 0.036461f
C4180 PAD.n4041 VSS 0.036461f
C4181 PAD.n4042 VSS 0.036461f
C4182 PAD.n4043 VSS 0.036461f
C4183 PAD.n4044 VSS 0.036461f
C4184 PAD.n4045 VSS 0.036461f
C4185 PAD.n4046 VSS 0.036461f
C4186 PAD.n4047 VSS 0.036461f
C4187 PAD.n4048 VSS 0.036461f
C4188 PAD.n4049 VSS 0.036461f
C4189 PAD.n4050 VSS 0.036461f
C4190 PAD.n4051 VSS 0.036461f
C4191 PAD.n4052 VSS 0.036461f
C4192 PAD.n4053 VSS 0.036461f
C4193 PAD.n4054 VSS 0.036461f
C4194 PAD.n4055 VSS 0.036461f
C4195 PAD.n4056 VSS 0.036461f
C4196 PAD.n4057 VSS 0.036461f
C4197 PAD.n4058 VSS 0.036461f
C4198 PAD.n4059 VSS 0.036461f
C4199 PAD.n4060 VSS 0.036461f
C4200 PAD.n4061 VSS 0.036461f
C4201 PAD.n4062 VSS 0.036461f
C4202 PAD.n4063 VSS 0.036461f
C4203 PAD.n4064 VSS 0.036461f
C4204 PAD.n4065 VSS 0.036461f
C4205 PAD.n4066 VSS 0.036461f
C4206 PAD.n4067 VSS 0.036461f
C4207 PAD.n4068 VSS 0.036461f
C4208 PAD.n4070 VSS 0.036461f
C4209 PAD.n4071 VSS 0.036461f
C4210 PAD.n4072 VSS 0.023109f
C4211 PAD.n4073 VSS 0.03338f
C4212 PAD.n4074 VSS 0.036461f
C4213 PAD.n4075 VSS 0.036461f
C4214 PAD.n4076 VSS 0.036461f
C4215 PAD.n4077 VSS 0.036461f
C4216 PAD.n4079 VSS 0.036461f
C4217 PAD.n4080 VSS 0.036461f
C4218 PAD.n4081 VSS 0.036461f
C4219 PAD.n4083 VSS 0.036461f
C4220 PAD.n4084 VSS 0.036461f
C4221 PAD.n4085 VSS 0.036461f
C4222 PAD.n4086 VSS 0.036461f
C4223 PAD.n4087 VSS 0.036461f
C4224 PAD.n4088 VSS 0.036461f
C4225 PAD.n4089 VSS 0.036461f
C4226 PAD.n4091 VSS 0.036461f
C4227 PAD.n4092 VSS 0.036461f
C4228 PAD.n4093 VSS 0.036461f
C4229 PAD.n4095 VSS 0.036461f
C4230 PAD.n4096 VSS 0.036461f
C4231 PAD.n4097 VSS 0.036461f
C4232 PAD.n4098 VSS 0.036461f
C4233 PAD.n4099 VSS 0.036461f
C4234 PAD.n4100 VSS 0.036461f
C4235 PAD.n4101 VSS 0.036461f
C4236 PAD.n4103 VSS 0.036461f
C4237 PAD.n4104 VSS 0.036461f
C4238 PAD.n4105 VSS 0.036461f
C4239 PAD.n4107 VSS 0.036461f
C4240 PAD.n4108 VSS 0.036461f
C4241 PAD.n4109 VSS 0.036461f
C4242 PAD.n4110 VSS 0.036461f
C4243 PAD.n4111 VSS 0.036461f
C4244 PAD.n4112 VSS 0.036461f
C4245 PAD.n4113 VSS 0.036461f
C4246 PAD.n4115 VSS 0.036461f
C4247 PAD.n4116 VSS 0.036461f
C4248 PAD.n4117 VSS 0.036461f
C4249 PAD.n4119 VSS 0.036461f
C4250 PAD.n4120 VSS 0.036461f
C4251 PAD.n4121 VSS 0.036461f
C4252 PAD.n4122 VSS 0.036461f
C4253 PAD.n4123 VSS 0.036461f
C4254 PAD.n4124 VSS 0.036461f
C4255 PAD.n4125 VSS 0.036461f
C4256 PAD.n4127 VSS 0.036461f
C4257 PAD.n4128 VSS 0.036461f
C4258 PAD.n4129 VSS 0.036461f
C4259 PAD.n4131 VSS 0.036461f
C4260 PAD.n4132 VSS 0.036461f
C4261 PAD.n4133 VSS 0.036461f
C4262 PAD.n4134 VSS 0.036461f
C4263 PAD.n4135 VSS 0.036461f
C4264 PAD.n4136 VSS 0.036461f
C4265 PAD.n4137 VSS 0.036461f
C4266 PAD.n4139 VSS 0.036461f
C4267 PAD.n4140 VSS 0.036461f
C4268 PAD.n4141 VSS 0.036461f
C4269 PAD.n4143 VSS 0.036461f
C4270 PAD.n4144 VSS 0.036461f
C4271 PAD.n4145 VSS 0.036461f
C4272 PAD.n4146 VSS 0.036461f
C4273 PAD.n4147 VSS 0.036461f
C4274 PAD.n4148 VSS 0.036461f
C4275 PAD.n4149 VSS 0.036461f
C4276 PAD.n4151 VSS 0.036461f
C4277 PAD.n4152 VSS 0.036461f
C4278 PAD.n4153 VSS 0.036461f
C4279 PAD.n4155 VSS 0.036461f
C4280 PAD.n4156 VSS 0.036461f
C4281 PAD.n4157 VSS 0.036461f
C4282 PAD.n4158 VSS 0.036461f
C4283 PAD.n4159 VSS 0.036461f
C4284 PAD.n4160 VSS 0.036461f
C4285 PAD.n4161 VSS 0.036461f
C4286 PAD.n4163 VSS 0.036461f
C4287 PAD.n4164 VSS 0.036461f
C4288 PAD.n4165 VSS 0.036461f
C4289 PAD.n4167 VSS 0.036461f
C4290 PAD.n4168 VSS 0.036461f
C4291 PAD.n4169 VSS 0.036461f
C4292 PAD.n4170 VSS 0.036461f
C4293 PAD.n4171 VSS 0.036461f
C4294 PAD.n4172 VSS 0.036461f
C4295 PAD.n4173 VSS 0.036461f
C4296 PAD.n4175 VSS 0.036461f
C4297 PAD.n4176 VSS 0.036461f
C4298 PAD.n4177 VSS 0.036461f
C4299 PAD.n4179 VSS 0.036461f
C4300 PAD.n4180 VSS 0.036461f
C4301 PAD.n4181 VSS 0.036461f
C4302 PAD.n4182 VSS 0.036461f
C4303 PAD.n4183 VSS 0.036461f
C4304 PAD.n4184 VSS 0.036461f
C4305 PAD.n4185 VSS 0.036461f
C4306 PAD.n4187 VSS 0.036461f
C4307 PAD.n4188 VSS 0.036461f
C4308 PAD.n4189 VSS 0.036461f
C4309 PAD.n4191 VSS 0.036461f
C4310 PAD.n4192 VSS 0.036461f
C4311 PAD.n4193 VSS 0.036461f
C4312 PAD.n4194 VSS 0.036461f
C4313 PAD.n4195 VSS 0.036461f
C4314 PAD.n4196 VSS 0.036461f
C4315 PAD.n4197 VSS 0.036461f
C4316 PAD.n4199 VSS 0.036461f
C4317 PAD.n4200 VSS 0.036461f
C4318 PAD.n4201 VSS 0.036461f
C4319 PAD.n4203 VSS 0.036461f
C4320 PAD.n4204 VSS 0.036461f
C4321 PAD.n4205 VSS 0.036461f
C4322 PAD.n4206 VSS 0.036461f
C4323 PAD.n4207 VSS 0.036461f
C4324 PAD.n4208 VSS 0.036461f
C4325 PAD.n4209 VSS 0.036461f
C4326 PAD.n4211 VSS 0.036461f
C4327 PAD.n4212 VSS 0.036461f
C4328 PAD.n4213 VSS 0.036461f
C4329 PAD.n4215 VSS 0.036461f
C4330 PAD.n4216 VSS 0.036461f
C4331 PAD.n4217 VSS 0.036461f
C4332 PAD.n4218 VSS 0.036461f
C4333 PAD.n4219 VSS 0.036461f
C4334 PAD.n4220 VSS 0.036461f
C4335 PAD.n4221 VSS 0.036461f
C4336 PAD.n4223 VSS 0.036461f
C4337 PAD.n4224 VSS 0.036461f
C4338 PAD.n4225 VSS 0.036461f
C4339 PAD.n4227 VSS 0.036461f
C4340 PAD.n4228 VSS 0.036461f
C4341 PAD.n4229 VSS 0.036461f
C4342 PAD.n4230 VSS 0.036461f
C4343 PAD.n4231 VSS 0.036461f
C4344 PAD.n4232 VSS 0.036461f
C4345 PAD.n4233 VSS 0.036461f
C4346 PAD.n4235 VSS 0.036461f
C4347 PAD.n4236 VSS 0.036461f
C4348 PAD.n4237 VSS 0.036461f
C4349 PAD.n4239 VSS 0.036461f
C4350 PAD.n4240 VSS 0.036461f
C4351 PAD.n4241 VSS 0.036461f
C4352 PAD.n4242 VSS 0.036461f
C4353 PAD.n4243 VSS 0.036461f
C4354 PAD.n4244 VSS 0.036461f
C4355 PAD.n4245 VSS 0.036461f
C4356 PAD.n4247 VSS 0.036461f
C4357 PAD.n4248 VSS 0.036461f
C4358 PAD.n4249 VSS 0.036461f
C4359 PAD.n4251 VSS 0.036461f
C4360 PAD.n4252 VSS 0.036461f
C4361 PAD.n4253 VSS 0.036461f
C4362 PAD.n4254 VSS 0.036461f
C4363 PAD.n4255 VSS 0.036461f
C4364 PAD.n4256 VSS 0.036461f
C4365 PAD.n4257 VSS 0.036461f
C4366 PAD.n4259 VSS 0.036461f
C4367 PAD.n4260 VSS 0.036461f
C4368 PAD.n4261 VSS 0.036461f
C4369 PAD.n4263 VSS 0.036461f
C4370 PAD.n4264 VSS 0.036461f
C4371 PAD.n4265 VSS 0.036461f
C4372 PAD.n4266 VSS 0.036461f
C4373 PAD.n4267 VSS 0.036461f
C4374 PAD.n4268 VSS 0.036461f
C4375 PAD.n4269 VSS 0.036461f
C4376 PAD.n4271 VSS 0.036461f
C4377 PAD.n4272 VSS 0.036461f
C4378 PAD.n4273 VSS 0.036461f
C4379 PAD.n4275 VSS 0.036461f
C4380 PAD.n4276 VSS 0.036461f
C4381 PAD.n4277 VSS 0.036461f
C4382 PAD.n4278 VSS 0.036461f
C4383 PAD.n4279 VSS 0.036461f
C4384 PAD.n4280 VSS 0.036461f
C4385 PAD.n4281 VSS 0.036461f
C4386 PAD.n4283 VSS 0.036461f
C4387 PAD.n4284 VSS 0.036461f
C4388 PAD.n4285 VSS 0.036461f
C4389 PAD.n4287 VSS 0.036461f
C4390 PAD.n4288 VSS 0.036461f
C4391 PAD.n4289 VSS 0.036461f
C4392 PAD.n4290 VSS 0.036461f
C4393 PAD.n4291 VSS 0.036461f
C4394 PAD.n4292 VSS 0.036461f
C4395 PAD.n4293 VSS 0.036461f
C4396 PAD.n4295 VSS 0.036461f
C4397 PAD.n4296 VSS 0.036461f
C4398 PAD.n4297 VSS 0.036461f
C4399 PAD.n4299 VSS 0.036461f
C4400 PAD.n4300 VSS 0.036461f
C4401 PAD.n4301 VSS 0.036461f
C4402 PAD.n4302 VSS 0.036461f
C4403 PAD.n4303 VSS 0.036461f
C4404 PAD.n4304 VSS 0.036461f
C4405 PAD.n4305 VSS 0.036461f
C4406 PAD.n4307 VSS 0.036461f
C4407 PAD.n4308 VSS 0.036461f
C4408 PAD.n4309 VSS 0.036461f
C4409 PAD.n4311 VSS 0.036461f
C4410 PAD.n4312 VSS 0.036461f
C4411 PAD.n4313 VSS 0.036461f
C4412 PAD.n4314 VSS 0.036461f
C4413 PAD.n4315 VSS 0.032474f
C4414 PAD.n4316 VSS 0.042895f
C4415 PAD.n4317 VSS 0.049115f
C4416 PAD.n4318 VSS 0.049115f
C4417 PAD.n4319 VSS 0.611734f
C4418 PAD.n4320 VSS 0.065264f
C4419 PAD.n4321 VSS 0.695601f
C4420 PAD.n4322 VSS 0.04726f
C4421 PAD.n4323 VSS 0.065264f
C4422 PAD.n4324 VSS 0.04726f
C4423 PAD.n4325 VSS 0.03338f
C4424 PAD.n4326 VSS 0.062274f
C4425 PAD.n4327 VSS 0.069765f
C4426 PAD.n4328 VSS 0.039761f
C4427 PAD.n4329 VSS 0.069765f
C4428 PAD.n4330 VSS 0.039761f
C4429 PAD.n4331 VSS 0.409467f
C4430 PAD.n4332 VSS 0.567334f
C4431 PAD.n4333 VSS 0.320667f
C4432 PAD.n4334 VSS 0.029436f
C4433 PAD.n4335 VSS 0.029436f
C4434 PAD.n4336 VSS 0.036461f
C4435 PAD.n4337 VSS 0.036461f
C4436 PAD.n4338 VSS 0.036461f
C4437 PAD.n4340 VSS 0.036461f
C4438 PAD.n4341 VSS 0.036461f
C4439 PAD.n4342 VSS 0.036461f
C4440 PAD.n4344 VSS 0.036461f
C4441 PAD.n4345 VSS 0.036461f
C4442 PAD.n4346 VSS 0.036461f
C4443 PAD.n4348 VSS 0.036461f
C4444 PAD.n4349 VSS 0.036461f
C4445 PAD.n4350 VSS 0.036461f
C4446 PAD.n4352 VSS 0.036461f
C4447 PAD.n4353 VSS 0.036461f
C4448 PAD.n4354 VSS 0.036461f
C4449 PAD.n4356 VSS 0.036461f
C4450 PAD.n4357 VSS 0.036461f
C4451 PAD.n4358 VSS 0.036461f
C4452 PAD.n4360 VSS 0.036461f
C4453 PAD.n4361 VSS 0.036461f
C4454 PAD.n4362 VSS 0.036461f
C4455 PAD.n4364 VSS 0.036461f
C4456 PAD.n4365 VSS 0.036461f
C4457 PAD.n4366 VSS 0.036461f
C4458 PAD.n4368 VSS 0.036461f
C4459 PAD.n4369 VSS 0.036461f
C4460 PAD.n4370 VSS 0.036461f
C4461 PAD.n4372 VSS 0.036461f
C4462 PAD.n4373 VSS 0.036461f
C4463 PAD.n4374 VSS 0.036461f
C4464 PAD.n4376 VSS 0.036461f
C4465 PAD.n4377 VSS 0.036461f
C4466 PAD.n4378 VSS 0.036461f
C4467 PAD.n4380 VSS 0.036461f
C4468 PAD.n4381 VSS 0.036461f
C4469 PAD.n4382 VSS 0.036461f
C4470 PAD.n4384 VSS 0.036461f
C4471 PAD.n4385 VSS 0.036461f
C4472 PAD.n4386 VSS 0.036461f
C4473 PAD.n4388 VSS 0.036461f
C4474 PAD.n4389 VSS 0.036461f
C4475 PAD.n4390 VSS 0.036461f
C4476 PAD.n4392 VSS 0.036461f
C4477 PAD.n4393 VSS 0.036461f
C4478 PAD.n4394 VSS 0.036461f
C4479 PAD.n4396 VSS 0.036461f
C4480 PAD.n4397 VSS 0.036461f
C4481 PAD.n4398 VSS 0.036461f
C4482 PAD.n4400 VSS 0.036461f
C4483 PAD.n4401 VSS 0.036461f
C4484 PAD.n4402 VSS 0.036461f
C4485 PAD.n4404 VSS 0.036461f
C4486 PAD.n4405 VSS 0.036461f
C4487 PAD.n4406 VSS 0.036461f
C4488 PAD.n4408 VSS 0.036461f
C4489 PAD.n4409 VSS 0.036461f
C4490 PAD.n4410 VSS 0.036461f
C4491 PAD.n4412 VSS 0.036461f
C4492 PAD.n4413 VSS 0.036461f
C4493 PAD.n4414 VSS 0.036461f
C4494 PAD.n4416 VSS 0.036461f
C4495 PAD.n4417 VSS 0.036461f
C4496 PAD.n4418 VSS 0.036461f
C4497 PAD.n4419 VSS 0.023109f
C4498 PAD.n4420 VSS 0.023109f
C4499 PAD.n4422 VSS 0.036461f
C4500 PAD.n4424 VSS 0.036461f
C4501 PAD.n4426 VSS 0.036461f
C4502 PAD.n4427 VSS 0.036461f
C4503 PAD.n4428 VSS 0.036461f
C4504 PAD.n4429 VSS 0.036461f
C4505 PAD.n4430 VSS 0.036461f
C4506 PAD.n4431 VSS 0.036461f
C4507 PAD.n4432 VSS 0.036461f
C4508 PAD.n4434 VSS 0.036461f
C4509 PAD.n4436 VSS 0.036461f
C4510 PAD.n4438 VSS 0.036461f
C4511 PAD.n4439 VSS 0.036461f
C4512 PAD.n4440 VSS 0.036461f
C4513 PAD.n4441 VSS 0.036461f
C4514 PAD.n4442 VSS 0.036461f
C4515 PAD.n4443 VSS 0.036461f
C4516 PAD.n4444 VSS 0.036461f
C4517 PAD.n4446 VSS 0.036461f
C4518 PAD.n4448 VSS 0.036461f
C4519 PAD.n4450 VSS 0.036461f
C4520 PAD.n4451 VSS 0.036461f
C4521 PAD.n4452 VSS 0.036461f
C4522 PAD.n4453 VSS 0.036461f
C4523 PAD.n4454 VSS 0.036461f
C4524 PAD.n4455 VSS 0.036461f
C4525 PAD.n4456 VSS 0.036461f
C4526 PAD.n4458 VSS 0.036461f
C4527 PAD.n4460 VSS 0.036461f
C4528 PAD.n4462 VSS 0.036461f
C4529 PAD.n4463 VSS 0.036461f
C4530 PAD.n4464 VSS 0.036461f
C4531 PAD.n4465 VSS 0.036461f
C4532 PAD.n4466 VSS 0.036461f
C4533 PAD.n4467 VSS 0.036461f
C4534 PAD.n4468 VSS 0.036461f
C4535 PAD.n4470 VSS 0.036461f
C4536 PAD.n4472 VSS 0.036461f
C4537 PAD.n4474 VSS 0.036461f
C4538 PAD.n4475 VSS 0.036461f
C4539 PAD.n4476 VSS 0.036461f
C4540 PAD.n4477 VSS 0.036461f
C4541 PAD.n4478 VSS 0.036461f
C4542 PAD.n4479 VSS 0.036461f
C4543 PAD.n4480 VSS 0.036461f
C4544 PAD.n4482 VSS 0.036461f
C4545 PAD.n4484 VSS 0.036461f
C4546 PAD.n4486 VSS 0.036461f
C4547 PAD.n4487 VSS 0.036461f
C4548 PAD.n4488 VSS 0.036461f
C4549 PAD.n4489 VSS 0.036461f
C4550 PAD.n4490 VSS 0.036461f
C4551 PAD.n4491 VSS 0.036461f
C4552 PAD.n4492 VSS 0.036461f
C4553 PAD.n4494 VSS 0.036461f
C4554 PAD.n4496 VSS 0.036461f
C4555 PAD.n4498 VSS 0.036461f
C4556 PAD.n4499 VSS 0.036461f
C4557 PAD.n4500 VSS 0.036461f
C4558 PAD.n4501 VSS 0.036461f
C4559 PAD.n4502 VSS 0.036461f
C4560 PAD.n4503 VSS 0.036461f
C4561 PAD.n4504 VSS 0.036461f
C4562 PAD.n4506 VSS 0.036461f
C4563 PAD.n4508 VSS 0.036461f
C4564 PAD.n4510 VSS 0.036461f
C4565 PAD.n4511 VSS 0.036461f
C4566 PAD.n4512 VSS 0.036461f
C4567 PAD.n4513 VSS 0.036461f
C4568 PAD.n4514 VSS 0.036461f
C4569 PAD.n4515 VSS 0.036461f
C4570 PAD.n4516 VSS 0.036461f
C4571 PAD.n4518 VSS 0.036461f
C4572 PAD.n4520 VSS 0.036461f
C4573 PAD.n4522 VSS 0.036461f
C4574 PAD.n4523 VSS 0.036461f
C4575 PAD.n4524 VSS 0.036461f
C4576 PAD.n4525 VSS 0.036461f
C4577 PAD.n4526 VSS 0.036461f
C4578 PAD.n4527 VSS 0.036461f
C4579 PAD.n4528 VSS 0.036461f
C4580 PAD.n4530 VSS 0.036461f
C4581 PAD.n4532 VSS 0.036461f
C4582 PAD.n4534 VSS 0.036461f
C4583 PAD.n4535 VSS 0.036461f
C4584 PAD.n4536 VSS 0.036461f
C4585 PAD.n4537 VSS 0.036461f
C4586 PAD.n4538 VSS 0.036461f
C4587 PAD.n4539 VSS 0.036461f
C4588 PAD.n4540 VSS 0.036461f
C4589 PAD.n4542 VSS 0.036461f
C4590 PAD.n4544 VSS 0.036461f
C4591 PAD.n4546 VSS 0.036461f
C4592 PAD.n4547 VSS 0.036461f
C4593 PAD.n4548 VSS 0.036461f
C4594 PAD.n4549 VSS 0.036461f
C4595 PAD.n4550 VSS 0.036461f
C4596 PAD.n4551 VSS 0.036461f
C4597 PAD.n4552 VSS 0.036461f
C4598 PAD.n4554 VSS 0.036461f
C4599 PAD.n4556 VSS 0.036461f
C4600 PAD.n4558 VSS 0.036461f
C4601 PAD.n4559 VSS 0.036461f
C4602 PAD.n4560 VSS 0.036461f
C4603 PAD.n4561 VSS 0.036461f
C4604 PAD.n4562 VSS 0.036461f
C4605 PAD.n4563 VSS 0.036461f
C4606 PAD.n4564 VSS 0.036461f
C4607 PAD.n4566 VSS 0.036461f
C4608 PAD.n4568 VSS 0.036461f
C4609 PAD.n4570 VSS 0.036461f
C4610 PAD.n4571 VSS 0.036461f
C4611 PAD.n4572 VSS 0.036461f
C4612 PAD.n4573 VSS 0.036461f
C4613 PAD.n4574 VSS 0.036461f
C4614 PAD.n4575 VSS 0.036461f
C4615 PAD.n4576 VSS 0.036461f
C4616 PAD.n4578 VSS 0.036461f
C4617 PAD.n4580 VSS 0.036461f
C4618 PAD.n4582 VSS 0.036461f
C4619 PAD.n4583 VSS 0.036461f
C4620 PAD.n4584 VSS 0.036461f
C4621 PAD.n4585 VSS 0.036461f
C4622 PAD.n4586 VSS 0.036461f
C4623 PAD.n4587 VSS 0.036461f
C4624 PAD.n4588 VSS 0.036461f
C4625 PAD.n4590 VSS 0.036461f
C4626 PAD.n4592 VSS 0.036461f
C4627 PAD.n4594 VSS 0.036461f
C4628 PAD.n4595 VSS 0.036461f
C4629 PAD.n4596 VSS 0.036461f
C4630 PAD.n4597 VSS 0.036461f
C4631 PAD.n4598 VSS 0.036461f
C4632 PAD.n4599 VSS 0.036461f
C4633 PAD.n4600 VSS 0.036461f
C4634 PAD.n4602 VSS 0.036461f
C4635 PAD.n4604 VSS 0.036461f
C4636 PAD.n4606 VSS 0.036461f
C4637 PAD.n4607 VSS 0.036461f
C4638 PAD.n4608 VSS 0.036461f
C4639 PAD.n4609 VSS 0.036461f
C4640 PAD.n4610 VSS 0.036461f
C4641 PAD.n4611 VSS 0.036461f
C4642 PAD.n4612 VSS 0.036461f
C4643 PAD.n4614 VSS 0.036461f
C4644 PAD.n4616 VSS 0.036461f
C4645 PAD.n4618 VSS 0.036461f
C4646 PAD.n4619 VSS 0.036461f
C4647 PAD.n4620 VSS 0.036461f
C4648 PAD.n4621 VSS 0.036461f
C4649 PAD.n4622 VSS 0.036461f
C4650 PAD.n4623 VSS 0.036461f
C4651 PAD.n4624 VSS 0.036461f
C4652 PAD.n4626 VSS 0.036461f
C4653 PAD.n4628 VSS 0.036461f
C4654 PAD.n4630 VSS 0.036461f
C4655 PAD.n4631 VSS 0.036461f
C4656 PAD.n4632 VSS 0.036461f
C4657 PAD.n4633 VSS 0.036461f
C4658 PAD.n4634 VSS 0.036461f
C4659 PAD.n4635 VSS 0.036461f
C4660 PAD.n4636 VSS 0.036461f
C4661 PAD.n4638 VSS 0.036461f
C4662 PAD.n4640 VSS 0.036461f
C4663 PAD.n4642 VSS 0.036461f
C4664 PAD.n4643 VSS 0.036461f
C4665 PAD.n4644 VSS 0.036461f
C4666 PAD.n4645 VSS 0.036461f
C4667 PAD.n4646 VSS 0.036461f
C4668 PAD.n4647 VSS 0.036461f
C4669 PAD.n4648 VSS 0.036461f
C4670 PAD.n4650 VSS 0.036461f
C4671 PAD.n4652 VSS 0.036461f
C4672 PAD.n4654 VSS 0.036461f
C4673 PAD.n4655 VSS 0.036461f
C4674 PAD.n4656 VSS 0.036461f
C4675 PAD.n4657 VSS 0.036461f
C4676 PAD.n4658 VSS 0.036461f
C4677 PAD.n4659 VSS 0.036461f
C4678 PAD.n4660 VSS 0.036461f
C4679 PAD.n4661 VSS 0.036461f
C4680 PAD.n4663 VSS 0.036461f
C4681 PAD.n4665 VSS 0.036461f
C4682 PAD.n4667 VSS 0.023109f
C4683 PAD.n4668 VSS 0.023109f
C4684 PAD.n4669 VSS 0.030555f
C4685 PAD.n4670 VSS 0.042895f
C4686 PAD.n4671 VSS 0.049115f
C4687 PAD.n4672 VSS 0.049115f
C4688 PAD.n4673 VSS 0.587068f
C4689 PAD.n4674 VSS 0.038258f
C4690 PAD.n4675 VSS 0.038258f
C4691 PAD.n4676 VSS 0.03338f
C4692 PAD.n4677 VSS 0.062274f
C4693 PAD.n4678 VSS 0.069765f
C4694 PAD.n4679 VSS 0.039761f
C4695 PAD.n4680 VSS 0.069765f
C4696 PAD.n4681 VSS 0.039761f
C4697 PAD.n4682 VSS 0.611734f
C4698 PAD.n4724 VSS 0.424267f
C4699 PAD.n4725 VSS 0.036461f
C4700 PAD.n4727 VSS 0.036461f
C4701 PAD.n4728 VSS 0.036461f
C4702 PAD.n4729 VSS 0.036461f
C4703 PAD.n4730 VSS 0.036461f
C4704 PAD.n4731 VSS 0.036461f
C4705 PAD.n4733 VSS 0.036461f
C4706 PAD.n4734 VSS 0.036461f
C4707 PAD.n4735 VSS 0.036461f
C4708 PAD.n4736 VSS 0.036461f
C4709 PAD.n4738 VSS 0.036461f
C4710 PAD.n4739 VSS 0.036461f
C4711 PAD.n4740 VSS 0.036461f
C4712 PAD.n4741 VSS 0.036461f
C4713 PAD.n4743 VSS 0.036461f
C4714 PAD.n4744 VSS 0.036461f
C4715 PAD.n4745 VSS 0.036461f
C4716 PAD.n4746 VSS 0.036461f
C4717 PAD.n4748 VSS 0.036461f
C4718 PAD.n4749 VSS 0.036461f
C4719 PAD.n4750 VSS 0.036461f
C4720 PAD.n4751 VSS 0.036461f
C4721 PAD.n4753 VSS 0.036461f
C4722 PAD.n4754 VSS 0.036461f
C4723 PAD.n4755 VSS 0.036461f
C4724 PAD.n4756 VSS 0.036461f
C4725 PAD.n4758 VSS 0.036461f
C4726 PAD.n4759 VSS 0.036461f
C4727 PAD.n4760 VSS 0.036461f
C4728 PAD.n4761 VSS 0.036461f
C4729 PAD.n4763 VSS 0.036461f
C4730 PAD.n4764 VSS 0.036461f
C4731 PAD.n4765 VSS 0.036461f
C4732 PAD.n4766 VSS 0.036461f
C4733 PAD.n4768 VSS 0.036461f
C4734 PAD.n4769 VSS 0.036461f
C4735 PAD.n4770 VSS 0.036461f
C4736 PAD.n4771 VSS 0.036461f
C4737 PAD.n4773 VSS 0.036461f
C4738 PAD.n4774 VSS 0.036461f
C4739 PAD.n4775 VSS 0.036461f
C4740 PAD.n4776 VSS 0.036461f
C4741 PAD.n4778 VSS 0.036461f
C4742 PAD.n4779 VSS 0.036461f
C4743 PAD.n4780 VSS 0.036461f
C4744 PAD.n4781 VSS 0.036461f
C4745 PAD.n4783 VSS 0.036461f
C4746 PAD.n4784 VSS 0.036461f
C4747 PAD.n4785 VSS 0.036461f
C4748 PAD.n4786 VSS 0.036461f
C4749 PAD.n4788 VSS 0.036461f
C4750 PAD.n4789 VSS 0.036461f
C4751 PAD.n4790 VSS 0.036461f
C4752 PAD.n4791 VSS 0.036461f
C4753 PAD.n4793 VSS 0.036461f
C4754 PAD.n4794 VSS 0.036461f
C4755 PAD.n4795 VSS 0.036461f
C4756 PAD.n4796 VSS 0.036461f
C4757 PAD.n4798 VSS 0.036461f
C4758 PAD.n4799 VSS 0.036461f
C4759 PAD.n4800 VSS 0.036461f
C4760 PAD.n4801 VSS 0.036461f
C4761 PAD.n4803 VSS 0.036461f
C4762 PAD.n4804 VSS 0.036461f
C4763 PAD.n4805 VSS 0.036461f
C4764 PAD.n4806 VSS 0.036461f
C4765 PAD.n4808 VSS 0.036461f
C4766 PAD.n4809 VSS 0.036461f
C4767 PAD.n4810 VSS 0.036461f
C4768 PAD.n4811 VSS 0.036461f
C4769 PAD.n4813 VSS 0.036461f
C4770 PAD.n4814 VSS 0.036461f
C4771 PAD.n4815 VSS 0.036461f
C4772 PAD.n4816 VSS 0.036461f
C4773 PAD.n4818 VSS 0.036461f
C4774 PAD.n4819 VSS 0.036461f
C4775 PAD.n4820 VSS 0.036461f
C4776 PAD.n4821 VSS 0.036461f
C4777 PAD.n4823 VSS 0.036461f
C4778 PAD.n4824 VSS 0.036461f
C4779 PAD.n4825 VSS 0.036461f
C4780 PAD.n4826 VSS 0.036461f
C4781 PAD.n4828 VSS 0.036461f
C4782 PAD.n4829 VSS 0.023109f
C4783 PAD.n4830 VSS 0.040328f
C4784 PAD.n4831 VSS 0.029436f
C4785 PAD.n4832 VSS 0.023109f
C4786 PAD.n4833 VSS 0.047559f
C4787 PAD.n4834 VSS 0.029436f
C4788 PAD.n4835 VSS 0.030555f
C4789 PAD.n4836 VSS 0.042895f
C4790 PAD.n4837 VSS 0.049115f
C4791 PAD.n4838 VSS 0.049115f
C4792 PAD.n4839 VSS 0.029436f
C4793 PAD.n4840 VSS 0.37f
C4794 PAD.n4841 VSS 0.700534f
C4795 PAD.n4842 VSS 0.434134f
C4796 PAD.n4843 VSS 0.458801f
C4797 PAD.n4844 VSS 0.039761f
C4798 PAD.n4845 VSS 0.039761f
C4799 PAD.n4846 VSS 0.036461f
C4800 PAD.n4847 VSS 0.023109f
C4801 PAD.n4848 VSS 0.036461f
C4802 PAD.n4851 VSS 0.036461f
C4803 PAD.n4852 VSS 0.036461f
C4804 PAD.n4853 VSS 0.036461f
C4805 PAD.n4854 VSS 0.036461f
C4806 PAD.n4856 VSS 0.036461f
C4807 PAD.n4857 VSS 0.036461f
C4808 PAD.n4858 VSS 0.036461f
C4809 PAD.n4860 VSS 0.036461f
C4810 PAD.n4861 VSS 0.036461f
C4811 PAD.n4862 VSS 0.036461f
C4812 PAD.n4864 VSS 0.036461f
C4813 PAD.n4865 VSS 0.036461f
C4814 PAD.n4866 VSS 0.036461f
C4815 PAD.n4868 VSS 0.036461f
C4816 PAD.n4869 VSS 0.036461f
C4817 PAD.n4870 VSS 0.036461f
C4818 PAD.n4872 VSS 0.036461f
C4819 PAD.n4873 VSS 0.036461f
C4820 PAD.n4874 VSS 0.036461f
C4821 PAD.n4876 VSS 0.036461f
C4822 PAD.n4877 VSS 0.036461f
C4823 PAD.n4878 VSS 0.036461f
C4824 PAD.n4880 VSS 0.036461f
C4825 PAD.n4881 VSS 0.036461f
C4826 PAD.n4882 VSS 0.036461f
C4827 PAD.n4884 VSS 0.036461f
C4828 PAD.n4885 VSS 0.036461f
C4829 PAD.n4886 VSS 0.036461f
C4830 PAD.n4888 VSS 0.036461f
C4831 PAD.n4889 VSS 0.036461f
C4832 PAD.n4890 VSS 0.036461f
C4833 PAD.n4892 VSS 0.036461f
C4834 PAD.n4893 VSS 0.036461f
C4835 PAD.n4894 VSS 0.036461f
C4836 PAD.n4896 VSS 0.036461f
C4837 PAD.n4897 VSS 0.036461f
C4838 PAD.n4898 VSS 0.036461f
C4839 PAD.n4900 VSS 0.036461f
C4840 PAD.n4901 VSS 0.036461f
C4841 PAD.n4902 VSS 0.036461f
C4842 PAD.n4904 VSS 0.036461f
C4843 PAD.n4905 VSS 0.036461f
C4844 PAD.n4906 VSS 0.036461f
C4845 PAD.n4908 VSS 0.036461f
C4846 PAD.n4909 VSS 0.036461f
C4847 PAD.n4910 VSS 0.036461f
C4848 PAD.n4912 VSS 0.036461f
C4849 PAD.n4913 VSS 0.036461f
C4850 PAD.n4914 VSS 0.036461f
C4851 PAD.n4916 VSS 0.036461f
C4852 PAD.n4917 VSS 0.036461f
C4853 PAD.n4918 VSS 0.036461f
C4854 PAD.n4920 VSS 0.036461f
C4855 PAD.n4921 VSS 0.036461f
C4856 PAD.n4922 VSS 0.036461f
C4857 PAD.n4924 VSS 0.036461f
C4858 PAD.n4925 VSS 0.036461f
C4859 PAD.n4926 VSS 0.036461f
C4860 PAD.n4928 VSS 0.036461f
C4861 PAD.n4929 VSS 0.036461f
C4862 PAD.n4930 VSS 0.036461f
C4863 PAD.n4931 VSS 0.023109f
C4864 PAD.n4932 VSS 0.023109f
C4865 PAD.n4934 VSS 0.036461f
C4866 PAD.n4936 VSS 0.036461f
C4867 PAD.n4938 VSS 0.036461f
C4868 PAD.n4939 VSS 0.036461f
C4869 PAD.n4940 VSS 0.036461f
C4870 PAD.n4941 VSS 0.036461f
C4871 PAD.n4942 VSS 0.036461f
C4872 PAD.n4943 VSS 0.036461f
C4873 PAD.n4944 VSS 0.036461f
C4874 PAD.n4946 VSS 0.036461f
C4875 PAD.n4948 VSS 0.036461f
C4876 PAD.n4950 VSS 0.036461f
C4877 PAD.n4951 VSS 0.036461f
C4878 PAD.n4952 VSS 0.036461f
C4879 PAD.n4953 VSS 0.036461f
C4880 PAD.n4954 VSS 0.036461f
C4881 PAD.n4955 VSS 0.036461f
C4882 PAD.n4956 VSS 0.036461f
C4883 PAD.n4958 VSS 0.036461f
C4884 PAD.n4960 VSS 0.036461f
C4885 PAD.n4962 VSS 0.036461f
C4886 PAD.n4963 VSS 0.036461f
C4887 PAD.n4964 VSS 0.036461f
C4888 PAD.n4965 VSS 0.036461f
C4889 PAD.n4966 VSS 0.036461f
C4890 PAD.n4967 VSS 0.036461f
C4891 PAD.n4968 VSS 0.036461f
C4892 PAD.n4970 VSS 0.036461f
C4893 PAD.n4972 VSS 0.036461f
C4894 PAD.n4974 VSS 0.036461f
C4895 PAD.n4975 VSS 0.036461f
C4896 PAD.n4976 VSS 0.036461f
C4897 PAD.n4977 VSS 0.036461f
C4898 PAD.n4978 VSS 0.036461f
C4899 PAD.n4979 VSS 0.036461f
C4900 PAD.n4980 VSS 0.036461f
C4901 PAD.n4982 VSS 0.036461f
C4902 PAD.n4984 VSS 0.036461f
C4903 PAD.n4986 VSS 0.036461f
C4904 PAD.n4987 VSS 0.036461f
C4905 PAD.n4988 VSS 0.036461f
C4906 PAD.n4989 VSS 0.036461f
C4907 PAD.n4990 VSS 0.036461f
C4908 PAD.n4991 VSS 0.036461f
C4909 PAD.n4992 VSS 0.036461f
C4910 PAD.n4994 VSS 0.036461f
C4911 PAD.n4996 VSS 0.036461f
C4912 PAD.n4998 VSS 0.036461f
C4913 PAD.n4999 VSS 0.036461f
C4914 PAD.n5000 VSS 0.036461f
C4915 PAD.n5001 VSS 0.036461f
C4916 PAD.n5002 VSS 0.036461f
C4917 PAD.n5003 VSS 0.036461f
C4918 PAD.n5004 VSS 0.036461f
C4919 PAD.n5006 VSS 0.036461f
C4920 PAD.n5008 VSS 0.036461f
C4921 PAD.n5010 VSS 0.036461f
C4922 PAD.n5011 VSS 0.036461f
C4923 PAD.n5012 VSS 0.036461f
C4924 PAD.n5013 VSS 0.036461f
C4925 PAD.n5014 VSS 0.036461f
C4926 PAD.n5015 VSS 0.036461f
C4927 PAD.n5016 VSS 0.036461f
C4928 PAD.n5018 VSS 0.036461f
C4929 PAD.n5020 VSS 0.036461f
C4930 PAD.n5022 VSS 0.036461f
C4931 PAD.n5023 VSS 0.036461f
C4932 PAD.n5024 VSS 0.036461f
C4933 PAD.n5025 VSS 0.036461f
C4934 PAD.n5026 VSS 0.036461f
C4935 PAD.n5027 VSS 0.036461f
C4936 PAD.n5028 VSS 0.036461f
C4937 PAD.n5030 VSS 0.036461f
C4938 PAD.n5032 VSS 0.036461f
C4939 PAD.n5034 VSS 0.036461f
C4940 PAD.n5035 VSS 0.036461f
C4941 PAD.n5036 VSS 0.036461f
C4942 PAD.n5037 VSS 0.036461f
C4943 PAD.n5038 VSS 0.036461f
C4944 PAD.n5039 VSS 0.036461f
C4945 PAD.n5040 VSS 0.036461f
C4946 PAD.n5042 VSS 0.036461f
C4947 PAD.n5044 VSS 0.036461f
C4948 PAD.n5046 VSS 0.036461f
C4949 PAD.n5047 VSS 0.036461f
C4950 PAD.n5048 VSS 0.036461f
C4951 PAD.n5049 VSS 0.036461f
C4952 PAD.n5050 VSS 0.036461f
C4953 PAD.n5051 VSS 0.036461f
C4954 PAD.n5052 VSS 0.036461f
C4955 PAD.n5054 VSS 0.036461f
C4956 PAD.n5056 VSS 0.036461f
C4957 PAD.n5058 VSS 0.036461f
C4958 PAD.n5059 VSS 0.036461f
C4959 PAD.n5060 VSS 0.036461f
C4960 PAD.n5061 VSS 0.036461f
C4961 PAD.n5062 VSS 0.036461f
C4962 PAD.n5063 VSS 0.036461f
C4963 PAD.n5064 VSS 0.036461f
C4964 PAD.n5066 VSS 0.036461f
C4965 PAD.n5068 VSS 0.036461f
C4966 PAD.n5070 VSS 0.036461f
C4967 PAD.n5071 VSS 0.036461f
C4968 PAD.n5072 VSS 0.036461f
C4969 PAD.n5073 VSS 0.036461f
C4970 PAD.n5074 VSS 0.036461f
C4971 PAD.n5075 VSS 0.036461f
C4972 PAD.n5076 VSS 0.036461f
C4973 PAD.n5078 VSS 0.036461f
C4974 PAD.n5080 VSS 0.036461f
C4975 PAD.n5082 VSS 0.036461f
C4976 PAD.n5083 VSS 0.036461f
C4977 PAD.n5084 VSS 0.036461f
C4978 PAD.n5085 VSS 0.036461f
C4979 PAD.n5086 VSS 0.036461f
C4980 PAD.n5087 VSS 0.036461f
C4981 PAD.n5088 VSS 0.036461f
C4982 PAD.n5090 VSS 0.036461f
C4983 PAD.n5092 VSS 0.036461f
C4984 PAD.n5094 VSS 0.036461f
C4985 PAD.n5095 VSS 0.036461f
C4986 PAD.n5096 VSS 0.036461f
C4987 PAD.n5097 VSS 0.036461f
C4988 PAD.n5098 VSS 0.036461f
C4989 PAD.n5099 VSS 0.036461f
C4990 PAD.n5100 VSS 0.036461f
C4991 PAD.n5102 VSS 0.036461f
C4992 PAD.n5104 VSS 0.036461f
C4993 PAD.n5106 VSS 0.036461f
C4994 PAD.n5107 VSS 0.036461f
C4995 PAD.n5108 VSS 0.036461f
C4996 PAD.n5109 VSS 0.036461f
C4997 PAD.n5110 VSS 0.036461f
C4998 PAD.n5111 VSS 0.036461f
C4999 PAD.n5112 VSS 0.036461f
C5000 PAD.n5114 VSS 0.036461f
C5001 PAD.n5116 VSS 0.036461f
C5002 PAD.n5118 VSS 0.036461f
C5003 PAD.n5119 VSS 0.036461f
C5004 PAD.n5120 VSS 0.036461f
C5005 PAD.n5121 VSS 0.036461f
C5006 PAD.n5122 VSS 0.036461f
C5007 PAD.n5123 VSS 0.036461f
C5008 PAD.n5124 VSS 0.036461f
C5009 PAD.n5126 VSS 0.036461f
C5010 PAD.n5128 VSS 0.036461f
C5011 PAD.n5130 VSS 0.036461f
C5012 PAD.n5131 VSS 0.036461f
C5013 PAD.n5132 VSS 0.036461f
C5014 PAD.n5133 VSS 0.036461f
C5015 PAD.n5134 VSS 0.036461f
C5016 PAD.n5135 VSS 0.036461f
C5017 PAD.n5136 VSS 0.036461f
C5018 PAD.n5138 VSS 0.036461f
C5019 PAD.n5140 VSS 0.036461f
C5020 PAD.n5142 VSS 0.036461f
C5021 PAD.n5143 VSS 0.036461f
C5022 PAD.n5144 VSS 0.036461f
C5023 PAD.n5145 VSS 0.036461f
C5024 PAD.n5146 VSS 0.036461f
C5025 PAD.n5147 VSS 0.036461f
C5026 PAD.n5148 VSS 0.036461f
C5027 PAD.n5150 VSS 0.036461f
C5028 PAD.n5152 VSS 0.036461f
C5029 PAD.n5154 VSS 0.036461f
C5030 PAD.n5155 VSS 0.036461f
C5031 PAD.n5156 VSS 0.036461f
C5032 PAD.n5157 VSS 0.036461f
C5033 PAD.n5158 VSS 0.036461f
C5034 PAD.n5159 VSS 0.036461f
C5035 PAD.n5160 VSS 0.036461f
C5036 PAD.n5162 VSS 0.036461f
C5037 PAD.n5164 VSS 0.036461f
C5038 PAD.n5166 VSS 0.036461f
C5039 PAD.n5167 VSS 0.036461f
C5040 PAD.n5168 VSS 0.036461f
C5041 PAD.n5169 VSS 0.036461f
C5042 PAD.n5170 VSS 0.036461f
C5043 PAD.n5171 VSS 0.036461f
C5044 PAD.n5172 VSS 0.036461f
C5045 PAD.n5174 VSS 0.036461f
C5046 PAD.n5176 VSS 0.036461f
C5047 PAD.n5177 VSS 0.036461f
C5048 PAD.n5178 VSS 0.023109f
C5049 PAD.n5179 VSS 0.03338f
C5050 PAD.n5180 VSS 0.062274f
C5051 PAD.n5181 VSS 0.069765f
C5052 PAD.n5182 VSS 0.069765f
C5053 PAD.n5183 VSS 0.1924f
C5054 PAD.n5184 VSS 0.029436f
C5055 PAD.n5185 VSS 0.029436f
C5056 PAD.n5186 VSS 0.030555f
C5057 PAD.n5187 VSS 0.042895f
C5058 PAD.n5188 VSS 0.049115f
C5059 PAD.n5189 VSS 0.049115f
C5060 PAD.n5190 VSS 0.172667f
C5061 PAD.n5191 VSS 0.039761f
C5062 PAD.n5192 VSS 0.039761f
C5063 PAD.n5193 VSS 0.03338f
C5064 PAD.n5194 VSS 0.051727f
C5065 PAD.n5195 VSS 0.069765f
C5066 PAD.n5196 VSS 0.061889f
C5067 PAD.n5197 VSS 0.537734f
C5068 PAD.n5198 VSS 0.029436f
C5069 PAD.n5199 VSS 0.029436f
C5070 PAD.n5200 VSS 0.030555f
C5071 PAD.n5201 VSS 0.042895f
C5072 PAD.n5202 VSS 0.049115f
C5073 PAD.n5203 VSS 0.049115f
C5074 PAD.n5204 VSS 0.448934f
C5075 PAD.n5205 VSS 0.069765f
C5076 PAD.n5206 VSS 0.039761f
C5077 PAD.n5207 VSS 0.069765f
C5078 PAD.n5208 VSS 0.039761f
C5079 PAD.n5209 VSS 0.062274f
C5080 PAD.n5210 VSS 0.036461f
C5081 PAD.n5211 VSS 0.023109f
C5082 PAD.n5212 VSS 0.036461f
C5083 PAD.n5215 VSS 0.036461f
C5084 PAD.n5216 VSS 0.036461f
C5085 PAD.n5217 VSS 0.036461f
C5086 PAD.n5218 VSS 0.036461f
C5087 PAD.n5220 VSS 0.036461f
C5088 PAD.n5221 VSS 0.036461f
C5089 PAD.n5222 VSS 0.036461f
C5090 PAD.n5224 VSS 0.036461f
C5091 PAD.n5225 VSS 0.036461f
C5092 PAD.n5226 VSS 0.036461f
C5093 PAD.n5228 VSS 0.036461f
C5094 PAD.n5229 VSS 0.036461f
C5095 PAD.n5230 VSS 0.036461f
C5096 PAD.n5232 VSS 0.036461f
C5097 PAD.n5233 VSS 0.036461f
C5098 PAD.n5234 VSS 0.036461f
C5099 PAD.n5236 VSS 0.036461f
C5100 PAD.n5237 VSS 0.036461f
C5101 PAD.n5238 VSS 0.036461f
C5102 PAD.n5240 VSS 0.036461f
C5103 PAD.n5241 VSS 0.036461f
C5104 PAD.n5242 VSS 0.036461f
C5105 PAD.n5244 VSS 0.036461f
C5106 PAD.n5245 VSS 0.036461f
C5107 PAD.n5246 VSS 0.036461f
C5108 PAD.n5248 VSS 0.036461f
C5109 PAD.n5249 VSS 0.036461f
C5110 PAD.n5250 VSS 0.036461f
C5111 PAD.n5252 VSS 0.036461f
C5112 PAD.n5253 VSS 0.036461f
C5113 PAD.n5254 VSS 0.036461f
C5114 PAD.n5256 VSS 0.036461f
C5115 PAD.n5257 VSS 0.036461f
C5116 PAD.n5258 VSS 0.036461f
C5117 PAD.n5260 VSS 0.036461f
C5118 PAD.n5261 VSS 0.036461f
C5119 PAD.n5262 VSS 0.036461f
C5120 PAD.n5264 VSS 0.036461f
C5121 PAD.n5265 VSS 0.036461f
C5122 PAD.n5266 VSS 0.036461f
C5123 PAD.n5268 VSS 0.036461f
C5124 PAD.n5269 VSS 0.036461f
C5125 PAD.n5270 VSS 0.036461f
C5126 PAD.n5272 VSS 0.036461f
C5127 PAD.n5273 VSS 0.036461f
C5128 PAD.n5274 VSS 0.036461f
C5129 PAD.n5276 VSS 0.036461f
C5130 PAD.n5277 VSS 0.036461f
C5131 PAD.n5278 VSS 0.036461f
C5132 PAD.n5280 VSS 0.036461f
C5133 PAD.n5281 VSS 0.036461f
C5134 PAD.n5282 VSS 0.036461f
C5135 PAD.n5284 VSS 0.036461f
C5136 PAD.n5285 VSS 0.036461f
C5137 PAD.n5286 VSS 0.036461f
C5138 PAD.n5288 VSS 0.036461f
C5139 PAD.n5289 VSS 0.036461f
C5140 PAD.n5290 VSS 0.036461f
C5141 PAD.n5292 VSS 0.036461f
C5142 PAD.n5293 VSS 0.036461f
C5143 PAD.n5294 VSS 0.036461f
C5144 PAD.n5295 VSS 0.023109f
C5145 PAD.n5296 VSS 0.023109f
C5146 PAD.n5298 VSS 0.036461f
C5147 PAD.n5300 VSS 0.036461f
C5148 PAD.n5302 VSS 0.036461f
C5149 PAD.n5303 VSS 0.036461f
C5150 PAD.n5304 VSS 0.036461f
C5151 PAD.n5305 VSS 0.036461f
C5152 PAD.n5306 VSS 0.036461f
C5153 PAD.n5307 VSS 0.036461f
C5154 PAD.n5308 VSS 0.036461f
C5155 PAD.n5310 VSS 0.036461f
C5156 PAD.n5312 VSS 0.036461f
C5157 PAD.n5314 VSS 0.036461f
C5158 PAD.n5315 VSS 0.036461f
C5159 PAD.n5316 VSS 0.036461f
C5160 PAD.n5317 VSS 0.036461f
C5161 PAD.n5318 VSS 0.036461f
C5162 PAD.n5319 VSS 0.036461f
C5163 PAD.n5320 VSS 0.036461f
C5164 PAD.n5322 VSS 0.036461f
C5165 PAD.n5324 VSS 0.036461f
C5166 PAD.n5326 VSS 0.036461f
C5167 PAD.n5327 VSS 0.036461f
C5168 PAD.n5328 VSS 0.036461f
C5169 PAD.n5329 VSS 0.036461f
C5170 PAD.n5330 VSS 0.036461f
C5171 PAD.n5331 VSS 0.036461f
C5172 PAD.n5332 VSS 0.036461f
C5173 PAD.n5334 VSS 0.036461f
C5174 PAD.n5336 VSS 0.036461f
C5175 PAD.n5338 VSS 0.036461f
C5176 PAD.n5339 VSS 0.036461f
C5177 PAD.n5340 VSS 0.036461f
C5178 PAD.n5341 VSS 0.036461f
C5179 PAD.n5342 VSS 0.036461f
C5180 PAD.n5343 VSS 0.036461f
C5181 PAD.n5344 VSS 0.036461f
C5182 PAD.n5346 VSS 0.036461f
C5183 PAD.n5348 VSS 0.036461f
C5184 PAD.n5350 VSS 0.036461f
C5185 PAD.n5351 VSS 0.036461f
C5186 PAD.n5352 VSS 0.036461f
C5187 PAD.n5353 VSS 0.036461f
C5188 PAD.n5354 VSS 0.036461f
C5189 PAD.n5355 VSS 0.036461f
C5190 PAD.n5356 VSS 0.036461f
C5191 PAD.n5358 VSS 0.036461f
C5192 PAD.n5360 VSS 0.036461f
C5193 PAD.n5362 VSS 0.036461f
C5194 PAD.n5363 VSS 0.036461f
C5195 PAD.n5364 VSS 0.036461f
C5196 PAD.n5365 VSS 0.036461f
C5197 PAD.n5366 VSS 0.036461f
C5198 PAD.n5367 VSS 0.036461f
C5199 PAD.n5368 VSS 0.036461f
C5200 PAD.n5370 VSS 0.036461f
C5201 PAD.n5372 VSS 0.036461f
C5202 PAD.n5374 VSS 0.036461f
C5203 PAD.n5375 VSS 0.036461f
C5204 PAD.n5376 VSS 0.036461f
C5205 PAD.n5377 VSS 0.036461f
C5206 PAD.n5378 VSS 0.036461f
C5207 PAD.n5379 VSS 0.036461f
C5208 PAD.n5380 VSS 0.036461f
C5209 PAD.n5382 VSS 0.036461f
C5210 PAD.n5384 VSS 0.036461f
C5211 PAD.n5386 VSS 0.036461f
C5212 PAD.n5387 VSS 0.036461f
C5213 PAD.n5388 VSS 0.036461f
C5214 PAD.n5389 VSS 0.036461f
C5215 PAD.n5390 VSS 0.036461f
C5216 PAD.n5391 VSS 0.036461f
C5217 PAD.n5392 VSS 0.036461f
C5218 PAD.n5394 VSS 0.036461f
C5219 PAD.n5396 VSS 0.036461f
C5220 PAD.n5398 VSS 0.036461f
C5221 PAD.n5399 VSS 0.036461f
C5222 PAD.n5400 VSS 0.036461f
C5223 PAD.n5401 VSS 0.036461f
C5224 PAD.n5402 VSS 0.036461f
C5225 PAD.n5403 VSS 0.036461f
C5226 PAD.n5404 VSS 0.036461f
C5227 PAD.n5406 VSS 0.036461f
C5228 PAD.n5408 VSS 0.036461f
C5229 PAD.n5410 VSS 0.036461f
C5230 PAD.n5411 VSS 0.036461f
C5231 PAD.n5412 VSS 0.036461f
C5232 PAD.n5413 VSS 0.036461f
C5233 PAD.n5414 VSS 0.036461f
C5234 PAD.n5415 VSS 0.036461f
C5235 PAD.n5416 VSS 0.036461f
C5236 PAD.n5418 VSS 0.036461f
C5237 PAD.n5420 VSS 0.036461f
C5238 PAD.n5422 VSS 0.036461f
C5239 PAD.n5423 VSS 0.036461f
C5240 PAD.n5424 VSS 0.036461f
C5241 PAD.n5425 VSS 0.036461f
C5242 PAD.n5426 VSS 0.036461f
C5243 PAD.n5427 VSS 0.036461f
C5244 PAD.n5428 VSS 0.036461f
C5245 PAD.n5430 VSS 0.036461f
C5246 PAD.n5432 VSS 0.036461f
C5247 PAD.n5434 VSS 0.036461f
C5248 PAD.n5435 VSS 0.036461f
C5249 PAD.n5436 VSS 0.036461f
C5250 PAD.n5437 VSS 0.036461f
C5251 PAD.n5438 VSS 0.036461f
C5252 PAD.n5439 VSS 0.036461f
C5253 PAD.n5440 VSS 0.036461f
C5254 PAD.n5442 VSS 0.036461f
C5255 PAD.n5444 VSS 0.036461f
C5256 PAD.n5446 VSS 0.036461f
C5257 PAD.n5447 VSS 0.036461f
C5258 PAD.n5448 VSS 0.036461f
C5259 PAD.n5449 VSS 0.036461f
C5260 PAD.n5450 VSS 0.036461f
C5261 PAD.n5451 VSS 0.036461f
C5262 PAD.n5452 VSS 0.036461f
C5263 PAD.n5454 VSS 0.036461f
C5264 PAD.n5456 VSS 0.036461f
C5265 PAD.n5458 VSS 0.036461f
C5266 PAD.n5459 VSS 0.036461f
C5267 PAD.n5460 VSS 0.036461f
C5268 PAD.n5461 VSS 0.036461f
C5269 PAD.n5462 VSS 0.036461f
C5270 PAD.n5463 VSS 0.036461f
C5271 PAD.n5464 VSS 0.036461f
C5272 PAD.n5466 VSS 0.036461f
C5273 PAD.n5468 VSS 0.036461f
C5274 PAD.n5470 VSS 0.036461f
C5275 PAD.n5471 VSS 0.036461f
C5276 PAD.n5472 VSS 0.036461f
C5277 PAD.n5473 VSS 0.036461f
C5278 PAD.n5474 VSS 0.036461f
C5279 PAD.n5475 VSS 0.036461f
C5280 PAD.n5476 VSS 0.036461f
C5281 PAD.n5478 VSS 0.036461f
C5282 PAD.n5480 VSS 0.036461f
C5283 PAD.n5482 VSS 0.036461f
C5284 PAD.n5483 VSS 0.036461f
C5285 PAD.n5484 VSS 0.036461f
C5286 PAD.n5485 VSS 0.036461f
C5287 PAD.n5486 VSS 0.036461f
C5288 PAD.n5487 VSS 0.036461f
C5289 PAD.n5488 VSS 0.036461f
C5290 PAD.n5490 VSS 0.036461f
C5291 PAD.n5492 VSS 0.036461f
C5292 PAD.n5494 VSS 0.036461f
C5293 PAD.n5495 VSS 0.036461f
C5294 PAD.n5496 VSS 0.036461f
C5295 PAD.n5497 VSS 0.036461f
C5296 PAD.n5498 VSS 0.036461f
C5297 PAD.n5499 VSS 0.036461f
C5298 PAD.n5500 VSS 0.036461f
C5299 PAD.n5502 VSS 0.036461f
C5300 PAD.n5504 VSS 0.036461f
C5301 PAD.n5506 VSS 0.036461f
C5302 PAD.n5507 VSS 0.036461f
C5303 PAD.n5508 VSS 0.036461f
C5304 PAD.n5509 VSS 0.036461f
C5305 PAD.n5510 VSS 0.036461f
C5306 PAD.n5511 VSS 0.036461f
C5307 PAD.n5512 VSS 0.036461f
C5308 PAD.n5514 VSS 0.036461f
C5309 PAD.n5516 VSS 0.036461f
C5310 PAD.n5518 VSS 0.036461f
C5311 PAD.n5519 VSS 0.036461f
C5312 PAD.n5520 VSS 0.036461f
C5313 PAD.n5521 VSS 0.036461f
C5314 PAD.n5522 VSS 0.036461f
C5315 PAD.n5523 VSS 0.036461f
C5316 PAD.n5524 VSS 0.036461f
C5317 PAD.n5526 VSS 0.036461f
C5318 PAD.n5528 VSS 0.036461f
C5319 PAD.n5530 VSS 0.036461f
C5320 PAD.n5531 VSS 0.036461f
C5321 PAD.n5532 VSS 0.036461f
C5322 PAD.n5533 VSS 0.036461f
C5323 PAD.n5534 VSS 0.036461f
C5324 PAD.n5535 VSS 0.036461f
C5325 PAD.n5536 VSS 0.036461f
C5326 PAD.n5538 VSS 0.036461f
C5327 PAD.n5540 VSS 0.036461f
C5328 PAD.n5541 VSS 0.036461f
C5329 PAD.n5542 VSS 0.023109f
C5330 PAD.n5543 VSS 0.03338f
C5331 PAD.n5544 VSS 0.035657f
C5332 PAD.n5545 VSS 0.03338f
C5333 PAD.n5546 VSS 0.062274f
C5334 PAD.n5547 VSS 0.039761f
C5335 PAD.n5548 VSS 0.069765f
C5336 PAD.n5549 VSS 0.039761f
C5337 PAD.n5550 VSS 0.069765f
C5338 PAD.n5551 VSS 0.527867f
C5339 PAD.n5552 VSS 0.700534f
C5340 PAD.n5553 VSS 0.029436f
C5341 PAD.n5554 VSS 0.048596f
C5342 PAD.n5555 VSS 0.029436f
C5343 PAD.n5556 VSS 0.048596f
C5344 PAD.n5557 VSS 0.030555f
C5345 PAD.n5558 VSS 0.042895f
C5346 PAD.n5559 VSS 0.049115f
C5347 PAD.n5560 VSS 0.049115f
C5348 PAD.n5602 VSS 0.036461f
C5349 PAD.n5604 VSS 0.036461f
C5350 PAD.n5605 VSS 0.036461f
C5351 PAD.n5606 VSS 0.036461f
C5352 PAD.n5607 VSS 0.036461f
C5353 PAD.n5608 VSS 0.036461f
C5354 PAD.n5610 VSS 0.036461f
C5355 PAD.n5611 VSS 0.036461f
C5356 PAD.n5612 VSS 0.036461f
C5357 PAD.n5613 VSS 0.036461f
C5358 PAD.n5615 VSS 0.036461f
C5359 PAD.n5616 VSS 0.036461f
C5360 PAD.n5617 VSS 0.036461f
C5361 PAD.n5618 VSS 0.036461f
C5362 PAD.n5620 VSS 0.036461f
C5363 PAD.n5621 VSS 0.036461f
C5364 PAD.n5622 VSS 0.036461f
C5365 PAD.n5623 VSS 0.036461f
C5366 PAD.n5625 VSS 0.036461f
C5367 PAD.n5626 VSS 0.036461f
C5368 PAD.n5627 VSS 0.036461f
C5369 PAD.n5628 VSS 0.036461f
C5370 PAD.n5630 VSS 0.036461f
C5371 PAD.n5631 VSS 0.036461f
C5372 PAD.n5632 VSS 0.036461f
C5373 PAD.n5633 VSS 0.036461f
C5374 PAD.n5635 VSS 0.036461f
C5375 PAD.n5636 VSS 0.036461f
C5376 PAD.n5637 VSS 0.036461f
C5377 PAD.n5638 VSS 0.036461f
C5378 PAD.n5640 VSS 0.036461f
C5379 PAD.n5641 VSS 0.036461f
C5380 PAD.n5642 VSS 0.036461f
C5381 PAD.n5643 VSS 0.036461f
C5382 PAD.n5645 VSS 0.036461f
C5383 PAD.n5646 VSS 0.036461f
C5384 PAD.n5647 VSS 0.036461f
C5385 PAD.n5648 VSS 0.036461f
C5386 PAD.n5650 VSS 0.036461f
C5387 PAD.n5651 VSS 0.036461f
C5388 PAD.n5652 VSS 0.036461f
C5389 PAD.n5653 VSS 0.036461f
C5390 PAD.n5655 VSS 0.036461f
C5391 PAD.n5656 VSS 0.036461f
C5392 PAD.n5657 VSS 0.036461f
C5393 PAD.n5658 VSS 0.036461f
C5394 PAD.n5660 VSS 0.036461f
C5395 PAD.n5661 VSS 0.036461f
C5396 PAD.n5662 VSS 0.036461f
C5397 PAD.n5663 VSS 0.036461f
C5398 PAD.n5665 VSS 0.036461f
C5399 PAD.n5666 VSS 0.036461f
C5400 PAD.n5667 VSS 0.036461f
C5401 PAD.n5668 VSS 0.036461f
C5402 PAD.n5670 VSS 0.036461f
C5403 PAD.n5671 VSS 0.036461f
C5404 PAD.n5672 VSS 0.036461f
C5405 PAD.n5673 VSS 0.036461f
C5406 PAD.n5675 VSS 0.036461f
C5407 PAD.n5676 VSS 0.036461f
C5408 PAD.n5677 VSS 0.036461f
C5409 PAD.n5678 VSS 0.036461f
C5410 PAD.n5680 VSS 0.036461f
C5411 PAD.n5681 VSS 0.036461f
C5412 PAD.n5682 VSS 0.036461f
C5413 PAD.n5683 VSS 0.036461f
C5414 PAD.n5685 VSS 0.036461f
C5415 PAD.n5686 VSS 0.036461f
C5416 PAD.n5687 VSS 0.036461f
C5417 PAD.n5688 VSS 0.036461f
C5418 PAD.n5690 VSS 0.036461f
C5419 PAD.n5691 VSS 0.036461f
C5420 PAD.n5692 VSS 0.036461f
C5421 PAD.n5693 VSS 0.036461f
C5422 PAD.n5695 VSS 0.036461f
C5423 PAD.n5696 VSS 0.036461f
C5424 PAD.n5697 VSS 0.036461f
C5425 PAD.n5698 VSS 0.036461f
C5426 PAD.n5700 VSS 0.036461f
C5427 PAD.n5701 VSS 0.036461f
C5428 PAD.n5702 VSS 0.023109f
C5429 PAD.n5703 VSS 0.023109f
C5430 PAD.n5704 VSS 0.036461f
C5431 PAD.n5705 VSS 0.036461f
C5432 PAD.n5707 VSS 0.036461f
C5433 PAD.n5708 VSS 0.036461f
C5434 PAD.n5709 VSS 0.036461f
C5435 PAD.n5710 VSS 0.036461f
C5436 PAD.n5711 VSS 0.036461f
C5437 PAD.n5712 VSS 0.036461f
C5438 PAD.n5714 VSS 0.036461f
C5439 PAD.n5715 VSS 0.036461f
C5440 PAD.n5716 VSS 0.036461f
C5441 PAD.n5717 VSS 0.036461f
C5442 PAD.n5718 VSS 0.036461f
C5443 PAD.n5719 VSS 0.036461f
C5444 PAD.n5720 VSS 0.036461f
C5445 PAD.n5721 VSS 0.036461f
C5446 PAD.n5723 VSS 0.036461f
C5447 PAD.n5724 VSS 0.036461f
C5448 PAD.n5725 VSS 0.036461f
C5449 PAD.n5726 VSS 0.036461f
C5450 PAD.n5727 VSS 0.036461f
C5451 PAD.n5728 VSS 0.036461f
C5452 PAD.n5729 VSS 0.036461f
C5453 PAD.n5730 VSS 0.036461f
C5454 PAD.n5732 VSS 0.036461f
C5455 PAD.n5733 VSS 0.036461f
C5456 PAD.n5734 VSS 0.036461f
C5457 PAD.n5735 VSS 0.036461f
C5458 PAD.n5736 VSS 0.036461f
C5459 PAD.n5737 VSS 0.036461f
C5460 PAD.n5738 VSS 0.036461f
C5461 PAD.n5739 VSS 0.036461f
C5462 PAD.n5741 VSS 0.036461f
C5463 PAD.n5742 VSS 0.036461f
C5464 PAD.n5743 VSS 0.036461f
C5465 PAD.n5744 VSS 0.036461f
C5466 PAD.n5745 VSS 0.036461f
C5467 PAD.n5746 VSS 0.036461f
C5468 PAD.n5747 VSS 0.036461f
C5469 PAD.n5748 VSS 0.036461f
C5470 PAD.n5750 VSS 0.036461f
C5471 PAD.n5751 VSS 0.036461f
C5472 PAD.n5752 VSS 0.036461f
C5473 PAD.n5753 VSS 0.036461f
C5474 PAD.n5754 VSS 0.036461f
C5475 PAD.n5755 VSS 0.036461f
C5476 PAD.n5756 VSS 0.036461f
C5477 PAD.n5757 VSS 0.036461f
C5478 PAD.n5759 VSS 0.036461f
C5479 PAD.n5760 VSS 0.036461f
C5480 PAD.n5761 VSS 0.036461f
C5481 PAD.n5762 VSS 0.036461f
C5482 PAD.n5763 VSS 0.036461f
C5483 PAD.n5764 VSS 0.036461f
C5484 PAD.n5765 VSS 0.036461f
C5485 PAD.n5766 VSS 0.036461f
C5486 PAD.n5768 VSS 0.036461f
C5487 PAD.n5769 VSS 0.036461f
C5488 PAD.n5770 VSS 0.036461f
C5489 PAD.n5771 VSS 0.036461f
C5490 PAD.n5772 VSS 0.036461f
C5491 PAD.n5773 VSS 0.036461f
C5492 PAD.n5774 VSS 0.036461f
C5493 PAD.n5775 VSS 0.036461f
C5494 PAD.n5777 VSS 0.036461f
C5495 PAD.n5778 VSS 0.036461f
C5496 PAD.n5779 VSS 0.036461f
C5497 PAD.n5780 VSS 0.036461f
C5498 PAD.n5781 VSS 0.036461f
C5499 PAD.n5782 VSS 0.036461f
C5500 PAD.n5783 VSS 0.036461f
C5501 PAD.n5784 VSS 0.036461f
C5502 PAD.n5786 VSS 0.036461f
C5503 PAD.n5787 VSS 0.036461f
C5504 PAD.n5788 VSS 0.036461f
C5505 PAD.n5789 VSS 0.036461f
C5506 PAD.n5790 VSS 0.036461f
C5507 PAD.n5791 VSS 0.036461f
C5508 PAD.n5792 VSS 0.036461f
C5509 PAD.n5793 VSS 0.036461f
C5510 PAD.n5795 VSS 0.036461f
C5511 PAD.n5796 VSS 0.036461f
C5512 PAD.n5797 VSS 0.036461f
C5513 PAD.n5798 VSS 0.036461f
C5514 PAD.n5799 VSS 0.036461f
C5515 PAD.n5800 VSS 0.036461f
C5516 PAD.n5801 VSS 0.036461f
C5517 PAD.n5802 VSS 0.036461f
C5518 PAD.n5804 VSS 0.036461f
C5519 PAD.n5805 VSS 0.036461f
C5520 PAD.n5806 VSS 0.036461f
C5521 PAD.n5807 VSS 0.036461f
C5522 PAD.n5808 VSS 0.036461f
C5523 PAD.n5809 VSS 0.036461f
C5524 PAD.n5810 VSS 0.036461f
C5525 PAD.n5811 VSS 0.036461f
C5526 PAD.n5813 VSS 0.036461f
C5527 PAD.n5814 VSS 0.036461f
C5528 PAD.n5815 VSS 0.036461f
C5529 PAD.n5816 VSS 0.036461f
C5530 PAD.n5817 VSS 0.036461f
C5531 PAD.n5818 VSS 0.036461f
C5532 PAD.n5819 VSS 0.036461f
C5533 PAD.n5820 VSS 0.036461f
C5534 PAD.n5822 VSS 0.036461f
C5535 PAD.n5823 VSS 0.036461f
C5536 PAD.n5824 VSS 0.036461f
C5537 PAD.n5825 VSS 0.036461f
C5538 PAD.n5826 VSS 0.036461f
C5539 PAD.n5827 VSS 0.036461f
C5540 PAD.n5828 VSS 0.036461f
C5541 PAD.n5829 VSS 0.036461f
C5542 PAD.n5831 VSS 0.036461f
C5543 PAD.n5832 VSS 0.036461f
C5544 PAD.n5833 VSS 0.036461f
C5545 PAD.n5834 VSS 0.036461f
C5546 PAD.n5835 VSS 0.036461f
C5547 PAD.n5836 VSS 0.036461f
C5548 PAD.n5837 VSS 0.036461f
C5549 PAD.n5838 VSS 0.036461f
C5550 PAD.n5840 VSS 0.036461f
C5551 PAD.n5841 VSS 0.036461f
C5552 PAD.n5842 VSS 0.036461f
C5553 PAD.n5843 VSS 0.036461f
C5554 PAD.n5844 VSS 0.036461f
C5555 PAD.n5845 VSS 0.036461f
C5556 PAD.n5846 VSS 0.036461f
C5557 PAD.n5847 VSS 0.036461f
C5558 PAD.n5849 VSS 0.036461f
C5559 PAD.n5850 VSS 0.036461f
C5560 PAD.n5851 VSS 0.036461f
C5561 PAD.n5852 VSS 0.036461f
C5562 PAD.n5853 VSS 0.036461f
C5563 PAD.n5854 VSS 0.036461f
C5564 PAD.n5855 VSS 0.036461f
C5565 PAD.n5856 VSS 0.036461f
C5566 PAD.n5858 VSS 0.036461f
C5567 PAD.n5859 VSS 0.036461f
C5568 PAD.n5860 VSS 0.036461f
C5569 PAD.n5861 VSS 0.036461f
C5570 PAD.n5862 VSS 0.036461f
C5571 PAD.n5863 VSS 0.036461f
C5572 PAD.n5864 VSS 0.036461f
C5573 PAD.n5865 VSS 0.036461f
C5574 PAD.n5867 VSS 0.036461f
C5575 PAD.n5868 VSS 0.036461f
C5576 PAD.n5869 VSS 0.036461f
C5577 PAD.n5870 VSS 0.036461f
C5578 PAD.n5871 VSS 0.036461f
C5579 PAD.n5872 VSS 0.036461f
C5580 PAD.n5873 VSS 0.036461f
C5581 PAD.n5874 VSS 0.036461f
C5582 PAD.n5876 VSS 0.036461f
C5583 PAD.n5877 VSS 0.036461f
C5584 PAD.n5878 VSS 0.036461f
C5585 PAD.n5879 VSS 0.036461f
C5586 PAD.n5880 VSS 0.036461f
C5587 PAD.n5881 VSS 0.036461f
C5588 PAD.n5882 VSS 0.036461f
C5589 PAD.n5883 VSS 0.036461f
C5590 PAD.n5885 VSS 0.036461f
C5591 PAD.n5886 VSS 0.036461f
C5592 PAD.n5887 VSS 0.036461f
C5593 PAD.n5888 VSS 0.036461f
C5594 PAD.n5889 VSS 0.036461f
C5595 PAD.n5890 VSS 0.036461f
C5596 PAD.n5891 VSS 0.023109f
C5597 PAD.n5892 VSS 0.023109f
C5598 PAD.n5894 VSS 0.611735f
C5599 PAD.n5895 VSS 0.069765f
C5600 PAD.n5896 VSS 0.06639f
C5601 PAD.n5897 VSS 0.03415f
C5602 PAD.n5898 VSS 0.036461f
C5603 PAD.n5899 VSS 0.039761f
C5604 PAD.n5900 VSS 0.036461f
C5605 PAD.n5901 VSS 0.039761f
C5606 PAD.n5903 VSS 0.582134f
C5607 PAD.n5904 VSS 0.300934f
C5608 PAD.n5905 VSS 0.036461f
C5609 PAD.n5948 VSS 0.029436f
C5610 PAD.n5949 VSS 0.036461f
C5611 PAD.n5950 VSS 0.036461f
C5612 PAD.n5951 VSS 0.030555f
C5613 PAD.n5952 VSS 0.033032f
C5614 PAD.n5953 VSS 0.035494f
C5615 PAD.n5954 VSS 0.069765f
C5616 PAD.n5955 VSS 0.063576f
C5617 PAD.n5956 VSS 0.128786f
C5618 PAD.n5957 VSS 0.103613f
C5619 PAD.n5958 VSS 0.066152f
C5620 PAD.n5959 VSS 0.103613f
C5621 PAD.n5960 VSS 0.066152f
C5622 PAD.n5962 VSS 0.611735f
C5623 PAD.n5963 VSS 0.611735f
C5624 PAD.n5964 VSS 0.611735f
C5625 PAD.n5965 VSS 0.611735f
C5626 PAD.n5966 VSS 0.651201f
C5627 PAD.n5967 VSS 0.069176f
C5628 PAD.n5968 VSS 0.069176f
C5629 PAD.n5969 VSS 0.103613f
C5630 PAD.n5970 VSS 0.063576f
C5631 PAD.n5971 VSS 0.700534f
C5632 PAD.n5972 VSS 0.042473f
C5633 PAD.n5973 VSS 0.033032f
C5634 PAD.n5974 VSS 0.611734f
C5635 PAD.n5975 VSS 0.049115f
C5636 PAD.n5976 VSS 0.042473f
C5637 PAD.n5977 VSS 0.049115f
C5638 PAD.n5978 VSS 0.06827f
C5639 PAD.n5979 VSS 0.611735f
C5640 PAD.n5980 VSS 0.611735f
C5641 PAD.n5981 VSS 0.611735f
C5642 PAD.n5982 VSS 0.611735f
C5643 PAD.n5983 VSS 0.074916f
C5644 PAD.n5984 VSS 0.074916f
C5645 PAD.n5985 VSS 0.074916f
C5646 PAD.n5986 VSS 0.074916f
C5647 PAD.n5987 VSS 0.074916f
C5648 PAD.n5988 VSS 0.074916f
C5649 PAD.n5989 VSS 0.074916f
C5650 PAD.n5990 VSS 0.074916f
C5651 PAD.n5991 VSS 0.074916f
C5652 PAD.n5992 VSS 0.074916f
C5653 PAD.n5993 VSS 0.074916f
C5654 PAD.n5994 VSS 0.074916f
C5655 PAD.n5995 VSS 0.074916f
C5656 PAD.n5996 VSS 0.074916f
C5657 PAD.n5997 VSS 0.074916f
C5658 PAD.n5998 VSS 0.074916f
C5659 PAD.n5999 VSS 0.074916f
C5660 PAD.n6000 VSS 0.074916f
C5661 PAD.n6001 VSS 0.074916f
C5662 PAD.n6002 VSS 0.074916f
C5663 PAD.n6003 VSS 0.074916f
C5664 PAD.n6004 VSS 0.074916f
C5665 PAD.n6005 VSS 0.074916f
C5666 PAD.n6006 VSS 0.074916f
C5667 PAD.n6007 VSS 0.074916f
C5668 PAD.n6008 VSS 0.074916f
C5669 PAD.n6009 VSS 0.074916f
C5670 PAD.n6010 VSS 0.074916f
C5671 PAD.n6011 VSS 0.074916f
C5672 PAD.n6012 VSS 0.074916f
C5673 PAD.n6013 VSS 0.074916f
C5674 PAD.n6014 VSS 0.074916f
C5675 PAD.n6015 VSS 0.074916f
C5676 PAD.n6016 VSS 0.074916f
C5677 PAD.n6017 VSS 0.074916f
C5678 PAD.n6018 VSS 0.074916f
C5679 PAD.n6019 VSS 0.074916f
C5680 PAD.n6020 VSS 0.074916f
C5681 PAD.n6021 VSS 0.074916f
C5682 PAD.n6022 VSS 0.074916f
C5683 PAD.n6023 VSS 0.074916f
C5684 PAD.n6024 VSS 0.074916f
C5685 PAD.n6025 VSS 0.074916f
C5686 PAD.n6026 VSS 0.074916f
C5687 PAD.n6027 VSS 0.074916f
C5688 PAD.n6028 VSS 0.074916f
C5689 PAD.n6029 VSS 0.074916f
C5690 PAD.n6030 VSS 0.074916f
C5691 PAD.n6032 VSS 0.074916f
C5692 PAD.n6034 VSS 0.103613f
C5693 PAD.n6037 VSS 0.074916f
C5694 PAD.n6040 VSS 0.074916f
C5695 PAD.n6043 VSS 0.074916f
C5696 PAD.n6046 VSS 0.074916f
C5697 PAD.n6049 VSS 0.074916f
C5698 PAD.n6052 VSS 0.074916f
C5699 PAD.n6055 VSS 0.074916f
C5700 PAD.n6058 VSS 0.074916f
C5701 PAD.n6061 VSS 0.074916f
C5702 PAD.n6064 VSS 0.074916f
C5703 PAD.n6067 VSS 0.074916f
C5704 PAD.n6070 VSS 0.074916f
C5705 PAD.n6073 VSS 0.074916f
C5706 PAD.n6076 VSS 0.074916f
C5707 PAD.n6079 VSS 0.074916f
C5708 PAD.n6082 VSS 0.074916f
C5709 PAD.n6085 VSS 0.074916f
C5710 PAD.n6088 VSS 0.074916f
C5711 PAD.n6091 VSS 0.074916f
C5712 PAD.n6094 VSS 0.074916f
C5713 PAD.n6097 VSS 0.074916f
C5714 PAD.n6100 VSS 0.074916f
C5715 PAD.n6103 VSS 0.074916f
C5716 PAD.n6106 VSS 0.074916f
C5717 PAD.n6109 VSS 0.074916f
C5718 PAD.n6112 VSS 0.074916f
C5719 PAD.n6115 VSS 0.074916f
C5720 PAD.n6118 VSS 0.074916f
C5721 PAD.n6121 VSS 0.074916f
C5722 PAD.n6124 VSS 0.074916f
C5723 PAD.n6127 VSS 0.074916f
C5724 PAD.n6130 VSS 0.074916f
C5725 PAD.n6133 VSS 0.074916f
C5726 PAD.n6136 VSS 0.074916f
C5727 PAD.n6139 VSS 0.074916f
C5728 PAD.n6142 VSS 0.074916f
C5729 PAD.n6145 VSS 0.074916f
C5730 PAD.n6148 VSS 0.074916f
C5731 PAD.n6151 VSS 0.074916f
C5732 PAD.n6154 VSS 0.074916f
C5733 PAD.n6157 VSS 0.074916f
C5734 PAD.n6160 VSS 0.074916f
C5735 PAD.n6163 VSS 0.074916f
C5736 PAD.n6166 VSS 0.074916f
C5737 PAD.n6169 VSS 0.074916f
C5738 PAD.n6172 VSS 0.074916f
C5739 PAD.n6175 VSS 0.074916f
C5740 PAD.n6177 VSS 0.074916f
C5741 PAD.n6178 VSS 0.074916f
C5742 PAD.n6179 VSS 0.074916f
C5743 PAD.n6180 VSS 0.074916f
C5744 PAD.n6181 VSS 0.074916f
C5745 PAD.n6182 VSS 0.074916f
C5746 PAD.n6183 VSS 0.074916f
C5747 PAD.n6184 VSS 0.074916f
C5748 PAD.n6185 VSS 0.074916f
C5749 PAD.n6186 VSS 0.074916f
C5750 PAD.n6187 VSS 0.074916f
C5751 PAD.n6188 VSS 0.074916f
C5752 PAD.n6189 VSS 0.074916f
C5753 PAD.n6190 VSS 0.074916f
C5754 PAD.n6191 VSS 0.074916f
C5755 PAD.n6192 VSS 0.074916f
C5756 PAD.n6193 VSS 0.074916f
C5757 PAD.n6194 VSS 0.074916f
C5758 PAD.n6195 VSS 0.074916f
C5759 PAD.n6196 VSS 0.074916f
C5760 PAD.n6197 VSS 0.074916f
C5761 PAD.n6198 VSS 0.074916f
C5762 PAD.n6199 VSS 0.074916f
C5763 PAD.n6200 VSS 0.074916f
C5764 PAD.n6201 VSS 0.074916f
C5765 PAD.n6202 VSS 0.074916f
C5766 PAD.n6203 VSS 0.074916f
C5767 PAD.n6204 VSS 0.074916f
C5768 PAD.n6205 VSS 0.074916f
C5769 PAD.n6206 VSS 0.074916f
C5770 PAD.n6207 VSS 0.074916f
C5771 PAD.n6208 VSS 0.074916f
C5772 PAD.n6209 VSS 0.074916f
C5773 PAD.n6210 VSS 0.074916f
C5774 PAD.n6211 VSS 0.074916f
C5775 PAD.n6212 VSS 0.074916f
C5776 PAD.n6213 VSS 0.074916f
C5777 PAD.n6214 VSS 0.074916f
C5778 PAD.n6215 VSS 0.074916f
C5779 PAD.n6216 VSS 0.074916f
C5780 PAD.n6217 VSS 0.074916f
C5781 PAD.n6218 VSS 0.074916f
C5782 PAD.n6219 VSS 0.074916f
C5783 PAD.n6220 VSS 0.074916f
C5784 PAD.n6221 VSS 0.074916f
C5785 PAD.n6222 VSS 0.074916f
C5786 PAD.n6223 VSS 0.074916f
C5787 PAD.n6224 VSS 0.074916f
C5788 PAD.n6225 VSS 0.103613f
C5789 PAD.n6226 VSS 0.103613f
C5790 PAD.n6227 VSS 0.074916f
C5791 PAD.n6228 VSS 0.074916f
C5792 PAD.n6229 VSS 0.074916f
C5793 PAD.n6230 VSS 0.074916f
C5794 PAD.n6231 VSS 0.074916f
C5795 PAD.n6232 VSS 0.074916f
C5796 PAD.n6233 VSS 0.074916f
C5797 PAD.n6234 VSS 0.074916f
C5798 PAD.n6235 VSS 0.074916f
C5799 PAD.n6236 VSS 0.074916f
C5800 PAD.n6237 VSS 0.074916f
C5801 PAD.n6238 VSS 0.074916f
C5802 PAD.n6239 VSS 0.074916f
C5803 PAD.n6240 VSS 0.074916f
C5804 PAD.n6241 VSS 0.074916f
C5805 PAD.n6242 VSS 0.074916f
C5806 PAD.n6243 VSS 0.074916f
C5807 PAD.n6244 VSS 0.074916f
C5808 PAD.n6245 VSS 0.074916f
C5809 PAD.n6246 VSS 0.074916f
C5810 PAD.n6247 VSS 0.074916f
C5811 PAD.n6248 VSS 0.074916f
C5812 PAD.n6249 VSS 0.074916f
C5813 PAD.n6250 VSS 0.074916f
C5814 PAD.n6251 VSS 0.074916f
C5815 PAD.n6252 VSS 0.074916f
C5816 PAD.n6253 VSS 0.074916f
C5817 PAD.n6254 VSS 0.074916f
C5818 PAD.n6255 VSS 0.074916f
C5819 PAD.n6256 VSS 0.074916f
C5820 PAD.n6257 VSS 0.074916f
C5821 PAD.n6258 VSS 0.074916f
C5822 PAD.n6259 VSS 0.074916f
C5823 PAD.n6260 VSS 0.074916f
C5824 PAD.n6261 VSS 0.074916f
C5825 PAD.n6262 VSS 0.074916f
C5826 PAD.n6263 VSS 0.074916f
C5827 PAD.n6264 VSS 0.074916f
C5828 PAD.n6265 VSS 0.074916f
C5829 PAD.n6266 VSS 0.074916f
C5830 PAD.n6267 VSS 0.074916f
C5831 PAD.n6268 VSS 0.074916f
C5832 PAD.n6269 VSS 0.074916f
C5833 PAD.n6270 VSS 0.074916f
C5834 PAD.n6271 VSS 0.074916f
C5835 PAD.n6272 VSS 0.074916f
C5836 PAD.n6273 VSS 0.074916f
C5837 PAD.n6274 VSS 0.074916f
C5838 PAD.n6275 VSS 0.074916f
C5839 PAD.n6276 VSS 0.074916f
C5840 PAD.n6277 VSS 0.074916f
C5841 PAD.n6278 VSS 0.074916f
C5842 PAD.n6279 VSS 0.074916f
C5843 PAD.n6280 VSS 0.074916f
C5844 PAD.n6281 VSS 0.074916f
C5845 PAD.n6282 VSS 0.074916f
C5846 PAD.n6283 VSS 0.074916f
C5847 PAD.n6284 VSS 0.074916f
C5848 PAD.n6285 VSS 0.074916f
C5849 PAD.n6286 VSS 0.074916f
C5850 PAD.n6287 VSS 0.074916f
C5851 PAD.n6288 VSS 0.074916f
C5852 PAD.n6289 VSS 0.074916f
C5853 PAD.n6290 VSS 0.074916f
C5854 PAD.n6291 VSS 0.074916f
C5855 PAD.n6292 VSS 0.074916f
C5856 PAD.n6293 VSS 0.074916f
C5857 PAD.n6294 VSS 0.074916f
C5858 PAD.n6295 VSS 0.074916f
C5859 PAD.n6296 VSS 0.074916f
C5860 PAD.n6297 VSS 0.074916f
C5861 PAD.n6298 VSS 0.074916f
C5862 PAD.n6299 VSS 0.074916f
C5863 PAD.n6300 VSS 0.074916f
C5864 PAD.n6301 VSS 0.074916f
C5865 PAD.n6302 VSS 0.074916f
C5866 PAD.n6303 VSS 0.074916f
C5867 PAD.n6304 VSS 0.074916f
C5868 PAD.n6305 VSS 0.074916f
C5869 PAD.n6306 VSS 0.074916f
C5870 PAD.n6307 VSS 0.074916f
C5871 PAD.n6308 VSS 0.074916f
C5872 PAD.n6309 VSS 0.074916f
C5873 PAD.n6310 VSS 0.074916f
C5874 PAD.n6311 VSS 0.074916f
C5875 PAD.n6312 VSS 0.074916f
C5876 PAD.n6313 VSS 0.074916f
C5877 PAD.n6314 VSS 0.074916f
C5878 PAD.n6315 VSS 0.074916f
C5879 PAD.n6316 VSS 0.074916f
C5880 PAD.n6317 VSS 0.074916f
C5881 PAD.n6318 VSS 0.074916f
C5882 PAD.n6319 VSS 0.074916f
C5883 PAD.n6320 VSS 0.074916f
C5884 PAD.n6321 VSS 0.074916f
C5885 PAD.n6322 VSS 0.074916f
C5886 PAD.n6323 VSS 0.074916f
C5887 PAD.n6324 VSS 0.074916f
C5888 PAD.n6325 VSS 0.074916f
C5889 PAD.n6326 VSS 0.074916f
C5890 PAD.n6327 VSS 0.074916f
C5891 PAD.n6328 VSS 0.074916f
C5892 PAD.n6329 VSS 0.074916f
C5893 PAD.n6330 VSS 0.074916f
C5894 PAD.n6331 VSS 0.074916f
C5895 PAD.n6332 VSS 0.074916f
C5896 PAD.n6333 VSS 0.074916f
C5897 PAD.n6334 VSS 0.074916f
C5898 PAD.n6335 VSS 0.074916f
C5899 PAD.n6336 VSS 0.074916f
C5900 PAD.n6337 VSS 0.074916f
C5901 PAD.n6338 VSS 0.074916f
C5902 PAD.n6339 VSS 0.074916f
C5903 PAD.n6340 VSS 0.074916f
C5904 PAD.n6341 VSS 0.074916f
C5905 PAD.n6342 VSS 0.074916f
C5906 PAD.n6343 VSS 0.074916f
C5907 PAD.n6344 VSS 0.074916f
C5908 PAD.n6345 VSS 0.074916f
C5909 PAD.n6346 VSS 0.074916f
C5910 PAD.n6347 VSS 0.074916f
C5911 PAD.n6348 VSS 0.074916f
C5912 PAD.n6349 VSS 0.074916f
C5913 PAD.n6350 VSS 0.074916f
C5914 PAD.n6351 VSS 0.074916f
C5915 PAD.n6352 VSS 0.074916f
C5916 PAD.n6353 VSS 0.074916f
C5917 PAD.n6354 VSS 0.074916f
C5918 PAD.n6355 VSS 0.074916f
C5919 PAD.n6356 VSS 0.074916f
C5920 PAD.n6357 VSS 0.074916f
C5921 PAD.n6358 VSS 0.074916f
C5922 PAD.n6359 VSS 0.074916f
C5923 PAD.n6360 VSS 0.074916f
C5924 PAD.n6361 VSS 0.074916f
C5925 PAD.n6362 VSS 0.074916f
C5926 PAD.n6363 VSS 0.074916f
C5927 PAD.n6364 VSS 0.074916f
C5928 PAD.n6365 VSS 0.074916f
C5929 PAD.n6366 VSS 0.074916f
C5930 PAD.n6367 VSS 0.074916f
C5931 PAD.n6368 VSS 0.074916f
C5932 PAD.n6369 VSS 0.074916f
C5933 PAD.n6370 VSS 0.074916f
C5934 PAD.n6371 VSS 0.05951f
C5935 PAD.n6372 VSS 0.05951f
C5936 PAD.n6373 VSS 1.51947f
C5937 PAD.n6374 VSS 0.122947f
C5938 PAD.n6375 VSS 0.12326f
C5939 PAD.n6376 VSS 0.155711f
C5940 PAD.n6377 VSS 0.033773f
C5941 PAD.n6378 VSS 0.028849f
C5942 PAD.n6379 VSS 0.042895f
C5943 PAD.n6380 VSS 0.025828f
C5944 PAD.n6381 VSS 0.029573f
C5945 PAD.n6382 VSS 0.029573f
C5946 PAD.n6383 VSS 0.611734f
C5947 PAD.n6385 VSS 0.125825f
C5948 PAD.n6386 VSS 0.863335f
C5949 PAD.n6387 VSS 0.043197f
C5950 PAD.n6388 VSS 0.043197f
C5951 PAD.n6389 VSS 0.055281f
C5952 PAD.n6390 VSS 0.238924f
C5953 PAD.n6391 VSS 0.05675f
C5954 PAD.n6392 VSS 0.062274f
C5955 PAD.n6393 VSS 0.069765f
C5956 PAD.n6394 VSS 0.038258f
C5957 PAD.n6395 VSS 0.038258f
C5958 PAD.n6396 VSS 0.582134f
C5959 PAD.n6436 VSS 0.036461f
C5960 PAD.n6437 VSS 0.036461f
C5961 PAD.n6438 VSS 0.036461f
C5962 PAD.n6439 VSS 0.036461f
C5963 PAD.n6440 VSS 0.036461f
C5964 PAD.n6441 VSS 0.036461f
C5965 PAD.n6442 VSS 0.036461f
C5966 PAD.n6443 VSS 0.036461f
C5967 PAD.n6444 VSS 0.036461f
C5968 PAD.n6445 VSS 0.036461f
C5969 PAD.n6446 VSS 0.036461f
C5970 PAD.n6447 VSS 0.036461f
C5971 PAD.n6448 VSS 0.036461f
C5972 PAD.n6449 VSS 0.036461f
C5973 PAD.n6450 VSS 0.036461f
C5974 PAD.n6451 VSS 0.036461f
C5975 PAD.n6452 VSS 0.036461f
C5976 PAD.n6453 VSS 0.036461f
C5977 PAD.n6454 VSS 0.036461f
C5978 PAD.n6455 VSS 0.036461f
C5979 PAD.n6456 VSS 0.036461f
C5980 PAD.n6457 VSS 0.036461f
C5981 PAD.n6458 VSS 0.036461f
C5982 PAD.n6459 VSS 0.036461f
C5983 PAD.n6460 VSS 0.036461f
C5984 PAD.n6461 VSS 0.036461f
C5985 PAD.n6462 VSS 0.036461f
C5986 PAD.n6463 VSS 0.036461f
C5987 PAD.n6464 VSS 0.036461f
C5988 PAD.n6465 VSS 0.036461f
C5989 PAD.n6466 VSS 0.036461f
C5990 PAD.n6467 VSS 0.036461f
C5991 PAD.n6468 VSS 0.036461f
C5992 PAD.n6469 VSS 0.036461f
C5993 PAD.n6470 VSS 0.036461f
C5994 PAD.n6471 VSS 0.036461f
C5995 PAD.n6472 VSS 0.036461f
C5996 PAD.n6473 VSS 0.036461f
C5997 PAD.n6474 VSS 0.036461f
C5998 PAD.n6475 VSS 0.036461f
C5999 PAD.n6476 VSS 0.036461f
C6000 PAD.n6477 VSS 0.036461f
C6001 PAD.n6478 VSS 0.036461f
C6002 PAD.n6479 VSS 0.036461f
C6003 PAD.n6480 VSS 0.036461f
C6004 PAD.n6481 VSS 0.036461f
C6005 PAD.n6482 VSS 0.036461f
C6006 PAD.n6483 VSS 0.036461f
C6007 PAD.n6484 VSS 0.036461f
C6008 PAD.n6485 VSS 0.036461f
C6009 PAD.n6486 VSS 0.036461f
C6010 PAD.n6487 VSS 0.036461f
C6011 PAD.n6488 VSS 0.036461f
C6012 PAD.n6489 VSS 0.036461f
C6013 PAD.n6490 VSS 0.036461f
C6014 PAD.n6491 VSS 0.036461f
C6015 PAD.n6492 VSS 0.036461f
C6016 PAD.n6493 VSS 0.036461f
C6017 PAD.n6494 VSS 0.036461f
C6018 PAD.n6495 VSS 0.036461f
C6019 PAD.n6496 VSS 0.036461f
C6020 PAD.n6497 VSS 0.036461f
C6021 PAD.n6498 VSS 0.036461f
C6022 PAD.n6499 VSS 0.036461f
C6023 PAD.n6500 VSS 0.036461f
C6024 PAD.n6501 VSS 0.036461f
C6025 PAD.n6502 VSS 0.036461f
C6026 PAD.n6503 VSS 0.036461f
C6027 PAD.n6504 VSS 0.036461f
C6028 PAD.n6505 VSS 0.036461f
C6029 PAD.n6506 VSS 0.036461f
C6030 PAD.n6507 VSS 0.036461f
C6031 PAD.n6508 VSS 0.036461f
C6032 PAD.n6509 VSS 0.036461f
C6033 PAD.n6510 VSS 0.036461f
C6034 PAD.n6511 VSS 0.036461f
C6035 PAD.n6512 VSS 0.036461f
C6036 PAD.n6513 VSS 0.036461f
C6037 PAD.n6514 VSS 0.036461f
C6038 PAD.n6515 VSS 0.036461f
C6039 PAD.n6516 VSS 0.036461f
C6040 PAD.n6517 VSS 0.036461f
C6041 PAD.n6518 VSS 0.036461f
C6042 PAD.n6519 VSS 0.036461f
C6043 PAD.n6520 VSS 0.036461f
C6044 PAD.n6521 VSS 0.036461f
C6045 PAD.n6522 VSS 0.036461f
C6046 PAD.n6523 VSS 0.036461f
C6047 PAD.n6524 VSS 0.036461f
C6048 PAD.n6525 VSS 0.036461f
C6049 PAD.n6526 VSS 0.036461f
C6050 PAD.n6527 VSS 0.036461f
C6051 PAD.n6528 VSS 0.036461f
C6052 PAD.n6529 VSS 0.036461f
C6053 PAD.n6530 VSS 0.036461f
C6054 PAD.n6531 VSS 0.036461f
C6055 PAD.n6532 VSS 0.036461f
C6056 PAD.n6533 VSS 0.036461f
C6057 PAD.n6534 VSS 0.036461f
C6058 PAD.n6535 VSS 0.036461f
C6059 PAD.n6536 VSS 0.036461f
C6060 PAD.n6537 VSS 0.036461f
C6061 PAD.n6538 VSS 0.036461f
C6062 PAD.n6539 VSS 0.036461f
C6063 PAD.n6540 VSS 0.036461f
C6064 PAD.n6541 VSS 0.036461f
C6065 PAD.n6542 VSS 0.036461f
C6066 PAD.n6543 VSS 0.036461f
C6067 PAD.n6544 VSS 0.036461f
C6068 PAD.n6545 VSS 0.036461f
C6069 PAD.n6546 VSS 0.036461f
C6070 PAD.n6547 VSS 0.036461f
C6071 PAD.n6548 VSS 0.036461f
C6072 PAD.n6549 VSS 0.036461f
C6073 PAD.n6550 VSS 0.036461f
C6074 PAD.n6551 VSS 0.036461f
C6075 PAD.n6552 VSS 0.036461f
C6076 PAD.n6553 VSS 0.036461f
C6077 PAD.n6554 VSS 0.036461f
C6078 PAD.n6555 VSS 0.036461f
C6079 PAD.n6556 VSS 0.036461f
C6080 PAD.n6557 VSS 0.036461f
C6081 PAD.n6558 VSS 0.036461f
C6082 PAD.n6559 VSS 0.036461f
C6083 PAD.n6560 VSS 0.036461f
C6084 PAD.n6561 VSS 0.036461f
C6085 PAD.n6562 VSS 0.036461f
C6086 PAD.n6563 VSS 0.036461f
C6087 PAD.n6564 VSS 0.036461f
C6088 PAD.n6565 VSS 0.036461f
C6089 PAD.n6566 VSS 0.036461f
C6090 PAD.n6567 VSS 0.036461f
C6091 PAD.n6568 VSS 0.036461f
C6092 PAD.n6569 VSS 0.036461f
C6093 PAD.n6570 VSS 0.036461f
C6094 PAD.n6571 VSS 0.036461f
C6095 PAD.n6572 VSS 0.036461f
C6096 PAD.n6573 VSS 0.036461f
C6097 PAD.n6574 VSS 0.036461f
C6098 PAD.n6575 VSS 0.036461f
C6099 PAD.n6576 VSS 0.036461f
C6100 PAD.n6577 VSS 0.036461f
C6101 PAD.n6578 VSS 0.036461f
C6102 PAD.n6579 VSS 0.036461f
C6103 PAD.n6580 VSS 0.036461f
C6104 PAD.n6581 VSS 0.036461f
C6105 PAD.n6582 VSS 0.036461f
C6106 PAD.n6583 VSS 0.036461f
C6107 PAD.n6584 VSS 0.036461f
C6108 PAD.n6585 VSS 0.036461f
C6109 PAD.n6586 VSS 0.036461f
C6110 PAD.n6587 VSS 0.036461f
C6111 PAD.n6588 VSS 0.036461f
C6112 PAD.n6589 VSS 0.036461f
C6113 PAD.n6590 VSS 0.036461f
C6114 PAD.n6591 VSS 0.036461f
C6115 PAD.n6592 VSS 0.036461f
C6116 PAD.n6593 VSS 0.036461f
C6117 PAD.n6594 VSS 0.036461f
C6118 PAD.n6595 VSS 0.036461f
C6119 PAD.n6596 VSS 0.036461f
C6120 PAD.n6597 VSS 0.036461f
C6121 PAD.n6598 VSS 0.036461f
C6122 PAD.n6599 VSS 0.036461f
C6123 PAD.n6600 VSS 0.036461f
C6124 PAD.n6601 VSS 0.036461f
C6125 PAD.n6602 VSS 0.036461f
C6126 PAD.n6603 VSS 0.036461f
C6127 PAD.n6604 VSS 0.036461f
C6128 PAD.n6605 VSS 0.036461f
C6129 PAD.n6606 VSS 0.036461f
C6130 PAD.n6607 VSS 0.036461f
C6131 PAD.n6608 VSS 0.036461f
C6132 PAD.n6609 VSS 0.036461f
C6133 PAD.n6610 VSS 0.036461f
C6134 PAD.n6611 VSS 0.036461f
C6135 PAD.n6612 VSS 0.036461f
C6136 PAD.n6613 VSS 0.036461f
C6137 PAD.n6614 VSS 0.036461f
C6138 PAD.n6615 VSS 0.036461f
C6139 PAD.n6616 VSS 0.036461f
C6140 PAD.n6617 VSS 0.036461f
C6141 PAD.n6618 VSS 0.036461f
C6142 PAD.n6619 VSS 0.036461f
C6143 PAD.n6620 VSS 0.036461f
C6144 PAD.n6621 VSS 0.036461f
C6145 PAD.n6622 VSS 0.036461f
C6146 PAD.n6623 VSS 0.036461f
C6147 PAD.n6624 VSS 0.036461f
C6148 PAD.n6625 VSS 0.036461f
C6149 PAD.n6626 VSS 0.036461f
C6150 PAD.n6627 VSS 0.036461f
C6151 PAD.n6628 VSS 0.036461f
C6152 PAD.n6629 VSS 0.036461f
C6153 PAD.n6630 VSS 0.036461f
C6154 PAD.n6631 VSS 0.036461f
C6155 PAD.n6632 VSS 0.036461f
C6156 PAD.n6633 VSS 0.036461f
C6157 PAD.n6634 VSS 0.036461f
C6158 PAD.n6635 VSS 0.036461f
C6159 PAD.n6636 VSS 0.036461f
C6160 PAD.n6637 VSS 0.036461f
C6161 PAD.n6638 VSS 0.036461f
C6162 PAD.n6639 VSS 0.036461f
C6163 PAD.n6640 VSS 0.036461f
C6164 PAD.n6641 VSS 0.036461f
C6165 PAD.n6642 VSS 0.036461f
C6166 PAD.n6643 VSS 0.036461f
C6167 PAD.n6644 VSS 0.036461f
C6168 PAD.n6645 VSS 0.036461f
C6169 PAD.n6646 VSS 0.036461f
C6170 PAD.n6647 VSS 0.036461f
C6171 PAD.n6648 VSS 0.036461f
C6172 PAD.n6649 VSS 0.036461f
C6173 PAD.n6650 VSS 0.036461f
C6174 PAD.n6651 VSS 0.036461f
C6175 PAD.n6652 VSS 0.036461f
C6176 PAD.n6653 VSS 0.036461f
C6177 PAD.n6654 VSS 0.036461f
C6178 PAD.n6655 VSS 0.036461f
C6179 PAD.n6656 VSS 0.036461f
C6180 PAD.n6657 VSS 0.036461f
C6181 PAD.n6658 VSS 0.036461f
C6182 PAD.n6659 VSS 0.036461f
C6183 PAD.n6660 VSS 0.036461f
C6184 PAD.n6661 VSS 0.036461f
C6185 PAD.n6662 VSS 0.036461f
C6186 PAD.n6663 VSS 0.036461f
C6187 PAD.n6664 VSS 0.036461f
C6188 PAD.n6665 VSS 0.036461f
C6189 PAD.n6666 VSS 0.036461f
C6190 PAD.n6667 VSS 0.036461f
C6191 PAD.n6668 VSS 0.036461f
C6192 PAD.n6669 VSS 0.036461f
C6193 PAD.n6670 VSS 0.036461f
C6194 PAD.n6671 VSS 0.036461f
C6195 PAD.n6672 VSS 0.036461f
C6196 PAD.n6673 VSS 0.036461f
C6197 PAD.n6674 VSS 0.036461f
C6198 PAD.n6675 VSS 0.036461f
C6199 PAD.n6676 VSS 0.036461f
C6200 PAD.n6678 VSS 0.518001f
C6201 PAD.n6679 VSS 0.478534f
C6202 PAD.n6680 VSS 0.611734f
C6203 PAD.n6681 VSS 0.06639f
C6204 PAD.n6682 VSS 0.700534f
C6205 PAD.n6683 VSS 0.212133f
C6206 PAD.n6684 VSS 0.040641f
C6207 PAD.n6685 VSS 0.040641f
C6208 PAD.n6686 VSS 0.029436f
C6209 PAD.n6687 VSS 0.023109f
C6210 PAD.n6688 VSS 0.023109f
C6211 PAD.n6689 VSS 0.429201f
C6212 PAD.n6690 VSS 0.023109f
C6213 PAD.n6691 VSS 0.023109f
C6214 PAD.n6692 VSS 0.03338f
C6215 PAD.n6693 VSS 0.046286f
C6216 PAD.n6694 VSS 0.059261f
C6217 PAD.n6695 VSS 0.062274f
C6218 PAD.n6696 VSS 0.069765f
C6219 PAD.n6697 VSS 0.046135f
C6220 PAD.n6698 VSS 0.046135f
C6221 PAD.n6699 VSS 0.222f
C6222 PAD.n6700 VSS 0.562401f
C6223 PAD.n6701 VSS 0.028535f
C6224 PAD.n6702 VSS 0.028535f
C6225 PAD.n6703 VSS 0.024922f
C6226 PAD.n6704 VSS 0.033773f
C6227 PAD.n6705 VSS 0.030555f
C6228 PAD.n6706 VSS 0.042895f
C6229 PAD.n6707 VSS 0.029436f
C6230 PAD.n6708 VSS 0.049115f
C6231 PAD.n6709 VSS 0.029436f
C6232 PAD.n6710 VSS 0.049115f
C6233 PAD.n6711 VSS 0.611734f
C6234 PAD.n6712 VSS 0.700534f
C6235 PAD.n6713 VSS 0.439067f
C6236 PAD.n6714 VSS 0.039761f
C6237 PAD.n6715 VSS 0.069765f
C6238 PAD.n6716 VSS 0.039761f
C6239 PAD.n6717 VSS 0.069765f
C6240 PAD.n6718 VSS 0.036461f
C6241 PAD.n6719 VSS 0.023109f
C6242 PAD.n6720 VSS 0.036461f
C6243 PAD.n6723 VSS 0.036461f
C6244 PAD.n6724 VSS 0.036461f
C6245 PAD.n6725 VSS 0.036461f
C6246 PAD.n6726 VSS 0.036461f
C6247 PAD.n6728 VSS 0.036461f
C6248 PAD.n6729 VSS 0.036461f
C6249 PAD.n6730 VSS 0.036461f
C6250 PAD.n6732 VSS 0.036461f
C6251 PAD.n6733 VSS 0.036461f
C6252 PAD.n6734 VSS 0.036461f
C6253 PAD.n6736 VSS 0.036461f
C6254 PAD.n6737 VSS 0.036461f
C6255 PAD.n6738 VSS 0.036461f
C6256 PAD.n6740 VSS 0.036461f
C6257 PAD.n6741 VSS 0.036461f
C6258 PAD.n6742 VSS 0.036461f
C6259 PAD.n6744 VSS 0.036461f
C6260 PAD.n6745 VSS 0.036461f
C6261 PAD.n6746 VSS 0.036461f
C6262 PAD.n6748 VSS 0.036461f
C6263 PAD.n6749 VSS 0.036461f
C6264 PAD.n6750 VSS 0.036461f
C6265 PAD.n6752 VSS 0.036461f
C6266 PAD.n6753 VSS 0.036461f
C6267 PAD.n6754 VSS 0.036461f
C6268 PAD.n6756 VSS 0.036461f
C6269 PAD.n6757 VSS 0.036461f
C6270 PAD.n6758 VSS 0.036461f
C6271 PAD.n6760 VSS 0.036461f
C6272 PAD.n6761 VSS 0.036461f
C6273 PAD.n6762 VSS 0.036461f
C6274 PAD.n6764 VSS 0.036461f
C6275 PAD.n6765 VSS 0.036461f
C6276 PAD.n6766 VSS 0.036461f
C6277 PAD.n6768 VSS 0.036461f
C6278 PAD.n6769 VSS 0.036461f
C6279 PAD.n6770 VSS 0.036461f
C6280 PAD.n6772 VSS 0.036461f
C6281 PAD.n6773 VSS 0.036461f
C6282 PAD.n6774 VSS 0.036461f
C6283 PAD.n6776 VSS 0.036461f
C6284 PAD.n6777 VSS 0.036461f
C6285 PAD.n6778 VSS 0.036461f
C6286 PAD.n6780 VSS 0.036461f
C6287 PAD.n6781 VSS 0.036461f
C6288 PAD.n6782 VSS 0.036461f
C6289 PAD.n6784 VSS 0.036461f
C6290 PAD.n6785 VSS 0.036461f
C6291 PAD.n6786 VSS 0.036461f
C6292 PAD.n6788 VSS 0.036461f
C6293 PAD.n6789 VSS 0.036461f
C6294 PAD.n6790 VSS 0.036461f
C6295 PAD.n6792 VSS 0.036461f
C6296 PAD.n6793 VSS 0.036461f
C6297 PAD.n6794 VSS 0.036461f
C6298 PAD.n6796 VSS 0.036461f
C6299 PAD.n6797 VSS 0.036461f
C6300 PAD.n6798 VSS 0.036461f
C6301 PAD.n6800 VSS 0.036461f
C6302 PAD.n6801 VSS 0.036461f
C6303 PAD.n6802 VSS 0.036461f
C6304 PAD.n6803 VSS 0.023109f
C6305 PAD.n6804 VSS 0.023109f
C6306 PAD.n6806 VSS 0.036461f
C6307 PAD.n6808 VSS 0.036461f
C6308 PAD.n6810 VSS 0.036461f
C6309 PAD.n6811 VSS 0.036461f
C6310 PAD.n6812 VSS 0.036461f
C6311 PAD.n6813 VSS 0.036461f
C6312 PAD.n6814 VSS 0.036461f
C6313 PAD.n6815 VSS 0.036461f
C6314 PAD.n6816 VSS 0.036461f
C6315 PAD.n6818 VSS 0.036461f
C6316 PAD.n6820 VSS 0.036461f
C6317 PAD.n6822 VSS 0.036461f
C6318 PAD.n6823 VSS 0.036461f
C6319 PAD.n6824 VSS 0.036461f
C6320 PAD.n6825 VSS 0.036461f
C6321 PAD.n6826 VSS 0.036461f
C6322 PAD.n6827 VSS 0.036461f
C6323 PAD.n6828 VSS 0.036461f
C6324 PAD.n6830 VSS 0.036461f
C6325 PAD.n6832 VSS 0.036461f
C6326 PAD.n6834 VSS 0.036461f
C6327 PAD.n6835 VSS 0.036461f
C6328 PAD.n6836 VSS 0.036461f
C6329 PAD.n6837 VSS 0.036461f
C6330 PAD.n6838 VSS 0.036461f
C6331 PAD.n6839 VSS 0.036461f
C6332 PAD.n6840 VSS 0.036461f
C6333 PAD.n6842 VSS 0.036461f
C6334 PAD.n6844 VSS 0.036461f
C6335 PAD.n6846 VSS 0.036461f
C6336 PAD.n6847 VSS 0.036461f
C6337 PAD.n6848 VSS 0.036461f
C6338 PAD.n6849 VSS 0.036461f
C6339 PAD.n6850 VSS 0.036461f
C6340 PAD.n6851 VSS 0.036461f
C6341 PAD.n6852 VSS 0.036461f
C6342 PAD.n6854 VSS 0.036461f
C6343 PAD.n6856 VSS 0.036461f
C6344 PAD.n6858 VSS 0.036461f
C6345 PAD.n6859 VSS 0.036461f
C6346 PAD.n6860 VSS 0.036461f
C6347 PAD.n6861 VSS 0.036461f
C6348 PAD.n6862 VSS 0.036461f
C6349 PAD.n6863 VSS 0.036461f
C6350 PAD.n6864 VSS 0.036461f
C6351 PAD.n6866 VSS 0.036461f
C6352 PAD.n6868 VSS 0.036461f
C6353 PAD.n6870 VSS 0.036461f
C6354 PAD.n6871 VSS 0.036461f
C6355 PAD.n6872 VSS 0.036461f
C6356 PAD.n6873 VSS 0.036461f
C6357 PAD.n6874 VSS 0.036461f
C6358 PAD.n6875 VSS 0.036461f
C6359 PAD.n6876 VSS 0.036461f
C6360 PAD.n6878 VSS 0.036461f
C6361 PAD.n6880 VSS 0.036461f
C6362 PAD.n6882 VSS 0.036461f
C6363 PAD.n6883 VSS 0.036461f
C6364 PAD.n6884 VSS 0.036461f
C6365 PAD.n6885 VSS 0.036461f
C6366 PAD.n6886 VSS 0.036461f
C6367 PAD.n6887 VSS 0.036461f
C6368 PAD.n6888 VSS 0.036461f
C6369 PAD.n6890 VSS 0.036461f
C6370 PAD.n6892 VSS 0.036461f
C6371 PAD.n6894 VSS 0.036461f
C6372 PAD.n6895 VSS 0.036461f
C6373 PAD.n6896 VSS 0.036461f
C6374 PAD.n6897 VSS 0.036461f
C6375 PAD.n6898 VSS 0.036461f
C6376 PAD.n6899 VSS 0.036461f
C6377 PAD.n6900 VSS 0.036461f
C6378 PAD.n6902 VSS 0.036461f
C6379 PAD.n6904 VSS 0.036461f
C6380 PAD.n6906 VSS 0.036461f
C6381 PAD.n6907 VSS 0.036461f
C6382 PAD.n6908 VSS 0.036461f
C6383 PAD.n6909 VSS 0.036461f
C6384 PAD.n6910 VSS 0.036461f
C6385 PAD.n6911 VSS 0.036461f
C6386 PAD.n6912 VSS 0.036461f
C6387 PAD.n6914 VSS 0.036461f
C6388 PAD.n6916 VSS 0.036461f
C6389 PAD.n6918 VSS 0.036461f
C6390 PAD.n6919 VSS 0.036461f
C6391 PAD.n6920 VSS 0.036461f
C6392 PAD.n6921 VSS 0.036461f
C6393 PAD.n6922 VSS 0.036461f
C6394 PAD.n6923 VSS 0.036461f
C6395 PAD.n6924 VSS 0.036461f
C6396 PAD.n6926 VSS 0.036461f
C6397 PAD.n6928 VSS 0.036461f
C6398 PAD.n6930 VSS 0.036461f
C6399 PAD.n6931 VSS 0.036461f
C6400 PAD.n6932 VSS 0.036461f
C6401 PAD.n6933 VSS 0.036461f
C6402 PAD.n6934 VSS 0.036461f
C6403 PAD.n6935 VSS 0.036461f
C6404 PAD.n6936 VSS 0.036461f
C6405 PAD.n6938 VSS 0.036461f
C6406 PAD.n6940 VSS 0.036461f
C6407 PAD.n6942 VSS 0.036461f
C6408 PAD.n6943 VSS 0.036461f
C6409 PAD.n6944 VSS 0.036461f
C6410 PAD.n6945 VSS 0.036461f
C6411 PAD.n6946 VSS 0.036461f
C6412 PAD.n6947 VSS 0.036461f
C6413 PAD.n6948 VSS 0.036461f
C6414 PAD.n6950 VSS 0.036461f
C6415 PAD.n6952 VSS 0.036461f
C6416 PAD.n6954 VSS 0.036461f
C6417 PAD.n6955 VSS 0.036461f
C6418 PAD.n6956 VSS 0.036461f
C6419 PAD.n6957 VSS 0.036461f
C6420 PAD.n6958 VSS 0.036461f
C6421 PAD.n6959 VSS 0.036461f
C6422 PAD.n6960 VSS 0.036461f
C6423 PAD.n6962 VSS 0.036461f
C6424 PAD.n6964 VSS 0.036461f
C6425 PAD.n6966 VSS 0.036461f
C6426 PAD.n6967 VSS 0.036461f
C6427 PAD.n6968 VSS 0.036461f
C6428 PAD.n6969 VSS 0.036461f
C6429 PAD.n6970 VSS 0.036461f
C6430 PAD.n6971 VSS 0.036461f
C6431 PAD.n6972 VSS 0.036461f
C6432 PAD.n6974 VSS 0.036461f
C6433 PAD.n6976 VSS 0.036461f
C6434 PAD.n6978 VSS 0.036461f
C6435 PAD.n6979 VSS 0.036461f
C6436 PAD.n6980 VSS 0.036461f
C6437 PAD.n6981 VSS 0.036461f
C6438 PAD.n6982 VSS 0.036461f
C6439 PAD.n6983 VSS 0.036461f
C6440 PAD.n6984 VSS 0.036461f
C6441 PAD.n6986 VSS 0.036461f
C6442 PAD.n6988 VSS 0.036461f
C6443 PAD.n6990 VSS 0.036461f
C6444 PAD.n6991 VSS 0.036461f
C6445 PAD.n6992 VSS 0.036461f
C6446 PAD.n6993 VSS 0.036461f
C6447 PAD.n6994 VSS 0.036461f
C6448 PAD.n6995 VSS 0.036461f
C6449 PAD.n6996 VSS 0.036461f
C6450 PAD.n6998 VSS 0.036461f
C6451 PAD.n7000 VSS 0.036461f
C6452 PAD.n7002 VSS 0.036461f
C6453 PAD.n7003 VSS 0.036461f
C6454 PAD.n7004 VSS 0.036461f
C6455 PAD.n7005 VSS 0.036461f
C6456 PAD.n7006 VSS 0.036461f
C6457 PAD.n7007 VSS 0.036461f
C6458 PAD.n7008 VSS 0.036461f
C6459 PAD.n7010 VSS 0.036461f
C6460 PAD.n7012 VSS 0.036461f
C6461 PAD.n7014 VSS 0.036461f
C6462 PAD.n7015 VSS 0.036461f
C6463 PAD.n7016 VSS 0.036461f
C6464 PAD.n7017 VSS 0.036461f
C6465 PAD.n7018 VSS 0.036461f
C6466 PAD.n7019 VSS 0.036461f
C6467 PAD.n7020 VSS 0.036461f
C6468 PAD.n7022 VSS 0.036461f
C6469 PAD.n7024 VSS 0.036461f
C6470 PAD.n7026 VSS 0.036461f
C6471 PAD.n7027 VSS 0.036461f
C6472 PAD.n7028 VSS 0.036461f
C6473 PAD.n7029 VSS 0.036461f
C6474 PAD.n7030 VSS 0.036461f
C6475 PAD.n7031 VSS 0.036461f
C6476 PAD.n7032 VSS 0.036461f
C6477 PAD.n7034 VSS 0.036461f
C6478 PAD.n7036 VSS 0.036461f
C6479 PAD.n7038 VSS 0.036461f
C6480 PAD.n7039 VSS 0.036461f
C6481 PAD.n7040 VSS 0.036461f
C6482 PAD.n7041 VSS 0.036461f
C6483 PAD.n7042 VSS 0.036461f
C6484 PAD.n7043 VSS 0.036461f
C6485 PAD.n7044 VSS 0.036461f
C6486 PAD.n7046 VSS 0.036461f
C6487 PAD.n7048 VSS 0.036461f
C6488 PAD.n7049 VSS 0.036461f
C6489 PAD.n7050 VSS 0.023109f
C6490 PAD.n7051 VSS 0.03338f
C6491 PAD.n7052 VSS 0.054012f
C6492 PAD.n7053 VSS 0.054012f
C6493 PAD.n7054 VSS 0.048212f
C6494 PAD.n7055 VSS 0.046286f
C6495 PAD.n7056 VSS 0.046286f
C6496 PAD.n7057 VSS 0.039761f
C6497 PAD.n7058 VSS 0.039761f
C6498 PAD.n7059 VSS 0.522934f
C6499 PAD.n7060 VSS 0.700534f
C6500 PAD.n7061 VSS 0.611734f
C6501 PAD.n7103 VSS 0.453867f
C6502 PAD.n7104 VSS 0.036461f
C6503 PAD.n7105 VSS 0.606801f
C6504 PAD.n7106 VSS 0.036461f
C6505 PAD.n7107 VSS 0.036461f
C6506 PAD.n7108 VSS 0.036461f
C6507 PAD.n7109 VSS 0.036461f
C6508 PAD.n7110 VSS 0.036461f
C6509 PAD.n7111 VSS 0.036461f
C6510 PAD.n7112 VSS 0.036461f
C6511 PAD.n7113 VSS 0.036461f
C6512 PAD.n7114 VSS 0.036461f
C6513 PAD.n7115 VSS 0.036461f
C6514 PAD.n7116 VSS 0.036461f
C6515 PAD.n7117 VSS 0.036461f
C6516 PAD.n7118 VSS 0.036461f
C6517 PAD.n7119 VSS 0.036461f
C6518 PAD.n7120 VSS 0.036461f
C6519 PAD.n7121 VSS 0.036461f
C6520 PAD.n7122 VSS 0.036461f
C6521 PAD.n7123 VSS 0.036461f
C6522 PAD.n7124 VSS 0.036461f
C6523 PAD.n7125 VSS 0.036461f
C6524 PAD.n7126 VSS 0.036461f
C6525 PAD.n7127 VSS 0.036461f
C6526 PAD.n7128 VSS 0.036461f
C6527 PAD.n7129 VSS 0.036461f
C6528 PAD.n7130 VSS 0.036461f
C6529 PAD.n7131 VSS 0.036461f
C6530 PAD.n7132 VSS 0.036461f
C6531 PAD.n7133 VSS 0.036461f
C6532 PAD.n7134 VSS 0.036461f
C6533 PAD.n7135 VSS 0.036461f
C6534 PAD.n7136 VSS 0.036461f
C6535 PAD.n7137 VSS 0.036461f
C6536 PAD.n7138 VSS 0.036461f
C6537 PAD.n7139 VSS 0.036461f
C6538 PAD.n7140 VSS 0.036461f
C6539 PAD.n7141 VSS 0.036461f
C6540 PAD.n7142 VSS 0.036461f
C6541 PAD.n7143 VSS 0.036461f
C6542 PAD.n7144 VSS 0.036461f
C6543 PAD.n7145 VSS 0.036461f
C6544 PAD.n7146 VSS 0.036461f
C6545 PAD.n7147 VSS 0.030555f
C6546 PAD.n7148 VSS 0.029436f
C6547 PAD.n7149 VSS 0.0441f
C6548 PAD.n7150 VSS 0.049115f
C6549 PAD.n7151 VSS 0.049115f
C6550 PAD.n7152 VSS 0.0441f
C6551 PAD.n7153 VSS 0.038515f
C6552 PAD.n7154 VSS 0.033773f
C6553 PAD.n7155 VSS 0.033773f
C6554 PAD.n7156 VSS 0.029436f
C6555 PAD.n7157 VSS 0.029436f
C6556 PAD.n7158 VSS 0.700534f
C6557 PAD.n7200 VSS 0.596934f
C6558 PAD.n7201 VSS 0.036461f
C6559 PAD.n7202 VSS 0.074644f
C6560 PAD.n7203 VSS 0.029755f
C6561 PAD.n7204 VSS 0.034069f
C6562 PAD.n7205 VSS 0.034069f
C6563 PAD.n7206 VSS 0.374933f
C6564 PAD.n7207 VSS 0.3404f
C6565 PAD.n7208 VSS 0.074644f
C6566 PAD.n7209 VSS 0.036461f
C6567 PAD.n7210 VSS 0.062274f
C6568 PAD.n7211 VSS 0.069765f
C6569 PAD.n7212 VSS 0.038168f
C6570 PAD.n7213 VSS 0.042759f
C6571 PAD.n7214 VSS 0.042759f
C6572 PAD.n7215 VSS 0.611734f
C6573 PAD.n7216 VSS 0.453867f
C6574 PAD.n7217 VSS 0.069765f
C6575 PAD.n7218 VSS 0.069765f
C6576 PAD.n7219 VSS 0.069765f
C6577 PAD.n7220 VSS 0.062274f
C6578 PAD.n7221 VSS 0.675868f
C6579 PAD.n7222 VSS 0.611734f
C6580 PAD.n7223 VSS 0.596934f
C6581 PAD.n7224 VSS 0.069765f
C6582 PAD.n7225 VSS 0.069765f
C6583 PAD.n7226 VSS 0.062274f
C6584 PAD.n7227 VSS 0.077423f
C6585 PAD.n7228 VSS 0.036461f
C6586 PAD.n7229 VSS 0.036461f
C6587 PAD.n7230 VSS 0.036461f
C6588 PAD.n7231 VSS 0.036461f
C6589 PAD.n7232 VSS 0.036461f
C6590 PAD.n7233 VSS 0.036461f
C6591 PAD.n7234 VSS 0.036461f
C6592 PAD.n7235 VSS 0.036461f
C6593 PAD.n7236 VSS 0.036461f
C6594 PAD.n7237 VSS 0.036461f
C6595 PAD.n7238 VSS 0.036461f
C6596 PAD.n7239 VSS 0.036461f
C6597 PAD.n7240 VSS 0.036461f
C6598 PAD.n7241 VSS 0.036461f
C6599 PAD.n7242 VSS 0.036461f
C6600 PAD.n7243 VSS 0.036461f
C6601 PAD.n7244 VSS 0.036461f
C6602 PAD.n7245 VSS 0.036461f
C6603 PAD.n7246 VSS 0.036461f
C6604 PAD.n7247 VSS 0.036461f
C6605 PAD.n7248 VSS 0.036461f
C6606 PAD.n7249 VSS 0.036461f
C6607 PAD.n7250 VSS 0.036461f
C6608 PAD.n7251 VSS 0.036461f
C6609 PAD.n7252 VSS 0.036461f
C6610 PAD.n7253 VSS 0.036461f
C6611 PAD.n7254 VSS 0.036461f
C6612 PAD.n7255 VSS 0.036461f
C6613 PAD.n7256 VSS 0.036461f
C6614 PAD.n7257 VSS 0.036461f
C6615 PAD.n7258 VSS 0.036461f
C6616 PAD.n7259 VSS 0.036461f
C6617 PAD.n7260 VSS 0.036461f
C6618 PAD.n7261 VSS 0.036461f
C6619 PAD.n7262 VSS 0.036461f
C6620 PAD.n7263 VSS 0.036461f
C6621 PAD.n7264 VSS 0.036461f
C6622 PAD.n7265 VSS 0.036461f
C6623 PAD.n7266 VSS 0.036461f
C6624 PAD.n7267 VSS 0.036461f
C6625 PAD.n7268 VSS 0.030555f
C6626 PAD.n7269 VSS 0.023109f
C6627 PAD.n7270 VSS 0.023109f
C6628 PAD.n7271 VSS 0.036461f
C6629 PAD.n7273 VSS 0.036461f
C6630 PAD.n7274 VSS 0.036461f
C6631 PAD.n7275 VSS 0.036461f
C6632 PAD.n7276 VSS 0.036461f
C6633 PAD.n7277 VSS 0.036461f
C6634 PAD.n7278 VSS 0.036461f
C6635 PAD.n7279 VSS 0.036461f
C6636 PAD.n7281 VSS 0.036461f
C6637 PAD.n7282 VSS 0.036461f
C6638 PAD.n7283 VSS 0.036461f
C6639 PAD.n7285 VSS 0.036461f
C6640 PAD.n7286 VSS 0.036461f
C6641 PAD.n7287 VSS 0.036461f
C6642 PAD.n7288 VSS 0.036461f
C6643 PAD.n7289 VSS 0.036461f
C6644 PAD.n7290 VSS 0.036461f
C6645 PAD.n7291 VSS 0.036461f
C6646 PAD.n7293 VSS 0.036461f
C6647 PAD.n7294 VSS 0.036461f
C6648 PAD.n7295 VSS 0.036461f
C6649 PAD.n7297 VSS 0.036461f
C6650 PAD.n7298 VSS 0.036461f
C6651 PAD.n7299 VSS 0.036461f
C6652 PAD.n7300 VSS 0.036461f
C6653 PAD.n7301 VSS 0.036461f
C6654 PAD.n7302 VSS 0.036461f
C6655 PAD.n7303 VSS 0.036461f
C6656 PAD.n7305 VSS 0.036461f
C6657 PAD.n7306 VSS 0.036461f
C6658 PAD.n7307 VSS 0.036461f
C6659 PAD.n7309 VSS 0.036461f
C6660 PAD.n7310 VSS 0.036461f
C6661 PAD.n7311 VSS 0.036461f
C6662 PAD.n7312 VSS 0.036461f
C6663 PAD.n7313 VSS 0.036461f
C6664 PAD.n7314 VSS 0.036461f
C6665 PAD.n7315 VSS 0.036461f
C6666 PAD.n7317 VSS 0.036461f
C6667 PAD.n7318 VSS 0.036461f
C6668 PAD.n7319 VSS 0.036461f
C6669 PAD.n7321 VSS 0.036461f
C6670 PAD.n7322 VSS 0.036461f
C6671 PAD.n7323 VSS 0.036461f
C6672 PAD.n7324 VSS 0.036461f
C6673 PAD.n7325 VSS 0.036461f
C6674 PAD.n7326 VSS 0.036461f
C6675 PAD.n7327 VSS 0.036461f
C6676 PAD.n7329 VSS 0.036461f
C6677 PAD.n7330 VSS 0.036461f
C6678 PAD.n7331 VSS 0.036461f
C6679 PAD.n7333 VSS 0.036461f
C6680 PAD.n7334 VSS 0.036461f
C6681 PAD.n7335 VSS 0.036461f
C6682 PAD.n7336 VSS 0.036461f
C6683 PAD.n7337 VSS 0.036461f
C6684 PAD.n7338 VSS 0.036461f
C6685 PAD.n7339 VSS 0.036461f
C6686 PAD.n7341 VSS 0.036461f
C6687 PAD.n7342 VSS 0.036461f
C6688 PAD.n7343 VSS 0.036461f
C6689 PAD.n7345 VSS 0.036461f
C6690 PAD.n7346 VSS 0.036461f
C6691 PAD.n7347 VSS 0.036461f
C6692 PAD.n7348 VSS 0.036461f
C6693 PAD.n7349 VSS 0.036461f
C6694 PAD.n7350 VSS 0.036461f
C6695 PAD.n7351 VSS 0.036461f
C6696 PAD.n7353 VSS 0.036461f
C6697 PAD.n7354 VSS 0.036461f
C6698 PAD.n7355 VSS 0.036461f
C6699 PAD.n7357 VSS 0.036461f
C6700 PAD.n7358 VSS 0.036461f
C6701 PAD.n7359 VSS 0.036461f
C6702 PAD.n7360 VSS 0.036461f
C6703 PAD.n7361 VSS 0.036461f
C6704 PAD.n7362 VSS 0.036461f
C6705 PAD.n7363 VSS 0.036461f
C6706 PAD.n7365 VSS 0.036461f
C6707 PAD.n7366 VSS 0.036461f
C6708 PAD.n7367 VSS 0.036461f
C6709 PAD.n7369 VSS 0.036461f
C6710 PAD.n7370 VSS 0.036461f
C6711 PAD.n7371 VSS 0.036461f
C6712 PAD.n7372 VSS 0.036461f
C6713 PAD.n7373 VSS 0.036461f
C6714 PAD.n7374 VSS 0.036461f
C6715 PAD.n7375 VSS 0.036461f
C6716 PAD.n7377 VSS 0.036461f
C6717 PAD.n7378 VSS 0.036461f
C6718 PAD.n7379 VSS 0.036461f
C6719 PAD.n7381 VSS 0.036461f
C6720 PAD.n7382 VSS 0.036461f
C6721 PAD.n7383 VSS 0.036461f
C6722 PAD.n7384 VSS 0.036461f
C6723 PAD.n7385 VSS 0.036461f
C6724 PAD.n7386 VSS 0.036461f
C6725 PAD.n7387 VSS 0.036461f
C6726 PAD.n7389 VSS 0.036461f
C6727 PAD.n7390 VSS 0.036461f
C6728 PAD.n7391 VSS 0.036461f
C6729 PAD.n7393 VSS 0.036461f
C6730 PAD.n7394 VSS 0.036461f
C6731 PAD.n7395 VSS 0.036461f
C6732 PAD.n7396 VSS 0.036461f
C6733 PAD.n7397 VSS 0.036461f
C6734 PAD.n7398 VSS 0.036461f
C6735 PAD.n7399 VSS 0.036461f
C6736 PAD.n7401 VSS 0.036461f
C6737 PAD.n7402 VSS 0.036461f
C6738 PAD.n7403 VSS 0.036461f
C6739 PAD.n7405 VSS 0.036461f
C6740 PAD.n7406 VSS 0.036461f
C6741 PAD.n7407 VSS 0.036461f
C6742 PAD.n7408 VSS 0.036461f
C6743 PAD.n7409 VSS 0.036461f
C6744 PAD.n7410 VSS 0.036461f
C6745 PAD.n7411 VSS 0.036461f
C6746 PAD.n7413 VSS 0.036461f
C6747 PAD.n7414 VSS 0.036461f
C6748 PAD.n7415 VSS 0.036461f
C6749 PAD.n7417 VSS 0.036461f
C6750 PAD.n7418 VSS 0.036461f
C6751 PAD.n7419 VSS 0.036461f
C6752 PAD.n7420 VSS 0.036461f
C6753 PAD.n7421 VSS 0.036461f
C6754 PAD.n7422 VSS 0.036461f
C6755 PAD.n7423 VSS 0.036461f
C6756 PAD.n7425 VSS 0.036461f
C6757 PAD.n7426 VSS 0.036461f
C6758 PAD.n7427 VSS 0.036461f
C6759 PAD.n7429 VSS 0.036461f
C6760 PAD.n7430 VSS 0.036461f
C6761 PAD.n7431 VSS 0.036461f
C6762 PAD.n7432 VSS 0.036461f
C6763 PAD.n7433 VSS 0.036461f
C6764 PAD.n7434 VSS 0.036461f
C6765 PAD.n7435 VSS 0.036461f
C6766 PAD.n7437 VSS 0.036461f
C6767 PAD.n7438 VSS 0.036461f
C6768 PAD.n7439 VSS 0.036461f
C6769 PAD.n7441 VSS 0.036461f
C6770 PAD.n7442 VSS 0.036461f
C6771 PAD.n7443 VSS 0.036461f
C6772 PAD.n7444 VSS 0.036461f
C6773 PAD.n7445 VSS 0.036461f
C6774 PAD.n7446 VSS 0.036461f
C6775 PAD.n7447 VSS 0.036461f
C6776 PAD.n7449 VSS 0.036461f
C6777 PAD.n7450 VSS 0.036461f
C6778 PAD.n7451 VSS 0.036461f
C6779 PAD.n7453 VSS 0.036461f
C6780 PAD.n7454 VSS 0.036461f
C6781 PAD.n7455 VSS 0.036461f
C6782 PAD.n7456 VSS 0.036461f
C6783 PAD.n7457 VSS 0.036461f
C6784 PAD.n7458 VSS 0.036461f
C6785 PAD.n7459 VSS 0.036461f
C6786 PAD.n7461 VSS 0.036461f
C6787 PAD.n7462 VSS 0.036461f
C6788 PAD.n7463 VSS 0.036461f
C6789 PAD.n7465 VSS 0.036461f
C6790 PAD.n7466 VSS 0.036461f
C6791 PAD.n7467 VSS 0.036461f
C6792 PAD.n7468 VSS 0.036461f
C6793 PAD.n7469 VSS 0.036461f
C6794 PAD.n7470 VSS 0.036461f
C6795 PAD.n7471 VSS 0.036461f
C6796 PAD.n7473 VSS 0.036461f
C6797 PAD.n7474 VSS 0.036461f
C6798 PAD.n7475 VSS 0.036461f
C6799 PAD.n7477 VSS 0.036461f
C6800 PAD.n7478 VSS 0.036461f
C6801 PAD.n7479 VSS 0.036461f
C6802 PAD.n7480 VSS 0.036461f
C6803 PAD.n7481 VSS 0.036461f
C6804 PAD.n7482 VSS 0.036461f
C6805 PAD.n7483 VSS 0.036461f
C6806 PAD.n7485 VSS 0.036461f
C6807 PAD.n7486 VSS 0.036461f
C6808 PAD.n7487 VSS 0.036461f
C6809 PAD.n7489 VSS 0.036461f
C6810 PAD.n7490 VSS 0.036461f
C6811 PAD.n7491 VSS 0.036461f
C6812 PAD.n7492 VSS 0.036461f
C6813 PAD.n7493 VSS 0.036461f
C6814 PAD.n7494 VSS 0.036461f
C6815 PAD.n7495 VSS 0.036461f
C6816 PAD.n7497 VSS 0.036461f
C6817 PAD.n7498 VSS 0.036461f
C6818 PAD.n7499 VSS 0.036461f
C6819 PAD.n7501 VSS 0.036461f
C6820 PAD.n7502 VSS 0.036461f
C6821 PAD.n7503 VSS 0.036461f
C6822 PAD.n7504 VSS 0.036461f
C6823 PAD.n7505 VSS 0.036461f
C6824 PAD.n7506 VSS 0.036461f
C6825 PAD.n7507 VSS 0.036461f
C6826 PAD.n7509 VSS 0.036461f
C6827 PAD.n7510 VSS 0.036461f
C6828 PAD.n7512 VSS 0.036461f
C6829 PAD.n7513 VSS 0.036461f
C6830 PAD.n7514 VSS 0.036461f
C6831 PAD.n7515 VSS 0.036461f
C6832 PAD.n7516 VSS 0.03338f
C6833 PAD.n7517 VSS 0.023109f
C6834 PAD.n7518 VSS 0.023109f
C6835 PAD.n7520 VSS 0.429201f
C6836 PAD.n7521 VSS 0.286133f
C6837 PAD.n7522 VSS 0.039603f
C6838 PAD.n7523 VSS 0.039603f
C6839 PAD.n7524 VSS 0.034588f
C6840 PAD.n7525 VSS 0.042895f
C6841 PAD.n7526 VSS 0.025828f
C6842 PAD.n7527 VSS 0.029573f
C6843 PAD.n7528 VSS 0.2516f
C6844 PAD.n7529 VSS 0.029573f
C6845 PAD.n7530 VSS 0.029436f
C6846 PAD.n7531 VSS 0.023109f
C6847 PAD.n7532 VSS 0.023109f
C6848 PAD.n7533 VSS 0.036461f
C6849 PAD.n7535 VSS 0.036461f
C6850 PAD.n7536 VSS 0.036461f
C6851 PAD.n7537 VSS 0.036461f
C6852 PAD.n7538 VSS 0.036461f
C6853 PAD.n7539 VSS 0.036461f
C6854 PAD.n7540 VSS 0.036461f
C6855 PAD.n7541 VSS 0.036461f
C6856 PAD.n7543 VSS 0.036461f
C6857 PAD.n7544 VSS 0.036461f
C6858 PAD.n7545 VSS 0.036461f
C6859 PAD.n7547 VSS 0.036461f
C6860 PAD.n7548 VSS 0.036461f
C6861 PAD.n7549 VSS 0.036461f
C6862 PAD.n7550 VSS 0.036461f
C6863 PAD.n7551 VSS 0.036461f
C6864 PAD.n7552 VSS 0.036461f
C6865 PAD.n7553 VSS 0.036461f
C6866 PAD.n7555 VSS 0.036461f
C6867 PAD.n7556 VSS 0.036461f
C6868 PAD.n7557 VSS 0.036461f
C6869 PAD.n7559 VSS 0.036461f
C6870 PAD.n7560 VSS 0.036461f
C6871 PAD.n7561 VSS 0.036461f
C6872 PAD.n7562 VSS 0.036461f
C6873 PAD.n7563 VSS 0.036461f
C6874 PAD.n7564 VSS 0.036461f
C6875 PAD.n7565 VSS 0.036461f
C6876 PAD.n7567 VSS 0.036461f
C6877 PAD.n7568 VSS 0.036461f
C6878 PAD.n7569 VSS 0.036461f
C6879 PAD.n7571 VSS 0.036461f
C6880 PAD.n7572 VSS 0.036461f
C6881 PAD.n7573 VSS 0.036461f
C6882 PAD.n7574 VSS 0.036461f
C6883 PAD.n7575 VSS 0.036461f
C6884 PAD.n7576 VSS 0.036461f
C6885 PAD.n7577 VSS 0.036461f
C6886 PAD.n7579 VSS 0.036461f
C6887 PAD.n7580 VSS 0.036461f
C6888 PAD.n7581 VSS 0.036461f
C6889 PAD.n7583 VSS 0.036461f
C6890 PAD.n7584 VSS 0.036461f
C6891 PAD.n7585 VSS 0.036461f
C6892 PAD.n7586 VSS 0.036461f
C6893 PAD.n7587 VSS 0.036461f
C6894 PAD.n7588 VSS 0.036461f
C6895 PAD.n7589 VSS 0.036461f
C6896 PAD.n7591 VSS 0.036461f
C6897 PAD.n7592 VSS 0.036461f
C6898 PAD.n7593 VSS 0.036461f
C6899 PAD.n7595 VSS 0.036461f
C6900 PAD.n7596 VSS 0.036461f
C6901 PAD.n7597 VSS 0.036461f
C6902 PAD.n7598 VSS 0.036461f
C6903 PAD.n7599 VSS 0.036461f
C6904 PAD.n7600 VSS 0.036461f
C6905 PAD.n7601 VSS 0.036461f
C6906 PAD.n7603 VSS 0.036461f
C6907 PAD.n7604 VSS 0.036461f
C6908 PAD.n7605 VSS 0.036461f
C6909 PAD.n7607 VSS 0.036461f
C6910 PAD.n7608 VSS 0.036461f
C6911 PAD.n7609 VSS 0.036461f
C6912 PAD.n7610 VSS 0.036461f
C6913 PAD.n7611 VSS 0.036461f
C6914 PAD.n7612 VSS 0.036461f
C6915 PAD.n7613 VSS 0.036461f
C6916 PAD.n7615 VSS 0.036461f
C6917 PAD.n7616 VSS 0.036461f
C6918 PAD.n7617 VSS 0.036461f
C6919 PAD.n7619 VSS 0.036461f
C6920 PAD.n7620 VSS 0.036461f
C6921 PAD.n7621 VSS 0.036461f
C6922 PAD.n7622 VSS 0.036461f
C6923 PAD.n7623 VSS 0.036461f
C6924 PAD.n7624 VSS 0.036461f
C6925 PAD.n7625 VSS 0.036461f
C6926 PAD.n7627 VSS 0.036461f
C6927 PAD.n7628 VSS 0.036461f
C6928 PAD.n7629 VSS 0.036461f
C6929 PAD.n7631 VSS 0.036461f
C6930 PAD.n7632 VSS 0.036461f
C6931 PAD.n7633 VSS 0.036461f
C6932 PAD.n7634 VSS 0.036461f
C6933 PAD.n7635 VSS 0.036461f
C6934 PAD.n7636 VSS 0.036461f
C6935 PAD.n7637 VSS 0.036461f
C6936 PAD.n7639 VSS 0.036461f
C6937 PAD.n7640 VSS 0.036461f
C6938 PAD.n7641 VSS 0.036461f
C6939 PAD.n7643 VSS 0.036461f
C6940 PAD.n7644 VSS 0.036461f
C6941 PAD.n7645 VSS 0.036461f
C6942 PAD.n7646 VSS 0.036461f
C6943 PAD.n7647 VSS 0.036461f
C6944 PAD.n7648 VSS 0.036461f
C6945 PAD.n7649 VSS 0.036461f
C6946 PAD.n7651 VSS 0.036461f
C6947 PAD.n7652 VSS 0.036461f
C6948 PAD.n7653 VSS 0.036461f
C6949 PAD.n7655 VSS 0.036461f
C6950 PAD.n7656 VSS 0.036461f
C6951 PAD.n7657 VSS 0.036461f
C6952 PAD.n7658 VSS 0.036461f
C6953 PAD.n7659 VSS 0.036461f
C6954 PAD.n7660 VSS 0.036461f
C6955 PAD.n7661 VSS 0.036461f
C6956 PAD.n7663 VSS 0.036461f
C6957 PAD.n7664 VSS 0.036461f
C6958 PAD.n7665 VSS 0.036461f
C6959 PAD.n7667 VSS 0.036461f
C6960 PAD.n7668 VSS 0.036461f
C6961 PAD.n7669 VSS 0.036461f
C6962 PAD.n7670 VSS 0.036461f
C6963 PAD.n7671 VSS 0.036461f
C6964 PAD.n7672 VSS 0.036461f
C6965 PAD.n7673 VSS 0.036461f
C6966 PAD.n7675 VSS 0.036461f
C6967 PAD.n7676 VSS 0.036461f
C6968 PAD.n7677 VSS 0.036461f
C6969 PAD.n7679 VSS 0.036461f
C6970 PAD.n7680 VSS 0.036461f
C6971 PAD.n7681 VSS 0.036461f
C6972 PAD.n7682 VSS 0.036461f
C6973 PAD.n7683 VSS 0.036461f
C6974 PAD.n7684 VSS 0.036461f
C6975 PAD.n7685 VSS 0.036461f
C6976 PAD.n7687 VSS 0.036461f
C6977 PAD.n7688 VSS 0.036461f
C6978 PAD.n7689 VSS 0.036461f
C6979 PAD.n7691 VSS 0.036461f
C6980 PAD.n7692 VSS 0.036461f
C6981 PAD.n7693 VSS 0.036461f
C6982 PAD.n7694 VSS 0.036461f
C6983 PAD.n7695 VSS 0.036461f
C6984 PAD.n7696 VSS 0.036461f
C6985 PAD.n7697 VSS 0.036461f
C6986 PAD.n7699 VSS 0.036461f
C6987 PAD.n7700 VSS 0.036461f
C6988 PAD.n7701 VSS 0.036461f
C6989 PAD.n7703 VSS 0.036461f
C6990 PAD.n7704 VSS 0.036461f
C6991 PAD.n7705 VSS 0.036461f
C6992 PAD.n7706 VSS 0.036461f
C6993 PAD.n7707 VSS 0.036461f
C6994 PAD.n7708 VSS 0.036461f
C6995 PAD.n7709 VSS 0.036461f
C6996 PAD.n7711 VSS 0.036461f
C6997 PAD.n7712 VSS 0.036461f
C6998 PAD.n7713 VSS 0.036461f
C6999 PAD.n7715 VSS 0.036461f
C7000 PAD.n7716 VSS 0.036461f
C7001 PAD.n7717 VSS 0.036461f
C7002 PAD.n7718 VSS 0.036461f
C7003 PAD.n7719 VSS 0.036461f
C7004 PAD.n7720 VSS 0.036461f
C7005 PAD.n7721 VSS 0.036461f
C7006 PAD.n7723 VSS 0.036461f
C7007 PAD.n7724 VSS 0.036461f
C7008 PAD.n7725 VSS 0.036461f
C7009 PAD.n7727 VSS 0.036461f
C7010 PAD.n7728 VSS 0.036461f
C7011 PAD.n7729 VSS 0.036461f
C7012 PAD.n7730 VSS 0.036461f
C7013 PAD.n7731 VSS 0.036461f
C7014 PAD.n7732 VSS 0.036461f
C7015 PAD.n7733 VSS 0.036461f
C7016 PAD.n7735 VSS 0.036461f
C7017 PAD.n7736 VSS 0.036461f
C7018 PAD.n7737 VSS 0.036461f
C7019 PAD.n7739 VSS 0.036461f
C7020 PAD.n7740 VSS 0.036461f
C7021 PAD.n7741 VSS 0.036461f
C7022 PAD.n7742 VSS 0.036461f
C7023 PAD.n7743 VSS 0.036461f
C7024 PAD.n7744 VSS 0.036461f
C7025 PAD.n7745 VSS 0.036461f
C7026 PAD.n7747 VSS 0.036461f
C7027 PAD.n7748 VSS 0.036461f
C7028 PAD.n7749 VSS 0.036461f
C7029 PAD.n7751 VSS 0.036461f
C7030 PAD.n7752 VSS 0.036461f
C7031 PAD.n7753 VSS 0.036461f
C7032 PAD.n7754 VSS 0.036461f
C7033 PAD.n7755 VSS 0.036461f
C7034 PAD.n7756 VSS 0.036461f
C7035 PAD.n7757 VSS 0.036461f
C7036 PAD.n7759 VSS 0.036461f
C7037 PAD.n7760 VSS 0.036461f
C7038 PAD.n7761 VSS 0.036461f
C7039 PAD.n7763 VSS 0.036461f
C7040 PAD.n7764 VSS 0.036461f
C7041 PAD.n7765 VSS 0.036461f
C7042 PAD.n7766 VSS 0.036461f
C7043 PAD.n7767 VSS 0.036461f
C7044 PAD.n7768 VSS 0.036461f
C7045 PAD.n7769 VSS 0.036461f
C7046 PAD.n7771 VSS 0.036461f
C7047 PAD.n7772 VSS 0.036461f
C7048 PAD.n7774 VSS 0.036461f
C7049 PAD.n7775 VSS 0.036461f
C7050 PAD.n7776 VSS 0.036461f
C7051 PAD.n7777 VSS 0.036461f
C7052 PAD.n7778 VSS 0.03338f
C7053 PAD.n7779 VSS 0.023109f
C7054 PAD.n7780 VSS 0.023109f
C7055 PAD.n7782 VSS 0.611734f
C7056 PAD.n7783 VSS 0.246666f
C7057 PAD.n7784 VSS 0.061889f
C7058 PAD.n7785 VSS 0.061889f
C7059 PAD.n7786 VSS 0.055243f
C7060 PAD.n7787 VSS 0.062274f
C7061 PAD.n7788 VSS 0.045199f
C7062 PAD.n7789 VSS 0.050636f
C7063 PAD.n7790 VSS 0.050636f
C7064 PAD.n7791 VSS 0.350267f
C7065 PAD.n7792 VSS 0.611734f
C7066 PAD.n7793 VSS 0.025076f
C7067 PAD.n7794 VSS 0.025076f
C7068 PAD.n7795 VSS 0.021901f
C7069 PAD.n7796 VSS 0.033773f
C7070 PAD.n7797 VSS 0.042442f
C7071 PAD.n7798 VSS 0.039421f
C7072 PAD.n7799 VSS 0.045138f
C7073 PAD.n7800 VSS 0.045138f
C7074 PAD.n7801 VSS 0.611734f
C7075 PAD.n7802 VSS 0.222f
C7076 PAD.n7803 VSS 0.058513f
C7077 PAD.n7804 VSS 0.058513f
C7078 PAD.n7805 VSS 0.05223f
C7079 PAD.n7806 VSS 0.041766f
C7080 PAD.n7807 VSS 1.26464f
C7081 PAD.n7808 VSS 16.0867f
C7082 PAD.n7809 VSS 19.374f
C7083 PAD.n7810 VSS 13.1453f
C7084 PAD.n7811 VSS 14.5427f
C7085 PAD.n7812 VSS 8.779059f
C7086 PAD.n7813 VSS 0.061889f
C7087 PAD.n7814 VSS 0.034652f
C7088 PAD.n7815 VSS 0.046286f
C7089 PAD.n7816 VSS 0.038168f
C7090 PAD.n7817 VSS 0.042759f
C7091 PAD.n7818 VSS 0.042759f
C7092 PAD.n7819 VSS 0.675868f
C7093 PAD.n7820 VSS 0.187466f
C7094 PAD.n7821 VSS 0.035107f
C7095 PAD.n7822 VSS 0.035107f
C7096 PAD.n7823 VSS 0.030661f
C7097 PAD.n7824 VSS 0.033773f
C7098 PAD.n7825 VSS 0.033682f
C7099 PAD.n7826 VSS 0.038566f
C7100 PAD.n7827 VSS 0.038566f
C7101 PAD.n7828 VSS 0.098666f
C7102 PAD.n7829 VSS 0.685734f
C7103 PAD.n7871 VSS 0.036461f
C7104 PAD.n7873 VSS 0.036461f
C7105 PAD.n7874 VSS 0.036461f
C7106 PAD.n7875 VSS 0.036461f
C7107 PAD.n7876 VSS 0.036461f
C7108 PAD.n7877 VSS 0.036461f
C7109 PAD.n7879 VSS 0.036461f
C7110 PAD.n7880 VSS 0.036461f
C7111 PAD.n7881 VSS 0.036461f
C7112 PAD.n7882 VSS 0.036461f
C7113 PAD.n7884 VSS 0.036461f
C7114 PAD.n7885 VSS 0.036461f
C7115 PAD.n7886 VSS 0.036461f
C7116 PAD.n7887 VSS 0.036461f
C7117 PAD.n7889 VSS 0.036461f
C7118 PAD.n7890 VSS 0.036461f
C7119 PAD.n7891 VSS 0.036461f
C7120 PAD.n7892 VSS 0.036461f
C7121 PAD.n7894 VSS 0.036461f
C7122 PAD.n7895 VSS 0.036461f
C7123 PAD.n7896 VSS 0.036461f
C7124 PAD.n7897 VSS 0.036461f
C7125 PAD.n7899 VSS 0.036461f
C7126 PAD.n7900 VSS 0.036461f
C7127 PAD.n7901 VSS 0.036461f
C7128 PAD.n7902 VSS 0.036461f
C7129 PAD.n7904 VSS 0.036461f
C7130 PAD.n7905 VSS 0.036461f
C7131 PAD.n7906 VSS 0.036461f
C7132 PAD.n7907 VSS 0.036461f
C7133 PAD.n7909 VSS 0.036461f
C7134 PAD.n7910 VSS 0.036461f
C7135 PAD.n7911 VSS 0.036461f
C7136 PAD.n7912 VSS 0.036461f
C7137 PAD.n7914 VSS 0.036461f
C7138 PAD.n7915 VSS 0.036461f
C7139 PAD.n7916 VSS 0.036461f
C7140 PAD.n7917 VSS 0.036461f
C7141 PAD.n7919 VSS 0.036461f
C7142 PAD.n7920 VSS 0.036461f
C7143 PAD.n7921 VSS 0.036461f
C7144 PAD.n7922 VSS 0.036461f
C7145 PAD.n7924 VSS 0.036461f
C7146 PAD.n7925 VSS 0.036461f
C7147 PAD.n7926 VSS 0.036461f
C7148 PAD.n7927 VSS 0.036461f
C7149 PAD.n7929 VSS 0.036461f
C7150 PAD.n7930 VSS 0.036461f
C7151 PAD.n7931 VSS 0.036461f
C7152 PAD.n7932 VSS 0.036461f
C7153 PAD.n7934 VSS 0.036461f
C7154 PAD.n7935 VSS 0.036461f
C7155 PAD.n7936 VSS 0.036461f
C7156 PAD.n7937 VSS 0.036461f
C7157 PAD.n7939 VSS 0.036461f
C7158 PAD.n7940 VSS 0.036461f
C7159 PAD.n7941 VSS 0.036461f
C7160 PAD.n7942 VSS 0.036461f
C7161 PAD.n7944 VSS 0.036461f
C7162 PAD.n7945 VSS 0.036461f
C7163 PAD.n7946 VSS 0.036461f
C7164 PAD.n7947 VSS 0.036461f
C7165 PAD.n7949 VSS 0.036461f
C7166 PAD.n7950 VSS 0.036461f
C7167 PAD.n7951 VSS 0.036461f
C7168 PAD.n7952 VSS 0.036461f
C7169 PAD.n7954 VSS 0.036461f
C7170 PAD.n7955 VSS 0.036461f
C7171 PAD.n7956 VSS 0.036461f
C7172 PAD.n7957 VSS 0.036461f
C7173 PAD.n7959 VSS 0.036461f
C7174 PAD.n7960 VSS 0.036461f
C7175 PAD.n7961 VSS 0.036461f
C7176 PAD.n7962 VSS 0.036461f
C7177 PAD.n7964 VSS 0.036461f
C7178 PAD.n7965 VSS 0.036461f
C7179 PAD.n7966 VSS 0.036461f
C7180 PAD.n7967 VSS 0.036461f
C7181 PAD.n7969 VSS 0.036461f
C7182 PAD.n7970 VSS 0.036461f
C7183 PAD.n7971 VSS 0.023109f
C7184 PAD.n7972 VSS 0.023109f
C7185 PAD.n7973 VSS 0.036461f
C7186 PAD.n7974 VSS 0.036461f
C7187 PAD.n7976 VSS 0.036461f
C7188 PAD.n7977 VSS 0.036461f
C7189 PAD.n7978 VSS 0.036461f
C7190 PAD.n7979 VSS 0.036461f
C7191 PAD.n7980 VSS 0.036461f
C7192 PAD.n7981 VSS 0.036461f
C7193 PAD.n7983 VSS 0.036461f
C7194 PAD.n7984 VSS 0.036461f
C7195 PAD.n7985 VSS 0.036461f
C7196 PAD.n7986 VSS 0.036461f
C7197 PAD.n7987 VSS 0.036461f
C7198 PAD.n7988 VSS 0.036461f
C7199 PAD.n7989 VSS 0.036461f
C7200 PAD.n7990 VSS 0.036461f
C7201 PAD.n7992 VSS 0.036461f
C7202 PAD.n7993 VSS 0.036461f
C7203 PAD.n7994 VSS 0.036461f
C7204 PAD.n7995 VSS 0.036461f
C7205 PAD.n7996 VSS 0.036461f
C7206 PAD.n7997 VSS 0.036461f
C7207 PAD.n7998 VSS 0.036461f
C7208 PAD.n7999 VSS 0.036461f
C7209 PAD.n8001 VSS 0.036461f
C7210 PAD.n8002 VSS 0.036461f
C7211 PAD.n8003 VSS 0.036461f
C7212 PAD.n8004 VSS 0.036461f
C7213 PAD.n8005 VSS 0.036461f
C7214 PAD.n8006 VSS 0.036461f
C7215 PAD.n8007 VSS 0.036461f
C7216 PAD.n8008 VSS 0.036461f
C7217 PAD.n8010 VSS 0.036461f
C7218 PAD.n8011 VSS 0.036461f
C7219 PAD.n8012 VSS 0.036461f
C7220 PAD.n8013 VSS 0.036461f
C7221 PAD.n8014 VSS 0.036461f
C7222 PAD.n8015 VSS 0.036461f
C7223 PAD.n8016 VSS 0.036461f
C7224 PAD.n8017 VSS 0.036461f
C7225 PAD.n8019 VSS 0.036461f
C7226 PAD.n8020 VSS 0.036461f
C7227 PAD.n8021 VSS 0.036461f
C7228 PAD.n8022 VSS 0.036461f
C7229 PAD.n8023 VSS 0.036461f
C7230 PAD.n8024 VSS 0.036461f
C7231 PAD.n8025 VSS 0.036461f
C7232 PAD.n8026 VSS 0.036461f
C7233 PAD.n8028 VSS 0.036461f
C7234 PAD.n8029 VSS 0.036461f
C7235 PAD.n8030 VSS 0.036461f
C7236 PAD.n8031 VSS 0.036461f
C7237 PAD.n8032 VSS 0.036461f
C7238 PAD.n8033 VSS 0.036461f
C7239 PAD.n8034 VSS 0.036461f
C7240 PAD.n8035 VSS 0.036461f
C7241 PAD.n8037 VSS 0.036461f
C7242 PAD.n8038 VSS 0.036461f
C7243 PAD.n8039 VSS 0.036461f
C7244 PAD.n8040 VSS 0.036461f
C7245 PAD.n8041 VSS 0.036461f
C7246 PAD.n8042 VSS 0.036461f
C7247 PAD.n8043 VSS 0.036461f
C7248 PAD.n8044 VSS 0.036461f
C7249 PAD.n8046 VSS 0.036461f
C7250 PAD.n8047 VSS 0.036461f
C7251 PAD.n8048 VSS 0.036461f
C7252 PAD.n8049 VSS 0.036461f
C7253 PAD.n8050 VSS 0.036461f
C7254 PAD.n8051 VSS 0.036461f
C7255 PAD.n8052 VSS 0.036461f
C7256 PAD.n8053 VSS 0.036461f
C7257 PAD.n8055 VSS 0.036461f
C7258 PAD.n8056 VSS 0.036461f
C7259 PAD.n8057 VSS 0.036461f
C7260 PAD.n8058 VSS 0.036461f
C7261 PAD.n8059 VSS 0.036461f
C7262 PAD.n8060 VSS 0.036461f
C7263 PAD.n8061 VSS 0.036461f
C7264 PAD.n8062 VSS 0.036461f
C7265 PAD.n8064 VSS 0.036461f
C7266 PAD.n8065 VSS 0.036461f
C7267 PAD.n8066 VSS 0.036461f
C7268 PAD.n8067 VSS 0.036461f
C7269 PAD.n8068 VSS 0.036461f
C7270 PAD.n8069 VSS 0.036461f
C7271 PAD.n8070 VSS 0.036461f
C7272 PAD.n8071 VSS 0.036461f
C7273 PAD.n8073 VSS 0.036461f
C7274 PAD.n8074 VSS 0.036461f
C7275 PAD.n8075 VSS 0.036461f
C7276 PAD.n8076 VSS 0.036461f
C7277 PAD.n8077 VSS 0.036461f
C7278 PAD.n8078 VSS 0.036461f
C7279 PAD.n8079 VSS 0.036461f
C7280 PAD.n8080 VSS 0.036461f
C7281 PAD.n8082 VSS 0.036461f
C7282 PAD.n8083 VSS 0.036461f
C7283 PAD.n8084 VSS 0.036461f
C7284 PAD.n8085 VSS 0.036461f
C7285 PAD.n8086 VSS 0.036461f
C7286 PAD.n8087 VSS 0.036461f
C7287 PAD.n8088 VSS 0.036461f
C7288 PAD.n8089 VSS 0.036461f
C7289 PAD.n8091 VSS 0.036461f
C7290 PAD.n8092 VSS 0.036461f
C7291 PAD.n8093 VSS 0.036461f
C7292 PAD.n8094 VSS 0.036461f
C7293 PAD.n8095 VSS 0.036461f
C7294 PAD.n8096 VSS 0.036461f
C7295 PAD.n8097 VSS 0.036461f
C7296 PAD.n8098 VSS 0.036461f
C7297 PAD.n8100 VSS 0.036461f
C7298 PAD.n8101 VSS 0.036461f
C7299 PAD.n8102 VSS 0.036461f
C7300 PAD.n8103 VSS 0.036461f
C7301 PAD.n8104 VSS 0.036461f
C7302 PAD.n8105 VSS 0.036461f
C7303 PAD.n8106 VSS 0.036461f
C7304 PAD.n8107 VSS 0.036461f
C7305 PAD.n8109 VSS 0.036461f
C7306 PAD.n8110 VSS 0.036461f
C7307 PAD.n8111 VSS 0.036461f
C7308 PAD.n8112 VSS 0.036461f
C7309 PAD.n8113 VSS 0.036461f
C7310 PAD.n8114 VSS 0.036461f
C7311 PAD.n8115 VSS 0.036461f
C7312 PAD.n8116 VSS 0.036461f
C7313 PAD.n8118 VSS 0.036461f
C7314 PAD.n8119 VSS 0.036461f
C7315 PAD.n8120 VSS 0.036461f
C7316 PAD.n8121 VSS 0.036461f
C7317 PAD.n8122 VSS 0.036461f
C7318 PAD.n8123 VSS 0.036461f
C7319 PAD.n8124 VSS 0.036461f
C7320 PAD.n8125 VSS 0.036461f
C7321 PAD.n8127 VSS 0.036461f
C7322 PAD.n8128 VSS 0.036461f
C7323 PAD.n8129 VSS 0.036461f
C7324 PAD.n8130 VSS 0.036461f
C7325 PAD.n8131 VSS 0.036461f
C7326 PAD.n8132 VSS 0.036461f
C7327 PAD.n8133 VSS 0.036461f
C7328 PAD.n8134 VSS 0.036461f
C7329 PAD.n8136 VSS 0.036461f
C7330 PAD.n8137 VSS 0.036461f
C7331 PAD.n8138 VSS 0.036461f
C7332 PAD.n8139 VSS 0.036461f
C7333 PAD.n8140 VSS 0.036461f
C7334 PAD.n8141 VSS 0.036461f
C7335 PAD.n8142 VSS 0.036461f
C7336 PAD.n8143 VSS 0.036461f
C7337 PAD.n8145 VSS 0.036461f
C7338 PAD.n8146 VSS 0.036461f
C7339 PAD.n8147 VSS 0.036461f
C7340 PAD.n8148 VSS 0.036461f
C7341 PAD.n8149 VSS 0.036461f
C7342 PAD.n8150 VSS 0.036461f
C7343 PAD.n8151 VSS 0.036461f
C7344 PAD.n8152 VSS 0.036461f
C7345 PAD.n8154 VSS 0.036461f
C7346 PAD.n8155 VSS 0.036461f
C7347 PAD.n8156 VSS 0.036461f
C7348 PAD.n8157 VSS 0.036461f
C7349 PAD.n8158 VSS 0.036461f
C7350 PAD.n8159 VSS 0.036461f
C7351 PAD.n8160 VSS 0.023109f
C7352 PAD.n8161 VSS 0.023109f
C7353 PAD.n8163 VSS 0.596934f
C7354 PAD.n8164 VSS 0.542667f
C7355 PAD.n8165 VSS 0.626534f
C7356 PAD.n8166 VSS 0.069765f
C7357 PAD.n8167 VSS 0.050636f
C7358 PAD.n8168 VSS 0.050636f
C7359 PAD.n8169 VSS 0.045199f
C7360 PAD.n8170 VSS 0.046286f
C7361 PAD.n8171 VSS 0.048212f
C7362 PAD.n8172 VSS 0.054012f
C7363 PAD.n8173 VSS 0.054012f
C7364 PAD.n8174 VSS 0.527867f
C7365 PAD.n8175 VSS 0.611734f
C7366 PAD.n8176 VSS 0.03061f
C7367 PAD.n8177 VSS 0.03061f
C7368 PAD.n8178 VSS 0.026734f
C7369 PAD.n8179 VSS 0.033773f
C7370 PAD.n8180 VSS 0.037609f
C7371 PAD.n8181 VSS 0.043062f
C7372 PAD.n8182 VSS 0.043062f
C7373 PAD.n8183 VSS 0.592001f
C7374 PAD.n8184 VSS 0.700534f
C7375 PAD.n8185 VSS 0.611734f
C7376 PAD.n8186 VSS 0.419334f
C7377 PAD.n8187 VSS 0.058513f
C7378 PAD.n8188 VSS 0.058513f
C7379 PAD.n8189 VSS 0.05223f
C7380 PAD.n8190 VSS 0.046286f
C7381 PAD.n8191 VSS 0.041181f
C7382 PAD.n8192 VSS 0.046135f
C7383 PAD.n8193 VSS 0.046135f
C7384 PAD.n8194 VSS 0.419334f
C7385 PAD.n8195 VSS 0.522934f
C7386 PAD.n8196 VSS 0.026114f
C7387 PAD.n8197 VSS 0.026114f
C7388 PAD.n8198 VSS 0.022807f
C7389 PAD.n8199 VSS 0.033773f
C7390 PAD.n8200 VSS 0.041536f
C7391 PAD.n8201 VSS 0.047559f
C7392 PAD.n8202 VSS 0.046175f
C7393 PAD.n8203 VSS 0.046175f
C7394 PAD.n8204 VSS 0.029436f
C7395 PAD.n8205 VSS 0.300934f
C7396 PAD.n8206 VSS 0.027498f
C7397 PAD.n8207 VSS 0.027498f
C7398 PAD.n8208 VSS 0.024015f
C7399 PAD.n8209 VSS 0.033773f
C7400 PAD.n8210 VSS 0.030555f
C7401 PAD.n8211 VSS 0.036461f
C7402 PAD.n8212 VSS 0.036461f
C7403 PAD.n8213 VSS 0.036461f
C7404 PAD.n8214 VSS 0.036461f
C7405 PAD.n8215 VSS 0.036461f
C7406 PAD.n8217 VSS 0.036461f
C7407 PAD.n8218 VSS 0.036461f
C7408 PAD.n8219 VSS 0.036461f
C7409 PAD.n8220 VSS 0.036461f
C7410 PAD.n8221 VSS 0.036461f
C7411 PAD.n8222 VSS 0.036461f
C7412 PAD.n8223 VSS 0.036461f
C7413 PAD.n8224 VSS 0.036461f
C7414 PAD.n8226 VSS 0.036461f
C7415 PAD.n8227 VSS 0.036461f
C7416 PAD.n8228 VSS 0.036461f
C7417 PAD.n8229 VSS 0.036461f
C7418 PAD.n8230 VSS 0.036461f
C7419 PAD.n8231 VSS 0.036461f
C7420 PAD.n8232 VSS 0.036461f
C7421 PAD.n8233 VSS 0.036461f
C7422 PAD.n8235 VSS 0.036461f
C7423 PAD.n8236 VSS 0.036461f
C7424 PAD.n8237 VSS 0.036461f
C7425 PAD.n8238 VSS 0.036461f
C7426 PAD.n8239 VSS 0.036461f
C7427 PAD.n8240 VSS 0.036461f
C7428 PAD.n8241 VSS 0.036461f
C7429 PAD.n8242 VSS 0.036461f
C7430 PAD.n8244 VSS 0.036461f
C7431 PAD.n8245 VSS 0.036461f
C7432 PAD.n8246 VSS 0.036461f
C7433 PAD.n8247 VSS 0.036461f
C7434 PAD.n8248 VSS 0.036461f
C7435 PAD.n8249 VSS 0.036461f
C7436 PAD.n8250 VSS 0.036461f
C7437 PAD.n8251 VSS 0.036461f
C7438 PAD.n8253 VSS 0.036461f
C7439 PAD.n8254 VSS 0.036461f
C7440 PAD.n8255 VSS 0.036461f
C7441 PAD.n8256 VSS 0.036461f
C7442 PAD.n8257 VSS 0.036461f
C7443 PAD.n8258 VSS 0.036461f
C7444 PAD.n8259 VSS 0.036461f
C7445 PAD.n8260 VSS 0.036461f
C7446 PAD.n8262 VSS 0.036461f
C7447 PAD.n8263 VSS 0.036461f
C7448 PAD.n8264 VSS 0.036461f
C7449 PAD.n8265 VSS 0.036461f
C7450 PAD.n8266 VSS 0.036461f
C7451 PAD.n8267 VSS 0.036461f
C7452 PAD.n8268 VSS 0.036461f
C7453 PAD.n8269 VSS 0.036461f
C7454 PAD.n8271 VSS 0.036461f
C7455 PAD.n8272 VSS 0.036461f
C7456 PAD.n8273 VSS 0.036461f
C7457 PAD.n8274 VSS 0.036461f
C7458 PAD.n8275 VSS 0.036461f
C7459 PAD.n8276 VSS 0.036461f
C7460 PAD.n8277 VSS 0.036461f
C7461 PAD.n8278 VSS 0.036461f
C7462 PAD.n8280 VSS 0.036461f
C7463 PAD.n8281 VSS 0.036461f
C7464 PAD.n8282 VSS 0.036461f
C7465 PAD.n8283 VSS 0.036461f
C7466 PAD.n8284 VSS 0.036461f
C7467 PAD.n8285 VSS 0.036461f
C7468 PAD.n8286 VSS 0.036461f
C7469 PAD.n8287 VSS 0.036461f
C7470 PAD.n8289 VSS 0.036461f
C7471 PAD.n8290 VSS 0.036461f
C7472 PAD.n8291 VSS 0.036461f
C7473 PAD.n8292 VSS 0.036461f
C7474 PAD.n8293 VSS 0.036461f
C7475 PAD.n8294 VSS 0.036461f
C7476 PAD.n8295 VSS 0.036461f
C7477 PAD.n8296 VSS 0.036461f
C7478 PAD.n8298 VSS 0.036461f
C7479 PAD.n8299 VSS 0.036461f
C7480 PAD.n8300 VSS 0.036461f
C7481 PAD.n8301 VSS 0.036461f
C7482 PAD.n8302 VSS 0.036461f
C7483 PAD.n8303 VSS 0.036461f
C7484 PAD.n8304 VSS 0.036461f
C7485 PAD.n8305 VSS 0.036461f
C7486 PAD.n8307 VSS 0.036461f
C7487 PAD.n8308 VSS 0.036461f
C7488 PAD.n8309 VSS 0.036461f
C7489 PAD.n8310 VSS 0.036461f
C7490 PAD.n8311 VSS 0.036461f
C7491 PAD.n8312 VSS 0.036461f
C7492 PAD.n8313 VSS 0.036461f
C7493 PAD.n8314 VSS 0.036461f
C7494 PAD.n8316 VSS 0.036461f
C7495 PAD.n8317 VSS 0.036461f
C7496 PAD.n8318 VSS 0.036461f
C7497 PAD.n8319 VSS 0.036461f
C7498 PAD.n8320 VSS 0.036461f
C7499 PAD.n8321 VSS 0.036461f
C7500 PAD.n8322 VSS 0.036461f
C7501 PAD.n8323 VSS 0.036461f
C7502 PAD.n8325 VSS 0.036461f
C7503 PAD.n8326 VSS 0.036461f
C7504 PAD.n8327 VSS 0.036461f
C7505 PAD.n8328 VSS 0.036461f
C7506 PAD.n8329 VSS 0.036461f
C7507 PAD.n8330 VSS 0.036461f
C7508 PAD.n8331 VSS 0.036461f
C7509 PAD.n8332 VSS 0.036461f
C7510 PAD.n8334 VSS 0.036461f
C7511 PAD.n8335 VSS 0.036461f
C7512 PAD.n8336 VSS 0.036461f
C7513 PAD.n8337 VSS 0.036461f
C7514 PAD.n8338 VSS 0.036461f
C7515 PAD.n8339 VSS 0.036461f
C7516 PAD.n8340 VSS 0.036461f
C7517 PAD.n8341 VSS 0.036461f
C7518 PAD.n8343 VSS 0.036461f
C7519 PAD.n8344 VSS 0.036461f
C7520 PAD.n8345 VSS 0.036461f
C7521 PAD.n8346 VSS 0.036461f
C7522 PAD.n8347 VSS 0.036461f
C7523 PAD.n8348 VSS 0.036461f
C7524 PAD.n8349 VSS 0.036461f
C7525 PAD.n8350 VSS 0.036461f
C7526 PAD.n8352 VSS 0.036461f
C7527 PAD.n8353 VSS 0.036461f
C7528 PAD.n8354 VSS 0.036461f
C7529 PAD.n8355 VSS 0.036461f
C7530 PAD.n8356 VSS 0.036461f
C7531 PAD.n8357 VSS 0.036461f
C7532 PAD.n8358 VSS 0.036461f
C7533 PAD.n8359 VSS 0.036461f
C7534 PAD.n8361 VSS 0.036461f
C7535 PAD.n8362 VSS 0.036461f
C7536 PAD.n8363 VSS 0.036461f
C7537 PAD.n8364 VSS 0.036461f
C7538 PAD.n8365 VSS 0.036461f
C7539 PAD.n8366 VSS 0.036461f
C7540 PAD.n8367 VSS 0.036461f
C7541 PAD.n8368 VSS 0.036461f
C7542 PAD.n8370 VSS 0.036461f
C7543 PAD.n8371 VSS 0.036461f
C7544 PAD.n8372 VSS 0.036461f
C7545 PAD.n8373 VSS 0.036461f
C7546 PAD.n8374 VSS 0.036461f
C7547 PAD.n8375 VSS 0.036461f
C7548 PAD.n8376 VSS 0.036461f
C7549 PAD.n8377 VSS 0.036461f
C7550 PAD.n8379 VSS 0.036461f
C7551 PAD.n8380 VSS 0.036461f
C7552 PAD.n8381 VSS 0.036461f
C7553 PAD.n8382 VSS 0.036461f
C7554 PAD.n8383 VSS 0.036461f
C7555 PAD.n8384 VSS 0.036461f
C7556 PAD.n8385 VSS 0.036461f
C7557 PAD.n8386 VSS 0.036461f
C7558 PAD.n8388 VSS 0.036461f
C7559 PAD.n8389 VSS 0.036461f
C7560 PAD.n8390 VSS 0.036461f
C7561 PAD.n8391 VSS 0.036461f
C7562 PAD.n8392 VSS 0.036461f
C7563 PAD.n8393 VSS 0.036461f
C7564 PAD.n8394 VSS 0.023109f
C7565 PAD.n8395 VSS 0.023109f
C7566 PAD.n8397 VSS 0.611734f
C7567 PAD.n8398 VSS 0.276267f
C7568 PAD.n8399 VSS 0.06639f
C7569 PAD.n8400 VSS 0.06639f
C7570 PAD.n8401 VSS 0.059261f
C7571 PAD.n8402 VSS 0.046286f
C7572 PAD.n8403 VSS 0.03415f
C7573 PAD.n8404 VSS 0.062274f
C7574 PAD.n8405 VSS 0.069765f
C7575 PAD.n8406 VSS 0.069765f
C7576 PAD.n8407 VSS 0.424267f
C7577 PAD.n8408 VSS 0.611734f
C7578 PAD.n8409 VSS 0.700534f
C7579 PAD.n8410 VSS 0.335467f
C7580 PAD.n8411 VSS 0.041679f
C7581 PAD.n8412 VSS 0.041679f
C7582 PAD.n8413 VSS 0.036401f
C7583 PAD.n8414 VSS 0.033773f
C7584 PAD.n8415 VSS 0.042895f
C7585 PAD.n8416 VSS 0.027942f
C7586 PAD.n8417 VSS 0.031994f
C7587 PAD.n8418 VSS 0.031994f
C7588 PAD.n8419 VSS 0.424267f
C7589 PAD.n8420 VSS 0.567334f
C7590 PAD.n8421 VSS 0.039384f
C7591 PAD.n8422 VSS 0.039384f
C7592 PAD.n8423 VSS 0.035155f
C7593 PAD.n8424 VSS 0.046286f
C7594 PAD.n8425 VSS 0.058256f
C7595 PAD.n8426 VSS 0.042186f
C7596 PAD.n8427 VSS 0.062274f
C7597 PAD.n8428 VSS 0.069765f
C7598 PAD.n8429 VSS 0.069765f
C7599 PAD.n8430 VSS 0.700534f
C7600 PAD.n8431 VSS 0.4736f
C7601 PAD.n8432 VSS 0.037182f
C7602 PAD.n8433 VSS 0.037182f
C7603 PAD.n8434 VSS 0.029436f
C7604 PAD.n8435 VSS 0.03649f
C7605 PAD.n8436 VSS 0.031869f
C7606 PAD.n8437 VSS 0.033773f
C7607 PAD.n8438 VSS 0.030555f
C7608 PAD.n8439 VSS 0.036461f
C7609 PAD.n8440 VSS 0.036461f
C7610 PAD.n8441 VSS 0.036461f
C7611 PAD.n8443 VSS 0.023109f
C7612 PAD.n8444 VSS 0.054266f
C7613 PAD.n8445 VSS 0.661068f
C7614 PAD.n8446 VSS 0.057388f
C7615 PAD.n8447 VSS 0.057388f
C7616 PAD.n8448 VSS 0.051225f
C7617 PAD.n8449 VSS 0.062274f
C7618 PAD.n8450 VSS 0.049216f
C7619 PAD.n8451 VSS 0.055137f
C7620 PAD.n8452 VSS 0.055137f
C7621 PAD.n8453 VSS 0.582134f
C7622 PAD.n8454 VSS 0.611734f
C7623 PAD.n8455 VSS 0.049115f
C7624 PAD.n8456 VSS 0.032686f
C7625 PAD.n8457 VSS 0.032686f
C7626 PAD.n8458 VSS 0.029436f
C7627 PAD.n8459 VSS 0.040987f
C7628 PAD.n8460 VSS 0.035797f
C7629 PAD.n8461 VSS 0.033773f
C7630 PAD.n8462 VSS 0.030555f
C7631 PAD.n8463 VSS 0.036461f
C7632 PAD.n8464 VSS 0.036461f
C7633 PAD.n8465 VSS 0.036461f
C7634 PAD.n8467 VSS 0.023109f
C7635 PAD.n8468 VSS 0.212133f
C7636 PAD.n8469 VSS 0.582134f
C7637 PAD.n8470 VSS 0.049511f
C7638 PAD.n8471 VSS 0.049511f
C7639 PAD.n8472 VSS 0.021343f
C7640 PAD.n8473 VSS 8.78048f
C7641 PAD.n8474 VSS 0.053987f
C7642 PAD.n8475 VSS 0.056247f
C7643 PAD.n8476 VSS 0.063014f
C7644 PAD.n8477 VSS 0.063014f
C7645 PAD.n8478 VSS 0.424267f
C7646 PAD.n8479 VSS 0.611734f
C7647 PAD.n8480 VSS 0.049115f
C7648 PAD.n8481 VSS 0.028189f
C7649 PAD.n8482 VSS 0.028189f
C7650 PAD.n8483 VSS 0.024619f
C7651 PAD.n8484 VSS 0.039724f
C7652 PAD.n8485 VSS 0.033773f
C7653 PAD.n8486 VSS 0.030555f
C7654 PAD.n8487 VSS 0.036461f
C7655 PAD.n8488 VSS 0.036461f
C7656 PAD.n8489 VSS 0.036461f
C7657 PAD.n8491 VSS 0.023109f
C7658 PAD.n8492 VSS 0.478534f
C7659 PAD.n8493 VSS 0.424267f
C7660 PAD.n8494 VSS 0.041634f
C7661 PAD.n8495 VSS 0.041634f
C7662 PAD.n8496 VSS 0.037163f
C7663 PAD.n8497 VSS 0.062274f
C7664 PAD.n8498 VSS 0.032141f
C7665 PAD.n8499 VSS 0.062274f
C7666 PAD.n8500 VSS 0.069765f
C7667 PAD.n8501 VSS 0.069765f
C7668 PAD.n8502 VSS 0.3108f
C7669 PAD.n8503 VSS 0.611734f
C7670 PAD.n8504 VSS 0.048251f
C7671 PAD.n8505 VSS 0.048251f
C7672 PAD.n8506 VSS 0.029436f
C7673 PAD.n8507 VSS 0.025422f
C7674 PAD.n8508 VSS 0.025422f
C7675 PAD.n8509 VSS 0.022203f
C7676 PAD.n8510 VSS 0.033773f
C7677 PAD.n8511 VSS 0.030555f
C7678 PAD.n8512 VSS 0.036461f
C7679 PAD.n8513 VSS 0.036461f
C7680 PAD.n8514 VSS 0.036461f
C7681 PAD.n8516 VSS 0.023109f
C7682 PAD.n8517 VSS 0.567334f
C7683 PAD.n8518 VSS 0.611734f
C7684 PAD.n8519 VSS 0.389734f
C7685 PAD.n8520 VSS 0.06864f
C7686 PAD.n8521 VSS 0.06864f
C7687 PAD.n8522 VSS 0.061269f
C7688 PAD.n8523 VSS 0.062274f
C7689 PAD.n8524 VSS 0.039172f
C7690 PAD.n8525 VSS 0.043885f
C7691 PAD.n8526 VSS 0.043885f
C7692 PAD.n8527 VSS 0.384801f
C7693 PAD.n8528 VSS 0.036461f
C7694 PAD.n8529 VSS 0.036461f
C7695 PAD.n8530 VSS 0.036461f
C7696 PAD.n8531 VSS 0.036461f
C7697 PAD.n8532 VSS 0.036461f
C7698 PAD.n8533 VSS 0.036461f
C7699 PAD.n8534 VSS 0.036461f
C7700 PAD.n8535 VSS 0.036461f
C7701 PAD.n8536 VSS 0.036461f
C7702 PAD.n8537 VSS 0.036461f
C7703 PAD.n8538 VSS 0.036461f
C7704 PAD.n8539 VSS 0.036461f
C7705 PAD.n8540 VSS 0.036461f
C7706 PAD.n8541 VSS 0.036461f
C7707 PAD.n8542 VSS 0.036461f
C7708 PAD.n8543 VSS 0.036461f
C7709 PAD.n8544 VSS 0.036461f
C7710 PAD.n8545 VSS 0.036461f
C7711 PAD.n8546 VSS 0.036461f
C7712 PAD.n8547 VSS 0.036461f
C7713 PAD.n8548 VSS 0.036461f
C7714 PAD.n8549 VSS 0.036461f
C7715 PAD.n8550 VSS 0.036461f
C7716 PAD.n8551 VSS 0.036461f
C7717 PAD.n8552 VSS 0.036461f
C7718 PAD.n8553 VSS 0.036461f
C7719 PAD.n8554 VSS 0.036461f
C7720 PAD.n8555 VSS 0.036461f
C7721 PAD.n8556 VSS 0.036461f
C7722 PAD.n8557 VSS 0.036461f
C7723 PAD.n8558 VSS 0.036461f
C7724 PAD.n8559 VSS 0.036461f
C7725 PAD.n8560 VSS 0.036461f
C7726 PAD.n8561 VSS 0.036461f
C7727 PAD.n8562 VSS 0.036461f
C7728 PAD.n8563 VSS 0.036461f
C7729 PAD.n8564 VSS 0.036461f
C7730 PAD.n8565 VSS 0.036461f
C7731 PAD.n8566 VSS 0.036461f
C7732 PAD.n8567 VSS 0.036461f
C7733 PAD.n8568 VSS 0.036461f
C7734 PAD.n8569 VSS 0.036461f
C7735 PAD.n8570 VSS 0.023109f
C7736 PAD.n8571 VSS 0.023109f
C7737 PAD.n8572 VSS 0.036461f
C7738 PAD.n8574 VSS 0.036461f
C7739 PAD.n8575 VSS 0.036461f
C7740 PAD.n8576 VSS 0.036461f
C7741 PAD.n8577 VSS 0.036461f
C7742 PAD.n8578 VSS 0.036461f
C7743 PAD.n8579 VSS 0.036461f
C7744 PAD.n8580 VSS 0.036461f
C7745 PAD.n8582 VSS 0.036461f
C7746 PAD.n8583 VSS 0.036461f
C7747 PAD.n8584 VSS 0.036461f
C7748 PAD.n8586 VSS 0.036461f
C7749 PAD.n8587 VSS 0.036461f
C7750 PAD.n8588 VSS 0.036461f
C7751 PAD.n8589 VSS 0.036461f
C7752 PAD.n8590 VSS 0.036461f
C7753 PAD.n8591 VSS 0.036461f
C7754 PAD.n8592 VSS 0.036461f
C7755 PAD.n8594 VSS 0.036461f
C7756 PAD.n8595 VSS 0.036461f
C7757 PAD.n8596 VSS 0.036461f
C7758 PAD.n8598 VSS 0.036461f
C7759 PAD.n8599 VSS 0.036461f
C7760 PAD.n8600 VSS 0.036461f
C7761 PAD.n8601 VSS 0.036461f
C7762 PAD.n8602 VSS 0.036461f
C7763 PAD.n8603 VSS 0.036461f
C7764 PAD.n8604 VSS 0.036461f
C7765 PAD.n8606 VSS 0.036461f
C7766 PAD.n8607 VSS 0.036461f
C7767 PAD.n8608 VSS 0.036461f
C7768 PAD.n8610 VSS 0.036461f
C7769 PAD.n8611 VSS 0.036461f
C7770 PAD.n8612 VSS 0.036461f
C7771 PAD.n8613 VSS 0.036461f
C7772 PAD.n8614 VSS 0.036461f
C7773 PAD.n8615 VSS 0.036461f
C7774 PAD.n8616 VSS 0.036461f
C7775 PAD.n8618 VSS 0.036461f
C7776 PAD.n8619 VSS 0.036461f
C7777 PAD.n8620 VSS 0.036461f
C7778 PAD.n8622 VSS 0.036461f
C7779 PAD.n8623 VSS 0.036461f
C7780 PAD.n8624 VSS 0.036461f
C7781 PAD.n8625 VSS 0.036461f
C7782 PAD.n8626 VSS 0.036461f
C7783 PAD.n8627 VSS 0.036461f
C7784 PAD.n8628 VSS 0.036461f
C7785 PAD.n8630 VSS 0.036461f
C7786 PAD.n8631 VSS 0.036461f
C7787 PAD.n8632 VSS 0.036461f
C7788 PAD.n8634 VSS 0.036461f
C7789 PAD.n8635 VSS 0.036461f
C7790 PAD.n8636 VSS 0.036461f
C7791 PAD.n8637 VSS 0.036461f
C7792 PAD.n8638 VSS 0.036461f
C7793 PAD.n8639 VSS 0.036461f
C7794 PAD.n8640 VSS 0.036461f
C7795 PAD.n8642 VSS 0.036461f
C7796 PAD.n8643 VSS 0.036461f
C7797 PAD.n8644 VSS 0.036461f
C7798 PAD.n8646 VSS 0.036461f
C7799 PAD.n8647 VSS 0.036461f
C7800 PAD.n8648 VSS 0.036461f
C7801 PAD.n8649 VSS 0.036461f
C7802 PAD.n8650 VSS 0.036461f
C7803 PAD.n8651 VSS 0.036461f
C7804 PAD.n8652 VSS 0.036461f
C7805 PAD.n8654 VSS 0.036461f
C7806 PAD.n8655 VSS 0.036461f
C7807 PAD.n8656 VSS 0.036461f
C7808 PAD.n8658 VSS 0.036461f
C7809 PAD.n8659 VSS 0.036461f
C7810 PAD.n8660 VSS 0.036461f
C7811 PAD.n8661 VSS 0.036461f
C7812 PAD.n8662 VSS 0.036461f
C7813 PAD.n8663 VSS 0.036461f
C7814 PAD.n8664 VSS 0.036461f
C7815 PAD.n8666 VSS 0.036461f
C7816 PAD.n8667 VSS 0.036461f
C7817 PAD.n8668 VSS 0.036461f
C7818 PAD.n8670 VSS 0.036461f
C7819 PAD.n8671 VSS 0.036461f
C7820 PAD.n8672 VSS 0.036461f
C7821 PAD.n8673 VSS 0.036461f
C7822 PAD.n8674 VSS 0.036461f
C7823 PAD.n8675 VSS 0.036461f
C7824 PAD.n8676 VSS 0.036461f
C7825 PAD.n8678 VSS 0.036461f
C7826 PAD.n8679 VSS 0.036461f
C7827 PAD.n8680 VSS 0.036461f
C7828 PAD.n8682 VSS 0.036461f
C7829 PAD.n8683 VSS 0.036461f
C7830 PAD.n8684 VSS 0.036461f
C7831 PAD.n8685 VSS 0.036461f
C7832 PAD.n8686 VSS 0.036461f
C7833 PAD.n8687 VSS 0.036461f
C7834 PAD.n8688 VSS 0.036461f
C7835 PAD.n8690 VSS 0.036461f
C7836 PAD.n8691 VSS 0.036461f
C7837 PAD.n8692 VSS 0.036461f
C7838 PAD.n8694 VSS 0.036461f
C7839 PAD.n8695 VSS 0.036461f
C7840 PAD.n8696 VSS 0.036461f
C7841 PAD.n8697 VSS 0.036461f
C7842 PAD.n8698 VSS 0.036461f
C7843 PAD.n8699 VSS 0.036461f
C7844 PAD.n8700 VSS 0.036461f
C7845 PAD.n8702 VSS 0.036461f
C7846 PAD.n8703 VSS 0.036461f
C7847 PAD.n8704 VSS 0.036461f
C7848 PAD.n8706 VSS 0.036461f
C7849 PAD.n8707 VSS 0.036461f
C7850 PAD.n8708 VSS 0.036461f
C7851 PAD.n8709 VSS 0.036461f
C7852 PAD.n8710 VSS 0.036461f
C7853 PAD.n8711 VSS 0.036461f
C7854 PAD.n8712 VSS 0.036461f
C7855 PAD.n8714 VSS 0.036461f
C7856 PAD.n8715 VSS 0.036461f
C7857 PAD.n8716 VSS 0.036461f
C7858 PAD.n8718 VSS 0.036461f
C7859 PAD.n8719 VSS 0.036461f
C7860 PAD.n8720 VSS 0.036461f
C7861 PAD.n8721 VSS 0.036461f
C7862 PAD.n8722 VSS 0.036461f
C7863 PAD.n8723 VSS 0.036461f
C7864 PAD.n8724 VSS 0.036461f
C7865 PAD.n8726 VSS 0.036461f
C7866 PAD.n8727 VSS 0.036461f
C7867 PAD.n8728 VSS 0.036461f
C7868 PAD.n8730 VSS 0.036461f
C7869 PAD.n8731 VSS 0.036461f
C7870 PAD.n8732 VSS 0.036461f
C7871 PAD.n8733 VSS 0.036461f
C7872 PAD.n8734 VSS 0.036461f
C7873 PAD.n8735 VSS 0.036461f
C7874 PAD.n8736 VSS 0.036461f
C7875 PAD.n8738 VSS 0.036461f
C7876 PAD.n8739 VSS 0.036461f
C7877 PAD.n8740 VSS 0.036461f
C7878 PAD.n8742 VSS 0.036461f
C7879 PAD.n8743 VSS 0.036461f
C7880 PAD.n8744 VSS 0.036461f
C7881 PAD.n8745 VSS 0.036461f
C7882 PAD.n8746 VSS 0.036461f
C7883 PAD.n8747 VSS 0.036461f
C7884 PAD.n8748 VSS 0.036461f
C7885 PAD.n8750 VSS 0.036461f
C7886 PAD.n8751 VSS 0.036461f
C7887 PAD.n8752 VSS 0.036461f
C7888 PAD.n8754 VSS 0.036461f
C7889 PAD.n8755 VSS 0.036461f
C7890 PAD.n8756 VSS 0.036461f
C7891 PAD.n8757 VSS 0.036461f
C7892 PAD.n8758 VSS 0.036461f
C7893 PAD.n8759 VSS 0.036461f
C7894 PAD.n8760 VSS 0.036461f
C7895 PAD.n8762 VSS 0.036461f
C7896 PAD.n8763 VSS 0.036461f
C7897 PAD.n8764 VSS 0.036461f
C7898 PAD.n8766 VSS 0.036461f
C7899 PAD.n8767 VSS 0.036461f
C7900 PAD.n8768 VSS 0.036461f
C7901 PAD.n8769 VSS 0.036461f
C7902 PAD.n8770 VSS 0.036461f
C7903 PAD.n8771 VSS 0.036461f
C7904 PAD.n8772 VSS 0.036461f
C7905 PAD.n8774 VSS 0.036461f
C7906 PAD.n8775 VSS 0.036461f
C7907 PAD.n8776 VSS 0.036461f
C7908 PAD.n8778 VSS 0.036461f
C7909 PAD.n8779 VSS 0.036461f
C7910 PAD.n8780 VSS 0.036461f
C7911 PAD.n8781 VSS 0.036461f
C7912 PAD.n8782 VSS 0.036461f
C7913 PAD.n8783 VSS 0.036461f
C7914 PAD.n8784 VSS 0.036461f
C7915 PAD.n8786 VSS 0.036461f
C7916 PAD.n8787 VSS 0.036461f
C7917 PAD.n8788 VSS 0.036461f
C7918 PAD.n8790 VSS 0.036461f
C7919 PAD.n8791 VSS 0.036461f
C7920 PAD.n8792 VSS 0.036461f
C7921 PAD.n8793 VSS 0.036461f
C7922 PAD.n8794 VSS 0.036461f
C7923 PAD.n8795 VSS 0.036461f
C7924 PAD.n8796 VSS 0.036461f
C7925 PAD.n8798 VSS 0.036461f
C7926 PAD.n8799 VSS 0.036461f
C7927 PAD.n8800 VSS 0.036461f
C7928 PAD.n8802 VSS 0.036461f
C7929 PAD.n8803 VSS 0.036461f
C7930 PAD.n8804 VSS 0.036461f
C7931 PAD.n8805 VSS 0.036461f
C7932 PAD.n8806 VSS 0.036461f
C7933 PAD.n8807 VSS 0.036461f
C7934 PAD.n8808 VSS 0.036461f
C7935 PAD.n8810 VSS 0.036461f
C7936 PAD.n8811 VSS 0.036461f
C7937 PAD.n8813 VSS 0.036461f
C7938 PAD.n8814 VSS 0.036461f
C7939 PAD.n8815 VSS 0.036461f
C7940 PAD.n8816 VSS 0.036461f
C7941 PAD.n8817 VSS 0.03338f
C7942 PAD.n8818 VSS 0.023109f
C7943 PAD.n8819 VSS 0.023109f
C7944 PAD.n8821 VSS 0.389734f
C7945 PAD.n8822 VSS 0.4144f
C7946 PAD.n8823 VSS 0.043754f
C7947 PAD.n8824 VSS 0.043754f
C7948 PAD.n8825 VSS 0.038213f
C7949 PAD.n8826 VSS 0.033773f
C7950 PAD.n8827 VSS 0.02613f
C7951 PAD.n8828 VSS 0.042895f
C7952 PAD.n8829 VSS 0.049115f
C7953 PAD.n8830 VSS 0.049115f
C7954 PAD.n8831 VSS 0.611734f
C7955 PAD.n8832 VSS 0.508134f
C7956 PAD.n8833 VSS 0.060763f
C7957 PAD.n8834 VSS 0.060763f
C7958 PAD.n8835 VSS 0.054238f
C7959 PAD.n8836 VSS 0.062274f
C7960 PAD.n8837 VSS 0.036461f
C7961 PAD.n8838 VSS 0.036461f
C7962 PAD.n8839 VSS 0.036461f
C7963 PAD.n8841 VSS 0.036461f
C7964 PAD.n8842 VSS 0.036461f
C7965 PAD.n8843 VSS 0.036461f
C7966 PAD.n8844 VSS 0.036461f
C7967 PAD.n8846 VSS 0.036461f
C7968 PAD.n8847 VSS 0.036461f
C7969 PAD.n8848 VSS 0.036461f
C7970 PAD.n8849 VSS 0.036461f
C7971 PAD.n8851 VSS 0.036461f
C7972 PAD.n8852 VSS 0.036461f
C7973 PAD.n8853 VSS 0.036461f
C7974 PAD.n8854 VSS 0.036461f
C7975 PAD.n8856 VSS 0.036461f
C7976 PAD.n8857 VSS 0.036461f
C7977 PAD.n8858 VSS 0.036461f
C7978 PAD.n8859 VSS 0.036461f
C7979 PAD.n8861 VSS 0.036461f
C7980 PAD.n8862 VSS 0.036461f
C7981 PAD.n8863 VSS 0.036461f
C7982 PAD.n8864 VSS 0.036461f
C7983 PAD.n8866 VSS 0.036461f
C7984 PAD.n8867 VSS 0.036461f
C7985 PAD.n8868 VSS 0.036461f
C7986 PAD.n8869 VSS 0.036461f
C7987 PAD.n8871 VSS 0.036461f
C7988 PAD.n8872 VSS 0.036461f
C7989 PAD.n8873 VSS 0.036461f
C7990 PAD.n8874 VSS 0.036461f
C7991 PAD.n8876 VSS 0.036461f
C7992 PAD.n8877 VSS 0.036461f
C7993 PAD.n8878 VSS 0.036461f
C7994 PAD.n8879 VSS 0.036461f
C7995 PAD.n8881 VSS 0.036461f
C7996 PAD.n8882 VSS 0.036461f
C7997 PAD.n8883 VSS 0.036461f
C7998 PAD.n8884 VSS 0.036461f
C7999 PAD.n8886 VSS 0.036461f
C8000 PAD.n8887 VSS 0.036461f
C8001 PAD.n8888 VSS 0.036461f
C8002 PAD.n8889 VSS 0.036461f
C8003 PAD.n8891 VSS 0.036461f
C8004 PAD.n8892 VSS 0.036461f
C8005 PAD.n8893 VSS 0.036461f
C8006 PAD.n8894 VSS 0.036461f
C8007 PAD.n8896 VSS 0.036461f
C8008 PAD.n8897 VSS 0.036461f
C8009 PAD.n8898 VSS 0.036461f
C8010 PAD.n8899 VSS 0.036461f
C8011 PAD.n8901 VSS 0.036461f
C8012 PAD.n8902 VSS 0.036461f
C8013 PAD.n8903 VSS 0.036461f
C8014 PAD.n8904 VSS 0.036461f
C8015 PAD.n8906 VSS 0.036461f
C8016 PAD.n8907 VSS 0.036461f
C8017 PAD.n8908 VSS 0.036461f
C8018 PAD.n8909 VSS 0.036461f
C8019 PAD.n8911 VSS 0.036461f
C8020 PAD.n8912 VSS 0.036461f
C8021 PAD.n8913 VSS 0.036461f
C8022 PAD.n8914 VSS 0.036461f
C8023 PAD.n8916 VSS 0.036461f
C8024 PAD.n8917 VSS 0.036461f
C8025 PAD.n8918 VSS 0.036461f
C8026 PAD.n8919 VSS 0.036461f
C8027 PAD.n8921 VSS 0.036461f
C8028 PAD.n8922 VSS 0.036461f
C8029 PAD.n8923 VSS 0.036461f
C8030 PAD.n8924 VSS 0.036461f
C8031 PAD.n8926 VSS 0.036461f
C8032 PAD.n8927 VSS 0.036461f
C8033 PAD.n8928 VSS 0.036461f
C8034 PAD.n8929 VSS 0.036461f
C8035 PAD.n8931 VSS 0.036461f
C8036 PAD.n8932 VSS 0.036461f
C8037 PAD.n8933 VSS 0.036461f
C8038 PAD.n8934 VSS 0.036461f
C8039 PAD.n8936 VSS 0.036461f
C8040 PAD.n8937 VSS 0.036461f
C8041 PAD.n8939 VSS 0.036461f
C8042 PAD.n8940 VSS 0.036461f
C8043 PAD.n8941 VSS 0.036461f
C8044 PAD.n8942 VSS 0.036461f
C8045 PAD.n8943 VSS 0.036461f
C8046 PAD.n8944 VSS 0.036461f
C8047 PAD.n8945 VSS 0.036461f
C8048 PAD.n8946 VSS 0.036461f
C8049 PAD.n8948 VSS 0.036461f
C8050 PAD.n8949 VSS 0.036461f
C8051 PAD.n8950 VSS 0.036461f
C8052 PAD.n8951 VSS 0.036461f
C8053 PAD.n8952 VSS 0.036461f
C8054 PAD.n8953 VSS 0.036461f
C8055 PAD.n8954 VSS 0.036461f
C8056 PAD.n8955 VSS 0.036461f
C8057 PAD.n8957 VSS 0.036461f
C8058 PAD.n8958 VSS 0.036461f
C8059 PAD.n8959 VSS 0.036461f
C8060 PAD.n8960 VSS 0.036461f
C8061 PAD.n8961 VSS 0.036461f
C8062 PAD.n8962 VSS 0.036461f
C8063 PAD.n8963 VSS 0.036461f
C8064 PAD.n8964 VSS 0.036461f
C8065 PAD.n8966 VSS 0.036461f
C8066 PAD.n8967 VSS 0.036461f
C8067 PAD.n8968 VSS 0.036461f
C8068 PAD.n8969 VSS 0.036461f
C8069 PAD.n8970 VSS 0.036461f
C8070 PAD.n8971 VSS 0.036461f
C8071 PAD.n8972 VSS 0.036461f
C8072 PAD.n8973 VSS 0.036461f
C8073 PAD.n8975 VSS 0.036461f
C8074 PAD.n8976 VSS 0.036461f
C8075 PAD.n8977 VSS 0.036461f
C8076 PAD.n8978 VSS 0.036461f
C8077 PAD.n8979 VSS 0.036461f
C8078 PAD.n8980 VSS 0.036461f
C8079 PAD.n8981 VSS 0.036461f
C8080 PAD.n8982 VSS 0.036461f
C8081 PAD.n8984 VSS 0.036461f
C8082 PAD.n8985 VSS 0.036461f
C8083 PAD.n8986 VSS 0.036461f
C8084 PAD.n8987 VSS 0.036461f
C8085 PAD.n8988 VSS 0.036461f
C8086 PAD.n8989 VSS 0.036461f
C8087 PAD.n8990 VSS 0.036461f
C8088 PAD.n8991 VSS 0.036461f
C8089 PAD.n8993 VSS 0.036461f
C8090 PAD.n8994 VSS 0.036461f
C8091 PAD.n8995 VSS 0.036461f
C8092 PAD.n8996 VSS 0.036461f
C8093 PAD.n8997 VSS 0.036461f
C8094 PAD.n8998 VSS 0.036461f
C8095 PAD.n8999 VSS 0.036461f
C8096 PAD.n9000 VSS 0.036461f
C8097 PAD.n9002 VSS 0.036461f
C8098 PAD.n9003 VSS 0.036461f
C8099 PAD.n9004 VSS 0.036461f
C8100 PAD.n9005 VSS 0.036461f
C8101 PAD.n9006 VSS 0.036461f
C8102 PAD.n9007 VSS 0.036461f
C8103 PAD.n9008 VSS 0.036461f
C8104 PAD.n9009 VSS 0.036461f
C8105 PAD.n9011 VSS 0.036461f
C8106 PAD.n9012 VSS 0.036461f
C8107 PAD.n9013 VSS 0.036461f
C8108 PAD.n9014 VSS 0.036461f
C8109 PAD.n9015 VSS 0.036461f
C8110 PAD.n9016 VSS 0.036461f
C8111 PAD.n9017 VSS 0.036461f
C8112 PAD.n9018 VSS 0.036461f
C8113 PAD.n9020 VSS 0.036461f
C8114 PAD.n9021 VSS 0.036461f
C8115 PAD.n9022 VSS 0.036461f
C8116 PAD.n9023 VSS 0.036461f
C8117 PAD.n9024 VSS 0.036461f
C8118 PAD.n9025 VSS 0.036461f
C8119 PAD.n9026 VSS 0.036461f
C8120 PAD.n9027 VSS 0.036461f
C8121 PAD.n9029 VSS 0.036461f
C8122 PAD.n9030 VSS 0.036461f
C8123 PAD.n9031 VSS 0.036461f
C8124 PAD.n9032 VSS 0.036461f
C8125 PAD.n9033 VSS 0.036461f
C8126 PAD.n9034 VSS 0.036461f
C8127 PAD.n9035 VSS 0.036461f
C8128 PAD.n9036 VSS 0.036461f
C8129 PAD.n9038 VSS 0.036461f
C8130 PAD.n9039 VSS 0.036461f
C8131 PAD.n9040 VSS 0.036461f
C8132 PAD.n9041 VSS 0.036461f
C8133 PAD.n9042 VSS 0.036461f
C8134 PAD.n9043 VSS 0.036461f
C8135 PAD.n9044 VSS 0.036461f
C8136 PAD.n9045 VSS 0.036461f
C8137 PAD.n9047 VSS 0.036461f
C8138 PAD.n9048 VSS 0.036461f
C8139 PAD.n9049 VSS 0.036461f
C8140 PAD.n9050 VSS 0.036461f
C8141 PAD.n9051 VSS 0.036461f
C8142 PAD.n9052 VSS 0.036461f
C8143 PAD.n9053 VSS 0.036461f
C8144 PAD.n9054 VSS 0.036461f
C8145 PAD.n9056 VSS 0.036461f
C8146 PAD.n9057 VSS 0.036461f
C8147 PAD.n9058 VSS 0.036461f
C8148 PAD.n9059 VSS 0.036461f
C8149 PAD.n9060 VSS 0.036461f
C8150 PAD.n9061 VSS 0.036461f
C8151 PAD.n9062 VSS 0.036461f
C8152 PAD.n9063 VSS 0.036461f
C8153 PAD.n9065 VSS 0.036461f
C8154 PAD.n9066 VSS 0.036461f
C8155 PAD.n9067 VSS 0.036461f
C8156 PAD.n9068 VSS 0.036461f
C8157 PAD.n9069 VSS 0.036461f
C8158 PAD.n9070 VSS 0.036461f
C8159 PAD.n9071 VSS 0.036461f
C8160 PAD.n9072 VSS 0.036461f
C8161 PAD.n9074 VSS 0.036461f
C8162 PAD.n9075 VSS 0.036461f
C8163 PAD.n9076 VSS 0.036461f
C8164 PAD.n9077 VSS 0.036461f
C8165 PAD.n9078 VSS 0.036461f
C8166 PAD.n9079 VSS 0.036461f
C8167 PAD.n9080 VSS 0.036461f
C8168 PAD.n9081 VSS 0.036461f
C8169 PAD.n9083 VSS 0.036461f
C8170 PAD.n9084 VSS 0.036461f
C8171 PAD.n9085 VSS 0.036461f
C8172 PAD.n9086 VSS 0.036461f
C8173 PAD.n9087 VSS 0.036461f
C8174 PAD.n9088 VSS 0.036461f
C8175 PAD.n9089 VSS 0.036461f
C8176 PAD.n9090 VSS 0.036461f
C8177 PAD.n9092 VSS 0.036461f
C8178 PAD.n9093 VSS 0.036461f
C8179 PAD.n9094 VSS 0.036461f
C8180 PAD.n9095 VSS 0.036461f
C8181 PAD.n9096 VSS 0.036461f
C8182 PAD.n9097 VSS 0.036461f
C8183 PAD.n9098 VSS 0.036461f
C8184 PAD.n9099 VSS 0.036461f
C8185 PAD.n9101 VSS 0.036461f
C8186 PAD.n9102 VSS 0.036461f
C8187 PAD.n9103 VSS 0.036461f
C8188 PAD.n9104 VSS 0.036461f
C8189 PAD.n9105 VSS 0.036461f
C8190 PAD.n9106 VSS 0.036461f
C8191 PAD.n9107 VSS 0.036461f
C8192 PAD.n9108 VSS 0.036461f
C8193 PAD.n9110 VSS 0.036461f
C8194 PAD.n9111 VSS 0.036461f
C8195 PAD.n9112 VSS 0.036461f
C8196 PAD.n9113 VSS 0.036461f
C8197 PAD.n9114 VSS 0.036461f
C8198 PAD.n9115 VSS 0.036461f
C8199 PAD.n9117 VSS 0.036461f
C8200 PAD.n9118 VSS 0.036461f
C8201 PAD.n9119 VSS 0.023109f
C8202 PAD.n9120 VSS 0.03338f
C8203 PAD.n9121 VSS 0.052887f
C8204 PAD.n9122 VSS 0.052887f
C8205 PAD.n9123 VSS 0.047208f
C8206 PAD.n9124 VSS 0.046286f
C8207 PAD.n9125 VSS 0.046203f
C8208 PAD.n9126 VSS 0.051761f
C8209 PAD.n9127 VSS 0.051761f
C8210 PAD.n9128 VSS 0.621601f
C8211 PAD.n9129 VSS 0.611734f
C8212 PAD.n9130 VSS 0.034415f
C8213 PAD.n9131 VSS 0.034415f
C8214 PAD.n9132 VSS 0.030057f
C8215 PAD.n9133 VSS 0.033773f
C8216 PAD.n9134 VSS 0.030555f
C8217 PAD.n9135 VSS 0.036461f
C8218 PAD.n9136 VSS 0.036461f
C8219 PAD.n9137 VSS 0.036461f
C8220 PAD.n9139 VSS 0.023109f
C8221 PAD.n9140 VSS 0.611734f
C8222 PAD.n9141 VSS 0.621601f
C8223 PAD.n9142 VSS 0.611734f
C8224 PAD.n9143 VSS 0.636401f
C8225 PAD.n9144 VSS 0.059638f
C8226 PAD.n9145 VSS 0.059638f
C8227 PAD.n9146 VSS 0.053234f
C8228 PAD.n9147 VSS 0.046286f
C8229 PAD.n9148 VSS 0.040177f
C8230 PAD.n9149 VSS 0.04501f
C8231 PAD.n9150 VSS 0.04501f
C8232 PAD.n9151 VSS 0.636401f
C8233 PAD.n9152 VSS 0.5328f
C8234 PAD.n9153 VSS 0.034761f
C8235 PAD.n9154 VSS 0.034761f
C8236 PAD.n9155 VSS 0.030359f
C8237 PAD.n9156 VSS 0.033773f
C8238 PAD.n9157 VSS 0.033984f
C8239 PAD.n9158 VSS 0.038912f
C8240 PAD.n9159 VSS 0.038912f
C8241 PAD.n9160 VSS 0.444f
C8242 PAD.n9161 VSS 0.700534f
C8243 PAD.n9162 VSS 0.611734f
C8244 PAD.n9163 VSS 0.493334f
C8245 PAD.n9164 VSS 0.067515f
C8246 PAD.n9165 VSS 0.067515f
C8247 PAD.n9166 VSS 0.060265f
C8248 PAD.n9167 VSS 0.046286f
C8249 PAD.n9168 VSS 14.5427f
C8250 PAD.n9169 VSS 0.062274f
C8251 PAD.n9170 VSS 0.055745f
C8252 PAD.n9171 VSS 8.779059f
C8253 PAD.n9172 VSS 0.008538f
C8254 PAD.n9173 VSS 0.037133f
C8255 PAD.n9174 VSS 0.037133f
C8256 PAD.n9175 VSS 0.493334f
C8257 PAD.n9176 VSS 0.409467f
C8258 PAD.n9177 VSS 0.030265f
C8259 PAD.n9178 VSS 0.030265f
C8260 PAD.n9179 VSS 0.026432f
C8261 PAD.n9180 VSS 0.033773f
C8262 PAD.n9181 VSS 0.037911f
C8263 PAD.n9182 VSS 0.043408f
C8264 PAD.n9183 VSS 0.043408f
C8265 PAD.n9184 VSS 0.320667f
C8266 PAD.n9185 VSS 0.700534f
C8267 PAD.n9186 VSS 0.611734f
C8268 PAD.n9187 VSS 0.389734f
C8269 PAD.n9188 VSS 0.069765f
C8270 PAD.n9189 VSS 0.039761f
C8271 PAD.n9190 VSS 0.040509f
C8272 PAD.n9191 VSS 0.040509f
C8273 PAD.n9192 VSS 0.04319f
C8274 PAD.n9193 VSS 0.062274f
C8275 PAD.n9194 VSS 0.057252f
C8276 PAD.n9195 VSS 0.064139f
C8277 PAD.n9196 VSS 0.039761f
C8278 PAD.n9197 VSS 0.023109f
C8279 PAD.n9198 VSS 0.03338f
C8280 PAD.n9199 VSS 0.036461f
C8281 PAD.n9200 VSS 0.036461f
C8282 PAD.n9201 VSS 0.036461f
C8283 PAD.n9202 VSS 0.036461f
C8284 PAD.n9204 VSS 0.036461f
C8285 PAD.n9205 VSS 0.036461f
C8286 PAD.n9206 VSS 0.036461f
C8287 PAD.n9208 VSS 0.036461f
C8288 PAD.n9209 VSS 0.036461f
C8289 PAD.n9210 VSS 0.036461f
C8290 PAD.n9211 VSS 0.036461f
C8291 PAD.n9212 VSS 0.036461f
C8292 PAD.n9213 VSS 0.036461f
C8293 PAD.n9214 VSS 0.036461f
C8294 PAD.n9216 VSS 0.036461f
C8295 PAD.n9217 VSS 0.036461f
C8296 PAD.n9218 VSS 0.036461f
C8297 PAD.n9220 VSS 0.036461f
C8298 PAD.n9221 VSS 0.036461f
C8299 PAD.n9222 VSS 0.036461f
C8300 PAD.n9223 VSS 0.036461f
C8301 PAD.n9224 VSS 0.036461f
C8302 PAD.n9225 VSS 0.036461f
C8303 PAD.n9226 VSS 0.036461f
C8304 PAD.n9228 VSS 0.036461f
C8305 PAD.n9229 VSS 0.036461f
C8306 PAD.n9230 VSS 0.036461f
C8307 PAD.n9232 VSS 0.036461f
C8308 PAD.n9233 VSS 0.036461f
C8309 PAD.n9234 VSS 0.036461f
C8310 PAD.n9235 VSS 0.036461f
C8311 PAD.n9236 VSS 0.036461f
C8312 PAD.n9237 VSS 0.036461f
C8313 PAD.n9238 VSS 0.036461f
C8314 PAD.n9240 VSS 0.036461f
C8315 PAD.n9241 VSS 0.036461f
C8316 PAD.n9242 VSS 0.036461f
C8317 PAD.n9244 VSS 0.036461f
C8318 PAD.n9245 VSS 0.036461f
C8319 PAD.n9246 VSS 0.036461f
C8320 PAD.n9247 VSS 0.036461f
C8321 PAD.n9248 VSS 0.036461f
C8322 PAD.n9249 VSS 0.036461f
C8323 PAD.n9250 VSS 0.036461f
C8324 PAD.n9252 VSS 0.036461f
C8325 PAD.n9253 VSS 0.036461f
C8326 PAD.n9254 VSS 0.036461f
C8327 PAD.n9256 VSS 0.036461f
C8328 PAD.n9257 VSS 0.036461f
C8329 PAD.n9258 VSS 0.036461f
C8330 PAD.n9259 VSS 0.036461f
C8331 PAD.n9260 VSS 0.036461f
C8332 PAD.n9261 VSS 0.036461f
C8333 PAD.n9262 VSS 0.036461f
C8334 PAD.n9264 VSS 0.036461f
C8335 PAD.n9265 VSS 0.036461f
C8336 PAD.n9266 VSS 0.036461f
C8337 PAD.n9268 VSS 0.036461f
C8338 PAD.n9269 VSS 0.036461f
C8339 PAD.n9270 VSS 0.036461f
C8340 PAD.n9271 VSS 0.036461f
C8341 PAD.n9272 VSS 0.036461f
C8342 PAD.n9273 VSS 0.036461f
C8343 PAD.n9274 VSS 0.036461f
C8344 PAD.n9276 VSS 0.036461f
C8345 PAD.n9277 VSS 0.036461f
C8346 PAD.n9278 VSS 0.036461f
C8347 PAD.n9280 VSS 0.036461f
C8348 PAD.n9281 VSS 0.036461f
C8349 PAD.n9282 VSS 0.036461f
C8350 PAD.n9283 VSS 0.036461f
C8351 PAD.n9284 VSS 0.036461f
C8352 PAD.n9285 VSS 0.036461f
C8353 PAD.n9286 VSS 0.036461f
C8354 PAD.n9288 VSS 0.036461f
C8355 PAD.n9289 VSS 0.036461f
C8356 PAD.n9290 VSS 0.036461f
C8357 PAD.n9292 VSS 0.036461f
C8358 PAD.n9293 VSS 0.036461f
C8359 PAD.n9294 VSS 0.036461f
C8360 PAD.n9295 VSS 0.036461f
C8361 PAD.n9296 VSS 0.036461f
C8362 PAD.n9297 VSS 0.036461f
C8363 PAD.n9298 VSS 0.036461f
C8364 PAD.n9300 VSS 0.036461f
C8365 PAD.n9301 VSS 0.036461f
C8366 PAD.n9302 VSS 0.036461f
C8367 PAD.n9304 VSS 0.036461f
C8368 PAD.n9305 VSS 0.036461f
C8369 PAD.n9306 VSS 0.036461f
C8370 PAD.n9307 VSS 0.036461f
C8371 PAD.n9308 VSS 0.036461f
C8372 PAD.n9309 VSS 0.036461f
C8373 PAD.n9310 VSS 0.036461f
C8374 PAD.n9312 VSS 0.036461f
C8375 PAD.n9313 VSS 0.036461f
C8376 PAD.n9314 VSS 0.036461f
C8377 PAD.n9316 VSS 0.036461f
C8378 PAD.n9317 VSS 0.036461f
C8379 PAD.n9318 VSS 0.036461f
C8380 PAD.n9319 VSS 0.036461f
C8381 PAD.n9320 VSS 0.036461f
C8382 PAD.n9321 VSS 0.036461f
C8383 PAD.n9322 VSS 0.036461f
C8384 PAD.n9324 VSS 0.036461f
C8385 PAD.n9325 VSS 0.036461f
C8386 PAD.n9326 VSS 0.036461f
C8387 PAD.n9328 VSS 0.036461f
C8388 PAD.n9329 VSS 0.036461f
C8389 PAD.n9330 VSS 0.036461f
C8390 PAD.n9331 VSS 0.036461f
C8391 PAD.n9332 VSS 0.036461f
C8392 PAD.n9333 VSS 0.036461f
C8393 PAD.n9334 VSS 0.036461f
C8394 PAD.n9336 VSS 0.036461f
C8395 PAD.n9337 VSS 0.036461f
C8396 PAD.n9338 VSS 0.036461f
C8397 PAD.n9340 VSS 0.036461f
C8398 PAD.n9341 VSS 0.036461f
C8399 PAD.n9342 VSS 0.036461f
C8400 PAD.n9343 VSS 0.036461f
C8401 PAD.n9344 VSS 0.036461f
C8402 PAD.n9345 VSS 0.036461f
C8403 PAD.n9346 VSS 0.036461f
C8404 PAD.n9348 VSS 0.036461f
C8405 PAD.n9349 VSS 0.036461f
C8406 PAD.n9350 VSS 0.036461f
C8407 PAD.n9352 VSS 0.036461f
C8408 PAD.n9353 VSS 0.036461f
C8409 PAD.n9354 VSS 0.036461f
C8410 PAD.n9355 VSS 0.036461f
C8411 PAD.n9356 VSS 0.036461f
C8412 PAD.n9357 VSS 0.036461f
C8413 PAD.n9358 VSS 0.036461f
C8414 PAD.n9360 VSS 0.036461f
C8415 PAD.n9361 VSS 0.036461f
C8416 PAD.n9362 VSS 0.036461f
C8417 PAD.n9364 VSS 0.036461f
C8418 PAD.n9365 VSS 0.036461f
C8419 PAD.n9366 VSS 0.036461f
C8420 PAD.n9367 VSS 0.036461f
C8421 PAD.n9368 VSS 0.036461f
C8422 PAD.n9369 VSS 0.036461f
C8423 PAD.n9370 VSS 0.036461f
C8424 PAD.n9372 VSS 0.036461f
C8425 PAD.n9373 VSS 0.036461f
C8426 PAD.n9374 VSS 0.036461f
C8427 PAD.n9376 VSS 0.036461f
C8428 PAD.n9377 VSS 0.036461f
C8429 PAD.n9378 VSS 0.036461f
C8430 PAD.n9379 VSS 0.036461f
C8431 PAD.n9380 VSS 0.036461f
C8432 PAD.n9381 VSS 0.036461f
C8433 PAD.n9382 VSS 0.036461f
C8434 PAD.n9384 VSS 0.036461f
C8435 PAD.n9385 VSS 0.036461f
C8436 PAD.n9386 VSS 0.036461f
C8437 PAD.n9388 VSS 0.036461f
C8438 PAD.n9389 VSS 0.036461f
C8439 PAD.n9390 VSS 0.036461f
C8440 PAD.n9391 VSS 0.036461f
C8441 PAD.n9392 VSS 0.036461f
C8442 PAD.n9393 VSS 0.036461f
C8443 PAD.n9394 VSS 0.036461f
C8444 PAD.n9396 VSS 0.036461f
C8445 PAD.n9397 VSS 0.036461f
C8446 PAD.n9398 VSS 0.036461f
C8447 PAD.n9400 VSS 0.036461f
C8448 PAD.n9401 VSS 0.036461f
C8449 PAD.n9402 VSS 0.036461f
C8450 PAD.n9403 VSS 0.036461f
C8451 PAD.n9404 VSS 0.036461f
C8452 PAD.n9405 VSS 0.036461f
C8453 PAD.n9406 VSS 0.036461f
C8454 PAD.n9408 VSS 0.036461f
C8455 PAD.n9409 VSS 0.036461f
C8456 PAD.n9410 VSS 0.036461f
C8457 PAD.n9412 VSS 0.036461f
C8458 PAD.n9413 VSS 0.036461f
C8459 PAD.n9414 VSS 0.036461f
C8460 PAD.n9415 VSS 0.036461f
C8461 PAD.n9416 VSS 0.036461f
C8462 PAD.n9417 VSS 0.036461f
C8463 PAD.n9418 VSS 0.036461f
C8464 PAD.n9420 VSS 0.036461f
C8465 PAD.n9421 VSS 0.036461f
C8466 PAD.n9422 VSS 0.036461f
C8467 PAD.n9424 VSS 0.036461f
C8468 PAD.n9425 VSS 0.036461f
C8469 PAD.n9426 VSS 0.036461f
C8470 PAD.n9427 VSS 0.036461f
C8471 PAD.n9428 VSS 0.036461f
C8472 PAD.n9429 VSS 0.036461f
C8473 PAD.n9430 VSS 0.036461f
C8474 PAD.n9432 VSS 0.036461f
C8475 PAD.n9433 VSS 0.036461f
C8476 PAD.n9434 VSS 0.036461f
C8477 PAD.n9436 VSS 0.036461f
C8478 PAD.n9437 VSS 0.036461f
C8479 PAD.n9438 VSS 0.036461f
C8480 PAD.n9439 VSS 0.036461f
C8481 PAD.n9440 VSS 0.036461f
C8482 PAD.n9441 VSS 0.036461f
C8483 PAD.n9442 VSS 0.036461f
C8484 PAD.n9444 VSS 0.023109f
C8485 PAD.n9445 VSS 0.547601f
C8486 PAD.n9446 VSS 0.453867f
C8487 PAD.n9447 VSS 0.025768f
C8488 PAD.n9448 VSS 0.025768f
C8489 PAD.n9449 VSS 0.022505f
C8490 PAD.n9450 VSS 0.033773f
C8491 PAD.n9451 VSS 0.041838f
C8492 PAD.n9452 VSS 0.040026f
C8493 PAD.n9453 VSS 0.045829f
C8494 PAD.n9454 VSS 0.045829f
C8495 PAD.n9455 VSS 0.5032f
C8496 PAD.n9456 VSS 0.700534f
C8497 PAD.n9457 VSS 0.069765f
C8498 PAD.n9458 VSS 0.048386f
C8499 PAD.n9459 VSS 0.039761f
C8500 PAD.n9460 VSS 0.056262f
C8501 PAD.n9461 VSS 0.056262f
C8502 PAD.n9462 VSS 0.039761f
C8503 PAD.n9463 VSS 0.023109f
C8504 PAD.n9464 VSS 0.03338f
C8505 PAD.n9465 VSS 0.036461f
C8506 PAD.n9466 VSS 0.036461f
C8507 PAD.n9467 VSS 0.036461f
C8508 PAD.n9468 VSS 0.036461f
C8509 PAD.n9470 VSS 0.036461f
C8510 PAD.n9471 VSS 0.036461f
C8511 PAD.n9472 VSS 0.036461f
C8512 PAD.n9474 VSS 0.036461f
C8513 PAD.n9475 VSS 0.036461f
C8514 PAD.n9476 VSS 0.036461f
C8515 PAD.n9477 VSS 0.036461f
C8516 PAD.n9478 VSS 0.036461f
C8517 PAD.n9479 VSS 0.036461f
C8518 PAD.n9480 VSS 0.036461f
C8519 PAD.n9482 VSS 0.036461f
C8520 PAD.n9483 VSS 0.036461f
C8521 PAD.n9484 VSS 0.036461f
C8522 PAD.n9486 VSS 0.036461f
C8523 PAD.n9487 VSS 0.036461f
C8524 PAD.n9488 VSS 0.036461f
C8525 PAD.n9489 VSS 0.036461f
C8526 PAD.n9490 VSS 0.036461f
C8527 PAD.n9491 VSS 0.036461f
C8528 PAD.n9492 VSS 0.036461f
C8529 PAD.n9494 VSS 0.036461f
C8530 PAD.n9495 VSS 0.036461f
C8531 PAD.n9496 VSS 0.036461f
C8532 PAD.n9498 VSS 0.036461f
C8533 PAD.n9499 VSS 0.036461f
C8534 PAD.n9500 VSS 0.036461f
C8535 PAD.n9501 VSS 0.036461f
C8536 PAD.n9502 VSS 0.036461f
C8537 PAD.n9503 VSS 0.036461f
C8538 PAD.n9504 VSS 0.036461f
C8539 PAD.n9506 VSS 0.036461f
C8540 PAD.n9507 VSS 0.036461f
C8541 PAD.n9508 VSS 0.036461f
C8542 PAD.n9510 VSS 0.036461f
C8543 PAD.n9511 VSS 0.036461f
C8544 PAD.n9512 VSS 0.036461f
C8545 PAD.n9513 VSS 0.036461f
C8546 PAD.n9514 VSS 0.036461f
C8547 PAD.n9515 VSS 0.036461f
C8548 PAD.n9516 VSS 0.036461f
C8549 PAD.n9518 VSS 0.036461f
C8550 PAD.n9519 VSS 0.036461f
C8551 PAD.n9520 VSS 0.036461f
C8552 PAD.n9522 VSS 0.036461f
C8553 PAD.n9523 VSS 0.036461f
C8554 PAD.n9524 VSS 0.036461f
C8555 PAD.n9525 VSS 0.036461f
C8556 PAD.n9526 VSS 0.036461f
C8557 PAD.n9527 VSS 0.036461f
C8558 PAD.n9528 VSS 0.036461f
C8559 PAD.n9530 VSS 0.036461f
C8560 PAD.n9531 VSS 0.036461f
C8561 PAD.n9532 VSS 0.036461f
C8562 PAD.n9534 VSS 0.036461f
C8563 PAD.n9535 VSS 0.036461f
C8564 PAD.n9536 VSS 0.036461f
C8565 PAD.n9537 VSS 0.036461f
C8566 PAD.n9538 VSS 0.036461f
C8567 PAD.n9539 VSS 0.036461f
C8568 PAD.n9540 VSS 0.036461f
C8569 PAD.n9542 VSS 0.036461f
C8570 PAD.n9543 VSS 0.036461f
C8571 PAD.n9544 VSS 0.036461f
C8572 PAD.n9546 VSS 0.036461f
C8573 PAD.n9547 VSS 0.036461f
C8574 PAD.n9548 VSS 0.036461f
C8575 PAD.n9549 VSS 0.036461f
C8576 PAD.n9550 VSS 0.036461f
C8577 PAD.n9551 VSS 0.036461f
C8578 PAD.n9552 VSS 0.036461f
C8579 PAD.n9554 VSS 0.036461f
C8580 PAD.n9555 VSS 0.036461f
C8581 PAD.n9556 VSS 0.036461f
C8582 PAD.n9558 VSS 0.036461f
C8583 PAD.n9559 VSS 0.036461f
C8584 PAD.n9560 VSS 0.036461f
C8585 PAD.n9561 VSS 0.036461f
C8586 PAD.n9562 VSS 0.036461f
C8587 PAD.n9563 VSS 0.036461f
C8588 PAD.n9564 VSS 0.036461f
C8589 PAD.n9566 VSS 0.036461f
C8590 PAD.n9567 VSS 0.036461f
C8591 PAD.n9568 VSS 0.036461f
C8592 PAD.n9570 VSS 0.036461f
C8593 PAD.n9571 VSS 0.036461f
C8594 PAD.n9572 VSS 0.036461f
C8595 PAD.n9573 VSS 0.036461f
C8596 PAD.n9574 VSS 0.036461f
C8597 PAD.n9575 VSS 0.036461f
C8598 PAD.n9576 VSS 0.036461f
C8599 PAD.n9578 VSS 0.036461f
C8600 PAD.n9579 VSS 0.036461f
C8601 PAD.n9580 VSS 0.036461f
C8602 PAD.n9582 VSS 0.036461f
C8603 PAD.n9583 VSS 0.036461f
C8604 PAD.n9584 VSS 0.036461f
C8605 PAD.n9585 VSS 0.036461f
C8606 PAD.n9586 VSS 0.036461f
C8607 PAD.n9587 VSS 0.036461f
C8608 PAD.n9588 VSS 0.036461f
C8609 PAD.n9590 VSS 0.036461f
C8610 PAD.n9591 VSS 0.036461f
C8611 PAD.n9592 VSS 0.036461f
C8612 PAD.n9594 VSS 0.036461f
C8613 PAD.n9595 VSS 0.036461f
C8614 PAD.n9596 VSS 0.036461f
C8615 PAD.n9597 VSS 0.036461f
C8616 PAD.n9598 VSS 0.036461f
C8617 PAD.n9599 VSS 0.036461f
C8618 PAD.n9600 VSS 0.036461f
C8619 PAD.n9602 VSS 0.036461f
C8620 PAD.n9603 VSS 0.036461f
C8621 PAD.n9604 VSS 0.036461f
C8622 PAD.n9606 VSS 0.036461f
C8623 PAD.n9607 VSS 0.036461f
C8624 PAD.n9608 VSS 0.036461f
C8625 PAD.n9609 VSS 0.036461f
C8626 PAD.n9610 VSS 0.036461f
C8627 PAD.n9611 VSS 0.036461f
C8628 PAD.n9612 VSS 0.036461f
C8629 PAD.n9614 VSS 0.036461f
C8630 PAD.n9615 VSS 0.036461f
C8631 PAD.n9616 VSS 0.036461f
C8632 PAD.n9618 VSS 0.036461f
C8633 PAD.n9619 VSS 0.036461f
C8634 PAD.n9620 VSS 0.036461f
C8635 PAD.n9621 VSS 0.036461f
C8636 PAD.n9622 VSS 0.036461f
C8637 PAD.n9623 VSS 0.036461f
C8638 PAD.n9624 VSS 0.036461f
C8639 PAD.n9626 VSS 0.036461f
C8640 PAD.n9627 VSS 0.036461f
C8641 PAD.n9628 VSS 0.036461f
C8642 PAD.n9630 VSS 0.036461f
C8643 PAD.n9631 VSS 0.036461f
C8644 PAD.n9632 VSS 0.036461f
C8645 PAD.n9633 VSS 0.036461f
C8646 PAD.n9634 VSS 0.036461f
C8647 PAD.n9635 VSS 0.036461f
C8648 PAD.n9636 VSS 0.036461f
C8649 PAD.n9638 VSS 0.036461f
C8650 PAD.n9639 VSS 0.036461f
C8651 PAD.n9640 VSS 0.036461f
C8652 PAD.n9642 VSS 0.036461f
C8653 PAD.n9643 VSS 0.036461f
C8654 PAD.n9644 VSS 0.036461f
C8655 PAD.n9645 VSS 0.036461f
C8656 PAD.n9646 VSS 0.036461f
C8657 PAD.n9647 VSS 0.036461f
C8658 PAD.n9648 VSS 0.036461f
C8659 PAD.n9650 VSS 0.036461f
C8660 PAD.n9651 VSS 0.036461f
C8661 PAD.n9652 VSS 0.036461f
C8662 PAD.n9654 VSS 0.036461f
C8663 PAD.n9655 VSS 0.036461f
C8664 PAD.n9656 VSS 0.036461f
C8665 PAD.n9657 VSS 0.036461f
C8666 PAD.n9658 VSS 0.036461f
C8667 PAD.n9659 VSS 0.036461f
C8668 PAD.n9660 VSS 0.036461f
C8669 PAD.n9662 VSS 0.036461f
C8670 PAD.n9663 VSS 0.036461f
C8671 PAD.n9664 VSS 0.036461f
C8672 PAD.n9666 VSS 0.036461f
C8673 PAD.n9667 VSS 0.036461f
C8674 PAD.n9668 VSS 0.036461f
C8675 PAD.n9669 VSS 0.036461f
C8676 PAD.n9670 VSS 0.036461f
C8677 PAD.n9671 VSS 0.036461f
C8678 PAD.n9672 VSS 0.036461f
C8679 PAD.n9674 VSS 0.036461f
C8680 PAD.n9675 VSS 0.036461f
C8681 PAD.n9676 VSS 0.036461f
C8682 PAD.n9678 VSS 0.036461f
C8683 PAD.n9679 VSS 0.036461f
C8684 PAD.n9680 VSS 0.036461f
C8685 PAD.n9681 VSS 0.036461f
C8686 PAD.n9682 VSS 0.036461f
C8687 PAD.n9683 VSS 0.036461f
C8688 PAD.n9684 VSS 0.036461f
C8689 PAD.n9686 VSS 0.036461f
C8690 PAD.n9687 VSS 0.036461f
C8691 PAD.n9688 VSS 0.036461f
C8692 PAD.n9690 VSS 0.036461f
C8693 PAD.n9691 VSS 0.036461f
C8694 PAD.n9692 VSS 0.036461f
C8695 PAD.n9693 VSS 0.036461f
C8696 PAD.n9694 VSS 0.036461f
C8697 PAD.n9695 VSS 0.036461f
C8698 PAD.n9696 VSS 0.036461f
C8699 PAD.n9698 VSS 0.036461f
C8700 PAD.n9699 VSS 0.036461f
C8701 PAD.n9700 VSS 0.036461f
C8702 PAD.n9702 VSS 0.036461f
C8703 PAD.n9703 VSS 0.036461f
C8704 PAD.n9704 VSS 0.036461f
C8705 PAD.n9705 VSS 0.036461f
C8706 PAD.n9706 VSS 0.030555f
C8707 PAD.n9707 VSS 0.036461f
C8708 PAD.n9708 VSS 0.036461f
C8709 PAD.n9709 VSS 0.036461f
C8710 PAD.n9711 VSS 0.023109f
C8711 PAD.n9712 VSS 0.2812f
C8712 PAD.n9713 VSS 0.592001f
C8713 PAD.n9714 VSS 0.027844f
C8714 PAD.n9715 VSS 0.027844f
C8715 PAD.n9716 VSS 0.024317f
C8716 PAD.n9717 VSS 0.042895f
C8717 PAD.n9718 VSS 0.036099f
C8718 PAD.n9719 VSS 0.041333f
C8719 PAD.n9720 VSS 0.041333f
C8720 PAD.n9721 VSS 0.611734f
C8721 PAD.n9722 VSS 0.157866f
C8722 PAD.n9723 VSS 0.056262f
C8723 PAD.n9724 VSS 0.056262f
C8724 PAD.n9725 VSS 0.050221f
C8725 PAD.n9726 VSS 0.046286f
C8726 PAD.n9727 VSS 0.057252f
C8727 PAD.n9728 VSS 0.062274f
C8728 PAD.n9729 VSS 0.04319f
C8729 PAD.n9730 VSS 0.048386f
C8730 PAD.n9731 VSS 0.048386f
C8731 PAD.n9732 VSS 0.157866f
C8732 PAD.n9733 VSS 0.557468f
C8733 PAD.n9734 VSS 0.03234f
C8734 PAD.n9735 VSS 0.03234f
C8735 PAD.n9736 VSS 0.028244f
C8736 PAD.n9737 VSS 0.042895f
C8737 PAD.n9738 VSS 0.032172f
C8738 PAD.n9739 VSS 0.036836f
C8739 PAD.n9740 VSS 0.036836f
C8740 PAD.n9741 VSS 0.1776f
C8741 PAD.n9742 VSS 0.700534f
C8742 PAD.n9743 VSS 0.064139f
C8743 PAD.n9744 VSS 0.039761f
C8744 PAD.n9745 VSS 0.069765f
C8745 PAD.n9746 VSS 0.040509f
C8746 PAD.n9747 VSS 0.040509f
C8747 PAD.n9748 VSS 0.039761f
C8748 PAD.n9749 VSS 0.023109f
C8749 PAD.n9750 VSS 0.03338f
C8750 PAD.n9751 VSS 0.036461f
C8751 PAD.n9752 VSS 0.036461f
C8752 PAD.n9753 VSS 0.036461f
C8753 PAD.n9754 VSS 0.036461f
C8754 PAD.n9756 VSS 0.036461f
C8755 PAD.n9757 VSS 0.036461f
C8756 PAD.n9758 VSS 0.036461f
C8757 PAD.n9760 VSS 0.036461f
C8758 PAD.n9761 VSS 0.036461f
C8759 PAD.n9762 VSS 0.036461f
C8760 PAD.n9763 VSS 0.036461f
C8761 PAD.n9764 VSS 0.036461f
C8762 PAD.n9765 VSS 0.036461f
C8763 PAD.n9766 VSS 0.036461f
C8764 PAD.n9768 VSS 0.036461f
C8765 PAD.n9769 VSS 0.036461f
C8766 PAD.n9770 VSS 0.036461f
C8767 PAD.n9772 VSS 0.036461f
C8768 PAD.n9773 VSS 0.036461f
C8769 PAD.n9774 VSS 0.036461f
C8770 PAD.n9775 VSS 0.036461f
C8771 PAD.n9776 VSS 0.036461f
C8772 PAD.n9777 VSS 0.036461f
C8773 PAD.n9778 VSS 0.036461f
C8774 PAD.n9780 VSS 0.036461f
C8775 PAD.n9781 VSS 0.036461f
C8776 PAD.n9782 VSS 0.036461f
C8777 PAD.n9784 VSS 0.036461f
C8778 PAD.n9785 VSS 0.036461f
C8779 PAD.n9786 VSS 0.036461f
C8780 PAD.n9787 VSS 0.036461f
C8781 PAD.n9788 VSS 0.036461f
C8782 PAD.n9789 VSS 0.036461f
C8783 PAD.n9790 VSS 0.036461f
C8784 PAD.n9792 VSS 0.036461f
C8785 PAD.n9793 VSS 0.036461f
C8786 PAD.n9794 VSS 0.036461f
C8787 PAD.n9796 VSS 0.036461f
C8788 PAD.n9797 VSS 0.036461f
C8789 PAD.n9798 VSS 0.036461f
C8790 PAD.n9799 VSS 0.036461f
C8791 PAD.n9800 VSS 0.036461f
C8792 PAD.n9801 VSS 0.036461f
C8793 PAD.n9802 VSS 0.036461f
C8794 PAD.n9804 VSS 0.036461f
C8795 PAD.n9805 VSS 0.036461f
C8796 PAD.n9806 VSS 0.036461f
C8797 PAD.n9808 VSS 0.036461f
C8798 PAD.n9809 VSS 0.036461f
C8799 PAD.n9810 VSS 0.036461f
C8800 PAD.n9811 VSS 0.036461f
C8801 PAD.n9812 VSS 0.036461f
C8802 PAD.n9813 VSS 0.036461f
C8803 PAD.n9814 VSS 0.036461f
C8804 PAD.n9816 VSS 0.036461f
C8805 PAD.n9817 VSS 0.036461f
C8806 PAD.n9818 VSS 0.036461f
C8807 PAD.n9820 VSS 0.036461f
C8808 PAD.n9821 VSS 0.036461f
C8809 PAD.n9822 VSS 0.036461f
C8810 PAD.n9823 VSS 0.036461f
C8811 PAD.n9824 VSS 0.036461f
C8812 PAD.n9825 VSS 0.036461f
C8813 PAD.n9826 VSS 0.036461f
C8814 PAD.n9828 VSS 0.036461f
C8815 PAD.n9829 VSS 0.036461f
C8816 PAD.n9830 VSS 0.036461f
C8817 PAD.n9832 VSS 0.036461f
C8818 PAD.n9833 VSS 0.036461f
C8819 PAD.n9834 VSS 0.036461f
C8820 PAD.n9835 VSS 0.036461f
C8821 PAD.n9836 VSS 0.036461f
C8822 PAD.n9837 VSS 0.036461f
C8823 PAD.n9838 VSS 0.036461f
C8824 PAD.n9840 VSS 0.036461f
C8825 PAD.n9841 VSS 0.036461f
C8826 PAD.n9842 VSS 0.036461f
C8827 PAD.n9844 VSS 0.036461f
C8828 PAD.n9845 VSS 0.036461f
C8829 PAD.n9846 VSS 0.036461f
C8830 PAD.n9847 VSS 0.036461f
C8831 PAD.n9848 VSS 0.036461f
C8832 PAD.n9849 VSS 0.036461f
C8833 PAD.n9850 VSS 0.036461f
C8834 PAD.n9852 VSS 0.036461f
C8835 PAD.n9853 VSS 0.036461f
C8836 PAD.n9854 VSS 0.036461f
C8837 PAD.n9856 VSS 0.036461f
C8838 PAD.n9857 VSS 0.036461f
C8839 PAD.n9858 VSS 0.036461f
C8840 PAD.n9859 VSS 0.036461f
C8841 PAD.n9860 VSS 0.036461f
C8842 PAD.n9861 VSS 0.036461f
C8843 PAD.n9862 VSS 0.036461f
C8844 PAD.n9864 VSS 0.036461f
C8845 PAD.n9865 VSS 0.036461f
C8846 PAD.n9866 VSS 0.036461f
C8847 PAD.n9868 VSS 0.036461f
C8848 PAD.n9869 VSS 0.036461f
C8849 PAD.n9870 VSS 0.036461f
C8850 PAD.n9871 VSS 0.036461f
C8851 PAD.n9872 VSS 0.036461f
C8852 PAD.n9873 VSS 0.036461f
C8853 PAD.n9874 VSS 0.036461f
C8854 PAD.n9876 VSS 0.036461f
C8855 PAD.n9877 VSS 0.036461f
C8856 PAD.n9878 VSS 0.036461f
C8857 PAD.n9880 VSS 0.036461f
C8858 PAD.n9881 VSS 0.036461f
C8859 PAD.n9882 VSS 0.036461f
C8860 PAD.n9883 VSS 0.036461f
C8861 PAD.n9884 VSS 0.036461f
C8862 PAD.n9885 VSS 0.036461f
C8863 PAD.n9886 VSS 0.036461f
C8864 PAD.n9888 VSS 0.036461f
C8865 PAD.n9889 VSS 0.036461f
C8866 PAD.n9890 VSS 0.036461f
C8867 PAD.n9892 VSS 0.036461f
C8868 PAD.n9893 VSS 0.036461f
C8869 PAD.n9894 VSS 0.036461f
C8870 PAD.n9895 VSS 0.036461f
C8871 PAD.n9896 VSS 0.036461f
C8872 PAD.n9897 VSS 0.036461f
C8873 PAD.n9898 VSS 0.036461f
C8874 PAD.n9900 VSS 0.036461f
C8875 PAD.n9901 VSS 0.036461f
C8876 PAD.n9902 VSS 0.036461f
C8877 PAD.n9904 VSS 0.036461f
C8878 PAD.n9905 VSS 0.036461f
C8879 PAD.n9906 VSS 0.036461f
C8880 PAD.n9907 VSS 0.036461f
C8881 PAD.n9908 VSS 0.036461f
C8882 PAD.n9909 VSS 0.036461f
C8883 PAD.n9910 VSS 0.036461f
C8884 PAD.n9912 VSS 0.036461f
C8885 PAD.n9913 VSS 0.036461f
C8886 PAD.n9914 VSS 0.036461f
C8887 PAD.n9916 VSS 0.036461f
C8888 PAD.n9917 VSS 0.036461f
C8889 PAD.n9918 VSS 0.036461f
C8890 PAD.n9919 VSS 0.036461f
C8891 PAD.n9920 VSS 0.036461f
C8892 PAD.n9921 VSS 0.036461f
C8893 PAD.n9922 VSS 0.036461f
C8894 PAD.n9924 VSS 0.036461f
C8895 PAD.n9925 VSS 0.036461f
C8896 PAD.n9926 VSS 0.036461f
C8897 PAD.n9928 VSS 0.036461f
C8898 PAD.n9929 VSS 0.036461f
C8899 PAD.n9930 VSS 0.036461f
C8900 PAD.n9931 VSS 0.036461f
C8901 PAD.n9932 VSS 0.036461f
C8902 PAD.n9933 VSS 0.036461f
C8903 PAD.n9934 VSS 0.036461f
C8904 PAD.n9936 VSS 0.036461f
C8905 PAD.n9937 VSS 0.036461f
C8906 PAD.n9938 VSS 0.036461f
C8907 PAD.n9940 VSS 0.036461f
C8908 PAD.n9941 VSS 0.036461f
C8909 PAD.n9942 VSS 0.036461f
C8910 PAD.n9943 VSS 0.036461f
C8911 PAD.n9944 VSS 0.036461f
C8912 PAD.n9945 VSS 0.036461f
C8913 PAD.n9946 VSS 0.036461f
C8914 PAD.n9948 VSS 0.036461f
C8915 PAD.n9949 VSS 0.036461f
C8916 PAD.n9950 VSS 0.036461f
C8917 PAD.n9952 VSS 0.036461f
C8918 PAD.n9953 VSS 0.036461f
C8919 PAD.n9954 VSS 0.036461f
C8920 PAD.n9955 VSS 0.036461f
C8921 PAD.n9956 VSS 0.036461f
C8922 PAD.n9957 VSS 0.036461f
C8923 PAD.n9958 VSS 0.036461f
C8924 PAD.n9960 VSS 0.036461f
C8925 PAD.n9961 VSS 0.036461f
C8926 PAD.n9962 VSS 0.036461f
C8927 PAD.n9964 VSS 0.036461f
C8928 PAD.n9965 VSS 0.036461f
C8929 PAD.n9966 VSS 0.036461f
C8930 PAD.n9967 VSS 0.036461f
C8931 PAD.n9968 VSS 0.036461f
C8932 PAD.n9969 VSS 0.036461f
C8933 PAD.n9970 VSS 0.036461f
C8934 PAD.n9972 VSS 0.036461f
C8935 PAD.n9973 VSS 0.036461f
C8936 PAD.n9974 VSS 0.036461f
C8937 PAD.n9976 VSS 0.036461f
C8938 PAD.n9977 VSS 0.036461f
C8939 PAD.n9978 VSS 0.036461f
C8940 PAD.n9979 VSS 0.036461f
C8941 PAD.n9980 VSS 0.036461f
C8942 PAD.n9981 VSS 0.036461f
C8943 PAD.n9982 VSS 0.036461f
C8944 PAD.n9984 VSS 0.036461f
C8945 PAD.n9985 VSS 0.036461f
C8946 PAD.n9986 VSS 0.036461f
C8947 PAD.n9988 VSS 0.036461f
C8948 PAD.n9989 VSS 0.036461f
C8949 PAD.n9990 VSS 0.036461f
C8950 PAD.n9991 VSS 0.036461f
C8951 PAD.n9992 VSS 0.030555f
C8952 PAD.n9993 VSS 0.036461f
C8953 PAD.n9994 VSS 0.036461f
C8954 PAD.n9995 VSS 0.036461f
C8955 PAD.n9997 VSS 0.023109f
C8956 PAD.n9998 VSS 0.360134f
C8957 PAD.n9999 VSS 0.2664f
C8958 PAD.n10000 VSS 0.036836f
C8959 PAD.n10001 VSS 0.036836f
C8960 PAD.n10002 VSS 0.032172f
C8961 PAD.n10003 VSS 0.042895f
C8962 PAD.n10004 VSS 0.028244f
C8963 PAD.n10005 VSS 0.03234f
C8964 PAD.n10006 VSS 0.03234f
C8965 PAD.n10007 VSS 0.296f
C8966 PAD.n10008 VSS 0.587068f
C8967 PAD.n10009 VSS 0.037133f
C8968 PAD.n10010 VSS 0.037133f
C8969 PAD.n10011 VSS 0.033146f
C8970 PAD.n10012 VSS 0.046286f
C8971 PAD.n10013 VSS 0.060265f
C8972 PAD.n10014 VSS 0.067515f
C8973 PAD.n10015 VSS 0.067515f
C8974 PAD.n10016 VSS 0.700534f
C8975 PAD.n10017 VSS 0.2072f
C8976 PAD.n10018 VSS 0.041333f
C8977 PAD.n10019 VSS 0.041333f
C8978 PAD.n10020 VSS 0.036099f
C8979 PAD.n10021 VSS 0.042895f
C8980 PAD.n10022 VSS 0.036461f
C8981 PAD.n10023 VSS 0.036461f
C8982 PAD.n10024 VSS 0.036461f
C8983 PAD.n10026 VSS 0.036461f
C8984 PAD.n10027 VSS 0.036461f
C8985 PAD.n10028 VSS 0.036461f
C8986 PAD.n10030 VSS 0.036461f
C8987 PAD.n10031 VSS 0.036461f
C8988 PAD.n10032 VSS 0.036461f
C8989 PAD.n10034 VSS 0.036461f
C8990 PAD.n10035 VSS 0.036461f
C8991 PAD.n10036 VSS 0.036461f
C8992 PAD.n10038 VSS 0.036461f
C8993 PAD.n10039 VSS 0.036461f
C8994 PAD.n10040 VSS 0.036461f
C8995 PAD.n10042 VSS 0.036461f
C8996 PAD.n10043 VSS 0.036461f
C8997 PAD.n10044 VSS 0.036461f
C8998 PAD.n10046 VSS 0.036461f
C8999 PAD.n10047 VSS 0.036461f
C9000 PAD.n10048 VSS 0.036461f
C9001 PAD.n10050 VSS 0.036461f
C9002 PAD.n10051 VSS 0.036461f
C9003 PAD.n10052 VSS 0.036461f
C9004 PAD.n10054 VSS 0.036461f
C9005 PAD.n10055 VSS 0.036461f
C9006 PAD.n10056 VSS 0.036461f
C9007 PAD.n10058 VSS 0.036461f
C9008 PAD.n10059 VSS 0.036461f
C9009 PAD.n10060 VSS 0.036461f
C9010 PAD.n10062 VSS 0.036461f
C9011 PAD.n10063 VSS 0.036461f
C9012 PAD.n10064 VSS 0.036461f
C9013 PAD.n10066 VSS 0.036461f
C9014 PAD.n10067 VSS 0.036461f
C9015 PAD.n10068 VSS 0.036461f
C9016 PAD.n10070 VSS 0.036461f
C9017 PAD.n10071 VSS 0.036461f
C9018 PAD.n10072 VSS 0.036461f
C9019 PAD.n10074 VSS 0.036461f
C9020 PAD.n10075 VSS 0.036461f
C9021 PAD.n10076 VSS 0.036461f
C9022 PAD.n10078 VSS 0.036461f
C9023 PAD.n10079 VSS 0.036461f
C9024 PAD.n10080 VSS 0.036461f
C9025 PAD.n10082 VSS 0.036461f
C9026 PAD.n10083 VSS 0.036461f
C9027 PAD.n10084 VSS 0.036461f
C9028 PAD.n10086 VSS 0.036461f
C9029 PAD.n10087 VSS 0.036461f
C9030 PAD.n10088 VSS 0.036461f
C9031 PAD.n10090 VSS 0.036461f
C9032 PAD.n10091 VSS 0.036461f
C9033 PAD.n10092 VSS 0.036461f
C9034 PAD.n10094 VSS 0.036461f
C9035 PAD.n10095 VSS 0.036461f
C9036 PAD.n10096 VSS 0.036461f
C9037 PAD.n10098 VSS 0.036461f
C9038 PAD.n10099 VSS 0.036461f
C9039 PAD.n10100 VSS 0.036461f
C9040 PAD.n10102 VSS 0.036461f
C9041 PAD.n10103 VSS 0.036461f
C9042 PAD.n10104 VSS 0.036461f
C9043 PAD.n10105 VSS 0.023109f
C9044 PAD.n10106 VSS 0.023109f
C9045 PAD.n10108 VSS 0.036461f
C9046 PAD.n10110 VSS 0.036461f
C9047 PAD.n10112 VSS 0.036461f
C9048 PAD.n10113 VSS 0.036461f
C9049 PAD.n10114 VSS 0.036461f
C9050 PAD.n10115 VSS 0.036461f
C9051 PAD.n10116 VSS 0.036461f
C9052 PAD.n10117 VSS 0.036461f
C9053 PAD.n10118 VSS 0.036461f
C9054 PAD.n10120 VSS 0.036461f
C9055 PAD.n10122 VSS 0.036461f
C9056 PAD.n10124 VSS 0.036461f
C9057 PAD.n10125 VSS 0.036461f
C9058 PAD.n10126 VSS 0.036461f
C9059 PAD.n10127 VSS 0.036461f
C9060 PAD.n10128 VSS 0.036461f
C9061 PAD.n10129 VSS 0.036461f
C9062 PAD.n10130 VSS 0.036461f
C9063 PAD.n10132 VSS 0.036461f
C9064 PAD.n10134 VSS 0.036461f
C9065 PAD.n10136 VSS 0.036461f
C9066 PAD.n10137 VSS 0.036461f
C9067 PAD.n10138 VSS 0.036461f
C9068 PAD.n10139 VSS 0.036461f
C9069 PAD.n10140 VSS 0.036461f
C9070 PAD.n10141 VSS 0.036461f
C9071 PAD.n10142 VSS 0.036461f
C9072 PAD.n10144 VSS 0.036461f
C9073 PAD.n10146 VSS 0.036461f
C9074 PAD.n10148 VSS 0.036461f
C9075 PAD.n10149 VSS 0.036461f
C9076 PAD.n10150 VSS 0.036461f
C9077 PAD.n10151 VSS 0.036461f
C9078 PAD.n10152 VSS 0.036461f
C9079 PAD.n10153 VSS 0.036461f
C9080 PAD.n10154 VSS 0.036461f
C9081 PAD.n10156 VSS 0.036461f
C9082 PAD.n10158 VSS 0.036461f
C9083 PAD.n10160 VSS 0.036461f
C9084 PAD.n10161 VSS 0.036461f
C9085 PAD.n10162 VSS 0.036461f
C9086 PAD.n10163 VSS 0.036461f
C9087 PAD.n10164 VSS 0.036461f
C9088 PAD.n10165 VSS 0.036461f
C9089 PAD.n10166 VSS 0.036461f
C9090 PAD.n10168 VSS 0.036461f
C9091 PAD.n10170 VSS 0.036461f
C9092 PAD.n10172 VSS 0.036461f
C9093 PAD.n10173 VSS 0.036461f
C9094 PAD.n10174 VSS 0.036461f
C9095 PAD.n10175 VSS 0.036461f
C9096 PAD.n10176 VSS 0.036461f
C9097 PAD.n10177 VSS 0.036461f
C9098 PAD.n10178 VSS 0.036461f
C9099 PAD.n10180 VSS 0.036461f
C9100 PAD.n10182 VSS 0.036461f
C9101 PAD.n10184 VSS 0.036461f
C9102 PAD.n10185 VSS 0.036461f
C9103 PAD.n10186 VSS 0.036461f
C9104 PAD.n10187 VSS 0.036461f
C9105 PAD.n10188 VSS 0.036461f
C9106 PAD.n10189 VSS 0.036461f
C9107 PAD.n10190 VSS 0.036461f
C9108 PAD.n10192 VSS 0.036461f
C9109 PAD.n10194 VSS 0.036461f
C9110 PAD.n10196 VSS 0.036461f
C9111 PAD.n10197 VSS 0.036461f
C9112 PAD.n10198 VSS 0.036461f
C9113 PAD.n10199 VSS 0.036461f
C9114 PAD.n10200 VSS 0.036461f
C9115 PAD.n10201 VSS 0.036461f
C9116 PAD.n10202 VSS 0.036461f
C9117 PAD.n10204 VSS 0.036461f
C9118 PAD.n10206 VSS 0.036461f
C9119 PAD.n10208 VSS 0.036461f
C9120 PAD.n10209 VSS 0.036461f
C9121 PAD.n10210 VSS 0.036461f
C9122 PAD.n10211 VSS 0.036461f
C9123 PAD.n10212 VSS 0.036461f
C9124 PAD.n10213 VSS 0.036461f
C9125 PAD.n10214 VSS 0.036461f
C9126 PAD.n10216 VSS 0.036461f
C9127 PAD.n10218 VSS 0.036461f
C9128 PAD.n10220 VSS 0.036461f
C9129 PAD.n10221 VSS 0.036461f
C9130 PAD.n10222 VSS 0.036461f
C9131 PAD.n10223 VSS 0.036461f
C9132 PAD.n10224 VSS 0.036461f
C9133 PAD.n10225 VSS 0.036461f
C9134 PAD.n10226 VSS 0.036461f
C9135 PAD.n10228 VSS 0.036461f
C9136 PAD.n10230 VSS 0.036461f
C9137 PAD.n10232 VSS 0.036461f
C9138 PAD.n10233 VSS 0.036461f
C9139 PAD.n10234 VSS 0.036461f
C9140 PAD.n10235 VSS 0.036461f
C9141 PAD.n10236 VSS 0.036461f
C9142 PAD.n10237 VSS 0.036461f
C9143 PAD.n10238 VSS 0.036461f
C9144 PAD.n10240 VSS 0.036461f
C9145 PAD.n10242 VSS 0.036461f
C9146 PAD.n10244 VSS 0.036461f
C9147 PAD.n10245 VSS 0.036461f
C9148 PAD.n10246 VSS 0.036461f
C9149 PAD.n10247 VSS 0.036461f
C9150 PAD.n10248 VSS 0.036461f
C9151 PAD.n10249 VSS 0.036461f
C9152 PAD.n10250 VSS 0.036461f
C9153 PAD.n10252 VSS 0.036461f
C9154 PAD.n10254 VSS 0.036461f
C9155 PAD.n10256 VSS 0.036461f
C9156 PAD.n10257 VSS 0.036461f
C9157 PAD.n10258 VSS 0.036461f
C9158 PAD.n10259 VSS 0.036461f
C9159 PAD.n10260 VSS 0.036461f
C9160 PAD.n10261 VSS 0.036461f
C9161 PAD.n10262 VSS 0.036461f
C9162 PAD.n10264 VSS 0.036461f
C9163 PAD.n10266 VSS 0.036461f
C9164 PAD.n10268 VSS 0.036461f
C9165 PAD.n10269 VSS 0.036461f
C9166 PAD.n10270 VSS 0.036461f
C9167 PAD.n10271 VSS 0.036461f
C9168 PAD.n10272 VSS 0.036461f
C9169 PAD.n10273 VSS 0.036461f
C9170 PAD.n10274 VSS 0.036461f
C9171 PAD.n10276 VSS 0.036461f
C9172 PAD.n10278 VSS 0.036461f
C9173 PAD.n10280 VSS 0.036461f
C9174 PAD.n10281 VSS 0.036461f
C9175 PAD.n10282 VSS 0.036461f
C9176 PAD.n10283 VSS 0.036461f
C9177 PAD.n10284 VSS 0.036461f
C9178 PAD.n10285 VSS 0.036461f
C9179 PAD.n10286 VSS 0.036461f
C9180 PAD.n10288 VSS 0.036461f
C9181 PAD.n10290 VSS 0.036461f
C9182 PAD.n10292 VSS 0.036461f
C9183 PAD.n10293 VSS 0.036461f
C9184 PAD.n10294 VSS 0.036461f
C9185 PAD.n10295 VSS 0.036461f
C9186 PAD.n10296 VSS 0.036461f
C9187 PAD.n10297 VSS 0.036461f
C9188 PAD.n10298 VSS 0.036461f
C9189 PAD.n10300 VSS 0.036461f
C9190 PAD.n10302 VSS 0.036461f
C9191 PAD.n10304 VSS 0.036461f
C9192 PAD.n10305 VSS 0.036461f
C9193 PAD.n10306 VSS 0.036461f
C9194 PAD.n10307 VSS 0.036461f
C9195 PAD.n10308 VSS 0.036461f
C9196 PAD.n10309 VSS 0.036461f
C9197 PAD.n10310 VSS 0.036461f
C9198 PAD.n10312 VSS 0.036461f
C9199 PAD.n10314 VSS 0.036461f
C9200 PAD.n10316 VSS 0.036461f
C9201 PAD.n10317 VSS 0.036461f
C9202 PAD.n10318 VSS 0.036461f
C9203 PAD.n10319 VSS 0.036461f
C9204 PAD.n10320 VSS 0.036461f
C9205 PAD.n10321 VSS 0.036461f
C9206 PAD.n10322 VSS 0.036461f
C9207 PAD.n10324 VSS 0.036461f
C9208 PAD.n10326 VSS 0.036461f
C9209 PAD.n10328 VSS 0.036461f
C9210 PAD.n10329 VSS 0.036461f
C9211 PAD.n10330 VSS 0.036461f
C9212 PAD.n10331 VSS 0.036461f
C9213 PAD.n10332 VSS 0.036461f
C9214 PAD.n10333 VSS 0.036461f
C9215 PAD.n10334 VSS 0.036461f
C9216 PAD.n10336 VSS 0.036461f
C9217 PAD.n10338 VSS 0.036461f
C9218 PAD.n10340 VSS 0.036461f
C9219 PAD.n10341 VSS 0.036461f
C9220 PAD.n10342 VSS 0.036461f
C9221 PAD.n10343 VSS 0.036461f
C9222 PAD.n10344 VSS 0.036461f
C9223 PAD.n10345 VSS 0.036461f
C9224 PAD.n10346 VSS 0.036461f
C9225 PAD.n10347 VSS 0.036461f
C9226 PAD.n10349 VSS 0.036461f
C9227 PAD.n10351 VSS 0.036461f
C9228 PAD.n10353 VSS 0.023109f
C9229 PAD.n10354 VSS 0.023109f
C9230 PAD.n10355 VSS 0.030555f
C9231 PAD.n10356 VSS 0.040026f
C9232 PAD.n10357 VSS 0.033773f
C9233 PAD.n10358 VSS 0.024317f
C9234 PAD.n10359 VSS 0.027844f
C9235 PAD.n10360 VSS 0.027844f
C9236 PAD.n10361 VSS 0.522934f
C9237 PAD.n10362 VSS 0.261467f
C9238 PAD.n10363 VSS 0.04501f
C9239 PAD.n10364 VSS 0.04501f
C9240 PAD.n10365 VSS 0.035657f
C9241 PAD.n10366 VSS 8.75696f
C9242 PAD.n10367 VSS 0.041766f
C9243 PAD.n10368 VSS 0.053234f
C9244 PAD.n10369 VSS 0.047208f
C9245 PAD.n10370 VSS 0.062274f
C9246 PAD.n10371 VSS 0.069765f
C9247 PAD.n10372 VSS 0.069765f
C9248 PAD.n10373 VSS 0.700534f
C9249 PAD.n10374 VSS 0.592001f
C9250 PAD.n10375 VSS 0.047905f
C9251 PAD.n10376 VSS 0.047905f
C9252 PAD.n10377 VSS 0.029436f
C9253 PAD.n10378 VSS 0.025768f
C9254 PAD.n10379 VSS 0.025768f
C9255 PAD.n10380 VSS 0.022505f
C9256 PAD.n10381 VSS 0.033773f
C9257 PAD.n10382 VSS 0.030555f
C9258 PAD.n10383 VSS 0.036461f
C9259 PAD.n10384 VSS 0.036461f
C9260 PAD.n10385 VSS 0.036461f
C9261 PAD.n10387 VSS 0.023109f
C9262 PAD.n10388 VSS 0.439067f
C9263 PAD.n10389 VSS 0.330534f
C9264 PAD.n10390 VSS 0.051761f
C9265 PAD.n10391 VSS 0.051761f
C9266 PAD.n10392 VSS 0.046203f
C9267 PAD.n10393 VSS 0.062274f
C9268 PAD.n10394 VSS 0.054238f
C9269 PAD.n10395 VSS 0.060763f
C9270 PAD.n10396 VSS 0.060763f
C9271 PAD.n10397 VSS 0.187466f
C9272 PAD.n10398 VSS 0.611734f
C9273 PAD.n10399 VSS 0.043408f
C9274 PAD.n10400 VSS 0.043408f
C9275 PAD.n10401 VSS 0.037911f
C9276 PAD.n10402 VSS 0.033773f
C9277 PAD.n10403 VSS 0.042895f
C9278 PAD.n10404 VSS 0.026432f
C9279 PAD.n10405 VSS 0.030265f
C9280 PAD.n10406 VSS 0.030265f
C9281 PAD.n10407 VSS 0.1924f
C9282 PAD.n10408 VSS 0.513067f
C9283 PAD.n10409 VSS 0.043885f
C9284 PAD.n10410 VSS 0.043885f
C9285 PAD.n10411 VSS 0.039172f
C9286 PAD.n10412 VSS 0.062274f
C9287 PAD.n10413 VSS 0.036461f
C9288 PAD.n10414 VSS 0.036461f
C9289 PAD.n10415 VSS 0.036461f
C9290 PAD.n10417 VSS 0.036461f
C9291 PAD.n10418 VSS 0.036461f
C9292 PAD.n10419 VSS 0.036461f
C9293 PAD.n10420 VSS 0.036461f
C9294 PAD.n10422 VSS 0.036461f
C9295 PAD.n10423 VSS 0.036461f
C9296 PAD.n10424 VSS 0.036461f
C9297 PAD.n10425 VSS 0.036461f
C9298 PAD.n10427 VSS 0.036461f
C9299 PAD.n10428 VSS 0.036461f
C9300 PAD.n10429 VSS 0.036461f
C9301 PAD.n10430 VSS 0.036461f
C9302 PAD.n10432 VSS 0.036461f
C9303 PAD.n10433 VSS 0.036461f
C9304 PAD.n10434 VSS 0.036461f
C9305 PAD.n10435 VSS 0.036461f
C9306 PAD.n10437 VSS 0.036461f
C9307 PAD.n10438 VSS 0.036461f
C9308 PAD.n10439 VSS 0.036461f
C9309 PAD.n10440 VSS 0.036461f
C9310 PAD.n10442 VSS 0.036461f
C9311 PAD.n10443 VSS 0.036461f
C9312 PAD.n10444 VSS 0.036461f
C9313 PAD.n10445 VSS 0.036461f
C9314 PAD.n10447 VSS 0.036461f
C9315 PAD.n10448 VSS 0.036461f
C9316 PAD.n10449 VSS 0.036461f
C9317 PAD.n10450 VSS 0.036461f
C9318 PAD.n10452 VSS 0.036461f
C9319 PAD.n10453 VSS 0.036461f
C9320 PAD.n10454 VSS 0.036461f
C9321 PAD.n10455 VSS 0.036461f
C9322 PAD.n10457 VSS 0.036461f
C9323 PAD.n10458 VSS 0.036461f
C9324 PAD.n10459 VSS 0.036461f
C9325 PAD.n10460 VSS 0.036461f
C9326 PAD.n10462 VSS 0.036461f
C9327 PAD.n10463 VSS 0.036461f
C9328 PAD.n10464 VSS 0.036461f
C9329 PAD.n10465 VSS 0.036461f
C9330 PAD.n10467 VSS 0.036461f
C9331 PAD.n10468 VSS 0.036461f
C9332 PAD.n10469 VSS 0.036461f
C9333 PAD.n10470 VSS 0.036461f
C9334 PAD.n10472 VSS 0.036461f
C9335 PAD.n10473 VSS 0.036461f
C9336 PAD.n10474 VSS 0.036461f
C9337 PAD.n10475 VSS 0.036461f
C9338 PAD.n10477 VSS 0.036461f
C9339 PAD.n10478 VSS 0.036461f
C9340 PAD.n10479 VSS 0.036461f
C9341 PAD.n10480 VSS 0.036461f
C9342 PAD.n10482 VSS 0.036461f
C9343 PAD.n10483 VSS 0.036461f
C9344 PAD.n10484 VSS 0.036461f
C9345 PAD.n10485 VSS 0.036461f
C9346 PAD.n10487 VSS 0.036461f
C9347 PAD.n10488 VSS 0.036461f
C9348 PAD.n10489 VSS 0.036461f
C9349 PAD.n10490 VSS 0.036461f
C9350 PAD.n10492 VSS 0.036461f
C9351 PAD.n10493 VSS 0.036461f
C9352 PAD.n10494 VSS 0.036461f
C9353 PAD.n10495 VSS 0.036461f
C9354 PAD.n10497 VSS 0.036461f
C9355 PAD.n10498 VSS 0.036461f
C9356 PAD.n10499 VSS 0.036461f
C9357 PAD.n10500 VSS 0.036461f
C9358 PAD.n10502 VSS 0.036461f
C9359 PAD.n10503 VSS 0.036461f
C9360 PAD.n10504 VSS 0.036461f
C9361 PAD.n10505 VSS 0.036461f
C9362 PAD.n10507 VSS 0.036461f
C9363 PAD.n10508 VSS 0.036461f
C9364 PAD.n10509 VSS 0.036461f
C9365 PAD.n10510 VSS 0.036461f
C9366 PAD.n10512 VSS 0.036461f
C9367 PAD.n10513 VSS 0.036461f
C9368 PAD.n10515 VSS 0.036461f
C9369 PAD.n10516 VSS 0.036461f
C9370 PAD.n10517 VSS 0.036461f
C9371 PAD.n10518 VSS 0.036461f
C9372 PAD.n10519 VSS 0.036461f
C9373 PAD.n10520 VSS 0.036461f
C9374 PAD.n10521 VSS 0.036461f
C9375 PAD.n10522 VSS 0.036461f
C9376 PAD.n10524 VSS 0.036461f
C9377 PAD.n10525 VSS 0.036461f
C9378 PAD.n10526 VSS 0.036461f
C9379 PAD.n10527 VSS 0.036461f
C9380 PAD.n10528 VSS 0.036461f
C9381 PAD.n10529 VSS 0.036461f
C9382 PAD.n10530 VSS 0.036461f
C9383 PAD.n10531 VSS 0.036461f
C9384 PAD.n10533 VSS 0.036461f
C9385 PAD.n10534 VSS 0.036461f
C9386 PAD.n10535 VSS 0.036461f
C9387 PAD.n10536 VSS 0.036461f
C9388 PAD.n10537 VSS 0.036461f
C9389 PAD.n10538 VSS 0.036461f
C9390 PAD.n10539 VSS 0.036461f
C9391 PAD.n10540 VSS 0.036461f
C9392 PAD.n10542 VSS 0.036461f
C9393 PAD.n10543 VSS 0.036461f
C9394 PAD.n10544 VSS 0.036461f
C9395 PAD.n10545 VSS 0.036461f
C9396 PAD.n10546 VSS 0.036461f
C9397 PAD.n10547 VSS 0.036461f
C9398 PAD.n10548 VSS 0.036461f
C9399 PAD.n10549 VSS 0.036461f
C9400 PAD.n10551 VSS 0.036461f
C9401 PAD.n10552 VSS 0.036461f
C9402 PAD.n10553 VSS 0.036461f
C9403 PAD.n10554 VSS 0.036461f
C9404 PAD.n10555 VSS 0.036461f
C9405 PAD.n10556 VSS 0.036461f
C9406 PAD.n10557 VSS 0.036461f
C9407 PAD.n10558 VSS 0.036461f
C9408 PAD.n10560 VSS 0.036461f
C9409 PAD.n10561 VSS 0.036461f
C9410 PAD.n10562 VSS 0.036461f
C9411 PAD.n10563 VSS 0.036461f
C9412 PAD.n10564 VSS 0.036461f
C9413 PAD.n10565 VSS 0.036461f
C9414 PAD.n10566 VSS 0.036461f
C9415 PAD.n10567 VSS 0.036461f
C9416 PAD.n10569 VSS 0.036461f
C9417 PAD.n10570 VSS 0.036461f
C9418 PAD.n10571 VSS 0.036461f
C9419 PAD.n10572 VSS 0.036461f
C9420 PAD.n10573 VSS 0.036461f
C9421 PAD.n10574 VSS 0.036461f
C9422 PAD.n10575 VSS 0.036461f
C9423 PAD.n10576 VSS 0.036461f
C9424 PAD.n10578 VSS 0.036461f
C9425 PAD.n10579 VSS 0.036461f
C9426 PAD.n10580 VSS 0.036461f
C9427 PAD.n10581 VSS 0.036461f
C9428 PAD.n10582 VSS 0.036461f
C9429 PAD.n10583 VSS 0.036461f
C9430 PAD.n10584 VSS 0.036461f
C9431 PAD.n10585 VSS 0.036461f
C9432 PAD.n10587 VSS 0.036461f
C9433 PAD.n10588 VSS 0.036461f
C9434 PAD.n10589 VSS 0.036461f
C9435 PAD.n10590 VSS 0.036461f
C9436 PAD.n10591 VSS 0.036461f
C9437 PAD.n10592 VSS 0.036461f
C9438 PAD.n10593 VSS 0.036461f
C9439 PAD.n10594 VSS 0.036461f
C9440 PAD.n10596 VSS 0.036461f
C9441 PAD.n10597 VSS 0.036461f
C9442 PAD.n10598 VSS 0.036461f
C9443 PAD.n10599 VSS 0.036461f
C9444 PAD.n10600 VSS 0.036461f
C9445 PAD.n10601 VSS 0.036461f
C9446 PAD.n10602 VSS 0.036461f
C9447 PAD.n10603 VSS 0.036461f
C9448 PAD.n10605 VSS 0.036461f
C9449 PAD.n10606 VSS 0.036461f
C9450 PAD.n10607 VSS 0.036461f
C9451 PAD.n10608 VSS 0.036461f
C9452 PAD.n10609 VSS 0.036461f
C9453 PAD.n10610 VSS 0.036461f
C9454 PAD.n10611 VSS 0.036461f
C9455 PAD.n10612 VSS 0.036461f
C9456 PAD.n10614 VSS 0.036461f
C9457 PAD.n10615 VSS 0.036461f
C9458 PAD.n10616 VSS 0.036461f
C9459 PAD.n10617 VSS 0.036461f
C9460 PAD.n10618 VSS 0.036461f
C9461 PAD.n10619 VSS 0.036461f
C9462 PAD.n10620 VSS 0.036461f
C9463 PAD.n10621 VSS 0.036461f
C9464 PAD.n10623 VSS 0.036461f
C9465 PAD.n10624 VSS 0.036461f
C9466 PAD.n10625 VSS 0.036461f
C9467 PAD.n10626 VSS 0.036461f
C9468 PAD.n10627 VSS 0.036461f
C9469 PAD.n10628 VSS 0.036461f
C9470 PAD.n10629 VSS 0.036461f
C9471 PAD.n10630 VSS 0.036461f
C9472 PAD.n10632 VSS 0.036461f
C9473 PAD.n10633 VSS 0.036461f
C9474 PAD.n10634 VSS 0.036461f
C9475 PAD.n10635 VSS 0.036461f
C9476 PAD.n10636 VSS 0.036461f
C9477 PAD.n10637 VSS 0.036461f
C9478 PAD.n10638 VSS 0.036461f
C9479 PAD.n10639 VSS 0.036461f
C9480 PAD.n10641 VSS 0.036461f
C9481 PAD.n10642 VSS 0.036461f
C9482 PAD.n10643 VSS 0.036461f
C9483 PAD.n10644 VSS 0.036461f
C9484 PAD.n10645 VSS 0.036461f
C9485 PAD.n10646 VSS 0.036461f
C9486 PAD.n10647 VSS 0.036461f
C9487 PAD.n10648 VSS 0.036461f
C9488 PAD.n10650 VSS 0.036461f
C9489 PAD.n10651 VSS 0.036461f
C9490 PAD.n10652 VSS 0.036461f
C9491 PAD.n10653 VSS 0.036461f
C9492 PAD.n10654 VSS 0.036461f
C9493 PAD.n10655 VSS 0.036461f
C9494 PAD.n10656 VSS 0.036461f
C9495 PAD.n10657 VSS 0.036461f
C9496 PAD.n10659 VSS 0.036461f
C9497 PAD.n10660 VSS 0.036461f
C9498 PAD.n10661 VSS 0.036461f
C9499 PAD.n10662 VSS 0.036461f
C9500 PAD.n10663 VSS 0.036461f
C9501 PAD.n10664 VSS 0.036461f
C9502 PAD.n10665 VSS 0.036461f
C9503 PAD.n10666 VSS 0.036461f
C9504 PAD.n10668 VSS 0.036461f
C9505 PAD.n10669 VSS 0.036461f
C9506 PAD.n10670 VSS 0.036461f
C9507 PAD.n10671 VSS 0.036461f
C9508 PAD.n10672 VSS 0.036461f
C9509 PAD.n10673 VSS 0.036461f
C9510 PAD.n10674 VSS 0.036461f
C9511 PAD.n10675 VSS 0.036461f
C9512 PAD.n10677 VSS 0.036461f
C9513 PAD.n10678 VSS 0.036461f
C9514 PAD.n10679 VSS 0.036461f
C9515 PAD.n10680 VSS 0.036461f
C9516 PAD.n10681 VSS 0.036461f
C9517 PAD.n10682 VSS 0.036461f
C9518 PAD.n10683 VSS 0.036461f
C9519 PAD.n10684 VSS 0.036461f
C9520 PAD.n10686 VSS 0.036461f
C9521 PAD.n10687 VSS 0.036461f
C9522 PAD.n10688 VSS 0.036461f
C9523 PAD.n10689 VSS 0.036461f
C9524 PAD.n10690 VSS 0.036461f
C9525 PAD.n10691 VSS 0.036461f
C9526 PAD.n10693 VSS 0.036461f
C9527 PAD.n10694 VSS 0.036461f
C9528 PAD.n10695 VSS 0.023109f
C9529 PAD.n10696 VSS 0.03338f
C9530 PAD.n10697 VSS 0.046286f
C9531 PAD.n10698 VSS 0.061269f
C9532 PAD.n10699 VSS 0.06864f
C9533 PAD.n10700 VSS 0.06864f
C9534 PAD.n10701 VSS 0.700534f
C9535 PAD.n10702 VSS 0.226933f
C9536 PAD.n10703 VSS 0.038912f
C9537 PAD.n10704 VSS 0.038912f
C9538 PAD.n10705 VSS 0.029436f
C9539 PAD.n10706 VSS 0.034761f
C9540 PAD.n10707 VSS 0.034761f
C9541 PAD.n10708 VSS 0.030359f
C9542 PAD.n10709 VSS 0.033773f
C9543 PAD.n10710 VSS 0.030555f
C9544 PAD.n10711 VSS 0.036461f
C9545 PAD.n10712 VSS 0.036461f
C9546 PAD.n10713 VSS 0.036461f
C9547 PAD.n10715 VSS 0.023109f
C9548 PAD.n10716 VSS 0.3404f
C9549 PAD.n10717 VSS 0.616668f
C9550 PAD.n10718 VSS 0.611734f
C9551 PAD.n10719 VSS 0.656134f
C9552 PAD.n10720 VSS 0.069765f
C9553 PAD.n10721 VSS 0.069765f
C9554 PAD.n10722 VSS 0.062274f
C9555 PAD.n10723 VSS 0.062274f
C9556 PAD.n10724 VSS 0.037163f
C9557 PAD.n10725 VSS 0.041634f
C9558 PAD.n10726 VSS 0.041634f
C9559 PAD.n10727 VSS 0.616668f
C9560 PAD.n10728 VSS 0.246666f
C9561 PAD.n10729 VSS 0.034415f
C9562 PAD.n10730 VSS 0.034415f
C9563 PAD.n10731 VSS 0.030057f
C9564 PAD.n10732 VSS 0.033773f
C9565 PAD.n10733 VSS 0.034286f
C9566 PAD.n10734 VSS 0.030555f
C9567 PAD.n10735 VSS 0.042895f
C9568 PAD.n10736 VSS 0.029436f
C9569 PAD.n10737 VSS 0.049115f
C9570 PAD.n10738 VSS 0.029436f
C9571 PAD.n10739 VSS 0.049115f
C9572 PAD.n10740 VSS 0.2072f
C9573 PAD.n10741 VSS 0.611734f
C9574 PAD.n10742 VSS 0.055137f
C9575 PAD.n10743 VSS 0.068077f
C9576 PAD.n10744 VSS 0.055137f
C9577 PAD.n10745 VSS 0.068077f
C9578 PAD.n10746 VSS 0.044194f
C9579 PAD.n10747 VSS 0.036461f
C9580 PAD.n10748 VSS 0.039761f
C9581 PAD.n10749 VSS 0.036461f
C9582 PAD.n10750 VSS 0.039761f
C9583 PAD.n10751 VSS 0.049511f
C9584 PAD.n10752 VSS 0.049511f
C9585 PAD.n10753 VSS 0.2072f
C9586 PAD.n10754 VSS 0.596934f
C9587 PAD.n10755 VSS 0.508134f
C9588 PAD.n10757 VSS 0.036461f
C9589 PAD.n10758 VSS 0.036461f
C9590 PAD.n10759 VSS 0.036461f
C9591 PAD.n10761 VSS 0.036461f
C9592 PAD.n10762 VSS 0.036461f
C9593 PAD.n10763 VSS 0.036461f
C9594 PAD.n10765 VSS 0.036461f
C9595 PAD.n10766 VSS 0.036461f
C9596 PAD.n10767 VSS 0.036461f
C9597 PAD.n10769 VSS 0.036461f
C9598 PAD.n10770 VSS 0.036461f
C9599 PAD.n10771 VSS 0.036461f
C9600 PAD.n10773 VSS 0.036461f
C9601 PAD.n10774 VSS 0.036461f
C9602 PAD.n10775 VSS 0.036461f
C9603 PAD.n10777 VSS 0.036461f
C9604 PAD.n10778 VSS 0.036461f
C9605 PAD.n10779 VSS 0.036461f
C9606 PAD.n10781 VSS 0.036461f
C9607 PAD.n10782 VSS 0.036461f
C9608 PAD.n10783 VSS 0.036461f
C9609 PAD.n10785 VSS 0.036461f
C9610 PAD.n10786 VSS 0.036461f
C9611 PAD.n10787 VSS 0.036461f
C9612 PAD.n10789 VSS 0.036461f
C9613 PAD.n10790 VSS 0.036461f
C9614 PAD.n10791 VSS 0.036461f
C9615 PAD.n10793 VSS 0.036461f
C9616 PAD.n10794 VSS 0.036461f
C9617 PAD.n10795 VSS 0.036461f
C9618 PAD.n10797 VSS 0.036461f
C9619 PAD.n10798 VSS 0.036461f
C9620 PAD.n10799 VSS 0.036461f
C9621 PAD.n10801 VSS 0.036461f
C9622 PAD.n10802 VSS 0.036461f
C9623 PAD.n10803 VSS 0.036461f
C9624 PAD.n10805 VSS 0.036461f
C9625 PAD.n10806 VSS 0.036461f
C9626 PAD.n10807 VSS 0.036461f
C9627 PAD.n10809 VSS 0.036461f
C9628 PAD.n10810 VSS 0.036461f
C9629 PAD.n10811 VSS 0.036461f
C9630 PAD.n10813 VSS 0.036461f
C9631 PAD.n10814 VSS 0.036461f
C9632 PAD.n10815 VSS 0.036461f
C9633 PAD.n10817 VSS 0.036461f
C9634 PAD.n10818 VSS 0.036461f
C9635 PAD.n10819 VSS 0.036461f
C9636 PAD.n10821 VSS 0.036461f
C9637 PAD.n10822 VSS 0.036461f
C9638 PAD.n10823 VSS 0.036461f
C9639 PAD.n10825 VSS 0.036461f
C9640 PAD.n10826 VSS 0.036461f
C9641 PAD.n10827 VSS 0.036461f
C9642 PAD.n10829 VSS 0.036461f
C9643 PAD.n10830 VSS 0.036461f
C9644 PAD.n10831 VSS 0.036461f
C9645 PAD.n10833 VSS 0.036461f
C9646 PAD.n10834 VSS 0.036461f
C9647 PAD.n10835 VSS 0.036461f
C9648 PAD.n10837 VSS 0.023109f
C9649 PAD.n10838 VSS 0.023109f
C9650 PAD.n10839 VSS 0.036461f
C9651 PAD.n10840 VSS 0.036461f
C9652 PAD.n10841 VSS 0.036461f
C9653 PAD.n10843 VSS 0.036461f
C9654 PAD.n10845 VSS 0.036461f
C9655 PAD.n10847 VSS 0.036461f
C9656 PAD.n10848 VSS 0.036461f
C9657 PAD.n10849 VSS 0.036461f
C9658 PAD.n10850 VSS 0.036461f
C9659 PAD.n10851 VSS 0.036461f
C9660 PAD.n10852 VSS 0.036461f
C9661 PAD.n10853 VSS 0.036461f
C9662 PAD.n10855 VSS 0.036461f
C9663 PAD.n10857 VSS 0.036461f
C9664 PAD.n10859 VSS 0.036461f
C9665 PAD.n10860 VSS 0.036461f
C9666 PAD.n10861 VSS 0.036461f
C9667 PAD.n10862 VSS 0.036461f
C9668 PAD.n10863 VSS 0.036461f
C9669 PAD.n10864 VSS 0.036461f
C9670 PAD.n10865 VSS 0.036461f
C9671 PAD.n10867 VSS 0.036461f
C9672 PAD.n10869 VSS 0.036461f
C9673 PAD.n10871 VSS 0.036461f
C9674 PAD.n10872 VSS 0.036461f
C9675 PAD.n10873 VSS 0.036461f
C9676 PAD.n10874 VSS 0.036461f
C9677 PAD.n10875 VSS 0.036461f
C9678 PAD.n10876 VSS 0.036461f
C9679 PAD.n10877 VSS 0.036461f
C9680 PAD.n10879 VSS 0.036461f
C9681 PAD.n10881 VSS 0.036461f
C9682 PAD.n10883 VSS 0.036461f
C9683 PAD.n10884 VSS 0.036461f
C9684 PAD.n10885 VSS 0.036461f
C9685 PAD.n10886 VSS 0.036461f
C9686 PAD.n10887 VSS 0.036461f
C9687 PAD.n10888 VSS 0.036461f
C9688 PAD.n10889 VSS 0.036461f
C9689 PAD.n10891 VSS 0.036461f
C9690 PAD.n10893 VSS 0.036461f
C9691 PAD.n10895 VSS 0.036461f
C9692 PAD.n10896 VSS 0.036461f
C9693 PAD.n10897 VSS 0.036461f
C9694 PAD.n10898 VSS 0.036461f
C9695 PAD.n10899 VSS 0.036461f
C9696 PAD.n10900 VSS 0.036461f
C9697 PAD.n10901 VSS 0.036461f
C9698 PAD.n10903 VSS 0.036461f
C9699 PAD.n10905 VSS 0.036461f
C9700 PAD.n10907 VSS 0.036461f
C9701 PAD.n10908 VSS 0.036461f
C9702 PAD.n10909 VSS 0.036461f
C9703 PAD.n10910 VSS 0.036461f
C9704 PAD.n10911 VSS 0.036461f
C9705 PAD.n10912 VSS 0.036461f
C9706 PAD.n10913 VSS 0.036461f
C9707 PAD.n10915 VSS 0.036461f
C9708 PAD.n10917 VSS 0.036461f
C9709 PAD.n10919 VSS 0.036461f
C9710 PAD.n10920 VSS 0.036461f
C9711 PAD.n10921 VSS 0.036461f
C9712 PAD.n10922 VSS 0.036461f
C9713 PAD.n10923 VSS 0.036461f
C9714 PAD.n10924 VSS 0.036461f
C9715 PAD.n10925 VSS 0.036461f
C9716 PAD.n10927 VSS 0.036461f
C9717 PAD.n10929 VSS 0.036461f
C9718 PAD.n10931 VSS 0.036461f
C9719 PAD.n10932 VSS 0.036461f
C9720 PAD.n10933 VSS 0.036461f
C9721 PAD.n10934 VSS 0.036461f
C9722 PAD.n10935 VSS 0.036461f
C9723 PAD.n10936 VSS 0.036461f
C9724 PAD.n10937 VSS 0.036461f
C9725 PAD.n10939 VSS 0.036461f
C9726 PAD.n10941 VSS 0.036461f
C9727 PAD.n10943 VSS 0.036461f
C9728 PAD.n10944 VSS 0.036461f
C9729 PAD.n10945 VSS 0.036461f
C9730 PAD.n10946 VSS 0.036461f
C9731 PAD.n10947 VSS 0.036461f
C9732 PAD.n10948 VSS 0.036461f
C9733 PAD.n10949 VSS 0.036461f
C9734 PAD.n10951 VSS 0.036461f
C9735 PAD.n10953 VSS 0.036461f
C9736 PAD.n10955 VSS 0.036461f
C9737 PAD.n10956 VSS 0.036461f
C9738 PAD.n10957 VSS 0.036461f
C9739 PAD.n10958 VSS 0.036461f
C9740 PAD.n10959 VSS 0.036461f
C9741 PAD.n10960 VSS 0.036461f
C9742 PAD.n10961 VSS 0.036461f
C9743 PAD.n10963 VSS 0.036461f
C9744 PAD.n10965 VSS 0.036461f
C9745 PAD.n10967 VSS 0.036461f
C9746 PAD.n10968 VSS 0.036461f
C9747 PAD.n10969 VSS 0.036461f
C9748 PAD.n10970 VSS 0.036461f
C9749 PAD.n10971 VSS 0.036461f
C9750 PAD.n10972 VSS 0.036461f
C9751 PAD.n10973 VSS 0.036461f
C9752 PAD.n10975 VSS 0.036461f
C9753 PAD.n10977 VSS 0.036461f
C9754 PAD.n10979 VSS 0.036461f
C9755 PAD.n10980 VSS 0.036461f
C9756 PAD.n10981 VSS 0.036461f
C9757 PAD.n10982 VSS 0.036461f
C9758 PAD.n10983 VSS 0.036461f
C9759 PAD.n10984 VSS 0.036461f
C9760 PAD.n10985 VSS 0.036461f
C9761 PAD.n10987 VSS 0.036461f
C9762 PAD.n10989 VSS 0.036461f
C9763 PAD.n10991 VSS 0.036461f
C9764 PAD.n10992 VSS 0.036461f
C9765 PAD.n10993 VSS 0.036461f
C9766 PAD.n10994 VSS 0.036461f
C9767 PAD.n10995 VSS 0.036461f
C9768 PAD.n10996 VSS 0.036461f
C9769 PAD.n10997 VSS 0.036461f
C9770 PAD.n10999 VSS 0.036461f
C9771 PAD.n11001 VSS 0.036461f
C9772 PAD.n11003 VSS 0.036461f
C9773 PAD.n11004 VSS 0.036461f
C9774 PAD.n11005 VSS 0.036461f
C9775 PAD.n11006 VSS 0.036461f
C9776 PAD.n11007 VSS 0.036461f
C9777 PAD.n11008 VSS 0.036461f
C9778 PAD.n11009 VSS 0.036461f
C9779 PAD.n11011 VSS 0.036461f
C9780 PAD.n11013 VSS 0.036461f
C9781 PAD.n11015 VSS 0.036461f
C9782 PAD.n11016 VSS 0.036461f
C9783 PAD.n11017 VSS 0.036461f
C9784 PAD.n11018 VSS 0.036461f
C9785 PAD.n11019 VSS 0.036461f
C9786 PAD.n11020 VSS 0.036461f
C9787 PAD.n11021 VSS 0.036461f
C9788 PAD.n11023 VSS 0.036461f
C9789 PAD.n11025 VSS 0.036461f
C9790 PAD.n11027 VSS 0.036461f
C9791 PAD.n11028 VSS 0.036461f
C9792 PAD.n11029 VSS 0.036461f
C9793 PAD.n11030 VSS 0.036461f
C9794 PAD.n11031 VSS 0.036461f
C9795 PAD.n11032 VSS 0.036461f
C9796 PAD.n11033 VSS 0.036461f
C9797 PAD.n11035 VSS 0.036461f
C9798 PAD.n11037 VSS 0.036461f
C9799 PAD.n11039 VSS 0.036461f
C9800 PAD.n11040 VSS 0.036461f
C9801 PAD.n11041 VSS 0.036461f
C9802 PAD.n11042 VSS 0.036461f
C9803 PAD.n11043 VSS 0.036461f
C9804 PAD.n11044 VSS 0.036461f
C9805 PAD.n11045 VSS 0.036461f
C9806 PAD.n11047 VSS 0.036461f
C9807 PAD.n11049 VSS 0.036461f
C9808 PAD.n11051 VSS 0.036461f
C9809 PAD.n11052 VSS 0.036461f
C9810 PAD.n11053 VSS 0.036461f
C9811 PAD.n11054 VSS 0.036461f
C9812 PAD.n11055 VSS 0.036461f
C9813 PAD.n11056 VSS 0.036461f
C9814 PAD.n11057 VSS 0.036461f
C9815 PAD.n11059 VSS 0.036461f
C9816 PAD.n11061 VSS 0.036461f
C9817 PAD.n11063 VSS 0.036461f
C9818 PAD.n11064 VSS 0.036461f
C9819 PAD.n11065 VSS 0.036461f
C9820 PAD.n11066 VSS 0.036461f
C9821 PAD.n11067 VSS 0.036461f
C9822 PAD.n11068 VSS 0.036461f
C9823 PAD.n11069 VSS 0.036461f
C9824 PAD.n11071 VSS 0.036461f
C9825 PAD.n11073 VSS 0.036461f
C9826 PAD.n11075 VSS 0.036461f
C9827 PAD.n11076 VSS 0.036461f
C9828 PAD.n11077 VSS 0.036461f
C9829 PAD.n11078 VSS 0.036461f
C9830 PAD.n11079 VSS 0.036461f
C9831 PAD.n11080 VSS 0.036461f
C9832 PAD.n11081 VSS 0.036461f
C9833 PAD.n11083 VSS 0.036461f
C9834 PAD.n11085 VSS 0.023109f
C9835 PAD.n11086 VSS 0.023109f
C9836 PAD.n11087 VSS 0.03338f
C9837 PAD.n11088 VSS 0.046286f
C9838 PAD.n11089 VSS 0.049216f
C9839 PAD.n11090 VSS 0.128378f
C9840 PAD.n11091 VSS 0.103613f
C9841 PAD.n11092 VSS 0.070653f
C9842 PAD.n11093 VSS 0.103613f
C9843 PAD.n11094 VSS 0.070653f
C9844 PAD.n11096 VSS 0.611735f
C9845 PAD.n11097 VSS 0.853468f
C9846 PAD.n11098 VSS 0.769602f
C9847 PAD.n11099 VSS 0.611735f
C9848 PAD.n11100 VSS 0.611735f
C9849 PAD.n11101 VSS 0.069176f
C9850 PAD.n11102 VSS 0.069176f
C9851 PAD.n11104 VSS 0.103613f
C9852 PAD.n11105 VSS 1.55894f
C9853 PAD.n11106 VSS 0.103613f
C9854 PAD.n11107 VSS 0.074916f
C9855 PAD.n11108 VSS 0.074916f
C9856 PAD.n11109 VSS 0.074916f
C9857 PAD.n11110 VSS 0.074916f
C9858 PAD.n11111 VSS 0.074916f
C9859 PAD.n11112 VSS 0.074916f
C9860 PAD.n11113 VSS 0.074916f
C9861 PAD.n11114 VSS 0.074916f
C9862 PAD.n11115 VSS 0.074916f
C9863 PAD.n11116 VSS 0.074916f
C9864 PAD.n11117 VSS 0.074916f
C9865 PAD.n11118 VSS 0.074916f
C9866 PAD.n11119 VSS 0.074916f
C9867 PAD.n11120 VSS 0.074916f
C9868 PAD.n11121 VSS 0.074916f
C9869 PAD.n11122 VSS 0.074916f
C9870 PAD.n11123 VSS 0.074916f
C9871 PAD.n11124 VSS 0.074916f
C9872 PAD.n11125 VSS 0.074916f
C9873 PAD.n11126 VSS 0.074916f
C9874 PAD.n11127 VSS 0.074916f
C9875 PAD.n11128 VSS 0.074916f
C9876 PAD.n11129 VSS 0.074916f
C9877 PAD.n11130 VSS 0.074916f
C9878 PAD.n11131 VSS 0.074916f
C9879 PAD.n11132 VSS 0.074916f
C9880 PAD.n11133 VSS 0.074916f
C9881 PAD.n11134 VSS 0.074916f
C9882 PAD.n11135 VSS 0.074916f
C9883 PAD.n11136 VSS 0.074916f
C9884 PAD.n11137 VSS 0.074916f
C9885 PAD.n11138 VSS 0.074916f
C9886 PAD.n11139 VSS 0.074916f
C9887 PAD.n11140 VSS 0.074916f
C9888 PAD.n11141 VSS 0.074916f
C9889 PAD.n11142 VSS 0.074916f
C9890 PAD.n11143 VSS 0.074916f
C9891 PAD.n11144 VSS 0.074916f
C9892 PAD.n11145 VSS 0.074916f
C9893 PAD.n11146 VSS 0.074916f
C9894 PAD.n11147 VSS 0.074916f
C9895 PAD.n11148 VSS 0.074916f
C9896 PAD.n11149 VSS 0.074916f
C9897 PAD.n11150 VSS 0.074916f
C9898 PAD.n11151 VSS 0.074916f
C9899 PAD.n11152 VSS 0.074916f
C9900 PAD.n11153 VSS 0.074916f
C9901 PAD.n11154 VSS 0.074916f
C9902 PAD.n11156 VSS 0.05951f
C9903 PAD.n11158 VSS 0.074916f
C9904 PAD.n11160 VSS 0.074916f
C9905 PAD.n11162 VSS 0.074916f
C9906 PAD.n11164 VSS 0.074916f
C9907 PAD.n11166 VSS 0.074916f
C9908 PAD.n11168 VSS 0.074916f
C9909 PAD.n11170 VSS 0.074916f
C9910 PAD.n11172 VSS 0.074916f
C9911 PAD.n11174 VSS 0.074916f
C9912 PAD.n11176 VSS 0.074916f
C9913 PAD.n11178 VSS 0.074916f
C9914 PAD.n11180 VSS 0.074916f
C9915 PAD.n11182 VSS 0.074916f
C9916 PAD.n11184 VSS 0.074916f
C9917 PAD.n11186 VSS 0.074916f
C9918 PAD.n11188 VSS 0.074916f
C9919 PAD.n11190 VSS 0.074916f
C9920 PAD.n11192 VSS 0.074916f
C9921 PAD.n11194 VSS 0.074916f
C9922 PAD.n11196 VSS 0.074916f
C9923 PAD.n11198 VSS 0.074916f
C9924 PAD.n11200 VSS 0.074916f
C9925 PAD.n11202 VSS 0.074916f
C9926 PAD.n11204 VSS 0.074916f
C9927 PAD.n11206 VSS 0.074916f
C9928 PAD.n11208 VSS 0.074916f
C9929 PAD.n11210 VSS 0.074916f
C9930 PAD.n11212 VSS 0.074916f
C9931 PAD.n11214 VSS 0.074916f
C9932 PAD.n11216 VSS 0.074916f
C9933 PAD.n11218 VSS 0.074916f
C9934 PAD.n11220 VSS 0.074916f
C9935 PAD.n11222 VSS 0.074916f
C9936 PAD.n11224 VSS 0.074916f
C9937 PAD.n11226 VSS 0.074916f
C9938 PAD.n11228 VSS 0.074916f
C9939 PAD.n11230 VSS 0.074916f
C9940 PAD.n11232 VSS 0.074916f
C9941 PAD.n11234 VSS 0.074916f
C9942 PAD.n11236 VSS 0.074916f
C9943 PAD.n11238 VSS 0.074916f
C9944 PAD.n11240 VSS 0.074916f
C9945 PAD.n11242 VSS 0.074916f
C9946 PAD.n11244 VSS 0.074916f
C9947 PAD.n11246 VSS 0.074916f
C9948 PAD.n11248 VSS 0.074916f
C9949 PAD.n11250 VSS 0.074916f
C9950 PAD.n11252 VSS 0.074916f
C9951 PAD.n11253 VSS 0.044894f
C9952 PAD.n11302 VSS 0.611735f
C9953 PAD.n11303 VSS 0.044894f
C9954 PAD.n11304 VSS 0.074916f
C9955 PAD.n11305 VSS 0.074916f
C9956 PAD.n11306 VSS 0.074916f
C9957 PAD.n11307 VSS 0.074916f
C9958 PAD.n11308 VSS 0.074916f
C9959 PAD.n11309 VSS 0.074916f
C9960 PAD.n11310 VSS 0.074916f
C9961 PAD.n11311 VSS 0.074916f
C9962 PAD.n11312 VSS 0.074916f
C9963 PAD.n11313 VSS 0.074916f
C9964 PAD.n11314 VSS 0.074916f
C9965 PAD.n11315 VSS 0.074916f
C9966 PAD.n11316 VSS 0.074916f
C9967 PAD.n11317 VSS 0.074916f
C9968 PAD.n11318 VSS 0.074916f
C9969 PAD.n11319 VSS 0.074916f
C9970 PAD.n11320 VSS 0.074916f
C9971 PAD.n11321 VSS 0.074916f
C9972 PAD.n11322 VSS 0.074916f
C9973 PAD.n11323 VSS 0.074916f
C9974 PAD.n11324 VSS 0.074916f
C9975 PAD.n11325 VSS 0.074916f
C9976 PAD.n11326 VSS 0.074916f
C9977 PAD.n11327 VSS 0.074916f
C9978 PAD.n11328 VSS 0.074916f
C9979 PAD.n11329 VSS 0.074916f
C9980 PAD.n11330 VSS 0.074916f
C9981 PAD.n11331 VSS 0.074916f
C9982 PAD.n11332 VSS 0.074916f
C9983 PAD.n11333 VSS 0.074916f
C9984 PAD.n11334 VSS 0.074916f
C9985 PAD.n11335 VSS 0.074916f
C9986 PAD.n11336 VSS 0.074916f
C9987 PAD.n11337 VSS 0.074916f
C9988 PAD.n11338 VSS 0.074916f
C9989 PAD.n11339 VSS 0.074916f
C9990 PAD.n11340 VSS 0.074916f
C9991 PAD.n11341 VSS 0.074916f
C9992 PAD.n11342 VSS 0.074916f
C9993 PAD.n11343 VSS 0.074916f
C9994 PAD.n11344 VSS 0.074916f
C9995 PAD.n11345 VSS 0.074916f
C9996 PAD.n11346 VSS 0.074916f
C9997 PAD.n11347 VSS 0.074916f
C9998 PAD.n11348 VSS 0.074916f
C9999 PAD.n11349 VSS 0.074916f
C10000 PAD.n11350 VSS 0.074916f
C10001 PAD.n11351 VSS 0.074916f
C10002 PAD.n11352 VSS 0.103613f
C10003 PAD.n11353 VSS 0.103613f
C10004 PAD.n11354 VSS 0.074916f
C10005 PAD.n11355 VSS 0.074916f
C10006 PAD.n11356 VSS 0.074916f
C10007 PAD.n11357 VSS 0.074916f
C10008 PAD.n11358 VSS 0.074916f
C10009 PAD.n11359 VSS 0.074916f
C10010 PAD.n11360 VSS 0.074916f
C10011 PAD.n11361 VSS 0.074916f
C10012 PAD.n11362 VSS 0.074916f
C10013 PAD.n11363 VSS 0.074916f
C10014 PAD.n11364 VSS 0.074916f
C10015 PAD.n11365 VSS 0.074916f
C10016 PAD.n11366 VSS 0.074916f
C10017 PAD.n11367 VSS 0.074916f
C10018 PAD.n11368 VSS 0.074916f
C10019 PAD.n11369 VSS 0.074916f
C10020 PAD.n11370 VSS 0.074916f
C10021 PAD.n11371 VSS 0.074916f
C10022 PAD.n11372 VSS 0.074916f
C10023 PAD.n11373 VSS 0.074916f
C10024 PAD.n11374 VSS 0.074916f
C10025 PAD.n11375 VSS 0.074916f
C10026 PAD.n11376 VSS 0.074916f
C10027 PAD.n11377 VSS 0.074916f
C10028 PAD.n11378 VSS 0.074916f
C10029 PAD.n11379 VSS 0.074916f
C10030 PAD.n11380 VSS 0.074916f
C10031 PAD.n11381 VSS 0.074916f
C10032 PAD.n11382 VSS 0.074916f
C10033 PAD.n11383 VSS 0.074916f
C10034 PAD.n11384 VSS 0.074916f
C10035 PAD.n11385 VSS 0.074916f
C10036 PAD.n11386 VSS 0.074916f
C10037 PAD.n11387 VSS 0.074916f
C10038 PAD.n11388 VSS 0.074916f
C10039 PAD.n11389 VSS 0.074916f
C10040 PAD.n11390 VSS 0.074916f
C10041 PAD.n11391 VSS 0.074916f
C10042 PAD.n11392 VSS 0.074916f
C10043 PAD.n11393 VSS 0.074916f
C10044 PAD.n11394 VSS 0.074916f
C10045 PAD.n11395 VSS 0.074916f
C10046 PAD.n11396 VSS 0.074916f
C10047 PAD.n11397 VSS 0.074916f
C10048 PAD.n11398 VSS 0.074916f
C10049 PAD.n11399 VSS 0.074916f
C10050 PAD.n11400 VSS 0.074916f
C10051 PAD.n11401 VSS 0.074916f
C10052 PAD.n11402 VSS 0.074916f
C10053 PAD.n11403 VSS 0.074916f
C10054 PAD.n11404 VSS 0.074916f
C10055 PAD.n11405 VSS 0.074916f
C10056 PAD.n11406 VSS 0.074916f
C10057 PAD.n11407 VSS 0.074916f
C10058 PAD.n11408 VSS 0.074916f
C10059 PAD.n11409 VSS 0.074916f
C10060 PAD.n11410 VSS 0.074916f
C10061 PAD.n11411 VSS 0.074916f
C10062 PAD.n11412 VSS 0.074916f
C10063 PAD.n11413 VSS 0.074916f
C10064 PAD.n11414 VSS 0.074916f
C10065 PAD.n11415 VSS 0.074916f
C10066 PAD.n11416 VSS 0.074916f
C10067 PAD.n11417 VSS 0.074916f
C10068 PAD.n11418 VSS 0.074916f
C10069 PAD.n11419 VSS 0.074916f
C10070 PAD.n11420 VSS 0.074916f
C10071 PAD.n11421 VSS 0.074916f
C10072 PAD.n11422 VSS 0.074916f
C10073 PAD.n11423 VSS 0.074916f
C10074 PAD.n11424 VSS 0.074916f
C10075 PAD.n11425 VSS 0.074916f
C10076 PAD.n11426 VSS 0.074916f
C10077 PAD.n11427 VSS 0.074916f
C10078 PAD.n11428 VSS 0.074916f
C10079 PAD.n11429 VSS 0.074916f
C10080 PAD.n11430 VSS 0.074916f
C10081 PAD.n11431 VSS 0.074916f
C10082 PAD.n11432 VSS 0.074916f
C10083 PAD.n11433 VSS 0.074916f
C10084 PAD.n11434 VSS 0.074916f
C10085 PAD.n11435 VSS 0.074916f
C10086 PAD.n11436 VSS 0.074916f
C10087 PAD.n11437 VSS 0.074916f
C10088 PAD.n11438 VSS 0.074916f
C10089 PAD.n11439 VSS 0.074916f
C10090 PAD.n11440 VSS 0.074916f
C10091 PAD.n11441 VSS 0.074916f
C10092 PAD.n11442 VSS 0.074916f
C10093 PAD.n11443 VSS 0.074916f
C10094 PAD.n11444 VSS 0.074916f
C10095 PAD.n11445 VSS 0.074916f
C10096 PAD.n11446 VSS 0.074916f
C10097 PAD.n11447 VSS 0.074916f
C10098 PAD.n11448 VSS 0.074916f
C10099 PAD.n11449 VSS 0.074916f
C10100 PAD.n11450 VSS 0.074916f
C10101 PAD.n11451 VSS 0.074916f
C10102 PAD.n11452 VSS 0.074916f
C10103 PAD.n11453 VSS 0.074916f
C10104 PAD.n11454 VSS 0.074916f
C10105 PAD.n11455 VSS 0.074916f
C10106 PAD.n11456 VSS 0.074916f
C10107 PAD.n11457 VSS 0.074916f
C10108 PAD.n11458 VSS 0.074916f
C10109 PAD.n11459 VSS 0.074916f
C10110 PAD.n11460 VSS 0.074916f
C10111 PAD.n11461 VSS 0.074916f
C10112 PAD.n11462 VSS 0.074916f
C10113 PAD.n11463 VSS 0.074916f
C10114 PAD.n11464 VSS 0.074916f
C10115 PAD.n11465 VSS 0.074916f
C10116 PAD.n11466 VSS 0.074916f
C10117 PAD.n11467 VSS 0.074916f
C10118 PAD.n11468 VSS 0.074916f
C10119 PAD.n11469 VSS 0.074916f
C10120 PAD.n11470 VSS 0.074916f
C10121 PAD.n11471 VSS 0.074916f
C10122 PAD.n11472 VSS 0.074916f
C10123 PAD.n11473 VSS 0.074916f
C10124 PAD.n11474 VSS 0.074916f
C10125 PAD.n11475 VSS 0.074916f
C10126 PAD.n11476 VSS 0.074916f
C10127 PAD.n11477 VSS 0.074916f
C10128 PAD.n11478 VSS 0.074916f
C10129 PAD.n11479 VSS 0.074916f
C10130 PAD.n11480 VSS 0.074916f
C10131 PAD.n11481 VSS 0.074916f
C10132 PAD.n11482 VSS 0.074916f
C10133 PAD.n11483 VSS 0.074916f
C10134 PAD.n11484 VSS 0.074916f
C10135 PAD.n11485 VSS 0.074916f
C10136 PAD.n11486 VSS 0.074916f
C10137 PAD.n11487 VSS 0.074916f
C10138 PAD.n11488 VSS 0.074916f
C10139 PAD.n11489 VSS 0.074916f
C10140 PAD.n11490 VSS 0.074916f
C10141 PAD.n11491 VSS 0.074916f
C10142 PAD.n11492 VSS 0.074916f
C10143 PAD.n11493 VSS 0.074916f
C10144 PAD.n11494 VSS 0.074916f
C10145 PAD.n11495 VSS 0.074916f
C10146 PAD.n11496 VSS 0.074916f
C10147 PAD.n11497 VSS 0.074916f
C10148 PAD.n11498 VSS 0.05951f
C10149 PAD.n11499 VSS 0.06827f
C10150 PAD.n11500 VSS 0.700534f
C10151 PAD.n11501 VSS 0.611734f
C10152 PAD.n11502 VSS 0.031994f
C10153 PAD.n11503 VSS 0.031994f
C10154 PAD.n11504 VSS 0.027942f
C10155 PAD.n11505 VSS 0.157826f
C10156 PAD.n11506 VSS 0.12326f
C10157 PAD.n11507 VSS 0.611735f
C10158 PAD.n11508 VSS 0.122947f
C10159 PAD.n11509 VSS 0.611735f
C10160 PAD.n11510 VSS 0.611735f
C10161 PAD.n11512 VSS 0.126224f
C10162 PAD.n11513 VSS 0.611735f
C10163 PAD.n11514 VSS 0.043197f
C10164 PAD.n11515 VSS 0.043197f
C10165 PAD.n11516 VSS 0.055281f
C10166 PAD.n11517 VSS 0.24295f
C10167 PAD.n11518 VSS 0.060767f
C10168 PAD.n11519 VSS 0.062274f
C10169 PAD.n11520 VSS 0.069765f
C10170 PAD.n11521 VSS 0.069765f
C10171 PAD.n11522 VSS 0.700534f
C10172 PAD.n11523 VSS 0.611734f
C10173 PAD.n11524 VSS 0.043754f
C10174 PAD.n11525 VSS 0.043754f
C10175 PAD.n11526 VSS 0.038213f
C10176 PAD.n11527 VSS 0.033773f
C10177 PAD.n11528 VSS 0.02613f
C10178 PAD.n11529 VSS 0.042895f
C10179 PAD.n11530 VSS 0.049115f
C10180 PAD.n11531 VSS 0.049115f
C10181 PAD.n11532 VSS 0.508134f
C10182 PAD.n11533 VSS 0.626534f
C10183 PAD.n11534 VSS 0.685734f
C10184 PAD.n11535 VSS 0.063014f
C10185 PAD.n11536 VSS 0.063014f
C10186 PAD.n11537 VSS 0.03415f
C10187 PAD.n11538 VSS 1.34014f
C10188 PAD.n11539 VSS 16.0798f
C10189 PAD.n11540 VSS 19.374f
C10190 PAD.n11541 VSS 10.1412f
C10191 PAD.n11542 VSS 0.182456f
C10192 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 VSS 3.15768f
C10193 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS VSS 82.8841f
C10194 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t5 VSS 0.254635f
C10195 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t1 VSS 0.25282f
C10196 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t12 VSS 0.25282f
C10197 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t3 VSS 0.25282f
C10198 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t6 VSS 0.179786f
C10199 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t11 VSS 0.176741f
C10200 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t8 VSS 0.162077f
C10201 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t7 VSS 0.158929f
C10202 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t10 VSS 0.279759f
C10203 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t9 VSS 0.279759f
C10204 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t4 VSS 0.279759f
C10205 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t2 VSS 0.279759f
C10206 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN.t0 VSS 0.048604f
C10207 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 VSS 2.03068f
C10208 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n1 VSS 0.72097f
C10209 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t2 VSS 0.355443f
C10210 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t9 VSS 0.201668f
C10211 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t1 VSS 0.355443f
C10212 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t8 VSS 0.201668f
C10213 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n2 VSS 0.515203f
C10214 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n3 VSS 0.511741f
C10215 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t0 VSS 0.128791f
C10216 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t4 VSS 0.31839f
C10217 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t3 VSS 0.2261f
C10218 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t10 VSS 0.226338f
C10219 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t5 VSS 0.22431f
C10220 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t11 VSS 0.317768f
C10221 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t12 VSS 0.317768f
C10222 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t6 VSS 0.317768f
C10223 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t7 VSS 0.317768f
C10224 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t2 VSS 0.978804f
C10225 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t4 VSS 0.098628f
C10226 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n0 VSS 0.719511f
C10227 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t5 VSS 11.609401f
C10228 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t1 VSS 1.09267f
C10229 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n1 VSS 1.57958f
C10230 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n2 VSS 0.77677f
C10231 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t3 VSS 2.47609f
C10232 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n3 VSS 1.22926f
C10233 GF_NI_BI_T_BASE_0.ndrive_y_<0>.t0 VSS 1.25612f
C10234 GF_NI_BI_T_BASE_0.ndrive_y_<0>.n4 VSS 1.15384f
C10235 GF_NI_BI_T_BASE_0.ndrive_x_<0>.t0 VSS 2.97732f
C10236 GF_NI_BI_T_BASE_0.ndrive_x_<0>.t1 VSS 0.736166f
C10237 GF_NI_BI_T_BASE_0.ndrive_x_<0>.t2 VSS 0.106531f
C10238 GF_NI_BI_T_BASE_0.ndrive_x_<0>.n0 VSS 1.72255f
C10239 GF_NI_BI_T_BASE_0.ndrive_x_<0>.t3 VSS 11.547501f
C10240 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t1 VSS 0.176762f
C10241 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t0 VSS 0.500068f
C10242 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t4 VSS 0.48626f
C10243 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t11 VSS 0.27589f
C10244 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t10 VSS 0.48626f
C10245 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t8 VSS 0.27589f
C10246 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n0 VSS 0.704818f
C10247 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n1 VSS 0.698682f
C10248 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t5 VSS 1.51298f
C10249 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t12 VSS 1.50265f
C10250 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n2 VSS 1.24529f
C10251 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t2 VSS 1.50265f
C10252 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t3 VSS 1.51298f
C10253 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n3 VSS 1.24529f
C10254 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t13 VSS 1.51298f
C10255 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t7 VSS 1.50265f
C10256 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n4 VSS 1.24529f
C10257 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n5 VSS 2.77844f
C10258 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t6 VSS 1.50265f
C10259 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.t9 VSS 1.51298f
C10260 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n6 VSS 1.24529f
C10261 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n7 VSS 2.28053f
C10262 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL.n8 VSS 2.53456f
C10263 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t0 VSS 0.924776f
C10264 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t1 VSS 0.146537f
C10265 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A VSS 0.561385f
C10266 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t3 VSS 0.134163f
C10267 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t2 VSS 0.089926f
C10268 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.n0 VSS 0.143212f
C10269 DVDD.n0 VSS 0.253338f
C10270 DVDD.n1 VSS 0.281047f
C10271 DVDD.n2 VSS 0.281047f
C10272 DVDD.n3 VSS 0.281047f
C10273 DVDD.n4 VSS 0.281047f
C10274 DVDD.n5 VSS 0.281047f
C10275 DVDD.n6 VSS 0.281047f
C10276 DVDD.n7 VSS 0.140524f
C10277 DVDD.n8 VSS 0.023765f
C10278 DVDD.n9 VSS 0.023765f
C10279 DVDD.n10 VSS 0.023765f
C10280 DVDD.n11 VSS 0.023765f
C10281 DVDD.n12 VSS 0.023765f
C10282 DVDD.n13 VSS 0.023765f
C10283 DVDD.n14 VSS 0.023765f
C10284 DVDD.n15 VSS 0.023765f
C10285 DVDD.n16 VSS 0.023765f
C10286 DVDD.n17 VSS 0.023765f
C10287 DVDD.n18 VSS 0.023765f
C10288 DVDD.n19 VSS 0.023765f
C10289 DVDD.n20 VSS 0.023765f
C10290 DVDD.n21 VSS 0.023765f
C10291 DVDD.n22 VSS 0.023765f
C10292 DVDD.n23 VSS 0.023765f
C10293 DVDD.n24 VSS 0.023765f
C10294 DVDD.n25 VSS 0.023765f
C10295 DVDD.n26 VSS 0.023765f
C10296 DVDD.n27 VSS 0.023765f
C10297 DVDD.n28 VSS 0.025004f
C10298 DVDD.n29 VSS 0.140524f
C10299 DVDD.n30 VSS 0.026448f
C10300 DVDD.n31 VSS 0.140524f
C10301 DVDD.n32 VSS 0.167243f
C10302 DVDD.n33 VSS 0.257297f
C10303 DVDD.n34 VSS 0.338444f
C10304 DVDD.n35 VSS 0.536365f
C10305 DVDD.n36 VSS 0.281047f
C10306 DVDD.n37 VSS 0.281047f
C10307 DVDD.n38 VSS 0.536365f
C10308 DVDD.n39 VSS 0.281047f
C10309 DVDD.n40 VSS 0.338444f
C10310 DVDD.n41 VSS 0.338444f
C10311 DVDD.n42 VSS 0.164274f
C10312 DVDD.n43 VSS 0.140524f
C10313 DVDD.n44 VSS 0.536365f
C10314 DVDD.n45 VSS 0.257297f
C10315 DVDD.n46 VSS 0.281047f
C10316 DVDD.n47 VSS 0.281047f
C10317 DVDD.n48 VSS 0.013032f
C10318 DVDD.n49 VSS 0.007282f
C10319 DVDD.n50 VSS 0.023764f
C10320 DVDD.n51 VSS 0.017248f
C10321 DVDD.n52 VSS 0.010349f
C10322 DVDD.n53 VSS 0.003449f
C10323 DVDD.n54 VSS 0.020315f
C10324 DVDD.n55 VSS 0.013415f
C10325 DVDD.n56 VSS 0.006516f
C10326 DVDD.n57 VSS 0.023381f
C10327 DVDD.n58 VSS 0.173181f
C10328 DVDD.n59 VSS 0.019931f
C10329 DVDD.n60 VSS 0.003066f
C10330 DVDD.n61 VSS 0.009965f
C10331 DVDD.n62 VSS 0.016865f
C10332 DVDD.n63 VSS 0.023764f
C10333 DVDD.n64 VSS 0.006899f
C10334 DVDD.n65 VSS 0.013798f
C10335 DVDD.n66 VSS 0.020698f
C10336 DVDD.n67 VSS 0.003832f
C10337 DVDD.n68 VSS 0.010732f
C10338 DVDD.n69 VSS 0.008241f
C10339 DVDD.n70 VSS 0.011691f
C10340 DVDD.n71 VSS 0.026256f
C10341 DVDD.n72 VSS 0.070927f
C10342 DVDD.n73 VSS 0.070927f
C10343 DVDD.n74 VSS 0.023765f
C10344 DVDD.n75 VSS 0.046045f
C10345 DVDD.n76 VSS 0.101929f
C10346 DVDD.n77 VSS 0.101929f
C10347 DVDD.n78 VSS 0.015524f
C10348 DVDD.n79 VSS 0.101929f
C10349 DVDD.n80 VSS 0.167243f
C10350 DVDD.n81 VSS 0.016673f
C10351 DVDD.n82 VSS 0.140524f
C10352 DVDD.n83 VSS 0.027215f
C10353 DVDD.n84 VSS 0.018781f
C10354 DVDD.n85 VSS 0.035463f
C10355 DVDD.n86 VSS 0.060345f
C10356 DVDD.n88 VSS 0.018046f
C10357 DVDD.n89 VSS 0.018174f
C10358 DVDD.n90 VSS 0.015999f
C10359 DVDD.n91 VSS 0.018174f
C10360 DVDD.n92 VSS 0.018174f
C10361 DVDD.n93 VSS 0.018174f
C10362 DVDD.n94 VSS 0.018174f
C10363 DVDD.n95 VSS 0.018174f
C10364 DVDD.n96 VSS 0.018174f
C10365 DVDD.n97 VSS 0.018174f
C10366 DVDD.n98 VSS 0.018046f
C10367 DVDD.n99 VSS 0.018174f
C10368 DVDD.n100 VSS 0.020862f
C10369 DVDD.n102 VSS 0.015871f
C10370 DVDD.n103 VSS 3.89787f
C10371 DVDD.n105 VSS 0.176949f
C10372 DVDD.n107 VSS 0.057397f
C10373 DVDD.n108 VSS 0.090054f
C10374 DVDD.n109 VSS 0.015871f
C10375 DVDD.n110 VSS 0.015871f
C10376 DVDD.n111 VSS 0.015871f
C10377 DVDD.n112 VSS 0.015871f
C10378 DVDD.n113 VSS 0.015871f
C10379 DVDD.n114 VSS 0.015871f
C10380 DVDD.n115 VSS 0.281047f
C10381 DVDD.n116 VSS 0.121721f
C10382 DVDD.n117 VSS 0.281047f
C10383 DVDD.n118 VSS 0.281047f
C10384 DVDD.n119 VSS 0.338444f
C10385 DVDD.n120 VSS 0.281047f
C10386 DVDD.n121 VSS 0.281047f
C10387 DVDD.n122 VSS 0.281047f
C10388 DVDD.n123 VSS 0.281047f
C10389 DVDD.n124 VSS 0.281047f
C10390 DVDD.n125 VSS 0.281047f
C10391 DVDD.n126 VSS 0.281047f
C10392 DVDD.n127 VSS 0.281047f
C10393 DVDD.n128 VSS 0.281047f
C10394 DVDD.n129 VSS 0.281047f
C10395 DVDD.n130 VSS 0.140524f
C10396 DVDD.n131 VSS 0.281047f
C10397 DVDD.n132 VSS 0.281047f
C10398 DVDD.n133 VSS 0.281047f
C10399 DVDD.n134 VSS 0.281047f
C10400 DVDD.n135 VSS 0.017881f
C10401 DVDD.n136 VSS 0.00998f
C10402 DVDD.n137 VSS 0.140524f
C10403 DVDD.n138 VSS 0.00998f
C10404 DVDD.n139 VSS 0.019961f
C10405 DVDD.n140 VSS 0.00998f
C10406 DVDD.n141 VSS 0.019961f
C10407 DVDD.n142 VSS 0.011429f
C10408 DVDD.n143 VSS 0.140524f
C10409 DVDD.n144 VSS 0.140524f
C10410 DVDD.n145 VSS 0.00998f
C10411 DVDD.n146 VSS 0.00998f
C10412 DVDD.n147 VSS 0.00998f
C10413 DVDD.n148 VSS 0.00998f
C10414 DVDD.n149 VSS 0.00998f
C10415 DVDD.n150 VSS 0.00998f
C10416 DVDD.n151 VSS 0.00998f
C10417 DVDD.n152 VSS 0.00998f
C10418 DVDD.n153 VSS 0.00998f
C10419 DVDD.n154 VSS 0.00998f
C10420 DVDD.n155 VSS 0.153388f
C10421 DVDD.n156 VSS 0.00998f
C10422 DVDD.n157 VSS 0.00998f
C10423 DVDD.n158 VSS 0.00998f
C10424 DVDD.n159 VSS 0.00998f
C10425 DVDD.n160 VSS 0.00998f
C10426 DVDD.n161 VSS 0.00998f
C10427 DVDD.n162 VSS 0.00998f
C10428 DVDD.n163 VSS 0.00998f
C10429 DVDD.n164 VSS 0.011429f
C10430 DVDD.n165 VSS -0.294669f
C10431 DVDD.n166 VSS 0.00998f
C10432 DVDD.n167 VSS 0.019961f
C10433 DVDD.n168 VSS 0.011429f
C10434 DVDD.n169 VSS 0.140524f
C10435 DVDD.n170 VSS 0.268182f
C10436 DVDD.n171 VSS 0.00998f
C10437 DVDD.n172 VSS 0.00998f
C10438 DVDD.n173 VSS 0.00998f
C10439 DVDD.n174 VSS 0.00998f
C10440 DVDD.n175 VSS 0.00998f
C10441 DVDD.n176 VSS 0.00998f
C10442 DVDD.n177 VSS 0.00998f
C10443 DVDD.n178 VSS 0.00998f
C10444 DVDD.n179 VSS 0.00998f
C10445 DVDD.n180 VSS 0.140524f
C10446 DVDD.n181 VSS 0.00998f
C10447 DVDD.n182 VSS 0.00998f
C10448 DVDD.n183 VSS 0.00998f
C10449 DVDD.n184 VSS 0.00998f
C10450 DVDD.n185 VSS 0.00998f
C10451 DVDD.n186 VSS 0.00998f
C10452 DVDD.n187 VSS 0.00998f
C10453 DVDD.n188 VSS 0.00998f
C10454 DVDD.n189 VSS 0.00998f
C10455 DVDD.n190 VSS 0.011429f
C10456 DVDD.n191 VSS 0.010624f
C10457 DVDD.n192 VSS 0.019961f
C10458 DVDD.n193 VSS 0.00998f
C10459 DVDD.n194 VSS 0.019961f
C10460 DVDD.n195 VSS 0.011429f
C10461 DVDD.n196 VSS 0.140524f
C10462 DVDD.n197 VSS 0.140524f
C10463 DVDD.n198 VSS 0.017326f
C10464 DVDD.n199 VSS 0.281047f
C10465 DVDD.n200 VSS 0.281047f
C10466 DVDD.n201 VSS 0.281047f
C10467 DVDD.n202 VSS 0.281047f
C10468 DVDD.n203 VSS 0.281047f
C10469 DVDD.n204 VSS 0.281047f
C10470 DVDD.n205 VSS 0.281047f
C10471 DVDD.n206 VSS 0.281047f
C10472 DVDD.n207 VSS 0.281047f
C10473 DVDD.n208 VSS 0.281047f
C10474 DVDD.n209 VSS 0.281047f
C10475 DVDD.n210 VSS 0.281047f
C10476 DVDD.n211 VSS 0.281047f
C10477 DVDD.n212 VSS 0.281047f
C10478 DVDD.n213 VSS 0.281047f
C10479 DVDD.n214 VSS 0.281047f
C10480 DVDD.n215 VSS 0.164274f
C10481 DVDD.n216 VSS 0.257297f
C10482 DVDD.n217 VSS 0.281047f
C10483 DVDD.n218 VSS 0.023764f
C10484 DVDD.n219 VSS 0.023764f
C10485 DVDD.n220 VSS 0.140524f
C10486 DVDD.n221 VSS 0.023764f
C10487 DVDD.n222 VSS 0.023764f
C10488 DVDD.n223 VSS 0.141142f
C10489 DVDD.n224 VSS 0.101929f
C10490 DVDD.n225 VSS 0.027214f
C10491 DVDD.n226 VSS 0.101929f
C10492 DVDD.n227 VSS 0.121721f
C10493 DVDD.n228 VSS 0.02675f
C10494 DVDD.n229 VSS 0.015871f
C10495 DVDD.n230 VSS 0.015871f
C10496 DVDD.n231 VSS 0.015871f
C10497 DVDD.n232 VSS 0.015871f
C10498 DVDD.n233 VSS 0.015871f
C10499 DVDD.n234 VSS 0.179118f
C10500 DVDD.n235 VSS 0.022142f
C10501 DVDD.n236 VSS 0.015871f
C10502 DVDD.n237 VSS 0.015871f
C10503 DVDD.n238 VSS 0.015871f
C10504 DVDD.n239 VSS 0.015871f
C10505 DVDD.n240 VSS 0.018174f
C10506 DVDD.n241 VSS 0.057397f
C10507 DVDD.n242 VSS 0.018046f
C10508 DVDD.n243 VSS 0.06111f
C10509 DVDD.n244 VSS 0.018174f
C10510 DVDD.n245 VSS 0.108697f
C10511 DVDD.n246 VSS 0.018174f
C10512 DVDD.n247 VSS 0.06111f
C10513 DVDD.n248 VSS 0.06111f
C10514 DVDD.n249 VSS 0.015999f
C10515 DVDD.n250 VSS 0.018046f
C10516 DVDD.n251 VSS 0.06111f
C10517 DVDD.n252 VSS 0.018174f
C10518 DVDD.n253 VSS 0.06111f
C10519 DVDD.n254 VSS 0.018174f
C10520 DVDD.n255 VSS 0.045832f
C10521 DVDD.n256 VSS 0.537986f
C10522 DVDD.n257 VSS 0.018174f
C10523 DVDD.n258 VSS 0.19988f
C10524 DVDD.n259 VSS 1.2609f
C10525 DVDD.t82 VSS 4.6783f
C10526 DVDD.n260 VSS 8.45063f
C10527 DVDD.n261 VSS 0.855461f
C10528 DVDD.t88 VSS 4.72285f
C10529 DVDD.n262 VSS 0.885587f
C10530 DVDD.t179 VSS 4.6783f
C10531 DVDD.n263 VSS 1.25662f
C10532 DVDD.n264 VSS 0.030269f
C10533 DVDD.n265 VSS 0.065912f
C10534 DVDD.n266 VSS -0.17236f
C10535 DVDD.n267 VSS 0.023765f
C10536 DVDD.n268 VSS 0.01399f
C10537 DVDD.n269 VSS 0.070763f
C10538 DVDD.n270 VSS 0.010732f
C10539 DVDD.n271 VSS 0.140524f
C10540 DVDD.n272 VSS 0.007282f
C10541 DVDD.n273 VSS 0.140524f
C10542 DVDD.n274 VSS 0.026256f
C10543 DVDD.n275 VSS 0.02089f
C10544 DVDD.n276 VSS 0.004024f
C10545 DVDD.n277 VSS 0.010924f
C10546 DVDD.n278 VSS 0.017823f
C10547 DVDD.n279 VSS 0.003258f
C10548 DVDD.n280 VSS 0.007857f
C10549 DVDD.n281 VSS 0.014757f
C10550 DVDD.n282 VSS 0.021657f
C10551 DVDD.n283 VSS 0.004791f
C10552 DVDD.n284 VSS 0.173181f
C10553 DVDD.n285 VSS 0.008241f
C10554 DVDD.n286 VSS 0.001341f
C10555 DVDD.n287 VSS 0.018207f
C10556 DVDD.n288 VSS 0.011307f
C10557 DVDD.n289 VSS 0.004408f
C10558 DVDD.n290 VSS 0.021273f
C10559 DVDD.n291 VSS 0.014374f
C10560 DVDD.n292 VSS 0.007474f
C10561 DVDD.n293 VSS 0.023765f
C10562 DVDD.n294 VSS 0.026256f
C10563 DVDD.n295 VSS 0.140524f
C10564 DVDD.n296 VSS 0.026211f
C10565 DVDD.n297 VSS 0.140524f
C10566 DVDD.n298 VSS 0.003832f
C10567 DVDD.n299 VSS 0.020698f
C10568 DVDD.n300 VSS 0.013798f
C10569 DVDD.n301 VSS 0.006899f
C10570 DVDD.n302 VSS 0.023764f
C10571 DVDD.n303 VSS 0.016865f
C10572 DVDD.n304 VSS 0.009965f
C10573 DVDD.n305 VSS 0.003066f
C10574 DVDD.n306 VSS 0.019931f
C10575 DVDD.n307 VSS 0.095991f
C10576 DVDD.n308 VSS 0.016482f
C10577 DVDD.n309 VSS 0.023381f
C10578 DVDD.n310 VSS 0.006516f
C10579 DVDD.n311 VSS 0.013415f
C10580 DVDD.n312 VSS 0.020315f
C10581 DVDD.n313 VSS 0.003449f
C10582 DVDD.n314 VSS 0.010349f
C10583 DVDD.n315 VSS 0.017248f
C10584 DVDD.n316 VSS 9.58e-19
C10585 DVDD.n317 VSS 0.026256f
C10586 DVDD.n318 VSS 0.070763f
C10587 DVDD.n319 VSS 0.070763f
C10588 DVDD.n320 VSS 0.070763f
C10589 DVDD.n321 VSS 0.091044f
C10590 DVDD.n322 VSS 0.140524f
C10591 DVDD.n323 VSS 0.027215f
C10592 DVDD.n324 VSS 0.091044f
C10593 DVDD.n325 VSS 0.059376f
C10594 DVDD.n326 VSS 0.023765f
C10595 DVDD.n327 VSS 0.05901f
C10596 DVDD.n328 VSS 0.130628f
C10597 DVDD.n329 VSS 0.018781f
C10598 DVDD.n330 VSS 0.070763f
C10599 DVDD.n331 VSS 0.015524f
C10600 DVDD.n332 VSS 0.045939f
C10601 DVDD.n333 VSS 0.035381f
C10602 DVDD.n334 VSS 0.018046f
C10603 DVDD.n335 VSS 0.018174f
C10604 DVDD.n336 VSS 0.018174f
C10605 DVDD.n337 VSS 0.018046f
C10606 DVDD.n338 VSS 0.018174f
C10607 DVDD.n339 VSS 0.020862f
C10608 DVDD.n341 VSS 0.020862f
C10609 DVDD.n342 VSS 0.018174f
C10610 DVDD.n343 VSS 0.018174f
C10611 DVDD.n344 VSS 0.015999f
C10612 DVDD.n345 VSS 0.018174f
C10613 DVDD.n346 VSS 0.018174f
C10614 DVDD.n347 VSS 0.018174f
C10615 DVDD.n349 VSS 0.015871f
C10616 DVDD.n350 VSS 0.176949f
C10617 DVDD.n352 VSS 0.015871f
C10618 DVDD.n353 VSS 0.059376f
C10619 DVDD.n354 VSS 0.281047f
C10620 DVDD.n355 VSS 0.281047f
C10621 DVDD.n356 VSS 0.281047f
C10622 DVDD.n357 VSS 0.188025f
C10623 DVDD.n358 VSS 0.338444f
C10624 DVDD.n359 VSS 0.536365f
C10625 DVDD.n360 VSS 0.281047f
C10626 DVDD.n361 VSS 0.233546f
C10627 DVDD.n362 VSS 0.281047f
C10628 DVDD.n363 VSS 0.281047f
C10629 DVDD.n364 VSS 0.281047f
C10630 DVDD.n365 VSS 0.281047f
C10631 DVDD.n366 VSS 0.281047f
C10632 DVDD.n367 VSS 0.281047f
C10633 DVDD.n368 VSS 0.281047f
C10634 DVDD.n369 VSS 0.281047f
C10635 DVDD.n370 VSS 0.281047f
C10636 DVDD.n371 VSS 0.281047f
C10637 DVDD.n372 VSS 0.281047f
C10638 DVDD.n373 VSS 0.281047f
C10639 DVDD.n374 VSS 0.281047f
C10640 DVDD.n375 VSS 0.281047f
C10641 DVDD.n376 VSS 0.281047f
C10642 DVDD.n377 VSS 0.017881f
C10643 DVDD.n378 VSS 0.00998f
C10644 DVDD.n379 VSS 0.140524f
C10645 DVDD.n380 VSS 0.00998f
C10646 DVDD.n381 VSS 0.005232f
C10647 DVDD.n382 VSS 0.281047f
C10648 DVDD.n383 VSS 0.281047f
C10649 DVDD.n384 VSS 0.281047f
C10650 DVDD.n385 VSS 0.281047f
C10651 DVDD.n386 VSS 0.281047f
C10652 DVDD.n387 VSS 0.281047f
C10653 DVDD.n388 VSS 0.281047f
C10654 DVDD.n389 VSS 0.281047f
C10655 DVDD.n390 VSS 0.281047f
C10656 DVDD.n391 VSS 0.281047f
C10657 DVDD.n392 VSS 0.281047f
C10658 DVDD.n393 VSS 0.281047f
C10659 DVDD.n394 VSS 0.281047f
C10660 DVDD.n395 VSS 0.281047f
C10661 DVDD.n396 VSS 0.281047f
C10662 DVDD.n397 VSS 0.281047f
C10663 DVDD.n398 VSS 0.281047f
C10664 DVDD.n399 VSS 0.180108f
C10665 DVDD.n400 VSS 0.017881f
C10666 DVDD.n401 VSS 0.00998f
C10667 DVDD.n402 VSS 0.101929f
C10668 DVDD.n403 VSS 0.00998f
C10669 DVDD.n404 VSS 0.005232f
C10670 DVDD.n405 VSS 0.276099f
C10671 DVDD.n406 VSS 0.281047f
C10672 DVDD.n407 VSS 0.338444f
C10673 DVDD.n408 VSS 0.241463f
C10674 DVDD.n409 VSS 0.281047f
C10675 DVDD.n410 VSS 0.281047f
C10676 DVDD.n411 VSS 0.281047f
C10677 DVDD.n412 VSS 0.281047f
C10678 DVDD.n413 VSS 0.281047f
C10679 DVDD.n414 VSS 0.281047f
C10680 DVDD.n415 VSS 0.281047f
C10681 DVDD.n416 VSS 0.281047f
C10682 DVDD.n417 VSS 0.281047f
C10683 DVDD.n418 VSS 0.281047f
C10684 DVDD.n419 VSS 0.281047f
C10685 DVDD.n420 VSS 0.281047f
C10686 DVDD.n421 VSS 0.281047f
C10687 DVDD.n422 VSS 0.281047f
C10688 DVDD.n423 VSS 0.281047f
C10689 DVDD.n424 VSS 0.017881f
C10690 DVDD.n425 VSS 0.00998f
C10691 DVDD.n426 VSS 0.140524f
C10692 DVDD.n427 VSS 0.00998f
C10693 DVDD.n428 VSS 0.005232f
C10694 DVDD.n429 VSS 0.281047f
C10695 DVDD.n430 VSS 0.281047f
C10696 DVDD.n431 VSS 0.281047f
C10697 DVDD.n432 VSS 0.281047f
C10698 DVDD.n433 VSS 0.281047f
C10699 DVDD.n434 VSS 0.281047f
C10700 DVDD.n435 VSS 0.281047f
C10701 DVDD.n436 VSS 0.281047f
C10702 DVDD.n437 VSS 0.281047f
C10703 DVDD.n438 VSS 0.281047f
C10704 DVDD.n439 VSS 0.281047f
C10705 DVDD.n440 VSS 0.281047f
C10706 DVDD.n441 VSS 0.281047f
C10707 DVDD.n442 VSS 0.281047f
C10708 DVDD.n443 VSS 0.281047f
C10709 DVDD.n444 VSS 0.281047f
C10710 DVDD.n445 VSS 0.281047f
C10711 DVDD.n446 VSS 0.281047f
C10712 DVDD.n447 VSS 0.172191f
C10713 DVDD.n448 VSS 0.338444f
C10714 DVDD.n449 VSS 0.108856f
C10715 DVDD.n450 VSS 0.460165f
C10716 DVDD.n451 VSS 0.172191f
C10717 DVDD.n452 VSS 0.00998f
C10718 DVDD.n453 VSS 0.00998f
C10719 DVDD.n454 VSS 0.00998f
C10720 DVDD.n455 VSS 0.00998f
C10721 DVDD.n456 VSS 0.00998f
C10722 DVDD.n457 VSS 0.00998f
C10723 DVDD.n458 VSS 0.00998f
C10724 DVDD.n459 VSS 0.00998f
C10725 DVDD.n460 VSS 0.00998f
C10726 DVDD.n461 VSS 0.00998f
C10727 DVDD.n462 VSS 0.140524f
C10728 DVDD.n463 VSS 0.00998f
C10729 DVDD.n464 VSS 0.00998f
C10730 DVDD.n465 VSS 0.00998f
C10731 DVDD.n466 VSS 0.00998f
C10732 DVDD.n467 VSS 0.00998f
C10733 DVDD.n468 VSS 0.00998f
C10734 DVDD.n469 VSS 0.00998f
C10735 DVDD.n470 VSS 0.00998f
C10736 DVDD.n471 VSS 0.00998f
C10737 DVDD.n472 VSS 0.00998f
C10738 DVDD.n473 VSS 0.011429f
C10739 DVDD.n474 VSS 0.011429f
C10740 DVDD.n475 VSS 0.281047f
C10741 DVDD.n476 VSS 0.24938f
C10742 DVDD.n477 VSS 0.536365f
C10743 DVDD.n478 VSS 0.338444f
C10744 DVDD.n479 VSS 0.281047f
C10745 DVDD.n480 VSS 0.281047f
C10746 DVDD.n481 VSS 0.338444f
C10747 DVDD.n482 VSS 0.172191f
C10748 DVDD.n483 VSS 0.24938f
C10749 DVDD.n484 VSS 0.281047f
C10750 DVDD.n485 VSS 0.108856f
C10751 DVDD.n486 VSS 0.00998f
C10752 DVDD.n487 VSS 0.00998f
C10753 DVDD.n488 VSS 0.00998f
C10754 DVDD.n489 VSS 0.00998f
C10755 DVDD.n490 VSS 0.00998f
C10756 DVDD.n491 VSS 0.00998f
C10757 DVDD.n492 VSS 0.00998f
C10758 DVDD.n493 VSS 0.00998f
C10759 DVDD.n494 VSS 0.00998f
C10760 DVDD.n495 VSS 0.00998f
C10761 DVDD.n496 VSS 0.281047f
C10762 DVDD.n497 VSS 0.281047f
C10763 DVDD.n498 VSS 0.281047f
C10764 DVDD.n499 VSS 0.281047f
C10765 DVDD.n500 VSS 0.281047f
C10766 DVDD.n501 VSS 0.281047f
C10767 DVDD.n502 VSS 0.281047f
C10768 DVDD.n503 VSS 0.281047f
C10769 DVDD.n504 VSS 0.281047f
C10770 DVDD.n505 VSS 0.281047f
C10771 DVDD.n506 VSS 0.281047f
C10772 DVDD.n507 VSS 0.281047f
C10773 DVDD.n508 VSS 0.281047f
C10774 DVDD.n509 VSS 0.281047f
C10775 DVDD.n510 VSS 0.281047f
C10776 DVDD.n511 VSS 0.281047f
C10777 DVDD.n512 VSS 0.281047f
C10778 DVDD.n513 VSS 0.281047f
C10779 DVDD.n514 VSS 0.281047f
C10780 DVDD.n515 VSS 0.281047f
C10781 DVDD.n516 VSS 0.281047f
C10782 DVDD.n517 VSS 0.281047f
C10783 DVDD.n518 VSS 0.281047f
C10784 DVDD.n519 VSS 0.281047f
C10785 DVDD.n520 VSS 0.281047f
C10786 DVDD.n521 VSS 0.281047f
C10787 DVDD.n522 VSS 0.281047f
C10788 DVDD.n523 VSS 0.281047f
C10789 DVDD.n524 VSS 0.281047f
C10790 DVDD.n525 VSS 0.281047f
C10791 DVDD.n526 VSS 0.281047f
C10792 DVDD.n527 VSS 0.281047f
C10793 DVDD.n528 VSS 0.281047f
C10794 DVDD.n529 VSS 0.281047f
C10795 DVDD.n530 VSS 0.281047f
C10796 DVDD.n531 VSS 0.281047f
C10797 DVDD.n532 VSS 0.281047f
C10798 DVDD.n533 VSS 0.281047f
C10799 DVDD.n534 VSS 0.281047f
C10800 DVDD.n535 VSS 0.281047f
C10801 DVDD.n536 VSS 0.281047f
C10802 DVDD.n537 VSS 0.153388f
C10803 DVDD.n538 VSS 0.281047f
C10804 DVDD.n539 VSS 0.281047f
C10805 DVDD.n540 VSS 0.281047f
C10806 DVDD.n541 VSS 0.281047f
C10807 DVDD.n542 VSS 0.281047f
C10808 DVDD.n543 VSS 0.281047f
C10809 DVDD.n544 VSS 0.281047f
C10810 DVDD.n545 VSS 0.281047f
C10811 DVDD.n546 VSS 0.281047f
C10812 DVDD.n547 VSS 0.281047f
C10813 DVDD.n548 VSS 0.281047f
C10814 DVDD.n549 VSS 0.281047f
C10815 DVDD.n550 VSS 0.281047f
C10816 DVDD.n551 VSS 0.281047f
C10817 DVDD.n552 VSS 0.281047f
C10818 DVDD.n553 VSS 0.281047f
C10819 DVDD.n554 VSS 0.281047f
C10820 DVDD.n555 VSS 0.216723f
C10821 DVDD.n556 VSS 0.00998f
C10822 DVDD.n557 VSS 0.00998f
C10823 DVDD.n558 VSS 0.00998f
C10824 DVDD.n559 VSS 0.00998f
C10825 DVDD.n560 VSS 0.00998f
C10826 DVDD.n561 VSS 0.00998f
C10827 DVDD.n562 VSS 0.00998f
C10828 DVDD.n563 VSS 0.00998f
C10829 DVDD.n564 VSS 0.00998f
C10830 DVDD.n565 VSS 0.00998f
C10831 DVDD.n566 VSS 0.018834f
C10832 DVDD.n567 VSS 0.010302f
C10833 DVDD.n568 VSS 0.019961f
C10834 DVDD.n569 VSS 0.011429f
C10835 DVDD.n570 VSS 0.140524f
C10836 DVDD.n571 VSS 0.262245f
C10837 DVDD.n572 VSS 0.027607f
C10838 DVDD.n573 VSS 0.00998f
C10839 DVDD.n574 VSS 0.281047f
C10840 DVDD.n575 VSS 0.281047f
C10841 DVDD.n576 VSS 0.281047f
C10842 DVDD.n577 VSS 0.281047f
C10843 DVDD.n578 VSS 0.281047f
C10844 DVDD.n579 VSS 0.281047f
C10845 DVDD.n580 VSS 0.281047f
C10846 DVDD.n581 VSS 0.281047f
C10847 DVDD.n582 VSS 0.281047f
C10848 DVDD.n583 VSS 0.281047f
C10849 DVDD.n584 VSS 0.140524f
C10850 DVDD.n585 VSS 0.281047f
C10851 DVDD.n586 VSS 0.281047f
C10852 DVDD.n587 VSS 0.281047f
C10853 DVDD.n588 VSS 0.281047f
C10854 DVDD.n589 VSS 0.027607f
C10855 DVDD.n590 VSS 0.00998f
C10856 DVDD.n591 VSS 0.140524f
C10857 DVDD.n592 VSS 0.00998f
C10858 DVDD.n593 VSS 0.017326f
C10859 DVDD.n594 VSS 0.011429f
C10860 DVDD.n595 VSS 0.019961f
C10861 DVDD.n596 VSS 0.00586f
C10862 DVDD.n597 VSS 0.011429f
C10863 DVDD.n598 VSS 0.063742f
C10864 DVDD.n599 VSS 0.011429f
C10865 DVDD.n600 VSS 0.019961f
C10866 DVDD.n601 VSS 0.019961f
C10867 DVDD.n602 VSS 0.019961f
C10868 DVDD.n603 VSS 0.140524f
C10869 DVDD.n604 VSS 0.011107f
C10870 DVDD.n605 VSS 0.141513f
C10871 DVDD.n606 VSS 0.00998f
C10872 DVDD.n607 VSS 0.00998f
C10873 DVDD.n608 VSS 0.00998f
C10874 DVDD.n609 VSS 0.00998f
C10875 DVDD.n610 VSS 0.00998f
C10876 DVDD.n611 VSS 0.00998f
C10877 DVDD.n612 VSS 0.00998f
C10878 DVDD.n613 VSS 0.00998f
C10879 DVDD.n614 VSS 0.00998f
C10880 DVDD.n615 VSS 0.00998f
C10881 DVDD.n616 VSS 0.140524f
C10882 DVDD.n617 VSS 0.00998f
C10883 DVDD.n618 VSS 0.00998f
C10884 DVDD.n619 VSS 0.00998f
C10885 DVDD.n620 VSS 0.00998f
C10886 DVDD.n621 VSS 0.00998f
C10887 DVDD.n622 VSS 0.00998f
C10888 DVDD.n623 VSS 0.00998f
C10889 DVDD.n624 VSS 0.00998f
C10890 DVDD.n625 VSS 0.00998f
C10891 DVDD.n626 VSS 0.011429f
C10892 DVDD.n627 VSS 0.019961f
C10893 DVDD.n628 VSS 0.010302f
C10894 DVDD.n629 VSS 0.019961f
C10895 DVDD.n630 VSS 0.011429f
C10896 DVDD.n631 VSS 0.019961f
C10897 DVDD.n632 VSS 0.011429f
C10898 DVDD.n633 VSS 0.019961f
C10899 DVDD.n634 VSS 0.011429f
C10900 DVDD.n635 VSS 0.019961f
C10901 DVDD.n636 VSS 0.011429f
C10902 DVDD.n637 VSS 0.019961f
C10903 DVDD.n638 VSS 0.011429f
C10904 DVDD.n639 VSS 0.019961f
C10905 DVDD.n640 VSS 0.011429f
C10906 DVDD.n641 VSS 0.019961f
C10907 DVDD.n642 VSS 0.019961f
C10908 DVDD.n643 VSS 0.010946f
C10909 DVDD.n644 VSS 0.010463f
C10910 DVDD.n645 VSS 0.019961f
C10911 DVDD.n646 VSS 0.011429f
C10912 DVDD.n647 VSS 0.019961f
C10913 DVDD.n648 VSS 0.011429f
C10914 DVDD.n649 VSS 0.019961f
C10915 DVDD.n650 VSS 0.011429f
C10916 DVDD.n651 VSS 0.019961f
C10917 DVDD.n652 VSS 0.011429f
C10918 DVDD.n653 VSS 0.019961f
C10919 DVDD.n654 VSS 0.011429f
C10920 DVDD.n655 VSS 0.019961f
C10921 DVDD.n656 VSS 0.011429f
C10922 DVDD.n657 VSS 0.019961f
C10923 DVDD.n658 VSS 0.019961f
C10924 DVDD.n659 VSS 0.010785f
C10925 DVDD.n660 VSS 0.010624f
C10926 DVDD.n661 VSS 0.019961f
C10927 DVDD.n662 VSS 0.011429f
C10928 DVDD.n663 VSS 0.019961f
C10929 DVDD.n664 VSS 0.011429f
C10930 DVDD.n665 VSS 0.019961f
C10931 DVDD.n666 VSS 0.011429f
C10932 DVDD.n667 VSS 0.019961f
C10933 DVDD.n668 VSS 0.011429f
C10934 DVDD.n669 VSS 0.019961f
C10935 DVDD.n670 VSS 0.019961f
C10936 DVDD.n671 VSS 0.019961f
C10937 DVDD.n672 VSS 0.140524f
C10938 DVDD.n673 VSS 0.011429f
C10939 DVDD.n674 VSS 0.141513f
C10940 DVDD.n675 VSS 0.00998f
C10941 DVDD.n676 VSS 0.00998f
C10942 DVDD.n677 VSS 0.00998f
C10943 DVDD.n678 VSS 0.00998f
C10944 DVDD.n679 VSS 0.00998f
C10945 DVDD.n680 VSS 0.00998f
C10946 DVDD.n681 VSS 0.00998f
C10947 DVDD.n682 VSS 0.00998f
C10948 DVDD.n683 VSS 0.00998f
C10949 DVDD.n684 VSS 0.281047f
C10950 DVDD.n685 VSS 0.281047f
C10951 DVDD.n686 VSS 0.281047f
C10952 DVDD.n687 VSS 0.281047f
C10953 DVDD.n688 VSS 0.281047f
C10954 DVDD.n689 VSS 0.281047f
C10955 DVDD.n690 VSS 0.281047f
C10956 DVDD.n691 VSS 0.281047f
C10957 DVDD.n692 VSS 0.281047f
C10958 DVDD.n693 VSS 0.281047f
C10959 DVDD.n694 VSS 0.281047f
C10960 DVDD.n695 VSS 0.10094f
C10961 DVDD.n696 VSS 0.536365f
C10962 DVDD.n697 VSS 0.536365f
C10963 DVDD.n698 VSS 0.180108f
C10964 DVDD.n699 VSS 0.338444f
C10965 DVDD.n700 VSS 0.281047f
C10966 DVDD.n701 VSS 0.281047f
C10967 DVDD.n702 VSS 0.140524f
C10968 DVDD.n703 VSS 0.276099f
C10969 DVDD.n704 VSS 0.101929f
C10970 DVDD.n705 VSS 0.00998f
C10971 DVDD.n706 VSS 0.00998f
C10972 DVDD.n707 VSS 0.00998f
C10973 DVDD.n708 VSS 0.00998f
C10974 DVDD.n709 VSS 0.00998f
C10975 DVDD.n710 VSS 0.00998f
C10976 DVDD.n711 VSS 0.00998f
C10977 DVDD.n712 VSS 0.00998f
C10978 DVDD.n713 VSS 0.00998f
C10979 DVDD.n714 VSS 0.00998f
C10980 DVDD.n715 VSS 0.202869f
C10981 DVDD.n716 VSS 0.00998f
C10982 DVDD.n717 VSS 0.00998f
C10983 DVDD.n718 VSS 0.00998f
C10984 DVDD.n719 VSS 0.00998f
C10985 DVDD.n720 VSS 0.00998f
C10986 DVDD.n721 VSS 0.00998f
C10987 DVDD.n722 VSS 0.00998f
C10988 DVDD.n723 VSS 0.00998f
C10989 DVDD.n724 VSS 0.00998f
C10990 DVDD.n725 VSS 0.00998f
C10991 DVDD.n726 VSS 0.018834f
C10992 DVDD.n727 VSS 0.011107f
C10993 DVDD.n728 VSS 0.281047f
C10994 DVDD.n729 VSS 0.281047f
C10995 DVDD.n730 VSS 0.281047f
C10996 DVDD.n731 VSS 0.180108f
C10997 DVDD.n732 VSS 0.180108f
C10998 DVDD.n733 VSS 0.241463f
C10999 DVDD.n734 VSS 0.281047f
C11000 DVDD.n735 VSS 0.017326f
C11001 DVDD.n736 VSS 0.00998f
C11002 DVDD.n737 VSS 0.00998f
C11003 DVDD.n738 VSS 0.00998f
C11004 DVDD.n739 VSS -0.294669f
C11005 DVDD.n740 VSS 0.00998f
C11006 DVDD.n741 VSS 0.019961f
C11007 DVDD.n742 VSS 0.010222f
C11008 DVDD.n743 VSS 0.019961f
C11009 DVDD.n744 VSS 0.00998f
C11010 DVDD.n745 VSS 0.00998f
C11011 DVDD.n746 VSS 0.019961f
C11012 DVDD.n747 VSS 0.00998f
C11013 DVDD.n748 VSS 0.019961f
C11014 DVDD.n749 VSS 0.00998f
C11015 DVDD.n750 VSS 0.019961f
C11016 DVDD.n751 VSS 0.00998f
C11017 DVDD.n752 VSS 0.019961f
C11018 DVDD.n753 VSS 0.010544f
C11019 DVDD.n754 VSS 0.019961f
C11020 DVDD.n755 VSS 0.00998f
C11021 DVDD.n756 VSS 0.00998f
C11022 DVDD.n757 VSS 0.019961f
C11023 DVDD.n758 VSS 0.011429f
C11024 DVDD.n759 VSS 0.061904f
C11025 DVDD.n760 VSS 0.011429f
C11026 DVDD.n761 VSS 0.019961f
C11027 DVDD.n762 VSS 0.019961f
C11028 DVDD.n763 VSS 0.014971f
C11029 DVDD.n764 VSS 0.019961f
C11030 DVDD.n765 VSS 0.015051f
C11031 DVDD.n766 VSS 0.019961f
C11032 DVDD.n767 VSS 0.019961f
C11033 DVDD.n768 VSS 0.011429f
C11034 DVDD.n769 VSS 0.00998f
C11035 DVDD.n770 VSS 0.011429f
C11036 DVDD.n771 VSS 0.00998f
C11037 DVDD.n772 VSS 0.011429f
C11038 DVDD.n773 VSS 0.019961f
C11039 DVDD.n774 VSS 0.019961f
C11040 DVDD.n775 VSS 0.019961f
C11041 DVDD.n776 VSS 0.010866f
C11042 DVDD.n777 VSS 0.00998f
C11043 DVDD.n778 VSS 0.011429f
C11044 DVDD.n779 VSS 0.00998f
C11045 DVDD.n780 VSS 0.011429f
C11046 DVDD.n781 VSS 0.019961f
C11047 DVDD.n782 VSS 0.019961f
C11048 DVDD.n783 VSS 0.011429f
C11049 DVDD.n784 VSS 0.00998f
C11050 DVDD.n785 VSS 0.011429f
C11051 DVDD.n786 VSS 0.00998f
C11052 DVDD.n787 VSS 0.011429f
C11053 DVDD.n788 VSS 0.019961f
C11054 DVDD.n789 VSS 0.019961f
C11055 DVDD.n790 VSS 0.011429f
C11056 DVDD.n791 VSS 0.00998f
C11057 DVDD.n792 VSS 0.010383f
C11058 DVDD.n793 VSS 0.011027f
C11059 DVDD.n794 VSS 0.019961f
C11060 DVDD.n795 VSS 0.019961f
C11061 DVDD.n796 VSS 0.011429f
C11062 DVDD.n797 VSS 0.00998f
C11063 DVDD.n798 VSS 0.011429f
C11064 DVDD.n799 VSS 0.00998f
C11065 DVDD.n800 VSS 0.011429f
C11066 DVDD.n801 VSS 0.019961f
C11067 DVDD.n802 VSS 0.019961f
C11068 DVDD.n803 VSS 0.011429f
C11069 DVDD.n804 VSS 0.00998f
C11070 DVDD.n805 VSS 0.011429f
C11071 DVDD.n806 VSS 0.00998f
C11072 DVDD.n807 VSS 0.011429f
C11073 DVDD.n808 VSS 0.019961f
C11074 DVDD.n809 VSS 0.019961f
C11075 DVDD.n810 VSS 0.019961f
C11076 DVDD.n811 VSS 0.011188f
C11077 DVDD.n812 VSS 0.00998f
C11078 DVDD.n813 VSS 0.011429f
C11079 DVDD.n814 VSS 0.00998f
C11080 DVDD.n815 VSS 0.011429f
C11081 DVDD.n816 VSS 0.019961f
C11082 DVDD.n817 VSS 0.019961f
C11083 DVDD.n818 VSS 0.015856f
C11084 DVDD.n819 VSS 0.019961f
C11085 DVDD.n820 VSS 0.012073f
C11086 DVDD.n821 VSS -0.36209f
C11087 DVDD.n822 VSS 0.011429f
C11088 DVDD.n823 VSS 0.019961f
C11089 DVDD.n824 VSS 0.011429f
C11090 DVDD.n825 VSS 0.019961f
C11091 DVDD.n826 VSS 0.011429f
C11092 DVDD.n827 VSS 0.019961f
C11093 DVDD.n828 VSS 0.011429f
C11094 DVDD.n829 VSS 0.019961f
C11095 DVDD.n830 VSS 0.011429f
C11096 DVDD.n831 VSS 0.019961f
C11097 DVDD.n832 VSS 0.019961f
C11098 DVDD.n833 VSS 0.010624f
C11099 DVDD.n834 VSS 0.010785f
C11100 DVDD.n835 VSS 0.019961f
C11101 DVDD.n836 VSS 0.011429f
C11102 DVDD.n837 VSS 0.019961f
C11103 DVDD.n838 VSS 0.011429f
C11104 DVDD.n839 VSS 0.019961f
C11105 DVDD.n840 VSS 0.011429f
C11106 DVDD.n841 VSS 0.019961f
C11107 DVDD.n842 VSS 0.011429f
C11108 DVDD.n843 VSS 0.019961f
C11109 DVDD.n844 VSS 0.011429f
C11110 DVDD.n845 VSS 0.019961f
C11111 DVDD.n846 VSS 0.011429f
C11112 DVDD.n847 VSS 0.019961f
C11113 DVDD.n848 VSS 0.019961f
C11114 DVDD.n849 VSS 0.010463f
C11115 DVDD.n850 VSS 0.010946f
C11116 DVDD.n851 VSS 0.019961f
C11117 DVDD.n852 VSS 0.011429f
C11118 DVDD.n853 VSS 0.019961f
C11119 DVDD.n854 VSS 0.011429f
C11120 DVDD.n855 VSS 0.019961f
C11121 DVDD.n856 VSS 0.011429f
C11122 DVDD.n857 VSS 0.019961f
C11123 DVDD.n858 VSS 0.011429f
C11124 DVDD.n859 VSS 0.019961f
C11125 DVDD.n860 VSS 0.011429f
C11126 DVDD.n861 VSS 0.019961f
C11127 DVDD.n862 VSS 0.011429f
C11128 DVDD.n863 VSS 0.019961f
C11129 DVDD.n864 VSS 0.010302f
C11130 DVDD.n865 VSS 0.019961f
C11131 DVDD.n866 VSS 0.019961f
C11132 DVDD.n867 VSS 0.019961f
C11133 DVDD.n868 VSS 0.019961f
C11134 DVDD.n869 VSS 0.019961f
C11135 DVDD.n870 VSS 0.01312f
C11136 DVDD.n871 VSS 0.019961f
C11137 DVDD.n872 VSS 0.011429f
C11138 DVDD.n873 VSS 0.019961f
C11139 DVDD.n874 VSS 0.011429f
C11140 DVDD.n875 VSS 0.019961f
C11141 DVDD.n876 VSS 0.011429f
C11142 DVDD.n877 VSS 0.063742f
C11143 DVDD.n878 VSS 0.00586f
C11144 DVDD.n879 VSS 0.281047f
C11145 DVDD.n880 VSS 0.281047f
C11146 DVDD.n881 VSS 0.281047f
C11147 DVDD.n882 VSS 0.281047f
C11148 DVDD.n883 VSS 0.281047f
C11149 DVDD.n884 VSS 0.281047f
C11150 DVDD.n885 VSS 0.281047f
C11151 DVDD.n886 VSS 0.281047f
C11152 DVDD.n887 VSS 0.281047f
C11153 DVDD.n888 VSS 0.281047f
C11154 DVDD.n889 VSS 0.281047f
C11155 DVDD.n890 VSS 0.281047f
C11156 DVDD.n891 VSS 0.140524f
C11157 DVDD.n892 VSS 0.017326f
C11158 DVDD.n893 VSS 0.00998f
C11159 DVDD.n894 VSS 0.00998f
C11160 DVDD.n895 VSS 0.00998f
C11161 DVDD.n896 VSS 0.00586f
C11162 DVDD.n897 VSS 0.281047f
C11163 DVDD.n898 VSS 0.281047f
C11164 DVDD.n899 VSS 0.281047f
C11165 DVDD.n900 VSS 0.281047f
C11166 DVDD.n901 VSS 0.281047f
C11167 DVDD.n902 VSS 0.281047f
C11168 DVDD.n903 VSS 0.281047f
C11169 DVDD.n904 VSS 0.281047f
C11170 DVDD.n905 VSS 0.281047f
C11171 DVDD.n906 VSS 0.281047f
C11172 DVDD.n907 VSS 0.338444f
C11173 DVDD.n908 VSS 0.338444f
C11174 DVDD.n909 VSS 0.536365f
C11175 DVDD.n910 VSS 0.140524f
C11176 DVDD.n911 VSS 0.281047f
C11177 DVDD.n912 VSS 0.281047f
C11178 DVDD.n913 VSS 0.281047f
C11179 DVDD.n914 VSS 0.091044f
C11180 DVDD.n915 VSS 0.022142f
C11181 DVDD.n916 VSS 0.015871f
C11182 DVDD.n917 VSS 0.015871f
C11183 DVDD.n918 VSS 0.015871f
C11184 DVDD.n919 VSS 0.015871f
C11185 DVDD.n920 VSS 0.015871f
C11186 DVDD.n921 VSS 0.140524f
C11187 DVDD.n922 VSS 0.091044f
C11188 DVDD.n923 VSS 0.015871f
C11189 DVDD.n924 VSS 0.015871f
C11190 DVDD.n925 VSS 0.015871f
C11191 DVDD.n926 VSS 0.015871f
C11192 DVDD.n927 VSS 0.018174f
C11193 DVDD.n928 VSS 0.197746f
C11194 DVDD.n929 VSS 0.018174f
C11195 DVDD.n930 VSS 0.045403f
C11196 DVDD.n931 VSS 0.018174f
C11197 DVDD.n932 VSS 0.060537f
C11198 DVDD.n933 VSS 0.018174f
C11199 DVDD.n934 VSS 0.060537f
C11200 DVDD.n935 VSS 0.060537f
C11201 DVDD.n936 VSS 0.018046f
C11202 DVDD.n937 VSS 0.015999f
C11203 DVDD.n938 VSS 0.060537f
C11204 DVDD.n939 VSS 0.060537f
C11205 DVDD.n940 VSS 0.018174f
C11206 DVDD.n941 VSS 0.015871f
C11207 DVDD.n942 VSS 0.018174f
C11208 DVDD.n943 VSS 0.059376f
C11209 DVDD.n944 VSS 0.06455f
C11210 DVDD.n945 VSS 0.023764f
C11211 DVDD.n946 VSS 0.023764f
C11212 DVDD.n947 VSS 0.023764f
C11213 DVDD.n948 VSS 0.027214f
C11214 DVDD.n949 VSS 0.020098f
C11215 DVDD.n950 VSS 0.018174f
C11216 DVDD.n951 VSS 0.045403f
C11217 DVDD.n952 VSS 0.018174f
C11218 DVDD.n953 VSS 0.060537f
C11219 DVDD.n954 VSS 0.060537f
C11220 DVDD.n955 VSS 0.018046f
C11221 DVDD.n956 VSS 0.015999f
C11222 DVDD.n957 VSS 0.060537f
C11223 DVDD.n958 VSS 0.018174f
C11224 DVDD.n959 VSS 0.060537f
C11225 DVDD.n960 VSS 0.108161f
C11226 DVDD.n961 VSS 0.140937f
C11227 DVDD.n962 VSS 0.027214f
C11228 DVDD.n963 VSS 0.070763f
C11229 DVDD.n964 VSS 0.027214f
C11230 DVDD.n965 VSS 0.049363f
C11231 DVDD.n966 VSS 0.035381f
C11232 DVDD.n967 VSS 0.027214f
C11233 DVDD.n968 VSS 0.056782f
C11234 DVDD.n969 VSS 0.070763f
C11235 DVDD.n970 VSS 0.070763f
C11236 DVDD.n971 VSS 0.140524f
C11237 DVDD.n972 VSS 0.140524f
C11238 DVDD.n973 VSS 0.026448f
C11239 DVDD.n974 VSS 0.140524f
C11240 DVDD.n975 VSS 0.1999f
C11241 DVDD.n976 VSS 0.023765f
C11242 DVDD.n977 VSS 0.023765f
C11243 DVDD.n978 VSS 0.023765f
C11244 DVDD.n979 VSS 0.023765f
C11245 DVDD.n980 VSS 0.023765f
C11246 DVDD.n981 VSS 0.023765f
C11247 DVDD.n982 VSS 0.023765f
C11248 DVDD.n983 VSS 0.023765f
C11249 DVDD.n984 VSS 0.023765f
C11250 DVDD.n985 VSS 0.281047f
C11251 DVDD.n986 VSS 0.281047f
C11252 DVDD.n987 VSS 0.281047f
C11253 DVDD.n988 VSS 0.281047f
C11254 DVDD.n989 VSS 0.188025f
C11255 DVDD.n990 VSS 0.536365f
C11256 DVDD.n991 VSS 0.233546f
C11257 DVDD.n992 VSS 0.281047f
C11258 DVDD.n993 VSS 0.281047f
C11259 DVDD.n994 VSS 0.281047f
C11260 DVDD.n995 VSS 0.281047f
C11261 DVDD.n996 VSS 0.281047f
C11262 DVDD.n997 VSS 0.281047f
C11263 DVDD.n998 VSS 0.281047f
C11264 DVDD.n999 VSS 0.281047f
C11265 DVDD.n1000 VSS 0.281047f
C11266 DVDD.n1001 VSS 0.281047f
C11267 DVDD.n1002 VSS 0.281047f
C11268 DVDD.n1003 VSS 0.281047f
C11269 DVDD.n1004 VSS 0.281047f
C11270 DVDD.n1005 VSS 0.140524f
C11271 DVDD.n1006 VSS 0.281047f
C11272 DVDD.n1007 VSS 0.281047f
C11273 DVDD.n1008 VSS 0.281047f
C11274 DVDD.n1009 VSS 0.281047f
C11275 DVDD.n1010 VSS 0.00998f
C11276 DVDD.n1011 VSS 0.00998f
C11277 DVDD.n1012 VSS 0.00998f
C11278 DVDD.n1013 VSS 0.00998f
C11279 DVDD.n1014 VSS 0.00998f
C11280 DVDD.n1015 VSS 0.00998f
C11281 DVDD.n1016 VSS 0.00998f
C11282 DVDD.n1017 VSS 0.00998f
C11283 DVDD.n1018 VSS 0.00998f
C11284 DVDD.n1019 VSS 0.00998f
C11285 DVDD.n1020 VSS 0.281047f
C11286 DVDD.n1021 VSS 0.281047f
C11287 DVDD.n1022 VSS 0.281047f
C11288 DVDD.n1023 VSS 0.281047f
C11289 DVDD.n1024 VSS 0.281047f
C11290 DVDD.n1025 VSS 0.281047f
C11291 DVDD.n1026 VSS 0.281047f
C11292 DVDD.n1027 VSS 0.281047f
C11293 DVDD.n1028 VSS 0.281047f
C11294 DVDD.n1029 VSS 0.281047f
C11295 DVDD.n1030 VSS 0.281047f
C11296 DVDD.n1031 VSS 0.281047f
C11297 DVDD.n1032 VSS 0.281047f
C11298 DVDD.n1033 VSS 0.281047f
C11299 DVDD.n1034 VSS 0.281047f
C11300 DVDD.n1035 VSS 0.281047f
C11301 DVDD.n1036 VSS 0.281047f
C11302 DVDD.n1037 VSS 0.281047f
C11303 DVDD.n1038 VSS 0.281047f
C11304 DVDD.n1039 VSS 0.281047f
C11305 DVDD.n1040 VSS 0.281047f
C11306 DVDD.n1041 VSS 0.281047f
C11307 DVDD.n1042 VSS 0.281047f
C11308 DVDD.n1043 VSS 0.281047f
C11309 DVDD.n1044 VSS 0.281047f
C11310 DVDD.n1045 VSS 0.281047f
C11311 DVDD.n1046 VSS 0.266203f
C11312 DVDD.n1047 VSS 0.00998f
C11313 DVDD.n1048 VSS 0.00998f
C11314 DVDD.n1049 VSS 0.00998f
C11315 DVDD.n1050 VSS 0.00998f
C11316 DVDD.n1051 VSS 0.00998f
C11317 DVDD.n1052 VSS 0.00998f
C11318 DVDD.n1053 VSS 0.00998f
C11319 DVDD.n1054 VSS 0.00998f
C11320 DVDD.n1055 VSS 0.00998f
C11321 DVDD.n1056 VSS 0.00998f
C11322 DVDD.n1057 VSS 0.018834f
C11323 DVDD.n1058 VSS 0.010302f
C11324 DVDD.n1059 VSS 0.011429f
C11325 DVDD.n1060 VSS 0.063742f
C11326 DVDD.n1061 VSS 0.011429f
C11327 DVDD.n1062 VSS 0.019961f
C11328 DVDD.n1063 VSS 0.011429f
C11329 DVDD.n1064 VSS 0.019961f
C11330 DVDD.n1065 VSS 0.019961f
C11331 DVDD.n1066 VSS 0.01312f
C11332 DVDD.n1067 VSS 0.019961f
C11333 DVDD.n1068 VSS 0.019961f
C11334 DVDD.n1069 VSS 0.019961f
C11335 DVDD.n1070 VSS -0.294669f
C11336 DVDD.n1071 VSS 0.00998f
C11337 DVDD.n1072 VSS 0.019961f
C11338 DVDD.n1073 VSS 0.140524f
C11339 DVDD.n1074 VSS 0.011429f
C11340 DVDD.n1075 VSS 0.155368f
C11341 DVDD.n1076 VSS 0.00998f
C11342 DVDD.n1077 VSS 0.00998f
C11343 DVDD.n1078 VSS 0.00998f
C11344 DVDD.n1079 VSS 0.00998f
C11345 DVDD.n1080 VSS 0.00998f
C11346 DVDD.n1081 VSS 0.00998f
C11347 DVDD.n1082 VSS 0.00998f
C11348 DVDD.n1083 VSS 0.00998f
C11349 DVDD.n1084 VSS 0.00998f
C11350 DVDD.n1085 VSS 0.281047f
C11351 DVDD.n1086 VSS 0.281047f
C11352 DVDD.n1087 VSS 0.281047f
C11353 DVDD.n1088 VSS 0.281047f
C11354 DVDD.n1089 VSS 0.281047f
C11355 DVDD.n1090 VSS 0.281047f
C11356 DVDD.n1091 VSS 0.281047f
C11357 DVDD.n1092 VSS 0.281047f
C11358 DVDD.n1093 VSS 0.281047f
C11359 DVDD.n1094 VSS 0.536365f
C11360 DVDD.n1095 VSS 0.338444f
C11361 DVDD.n1096 VSS 0.281047f
C11362 DVDD.n1097 VSS 0.281047f
C11363 DVDD.n1098 VSS 0.281047f
C11364 DVDD.n1099 VSS 0.281047f
C11365 DVDD.n1100 VSS 0.281047f
C11366 DVDD.n1101 VSS 0.281047f
C11367 DVDD.n1102 VSS 0.281047f
C11368 DVDD.n1103 VSS 0.281047f
C11369 DVDD.n1104 VSS 0.281047f
C11370 DVDD.n1105 VSS 0.281047f
C11371 DVDD.n1106 VSS 1.042f
C11372 DVDD.n1107 VSS 0.281047f
C11373 DVDD.n1108 VSS 0.140524f
C11374 DVDD.n1109 VSS 0.037473f
C11375 DVDD.n1110 VSS 0.037473f
C11376 DVDD.n1111 VSS 0.037473f
C11377 DVDD.n1112 VSS 0.037473f
C11378 DVDD.n1113 VSS 0.037473f
C11379 DVDD.n1114 VSS 0.037473f
C11380 DVDD.n1115 VSS 0.037473f
C11381 DVDD.n1116 VSS 0.037473f
C11382 DVDD.n1117 VSS 0.037473f
C11383 DVDD.n1118 VSS 0.037473f
C11384 DVDD.n1120 VSS 0.628154f
C11385 DVDD.n1121 VSS 0.140524f
C11386 DVDD.n1122 VSS 0.042532f
C11387 DVDD.n1123 VSS 0.042532f
C11388 DVDD.n1124 VSS 0.042532f
C11389 DVDD.n1125 VSS 0.042532f
C11390 DVDD.n1126 VSS 0.042532f
C11391 DVDD.n1127 VSS 0.042532f
C11392 DVDD.n1128 VSS 0.042532f
C11393 DVDD.n1129 VSS 0.042532f
C11394 DVDD.n1130 VSS 0.042532f
C11395 DVDD.n1131 VSS 0.157347f
C11396 DVDD.n1134 VSS 0.042532f
C11397 DVDD.n1136 VSS 0.042532f
C11398 DVDD.n1138 VSS 0.042532f
C11399 DVDD.n1140 VSS 0.042532f
C11400 DVDD.n1142 VSS 0.042532f
C11401 DVDD.n1144 VSS 0.042532f
C11402 DVDD.n1146 VSS 0.042532f
C11403 DVDD.n1148 VSS 0.042532f
C11404 DVDD.n1150 VSS 0.535669f
C11405 DVDD.n1151 VSS 1.042f
C11406 DVDD.n1152 VSS 0.281047f
C11407 DVDD.n1153 VSS 0.281047f
C11408 DVDD.n1154 VSS 0.281047f
C11409 DVDD.n1155 VSS 0.281047f
C11410 DVDD.n1156 VSS 0.281047f
C11411 DVDD.n1157 VSS 0.281047f
C11412 DVDD.n1158 VSS 0.281047f
C11413 DVDD.n1159 VSS 0.281047f
C11414 DVDD.n1160 VSS 0.281047f
C11415 DVDD.n1161 VSS 0.190004f
C11416 DVDD.n1162 VSS 0.281047f
C11417 DVDD.n1163 VSS 0.281047f
C11418 DVDD.n1164 VSS 0.281047f
C11419 DVDD.n1165 VSS 0.281047f
C11420 DVDD.n1166 VSS 0.281047f
C11421 DVDD.n1167 VSS 0.281047f
C11422 DVDD.n1168 VSS 0.281047f
C11423 DVDD.n1169 VSS 0.281047f
C11424 DVDD.n1170 VSS 0.281047f
C11425 DVDD.n1171 VSS 0.281047f
C11426 DVDD.n1172 VSS 0.281047f
C11427 DVDD.n1173 VSS 0.281047f
C11428 DVDD.n1174 VSS 0.281047f
C11429 DVDD.n1175 VSS 0.281047f
C11430 DVDD.n1176 VSS 0.281047f
C11431 DVDD.n1177 VSS 0.281047f
C11432 DVDD.n1178 VSS 0.281047f
C11433 DVDD.n1179 VSS 0.281047f
C11434 DVDD.n1180 VSS 0.281047f
C11435 DVDD.n1181 VSS 0.140524f
C11436 DVDD.n1189 VSS 0.042532f
C11437 DVDD.n1192 VSS 0.065578f
C11438 DVDD.n1193 VSS 0.489671f
C11439 DVDD.n1194 VSS 0.062299f
C11440 DVDD.n1195 VSS 0.041679f
C11441 DVDD.n1196 VSS 0.062299f
C11442 DVDD.n1197 VSS 0.065578f
C11443 DVDD.n1199 VSS 0.062299f
C11444 DVDD.n1200 VSS 0.051769f
C11445 DVDD.n1202 VSS 0.062299f
C11446 DVDD.n1205 VSS 0.194805f
C11447 DVDD.n1206 VSS 0.131155f
C11448 DVDD.n1207 VSS 0.131155f
C11449 DVDD.n1208 VSS 0.131155f
C11450 DVDD.n1209 VSS 0.113145f
C11451 DVDD.n1210 VSS 0.131155f
C11452 DVDD.n1211 VSS 0.131155f
C11453 DVDD.n1212 VSS 0.131155f
C11454 DVDD.n1213 VSS 0.131155f
C11455 DVDD.n1214 VSS 0.016868f
C11456 DVDD.n1215 VSS 0.008917f
C11457 DVDD.n1216 VSS 0.008917f
C11458 DVDD.n1217 VSS 0.008917f
C11459 DVDD.n1218 VSS 0.065578f
C11460 DVDD.n1219 VSS 0.008917f
C11461 DVDD.n1220 VSS 0.005537f
C11462 DVDD.n1221 VSS 0.008917f
C11463 DVDD.n1222 VSS 0.003713f
C11464 DVDD.n1223 VSS 0.131155f
C11465 DVDD.n1224 VSS 0.131155f
C11466 DVDD.n1225 VSS 0.131155f
C11467 DVDD.n1226 VSS 0.131155f
C11468 DVDD.n1227 VSS 0.131155f
C11469 DVDD.n1228 VSS 0.131155f
C11470 DVDD.n1229 VSS 0.131155f
C11471 DVDD.n1230 VSS 0.131155f
C11472 DVDD.n1231 VSS 0.131155f
C11473 DVDD.n1232 VSS 0.131155f
C11474 DVDD.n1233 VSS 0.131155f
C11475 DVDD.n1234 VSS 0.131155f
C11476 DVDD.n1235 VSS 0.131155f
C11477 DVDD.n1236 VSS 0.131155f
C11478 DVDD.n1237 VSS 0.131155f
C11479 DVDD.n1238 VSS 0.131155f
C11480 DVDD.n1239 VSS 0.131155f
C11481 DVDD.n1240 VSS 0.131155f
C11482 DVDD.n1241 VSS 0.131155f
C11483 DVDD.n1242 VSS 0.131155f
C11484 DVDD.n1243 VSS 0.131155f
C11485 DVDD.n1244 VSS 0.131155f
C11486 DVDD.n1245 VSS 0.131155f
C11487 DVDD.n1246 VSS 0.131155f
C11488 DVDD.n1247 VSS 0.131155f
C11489 DVDD.n1248 VSS 0.131155f
C11490 DVDD.n1249 VSS 0.131155f
C11491 DVDD.n1250 VSS 0.131155f
C11492 DVDD.n1251 VSS 0.131155f
C11493 DVDD.n1252 VSS 0.131155f
C11494 DVDD.n1253 VSS 0.131155f
C11495 DVDD.n1254 VSS 0.131155f
C11496 DVDD.n1255 VSS 0.131155f
C11497 DVDD.n1256 VSS 0.131155f
C11498 DVDD.n1257 VSS 0.131155f
C11499 DVDD.n1258 VSS 0.131155f
C11500 DVDD.n1259 VSS 0.131155f
C11501 DVDD.n1260 VSS 0.131155f
C11502 DVDD.n1261 VSS 0.131155f
C11503 DVDD.n1262 VSS 0.131155f
C11504 DVDD.n1263 VSS 0.131155f
C11505 DVDD.n1264 VSS 0.131155f
C11506 DVDD.n1265 VSS 0.131155f
C11507 DVDD.n1266 VSS 0.131155f
C11508 DVDD.n1267 VSS 0.131155f
C11509 DVDD.n1268 VSS 0.131155f
C11510 DVDD.n1269 VSS 0.131155f
C11511 DVDD.n1270 VSS 0.131155f
C11512 DVDD.n1271 VSS 0.131155f
C11513 DVDD.n1272 VSS 0.131155f
C11514 DVDD.n1273 VSS 0.131155f
C11515 DVDD.n1274 VSS 0.131155f
C11516 DVDD.n1275 VSS 0.131155f
C11517 DVDD.n1276 VSS 0.131155f
C11518 DVDD.n1277 VSS 0.131155f
C11519 DVDD.n1278 VSS 0.131155f
C11520 DVDD.n1279 VSS 0.131155f
C11521 DVDD.n1280 VSS 0.131155f
C11522 DVDD.n1281 VSS 0.131155f
C11523 DVDD.n1282 VSS 0.131155f
C11524 DVDD.n1283 VSS 0.131155f
C11525 DVDD.n1284 VSS 0.131155f
C11526 DVDD.n1285 VSS 0.131155f
C11527 DVDD.n1286 VSS 0.131155f
C11528 DVDD.n1287 VSS 0.131155f
C11529 DVDD.n1288 VSS 0.131155f
C11530 DVDD.n1289 VSS 0.131155f
C11531 DVDD.n1290 VSS 0.131155f
C11532 DVDD.n1291 VSS 0.131155f
C11533 DVDD.n1292 VSS 0.131155f
C11534 DVDD.n1293 VSS 0.131155f
C11535 DVDD.n1294 VSS 0.131155f
C11536 DVDD.n1295 VSS 0.131155f
C11537 DVDD.n1296 VSS 0.131155f
C11538 DVDD.n1297 VSS 0.131155f
C11539 DVDD.n1298 VSS 0.131155f
C11540 DVDD.n1299 VSS 0.131155f
C11541 DVDD.n1300 VSS 0.131155f
C11542 DVDD.n1301 VSS 0.117763f
C11543 DVDD.n1302 VSS 0.131155f
C11544 DVDD.n1303 VSS 0.131155f
C11545 DVDD.n1304 VSS 0.131155f
C11546 DVDD.n1305 VSS 0.065578f
C11547 DVDD.n1306 VSS 0.005537f
C11548 DVDD.n1307 VSS 0.008917f
C11549 DVDD.n1308 VSS 0.008917f
C11550 DVDD.n1309 VSS 0.016868f
C11551 DVDD.n1310 VSS 0.07897f
C11552 DVDD.n1311 VSS 0.008917f
C11553 DVDD.n1312 VSS 0.008917f
C11554 DVDD.n1313 VSS 0.008917f
C11555 DVDD.n1314 VSS 0.010211f
C11556 DVDD.n1315 VSS 0.036896f
C11557 DVDD.n1316 VSS 0.033417f
C11558 DVDD.n1317 VSS 0.010211f
C11559 DVDD.n1318 VSS 0.010211f
C11560 DVDD.n1320 VSS 0.010211f
C11561 DVDD.n1321 VSS 0.008989f
C11562 DVDD.n1322 VSS 0.010139f
C11563 DVDD.n1323 VSS 0.138114f
C11564 DVDD.n1324 VSS 0.010211f
C11565 DVDD.n1325 VSS 1.48827f
C11566 DVDD.n1326 VSS 8.59664f
C11567 DVDD.n1327 VSS 3.64002f
C11568 DVDD.n1328 VSS 2.54694f
C11569 DVDD.n1329 VSS 0.028026f
C11570 DVDD.n1331 VSS 0.065578f
C11571 DVDD.n1332 VSS 0.033726f
C11572 DVDD.n1335 VSS 0.033726f
C11573 DVDD.n1336 VSS 0.025888f
C11574 DVDD.n1337 VSS 0.065578f
C11575 DVDD.n1339 VSS 0.033726f
C11576 DVDD.n1340 VSS 0.065578f
C11577 DVDD.n1342 VSS 0.131155f
C11578 DVDD.n1343 VSS 0.131155f
C11579 DVDD.n1344 VSS 0.131155f
C11580 DVDD.n1345 VSS 0.131155f
C11581 DVDD.n1346 VSS 0.131155f
C11582 DVDD.n1347 VSS 0.131155f
C11583 DVDD.n1348 VSS 0.131155f
C11584 DVDD.n1349 VSS 0.131155f
C11585 DVDD.n1350 VSS 0.131155f
C11586 DVDD.n1351 VSS 0.131155f
C11587 DVDD.n1352 VSS 0.131155f
C11588 DVDD.n1353 VSS 0.131155f
C11589 DVDD.n1354 VSS 0.131155f
C11590 DVDD.n1355 VSS 0.131155f
C11591 DVDD.n1356 VSS 0.131155f
C11592 DVDD.n1357 VSS 0.118225f
C11593 DVDD.n1358 VSS 0.118225f
C11594 DVDD.n1359 VSS 0.131155f
C11595 DVDD.n1360 VSS 0.067425f
C11596 DVDD.n1361 VSS 0.078508f
C11597 DVDD.n1362 VSS 0.21425f
C11598 DVDD.n1363 VSS 0.453156f
C11599 DVDD.n1364 VSS 0.507717f
C11600 DVDD.n1365 VSS 0.033726f
C11601 DVDD.n1367 VSS 0.025888f
C11602 DVDD.n1368 VSS 0.012931f
C11603 DVDD.n1369 VSS 0.022563f
C11604 DVDD.n1370 VSS 1.14562f
C11605 DVDD.n1371 VSS 1.16514f
C11606 DVDD.n1372 VSS 7.6398f
C11607 DVDD.n1373 VSS 5.65298f
C11608 DVDD.n1374 VSS 2.40462f
C11609 DVDD.n1375 VSS 5.66119f
C11610 DVDD.n1376 VSS 7.90719f
C11611 DVDD.n1377 VSS 8.86412f
C11612 DVDD.n1378 VSS 10.9093f
C11613 DVDD.n1379 VSS 5.88404f
C11614 DVDD.n1380 VSS 1.48355f
C11615 DVDD.n1381 VSS 0.010211f
C11616 DVDD.n1382 VSS 0.010211f
C11617 DVDD.n1383 VSS 0.008989f
C11618 DVDD.n1385 VSS 0.010139f
C11619 DVDD.n1386 VSS 0.010211f
C11620 DVDD.n1387 VSS 0.010211f
C11621 DVDD.n1388 VSS 0.112907f
C11622 DVDD.n1389 VSS 0.033417f
C11623 DVDD.n1390 VSS 0.010211f
C11624 DVDD.n1391 VSS 0.036896f
C11625 DVDD.n1392 VSS 0.003713f
C11626 DVDD.n1393 VSS 0.014701f
C11627 DVDD.n1394 VSS 0.065578f
C11628 DVDD.n1395 VSS 0.065578f
C11629 DVDD.n1396 VSS 0.131155f
C11630 DVDD.n1397 VSS 0.131155f
C11631 DVDD.n1398 VSS 0.131155f
C11632 DVDD.n1399 VSS 0.131155f
C11633 DVDD.n1400 VSS 0.131155f
C11634 DVDD.n1401 VSS 0.131155f
C11635 DVDD.n1402 VSS 0.131155f
C11636 DVDD.n1403 VSS 0.131155f
C11637 DVDD.n1404 VSS 0.131155f
C11638 DVDD.n1405 VSS 0.131155f
C11639 DVDD.n1406 VSS 0.131155f
C11640 DVDD.n1407 VSS 0.131155f
C11641 DVDD.n1408 VSS 0.131155f
C11642 DVDD.n1409 VSS 0.131155f
C11643 DVDD.n1410 VSS 0.131155f
C11644 DVDD.n1411 VSS 0.131155f
C11645 DVDD.n1412 VSS 0.131155f
C11646 DVDD.n1413 VSS 0.131155f
C11647 DVDD.n1414 VSS 0.131155f
C11648 DVDD.n1415 VSS 0.131155f
C11649 DVDD.n1416 VSS 0.131155f
C11650 DVDD.n1417 VSS 0.131155f
C11651 DVDD.n1418 VSS 0.131155f
C11652 DVDD.n1419 VSS 0.131155f
C11653 DVDD.n1420 VSS 0.131155f
C11654 DVDD.n1421 VSS 0.131155f
C11655 DVDD.n1422 VSS 0.131155f
C11656 DVDD.n1423 VSS 0.131155f
C11657 DVDD.n1424 VSS 0.131155f
C11658 DVDD.n1425 VSS 0.131155f
C11659 DVDD.n1426 VSS 0.131155f
C11660 DVDD.n1427 VSS 0.131155f
C11661 DVDD.n1428 VSS 0.131155f
C11662 DVDD.n1429 VSS 0.131155f
C11663 DVDD.n1430 VSS 0.131155f
C11664 DVDD.n1431 VSS 0.131155f
C11665 DVDD.n1432 VSS 0.131155f
C11666 DVDD.n1433 VSS 0.131155f
C11667 DVDD.n1434 VSS 0.131155f
C11668 DVDD.n1435 VSS 0.131155f
C11669 DVDD.n1436 VSS 0.131155f
C11670 DVDD.n1437 VSS 0.131155f
C11671 DVDD.n1438 VSS 0.131155f
C11672 DVDD.n1439 VSS 0.131155f
C11673 DVDD.n1440 VSS 0.131155f
C11674 DVDD.n1441 VSS 0.131155f
C11675 DVDD.n1442 VSS 0.131155f
C11676 DVDD.n1443 VSS 0.131155f
C11677 DVDD.n1444 VSS 0.131155f
C11678 DVDD.n1445 VSS 0.131155f
C11679 DVDD.n1446 VSS 0.131155f
C11680 DVDD.n1447 VSS 0.131155f
C11681 DVDD.n1448 VSS 0.131155f
C11682 DVDD.n1449 VSS 0.131155f
C11683 DVDD.n1450 VSS 0.131155f
C11684 DVDD.n1451 VSS 0.131155f
C11685 DVDD.n1452 VSS 0.131155f
C11686 DVDD.n1453 VSS 0.131155f
C11687 DVDD.n1454 VSS 0.131155f
C11688 DVDD.n1455 VSS 0.131155f
C11689 DVDD.n1456 VSS 0.131155f
C11690 DVDD.n1457 VSS 0.131155f
C11691 DVDD.n1458 VSS 0.131155f
C11692 DVDD.n1459 VSS 0.131155f
C11693 DVDD.n1460 VSS 0.131155f
C11694 DVDD.n1461 VSS 0.131155f
C11695 DVDD.n1462 VSS 0.131155f
C11696 DVDD.n1463 VSS 0.131155f
C11697 DVDD.n1464 VSS 0.131155f
C11698 DVDD.n1465 VSS 0.131155f
C11699 DVDD.n1466 VSS 0.131155f
C11700 DVDD.n1467 VSS 0.131155f
C11701 DVDD.n1468 VSS 0.131155f
C11702 DVDD.n1469 VSS 0.131155f
C11703 DVDD.n1470 VSS 0.131155f
C11704 DVDD.n1471 VSS 0.131155f
C11705 DVDD.n1472 VSS 0.131155f
C11706 DVDD.n1473 VSS 0.131155f
C11707 DVDD.n1474 VSS 0.131155f
C11708 DVDD.n1475 VSS 0.131155f
C11709 DVDD.n1476 VSS 0.131155f
C11710 DVDD.n1477 VSS 0.131155f
C11711 DVDD.n1478 VSS 0.131155f
C11712 DVDD.n1479 VSS 0.131155f
C11713 DVDD.n1480 VSS 0.131155f
C11714 DVDD.n1481 VSS 0.131155f
C11715 DVDD.n1482 VSS 0.131155f
C11716 DVDD.n1483 VSS 0.131155f
C11717 DVDD.n1484 VSS 0.131155f
C11718 DVDD.n1485 VSS 0.131155f
C11719 DVDD.n1486 VSS 0.131155f
C11720 DVDD.n1487 VSS 0.131155f
C11721 DVDD.n1488 VSS 0.131155f
C11722 DVDD.n1489 VSS 0.131155f
C11723 DVDD.n1490 VSS 0.131155f
C11724 DVDD.n1491 VSS 0.131155f
C11725 DVDD.n1492 VSS 0.131155f
C11726 DVDD.n1493 VSS 0.131155f
C11727 DVDD.n1494 VSS 0.131155f
C11728 DVDD.n1495 VSS 0.131155f
C11729 DVDD.n1496 VSS 0.131155f
C11730 DVDD.n1497 VSS 0.131155f
C11731 DVDD.n1498 VSS 0.131155f
C11732 DVDD.n1499 VSS 0.131155f
C11733 DVDD.n1500 VSS 0.131155f
C11734 DVDD.n1501 VSS 0.131155f
C11735 DVDD.n1502 VSS 0.131155f
C11736 DVDD.n1503 VSS 0.131155f
C11737 DVDD.n1504 VSS 0.131155f
C11738 DVDD.n1505 VSS 0.131155f
C11739 DVDD.n1506 VSS 0.131155f
C11740 DVDD.n1507 VSS 0.131155f
C11741 DVDD.n1508 VSS 0.131155f
C11742 DVDD.n1509 VSS 0.131155f
C11743 DVDD.n1510 VSS 0.131155f
C11744 DVDD.n1511 VSS 0.131155f
C11745 DVDD.n1512 VSS 0.131155f
C11746 DVDD.n1513 VSS 0.131155f
C11747 DVDD.n1514 VSS 0.131155f
C11748 DVDD.n1515 VSS 0.131155f
C11749 DVDD.n1516 VSS 0.131155f
C11750 DVDD.n1517 VSS 0.131155f
C11751 DVDD.n1518 VSS 0.131155f
C11752 DVDD.n1519 VSS 0.131155f
C11753 DVDD.n1520 VSS 0.131155f
C11754 DVDD.n1521 VSS 0.131155f
C11755 DVDD.n1522 VSS 0.131155f
C11756 DVDD.n1523 VSS 0.131155f
C11757 DVDD.n1524 VSS 0.131155f
C11758 DVDD.n1525 VSS 0.131155f
C11759 DVDD.n1526 VSS 0.131155f
C11760 DVDD.n1527 VSS 0.131155f
C11761 DVDD.n1528 VSS 0.131155f
C11762 DVDD.n1529 VSS 0.131155f
C11763 DVDD.n1530 VSS 0.131155f
C11764 DVDD.n1531 VSS 0.131155f
C11765 DVDD.n1532 VSS 0.131155f
C11766 DVDD.n1533 VSS 0.131155f
C11767 DVDD.n1534 VSS 0.131155f
C11768 DVDD.n1535 VSS 0.131155f
C11769 DVDD.n1536 VSS 0.131155f
C11770 DVDD.n1537 VSS 0.131155f
C11771 DVDD.n1538 VSS 0.131155f
C11772 DVDD.n1539 VSS 0.131155f
C11773 DVDD.n1540 VSS 0.131155f
C11774 DVDD.n1541 VSS 0.131155f
C11775 DVDD.n1542 VSS 0.131155f
C11776 DVDD.n1543 VSS 0.131155f
C11777 DVDD.n1544 VSS 0.131155f
C11778 DVDD.n1545 VSS 0.131155f
C11779 DVDD.n1546 VSS 0.131155f
C11780 DVDD.n1547 VSS 0.131155f
C11781 DVDD.n1548 VSS 0.131155f
C11782 DVDD.n1549 VSS 0.131155f
C11783 DVDD.n1550 VSS 0.131155f
C11784 DVDD.n1551 VSS 0.131155f
C11785 DVDD.n1552 VSS 0.131155f
C11786 DVDD.n1553 VSS 0.125152f
C11787 DVDD.n1554 VSS 0.065578f
C11788 DVDD.n1555 VSS 0.014701f
C11789 DVDD.n1556 VSS 0.065578f
C11790 DVDD.n1557 VSS 0.071581f
C11791 DVDD.n1558 VSS 0.131155f
C11792 DVDD.n1559 VSS 0.131155f
C11793 DVDD.n1560 VSS 0.131155f
C11794 DVDD.n1561 VSS 0.131155f
C11795 DVDD.n1562 VSS 0.131155f
C11796 DVDD.n1563 VSS 0.131155f
C11797 DVDD.n1564 VSS 0.131155f
C11798 DVDD.n1565 VSS 0.131155f
C11799 DVDD.n1566 VSS 0.131155f
C11800 DVDD.n1567 VSS 0.131155f
C11801 DVDD.n1568 VSS 0.131155f
C11802 DVDD.n1569 VSS 0.131155f
C11803 DVDD.n1570 VSS 0.710188f
C11804 DVDD.n1571 VSS 0.131155f
C11805 DVDD.n1572 VSS 0.065578f
C11806 DVDD.n1573 VSS 0.065578f
C11807 DVDD.n1575 VSS 0.047821f
C11808 DVDD.n1576 VSS 0.513093f
C11809 DVDD.n1577 VSS 0.188516f
C11810 DVDD.n1578 VSS 0.182545f
C11811 DVDD.n1579 VSS 0.140524f
C11812 DVDD.n1581 VSS 0.042532f
C11813 DVDD.n1582 VSS 0.140524f
C11814 DVDD.n1583 VSS 0.072333f
C11815 DVDD.n1584 VSS 0.065521f
C11816 DVDD.n1585 VSS 0.037473f
C11817 DVDD.n1586 VSS 0.037473f
C11818 DVDD.n1587 VSS 0.037473f
C11819 DVDD.n1588 VSS 0.037473f
C11820 DVDD.n1589 VSS 0.037473f
C11821 DVDD.n1590 VSS 0.037473f
C11822 DVDD.n1591 VSS 0.037473f
C11823 DVDD.n1592 VSS 0.037473f
C11824 DVDD.n1593 VSS 0.037473f
C11825 DVDD.n1595 VSS 0.628154f
C11826 DVDD.n1596 VSS 0.140524f
C11827 DVDD.n1597 VSS 0.037473f
C11828 DVDD.n1598 VSS 0.037473f
C11829 DVDD.n1599 VSS 0.037473f
C11830 DVDD.n1600 VSS 0.037473f
C11831 DVDD.n1601 VSS 0.037473f
C11832 DVDD.n1602 VSS 0.037473f
C11833 DVDD.n1603 VSS 0.037473f
C11834 DVDD.n1604 VSS 0.037473f
C11835 DVDD.n1605 VSS 0.037473f
C11836 DVDD.n1606 VSS 0.037473f
C11837 DVDD.n1607 VSS 0.157347f
C11838 DVDD.n1609 VSS 0.037473f
C11839 DVDD.n1611 VSS 0.037473f
C11840 DVDD.n1613 VSS 0.037473f
C11841 DVDD.n1615 VSS 0.037473f
C11842 DVDD.n1617 VSS 0.037473f
C11843 DVDD.n1619 VSS 0.037473f
C11844 DVDD.n1621 VSS 0.037473f
C11845 DVDD.n1623 VSS 0.037473f
C11846 DVDD.n1625 VSS 0.037473f
C11847 DVDD.n1627 VSS 0.628154f
C11848 DVDD.n1628 VSS 0.140524f
C11849 DVDD.n1629 VSS 0.037473f
C11850 DVDD.n1630 VSS 0.037473f
C11851 DVDD.n1631 VSS 0.037473f
C11852 DVDD.n1632 VSS 0.037473f
C11853 DVDD.n1633 VSS 0.037473f
C11854 DVDD.n1634 VSS 0.037473f
C11855 DVDD.n1635 VSS 0.037473f
C11856 DVDD.n1636 VSS 0.037473f
C11857 DVDD.n1637 VSS 0.037473f
C11858 DVDD.n1638 VSS 0.037473f
C11859 DVDD.n1639 VSS 0.157347f
C11860 DVDD.n1641 VSS 0.037473f
C11861 DVDD.n1643 VSS 0.037473f
C11862 DVDD.n1645 VSS 0.037473f
C11863 DVDD.n1647 VSS 0.037473f
C11864 DVDD.n1649 VSS 0.037473f
C11865 DVDD.n1651 VSS 0.037473f
C11866 DVDD.n1653 VSS 0.037473f
C11867 DVDD.n1655 VSS 0.037473f
C11868 DVDD.n1657 VSS 0.037473f
C11869 DVDD.n1658 VSS 0.037473f
C11870 DVDD.n1659 VSS 0.040424f
C11871 DVDD.n1660 VSS 0.080848f
C11872 DVDD.n1661 VSS 0.080848f
C11873 DVDD.n1662 VSS 0.080848f
C11874 DVDD.n1663 VSS 0.040424f
C11875 DVDD.n1664 VSS 0.037473f
C11876 DVDD.n1665 VSS 0.02135f
C11877 DVDD.n1666 VSS 0.057312f
C11878 DVDD.n1667 VSS 0.059497f
C11879 DVDD.n1668 VSS 0.149892f
C11880 DVDD.n1669 VSS 0.149892f
C11881 DVDD.n1670 VSS 0.047634f
C11882 DVDD.n1671 VSS 0.149892f
C11883 DVDD.n1672 VSS 0.149892f
C11884 DVDD.n1673 VSS 0.149892f
C11885 DVDD.n1674 VSS 0.149892f
C11886 DVDD.n1675 VSS 0.075143f
C11887 DVDD.n1676 VSS 0.149892f
C11888 DVDD.n1677 VSS 0.149892f
C11889 DVDD.n1678 VSS 0.149892f
C11890 DVDD.n1679 VSS 0.074946f
C11891 DVDD.n1680 VSS 0.074946f
C11892 DVDD.n1681 VSS 0.074946f
C11893 DVDD.n1682 VSS 0.012388f
C11894 DVDD.n1683 VSS 0.00534f
C11895 DVDD.n1684 VSS 0.025334f
C11896 DVDD.n1685 VSS 0.21547f
C11897 DVDD.n1686 VSS 0.124558f
C11898 DVDD.n1687 VSS 0.188025f
C11899 DVDD.n1688 VSS 0.281047f
C11900 DVDD.n1689 VSS 0.281047f
C11901 DVDD.n1690 VSS 0.170572f
C11902 DVDD.n1691 VSS 0.218072f
C11903 DVDD.n1692 VSS 0.281047f
C11904 DVDD.n1693 VSS 0.281047f
C11905 DVDD.n1694 VSS 0.281047f
C11906 DVDD.n1695 VSS 0.216021f
C11907 DVDD.n1696 VSS 0.281047f
C11908 DVDD.n1697 VSS 0.281047f
C11909 DVDD.n1698 VSS 0.281047f
C11910 DVDD.n1699 VSS 0.281047f
C11911 DVDD.n1700 VSS 0.163285f
C11912 DVDD.n1701 VSS 0.281047f
C11913 DVDD.n1702 VSS 0.281047f
C11914 DVDD.n1703 VSS 0.281047f
C11915 DVDD.n1704 VSS 0.281047f
C11916 DVDD.n1705 VSS 0.281047f
C11917 DVDD.n1706 VSS 0.152357f
C11918 DVDD.n1707 VSS 0.163285f
C11919 DVDD.n1708 VSS 0.038425f
C11920 DVDD.t29 VSS 0.594134f
C11921 DVDD.n1709 VSS -0.068036f
C11922 DVDD.t184 VSS 0.435346f
C11923 DVDD.t183 VSS 0.435346f
C11924 DVDD.n1710 VSS 0.055284f
C11925 DVDD.n1711 VSS -0.068036f
C11926 DVDD.t170 VSS 0.594134f
C11927 DVDD.n1712 VSS 0.237835f
C11928 DVDD.n1713 VSS 0.051157f
C11929 DVDD.t171 VSS 0.09794f
C11930 DVDD.n1714 VSS 0.125601f
C11931 DVDD.t72 VSS 0.041167f
C11932 DVDD.t74 VSS 0.041167f
C11933 DVDD.n1715 VSS 0.082335f
C11934 DVDD.n1716 VSS 0.101471f
C11935 DVDD.t70 VSS 0.09794f
C11936 DVDD.n1717 VSS 0.172003f
C11937 DVDD.n1718 VSS 0.044349f
C11938 DVDD.n1719 VSS 0.00534f
C11939 DVDD.n1720 VSS 0.00712f
C11940 DVDD.n1721 VSS 0.074946f
C11941 DVDD.n1722 VSS 0.117235f
C11942 DVDD.n1723 VSS 0.149892f
C11943 DVDD.n1724 VSS 0.21547f
C11944 DVDD.n1725 VSS 0.149892f
C11945 DVDD.n1726 VSS 0.149892f
C11946 DVDD.n1727 VSS 0.149892f
C11947 DVDD.n1728 VSS 0.062279f
C11948 DVDD.n1729 VSS 0.074946f
C11949 DVDD.n1730 VSS 0.075143f
C11950 DVDD.n1731 VSS 0.149892f
C11951 DVDD.n1732 VSS 0.149892f
C11952 DVDD.n1733 VSS 0.149892f
C11953 DVDD.n1734 VSS 0.126669f
C11954 DVDD.n1735 VSS 0.149892f
C11955 DVDD.n1736 VSS 0.149892f
C11956 DVDD.n1737 VSS 0.129836f
C11957 DVDD.n1738 VSS 0.129836f
C11958 DVDD.n1739 VSS 0.377065f
C11959 DVDD.n1740 VSS 0.472616f
C11960 DVDD.n1741 VSS 0.170869f
C11961 DVDD.n1742 VSS 0.371442f
C11962 DVDD.n1743 VSS 0.453406f
C11963 DVDD.n1744 VSS 0.129836f
C11964 DVDD.n1745 VSS 0.149892f
C11965 DVDD.n1746 VSS 0.149892f
C11966 DVDD.n1747 VSS 0.149892f
C11967 DVDD.n1748 VSS 0.149892f
C11968 DVDD.n1749 VSS 0.149892f
C11969 DVDD.n1750 VSS 0.149892f
C11970 DVDD.n1751 VSS 0.149892f
C11971 DVDD.n1752 VSS 0.149892f
C11972 DVDD.n1753 VSS 0.149892f
C11973 DVDD.n1754 VSS 0.149892f
C11974 DVDD.n1755 VSS 0.149892f
C11975 DVDD.n1756 VSS 0.149892f
C11976 DVDD.n1757 VSS 0.149892f
C11977 DVDD.n1758 VSS 0.149892f
C11978 DVDD.n1759 VSS 0.074946f
C11979 DVDD.n1760 VSS 0.074946f
C11980 DVDD.n1761 VSS 0.012388f
C11981 DVDD.n1762 VSS 0.00712f
C11982 DVDD.n1763 VSS 0.074946f
C11983 DVDD.n1764 VSS 0.074946f
C11984 DVDD.n1765 VSS 0.137225f
C11985 DVDD.n1766 VSS 0.137225f
C11986 DVDD.n1767 VSS 0.281047f
C11987 DVDD.n1768 VSS 0.281047f
C11988 DVDD.n1769 VSS 0.218072f
C11989 DVDD.n1770 VSS 0.281047f
C11990 DVDD.n1771 VSS 0.281047f
C11991 DVDD.n1772 VSS 0.281047f
C11992 DVDD.n1773 VSS 0.281047f
C11993 DVDD.n1774 VSS 0.281047f
C11994 DVDD.n1775 VSS 0.281047f
C11995 DVDD.n1776 VSS 0.281047f
C11996 DVDD.n1777 VSS 0.281047f
C11997 DVDD.n1778 VSS 0.281047f
C11998 DVDD.n1779 VSS 0.281047f
C11999 DVDD.n1780 VSS 0.270162f
C12000 DVDD.n1781 VSS 0.281047f
C12001 DVDD.n1782 VSS 0.281047f
C12002 DVDD.n1783 VSS 0.281047f
C12003 DVDD.n1784 VSS 0.281047f
C12004 DVDD.t136 VSS 0.09794f
C12005 DVDD.n1785 VSS 0.143921f
C12006 DVDD.n1786 VSS 0.208806f
C12007 DVDD.n1787 VSS 0.281047f
C12008 DVDD.n1788 VSS 0.24938f
C12009 DVDD.n1789 VSS 0.172191f
C12010 DVDD.n1790 VSS 0.091835f
C12011 DVDD.n1791 VSS 0.149892f
C12012 DVDD.n1792 VSS 0.21547f
C12013 DVDD.n1793 VSS 0.149892f
C12014 DVDD.n1794 VSS 0.091835f
C12015 DVDD.n1795 VSS 0.281047f
C12016 DVDD.n1796 VSS 0.281047f
C12017 DVDD.n1797 VSS 0.281047f
C12018 DVDD.n1798 VSS 0.281047f
C12019 DVDD.n1799 VSS 0.281047f
C12020 DVDD.n1800 VSS 0.281047f
C12021 DVDD.n1801 VSS 0.281047f
C12022 DVDD.n1802 VSS 0.281047f
C12023 DVDD.n1803 VSS 0.281047f
C12024 DVDD.n1804 VSS 0.281047f
C12025 DVDD.n1805 VSS 0.281047f
C12026 DVDD.n1806 VSS 0.281047f
C12027 DVDD.n1807 VSS 0.264224f
C12028 DVDD.n1808 VSS 0.281047f
C12029 DVDD.n1809 VSS 0.281047f
C12030 DVDD.n1810 VSS 0.281047f
C12031 DVDD.n1811 VSS 0.281047f
C12032 DVDD.n1812 VSS 0.281047f
C12033 DVDD.n1813 VSS 0.281047f
C12034 DVDD.n1814 VSS 0.281047f
C12035 DVDD.n1815 VSS 0.281047f
C12036 DVDD.n1816 VSS 0.281047f
C12037 DVDD.n1817 VSS 0.21547f
C12038 DVDD.n1818 VSS 0.21547f
C12039 DVDD.n1819 VSS 0.149892f
C12040 DVDD.n1820 VSS 0.149892f
C12041 DVDD.n1821 VSS 0.149892f
C12042 DVDD.n1822 VSS 0.149892f
C12043 DVDD.n1823 VSS 0.149892f
C12044 DVDD.n1824 VSS 0.149892f
C12045 DVDD.n1825 VSS 0.149892f
C12046 DVDD.n1826 VSS 0.149892f
C12047 DVDD.n1827 VSS 0.149892f
C12048 DVDD.n1828 VSS 0.149892f
C12049 DVDD.n1829 VSS 0.437123f
C12050 DVDD.n1830 VSS 0.178748f
C12051 DVDD.n1831 VSS 0.169208f
C12052 DVDD.n1832 VSS 0.149892f
C12053 DVDD.n1833 VSS 0.149892f
C12054 DVDD.n1834 VSS 0.149892f
C12055 DVDD.n1835 VSS 0.149892f
C12056 DVDD.n1836 VSS 0.075143f
C12057 DVDD.n1837 VSS 0.149892f
C12058 DVDD.n1838 VSS 0.149892f
C12059 DVDD.n1839 VSS 0.149892f
C12060 DVDD.n1840 VSS 0.074946f
C12061 DVDD.n1841 VSS 0.074946f
C12062 DVDD.n1842 VSS 0.00534f
C12063 DVDD.n1843 VSS 0.074946f
C12064 DVDD.n1844 VSS 0.281047f
C12065 DVDD.n1845 VSS 0.281047f
C12066 DVDD.n1846 VSS 0.281047f
C12067 DVDD.n1847 VSS 0.281047f
C12068 DVDD.n1848 VSS 0.281047f
C12069 DVDD.n1849 VSS 0.281047f
C12070 DVDD.n1850 VSS 0.281047f
C12071 DVDD.n1851 VSS 0.281047f
C12072 DVDD.n1852 VSS 0.218072f
C12073 DVDD.n1853 VSS 0.281047f
C12074 DVDD.n1854 VSS 0.281047f
C12075 DVDD.n1855 VSS 0.281047f
C12076 DVDD.n1856 VSS 0.140524f
C12077 DVDD.n1861 VSS 0.03048f
C12078 DVDD.t185 VSS 0.517068f
C12079 DVDD.t97 VSS 0.041167f
C12080 DVDD.t143 VSS 0.041167f
C12081 DVDD.n1867 VSS 0.082335f
C12082 DVDD.n1868 VSS 0.13166f
C12083 DVDD.n1869 VSS 0.068024f
C12084 DVDD.t190 VSS 0.041167f
C12085 DVDD.t151 VSS 0.041167f
C12086 DVDD.n1870 VSS 0.082335f
C12087 DVDD.n1871 VSS 0.130607f
C12088 DVDD.t32 VSS 0.09794f
C12089 DVDD.n1872 VSS 0.172003f
C12090 DVDD.t213 VSS 0.032179f
C12091 DVDD.n1873 VSS 0.163921f
C12092 DVDD.t30 VSS 0.09794f
C12093 DVDD.n1874 VSS 0.125601f
C12094 DVDD.n1875 VSS 0.051157f
C12095 DVDD.t34 VSS 0.041167f
C12096 DVDD.t28 VSS 0.041167f
C12097 DVDD.n1876 VSS 0.082335f
C12098 DVDD.n1877 VSS 0.102524f
C12099 DVDD.n1878 VSS 0.057077f
C12100 DVDD.n1879 VSS 0.054855f
C12101 DVDD.n1880 VSS 0.00356f
C12102 DVDD.n1881 VSS 0.010429f
C12103 DVDD.n1882 VSS 0.03941f
C12104 DVDD.n1883 VSS -0.064095f
C12105 DVDD.t27 VSS 0.480029f
C12106 DVDD.t33 VSS 0.480029f
C12107 DVDD.t31 VSS 0.649219f
C12108 DVDD.t150 VSS 0.649219f
C12109 DVDD.t189 VSS 0.382474f
C12110 DVDD.t93 VSS 0.649219f
C12111 DVDD.t0 VSS 0.649219f
C12112 DVDD.t21 VSS 0.480029f
C12113 DVDD.t142 VSS 0.343299f
C12114 DVDD.n1884 VSS 0.500617f
C12115 DVDD.t96 VSS 0.492136f
C12116 DVDD.n1885 VSS 0.504304f
C12117 DVDD.n1886 VSS 0.047318f
C12118 DVDD.n1887 VSS 0.02573f
C12119 DVDD.n1888 VSS 0.037473f
C12120 DVDD.n1889 VSS 0.040423f
C12121 DVDD.n1890 VSS 0.080848f
C12122 DVDD.n1891 VSS 0.080848f
C12123 DVDD.n1892 VSS 0.080848f
C12124 DVDD.n1893 VSS 0.040423f
C12125 DVDD.n1894 VSS 0.037473f
C12126 DVDD.n1895 VSS 0.019073f
C12127 DVDD.n1896 VSS 0.958252f
C12128 DVDD.n1897 VSS 0.169751f
C12129 DVDD.n1898 VSS 0.380569f
C12130 DVDD.n1899 VSS 0.206827f
C12131 DVDD.n1900 VSS 0.214744f
C12132 DVDD.n1901 VSS 0.027577f
C12133 DVDD.n1902 VSS 0.168394f
C12134 DVDD.n1903 VSS 0.206827f
C12135 DVDD.n1904 VSS 0.214744f
C12136 DVDD.n1905 VSS 0.1692f
C12137 DVDD.n1906 VSS 0.168394f
C12138 DVDD.n1907 VSS 0.206827f
C12139 DVDD.n1908 VSS 0.214744f
C12140 DVDD.n1909 VSS 0.1692f
C12141 DVDD.n1910 VSS 0.061774f
C12142 DVDD.n1911 VSS 0.214744f
C12143 DVDD.n1912 VSS 1.0686f
C12144 DVDD.n1913 VSS 0.281047f
C12145 DVDD.n1914 VSS 0.206827f
C12146 DVDD.n1915 VSS 0.214744f
C12147 DVDD.n1916 VSS 0.027577f
C12148 DVDD.n1917 VSS 0.214744f
C12149 DVDD.n1918 VSS 0.281047f
C12150 DVDD.n1919 VSS 1.0686f
C12151 DVDD.n1920 VSS 0.517784f
C12152 DVDD.n1921 VSS 0.022827f
C12153 DVDD.n1922 VSS 0.14181f
C12154 DVDD.n1923 VSS 0.027577f
C12155 DVDD.n1924 VSS 0.037473f
C12156 DVDD.n1925 VSS 0.037473f
C12157 DVDD.n1926 VSS 0.045294f
C12158 DVDD.n1927 VSS 0.073355f
C12159 DVDD.n1928 VSS 0.086693f
C12160 DVDD.n1929 VSS 0.026554f
C12161 DVDD.t118 VSS 0.020584f
C12162 DVDD.t175 VSS 0.020584f
C12163 DVDD.n1930 VSS 0.077533f
C12164 DVDD.t174 VSS 0.299967f
C12165 DVDD.t91 VSS 0.299959f
C12166 DVDD.t92 VSS 0.020584f
C12167 DVDD.t140 VSS 0.020584f
C12168 DVDD.n1931 VSS 0.077533f
C12169 DVDD.n1932 VSS 0.395692f
C12170 DVDD.n1933 VSS 0.130328f
C12171 DVDD.t139 VSS 0.297053f
C12172 DVDD.n1934 VSS 0.353976f
C12173 DVDD.t117 VSS 0.297053f
C12174 DVDD.n1935 VSS 0.130331f
C12175 DVDD.n1936 VSS 0.395744f
C12176 DVDD.n1937 VSS 0.025466f
C12177 DVDD.n1938 VSS 0.171201f
C12178 DVDD.n1939 VSS 1.06722f
C12179 DVDD.n1940 VSS 0.206827f
C12180 DVDD.n1941 VSS 0.281047f
C12181 DVDD.n1942 VSS 0.281047f
C12182 DVDD.n1943 VSS 0.363555f
C12183 DVDD.n1944 VSS 0.517952f
C12184 DVDD.n1945 VSS 0.677237f
C12185 DVDD.n1946 VSS 0.037717f
C12186 DVDD.n1947 VSS 0.033079f
C12187 DVDD.n1948 VSS 0.655388f
C12188 DVDD.n1949 VSS 0.171201f
C12189 DVDD.n1950 VSS 0.36353f
C12190 DVDD.n1951 VSS 0.281047f
C12191 DVDD.n1952 VSS 0.206827f
C12192 DVDD.n1953 VSS 0.206827f
C12193 DVDD.n1954 VSS 0.348732f
C12194 DVDD.n1955 VSS 0.281047f
C12195 DVDD.n1956 VSS 0.363555f
C12196 DVDD.n1957 VSS 0.171201f
C12197 DVDD.t131 VSS 0.299943f
C12198 DVDD.t132 VSS 0.020584f
C12199 DVDD.t149 VSS 0.020584f
C12200 DVDD.n1958 VSS 0.077533f
C12201 DVDD.n1959 VSS 0.399479f
C12202 DVDD.n1960 VSS 0.132913f
C12203 DVDD.t148 VSS 0.297023f
C12204 DVDD.n1961 VSS 0.349495f
C12205 DVDD.t188 VSS 0.020584f
C12206 DVDD.t165 VSS 0.020584f
C12207 DVDD.n1962 VSS 0.077533f
C12208 DVDD.t164 VSS 0.299996f
C12209 DVDD.t187 VSS 0.297053f
C12210 DVDD.n1963 VSS 0.130274f
C12211 DVDD.n1964 VSS 0.394659f
C12212 DVDD.n1965 VSS 0.028936f
C12213 DVDD.n1966 VSS 0.050816f
C12214 DVDD.n1967 VSS 0.706313f
C12215 DVDD.n1968 VSS 0.517952f
C12216 DVDD.n1969 VSS 1.06722f
C12217 DVDD.n1970 VSS 0.281047f
C12218 DVDD.n1971 VSS 0.206827f
C12219 DVDD.n1972 VSS 0.206827f
C12220 DVDD.n1973 VSS 0.214744f
C12221 DVDD.n1974 VSS 0.214744f
C12222 DVDD.n1975 VSS 0.040423f
C12223 DVDD.n1976 VSS 0.080848f
C12224 DVDD.n1977 VSS 0.080848f
C12225 DVDD.n1978 VSS 0.040423f
C12226 DVDD.n1979 VSS 0.037473f
C12227 DVDD.n1980 VSS 0.040423f
C12228 DVDD.n1982 VSS 0.292822f
C12229 DVDD.n1983 VSS 0.065578f
C12230 DVDD.n1984 VSS 0.037473f
C12231 DVDD.n1985 VSS 0.037473f
C12232 DVDD.n1986 VSS 0.037473f
C12233 DVDD.n1987 VSS 0.037473f
C12234 DVDD.n1988 VSS 0.073429f
C12235 DVDD.n1990 VSS 0.037473f
C12236 DVDD.n1992 VSS 0.037473f
C12237 DVDD.n1994 VSS 0.037473f
C12238 DVDD.n1996 VSS 0.037473f
C12239 DVDD.n1997 VSS 0.065578f
C12240 DVDD.n1999 VSS 0.065578f
C12241 DVDD.n2000 VSS 0.037473f
C12242 DVDD.n2001 VSS 0.037473f
C12243 DVDD.n2002 VSS 0.037473f
C12244 DVDD.n2003 VSS 0.037473f
C12245 DVDD.n2004 VSS 0.073429f
C12246 DVDD.n2006 VSS 0.037473f
C12247 DVDD.n2008 VSS 0.037473f
C12248 DVDD.n2010 VSS 0.037473f
C12249 DVDD.n2012 VSS 0.037473f
C12250 DVDD.t222 VSS 0.143902f
C12251 DVDD.n2013 VSS 0.065267f
C12252 DVDD.n2014 VSS 0.229669f
C12253 DVDD.t209 VSS 0.143902f
C12254 DVDD.n2015 VSS 0.075241f
C12255 DVDD.n2016 VSS 0.075241f
C12256 DVDD.n2017 VSS 0.106877f
C12257 DVDD.n2018 VSS 0.106877f
C12258 DVDD.t219 VSS 0.143902f
C12259 DVDD.n2019 VSS 0.075241f
C12260 DVDD.n2020 VSS 0.075241f
C12261 DVDD.n2021 VSS 0.106877f
C12262 DVDD.n2022 VSS 0.106877f
C12263 DVDD.t207 VSS 0.143902f
C12264 DVDD.n2023 VSS 0.075241f
C12265 DVDD.n2024 VSS 0.075241f
C12266 DVDD.n2025 VSS 0.106877f
C12267 DVDD.n2026 VSS 0.106877f
C12268 DVDD.t218 VSS 0.143902f
C12269 DVDD.n2027 VSS 0.075241f
C12270 DVDD.n2028 VSS 0.075241f
C12271 DVDD.n2029 VSS 0.106877f
C12272 DVDD.n2030 VSS 0.106877f
C12273 DVDD.t211 VSS 0.143902f
C12274 DVDD.n2031 VSS 0.075241f
C12275 DVDD.n2032 VSS 0.075241f
C12276 DVDD.n2033 VSS 0.106877f
C12277 DVDD.n2034 VSS 0.106877f
C12278 DVDD.t221 VSS 0.143902f
C12279 DVDD.n2035 VSS 0.075241f
C12280 DVDD.n2036 VSS 0.075241f
C12281 DVDD.n2037 VSS 0.147758f
C12282 DVDD.n2038 VSS 0.086802f
C12283 DVDD.t208 VSS 0.143902f
C12284 DVDD.n2039 VSS 0.250567f
C12285 DVDD.n2043 VSS 0.131155f
C12286 DVDD.n2044 VSS 0.131155f
C12287 DVDD.n2045 VSS 0.131155f
C12288 DVDD.n2046 VSS 0.131155f
C12289 DVDD.n2047 VSS 0.131155f
C12290 DVDD.n2048 VSS 0.131155f
C12291 DVDD.n2049 VSS 0.131155f
C12292 DVDD.n2050 VSS 0.131155f
C12293 DVDD.n2051 VSS 0.131155f
C12294 DVDD.n2052 VSS 0.131155f
C12295 DVDD.n2053 VSS 0.131155f
C12296 DVDD.n2054 VSS 0.089971f
C12297 DVDD.n2055 VSS 0.131155f
C12298 DVDD.n2056 VSS 0.131155f
C12299 DVDD.n2057 VSS 0.131155f
C12300 DVDD.n2058 VSS 0.06881f
C12301 DVDD.n2059 VSS 0.113145f
C12302 DVDD.n2060 VSS -0.005459f
C12303 DVDD.t67 VSS 0.233913f
C12304 DVDD.n2061 VSS 0.018243f
C12305 DVDD.n2062 VSS 0.08405f
C12306 DVDD.n2063 VSS 0.08556f
C12307 DVDD.n2064 VSS 0.131155f
C12308 DVDD.n2065 VSS 0.131155f
C12309 DVDD.n2066 VSS 0.131155f
C12310 DVDD.n2067 VSS 0.131155f
C12311 DVDD.n2068 VSS 0.084512f
C12312 DVDD.n2069 VSS 0.131155f
C12313 DVDD.n2070 VSS 0.131155f
C12314 DVDD.n2071 VSS 0.131155f
C12315 DVDD.n2072 VSS 0.131155f
C12316 DVDD.t173 VSS 0.010292f
C12317 DVDD.t112 VSS 0.010292f
C12318 DVDD.n2073 VSS 0.022718f
C12319 DVDD.n2074 VSS 0.049968f
C12320 DVDD.n2075 VSS 0.085561f
C12321 DVDD.n2076 VSS 0.112221f
C12322 DVDD.n2077 VSS 0.131155f
C12323 DVDD.n2078 VSS 0.131155f
C12324 DVDD.n2079 VSS 0.131155f
C12325 DVDD.n2080 VSS 0.131155f
C12326 DVDD.n2081 VSS 0.131155f
C12327 DVDD.n2082 VSS 0.131155f
C12328 DVDD.n2083 VSS 0.131155f
C12329 DVDD.n2084 VSS 0.016247f
C12330 DVDD.t114 VSS 0.02622f
C12331 DVDD.n2085 VSS 0.060717f
C12332 DVDD.n2086 VSS 0.08556f
C12333 DVDD.n2087 VSS 0.075276f
C12334 DVDD.n2088 VSS 0.131155f
C12335 DVDD.n2089 VSS 0.131155f
C12336 DVDD.n2090 VSS 0.131155f
C12337 DVDD.n2091 VSS 0.131155f
C12338 DVDD.n2092 VSS 0.131155f
C12339 DVDD.n2093 VSS 0.084512f
C12340 DVDD.n2094 VSS 0.085561f
C12341 DVDD.n2095 VSS 0.131155f
C12342 DVDD.n2096 VSS 0.131155f
C12343 DVDD.n2097 VSS 0.131155f
C12344 DVDD.n2098 VSS 0.121457f
C12345 DVDD.n2099 VSS 0.086821f
C12346 DVDD.n2100 VSS 0.131155f
C12347 DVDD.n2101 VSS 0.131155f
C12348 DVDD.n2102 VSS 0.131155f
C12349 DVDD.n2103 VSS 0.131155f
C12350 DVDD.n2104 VSS 0.131155f
C12351 DVDD.n2105 VSS 0.131155f
C12352 DVDD.n2106 VSS 0.131155f
C12353 DVDD.n2107 VSS 0.131155f
C12354 DVDD.n2108 VSS 0.131155f
C12355 DVDD.n2109 VSS 0.131155f
C12356 DVDD.n2110 VSS 0.131155f
C12357 DVDD.n2111 VSS 0.131155f
C12358 DVDD.n2112 VSS 0.131155f
C12359 DVDD.n2113 VSS 0.131155f
C12360 DVDD.n2114 VSS 0.131155f
C12361 DVDD.n2115 VSS 0.131155f
C12362 DVDD.n2116 VSS 0.131155f
C12363 DVDD.n2117 VSS 0.131155f
C12364 DVDD.n2118 VSS 0.123305f
C12365 DVDD.n2119 VSS 0.131155f
C12366 DVDD.n2120 VSS 0.131155f
C12367 DVDD.n2121 VSS 0.131155f
C12368 DVDD.n2122 VSS 0.089971f
C12369 DVDD.n2123 VSS 0.117763f
C12370 DVDD.n2124 VSS -0.005459f
C12371 DVDD.t193 VSS 0.233913f
C12372 DVDD.n2125 VSS 0.018243f
C12373 DVDD.n2126 VSS 0.08405f
C12374 DVDD.n2127 VSS 0.08556f
C12375 DVDD.n2128 VSS 0.131155f
C12376 DVDD.n2129 VSS 0.131155f
C12377 DVDD.n2130 VSS 0.131155f
C12378 DVDD.n2131 VSS 0.131155f
C12379 DVDD.n2132 VSS 0.08913f
C12380 DVDD.n2133 VSS 0.131155f
C12381 DVDD.n2134 VSS 0.131155f
C12382 DVDD.n2135 VSS 0.131155f
C12383 DVDD.n2136 VSS 0.131155f
C12384 DVDD.n2137 VSS 0.131155f
C12385 DVDD.n2138 VSS 0.131155f
C12386 DVDD.t147 VSS 0.010292f
C12387 DVDD.t56 VSS 0.010292f
C12388 DVDD.n2139 VSS 0.022718f
C12389 DVDD.n2140 VSS 0.049968f
C12390 DVDD.n2141 VSS 0.085561f
C12391 DVDD.n2142 VSS 0.107603f
C12392 DVDD.n2143 VSS 0.131155f
C12393 DVDD.n2144 VSS 0.131155f
C12394 DVDD.n2145 VSS 0.131155f
C12395 DVDD.n2146 VSS 0.131155f
C12396 DVDD.n2147 VSS 0.131155f
C12397 DVDD.n2148 VSS 0.131155f
C12398 DVDD.n2149 VSS 0.131155f
C12399 DVDD.n2150 VSS 0.016247f
C12400 DVDD.t50 VSS 0.02622f
C12401 DVDD.n2151 VSS 0.060717f
C12402 DVDD.n2152 VSS 0.08556f
C12403 DVDD.n2153 VSS 0.070658f
C12404 DVDD.n2154 VSS 0.131155f
C12405 DVDD.n2155 VSS 0.131155f
C12406 DVDD.n2156 VSS 0.131155f
C12407 DVDD.n2157 VSS 0.131155f
C12408 DVDD.n2158 VSS 0.131155f
C12409 DVDD.n2159 VSS 0.08913f
C12410 DVDD.n2160 VSS 0.085561f
C12411 DVDD.n2161 VSS 0.131155f
C12412 DVDD.n2162 VSS 0.131155f
C12413 DVDD.n2163 VSS 0.131155f
C12414 DVDD.n2164 VSS 0.126075f
C12415 DVDD.n2165 VSS 0.086821f
C12416 DVDD.n2166 VSS 0.131155f
C12417 DVDD.n2167 VSS 0.131155f
C12418 DVDD.n2168 VSS 0.131155f
C12419 DVDD.n2169 VSS 0.131155f
C12420 DVDD.n2170 VSS 0.131155f
C12421 DVDD.n2171 VSS 0.131155f
C12422 DVDD.n2172 VSS 0.131155f
C12423 DVDD.n2173 VSS 0.131155f
C12424 DVDD.n2174 VSS 0.131155f
C12425 DVDD.n2175 VSS 0.131155f
C12426 DVDD.n2176 VSS 0.131155f
C12427 DVDD.n2177 VSS 0.131155f
C12428 DVDD.n2178 VSS 0.131155f
C12429 DVDD.n2179 VSS 0.131155f
C12430 DVDD.n2180 VSS 0.131155f
C12431 DVDD.n2181 VSS 0.131155f
C12432 DVDD.n2182 VSS 0.131155f
C12433 DVDD.n2183 VSS 0.131155f
C12434 DVDD.n2184 VSS 0.131155f
C12435 DVDD.n2185 VSS 0.131155f
C12436 DVDD.n2186 VSS 0.131155f
C12437 DVDD.n2187 VSS 0.131155f
C12438 DVDD.n2188 VSS 0.131155f
C12439 DVDD.n2189 VSS 0.131155f
C12440 DVDD.n2190 VSS 0.131155f
C12441 DVDD.n2191 VSS 0.131155f
C12442 DVDD.n2192 VSS 0.131155f
C12443 DVDD.n2193 VSS 0.131155f
C12444 DVDD.n2194 VSS 0.131155f
C12445 DVDD.n2195 VSS 0.118225f
C12446 DVDD.n2196 VSS 0.067425f
C12447 DVDD.n2197 VSS 0.172652f
C12448 DVDD.n2198 VSS 0.63196f
C12449 DVDD.n2199 VSS 0.096981f
C12450 DVDD.t206 VSS 0.143902f
C12451 DVDD.n2200 VSS 0.08914f
C12452 DVDD.t212 VSS 0.143902f
C12453 DVDD.n2201 VSS 0.079113f
C12454 DVDD.n2202 VSS 0.202208f
C12455 DVDD.n2203 VSS 0.147146f
C12456 DVDD.n2204 VSS 0.086821f
C12457 DVDD.n2205 VSS 0.131155f
C12458 DVDD.n2206 VSS 0.131155f
C12459 DVDD.n2207 VSS 0.131155f
C12460 DVDD.n2208 VSS 0.131155f
C12461 DVDD.n2209 VSS 0.131155f
C12462 DVDD.n2210 VSS 0.131155f
C12463 DVDD.n2211 VSS 0.131155f
C12464 DVDD.n2212 VSS 0.131155f
C12465 DVDD.n2213 VSS 0.131155f
C12466 DVDD.n2214 VSS 0.131155f
C12467 DVDD.n2215 VSS 0.131155f
C12468 DVDD.n2216 VSS 0.131155f
C12469 DVDD.n2217 VSS 0.131155f
C12470 DVDD.n2218 VSS 0.131155f
C12471 DVDD.n2219 VSS 0.131155f
C12472 DVDD.n2220 VSS 0.131155f
C12473 DVDD.n2221 VSS 0.131155f
C12474 DVDD.n2222 VSS 0.131155f
C12475 DVDD.n2223 VSS 0.131155f
C12476 DVDD.n2224 VSS 0.131155f
C12477 DVDD.n2225 VSS 0.131155f
C12478 DVDD.n2226 VSS 0.131155f
C12479 DVDD.n2227 VSS 0.131155f
C12480 DVDD.n2228 VSS 0.131155f
C12481 DVDD.n2229 VSS 0.131155f
C12482 DVDD.n2230 VSS 0.131155f
C12483 DVDD.n2231 VSS 0.131155f
C12484 DVDD.n2232 VSS 0.131155f
C12485 DVDD.n2233 VSS 0.131155f
C12486 DVDD.n2234 VSS 0.131155f
C12487 DVDD.n2235 VSS 0.131155f
C12488 DVDD.n2236 VSS 0.131155f
C12489 DVDD.n2237 VSS 0.131155f
C12490 DVDD.n2238 VSS 0.131155f
C12491 DVDD.n2239 VSS 0.131155f
C12492 DVDD.n2240 VSS 0.131155f
C12493 DVDD.n2241 VSS 0.131155f
C12494 DVDD.n2242 VSS 0.131155f
C12495 DVDD.n2243 VSS 0.131155f
C12496 DVDD.n2244 VSS 0.131155f
C12497 DVDD.n2245 VSS 0.131155f
C12498 DVDD.n2246 VSS 0.131155f
C12499 DVDD.n2247 VSS 0.131155f
C12500 DVDD.n2248 VSS 0.131155f
C12501 DVDD.n2249 VSS 0.131155f
C12502 DVDD.n2250 VSS 0.131155f
C12503 DVDD.n2251 VSS 0.131155f
C12504 DVDD.n2252 VSS 0.131155f
C12505 DVDD.n2253 VSS 0.131155f
C12506 DVDD.n2254 VSS 0.131155f
C12507 DVDD.n2255 VSS 0.131155f
C12508 DVDD.n2256 VSS 0.131155f
C12509 DVDD.n2257 VSS 0.131155f
C12510 DVDD.n2258 VSS 0.076199f
C12511 DVDD.n2259 VSS 0.089971f
C12512 DVDD.n2260 VSS 0.24033f
C12513 DVDD.t62 VSS 0.156654f
C12514 DVDD.t77 VSS 0.235776f
C12515 DVDD.t59 VSS 0.1558f
C12516 DVDD.n2261 VSS 0.070782f
C12517 DVDD.t63 VSS 0.010292f
C12518 DVDD.t60 VSS 0.010292f
C12519 DVDD.n2262 VSS 0.022718f
C12520 DVDD.n2263 VSS 0.049968f
C12521 DVDD.t194 VSS 0.02622f
C12522 DVDD.n2264 VSS 0.060717f
C12523 DVDD.n2265 VSS 0.016247f
C12524 DVDD.n2266 VSS -0.005459f
C12525 DVDD.n2267 VSS 0.035625f
C12526 DVDD.t78 VSS 0.026135f
C12527 DVDD.n2268 VSS 0.060979f
C12528 DVDD.n2269 VSS 0.085666f
C12529 DVDD.n2270 VSS 0.09929f
C12530 DVDD.n2271 VSS 0.131155f
C12531 DVDD.n2272 VSS 0.131155f
C12532 DVDD.n2273 VSS 0.131155f
C12533 DVDD.n2274 VSS 0.131155f
C12534 DVDD.n2275 VSS 0.131155f
C12535 DVDD.n2276 VSS 0.131155f
C12536 DVDD.n2277 VSS 0.070658f
C12537 DVDD.n2278 VSS 0.131155f
C12538 DVDD.n2279 VSS 0.131155f
C12539 DVDD.n2280 VSS 0.131155f
C12540 DVDD.n2281 VSS 0.131155f
C12541 DVDD.n2282 VSS 0.131155f
C12542 DVDD.n2283 VSS 0.131155f
C12543 DVDD.n2284 VSS 0.131155f
C12544 DVDD.n2285 VSS 0.08405f
C12545 DVDD.n2286 VSS 0.089971f
C12546 DVDD.n2287 VSS 0.028611f
C12547 DVDD.n2288 VSS 0.228945f
C12548 DVDD.t49 VSS 0.233913f
C12549 DVDD.t55 VSS 0.156654f
C12550 DVDD.n2289 VSS 0.070782f
C12551 DVDD.t146 VSS 0.1558f
C12552 DVDD.t168 VSS 0.235776f
C12553 DVDD.n2290 VSS 0.24033f
C12554 DVDD.n2291 VSS 0.035457f
C12555 DVDD.t169 VSS 0.02622f
C12556 DVDD.n2292 VSS 0.060717f
C12557 DVDD.n2293 VSS 0.08556f
C12558 DVDD.n2294 VSS 0.07897f
C12559 DVDD.n2295 VSS 0.073429f
C12560 DVDD.n2296 VSS 0.131155f
C12561 DVDD.n2297 VSS 0.131155f
C12562 DVDD.n2298 VSS 0.131155f
C12563 DVDD.n2299 VSS 0.131155f
C12564 DVDD.n2300 VSS 0.131155f
C12565 DVDD.n2301 VSS 0.131155f
C12566 DVDD.n2302 VSS 0.131155f
C12567 DVDD.n2303 VSS 0.131155f
C12568 DVDD.n2304 VSS 0.131155f
C12569 DVDD.n2305 VSS 0.131155f
C12570 DVDD.n2306 VSS 0.131155f
C12571 DVDD.n2307 VSS 0.131155f
C12572 DVDD.n2308 VSS 0.131155f
C12573 DVDD.n2309 VSS 0.131155f
C12574 DVDD.n2310 VSS 0.131155f
C12575 DVDD.n2311 VSS 0.131155f
C12576 DVDD.n2312 VSS 0.131155f
C12577 DVDD.n2313 VSS 0.131155f
C12578 DVDD.n2314 VSS 0.131155f
C12579 DVDD.n2315 VSS 0.131155f
C12580 DVDD.n2316 VSS 0.131155f
C12581 DVDD.n2317 VSS 0.131155f
C12582 DVDD.n2318 VSS 0.131155f
C12583 DVDD.n2319 VSS 0.131155f
C12584 DVDD.n2320 VSS 0.131155f
C12585 DVDD.n2321 VSS 0.131155f
C12586 DVDD.n2322 VSS 0.131155f
C12587 DVDD.n2323 VSS 0.131155f
C12588 DVDD.n2324 VSS 0.131155f
C12589 DVDD.n2325 VSS 0.131155f
C12590 DVDD.n2326 VSS 0.131155f
C12591 DVDD.n2327 VSS 0.131155f
C12592 DVDD.n2328 VSS 0.131155f
C12593 DVDD.n2329 VSS 0.131155f
C12594 DVDD.n2330 VSS 0.131155f
C12595 DVDD.n2331 VSS 0.131155f
C12596 DVDD.n2332 VSS 0.131155f
C12597 DVDD.n2333 VSS 0.071581f
C12598 DVDD.n2334 VSS 0.089971f
C12599 DVDD.n2335 VSS 0.24033f
C12600 DVDD.t162 VSS 0.156654f
C12601 DVDD.t133 VSS 0.235776f
C12602 DVDD.t166 VSS 0.1558f
C12603 DVDD.n2336 VSS 0.070782f
C12604 DVDD.t163 VSS 0.010292f
C12605 DVDD.t167 VSS 0.010292f
C12606 DVDD.n2337 VSS 0.022718f
C12607 DVDD.n2338 VSS 0.049968f
C12608 DVDD.t68 VSS 0.02622f
C12609 DVDD.n2339 VSS 0.060717f
C12610 DVDD.n2340 VSS 0.016247f
C12611 DVDD.n2341 VSS -0.005459f
C12612 DVDD.n2342 VSS 0.035457f
C12613 DVDD.t134 VSS 0.02622f
C12614 DVDD.n2343 VSS 0.060717f
C12615 DVDD.n2344 VSS 0.08556f
C12616 DVDD.n2345 VSS 0.103908f
C12617 DVDD.n2346 VSS 0.131155f
C12618 DVDD.n2347 VSS 0.131155f
C12619 DVDD.n2348 VSS 0.131155f
C12620 DVDD.n2349 VSS 0.131155f
C12621 DVDD.n2350 VSS 0.131155f
C12622 DVDD.n2351 VSS 0.131155f
C12623 DVDD.n2352 VSS 0.075276f
C12624 DVDD.n2353 VSS 0.131155f
C12625 DVDD.n2354 VSS 0.131155f
C12626 DVDD.n2355 VSS 0.131155f
C12627 DVDD.n2356 VSS 0.131155f
C12628 DVDD.n2357 VSS 0.131155f
C12629 DVDD.n2358 VSS 0.131155f
C12630 DVDD.n2359 VSS 0.131155f
C12631 DVDD.n2360 VSS 0.08405f
C12632 DVDD.n2361 VSS 0.089971f
C12633 DVDD.n2362 VSS 0.028611f
C12634 DVDD.n2363 VSS 0.228945f
C12635 DVDD.t113 VSS 0.233913f
C12636 DVDD.t111 VSS 0.156654f
C12637 DVDD.n2364 VSS 0.070782f
C12638 DVDD.t172 VSS 0.1558f
C12639 DVDD.t129 VSS 0.235776f
C12640 DVDD.n2365 VSS 0.24033f
C12641 DVDD.n2366 VSS 0.035457f
C12642 DVDD.t130 VSS 0.02622f
C12643 DVDD.n2367 VSS 0.060717f
C12644 DVDD.n2368 VSS 0.08556f
C12645 DVDD.n2369 VSS 0.083589f
C12646 DVDD.n2370 VSS 0.131155f
C12647 DVDD.n2371 VSS 0.131155f
C12648 DVDD.n2372 VSS 0.131155f
C12649 DVDD.n2373 VSS 0.131155f
C12650 DVDD.n2374 VSS 0.131155f
C12651 DVDD.n2375 VSS 0.127923f
C12652 DVDD.n2376 VSS 0.131155f
C12653 DVDD.n2377 VSS 0.131155f
C12654 DVDD.n2378 VSS 0.131155f
C12655 DVDD.n2379 VSS 0.131155f
C12656 DVDD.n2380 VSS 0.131155f
C12657 DVDD.n2381 VSS 0.131155f
C12658 DVDD.n2382 VSS 0.131155f
C12659 DVDD.n2383 VSS 0.131155f
C12660 DVDD.n2384 VSS 0.131155f
C12661 DVDD.n2385 VSS 0.131155f
C12662 DVDD.n2386 VSS 0.131155f
C12663 DVDD.n2387 VSS 0.131155f
C12664 DVDD.n2388 VSS 0.131155f
C12665 DVDD.n2389 VSS 0.131155f
C12666 DVDD.n2390 VSS 0.131155f
C12667 DVDD.n2391 VSS 0.131155f
C12668 DVDD.n2392 VSS 0.131155f
C12669 DVDD.n2393 VSS 0.131155f
C12670 DVDD.n2394 VSS 0.131155f
C12671 DVDD.n2395 VSS 0.131155f
C12672 DVDD.n2396 VSS 0.131155f
C12673 DVDD.n2397 VSS 0.485997f
C12674 DVDD.n2398 VSS 0.131155f
C12675 DVDD.n2399 VSS 0.131155f
C12676 DVDD.n2400 VSS 0.065578f
C12677 DVDD.n2401 VSS 0.292822f
C12678 DVDD.n2403 VSS 0.265984f
C12679 DVDD.n2404 VSS 0.065578f
C12680 DVDD.n2405 VSS 0.923125f
C12681 DVDD.n2406 VSS 0.131155f
C12682 DVDD.n2407 VSS 0.131155f
C12683 DVDD.n2408 VSS 0.131155f
C12684 DVDD.n2409 VSS 0.131155f
C12685 DVDD.n2410 VSS 0.131155f
C12686 DVDD.n2411 VSS 0.131155f
C12687 DVDD.n2412 VSS 0.131155f
C12688 DVDD.n2413 VSS 0.131155f
C12689 DVDD.n2414 VSS 0.131155f
C12690 DVDD.n2415 VSS 0.131155f
C12691 DVDD.n2416 VSS 0.131155f
C12692 DVDD.n2417 VSS 0.131155f
C12693 DVDD.n2418 VSS 0.131155f
C12694 DVDD.n2419 VSS 0.131155f
C12695 DVDD.n2420 VSS 0.131155f
C12696 DVDD.n2421 VSS 0.131155f
C12697 DVDD.n2422 VSS 0.131155f
C12698 DVDD.n2423 VSS 0.131155f
C12699 DVDD.n2424 VSS 0.131155f
C12700 DVDD.n2425 VSS 0.131155f
C12701 DVDD.n2426 VSS 0.131155f
C12702 DVDD.n2427 VSS 0.131155f
C12703 DVDD.n2428 VSS 0.131155f
C12704 DVDD.n2429 VSS 0.131155f
C12705 DVDD.t110 VSS 0.026836f
C12706 DVDD.t109 VSS 0.297789f
C12707 DVDD.n2430 VSS 0.27409f
C12708 DVDD.n2431 VSS 0.05429f
C12709 DVDD.n2432 VSS 0.056574f
C12710 DVDD.n2433 VSS 0.081547f
C12711 DVDD.n2434 VSS 0.131155f
C12712 DVDD.n2435 VSS 0.131155f
C12713 DVDD.n2436 VSS 0.131155f
C12714 DVDD.n2437 VSS 0.077585f
C12715 DVDD.n2438 VSS 0.073429f
C12716 DVDD.n2439 VSS 0.131155f
C12717 DVDD.n2440 VSS 0.131155f
C12718 DVDD.n2441 VSS 0.131155f
C12719 DVDD.n2442 VSS 0.065578f
C12720 DVDD.n2443 VSS 0.01311f
C12721 DVDD.n2444 VSS 0.01311f
C12722 DVDD.n2445 VSS 0.01311f
C12723 DVDD.n2446 VSS 0.01311f
C12724 DVDD.n2447 VSS 0.01311f
C12725 DVDD.n2448 VSS 0.065578f
C12726 DVDD.n2449 VSS 0.01311f
C12727 DVDD.n2450 VSS 0.01311f
C12728 DVDD.n2451 VSS 0.01311f
C12729 DVDD.n2452 VSS 0.01311f
C12730 DVDD.n2453 VSS -0.348668f
C12731 DVDD.n2454 VSS 0.017238f
C12732 DVDD.n2455 VSS 0.131155f
C12733 DVDD.n2456 VSS 0.131155f
C12734 DVDD.n2457 VSS 0.131155f
C12735 DVDD.n2458 VSS 0.131155f
C12736 DVDD.n2459 VSS 0.131155f
C12737 DVDD.n2460 VSS 0.131155f
C12738 DVDD.n2461 VSS 0.131155f
C12739 DVDD.n2462 VSS 0.131155f
C12740 DVDD.n2463 VSS 0.131155f
C12741 DVDD.n2464 VSS 0.131155f
C12742 DVDD.n2465 VSS 0.131155f
C12743 DVDD.n2466 VSS 0.131155f
C12744 DVDD.n2467 VSS 0.131155f
C12745 DVDD.n2468 VSS 0.131155f
C12746 DVDD.n2469 VSS 0.131155f
C12747 DVDD.n2470 VSS 0.131155f
C12748 DVDD.n2471 VSS 0.131155f
C12749 DVDD.n2472 VSS 0.131155f
C12750 DVDD.n2473 VSS 0.131155f
C12751 DVDD.n2474 VSS 0.131155f
C12752 DVDD.n2475 VSS 0.131155f
C12753 DVDD.n2476 VSS 0.131155f
C12754 DVDD.n2477 VSS 0.131155f
C12755 DVDD.n2478 VSS 0.131155f
C12756 DVDD.n2479 VSS 0.131155f
C12757 DVDD.n2480 VSS 0.131155f
C12758 DVDD.n2481 VSS 0.131155f
C12759 DVDD.n2482 VSS 0.131155f
C12760 DVDD.n2483 VSS 0.131155f
C12761 DVDD.n2484 VSS 0.131155f
C12762 DVDD.n2485 VSS 0.131155f
C12763 DVDD.n2486 VSS 0.131155f
C12764 DVDD.n2487 VSS 0.131155f
C12765 DVDD.n2488 VSS 0.131155f
C12766 DVDD.n2489 VSS 0.131155f
C12767 DVDD.n2490 VSS 0.131155f
C12768 DVDD.n2491 VSS 0.031743f
C12769 DVDD.n2492 VSS 0.01425f
C12770 DVDD.n2493 VSS 0.01425f
C12771 DVDD.n2494 VSS 0.01425f
C12772 DVDD.n2495 VSS 0.065578f
C12773 DVDD.n2496 VSS 0.01425f
C12774 DVDD.n2497 VSS 0.01425f
C12775 DVDD.n2498 VSS 0.01425f
C12776 DVDD.n2499 VSS 0.027445f
C12777 DVDD.n2500 VSS 0.065578f
C12778 DVDD.n2501 VSS 0.004458f
C12779 DVDD.n2502 VSS 0.032723f
C12780 DVDD.n2503 VSS 0.030105f
C12781 DVDD.n2504 VSS 0.032723f
C12782 DVDD.n2505 VSS 0.021608f
C12783 DVDD.n2507 VSS 0.180438f
C12784 DVDD.n2508 VSS 0.021608f
C12785 DVDD.n2509 VSS 0.032723f
C12786 DVDD.n2510 VSS 0.11263f
C12787 DVDD.n2511 VSS 0.65561f
C12788 DVDD.t182 VSS 0.0102f
C12789 DVDD.n2512 VSS 0.032309f
C12790 DVDD.n2513 VSS 0.116121f
C12791 DVDD.t11 VSS 0.006518f
C12792 DVDD.t24 VSS 0.006518f
C12793 DVDD.n2514 VSS 0.019862f
C12794 DVDD.t9 VSS 0.009408f
C12795 DVDD.t192 VSS 0.006861f
C12796 DVDD.t13 VSS 0.006861f
C12797 DVDD.n2515 VSS 0.029349f
C12798 DVDD.n2516 VSS 0.049378f
C12799 DVDD.t54 VSS 0.016195f
C12800 DVDD.n2517 VSS 0.029042f
C12801 DVDD.n2518 VSS 0.043596f
C12802 DVDD.n2519 VSS 0.143921f
C12803 DVDD.t94 VSS 0.182006f
C12804 DVDD.n2520 VSS 0.111624f
C12805 DVDD.t95 VSS 0.0131f
C12806 DVDD.n2521 VSS 0.324777f
C12807 DVDD.n2522 VSS 0.279548f
C12808 DVDD.n2523 VSS 0.305779f
C12809 DVDD.t141 VSS 0.361167f
C12810 DVDD.t204 VSS 0.495145f
C12811 DVDD.t18 VSS 0.433678f
C12812 DVDD.t17 VSS 0.269768f
C12813 DVDD.t2 VSS 0.269768f
C12814 DVDD.t3 VSS 0.370505f
C12815 DVDD.t10 VSS 0.346601f
C12816 DVDD.n2524 VSS 0.07465f
C12817 DVDD.n2525 VSS 0.047343f
C12818 DVDD.n2526 VSS 0.047343f
C12819 DVDD.n2527 VSS 0.035052f
C12820 DVDD.n2528 VSS 0.047343f
C12821 DVDD.n2530 VSS 0.047343f
C12822 DVDD.n2531 VSS 0.023671f
C12823 DVDD.n2532 VSS 0.08948f
C12824 DVDD.n2533 VSS 0.047343f
C12825 DVDD.n2538 VSS 0.063261f
C12826 DVDD.t52 VSS 0.051913f
C12827 DVDD.t48 VSS 0.051913f
C12828 DVDD.t58 VSS 0.016195f
C12829 DVDD.n2539 VSS 0.046465f
C12830 DVDD.n2540 VSS 0.045624f
C12831 DVDD.n2541 VSS 0.045391f
C12832 DVDD.n2542 VSS 0.063261f
C12833 DVDD.n2545 VSS 0.034304f
C12834 DVDD.n2547 VSS 0.07465f
C12835 DVDD.n2548 VSS 0.053518f
C12836 DVDD.n2549 VSS 0.053518f
C12837 DVDD.n2550 VSS 0.053518f
C12838 DVDD.n2551 VSS 0.053518f
C12839 DVDD.n2553 VSS 0.053518f
C12840 DVDD.n2554 VSS 0.053518f
C12841 DVDD.n2556 VSS 0.063261f
C12842 DVDD.n2557 VSS 0.063261f
C12843 DVDD.n2560 VSS 0.063261f
C12844 DVDD.n2564 VSS 0.063261f
C12845 DVDD.n2569 VSS 0.187266f
C12846 DVDD.n2573 VSS 0.044255f
C12847 DVDD.n2574 VSS 0.063261f
C12848 DVDD.n2575 VSS 0.07559f
C12849 DVDD.n2576 VSS 0.07465f
C12850 DVDD.n2577 VSS 0.07465f
C12851 DVDD.n2578 VSS 0.07465f
C12852 DVDD.n2579 VSS 0.07465f
C12853 DVDD.n2580 VSS 0.063261f
C12854 DVDD.n2581 VSS 0.044255f
C12855 DVDD.n2582 VSS 0.063261f
C12856 DVDD.n2583 VSS 0.07465f
C12857 DVDD.n2584 VSS 0.07465f
C12858 DVDD.n2588 VSS 0.063261f
C12859 DVDD.n2589 VSS 0.07465f
C12860 DVDD.n2590 VSS 0.07465f
C12861 DVDD.n2591 VSS 0.063261f
C12862 DVDD.n2592 VSS 0.048889f
C12863 DVDD.n2593 VSS 0.059003f
C12864 DVDD.n2594 VSS 0.098178f
C12865 DVDD.n2595 VSS 0.23825f
C12866 DVDD.t51 VSS 0.2579f
C12867 DVDD.t47 VSS 0.49907f
C12868 DVDD.t57 VSS 0.516487f
C12869 DVDD.t53 VSS 0.297087f
C12870 DVDD.t8 VSS 0.297087f
C12871 DVDD.t12 VSS 0.208302f
C12872 DVDD.t191 VSS 0.301355f
C12873 DVDD.t23 VSS 0.221108f
C12874 DVDD.n2596 VSS 0.104151f
C12875 DVDD.n2597 VSS 0.300925f
C12876 DVDD.n2598 VSS 0.029808f
C12877 DVDD.n2599 VSS 0.079246f
C12878 DVDD.n2600 VSS 0.063461f
C12879 DVDD.n2601 VSS 0.321965f
C12880 DVDD.n2602 VSS -0.571949f
C12881 DVDD.n2603 VSS 0.524053f
C12882 DVDD.n2604 VSS 0.320714f
C12883 DVDD.n2605 VSS 0.016995f
C12884 DVDD.n2607 VSS 0.127857f
C12885 DVDD.n2608 VSS 0.031562f
C12886 DVDD.n2609 VSS 0.032723f
C12887 DVDD.n2610 VSS 0.032723f
C12888 DVDD.n2611 VSS 0.032723f
C12889 DVDD.n2612 VSS 0.030105f
C12890 DVDD.n2613 VSS 0.030105f
C12891 DVDD.n2614 VSS 0.030105f
C12892 DVDD.n2615 VSS 0.032723f
C12893 DVDD.n2616 VSS 0.032723f
C12894 DVDD.n2617 VSS 0.032723f
C12895 DVDD.n2618 VSS 0.030105f
C12896 DVDD.n2619 VSS 0.030105f
C12897 DVDD.n2620 VSS 0.030105f
C12898 DVDD.n2621 VSS 0.032723f
C12899 DVDD.n2622 VSS 0.032723f
C12900 DVDD.n2623 VSS 0.038265f
C12901 DVDD.n2624 VSS -0.734197f
C12902 DVDD.n2625 VSS 0.033261f
C12903 DVDD.n2626 VSS 0.017238f
C12904 DVDD.n2628 VSS 0.026221f
C12905 DVDD.n2629 VSS 0.017238f
C12906 DVDD.n2630 VSS 0.026221f
C12907 DVDD.n2631 VSS 0.026221f
C12908 DVDD.n2632 VSS 0.016024f
C12909 DVDD.n2633 VSS 0.014324f
C12910 DVDD.n2634 VSS 0.026221f
C12911 DVDD.n2635 VSS 0.017238f
C12912 DVDD.n2636 VSS 0.026221f
C12913 DVDD.n2637 VSS 0.017238f
C12914 DVDD.n2638 VSS 0.026221f
C12915 DVDD.n2639 VSS 0.026221f
C12916 DVDD.n2640 VSS 0.016752f
C12917 DVDD.n2641 VSS 0.013596f
C12918 DVDD.n2642 VSS 0.026221f
C12919 DVDD.n2643 VSS 0.017238f
C12920 DVDD.n2644 VSS 0.016509f
C12921 DVDD.n2645 VSS 0.029619f
C12922 DVDD.n2646 VSS 0.012868f
C12923 DVDD.n2647 VSS 0.031562f
C12924 DVDD.n2649 VSS 0.017238f
C12925 DVDD.n2650 VSS 0.013744f
C12926 DVDD.n2651 VSS 0.036914f
C12927 DVDD.n2652 VSS 0.018737f
C12928 DVDD.n2653 VSS 0.053101f
C12929 DVDD.n2654 VSS 0.026221f
C12930 DVDD.n2655 VSS 0.018209f
C12931 DVDD.n2656 VSS 0.014778f
C12932 DVDD.n2657 VSS 0.026221f
C12933 DVDD.n2658 VSS 0.018737f
C12934 DVDD.n2659 VSS 0.026221f
C12935 DVDD.n2660 VSS 0.018737f
C12936 DVDD.n2661 VSS 0.026221f
C12937 DVDD.n2662 VSS 0.018737f
C12938 DVDD.n2663 VSS 0.026221f
C12939 DVDD.n2664 VSS 0.026221f
C12940 DVDD.n2665 VSS 0.014514f
C12941 DVDD.n2666 VSS 0.018473f
C12942 DVDD.n2667 VSS 0.026221f
C12943 DVDD.n2668 VSS 0.026221f
C12944 DVDD.n2669 VSS 0.018737f
C12945 DVDD.n2670 VSS 0.065578f
C12946 DVDD.n2671 VSS 0.131155f
C12947 DVDD.n2672 VSS 0.131155f
C12948 DVDD.n2673 VSS 0.131155f
C12949 DVDD.n2674 VSS 0.131155f
C12950 DVDD.n2675 VSS 0.131155f
C12951 DVDD.n2676 VSS 0.131155f
C12952 DVDD.n2677 VSS 0.131155f
C12953 DVDD.n2678 VSS 0.131155f
C12954 DVDD.n2679 VSS 0.131155f
C12955 DVDD.n2680 VSS 0.131155f
C12956 DVDD.n2681 VSS 0.123305f
C12957 DVDD.n2682 VSS 0.131155f
C12958 DVDD.n2683 VSS 0.131155f
C12959 DVDD.n2684 VSS 0.131155f
C12960 DVDD.n2685 VSS 4.71774f
C12961 DVDD.n2686 VSS 0.071912f
C12962 DVDD.n2687 VSS 0.607409f
C12963 DVDD.n2688 VSS 0.090936f
C12964 DVDD.n2689 VSS 0.266203f
C12965 DVDD.n2690 VSS 0.281047f
C12966 DVDD.n2691 VSS 0.281047f
C12967 DVDD.n2692 VSS 0.214744f
C12968 DVDD.n2693 VSS 0.281047f
C12969 DVDD.n2694 VSS 0.451259f
C12970 DVDD.n2695 VSS 0.451259f
C12971 DVDD.n2696 VSS 0.140524f
C12972 DVDD.n2697 VSS 0.00712f
C12973 DVDD.n2698 VSS 0.140524f
C12974 DVDD.n2699 VSS 0.281047f
C12975 DVDD.n2700 VSS 0.281047f
C12976 DVDD.n2701 VSS 2.80563f
C12977 DVDD.n2702 VSS 1.17847f
C12978 DVDD.n2703 VSS 0.07422f
C12979 DVDD.n2704 VSS 0.140524f
C12980 DVDD.n2705 VSS 0.00712f
C12981 DVDD.n2706 VSS 0.140524f
C12982 DVDD.n2707 VSS 0.167747f
C12983 DVDD.n2708 VSS 0.34739f
C12984 DVDD.n2709 VSS 0.336402f
C12985 DVDD.n2710 VSS 0.169743f
C12986 DVDD.n2711 VSS 0.167747f
C12987 DVDD.n2712 VSS 0.169743f
C12988 DVDD.n2713 VSS 0.167747f
C12989 DVDD.n2714 VSS 0.169743f
C12990 DVDD.n2715 VSS 0.377053f
C12991 DVDD.n2716 VSS 0.295314f
C12992 DVDD.n2717 VSS 0.04049f
C12993 DVDD.n2718 VSS 0.04049f
C12994 DVDD.n2719 VSS 0.04049f
C12995 DVDD.n2720 VSS 2.56448f
C12996 DVDD.n2721 VSS 0.281047f
C12997 DVDD.n2722 VSS 0.281047f
C12998 DVDD.n2723 VSS 0.281047f
C12999 DVDD.n2724 VSS 0.140524f
C13000 DVDD.n2725 VSS 0.326766f
C13001 DVDD.n2726 VSS 0.467093f
C13002 DVDD.n2727 VSS 0.281047f
C13003 DVDD.n2728 VSS 0.281047f
C13004 DVDD.n2729 VSS 0.140524f
C13005 DVDD.n2730 VSS 0.318652f
C13006 DVDD.n2731 VSS 0.00712f
C13007 DVDD.n2732 VSS 0.140524f
C13008 DVDD.n2733 VSS 0.206827f
C13009 DVDD.n2734 VSS 0.347418f
C13010 DVDD.n2735 VSS 0.346681f
C13011 DVDD.n2736 VSS 1.15913f
C13012 DVDD.n2737 VSS 0.206827f
C13013 DVDD.n2738 VSS 0.028632f
C13014 DVDD.n2739 VSS 0.214744f
C13015 DVDD.n2740 VSS 0.169208f
C13016 DVDD.n2741 VSS 0.169748f
C13017 DVDD.n2742 VSS 0.380561f
C13018 DVDD.n2743 VSS 0.206827f
C13019 DVDD.n2744 VSS 0.214744f
C13020 DVDD.n2745 VSS 0.150773f
C13021 DVDD.n2746 VSS 0.169751f
C13022 DVDD.n2747 VSS 0.169208f
C13023 DVDD.n2748 VSS 0.214744f
C13024 DVDD.n2749 VSS 0.281047f
C13025 DVDD.n2750 VSS 1.40791f
C13026 DVDD.n2751 VSS 0.070262f
C13027 DVDD.n2752 VSS 0.277089f
C13028 DVDD.n2753 VSS 0.281047f
C13029 DVDD.n2754 VSS 0.281047f
C13030 DVDD.n2755 VSS 0.467093f
C13031 DVDD.n2756 VSS 0.281047f
C13032 DVDD.n2757 VSS 0.442353f
C13033 DVDD.n2758 VSS 0.140524f
C13034 DVDD.n2759 VSS 0.140524f
C13035 DVDD.n2760 VSS 0.281047f
C13036 DVDD.n2761 VSS 0.206827f
C13037 DVDD.n2762 VSS 0.140524f
C13038 DVDD.n2763 VSS 0.013839f
C13039 DVDD.n2764 VSS 0.01311f
C13040 DVDD.n2765 VSS 0.026221f
C13041 DVDD.n2766 VSS -0.22979f
C13042 DVDD.n2767 VSS 0.017238f
C13043 DVDD.n2768 VSS 0.07422f
C13044 DVDD.n2769 VSS 0.140524f
C13045 DVDD.n2770 VSS 0.140524f
C13046 DVDD.n2771 VSS 0.214744f
C13047 DVDD.n2772 VSS 0.281047f
C13048 DVDD.n2773 VSS 0.214744f
C13049 DVDD.n2774 VSS 0.451259f
C13050 DVDD.n2775 VSS 0.140524f
C13051 DVDD.n2776 VSS 0.316673f
C13052 DVDD.n2777 VSS 0.140524f
C13053 DVDD.n2778 VSS 0.281047f
C13054 DVDD.n2779 VSS 0.281047f
C13055 DVDD.n2780 VSS 0.140524f
C13056 DVDD.n2781 VSS 0.01311f
C13057 DVDD.n2782 VSS 0.01311f
C13058 DVDD.n2783 VSS 0.01311f
C13059 DVDD.n2784 VSS 0.01311f
C13060 DVDD.n2785 VSS 0.01311f
C13061 DVDD.n2786 VSS 0.01311f
C13062 DVDD.n2787 VSS 0.01311f
C13063 DVDD.n2788 VSS 0.021365f
C13064 DVDD.n2789 VSS 0.025393f
C13065 DVDD.n2790 VSS 0.028891f
C13066 DVDD.n2791 VSS 0.018816f
C13067 DVDD.n2792 VSS 0.01311f
C13068 DVDD.n2793 VSS 0.01311f
C13069 DVDD.n2794 VSS 0.01311f
C13070 DVDD.n2795 VSS 0.01311f
C13071 DVDD.n2796 VSS 0.01311f
C13072 DVDD.n2797 VSS 0.01311f
C13073 DVDD.n2798 VSS 0.016873f
C13074 DVDD.n2799 VSS 0.140524f
C13075 DVDD.n2800 VSS 0.026221f
C13076 DVDD.n2801 VSS 0.140524f
C13077 DVDD.n2802 VSS 0.01311f
C13078 DVDD.n2803 VSS 0.026221f
C13079 DVDD.n2804 VSS -0.22979f
C13080 DVDD.n2805 VSS 0.026221f
C13081 DVDD.n2806 VSS 0.017238f
C13082 DVDD.n2807 VSS 0.140524f
C13083 DVDD.n2808 VSS 0.140524f
C13084 DVDD.n2809 VSS 0.01311f
C13085 DVDD.n2810 VSS 0.017238f
C13086 DVDD.n2811 VSS 0.026221f
C13087 DVDD.n2812 VSS 0.026221f
C13088 DVDD.n2813 VSS 0.017966f
C13089 DVDD.n2814 VSS 0.026221f
C13090 DVDD.n2815 VSS 0.015781f
C13091 DVDD.n2816 VSS 0.015781f
C13092 DVDD.n2817 VSS 0.006715f
C13093 DVDD.n2818 VSS 0.059907f
C13094 DVDD.n2819 VSS 0.017238f
C13095 DVDD.n2820 VSS 0.036053f
C13096 DVDD.n2821 VSS 0.036053f
C13097 DVDD.n2822 VSS 0.014688f
C13098 DVDD.n2823 VSS 0.015659f
C13099 DVDD.n2824 VSS 0.026221f
C13100 DVDD.n2825 VSS 0.017238f
C13101 DVDD.n2826 VSS 0.026221f
C13102 DVDD.n2827 VSS 0.017238f
C13103 DVDD.n2828 VSS 0.026221f
C13104 DVDD.n2829 VSS 0.026221f
C13105 DVDD.n2830 VSS 0.015417f
C13106 DVDD.n2831 VSS 0.014931f
C13107 DVDD.n2832 VSS 0.026221f
C13108 DVDD.n2833 VSS 0.017238f
C13109 DVDD.n2834 VSS 0.026221f
C13110 DVDD.n2835 VSS 0.017238f
C13111 DVDD.n2836 VSS 0.026221f
C13112 DVDD.n2837 VSS 0.026221f
C13113 DVDD.n2838 VSS 0.016145f
C13114 DVDD.n2839 VSS 0.014203f
C13115 DVDD.n2840 VSS 0.026221f
C13116 DVDD.n2841 VSS 0.017238f
C13117 DVDD.n2842 VSS 0.026221f
C13118 DVDD.n2843 VSS 0.017238f
C13119 DVDD.n2844 VSS 0.026221f
C13120 DVDD.n2845 VSS 0.026221f
C13121 DVDD.n2846 VSS 0.016873f
C13122 DVDD.n2847 VSS 0.013474f
C13123 DVDD.n2848 VSS 0.026221f
C13124 DVDD.n2849 VSS 0.017238f
C13125 DVDD.n2850 VSS 0.026221f
C13126 DVDD.n2851 VSS 0.017238f
C13127 DVDD.n2852 VSS 0.026221f
C13128 DVDD.n2853 VSS 0.017238f
C13129 DVDD.n2854 VSS 0.026221f
C13130 DVDD.n2855 VSS 0.013474f
C13131 DVDD.n2856 VSS 0.026221f
C13132 DVDD.n2857 VSS 0.026221f
C13133 DVDD.n2858 VSS 0.026221f
C13134 DVDD.n2859 VSS 0.140524f
C13135 DVDD.n2860 VSS 0.016873f
C13136 DVDD.n2861 VSS 0.310735f
C13137 DVDD.n2862 VSS 0.140524f
C13138 DVDD.n2863 VSS 0.01311f
C13139 DVDD.n2864 VSS 0.01311f
C13140 DVDD.n2865 VSS 0.01311f
C13141 DVDD.n2866 VSS 0.01311f
C13142 DVDD.n2867 VSS 0.01311f
C13143 DVDD.n2868 VSS 0.01311f
C13144 DVDD.n2869 VSS 0.01311f
C13145 DVDD.n2870 VSS 0.025393f
C13146 DVDD.n2871 VSS 0.021365f
C13147 DVDD.n2872 VSS 0.140524f
C13148 DVDD.n2873 VSS 0.028891f
C13149 DVDD.n2874 VSS 0.01311f
C13150 DVDD.n2875 VSS 0.01311f
C13151 DVDD.n2876 VSS 0.01311f
C13152 DVDD.n2877 VSS 0.01311f
C13153 DVDD.n2878 VSS 0.01311f
C13154 DVDD.n2879 VSS 0.01311f
C13155 DVDD.n2880 VSS 0.015659f
C13156 DVDD.n2881 VSS 0.013474f
C13157 DVDD.n2882 VSS 0.026221f
C13158 DVDD.n2883 VSS 0.017238f
C13159 DVDD.n2884 VSS 0.026221f
C13160 DVDD.n2885 VSS 0.017238f
C13161 DVDD.n2886 VSS 0.026221f
C13162 DVDD.n2887 VSS 0.017238f
C13163 DVDD.n2888 VSS 0.026221f
C13164 DVDD.n2889 VSS 0.026221f
C13165 DVDD.n2890 VSS 0.013474f
C13166 DVDD.n2891 VSS 0.016873f
C13167 DVDD.n2892 VSS 0.026221f
C13168 DVDD.n2893 VSS 0.017238f
C13169 DVDD.n2894 VSS 0.026221f
C13170 DVDD.n2895 VSS 0.017238f
C13171 DVDD.n2896 VSS 0.026221f
C13172 DVDD.n2897 VSS 0.026221f
C13173 DVDD.n2898 VSS 0.014203f
C13174 DVDD.n2899 VSS 0.016145f
C13175 DVDD.n2900 VSS 0.026221f
C13176 DVDD.n2901 VSS 0.017238f
C13177 DVDD.n2902 VSS 0.026221f
C13178 DVDD.n2903 VSS 0.017238f
C13179 DVDD.n2904 VSS 0.026221f
C13180 DVDD.n2905 VSS 0.026221f
C13181 DVDD.n2906 VSS 0.014931f
C13182 DVDD.n2907 VSS 0.015417f
C13183 DVDD.n2908 VSS 0.026221f
C13184 DVDD.n2909 VSS 0.017238f
C13185 DVDD.n2910 VSS 0.026221f
C13186 DVDD.n2911 VSS 0.017238f
C13187 DVDD.n2912 VSS 0.026221f
C13188 DVDD.n2913 VSS 0.025978f
C13189 DVDD.n2914 VSS 0.026221f
C13190 DVDD.n2915 VSS 0.01311f
C13191 DVDD.n2916 VSS 0.026221f
C13192 DVDD.n2917 VSS 0.017238f
C13193 DVDD.n2918 VSS 0.140524f
C13194 DVDD.n2919 VSS 0.140524f
C13195 DVDD.n2920 VSS 0.281047f
C13196 DVDD.n2921 VSS 0.214744f
C13197 DVDD.n2922 VSS 0.214744f
C13198 DVDD.n2923 VSS 0.140524f
C13199 DVDD.n2924 VSS 0.017238f
C13200 DVDD.n2925 VSS 0.026221f
C13201 DVDD.n2926 VSS 0.013839f
C13202 DVDD.n2927 VSS 0.140524f
C13203 DVDD.n2928 VSS 0.281047f
C13204 DVDD.n2929 VSS 0.281047f
C13205 DVDD.n2930 VSS 0.281047f
C13206 DVDD.n2931 VSS 0.140524f
C13207 DVDD.n2932 VSS 0.017238f
C13208 DVDD.n2934 VSS 0.014567f
C13209 DVDD.n2935 VSS 0.326617f
C13210 DVDD.n2937 VSS 0.028891f
C13211 DVDD.n2938 VSS 0.140524f
C13212 DVDD.n2939 VSS 0.01311f
C13213 DVDD.n2940 VSS 0.017238f
C13214 DVDD.n2941 VSS 0.015781f
C13215 DVDD.n2942 VSS 0.026221f
C13216 DVDD.n2943 VSS 0.016509f
C13217 DVDD.n2944 VSS 0.01311f
C13218 DVDD.n2945 VSS 0.140524f
C13219 DVDD.n2946 VSS 0.140524f
C13220 DVDD.n2947 VSS 0.140524f
C13221 DVDD.n2948 VSS 0.01311f
C13222 DVDD.n2949 VSS 0.017238f
C13223 DVDD.n2950 VSS 0.031562f
C13224 DVDD.n2951 VSS 0.029086f
C13225 DVDD.n2952 VSS 0.013558f
C13226 DVDD.n2953 VSS 0.013558f
C13227 DVDD.n2955 VSS 0.031562f
C13228 DVDD.n2956 VSS 0.014567f
C13229 DVDD.n2957 VSS 0.029086f
C13230 DVDD.n2958 VSS 0.326617f
C13231 DVDD.n2959 VSS 0.467093f
C13232 DVDD.n2960 VSS 0.281047f
C13233 DVDD.n2961 VSS 0.281047f
C13234 DVDD.n2962 VSS 0.140607f
C13235 DVDD.n2963 VSS 0.352374f
C13236 DVDD.n2964 VSS 0.093023f
C13237 DVDD.n2965 VSS 0.140524f
C13238 DVDD.n2966 VSS 0.00712f
C13239 DVDD.n2967 VSS 0.140524f
C13240 DVDD.n2968 VSS 0.281047f
C13241 DVDD.n2969 VSS 0.214744f
C13242 DVDD.n2970 VSS 0.263903f
C13243 DVDD.n2971 VSS 0.140524f
C13244 DVDD.n2972 VSS 0.018672f
C13245 DVDD.n2973 VSS 0.140524f
C13246 DVDD.n2974 VSS 0.253238f
C13247 DVDD.n2975 VSS 0.281047f
C13248 DVDD.n2976 VSS 0.269822f
C13249 DVDD.n2977 VSS 0.798425f
C13250 DVDD.n2978 VSS 0.281047f
C13251 DVDD.n2979 VSS 0.281047f
C13252 DVDD.n2980 VSS 0.140524f
C13253 DVDD.n2981 VSS 0.140524f
C13254 DVDD.n2982 VSS 0.00534f
C13255 DVDD.n2983 VSS 0.00356f
C13256 DVDD.n2984 VSS 0.00534f
C13257 DVDD.n2985 VSS 0.066303f
C13258 DVDD.n2986 VSS 0.009896f
C13259 DVDD.n2987 VSS 0.281047f
C13260 DVDD.n2988 VSS 0.281047f
C13261 DVDD.n2989 VSS 0.281047f
C13262 DVDD.n2990 VSS 0.281047f
C13263 DVDD.n2991 VSS 0.327059f
C13264 DVDD.n2992 VSS 0.281047f
C13265 DVDD.n2993 VSS 0.467093f
C13266 DVDD.n2994 VSS 0.467093f
C13267 DVDD.n2995 VSS 0.281047f
C13268 DVDD.n2996 VSS 0.110836f
C13269 DVDD.n2997 VSS 0.00906f
C13270 DVDD.n2998 VSS 0.070192f
C13271 DVDD.t216 VSS 0.156498f
C13272 DVDD.n2999 VSS 0.121191f
C13273 DVDD.n3000 VSS 0.037832f
C13274 DVDD.n3001 VSS 0.127659f
C13275 DVDD.n3002 VSS 0.281047f
C13276 DVDD.n3003 VSS 0.281047f
C13277 DVDD.n3004 VSS 0.281047f
C13278 DVDD.n3005 VSS 0.206827f
C13279 DVDD.n3006 VSS 0.206827f
C13280 DVDD.n3007 VSS 0.1237f
C13281 DVDD.n3008 VSS 0.108856f
C13282 DVDD.n3009 VSS 0.037832f
C13283 DVDD.n3010 VSS 0.037832f
C13284 DVDD.n3011 VSS 0.140524f
C13285 DVDD.n3012 VSS 0.214744f
C13286 DVDD.n3013 VSS 0.281047f
C13287 DVDD.n3014 VSS 0.281047f
C13288 DVDD.n3015 VSS 0.131617f
C13289 DVDD.n3016 VSS 0.00906f
C13290 DVDD.n3017 VSS 0.070192f
C13291 DVDD.t214 VSS 0.156498f
C13292 DVDD.n3018 VSS 0.121191f
C13293 DVDD.n3019 VSS 0.110836f
C13294 DVDD.n3020 VSS 0.451259f
C13295 DVDD.n3021 VSS 0.281047f
C13296 DVDD.n3022 VSS 0.281047f
C13297 DVDD.n3023 VSS 0.451259f
C13298 DVDD.n3024 VSS 0.451259f
C13299 DVDD.n3025 VSS 0.281047f
C13300 DVDD.n3026 VSS 0.281047f
C13301 DVDD.n3027 VSS 0.281047f
C13302 DVDD.n3028 VSS 0.281047f
C13303 DVDD.n3029 VSS 0.281047f
C13304 DVDD.n3030 VSS 0.214744f
C13305 DVDD.n3031 VSS 0.281047f
C13306 DVDD.n3032 VSS 0.281047f
C13307 DVDD.n3033 VSS 0.281047f
C13308 DVDD.n3034 VSS 0.281047f
C13309 DVDD.n3035 VSS 0.451259f
C13310 DVDD.n3036 VSS 0.451259f
C13311 DVDD.n3037 VSS 0.451259f
C13312 DVDD.n3038 VSS 0.281047f
C13313 DVDD.n3039 VSS 0.190993f
C13314 DVDD.n3040 VSS 0.14064f
C13315 DVDD.n3041 VSS 0.00906f
C13316 DVDD.n3042 VSS 0.070192f
C13317 DVDD.t215 VSS 0.156498f
C13318 DVDD.n3043 VSS 0.121191f
C13319 DVDD.n3044 VSS 0.041938f
C13320 DVDD.n3045 VSS 0.030569f
C13321 DVDD.n3046 VSS 0.037832f
C13322 DVDD.n3047 VSS 0.119742f
C13323 DVDD.n3048 VSS 0.110836f
C13324 DVDD.n3049 VSS 0.281047f
C13325 DVDD.n3050 VSS 0.214744f
C13326 DVDD.n3051 VSS 0.110836f
C13327 DVDD.n3052 VSS 0.07422f
C13328 DVDD.n3053 VSS 0.037832f
C13329 DVDD.n3054 VSS 0.037832f
C13330 DVDD.n3055 VSS 0.140524f
C13331 DVDD.n3056 VSS 0.110836f
C13332 DVDD.n3057 VSS 0.281047f
C13333 DVDD.n3058 VSS 0.281047f
C13334 DVDD.n3059 VSS 0.110836f
C13335 DVDD.n3060 VSS 0.140524f
C13336 DVDD.n3061 VSS 0.031414f
C13337 DVDD.n3062 VSS 0.00906f
C13338 DVDD.n3063 VSS 0.070192f
C13339 DVDD.t220 VSS 0.156498f
C13340 DVDD.n3064 VSS 0.121191f
C13341 DVDD.n3065 VSS 0.018916f
C13342 DVDD.n3066 VSS 0.062676f
C13343 DVDD.n3067 VSS 0.140524f
C13344 DVDD.n3068 VSS 0.110836f
C13345 DVDD.n3069 VSS 0.467093f
C13346 DVDD.n3070 VSS 0.467093f
C13347 DVDD.n3071 VSS 0.432457f
C13348 DVDD.n3072 VSS 0.281047f
C13349 DVDD.n3073 VSS 0.281047f
C13350 DVDD.n3074 VSS 0.281047f
C13351 DVDD.n3075 VSS 0.281047f
C13352 DVDD.n3076 VSS 0.206827f
C13353 DVDD.n3077 VSS 0.206827f
C13354 DVDD.n3078 VSS 0.07422f
C13355 DVDD.n3079 VSS 0.051795f
C13356 DVDD.n3080 VSS 0.009368f
C13357 DVDD.n3081 VSS 0.140524f
C13358 DVDD.n3082 VSS 0.038693f
C13359 DVDD.n3083 VSS 0.038693f
C13360 DVDD.n3084 VSS 0.010399f
C13361 DVDD.n3085 VSS 0.074622f
C13362 DVDD.n3086 VSS 0.007909f
C13363 DVDD.n3087 VSS 0.007909f
C13364 DVDD.n3088 VSS 0.009081f
C13365 DVDD.n3089 VSS 0.140524f
C13366 DVDD.n3090 VSS 0.041782f
C13367 DVDD.n3091 VSS 0.041782f
C13368 DVDD.n3092 VSS 0.140524f
C13369 DVDD.n3093 VSS 0.041782f
C13370 DVDD.n3094 VSS 0.007909f
C13371 DVDD.n3095 VSS 0.038294f
C13372 DVDD.n3096 VSS 0.01157f
C13373 DVDD.n3097 VSS 0.267309f
C13374 DVDD.n3098 VSS 0.045607f
C13375 DVDD.n3099 VSS 0.798425f
C13376 DVDD.n3100 VSS 0.281047f
C13377 DVDD.n3101 VSS 0.214744f
C13378 DVDD.n3102 VSS 0.281047f
C13379 DVDD.n3103 VSS 0.281047f
C13380 DVDD.n3104 VSS 0.281047f
C13381 DVDD.n3105 VSS 0.140524f
C13382 DVDD.n3106 VSS 0.210235f
C13383 DVDD.n3107 VSS 0.064248f
C13384 DVDD.n3108 VSS 0.130405f
C13385 DVDD.n3109 VSS 0.250777f
C13386 DVDD.n3110 VSS 0.022624f
C13387 DVDD.n3111 VSS 0.110619f
C13388 DVDD.n3112 VSS 0.083329f
C13389 DVDD.n3113 VSS 0.005003f
C13390 DVDD.n3114 VSS 0.020672f
C13391 DVDD.n3115 VSS 0.037528f
C13392 DVDD.n3116 VSS 0.249487f
C13393 DVDD.n3117 VSS 0.093076f
C13394 DVDD.n3118 VSS 0.050379f
C13395 DVDD.n3119 VSS 0.144777f
C13396 DVDD.n3120 VSS 0.020891f
C13397 DVDD.n3121 VSS 0.050379f
C13398 DVDD.n3122 VSS 0.010399f
C13399 DVDD.n3123 VSS 0.012303f
C13400 DVDD.n3124 VSS 0.015671f
C13401 DVDD.n3125 VSS 0.009227f
C13402 DVDD.n3126 VSS 0.140524f
C13403 DVDD.n3127 VSS 0.140524f
C13404 DVDD.n3128 VSS 0.038693f
C13405 DVDD.n3129 VSS 0.041782f
C13406 DVDD.n3130 VSS 0.041782f
C13407 DVDD.n3131 VSS 0.038693f
C13408 DVDD.n3132 VSS 0.018737f
C13409 DVDD.n3133 VSS 0.037473f
C13410 DVDD.n3134 VSS 0.034668f
C13411 DVDD.n3135 VSS 0.045607f
C13412 DVDD.n3136 VSS 0.140524f
C13413 DVDD.n3137 VSS 0.140524f
C13414 DVDD.n3138 VSS 0.041782f
C13415 DVDD.n3139 VSS 0.010399f
C13416 DVDD.n3140 VSS 0.041782f
C13417 DVDD.n3141 VSS 0.140524f
C13418 DVDD.n3142 VSS 0.007909f
C13419 DVDD.n3143 VSS 0.022624f
C13420 DVDD.n3144 VSS 0.071492f
C13421 DVDD.n3145 VSS 0.004906f
C13422 DVDD.n3146 VSS 0.040299f
C13423 DVDD.n3147 VSS 0.080571f
C13424 DVDD.n3148 VSS 0.564594f
C13425 DVDD.n3149 VSS 0.110619f
C13426 DVDD.n3150 VSS 0.010225f
C13427 DVDD.n3151 VSS 0.005036f
C13428 DVDD.n3152 VSS 0.023207f
C13429 DVDD.n3153 VSS 0.013485f
C13430 DVDD.n3154 VSS 0.020672f
C13431 DVDD.n3155 VSS 0.126387f
C13432 DVDD.n3156 VSS 0.281047f
C13433 DVDD.n3157 VSS 0.281047f
C13434 DVDD.n3158 VSS 0.214744f
C13435 DVDD.n3159 VSS 0.281047f
C13436 DVDD.n3160 VSS 0.281047f
C13437 DVDD.n3161 VSS 0.798425f
C13438 DVDD.n3162 VSS 0.267309f
C13439 DVDD.n3163 VSS 0.01157f
C13440 DVDD.n3164 VSS 0.007909f
C13441 DVDD.n3165 VSS 0.260334f
C13442 DVDD.n3166 VSS 0.045607f
C13443 DVDD.n3167 VSS 0.272214f
C13444 DVDD.n3168 VSS 0.157642f
C13445 DVDD.n3169 VSS 0.245208f
C13446 DVDD.n3170 VSS 0.272214f
C13447 DVDD.n3171 VSS 0.210235f
C13448 DVDD.n3172 VSS 0.128218f
C13449 DVDD.n3173 VSS 0.038294f
C13450 DVDD.n3174 VSS 0.012596f
C13451 DVDD.n3175 VSS 0.007909f
C13452 DVDD.n3176 VSS 0.009081f
C13453 DVDD.n3177 VSS 0.008055f
C13454 DVDD.n3178 VSS 0.015818f
C13455 DVDD.n3179 VSS 0.010399f
C13456 DVDD.n3180 VSS 0.007909f
C13457 DVDD.n3181 VSS 0.140524f
C13458 DVDD.n3182 VSS 0.041782f
C13459 DVDD.n3183 VSS 0.018737f
C13460 DVDD.n3184 VSS 0.018737f
C13461 DVDD.n3185 VSS 0.140524f
C13462 DVDD.n3186 VSS 0.041782f
C13463 DVDD.n3187 VSS 0.018737f
C13464 DVDD.n3188 VSS 0.018737f
C13465 DVDD.n3189 VSS 0.037473f
C13466 DVDD.n3190 VSS 0.03585f
C13467 DVDD.n3191 VSS 0.106291f
C13468 DVDD.n3192 VSS 0.037473f
C13469 DVDD.n3193 VSS 0.037473f
C13470 DVDD.n3194 VSS 0.028632f
C13471 DVDD.n3195 VSS 0.018737f
C13472 DVDD.n3196 VSS 0.018737f
C13473 DVDD.n3197 VSS 0.041782f
C13474 DVDD.n3198 VSS 0.140524f
C13475 DVDD.n3199 VSS 0.007909f
C13476 DVDD.n3200 VSS 0.007909f
C13477 DVDD.n3201 VSS 0.010399f
C13478 DVDD.n3202 VSS 0.012449f
C13479 DVDD.n3203 VSS 0.012449f
C13480 DVDD.n3204 VSS 0.144777f
C13481 DVDD.n3205 VSS 0.074622f
C13482 DVDD.n3206 VSS 0.01157f
C13483 DVDD.n3207 VSS 0.007909f
C13484 DVDD.n3208 VSS 0.140607f
C13485 DVDD.n3209 VSS 0.029571f
C13486 DVDD.n3210 VSS 0.154817f
C13487 DVDD.n3211 VSS 0.029571f
C13488 DVDD.n3212 VSS 0.020891f
C13489 DVDD.n3213 VSS 0.093076f
C13490 DVDD.n3214 VSS 0.037933f
C13491 DVDD.n3215 VSS 0.41812f
C13492 DVDD.n3216 VSS 0.249497f
C13493 DVDD.n3217 VSS 0.023207f
C13494 DVDD.n3218 VSS 0.013455f
C13495 DVDD.n3219 VSS 0.07143f
C13496 DVDD.n3220 VSS 0.004876f
C13497 DVDD.n3221 VSS 0.01026f
C13498 DVDD.n3222 VSS 0.128218f
C13499 DVDD.n3223 VSS 0.250785f
C13500 DVDD.n3224 VSS 0.417154f
C13501 DVDD.n3225 VSS 0.037933f
C13502 DVDD.n3226 VSS 0.130405f
C13503 DVDD.n3227 VSS 0.272214f
C13504 DVDD.n3228 VSS 0.157642f
C13505 DVDD.n3229 VSS 0.126387f
C13506 DVDD.n3230 VSS 0.245208f
C13507 DVDD.n3231 VSS 0.272214f
C13508 DVDD.n3232 VSS 0.045607f
C13509 DVDD.n3233 VSS 0.260334f
C13510 DVDD.n3234 VSS 0.007909f
C13511 DVDD.n3235 VSS 0.010399f
C13512 DVDD.n3236 VSS 0.012596f
C13513 DVDD.n3237 VSS 0.008055f
C13514 DVDD.n3238 VSS 0.015818f
C13515 DVDD.n3239 VSS 0.010399f
C13516 DVDD.n3240 VSS 0.007909f
C13517 DVDD.n3241 VSS 0.140524f
C13518 DVDD.n3242 VSS 0.041782f
C13519 DVDD.n3243 VSS 0.041782f
C13520 DVDD.n3244 VSS 0.140524f
C13521 DVDD.n3245 VSS 0.007909f
C13522 DVDD.n3246 VSS 0.009227f
C13523 DVDD.n3247 VSS 0.015671f
C13524 DVDD.n3248 VSS 0.012449f
C13525 DVDD.n3249 VSS 0.012449f
C13526 DVDD.n3250 VSS 0.01157f
C13527 DVDD.n3251 VSS 0.012303f
C13528 DVDD.n3252 VSS 0.010399f
C13529 DVDD.n3253 VSS 0.007909f
C13530 DVDD.n3254 VSS 0.07422f
C13531 DVDD.n3255 VSS 3.54248f
C13532 DVDD.n3256 VSS 0.070262f
C13533 DVDD.n3257 VSS 0.206827f
C13534 DVDD.n3258 VSS 0.281047f
C13535 DVDD.n3259 VSS 0.281047f
C13536 DVDD.n3260 VSS 0.277089f
C13537 DVDD.n3261 VSS 0.281047f
C13538 DVDD.n3262 VSS 0.442353f
C13539 DVDD.n3263 VSS 0.281047f
C13540 DVDD.n3264 VSS 0.281047f
C13541 DVDD.n3265 VSS 0.281047f
C13542 DVDD.n3266 VSS 0.467093f
C13543 DVDD.n3267 VSS 0.467093f
C13544 DVDD.n3268 VSS 0.467093f
C13545 DVDD.n3269 VSS 0.140524f
C13546 DVDD.n3270 VSS 0.140524f
C13547 DVDD.n3271 VSS 0.140524f
C13548 DVDD.n3272 VSS 0.01311f
C13549 DVDD.n3273 VSS 0.01311f
C13550 DVDD.n3274 VSS 0.017238f
C13551 DVDD.n3276 VSS 0.028891f
C13552 DVDD.n3277 VSS 0.015781f
C13553 DVDD.n3278 VSS 0.026221f
C13554 DVDD.n3279 VSS 0.026221f
C13555 DVDD.n3280 VSS 0.016509f
C13556 DVDD.n3281 VSS 0.01311f
C13557 DVDD.n3282 VSS 0.140524f
C13558 DVDD.n3283 VSS 0.140524f
C13559 DVDD.n3284 VSS 0.281047f
C13560 DVDD.n3285 VSS 0.281047f
C13561 DVDD.n3286 VSS 0.281047f
C13562 DVDD.n3287 VSS 0.206827f
C13563 DVDD.n3288 VSS 0.206827f
C13564 DVDD.n3289 VSS 0.091044f
C13565 DVDD.n3290 VSS 0.140524f
C13566 DVDD.n3291 VSS 0.01311f
C13567 DVDD.n3292 VSS 0.017238f
C13568 DVDD.n3293 VSS 0.140524f
C13569 DVDD.n3294 VSS 0.07422f
C13570 DVDD.n3295 VSS 0.01311f
C13571 DVDD.n3296 VSS 0.01311f
C13572 DVDD.n3297 VSS 0.017238f
C13573 DVDD.n3298 VSS 0.026221f
C13574 DVDD.n3299 VSS -0.22979f
C13575 DVDD.n3300 VSS -0.22979f
C13576 DVDD.n3301 VSS 0.026221f
C13577 DVDD.n3302 VSS 0.140524f
C13578 DVDD.n3303 VSS 0.140524f
C13579 DVDD.n3304 VSS 0.281047f
C13580 DVDD.n3305 VSS 0.281047f
C13581 DVDD.n3306 VSS 0.281047f
C13582 DVDD.n3307 VSS 0.281047f
C13583 DVDD.n3308 VSS 0.451259f
C13584 DVDD.n3309 VSS 0.451259f
C13585 DVDD.n3310 VSS 0.281047f
C13586 DVDD.n3311 VSS 0.281047f
C13587 DVDD.n3312 VSS 0.281047f
C13588 DVDD.n3313 VSS 0.214744f
C13589 DVDD.n3314 VSS 0.281047f
C13590 DVDD.n3315 VSS 0.281047f
C13591 DVDD.n3316 VSS 0.159326f
C13592 DVDD.n3317 VSS 0.281047f
C13593 DVDD.n3318 VSS 0.281047f
C13594 DVDD.n3319 VSS 0.451259f
C13595 DVDD.n3320 VSS 0.316673f
C13596 DVDD.n3321 VSS 0.451259f
C13597 DVDD.n3322 VSS 0.281047f
C13598 DVDD.n3323 VSS 0.140524f
C13599 DVDD.n3324 VSS 0.140524f
C13600 DVDD.n3325 VSS 0.01311f
C13601 DVDD.n3326 VSS 0.017238f
C13602 DVDD.n3327 VSS 0.026221f
C13603 DVDD.n3328 VSS 0.026221f
C13604 DVDD.n3329 VSS 0.017966f
C13605 DVDD.n3330 VSS 0.026221f
C13606 DVDD.n3331 VSS 0.015781f
C13607 DVDD.n3332 VSS 0.015781f
C13608 DVDD.n3333 VSS 0.006715f
C13609 DVDD.n3334 VSS 0.059907f
C13610 DVDD.n3335 VSS 0.017238f
C13611 DVDD.n3336 VSS 0.036053f
C13612 DVDD.n3337 VSS 0.023186f
C13613 DVDD.n3338 VSS 0.014688f
C13614 DVDD.n3340 VSS 0.018816f
C13615 DVDD.n3341 VSS 0.140524f
C13616 DVDD.n3342 VSS 0.031453f
C13617 DVDD.n3343 VSS -0.530288f
C13618 DVDD.n3344 VSS -0.530288f
C13619 DVDD.n3346 VSS 0.310735f
C13620 DVDD.n3347 VSS 0.031453f
C13621 DVDD.n3348 VSS 0.140524f
C13622 DVDD.n3349 VSS 0.159326f
C13623 DVDD.n3350 VSS 0.281047f
C13624 DVDD.n3351 VSS 0.214744f
C13625 DVDD.n3352 VSS 0.281047f
C13626 DVDD.n3353 VSS 0.281047f
C13627 DVDD.n3354 VSS 0.281047f
C13628 DVDD.n3355 VSS 0.281047f
C13629 DVDD.n3356 VSS 0.451259f
C13630 DVDD.n3357 VSS 0.451259f
C13631 DVDD.n3358 VSS 0.451259f
C13632 DVDD.n3359 VSS 0.281047f
C13633 DVDD.n3360 VSS 0.281047f
C13634 DVDD.n3361 VSS 0.281047f
C13635 DVDD.n3362 VSS 0.281047f
C13636 DVDD.n3363 VSS 0.281047f
C13637 DVDD.n3364 VSS 0.140524f
C13638 DVDD.n3365 VSS 0.140524f
C13639 DVDD.n3366 VSS 0.01311f
C13640 DVDD.n3367 VSS 0.017238f
C13641 DVDD.n3368 VSS 0.026221f
C13642 DVDD.n3369 VSS 0.026221f
C13643 DVDD.n3370 VSS 0.017238f
C13644 DVDD.n3371 VSS 0.01311f
C13645 DVDD.n3372 VSS 0.140524f
C13646 DVDD.n3373 VSS 0.091044f
C13647 DVDD.n3374 VSS 0.206827f
C13648 DVDD.n3375 VSS 0.281047f
C13649 DVDD.n3376 VSS 0.281047f
C13650 DVDD.n3377 VSS 0.281047f
C13651 DVDD.n3378 VSS 0.281047f
C13652 DVDD.n3379 VSS 0.281047f
C13653 DVDD.n3380 VSS 0.467093f
C13654 DVDD.n3381 VSS 0.467093f
C13655 DVDD.n3382 VSS 0.467093f
C13656 DVDD.n3383 VSS 0.281047f
C13657 DVDD.n3384 VSS 0.281047f
C13658 DVDD.n3385 VSS 0.281047f
C13659 DVDD.n3386 VSS 0.281047f
C13660 DVDD.n3387 VSS 0.206827f
C13661 DVDD.n3388 VSS 0.206827f
C13662 DVDD.n3389 VSS 3.8854f
C13663 DVDD.n3390 VSS 0.206827f
C13664 DVDD.n3391 VSS 0.281047f
C13665 DVDD.n3392 VSS 0.281047f
C13666 DVDD.n3393 VSS 0.140524f
C13667 DVDD.n3394 VSS 0.140524f
C13668 DVDD.n3395 VSS 0.140524f
C13669 DVDD.n3396 VSS 0.00712f
C13670 DVDD.n3397 VSS 0.012388f
C13671 DVDD.n3398 VSS 0.140721f
C13672 DVDD.n3399 VSS 0.140524f
C13673 DVDD.n3400 VSS 0.281047f
C13674 DVDD.n3401 VSS 0.281047f
C13675 DVDD.n3402 VSS 0.467093f
C13676 DVDD.n3403 VSS 0.467093f
C13677 DVDD.n3404 VSS 0.467093f
C13678 DVDD.n3405 VSS 0.140524f
C13679 DVDD.n3406 VSS 0.140524f
C13680 DVDD.n3407 VSS 0.012388f
C13681 DVDD.n3408 VSS 0.00712f
C13682 DVDD.n3409 VSS 0.140524f
C13683 DVDD.n3410 VSS 0.140524f
C13684 DVDD.n3411 VSS 0.140524f
C13685 DVDD.n3412 VSS 0.281047f
C13686 DVDD.n3413 VSS 0.281047f
C13687 DVDD.n3414 VSS 0.281047f
C13688 DVDD.n3415 VSS 0.206827f
C13689 DVDD.n3416 VSS 0.206827f
C13690 DVDD.n3417 VSS 0.093023f
C13691 DVDD.n3418 VSS 0.140524f
C13692 DVDD.n3419 VSS 0.00534f
C13693 DVDD.n3420 VSS 0.00356f
C13694 DVDD.n3421 VSS 0.00534f
C13695 DVDD.n3422 VSS 0.00712f
C13696 DVDD.n3423 VSS 0.140524f
C13697 DVDD.n3424 VSS 0.140524f
C13698 DVDD.n3425 VSS 0.214744f
C13699 DVDD.n3426 VSS 0.214744f
C13700 DVDD.n3427 VSS 0.281047f
C13701 DVDD.n3428 VSS 0.281047f
C13702 DVDD.n3429 VSS 0.281047f
C13703 DVDD.n3430 VSS 0.281047f
C13704 DVDD.n3431 VSS 0.140524f
C13705 DVDD.n3432 VSS 0.140524f
C13706 DVDD.n3433 VSS 0.012388f
C13707 DVDD.n3434 VSS 0.140721f
C13708 DVDD.n3435 VSS 0.337455f
C13709 DVDD.n3436 VSS 0.451259f
C13710 DVDD.n3437 VSS 0.451259f
C13711 DVDD.n3438 VSS 0.451259f
C13712 DVDD.n3439 VSS 0.281047f
C13713 DVDD.n3440 VSS 0.281047f
C13714 DVDD.n3441 VSS 0.281047f
C13715 DVDD.n3442 VSS 0.281047f
C13716 DVDD.n3443 VSS 0.155368f
C13717 DVDD.n3444 VSS 0.194943f
C13718 DVDD.n3445 VSS 0.106356f
C13719 DVDD.n3446 VSS 2.93858f
C13720 DVDD.t61 VSS 3.96646f
C13721 DVDD.t26 VSS 1.36533f
C13722 DVDD.n3447 VSS 4.37787f
C13723 DVDD.n3448 VSS 0.392955f
C13724 DVDD.n3449 VSS 0.074538f
C13725 DVDD.n3450 VSS 0.160292f
C13726 DVDD.n3451 VSS 0.09228f
C13727 DVDD.n3452 VSS 0.131155f
C13728 DVDD.n3453 VSS 0.131155f
C13729 DVDD.n3454 VSS 0.131155f
C13730 DVDD.n3455 VSS 0.131155f
C13731 DVDD.n3456 VSS 0.131155f
C13732 DVDD.n3457 VSS 0.131155f
C13733 DVDD.n3458 VSS 0.131155f
C13734 DVDD.n3459 VSS 0.131155f
C13735 DVDD.n3460 VSS 0.131155f
C13736 DVDD.n3461 VSS 0.131155f
C13737 DVDD.n3462 VSS 0.131155f
C13738 DVDD.n3463 VSS 0.131155f
C13739 DVDD.n3464 VSS 0.131155f
C13740 DVDD.n3465 VSS 0.131155f
C13741 DVDD.n3466 VSS 0.131155f
C13742 DVDD.n3467 VSS 0.131155f
C13743 DVDD.n3468 VSS 0.118225f
C13744 DVDD.n3469 VSS 0.118225f
C13745 DVDD.n3470 VSS 0.63196f
C13746 DVDD.n3471 VSS 0.172652f
C13747 DVDD.n3472 VSS 0.067425f
C13748 DVDD.n3473 VSS 0.131155f
C13749 DVDD.n3474 VSS 0.131155f
C13750 DVDD.n3475 VSS 0.131155f
C13751 DVDD.n3476 VSS 0.131155f
C13752 DVDD.n3477 VSS 0.131155f
C13753 DVDD.n3478 VSS 0.131155f
C13754 DVDD.n3479 VSS 0.131155f
C13755 DVDD.n3480 VSS 0.131155f
C13756 DVDD.n3481 VSS 0.131155f
C13757 DVDD.n3482 VSS 0.131155f
C13758 DVDD.n3483 VSS 0.131155f
C13759 DVDD.n3484 VSS 0.131155f
C13760 DVDD.n3485 VSS 0.131155f
C13761 DVDD.n3486 VSS 0.131155f
C13762 DVDD.n3487 VSS 0.131155f
C13763 DVDD.n3488 VSS 0.131155f
C13764 DVDD.n3489 VSS 0.131155f
C13765 DVDD.n3490 VSS 0.131155f
C13766 DVDD.n3491 VSS 0.131155f
C13767 DVDD.n3492 VSS 0.131155f
C13768 DVDD.n3493 VSS 0.131155f
C13769 DVDD.n3494 VSS 0.131155f
C13770 DVDD.n3495 VSS 0.131155f
C13771 DVDD.n3496 VSS 0.131155f
C13772 DVDD.n3497 VSS 0.131155f
C13773 DVDD.n3498 VSS 0.131155f
C13774 DVDD.n3499 VSS 0.131155f
C13775 DVDD.n3500 VSS 0.131155f
C13776 DVDD.n3501 VSS 0.131155f
C13777 DVDD.n3502 VSS 0.131155f
C13778 DVDD.n3503 VSS 0.131155f
C13779 DVDD.n3504 VSS 0.131155f
C13780 DVDD.n3505 VSS 0.131155f
C13781 DVDD.n3506 VSS 0.131155f
C13782 DVDD.n3507 VSS 0.131155f
C13783 DVDD.n3508 VSS 0.131155f
C13784 DVDD.n3509 VSS 0.131155f
C13785 DVDD.n3510 VSS 0.073429f
C13786 DVDD.n3511 VSS 0.131155f
C13787 DVDD.n3512 VSS 0.131155f
C13788 DVDD.n3513 VSS 0.131155f
C13789 DVDD.n3514 VSS 0.131155f
C13790 DVDD.n3515 VSS 0.131155f
C13791 DVDD.n3516 VSS 0.131155f
C13792 DVDD.n3517 VSS 0.131155f
C13793 DVDD.n3518 VSS 0.131155f
C13794 DVDD.n3519 VSS 0.131155f
C13795 DVDD.n3520 VSS 0.131155f
C13796 DVDD.n3521 VSS 0.131155f
C13797 DVDD.n3522 VSS 0.131155f
C13798 DVDD.n3523 VSS 0.131155f
C13799 DVDD.n3524 VSS 0.131155f
C13800 DVDD.n3525 VSS 0.071581f
C13801 DVDD.n3526 VSS 0.065578f
C13802 DVDD.n3527 VSS 0.01425f
C13803 DVDD.n3528 VSS 0.065578f
C13804 DVDD.n3529 VSS 0.125152f
C13805 DVDD.n3530 VSS 0.131155f
C13806 DVDD.n3531 VSS 0.131155f
C13807 DVDD.n3532 VSS 0.131155f
C13808 DVDD.n3533 VSS 0.131155f
C13809 DVDD.n3534 VSS 0.131155f
C13810 DVDD.n3535 VSS 0.131155f
C13811 DVDD.n3536 VSS 0.131155f
C13812 DVDD.n3537 VSS 0.131155f
C13813 DVDD.n3538 VSS 0.131155f
C13814 DVDD.n3539 VSS 0.131155f
C13815 DVDD.n3540 VSS 0.131155f
C13816 DVDD.n3541 VSS 0.131155f
C13817 DVDD.n3542 VSS 0.131155f
C13818 DVDD.n3543 VSS 0.131155f
C13819 DVDD.n3544 VSS 0.131155f
C13820 DVDD.n3545 VSS 0.131155f
C13821 DVDD.n3546 VSS 0.131155f
C13822 DVDD.n3547 VSS 0.131155f
C13823 DVDD.n3548 VSS 0.131155f
C13824 DVDD.n3549 VSS 0.131155f
C13825 DVDD.n3550 VSS 0.131155f
C13826 DVDD.n3551 VSS 0.131155f
C13827 DVDD.n3552 VSS 0.131155f
C13828 DVDD.n3553 VSS 0.131155f
C13829 DVDD.n3554 VSS 0.131155f
C13830 DVDD.n3555 VSS 0.131155f
C13831 DVDD.n3556 VSS 0.131155f
C13832 DVDD.n3557 VSS 0.131155f
C13833 DVDD.n3558 VSS 0.131155f
C13834 DVDD.n3559 VSS 0.131155f
C13835 DVDD.n3560 VSS 0.131155f
C13836 DVDD.n3561 VSS 0.131155f
C13837 DVDD.n3562 VSS 0.131155f
C13838 DVDD.n3563 VSS 0.131155f
C13839 DVDD.n3564 VSS 0.131155f
C13840 DVDD.n3565 VSS 0.131155f
C13841 DVDD.n3566 VSS 0.131155f
C13842 DVDD.n3567 VSS 0.131155f
C13843 DVDD.n3568 VSS 0.131155f
C13844 DVDD.n3569 VSS 0.131155f
C13845 DVDD.n3570 VSS 0.131155f
C13846 DVDD.n3571 VSS 0.131155f
C13847 DVDD.n3572 VSS 0.131155f
C13848 DVDD.n3573 VSS 0.131155f
C13849 DVDD.n3574 VSS 0.131155f
C13850 DVDD.n3575 VSS 0.131155f
C13851 DVDD.n3576 VSS 0.131155f
C13852 DVDD.n3577 VSS 0.131155f
C13853 DVDD.n3578 VSS 0.131155f
C13854 DVDD.n3579 VSS 0.131155f
C13855 DVDD.n3580 VSS 0.131155f
C13856 DVDD.n3581 VSS 0.131155f
C13857 DVDD.n3582 VSS 0.131155f
C13858 DVDD.n3583 VSS 0.131155f
C13859 DVDD.n3584 VSS 0.131155f
C13860 DVDD.n3585 VSS 0.131155f
C13861 DVDD.n3586 VSS 0.131155f
C13862 DVDD.n3587 VSS 0.131155f
C13863 DVDD.n3588 VSS 0.131155f
C13864 DVDD.n3589 VSS 0.131155f
C13865 DVDD.n3590 VSS 0.131155f
C13866 DVDD.n3591 VSS 0.131155f
C13867 DVDD.n3592 VSS 0.131155f
C13868 DVDD.n3593 VSS 0.131155f
C13869 DVDD.n3594 VSS 0.131155f
C13870 DVDD.n3595 VSS 0.131155f
C13871 DVDD.n3596 VSS 0.131155f
C13872 DVDD.n3597 VSS 0.131155f
C13873 DVDD.n3598 VSS 0.131155f
C13874 DVDD.n3599 VSS 0.131155f
C13875 DVDD.n3600 VSS 0.123305f
C13876 DVDD.n3601 VSS 0.065578f
C13877 DVDD.n3602 VSS 0.027639f
C13878 DVDD.n3603 VSS 0.065578f
C13879 DVDD.n3604 VSS 0.065578f
C13880 DVDD.n3605 VSS 0.131155f
C13881 DVDD.n3606 VSS 0.131155f
C13882 DVDD.n3607 VSS 0.131155f
C13883 DVDD.n3608 VSS 0.131155f
C13884 DVDD.n3609 VSS 0.131155f
C13885 DVDD.n3610 VSS 0.131155f
C13886 DVDD.n3611 VSS 0.131155f
C13887 DVDD.n3612 VSS 0.131155f
C13888 DVDD.n3613 VSS 0.131155f
C13889 DVDD.n3614 VSS 0.131155f
C13890 DVDD.n3615 VSS 0.131155f
C13891 DVDD.n3616 VSS 0.131155f
C13892 DVDD.n3617 VSS 0.131155f
C13893 DVDD.n3618 VSS 0.119148f
C13894 DVDD.n3619 VSS 0.131155f
C13895 DVDD.n3620 VSS 0.131155f
C13896 DVDD.n3621 VSS 0.131155f
C13897 DVDD.n3622 VSS 0.131155f
C13898 DVDD.n3623 VSS 0.131155f
C13899 DVDD.n3624 VSS 0.131155f
C13900 DVDD.n3625 VSS 0.131155f
C13901 DVDD.n3626 VSS 0.131155f
C13902 DVDD.n3627 VSS 0.131155f
C13903 DVDD.n3628 VSS 0.131155f
C13904 DVDD.n3629 VSS 0.131155f
C13905 DVDD.n3630 VSS 0.131155f
C13906 DVDD.n3631 VSS 0.131155f
C13907 DVDD.n3632 VSS 0.131155f
C13908 DVDD.n3633 VSS 0.131155f
C13909 DVDD.n3634 VSS 0.131155f
C13910 DVDD.n3635 VSS 0.131155f
C13911 DVDD.n3636 VSS 0.131155f
C13912 DVDD.n3637 VSS 0.131155f
C13913 DVDD.n3638 VSS 0.131155f
C13914 DVDD.n3639 VSS 0.131155f
C13915 DVDD.n3640 VSS 0.131155f
C13916 DVDD.n3641 VSS 0.131155f
C13917 DVDD.n3642 VSS 0.131155f
C13918 DVDD.n3643 VSS 0.131155f
C13919 DVDD.n3644 VSS 0.131155f
C13920 DVDD.n3645 VSS 0.131155f
C13921 DVDD.n3646 VSS 0.131155f
C13922 DVDD.n3647 VSS 0.131155f
C13923 DVDD.n3648 VSS 0.131155f
C13924 DVDD.n3649 VSS 0.131155f
C13925 DVDD.n3650 VSS 0.131155f
C13926 DVDD.n3651 VSS 0.131155f
C13927 DVDD.n3652 VSS 0.131155f
C13928 DVDD.n3653 VSS 0.131155f
C13929 DVDD.n3654 VSS 0.131155f
C13930 DVDD.n3655 VSS 0.131155f
C13931 DVDD.n3656 VSS 0.131155f
C13932 DVDD.n3657 VSS 0.131155f
C13933 DVDD.n3658 VSS 0.131155f
C13934 DVDD.n3659 VSS 0.131155f
C13935 DVDD.n3660 VSS 0.131155f
C13936 DVDD.n3661 VSS 0.131155f
C13937 DVDD.n3662 VSS 0.131155f
C13938 DVDD.n3663 VSS 0.131155f
C13939 DVDD.n3664 VSS 0.485997f
C13940 DVDD.n3665 VSS 0.250567f
C13941 DVDD.n3666 VSS 0.131155f
C13942 DVDD.n3667 VSS 0.065578f
C13943 DVDD.n3671 VSS 0.065578f
C13944 DVDD.n3673 VSS 1.00993f
C13945 DVDD.n3674 VSS 0.065578f
C13946 DVDD.n3675 VSS 0.69457f
C13947 DVDD.n3676 VSS 0.694605f
C13948 DVDD.n3677 VSS 0.068071f
C13949 DVDD.n3678 VSS 0.230494f
C13950 DVDD.n3679 VSS 0.076316f
C13951 DVDD.n3680 VSS 0.080848f
C13952 DVDD.n3681 VSS 0.040423f
C13953 DVDD.n3682 VSS 0.040423f
C13954 DVDD.n3683 VSS 0.037473f
C13955 DVDD.n3684 VSS 0.037473f
C13956 DVDD.n3685 VSS 0.037473f
C13957 DVDD.n3686 VSS 0.040423f
C13958 DVDD.n3687 VSS 0.040423f
C13959 DVDD.n3688 VSS 0.080848f
C13960 DVDD.n3689 VSS 0.061774f
C13961 DVDD.n3690 VSS 0.026759f
C13962 DVDD.n3691 VSS 1.84025f
C13963 DVDD.t16 VSS 0.010292f
C13964 DVDD.t161 VSS 0.010292f
C13965 DVDD.n3692 VSS 0.040258f
C13966 DVDD.n3693 VSS 0.047824f
C13967 DVDD.t5 VSS 0.042949f
C13968 DVDD.n3694 VSS 0.375287f
C13969 DVDD.t4 VSS 0.337801f
C13970 DVDD.t15 VSS 0.203882f
C13971 DVDD.t159 VSS 0.042949f
C13972 DVDD.n3695 VSS 0.381859f
C13973 DVDD.t158 VSS 0.335563f
C13974 DVDD.t160 VSS 0.206122f
C13975 DVDD.n3696 VSS 0.100508f
C13976 DVDD.n3697 VSS -0.035151f
C13977 DVDD.n3698 VSS 0.030756f
C13978 DVDD.n3699 VSS 0.680236f
C13979 DVDD.n3700 VSS 0.517784f
C13980 DVDD.n3701 VSS 0.36353f
C13981 DVDD.n3702 VSS 0.171201f
C13982 DVDD.n3703 VSS 0.281047f
C13983 DVDD.n3704 VSS 0.206827f
C13984 DVDD.n3705 VSS 0.206827f
C13985 DVDD.n3706 VSS 0.206827f
C13986 DVDD.n3707 VSS 1.90523f
C13987 DVDD.n3708 VSS 0.059497f
C13988 DVDD.n3709 VSS 0.059497f
C13989 DVDD.n3710 VSS 0.040423f
C13990 DVDD.n3711 VSS 0.040423f
C13991 DVDD.n3712 VSS 0.037473f
C13992 DVDD.n3713 VSS 0.037473f
C13993 DVDD.n3714 VSS 0.040423f
C13994 DVDD.n3715 VSS 0.040423f
C13995 DVDD.n3716 VSS 0.040423f
C13996 DVDD.n3717 VSS 0.080848f
C13997 DVDD.n3718 VSS 0.234902f
C13998 DVDD.n3719 VSS 0.081071f
C13999 DVDD.n3720 VSS 0.083426f
C14000 DVDD.n3721 VSS 0.907268f
C14001 DVDD.n3723 VSS 0.535669f
C14002 DVDD.n3724 VSS 0.037473f
C14003 DVDD.n3725 VSS 0.037473f
C14004 DVDD.n3726 VSS 0.037473f
C14005 DVDD.n3727 VSS 0.037473f
C14006 DVDD.n3728 VSS 0.037473f
C14007 DVDD.n3729 VSS 0.037473f
C14008 DVDD.n3730 VSS 0.037473f
C14009 DVDD.n3731 VSS 0.037473f
C14010 DVDD.n3732 VSS 0.037473f
C14011 DVDD.n3733 VSS 1.042f
C14012 DVDD.n3734 VSS 0.281047f
C14013 DVDD.n3735 VSS 0.281047f
C14014 DVDD.n3736 VSS 0.140524f
C14015 DVDD.n3737 VSS 0.037473f
C14016 DVDD.n3738 VSS 0.037473f
C14017 DVDD.n3739 VSS 0.037473f
C14018 DVDD.n3740 VSS 0.037473f
C14019 DVDD.n3741 VSS 0.037473f
C14020 DVDD.n3742 VSS 0.037473f
C14021 DVDD.n3743 VSS 0.037473f
C14022 DVDD.n3744 VSS 0.037473f
C14023 DVDD.n3754 VSS 0.140524f
C14024 DVDD.n3755 VSS 0.037473f
C14025 DVDD.n3756 VSS 0.040424f
C14026 DVDD.n3757 VSS 0.080848f
C14027 DVDD.n3758 VSS 0.080848f
C14028 DVDD.n3759 VSS 0.080848f
C14029 DVDD.n3760 VSS 0.040424f
C14030 DVDD.n3761 VSS 0.040424f
C14031 DVDD.n3762 VSS 0.040424f
C14032 DVDD.n3763 VSS 0.037473f
C14033 DVDD.n3764 VSS 0.059497f
C14034 DVDD.n3765 VSS 0.028752f
C14035 DVDD.n3766 VSS 0.040424f
C14036 DVDD.n3767 VSS 0.037473f
C14037 DVDD.n3768 VSS 0.037473f
C14038 DVDD.n3769 VSS 0.040424f
C14039 DVDD.n3770 VSS 0.040424f
C14040 DVDD.n3771 VSS 0.080848f
C14041 DVDD.n3772 VSS 0.234902f
C14042 DVDD.n3773 VSS 0.080977f
C14043 DVDD.n3774 VSS 0.066709f
C14044 DVDD.n3775 VSS 0.063791f
C14045 DVDD.n3776 VSS 0.06373f
C14046 DVDD.n3777 VSS 0.628154f
C14047 DVDD.n3778 VSS 0.907268f
C14048 DVDD.n3779 VSS 0.140524f
C14049 DVDD.n3780 VSS 0.157347f
C14050 DVDD.n3781 VSS 0.218702f
C14051 DVDD.n3782 VSS 0.281047f
C14052 DVDD.n3783 VSS 0.281047f
C14053 DVDD.n3784 VSS 0.281047f
C14054 DVDD.n3785 VSS 0.281047f
C14055 DVDD.n3786 VSS 0.281047f
C14056 DVDD.n3787 VSS 0.281047f
C14057 DVDD.n3788 VSS 0.202869f
C14058 DVDD.n3789 VSS 0.281047f
C14059 DVDD.n3790 VSS 0.281047f
C14060 DVDD.n3791 VSS 0.281047f
C14061 DVDD.n3792 VSS 0.281047f
C14062 DVDD.n3793 VSS 0.281047f
C14063 DVDD.n3794 VSS 0.281047f
C14064 DVDD.n3795 VSS 0.281047f
C14065 DVDD.n3796 VSS 0.281047f
C14066 DVDD.n3797 VSS 0.281047f
C14067 DVDD.n3798 VSS 0.281047f
C14068 DVDD.n3799 VSS 0.281047f
C14069 DVDD.n3800 VSS 0.281047f
C14070 DVDD.n3801 VSS 0.281047f
C14071 DVDD.n3802 VSS 0.281047f
C14072 DVDD.n3803 VSS 0.281047f
C14073 DVDD.n3804 VSS 0.281047f
C14074 DVDD.n3805 VSS 0.188025f
C14075 DVDD.n3806 VSS 0.188025f
C14076 DVDD.n3807 VSS 0.10061f
C14077 DVDD.n3808 VSS 0.074418f
C14078 DVDD.n3809 VSS 0.124558f
C14079 DVDD.n3810 VSS 0.149892f
C14080 DVDD.n3811 VSS 0.149892f
C14081 DVDD.n3812 VSS 0.074946f
C14082 DVDD.n3813 VSS 0.074946f
C14083 DVDD.n3814 VSS 0.074946f
C14084 DVDD.n3815 VSS 0.00712f
C14085 DVDD.n3816 VSS 0.00712f
C14086 DVDD.n3817 VSS 0.012388f
C14087 DVDD.n3818 VSS 0.074946f
C14088 DVDD.n3819 VSS 0.074946f
C14089 DVDD.n3820 VSS 0.149892f
C14090 DVDD.n3821 VSS 0.149892f
C14091 DVDD.n3822 VSS 0.149892f
C14092 DVDD.n3823 VSS 0.149892f
C14093 DVDD.n3824 VSS 0.149892f
C14094 DVDD.n3825 VSS 0.125086f
C14095 DVDD.n3826 VSS 0.149892f
C14096 DVDD.n3827 VSS 0.149892f
C14097 DVDD.n3828 VSS 0.149892f
C14098 DVDD.n3829 VSS 0.149892f
C14099 DVDD.n3830 VSS 0.149892f
C14100 DVDD.n3831 VSS 0.142503f
C14101 DVDD.n3832 VSS 0.142503f
C14102 DVDD.n3833 VSS 0.142503f
C14103 DVDD.n3834 VSS 0.169751f
C14104 DVDD.n3835 VSS 0.419531f
C14105 DVDD.n3836 VSS 0.096057f
C14106 DVDD.n3837 VSS 0.096057f
C14107 DVDD.n3838 VSS 0.096057f
C14108 DVDD.n3839 VSS 0.149892f
C14109 DVDD.n3840 VSS 0.149892f
C14110 DVDD.n3841 VSS 0.149892f
C14111 DVDD.n3842 VSS 0.149892f
C14112 DVDD.n3843 VSS 0.149892f
C14113 DVDD.n3844 VSS 0.149892f
C14114 DVDD.n3845 VSS 0.149892f
C14115 DVDD.n3846 VSS 0.149892f
C14116 DVDD.n3847 VSS 0.149892f
C14117 DVDD.n3848 VSS 0.149892f
C14118 DVDD.n3849 VSS 0.149892f
C14119 DVDD.n3850 VSS 0.149892f
C14120 DVDD.n3851 VSS 0.149892f
C14121 DVDD.n3852 VSS 0.149892f
C14122 DVDD.n3853 VSS 0.149892f
C14123 DVDD.n3854 VSS 0.149892f
C14124 DVDD.n3855 VSS 0.149892f
C14125 DVDD.n3856 VSS 0.096057f
C14126 DVDD.n3857 VSS 0.096057f
C14127 DVDD.n3858 VSS 0.096057f
C14128 DVDD.n3859 VSS 0.149892f
C14129 DVDD.n3860 VSS 0.149892f
C14130 DVDD.n3861 VSS 0.149892f
C14131 DVDD.n3862 VSS 0.149892f
C14132 DVDD.n3863 VSS 0.149892f
C14133 DVDD.n3864 VSS 0.149892f
C14134 DVDD.n3865 VSS 0.149892f
C14135 DVDD.n3866 VSS 0.149892f
C14136 DVDD.n3867 VSS 0.138281f
C14137 DVDD.n3868 VSS 0.138281f
C14138 DVDD.n3869 VSS 0.10028f
C14139 DVDD.n3870 VSS 0.167747f
C14140 DVDD.n3871 VSS 0.42034f
C14141 DVDD.n3872 VSS 0.149892f
C14142 DVDD.n3873 VSS 0.149892f
C14143 DVDD.n3874 VSS 0.149892f
C14144 DVDD.n3875 VSS 0.149892f
C14145 DVDD.n3876 VSS 0.149892f
C14146 DVDD.n3877 VSS 0.149892f
C14147 DVDD.n3878 VSS 0.149892f
C14148 DVDD.n3879 VSS 0.149892f
C14149 DVDD.n3880 VSS 0.149892f
C14150 DVDD.n3881 VSS 0.091835f
C14151 DVDD.n3882 VSS 0.149892f
C14152 DVDD.n3883 VSS 0.149892f
C14153 DVDD.n3884 VSS 0.149892f
C14154 DVDD.n3885 VSS 0.149892f
C14155 DVDD.n3886 VSS 0.149892f
C14156 DVDD.n3887 VSS 0.149892f
C14157 DVDD.n3888 VSS 0.149892f
C14158 DVDD.n3889 VSS 0.149892f
C14159 DVDD.n3890 VSS 0.149892f
C14160 DVDD.n3891 VSS 0.149892f
C14161 DVDD.n3892 VSS 0.149892f
C14162 DVDD.n3893 VSS 0.149892f
C14163 DVDD.n3894 VSS 0.149892f
C14164 DVDD.n3895 VSS 0.149892f
C14165 DVDD.n3896 VSS 0.149892f
C14166 DVDD.n3897 VSS 0.149892f
C14167 DVDD.n3898 VSS 0.149892f
C14168 DVDD.n3899 VSS 0.149892f
C14169 DVDD.n3900 VSS 0.10028f
C14170 DVDD.n3901 VSS 0.10028f
C14171 DVDD.n3902 VSS 0.179572f
C14172 DVDD.n3903 VSS 0.169743f
C14173 DVDD.n3904 VSS 0.436959f
C14174 DVDD.n3905 VSS 0.138281f
C14175 DVDD.n3906 VSS 0.149892f
C14176 DVDD.n3907 VSS 0.149892f
C14177 DVDD.n3908 VSS 0.149892f
C14178 DVDD.n3909 VSS 0.149892f
C14179 DVDD.n3910 VSS 0.149892f
C14180 DVDD.n3911 VSS 0.149892f
C14181 DVDD.n3912 VSS 0.149892f
C14182 DVDD.n3913 VSS 0.149892f
C14183 DVDD.n3914 VSS 0.149892f
C14184 DVDD.n3915 VSS 0.149892f
C14185 DVDD.n3916 VSS 0.149892f
C14186 DVDD.n3917 VSS 0.149892f
C14187 DVDD.n3918 VSS 0.149892f
C14188 DVDD.n3919 VSS 0.149892f
C14189 DVDD.n3920 VSS 0.149892f
C14190 DVDD.n3921 VSS 0.149892f
C14191 DVDD.n3922 VSS 0.12878f
C14192 DVDD.n3923 VSS 0.12878f
C14193 DVDD.n3924 VSS 0.12878f
C14194 DVDD.n3925 VSS 0.216021f
C14195 DVDD.n3926 VSS 0.281047f
C14196 DVDD.n3927 VSS 0.281047f
C14197 DVDD.n3928 VSS 0.281047f
C14198 DVDD.n3929 VSS 0.194952f
C14199 DVDD.t157 VSS 0.041167f
C14200 DVDD.t120 VSS 0.041167f
C14201 DVDD.n3930 VSS 0.082335f
C14202 DVDD.n3931 VSS 0.102524f
C14203 DVDD.n3932 VSS 0.04694f
C14204 DVDD.t36 VSS 0.041167f
C14205 DVDD.t42 VSS 0.041167f
C14206 DVDD.n3933 VSS 0.082335f
C14207 DVDD.n3934 VSS 0.102524f
C14208 DVDD.t217 VSS 0.032179f
C14209 DVDD.n3935 VSS 0.212765f
C14210 DVDD.n3936 VSS 0.281047f
C14211 DVDD.n3937 VSS 0.281047f
C14212 DVDD.n3938 VSS 0.281047f
C14213 DVDD.n3939 VSS 0.281047f
C14214 DVDD.n3940 VSS 0.281047f
C14215 DVDD.n3941 VSS 0.281047f
C14216 DVDD.n3942 VSS 0.281047f
C14217 DVDD.n3943 VSS 0.281047f
C14218 DVDD.n3944 VSS 0.281047f
C14219 DVDD.n3945 VSS 0.281047f
C14220 DVDD.n3946 VSS 0.281047f
C14221 DVDD.n3947 VSS 0.281047f
C14222 DVDD.n3948 VSS 0.281047f
C14223 DVDD.n3949 VSS 0.281047f
C14224 DVDD.n3950 VSS 0.281047f
C14225 DVDD.n3951 VSS 0.281047f
C14226 DVDD.n3952 VSS 0.281047f
C14227 DVDD.n3953 VSS 0.147451f
C14228 DVDD.n3954 VSS 0.216021f
C14229 DVDD.n3955 VSS 0.27412f
C14230 DVDD.n3956 VSS 0.281047f
C14231 DVDD.n3957 VSS 0.281047f
C14232 DVDD.n3958 VSS 0.281047f
C14233 DVDD.n3959 VSS 0.208806f
C14234 DVDD.n3960 VSS 0.152357f
C14235 DVDD.n3961 VSS 0.163921f
C14236 DVDD.t38 VSS 0.09794f
C14237 DVDD.n3962 VSS 0.125601f
C14238 DVDD.n3963 VSS 0.051157f
C14239 DVDD.n3964 VSS 0.055913f
C14240 DVDD.n3965 VSS 0.054298f
C14241 DVDD.t40 VSS 0.09794f
C14242 DVDD.n3966 VSS 0.143921f
C14243 DVDD.n3967 VSS 0.216021f
C14244 DVDD.n3968 VSS 0.226619f
C14245 DVDD.n3969 VSS 0.185056f
C14246 DVDD.n3970 VSS 0.281047f
C14247 DVDD.n3971 VSS 0.281047f
C14248 DVDD.n3972 VSS 0.281047f
C14249 DVDD.n3973 VSS 0.281047f
C14250 DVDD.n3974 VSS 0.180108f
C14251 DVDD.n3975 VSS 0.180108f
C14252 DVDD.n3976 VSS 0.135576f
C14253 DVDD.n3977 VSS 0.21547f
C14254 DVDD.n3978 VSS 0.241463f
C14255 DVDD.n3979 VSS 0.241463f
C14256 DVDD.n3980 VSS 0.241463f
C14257 DVDD.n3981 VSS 0.281047f
C14258 DVDD.n3982 VSS 0.281047f
C14259 DVDD.n3983 VSS 0.281047f
C14260 DVDD.n3984 VSS 0.281047f
C14261 DVDD.n3985 VSS 0.281047f
C14262 DVDD.n3986 VSS 0.281047f
C14263 DVDD.n3987 VSS 0.281047f
C14264 DVDD.n3988 VSS 0.281047f
C14265 DVDD.n3989 VSS 0.281047f
C14266 DVDD.n3990 VSS 0.281047f
C14267 DVDD.n3991 VSS 0.281047f
C14268 DVDD.n3992 VSS 0.281047f
C14269 DVDD.n3993 VSS 0.281047f
C14270 DVDD.n3994 VSS 0.068295f
C14271 DVDD.t46 VSS 0.041167f
C14272 DVDD.t44 VSS 0.041167f
C14273 DVDD.n3995 VSS 0.082335f
C14274 DVDD.n3996 VSS 0.13166f
C14275 DVDD.n3997 VSS 0.218072f
C14276 DVDD.n3998 VSS 0.157347f
C14277 DVDD.n3999 VSS 0.281047f
C14278 DVDD.n4000 VSS 0.281047f
C14279 DVDD.n4001 VSS 0.281047f
C14280 DVDD.n4002 VSS 0.281047f
C14281 DVDD.n4003 VSS 0.281047f
C14282 DVDD.n4004 VSS 0.281047f
C14283 DVDD.n4005 VSS 0.281047f
C14284 DVDD.n4006 VSS 0.281047f
C14285 DVDD.n4007 VSS 0.281047f
C14286 DVDD.n4008 VSS 0.281047f
C14287 DVDD.n4009 VSS 0.281047f
C14288 DVDD.n4010 VSS 0.281047f
C14289 DVDD.n4011 VSS 0.281047f
C14290 DVDD.n4012 VSS 0.268182f
C14291 DVDD.n4013 VSS 0.068295f
C14292 DVDD.t203 VSS 0.041167f
C14293 DVDD.t99 VSS 0.041167f
C14294 DVDD.n4014 VSS 0.082335f
C14295 DVDD.n4015 VSS 0.13166f
C14296 DVDD.n4016 VSS 0.218072f
C14297 DVDD.n4017 VSS 0.153388f
C14298 DVDD.n4018 VSS 0.281047f
C14299 DVDD.n4019 VSS 0.281047f
C14300 DVDD.n4020 VSS 0.281047f
C14301 DVDD.n4021 VSS 0.281047f
C14302 DVDD.n4022 VSS 0.281047f
C14303 DVDD.n4023 VSS 0.281047f
C14304 DVDD.n4024 VSS 0.281047f
C14305 DVDD.n4025 VSS 0.281047f
C14306 DVDD.n4026 VSS 0.281047f
C14307 DVDD.n4027 VSS 0.281047f
C14308 DVDD.n4028 VSS 0.281047f
C14309 DVDD.n4029 VSS 0.281047f
C14310 DVDD.n4030 VSS 0.281047f
C14311 DVDD.n4031 VSS 0.281047f
C14312 DVDD.n4032 VSS 0.281047f
C14313 DVDD.n4033 VSS 0.172191f
C14314 DVDD.n4034 VSS 0.172191f
C14315 DVDD.n4035 VSS 0.21547f
C14316 DVDD.n4036 VSS 0.149892f
C14317 DVDD.n4037 VSS 0.149892f
C14318 DVDD.n4038 VSS 0.149892f
C14319 DVDD.n4039 VSS 0.149892f
C14320 DVDD.n4040 VSS 0.149892f
C14321 DVDD.n4041 VSS 0.149892f
C14322 DVDD.n4042 VSS 0.134058f
C14323 DVDD.n4043 VSS 0.134058f
C14324 DVDD.n4044 VSS 0.104502f
C14325 DVDD.n4045 VSS 0.167854f
C14326 DVDD.n4046 VSS 0.179314f
C14327 DVDD.n4047 VSS 0.149892f
C14328 DVDD.n4048 VSS 0.149892f
C14329 DVDD.n4049 VSS 0.098169f
C14330 DVDD.n4050 VSS 0.149892f
C14331 DVDD.n4051 VSS 0.149892f
C14332 DVDD.n4052 VSS 0.149892f
C14333 DVDD.n4053 VSS 0.149892f
C14334 DVDD.n4054 VSS 0.075143f
C14335 DVDD.n4055 VSS 0.074946f
C14336 DVDD.n4056 VSS 0.00712f
C14337 DVDD.n4057 VSS 0.074946f
C14338 DVDD.n4058 VSS 0.074946f
C14339 DVDD.n4059 VSS 0.074946f
C14340 DVDD.n4060 VSS 0.149892f
C14341 DVDD.n4061 VSS 0.149892f
C14342 DVDD.n4062 VSS 0.149892f
C14343 DVDD.n4063 VSS 0.149892f
C14344 DVDD.n4064 VSS 0.074946f
C14345 DVDD.n4065 VSS 0.074946f
C14346 DVDD.n4066 VSS 0.00712f
C14347 DVDD.n4067 VSS 0.012388f
C14348 DVDD.n4068 VSS 0.074946f
C14349 DVDD.n4069 VSS 0.074946f
C14350 DVDD.n4070 VSS 0.149892f
C14351 DVDD.n4071 VSS 0.149892f
C14352 DVDD.n4072 VSS 0.149892f
C14353 DVDD.n4073 VSS 0.149892f
C14354 DVDD.n4074 VSS 0.149892f
C14355 DVDD.n4075 VSS 0.149892f
C14356 DVDD.n4076 VSS 0.149892f
C14357 DVDD.n4077 VSS 0.149892f
C14358 DVDD.n4078 VSS 0.149892f
C14359 DVDD.n4079 VSS 0.104502f
C14360 DVDD.n4080 VSS 0.104502f
C14361 DVDD.n4081 VSS 0.436898f
C14362 DVDD.n4082 VSS 0.169743f
C14363 DVDD.n4083 VSS 0.420551f
C14364 DVDD.n4084 VSS 0.134058f
C14365 DVDD.n4085 VSS 0.149892f
C14366 DVDD.n4086 VSS 0.149892f
C14367 DVDD.n4087 VSS 0.149892f
C14368 DVDD.n4088 VSS 0.149892f
C14369 DVDD.n4089 VSS 0.149892f
C14370 DVDD.n4090 VSS 0.149892f
C14371 DVDD.n4091 VSS 0.149892f
C14372 DVDD.n4092 VSS 0.149892f
C14373 DVDD.n4093 VSS 0.149892f
C14374 DVDD.n4094 VSS 0.149892f
C14375 DVDD.n4095 VSS 0.149892f
C14376 DVDD.n4096 VSS 0.149892f
C14377 DVDD.n4097 VSS 0.149892f
C14378 DVDD.n4098 VSS 0.149892f
C14379 DVDD.n4099 VSS 0.149892f
C14380 DVDD.n4100 VSS 0.149892f
C14381 DVDD.n4101 VSS 0.133003f
C14382 DVDD.n4102 VSS 0.133003f
C14383 DVDD.n4103 VSS 0.133003f
C14384 DVDD.n4104 VSS 0.21547f
C14385 DVDD.n4105 VSS 0.24938f
C14386 DVDD.n4106 VSS 0.281047f
C14387 DVDD.n4107 VSS 0.281047f
C14388 DVDD.n4108 VSS 0.281047f
C14389 DVDD.n4109 VSS 0.281047f
C14390 DVDD.n4110 VSS 0.281047f
C14391 DVDD.n4111 VSS 0.281047f
C14392 DVDD.n4112 VSS 0.281047f
C14393 DVDD.n4113 VSS 0.281047f
C14394 DVDD.n4114 VSS 0.190993f
C14395 DVDD.n4115 VSS 0.216021f
C14396 DVDD.n4116 VSS 0.230578f
C14397 DVDD.n4117 VSS 0.281047f
C14398 DVDD.n4118 VSS 0.281047f
C14399 DVDD.n4119 VSS 0.281047f
C14400 DVDD.n4120 VSS 0.181097f
C14401 DVDD.n4121 VSS 0.216021f
C14402 DVDD.t128 VSS 0.041167f
C14403 DVDD.t155 VSS 0.041167f
C14404 DVDD.n4122 VSS 0.082335f
C14405 DVDD.n4123 VSS 0.102524f
C14406 DVDD.n4124 VSS 0.04694f
C14407 DVDD.n4125 VSS 0.054298f
C14408 DVDD.n4126 VSS 0.055913f
C14409 DVDD.t138 VSS 0.041167f
C14410 DVDD.t122 VSS 0.041167f
C14411 DVDD.n4127 VSS 0.082335f
C14412 DVDD.n4128 VSS 0.102524f
C14413 DVDD.n4129 VSS 0.216021f
C14414 DVDD.n4130 VSS 0.151409f
C14415 DVDD.n4131 VSS 0.281047f
C14416 DVDD.n4132 VSS 0.281047f
C14417 DVDD.n4133 VSS 0.281047f
C14418 DVDD.n4134 VSS 0.281047f
C14419 DVDD.n4135 VSS 0.281047f
C14420 DVDD.n4136 VSS 0.281047f
C14421 DVDD.n4137 VSS 0.212765f
C14422 DVDD.t124 VSS 0.09794f
C14423 DVDD.n4138 VSS 0.125601f
C14424 DVDD.t205 VSS 0.032179f
C14425 DVDD.n4139 VSS 0.163921f
C14426 DVDD.n4140 VSS 0.152357f
C14427 DVDD.n4141 VSS 0.167243f
C14428 DVDD.n4142 VSS 0.208806f
C14429 DVDD.n4143 VSS 0.281047f
C14430 DVDD.n4144 VSS 0.281047f
C14431 DVDD.n4145 VSS 0.281047f
C14432 DVDD.n4146 VSS 0.281047f
C14433 DVDD.n4147 VSS 0.281047f
C14434 DVDD.n4148 VSS 0.235526f
C14435 DVDD.t210 VSS 0.032179f
C14436 DVDD.n4149 VSS 0.163921f
C14437 DVDD.n4150 VSS 0.152357f
C14438 DVDD.n4151 VSS 0.159326f
C14439 DVDD.n4152 VSS 0.281047f
C14440 DVDD.n4153 VSS 0.281047f
C14441 DVDD.n4154 VSS 0.281047f
C14442 DVDD.n4155 VSS 0.281047f
C14443 DVDD.n4156 VSS 0.281047f
C14444 DVDD.n4157 VSS 0.281047f
C14445 DVDD.n4158 VSS 0.183077f
C14446 DVDD.n4159 VSS 0.216021f
C14447 DVDD.n4160 VSS 0.238494f
C14448 DVDD.n4161 VSS 0.244432f
C14449 DVDD.n4162 VSS 0.281047f
C14450 DVDD.n4163 VSS 0.281047f
C14451 DVDD.n4164 VSS 0.281047f
C14452 DVDD.n4165 VSS 0.281047f
C14453 DVDD.n4166 VSS 0.281047f
C14454 DVDD.n4167 VSS 0.281047f
C14455 DVDD.n4168 VSS 0.177139f
C14456 DVDD.n4169 VSS 0.281047f
C14457 DVDD.n4170 VSS 0.164274f
C14458 DVDD.n4171 VSS 0.164274f
C14459 DVDD.n4172 VSS 0.164274f
C14460 DVDD.n4173 VSS 0.281047f
C14461 DVDD.n4174 VSS 0.281047f
C14462 DVDD.t153 VSS 0.041167f
C14463 DVDD.t145 VSS 0.041167f
C14464 DVDD.n4175 VSS 0.082335f
C14465 DVDD.n4176 VSS 0.130607f
C14466 DVDD.n4177 VSS 0.194322f
C14467 DVDD.n4178 VSS 0.281047f
C14468 DVDD.n4179 VSS 0.281047f
C14469 DVDD.n4180 VSS 0.281047f
C14470 DVDD.n4181 VSS 0.281047f
C14471 DVDD.n4182 VSS 0.281047f
C14472 DVDD.n4183 VSS 0.281047f
C14473 DVDD.n4184 VSS 0.281047f
C14474 DVDD.n4185 VSS 0.281047f
C14475 DVDD.n4186 VSS 0.281047f
C14476 DVDD.n4187 VSS 0.281047f
C14477 DVDD.n4188 VSS 0.281047f
C14478 DVDD.n4189 VSS 0.187035f
C14479 DVDD.n4190 VSS -0.065036f
C14480 DVDD.n4191 VSS 0.262245f
C14481 DVDD.n4192 VSS 0.281047f
C14482 DVDD.n4193 VSS 0.253338f
C14483 DVDD.n4194 VSS 0.281047f
C14484 DVDD.n4195 VSS 0.144482f
C14485 DVDD.n4196 VSS 0.168233f
C14486 DVDD.n4197 VSS 0.168233f
C14487 DVDD.n4198 VSS 0.440119f
C14488 DVDD.n4199 VSS 1.00987f
C14489 DVDD.n4200 VSS 1.24213f
C14490 DVDD.t186 VSS 0.517068f
C14491 DVDD.t71 VSS 0.480029f
C14492 DVDD.t73 VSS 0.480029f
C14493 DVDD.t69 VSS 0.649219f
C14494 DVDD.t152 VSS 0.649219f
C14495 DVDD.t144 VSS 0.382474f
C14496 DVDD.t198 VSS 0.649219f
C14497 DVDD.t25 VSS 0.649219f
C14498 DVDD.t22 VSS 0.480029f
C14499 DVDD.t125 VSS 0.343299f
C14500 DVDD.n4201 VSS 0.500617f
C14501 DVDD.t115 VSS 0.492136f
C14502 DVDD.n4202 VSS 0.584907f
C14503 DVDD.n4203 VSS 0.067926f
C14504 DVDD.t126 VSS 0.041167f
C14505 DVDD.t116 VSS 0.041167f
C14506 DVDD.n4204 VSS 0.082335f
C14507 DVDD.n4205 VSS 0.13166f
C14508 DVDD.n4206 VSS 0.218072f
C14509 DVDD.n4207 VSS 0.206827f
C14510 DVDD.n4208 VSS 0.281047f
C14511 DVDD.n4209 VSS 0.281047f
C14512 DVDD.n4210 VSS 0.281047f
C14513 DVDD.n4211 VSS 0.281047f
C14514 DVDD.n4212 VSS 0.281047f
C14515 DVDD.n4213 VSS 0.281047f
C14516 DVDD.n4214 VSS 0.281047f
C14517 DVDD.n4215 VSS 0.281047f
C14518 DVDD.n4216 VSS 0.281047f
C14519 DVDD.n4217 VSS 0.281047f
C14520 DVDD.n4218 VSS 0.281047f
C14521 DVDD.n4219 VSS 0.281047f
C14522 DVDD.n4220 VSS 0.187035f
C14523 DVDD.n4221 VSS 0.257297f
C14524 DVDD.n4222 VSS 0.257297f
C14525 DVDD.n4223 VSS 0.21547f
C14526 DVDD.n4224 VSS 0.087613f
C14527 DVDD.n4225 VSS 0.087613f
C14528 DVDD.n4226 VSS 0.06439f
C14529 DVDD.n4227 VSS 0.074946f
C14530 DVDD.n4228 VSS 0.00534f
C14531 DVDD.n4229 VSS 0.00356f
C14532 DVDD.n4230 VSS 0.010429f
C14533 DVDD.n4231 VSS 0.050716f
C14534 DVDD.n4232 VSS 0.057276f
C14535 DVDD.n4233 VSS 0.051934f
C14536 DVDD.n4234 VSS 0.038425f
C14537 DVDD.n4235 VSS 0.018029f
C14538 DVDD.n4236 VSS 0.624638f
C14539 DVDD.t123 VSS 0.594134f
C14540 DVDD.t121 VSS 0.480029f
C14541 DVDD.t137 VSS 0.480029f
C14542 DVDD.t135 VSS 0.649219f
C14543 DVDD.t154 VSS 0.649219f
C14544 DVDD.t127 VSS 0.382474f
C14545 DVDD.t76 VSS 0.649219f
C14546 DVDD.t20 VSS 0.649219f
C14547 DVDD.t1 VSS 0.480029f
C14548 DVDD.t98 VSS 0.480029f
C14549 DVDD.t202 VSS 0.594134f
C14550 DVDD.n4237 VSS 1.13375f
C14551 DVDD.t43 VSS 0.594134f
C14552 DVDD.t45 VSS 0.480029f
C14553 DVDD.t14 VSS 0.480029f
C14554 DVDD.t19 VSS 0.649219f
C14555 DVDD.t75 VSS 0.649219f
C14556 DVDD.t119 VSS 0.382474f
C14557 DVDD.t156 VSS 0.649219f
C14558 DVDD.t39 VSS 0.649219f
C14559 DVDD.t41 VSS 0.480029f
C14560 DVDD.t35 VSS 0.480029f
C14561 DVDD.t37 VSS 0.594134f
C14562 DVDD.n4238 VSS 0.624638f
C14563 DVDD.n4239 VSS 0.018029f
C14564 DVDD.n4240 VSS 0.237835f
C14565 DVDD.n4241 VSS 0.235526f
C14566 DVDD.n4242 VSS 0.281047f
C14567 DVDD.n4243 VSS 0.281047f
C14568 DVDD.n4244 VSS 0.281047f
C14569 DVDD.n4245 VSS 0.281047f
C14570 DVDD.n4246 VSS 0.281047f
C14571 DVDD.n4247 VSS 0.179118f
C14572 DVDD.n4248 VSS 0.281047f
C14573 DVDD.n4249 VSS 0.281047f
C14574 DVDD.n4250 VSS 0.242453f
C14575 DVDD.n4251 VSS 0.281047f
C14576 DVDD.n4252 VSS 0.240474f
C14577 DVDD.n4253 VSS 0.281047f
C14578 DVDD.n4254 VSS 0.281047f
C14579 DVDD.n4255 VSS 0.181097f
C14580 DVDD.n4256 VSS 0.281047f
C14581 DVDD.n4257 VSS 0.230578f
C14582 DVDD.n4258 VSS 0.233546f
C14583 DVDD.n4259 VSS 0.233546f
C14584 DVDD.n4260 VSS 0.21547f
C14585 DVDD.n4261 VSS 0.10028f
C14586 DVDD.n4262 VSS 0.10028f
C14587 DVDD.n4263 VSS 0.074946f
C14588 DVDD.n4264 VSS 0.074946f
C14589 DVDD.n4265 VSS 0.00712f
C14590 DVDD.n4266 VSS 0.00712f
C14591 DVDD.n4267 VSS 0.074946f
C14592 DVDD.n4268 VSS 0.074946f
C14593 DVDD.n4269 VSS 0.149892f
C14594 DVDD.n4270 VSS 0.149892f
C14595 DVDD.n4271 VSS 0.149892f
C14596 DVDD.n4272 VSS 0.149892f
C14597 DVDD.n4273 VSS 0.149892f
C14598 DVDD.n4274 VSS 0.099752f
C14599 DVDD.n4275 VSS 0.149892f
C14600 DVDD.n4276 VSS 0.149892f
C14601 DVDD.n4277 VSS 0.149892f
C14602 DVDD.n4278 VSS 0.149892f
C14603 DVDD.n4279 VSS 0.149892f
C14604 DVDD.n4280 VSS 0.149892f
C14605 DVDD.n4281 VSS 0.149892f
C14606 DVDD.n4282 VSS 0.149892f
C14607 DVDD.n4283 VSS 0.149892f
C14608 DVDD.n4284 VSS 0.091835f
C14609 DVDD.n4285 VSS 0.091835f
C14610 DVDD.n4286 VSS 0.091835f
C14611 DVDD.n4287 VSS 0.057312f
C14612 DVDD.n4288 VSS 0.061774f
C14613 DVDD.n4289 VSS 0.061774f
C14614 DVDD.n4290 VSS 0.040424f
C14615 DVDD.n4291 VSS 0.040424f
C14616 DVDD.n4292 VSS 0.037473f
C14617 DVDD.n4293 VSS 0.037473f
C14618 DVDD.n4294 VSS 0.040424f
C14619 DVDD.n4295 VSS 0.040424f
C14620 DVDD.n4296 VSS 0.040424f
C14621 DVDD.n4297 VSS 0.080848f
C14622 DVDD.n4298 VSS 0.230494f
C14623 DVDD.n4299 VSS 0.076483f
C14624 DVDD.n4300 VSS 0.083029f
C14625 DVDD.n4301 VSS 0.274846f
C14626 DVDD.n4302 VSS 0.535669f
C14627 DVDD.n4303 VSS 1.042f
C14628 DVDD.n4304 VSS 0.281047f
C14629 DVDD.n4305 VSS 0.281047f
C14630 DVDD.n4306 VSS 0.281047f
C14631 DVDD.n4307 VSS 0.281047f
C14632 DVDD.n4308 VSS 0.281047f
C14633 DVDD.n4309 VSS 0.281047f
C14634 DVDD.n4310 VSS 0.281047f
C14635 DVDD.n4311 VSS 0.281047f
C14636 DVDD.n4312 VSS 0.281047f
C14637 DVDD.n4313 VSS 0.190004f
C14638 DVDD.n4314 VSS 0.281047f
C14639 DVDD.n4315 VSS 0.281047f
C14640 DVDD.n4316 VSS 0.281047f
C14641 DVDD.n4317 VSS 0.281047f
C14642 DVDD.n4318 VSS 0.281047f
C14643 DVDD.n4319 VSS 0.281047f
C14644 DVDD.n4320 VSS 0.281047f
C14645 DVDD.n4321 VSS 0.281047f
C14646 DVDD.n4322 VSS 0.281047f
C14647 DVDD.n4323 VSS 0.281047f
C14648 DVDD.n4324 VSS 0.281047f
C14649 DVDD.n4325 VSS 0.281047f
C14650 DVDD.n4326 VSS 0.281047f
C14651 DVDD.n4327 VSS 0.281047f
C14652 DVDD.n4328 VSS 0.281047f
C14653 DVDD.n4329 VSS 0.281047f
C14654 DVDD.n4330 VSS 0.281047f
C14655 DVDD.n4331 VSS 0.281047f
C14656 DVDD.n4332 VSS 0.140524f
C14657 DVDD.n4342 VSS 0.140524f
C14658 DVDD.n4344 VSS 0.274846f
C14659 DVDD.n4345 VSS 0.140524f
C14660 DVDD.n4346 VSS 0.066237f
C14661 DVDD.n4347 VSS 0.535669f
C14662 DVDD.n4348 VSS 1.042f
C14663 DVDD.n4349 VSS 0.281047f
C14664 DVDD.n4350 VSS 0.281047f
C14665 DVDD.n4351 VSS 0.281047f
C14666 DVDD.n4352 VSS 0.281047f
C14667 DVDD.n4353 VSS 0.281047f
C14668 DVDD.n4354 VSS 0.281047f
C14669 DVDD.n4355 VSS 0.281047f
C14670 DVDD.n4356 VSS 0.281047f
C14671 DVDD.n4357 VSS 0.281047f
C14672 DVDD.n4358 VSS 0.281047f
C14673 DVDD.n4359 VSS 0.281047f
C14674 DVDD.n4360 VSS 0.281047f
C14675 DVDD.n4361 VSS 0.281047f
C14676 DVDD.n4362 VSS 0.281047f
C14677 DVDD.n4363 VSS 0.281047f
C14678 DVDD.n4364 VSS 0.281047f
C14679 DVDD.n4365 VSS 0.281047f
C14680 DVDD.n4366 VSS 0.281047f
C14681 DVDD.n4367 VSS 0.281047f
C14682 DVDD.n4368 VSS 0.281047f
C14683 DVDD.n4369 VSS 0.281047f
C14684 DVDD.n4370 VSS 0.281047f
C14685 DVDD.n4371 VSS 0.281047f
C14686 DVDD.n4372 VSS 0.281047f
C14687 DVDD.n4373 VSS 0.281047f
C14688 DVDD.n4374 VSS 0.281047f
C14689 DVDD.n4375 VSS 0.140524f
C14690 DVDD.n4385 VSS 0.140524f
C14691 DVDD.n4387 VSS 0.066237f
C14692 DVDD.n4388 VSS 0.140524f
C14693 DVDD.n4389 VSS 0.066237f
C14694 DVDD.n4400 VSS 0.140524f
C14695 DVDD.n4401 VSS 0.535669f
C14696 DVDD.n4411 VSS 0.281047f
C14697 DVDD.n4412 VSS 0.140524f
C14698 DVDD.n4413 VSS 0.628154f
C14699 DVDD.n4415 VSS 0.066237f
C14700 DVDD.n4416 VSS 0.140524f
C14701 DVDD.n4417 VSS 0.157347f
C14702 DVDD.n4418 VSS 0.281047f
C14703 DVDD.n4419 VSS 0.281047f
C14704 DVDD.n4420 VSS 0.281047f
C14705 DVDD.n4421 VSS 0.281047f
C14706 DVDD.n4422 VSS 0.281047f
C14707 DVDD.n4423 VSS 0.281047f
C14708 DVDD.n4424 VSS 0.281047f
C14709 DVDD.n4425 VSS 0.281047f
C14710 DVDD.n4426 VSS 0.281047f
C14711 DVDD.n4427 VSS 0.281047f
C14712 DVDD.n4428 VSS 0.281047f
C14713 DVDD.n4429 VSS 0.281047f
C14714 DVDD.n4430 VSS 0.281047f
C14715 DVDD.n4431 VSS 0.281047f
C14716 DVDD.n4432 VSS 0.281047f
C14717 DVDD.n4433 VSS 0.1999f
C14718 DVDD.n4434 VSS 0.281047f
C14719 DVDD.n4435 VSS 0.281047f
C14720 DVDD.n4436 VSS 0.281047f
C14721 DVDD.n4437 VSS 0.281047f
C14722 DVDD.n4438 VSS 0.281047f
C14723 DVDD.n4439 VSS 0.281047f
C14724 DVDD.n4440 VSS 0.188025f
C14725 DVDD.n4441 VSS 0.188025f
C14726 DVDD.n4442 VSS 0.536365f
C14727 DVDD.n4443 VSS 0.233546f
C14728 DVDD.n4444 VSS 0.233546f
C14729 DVDD.n4445 VSS 0.233546f
C14730 DVDD.n4446 VSS 0.281047f
C14731 DVDD.n4447 VSS 0.281047f
C14732 DVDD.n4448 VSS 0.281047f
C14733 DVDD.n4449 VSS 0.281047f
C14734 DVDD.n4450 VSS 0.281047f
C14735 DVDD.n4451 VSS 0.281047f
C14736 DVDD.n4452 VSS 0.281047f
C14737 DVDD.n4453 VSS 0.281047f
C14738 DVDD.n4454 VSS 0.281047f
C14739 DVDD.n4455 VSS 0.281047f
C14740 DVDD.n4456 VSS 0.281047f
C14741 DVDD.n4457 VSS 0.281047f
C14742 DVDD.n4458 VSS 0.281047f
C14743 DVDD.n4459 VSS 0.281047f
C14744 DVDD.n4460 VSS 0.281047f
C14745 DVDD.n4461 VSS 0.281047f
C14746 DVDD.n4462 VSS 0.281047f
C14747 DVDD.n4463 VSS 0.281047f
C14748 DVDD.n4464 VSS 0.281047f
C14749 DVDD.n4465 VSS 0.281047f
C14750 DVDD.n4466 VSS 0.281047f
C14751 DVDD.n4467 VSS 0.281047f
C14752 DVDD.n4468 VSS 0.281047f
C14753 DVDD.n4469 VSS 0.281047f
C14754 DVDD.n4470 VSS 0.281047f
C14755 DVDD.n4471 VSS 0.281047f
C14756 DVDD.n4472 VSS 0.281047f
C14757 DVDD.n4473 VSS 0.281047f
C14758 DVDD.n4474 VSS 0.281047f
C14759 DVDD.n4475 VSS 0.281047f
C14760 DVDD.n4476 VSS 0.281047f
C14761 DVDD.n4477 VSS 0.281047f
C14762 DVDD.n4478 VSS 0.281047f
C14763 DVDD.n4479 VSS 0.281047f
C14764 DVDD.n4480 VSS 0.281047f
C14765 DVDD.n4481 VSS 0.281047f
C14766 DVDD.n4482 VSS 0.218702f
C14767 DVDD.n4483 VSS 0.281047f
C14768 DVDD.n4484 VSS 0.281047f
C14769 DVDD.n4485 VSS 0.281047f
C14770 DVDD.n4486 VSS 0.281047f
C14771 DVDD.n4487 VSS 0.281047f
C14772 DVDD.n4488 VSS 0.281047f
C14773 DVDD.n4489 VSS 0.281047f
C14774 DVDD.n4490 VSS 0.281047f
C14775 DVDD.n4491 VSS 0.281047f
C14776 DVDD.n4492 VSS 0.281047f
C14777 DVDD.n4493 VSS 0.281047f
C14778 DVDD.n4494 VSS 0.281047f
C14779 DVDD.n4495 VSS 0.281047f
C14780 DVDD.n4496 VSS 0.266203f
C14781 DVDD.n4497 VSS 0.281047f
C14782 DVDD.n4498 VSS 0.281047f
C14783 DVDD.n4499 VSS 0.140524f
C14784 DVDD.n4500 VSS 0.00998f
C14785 DVDD.n4501 VSS 0.00998f
C14786 DVDD.n4502 VSS 0.00998f
C14787 DVDD.n4503 VSS 0.00998f
C14788 DVDD.n4504 VSS 0.00998f
C14789 DVDD.n4505 VSS 0.00998f
C14790 DVDD.n4506 VSS 0.00998f
C14791 DVDD.n4507 VSS 0.00998f
C14792 DVDD.n4508 VSS 0.00998f
C14793 DVDD.n4509 VSS 0.011429f
C14794 DVDD.n4510 VSS 0.019961f
C14795 DVDD.n4511 VSS 0.011188f
C14796 DVDD.n4512 VSS 0.010222f
C14797 DVDD.n4513 VSS 0.019961f
C14798 DVDD.n4514 VSS 0.011429f
C14799 DVDD.n4515 VSS 0.019961f
C14800 DVDD.n4516 VSS 0.011429f
C14801 DVDD.n4517 VSS 0.019961f
C14802 DVDD.n4518 VSS 0.011429f
C14803 DVDD.n4519 VSS 0.019961f
C14804 DVDD.n4520 VSS 0.011429f
C14805 DVDD.n4521 VSS 0.019961f
C14806 DVDD.n4522 VSS 0.011429f
C14807 DVDD.n4523 VSS 0.019961f
C14808 DVDD.n4524 VSS 0.011429f
C14809 DVDD.n4525 VSS 0.019961f
C14810 DVDD.n4526 VSS 0.019961f
C14811 DVDD.n4527 VSS 0.011027f
C14812 DVDD.n4528 VSS 0.010383f
C14813 DVDD.n4529 VSS 0.019961f
C14814 DVDD.n4530 VSS 0.011429f
C14815 DVDD.n4531 VSS 0.019961f
C14816 DVDD.n4532 VSS 0.011429f
C14817 DVDD.n4533 VSS 0.019961f
C14818 DVDD.n4534 VSS 0.011429f
C14819 DVDD.n4535 VSS 0.019961f
C14820 DVDD.n4536 VSS 0.011429f
C14821 DVDD.n4537 VSS 0.019961f
C14822 DVDD.n4538 VSS 0.011429f
C14823 DVDD.n4539 VSS 0.019961f
C14824 DVDD.n4540 VSS 0.011429f
C14825 DVDD.n4541 VSS 0.019961f
C14826 DVDD.n4542 VSS 0.019961f
C14827 DVDD.n4543 VSS 0.010866f
C14828 DVDD.n4544 VSS 0.010544f
C14829 DVDD.n4545 VSS 0.019961f
C14830 DVDD.n4546 VSS 0.011429f
C14831 DVDD.n4547 VSS 0.019961f
C14832 DVDD.n4548 VSS 0.019961f
C14833 DVDD.n4549 VSS 0.019961f
C14834 DVDD.n4550 VSS 0.011429f
C14835 DVDD.n4551 VSS 0.061904f
C14836 DVDD.n4552 VSS 0.011429f
C14837 DVDD.n4553 VSS 0.019961f
C14838 DVDD.n4554 VSS 0.019961f
C14839 DVDD.n4555 VSS 0.014971f
C14840 DVDD.n4556 VSS 0.019961f
C14841 DVDD.n4557 VSS 0.015051f
C14842 DVDD.n4558 VSS 0.019961f
C14843 DVDD.n4559 VSS 0.019961f
C14844 DVDD.n4560 VSS 0.011429f
C14845 DVDD.n4561 VSS 0.00998f
C14846 DVDD.n4562 VSS 0.140524f
C14847 DVDD.n4563 VSS 0.00998f
C14848 DVDD.n4564 VSS 0.011429f
C14849 DVDD.n4565 VSS 0.019961f
C14850 DVDD.n4566 VSS 0.019961f
C14851 DVDD.n4567 VSS 0.015856f
C14852 DVDD.n4568 VSS 0.019961f
C14853 DVDD.n4569 VSS 0.012073f
C14854 DVDD.n4570 VSS -0.36209f
C14855 DVDD.n4571 VSS 0.011429f
C14856 DVDD.n4572 VSS 0.019961f
C14857 DVDD.n4573 VSS 0.011429f
C14858 DVDD.n4574 VSS 0.019961f
C14859 DVDD.n4575 VSS 0.011429f
C14860 DVDD.n4576 VSS 0.019961f
C14861 DVDD.n4577 VSS 0.011429f
C14862 DVDD.n4578 VSS 0.019961f
C14863 DVDD.n4579 VSS 0.011429f
C14864 DVDD.n4580 VSS 0.019961f
C14865 DVDD.n4581 VSS 0.019961f
C14866 DVDD.n4582 VSS 0.010624f
C14867 DVDD.n4583 VSS 0.010785f
C14868 DVDD.n4584 VSS 0.019961f
C14869 DVDD.n4585 VSS 0.011429f
C14870 DVDD.n4586 VSS 0.019961f
C14871 DVDD.n4587 VSS 0.011429f
C14872 DVDD.n4588 VSS 0.019961f
C14873 DVDD.n4589 VSS 0.011429f
C14874 DVDD.n4590 VSS 0.019961f
C14875 DVDD.n4591 VSS 0.011429f
C14876 DVDD.n4592 VSS 0.019961f
C14877 DVDD.n4593 VSS 0.011429f
C14878 DVDD.n4594 VSS 0.019961f
C14879 DVDD.n4595 VSS 0.011429f
C14880 DVDD.n4596 VSS 0.019961f
C14881 DVDD.n4597 VSS 0.019961f
C14882 DVDD.n4598 VSS 0.010463f
C14883 DVDD.n4599 VSS 0.010946f
C14884 DVDD.n4600 VSS 0.019961f
C14885 DVDD.n4601 VSS 0.011429f
C14886 DVDD.n4602 VSS 0.019961f
C14887 DVDD.n4603 VSS 0.011429f
C14888 DVDD.n4604 VSS 0.019961f
C14889 DVDD.n4605 VSS 0.011429f
C14890 DVDD.n4606 VSS 0.019961f
C14891 DVDD.n4607 VSS 0.011429f
C14892 DVDD.n4608 VSS 0.019961f
C14893 DVDD.n4609 VSS 0.011429f
C14894 DVDD.n4610 VSS 0.019961f
C14895 DVDD.n4611 VSS 0.011429f
C14896 DVDD.n4612 VSS 0.019961f
C14897 DVDD.n4613 VSS 0.019961f
C14898 DVDD.n4614 VSS 0.019961f
C14899 DVDD.n4615 VSS 0.011107f
C14900 DVDD.n4616 VSS 0.00998f
C14901 DVDD.n4617 VSS 0.140524f
C14902 DVDD.n4618 VSS 0.140524f
C14903 DVDD.n4619 VSS 0.281047f
C14904 DVDD.n4620 VSS 0.281047f
C14905 DVDD.n4621 VSS 0.155368f
C14906 DVDD.n4622 VSS 0.281047f
C14907 DVDD.n4623 VSS 0.281047f
C14908 DVDD.n4624 VSS 0.281047f
C14909 DVDD.n4625 VSS 0.281047f
C14910 DVDD.n4626 VSS 0.281047f
C14911 DVDD.n4627 VSS 0.281047f
C14912 DVDD.n4628 VSS 0.281047f
C14913 DVDD.n4629 VSS 0.281047f
C14914 DVDD.n4630 VSS 0.281047f
C14915 DVDD.n4631 VSS 0.281047f
C14916 DVDD.n4632 VSS 0.281047f
C14917 DVDD.n4633 VSS 0.281047f
C14918 DVDD.n4634 VSS 0.281047f
C14919 DVDD.n4635 VSS 0.233546f
C14920 DVDD.n4636 VSS 0.233546f
C14921 DVDD.n4637 VSS 0.536365f
C14922 DVDD.n4638 VSS 0.095991f
C14923 DVDD.n4639 VSS 0.188025f
C14924 DVDD.n4640 VSS 0.140524f
C14925 DVDD.n4641 VSS 0.281047f
C14926 DVDD.n4642 VSS 0.173181f
C14927 DVDD.n4643 VSS 0.281047f
C14928 DVDD.n4644 VSS 0.281047f
C14929 DVDD.n4645 VSS 0.140524f
C14930 DVDD.n4646 VSS 0.027215f
C14931 DVDD.n4647 VSS 0.023765f
C14932 DVDD.n4648 VSS 0.023765f
C14933 DVDD.n4649 VSS 0.023765f
C14934 DVDD.n4650 VSS 0.023765f
C14935 DVDD.n4651 VSS 0.023765f
C14936 DVDD.n4652 VSS 0.023765f
C14937 DVDD.n4653 VSS 0.023765f
C14938 DVDD.n4654 VSS 0.023765f
C14939 DVDD.n4655 VSS 0.023765f
C14940 DVDD.n4656 VSS 0.024532f
C14941 DVDD.n4657 VSS 0.070763f
C14942 DVDD.n4658 VSS 0.027215f
C14943 DVDD.n4659 VSS 0.070763f
C14944 DVDD.n4660 VSS 0.027215f
C14945 DVDD.n4661 VSS 0.070763f
C14946 DVDD.n4662 VSS 0.027215f
C14947 DVDD.n4663 VSS 0.070763f
C14948 DVDD.n4664 VSS 0.027215f
C14949 DVDD.n4665 VSS 0.070763f
C14950 DVDD.n4666 VSS 0.070763f
C14951 DVDD.n4667 VSS 0.025298f
C14952 DVDD.n4668 VSS 0.025681f
C14953 DVDD.n4669 VSS 0.070763f
C14954 DVDD.n4670 VSS 0.027215f
C14955 DVDD.n4671 VSS 0.070763f
C14956 DVDD.n4672 VSS 0.027215f
C14957 DVDD.n4673 VSS 0.070763f
C14958 DVDD.n4674 VSS 0.027215f
C14959 DVDD.n4675 VSS 0.070763f
C14960 DVDD.n4676 VSS 0.027215f
C14961 DVDD.n4677 VSS 0.058779f
C14962 DVDD.n4678 VSS 0.035382f
C14963 DVDD.n4679 VSS 0.027215f
C14964 DVDD.n4680 VSS 0.047366f
C14965 DVDD.n4681 VSS 0.027215f
C14966 DVDD.n4682 VSS 0.070763f
C14967 DVDD.n4683 VSS 0.070763f
C14968 DVDD.n4684 VSS 0.024915f
C14969 DVDD.n4685 VSS 0.026065f
C14970 DVDD.n4686 VSS 0.070763f
C14971 DVDD.n4687 VSS 0.027215f
C14972 DVDD.n4688 VSS 0.070763f
C14973 DVDD.n4689 VSS 0.027215f
C14974 DVDD.n4690 VSS 0.070763f
C14975 DVDD.n4691 VSS 0.027215f
C14976 DVDD.n4692 VSS 0.070763f
C14977 DVDD.n4693 VSS 0.027215f
C14978 DVDD.n4694 VSS 0.070763f
C14979 DVDD.n4695 VSS 0.027215f
C14980 DVDD.n4696 VSS 0.070763f
C14981 DVDD.n4697 VSS 0.070763f
C14982 DVDD.n4698 VSS 0.027215f
C14983 DVDD.n4699 VSS 0.023765f
C14984 DVDD.n4700 VSS 0.140524f
C14985 DVDD.n4701 VSS 0.026266f
C14986 DVDD.n4702 VSS 0.025004f
C14987 DVDD.n4703 VSS 0.070763f
C14988 DVDD.n4704 VSS 0.070763f
C14989 DVDD.n4705 VSS 0.070763f
C14990 DVDD.n4706 VSS 0.031546f
C14991 DVDD.n4707 VSS 0.023764f
C14992 DVDD.n4708 VSS 0.091044f
C14993 DVDD.n4709 VSS 0.130628f
C14994 DVDD.n4710 VSS 0.059376f
C14995 DVDD.n4711 VSS 0.02675f
C14996 DVDD.n4712 VSS 0.092033f
C14997 DVDD.n4713 VSS 0.130628f
C14998 DVDD.n4714 VSS 0.281047f
C14999 DVDD.n4715 VSS 0.281047f
C15000 DVDD.n4716 VSS 0.281047f
C15001 DVDD.n4717 VSS 0.188025f
C15002 DVDD.n4718 VSS 0.188025f
C15003 DVDD.n4719 VSS 0.095991f
C15004 DVDD.n4720 VSS 0.338444f
C15005 DVDD.n4721 VSS 0.233546f
C15006 DVDD.n4722 VSS 0.233546f
C15007 DVDD.n4723 VSS 0.233546f
C15008 DVDD.n4724 VSS 0.281047f
C15009 DVDD.n4725 VSS 0.281047f
C15010 DVDD.n4726 VSS 0.281047f
C15011 DVDD.n4727 VSS 0.281047f
C15012 DVDD.n4728 VSS 0.281047f
C15013 DVDD.n4729 VSS 0.281047f
C15014 DVDD.n4730 VSS 0.281047f
C15015 DVDD.n4731 VSS 0.281047f
C15016 DVDD.n4732 VSS 0.281047f
C15017 DVDD.n4733 VSS 0.281047f
C15018 DVDD.n4734 VSS 0.281047f
C15019 DVDD.n4735 VSS 0.281047f
C15020 DVDD.n4736 VSS 0.281047f
C15021 DVDD.n4737 VSS 0.281047f
C15022 DVDD.n4738 VSS 0.281047f
C15023 DVDD.n4739 VSS 0.281047f
C15024 DVDD.n4740 VSS 0.281047f
C15025 DVDD.n4741 VSS 0.281047f
C15026 DVDD.n4742 VSS 0.281047f
C15027 DVDD.n4743 VSS 0.155368f
C15028 DVDD.n4744 VSS 0.140524f
C15029 DVDD.n4745 VSS 0.027607f
C15030 DVDD.n4746 VSS 0.140524f
C15031 DVDD.n4747 VSS 0.266203f
C15032 DVDD.n4748 VSS 0.281047f
C15033 DVDD.n4749 VSS 0.281047f
C15034 DVDD.n4750 VSS 0.281047f
C15035 DVDD.n4751 VSS 0.281047f
C15036 DVDD.n4752 VSS 0.281047f
C15037 DVDD.n4753 VSS 0.281047f
C15038 DVDD.n4754 VSS 0.281047f
C15039 DVDD.n4755 VSS 0.281047f
C15040 DVDD.n4756 VSS 0.281047f
C15041 DVDD.n4757 VSS 0.281047f
C15042 DVDD.n4758 VSS 0.281047f
C15043 DVDD.n4759 VSS 0.281047f
C15044 DVDD.n4760 VSS 0.281047f
C15045 DVDD.n4761 VSS 0.281047f
C15046 DVDD.n4762 VSS 0.281047f
C15047 DVDD.n4763 VSS 0.281047f
C15048 DVDD.n4764 VSS 0.281047f
C15049 DVDD.n4765 VSS 0.281047f
C15050 DVDD.n4766 VSS 0.281047f
C15051 DVDD.n4767 VSS 0.338444f
C15052 DVDD.n4768 VSS 0.180108f
C15053 DVDD.n4769 VSS 0.281047f
C15054 DVDD.n4770 VSS 0.281047f
C15055 DVDD.n4771 VSS 0.218702f
C15056 DVDD.n4772 VSS 0.101929f
C15057 DVDD.n4773 VSS 0.140524f
C15058 DVDD.n4774 VSS 0.027607f
C15059 DVDD.n4775 VSS 0.10094f
C15060 DVDD.n4776 VSS 0.281047f
C15061 DVDD.n4777 VSS 0.281047f
C15062 DVDD.n4778 VSS 0.281047f
C15063 DVDD.n4779 VSS 0.281047f
C15064 DVDD.n4780 VSS 0.281047f
C15065 DVDD.n4781 VSS 0.281047f
C15066 DVDD.n4782 VSS 0.281047f
C15067 DVDD.n4783 VSS 0.281047f
C15068 DVDD.n4784 VSS 0.281047f
C15069 DVDD.n4785 VSS 0.281047f
C15070 DVDD.n4786 VSS 0.281047f
C15071 DVDD.n4787 VSS 0.281047f
C15072 DVDD.n4788 VSS 0.281047f
C15073 DVDD.n4789 VSS 0.281047f
C15074 DVDD.n4790 VSS 0.281047f
C15075 DVDD.n4791 VSS 0.281047f
C15076 DVDD.n4792 VSS 0.281047f
C15077 DVDD.n4793 VSS 0.281047f
C15078 DVDD.n4794 VSS 0.281047f
C15079 DVDD.n4795 VSS 0.281047f
C15080 DVDD.n4796 VSS 0.281047f
C15081 DVDD.n4797 VSS 0.281047f
C15082 DVDD.n4798 VSS 0.281047f
C15083 DVDD.n4799 VSS 0.281047f
C15084 DVDD.n4800 VSS 0.281047f
C15085 DVDD.n4801 VSS 0.281047f
C15086 DVDD.n4802 VSS 0.202869f
C15087 DVDD.n4803 VSS 0.241463f
C15088 DVDD.n4804 VSS 0.338444f
C15089 DVDD.n4805 VSS 0.241463f
C15090 DVDD.n4806 VSS 0.281047f
C15091 DVDD.n4807 VSS 0.281047f
C15092 DVDD.n4808 VSS 0.281047f
C15093 DVDD.n4809 VSS 0.281047f
C15094 DVDD.n4810 VSS 0.281047f
C15095 DVDD.n4811 VSS 0.281047f
C15096 DVDD.n4812 VSS 0.281047f
C15097 DVDD.n4813 VSS 0.281047f
C15098 DVDD.n4814 VSS 0.281047f
C15099 DVDD.n4815 VSS 0.281047f
C15100 DVDD.n4816 VSS 0.281047f
C15101 DVDD.n4817 VSS 0.281047f
C15102 DVDD.n4818 VSS 0.281047f
C15103 DVDD.n4819 VSS 0.281047f
C15104 DVDD.n4820 VSS 0.281047f
C15105 DVDD.n4821 VSS 0.281047f
C15106 DVDD.n4822 VSS 0.281047f
C15107 DVDD.n4823 VSS 0.281047f
C15108 DVDD.n4824 VSS 0.281047f
C15109 DVDD.n4825 VSS 0.281047f
C15110 DVDD.n4826 VSS 0.281047f
C15111 DVDD.n4827 VSS 0.281047f
C15112 DVDD.n4828 VSS 0.281047f
C15113 DVDD.n4829 VSS 0.281047f
C15114 DVDD.n4830 VSS 0.281047f
C15115 DVDD.n4831 VSS 0.281047f
C15116 DVDD.n4832 VSS 0.281047f
C15117 DVDD.n4833 VSS 0.281047f
C15118 DVDD.n4834 VSS 0.281047f
C15119 DVDD.n4835 VSS 0.172191f
C15120 DVDD.n4836 VSS 0.281047f
C15121 DVDD.n4837 VSS 0.281047f
C15122 DVDD.n4838 VSS 0.172191f
C15123 DVDD.n4839 VSS 0.281047f
C15124 DVDD.n4840 VSS 0.281047f
C15125 DVDD.n4841 VSS 0.281047f
C15126 DVDD.n4842 VSS 0.281047f
C15127 DVDD.n4843 VSS 0.281047f
C15128 DVDD.n4844 VSS 0.281047f
C15129 DVDD.n4845 VSS 0.281047f
C15130 DVDD.n4846 VSS 0.281047f
C15131 DVDD.n4847 VSS 0.281047f
C15132 DVDD.n4848 VSS 0.281047f
C15133 DVDD.n4849 VSS 0.281047f
C15134 DVDD.n4850 VSS 0.281047f
C15135 DVDD.n4851 VSS 0.281047f
C15136 DVDD.n4852 VSS 0.280058f
C15137 DVDD.n4853 VSS 0.281047f
C15138 DVDD.n4854 VSS 0.281047f
C15139 DVDD.n4855 VSS 0.281047f
C15140 DVDD.n4856 VSS 0.281047f
C15141 DVDD.n4857 VSS 0.281047f
C15142 DVDD.n4858 VSS 0.281047f
C15143 DVDD.n4859 VSS 0.281047f
C15144 DVDD.n4860 VSS 0.281047f
C15145 DVDD.n4861 VSS 0.281047f
C15146 DVDD.n4862 VSS 0.281047f
C15147 DVDD.n4863 VSS 0.281047f
C15148 DVDD.n4864 VSS 0.281047f
C15149 DVDD.n4865 VSS 0.281047f
C15150 DVDD.n4866 VSS 0.281047f
C15151 DVDD.n4867 VSS 0.281047f
C15152 DVDD.n4868 VSS 0.281047f
C15153 DVDD.n4869 VSS 0.281047f
C15154 DVDD.n4870 VSS 0.281047f
C15155 DVDD.n4871 VSS 0.281047f
C15156 DVDD.n4872 VSS 0.241463f
C15157 DVDD.n4873 VSS 0.536365f
C15158 DVDD.n4874 VSS 0.180108f
C15159 DVDD.n4875 VSS 0.281047f
C15160 DVDD.n4876 VSS 0.218702f
C15161 DVDD.n4877 VSS 0.140524f
C15162 DVDD.n4878 VSS 0.00998f
C15163 DVDD.n4879 VSS 0.10094f
C15164 DVDD.n4880 VSS 0.47402f
C15165 DVDD.n4881 VSS 0.47402f
C15166 DVDD.n4882 VSS 0.101929f
C15167 DVDD.n4883 VSS 0.180108f
C15168 DVDD.n4884 VSS 0.180108f
C15169 DVDD.n4885 VSS 0.536365f
C15170 DVDD.n4886 VSS 0.241463f
C15171 DVDD.n4887 VSS 0.241463f
C15172 DVDD.n4888 VSS 0.202869f
C15173 DVDD.n4889 VSS 0.281047f
C15174 DVDD.n4890 VSS 0.281047f
C15175 DVDD.n4891 VSS 0.281047f
C15176 DVDD.n4892 VSS 0.281047f
C15177 DVDD.n4893 VSS 0.281047f
C15178 DVDD.n4894 VSS 0.281047f
C15179 DVDD.n4895 VSS 0.281047f
C15180 DVDD.n4896 VSS 0.281047f
C15181 DVDD.n4897 VSS 0.281047f
C15182 DVDD.n4898 VSS 0.281047f
C15183 DVDD.n4899 VSS 0.281047f
C15184 DVDD.n4900 VSS 0.281047f
C15185 DVDD.n4901 VSS 0.281047f
C15186 DVDD.n4902 VSS 0.281047f
C15187 DVDD.n4903 VSS 0.281047f
C15188 DVDD.n4904 VSS 0.281047f
C15189 DVDD.n4905 VSS 0.281047f
C15190 DVDD.n4906 VSS 0.281047f
C15191 DVDD.n4907 VSS 0.281047f
C15192 DVDD.n4908 VSS 0.281047f
C15193 DVDD.n4909 VSS 0.281047f
C15194 DVDD.n4910 VSS 0.281047f
C15195 DVDD.n4911 VSS 0.281047f
C15196 DVDD.n4912 VSS 0.281047f
C15197 DVDD.n4913 VSS 0.281047f
C15198 DVDD.n4914 VSS 0.281047f
C15199 DVDD.n4915 VSS 0.281047f
C15200 DVDD.n4916 VSS 0.281047f
C15201 DVDD.n4917 VSS 0.281047f
C15202 DVDD.n4918 VSS 0.281047f
C15203 DVDD.n4919 VSS 0.281047f
C15204 DVDD.n4920 VSS 0.281047f
C15205 DVDD.n4921 VSS 0.281047f
C15206 DVDD.n4922 VSS 0.281047f
C15207 DVDD.n4923 VSS 0.281047f
C15208 DVDD.n4924 VSS 0.281047f
C15209 DVDD.n4925 VSS 0.281047f
C15210 DVDD.n4926 VSS 0.281047f
C15211 DVDD.n4927 VSS 0.281047f
C15212 DVDD.n4928 VSS 0.281047f
C15213 DVDD.n4929 VSS 0.281047f
C15214 DVDD.n4930 VSS 0.281047f
C15215 DVDD.n4931 VSS 0.281047f
C15216 DVDD.n4932 VSS 0.281047f
C15217 DVDD.n4933 VSS 0.281047f
C15218 DVDD.n4934 VSS 0.281047f
C15219 DVDD.n4935 VSS 0.281047f
C15220 DVDD.n4936 VSS 0.281047f
C15221 DVDD.n4937 VSS 0.280058f
C15222 DVDD.n4938 VSS 0.281047f
C15223 DVDD.n4939 VSS 0.281047f
C15224 DVDD.n4940 VSS 0.140524f
C15225 DVDD.n4941 VSS 0.00998f
C15226 DVDD.n4942 VSS 0.00998f
C15227 DVDD.n4943 VSS 0.00998f
C15228 DVDD.n4944 VSS 0.00998f
C15229 DVDD.n4945 VSS 0.00998f
C15230 DVDD.n4946 VSS 0.00998f
C15231 DVDD.n4947 VSS 0.00998f
C15232 DVDD.n4948 VSS 0.00998f
C15233 DVDD.n4949 VSS 0.00998f
C15234 DVDD.n4950 VSS 0.00998f
C15235 DVDD.n4951 VSS 0.011429f
C15236 DVDD.n4952 VSS 0.011429f
C15237 DVDD.n4953 VSS 0.019961f
C15238 DVDD.n4954 VSS 0.019961f
C15239 DVDD.n4955 VSS 0.011188f
C15240 DVDD.n4956 VSS 0.010222f
C15241 DVDD.n4957 VSS 0.019961f
C15242 DVDD.n4958 VSS 0.011429f
C15243 DVDD.n4959 VSS 0.019961f
C15244 DVDD.n4960 VSS 0.011429f
C15245 DVDD.n4961 VSS 0.019961f
C15246 DVDD.n4962 VSS 0.011429f
C15247 DVDD.n4963 VSS 0.019961f
C15248 DVDD.n4964 VSS 0.011429f
C15249 DVDD.n4965 VSS 0.019961f
C15250 DVDD.n4966 VSS 0.011429f
C15251 DVDD.n4967 VSS 0.019961f
C15252 DVDD.n4968 VSS 0.011429f
C15253 DVDD.n4969 VSS 0.019961f
C15254 DVDD.n4970 VSS 0.019961f
C15255 DVDD.n4971 VSS 0.011027f
C15256 DVDD.n4972 VSS 0.010383f
C15257 DVDD.n4973 VSS 0.019961f
C15258 DVDD.n4974 VSS 0.011429f
C15259 DVDD.n4975 VSS 0.019961f
C15260 DVDD.n4976 VSS 0.011429f
C15261 DVDD.n4977 VSS 0.019961f
C15262 DVDD.n4978 VSS 0.011429f
C15263 DVDD.n4979 VSS 0.019961f
C15264 DVDD.n4980 VSS 0.011429f
C15265 DVDD.n4981 VSS 0.019961f
C15266 DVDD.n4982 VSS 0.011429f
C15267 DVDD.n4983 VSS 0.019961f
C15268 DVDD.n4984 VSS 0.011429f
C15269 DVDD.n4985 VSS 0.019961f
C15270 DVDD.n4986 VSS 0.019961f
C15271 DVDD.n4987 VSS 0.010866f
C15272 DVDD.n4988 VSS 0.010544f
C15273 DVDD.n4989 VSS 0.019961f
C15274 DVDD.n4990 VSS 0.011429f
C15275 DVDD.n4991 VSS 0.019961f
C15276 DVDD.n4992 VSS 0.019961f
C15277 DVDD.n4993 VSS 0.019961f
C15278 DVDD.n4994 VSS 0.011429f
C15279 DVDD.n4995 VSS 0.061904f
C15280 DVDD.n4996 VSS 0.011429f
C15281 DVDD.n4997 VSS 0.019961f
C15282 DVDD.n4998 VSS 0.019961f
C15283 DVDD.n4999 VSS 0.014971f
C15284 DVDD.n5000 VSS 0.019961f
C15285 DVDD.n5001 VSS 0.015051f
C15286 DVDD.n5002 VSS 0.019961f
C15287 DVDD.n5003 VSS 0.019961f
C15288 DVDD.n5004 VSS 0.011429f
C15289 DVDD.n5005 VSS 0.00998f
C15290 DVDD.n5006 VSS 0.140524f
C15291 DVDD.n5007 VSS 0.00998f
C15292 DVDD.n5008 VSS 0.015856f
C15293 DVDD.n5009 VSS 0.019961f
C15294 DVDD.n5010 VSS -0.294669f
C15295 DVDD.n5011 VSS -0.36209f
C15296 DVDD.n5012 VSS 0.012073f
C15297 DVDD.n5013 VSS 0.00998f
C15298 DVDD.n5014 VSS 0.140524f
C15299 DVDD.n5015 VSS 0.00998f
C15300 DVDD.n5016 VSS 0.018834f
C15301 DVDD.n5017 VSS 0.019961f
C15302 DVDD.n5018 VSS 0.019961f
C15303 DVDD.n5019 VSS 0.019961f
C15304 DVDD.n5020 VSS 0.01312f
C15305 DVDD.n5021 VSS 0.00998f
C15306 DVDD.n5022 VSS 0.140524f
C15307 DVDD.n5023 VSS 0.141513f
C15308 DVDD.n5024 VSS 0.281047f
C15309 DVDD.n5025 VSS 0.281047f
C15310 DVDD.n5026 VSS 0.281047f
C15311 DVDD.n5027 VSS 0.281047f
C15312 DVDD.n5028 VSS 0.281047f
C15313 DVDD.n5029 VSS 0.280058f
C15314 DVDD.n5030 VSS 0.281047f
C15315 DVDD.n5031 VSS 0.281047f
C15316 DVDD.n5032 VSS 0.281047f
C15317 DVDD.n5033 VSS 0.281047f
C15318 DVDD.n5034 VSS 0.281047f
C15319 DVDD.n5035 VSS 0.281047f
C15320 DVDD.n5036 VSS 0.281047f
C15321 DVDD.n5037 VSS 0.281047f
C15322 DVDD.n5038 VSS 0.281047f
C15323 DVDD.n5039 VSS 0.281047f
C15324 DVDD.n5040 VSS 0.281047f
C15325 DVDD.n5041 VSS 0.281047f
C15326 DVDD.n5042 VSS 0.281047f
C15327 DVDD.n5043 VSS 0.281047f
C15328 DVDD.n5044 VSS 0.281047f
C15329 DVDD.n5045 VSS 0.281047f
C15330 DVDD.n5046 VSS 0.281047f
C15331 DVDD.n5047 VSS 0.172191f
C15332 DVDD.n5048 VSS 0.172191f
C15333 DVDD.n5049 VSS 0.172191f
C15334 DVDD.n5050 VSS 0.338444f
C15335 DVDD.n5051 VSS 0.24938f
C15336 DVDD.n5052 VSS 0.281047f
C15337 DVDD.n5053 VSS 0.281047f
C15338 DVDD.n5054 VSS 0.281047f
C15339 DVDD.n5055 VSS 0.281047f
C15340 DVDD.n5056 VSS 0.281047f
C15341 DVDD.n5057 VSS 0.281047f
C15342 DVDD.n5058 VSS 0.281047f
C15343 DVDD.n5059 VSS 0.281047f
C15344 DVDD.n5060 VSS 0.281047f
C15345 DVDD.n5061 VSS 0.281047f
C15346 DVDD.n5062 VSS 0.281047f
C15347 DVDD.n5063 VSS 0.281047f
C15348 DVDD.n5064 VSS 0.281047f
C15349 DVDD.n5065 VSS 0.281047f
C15350 DVDD.n5066 VSS 0.281047f
C15351 DVDD.n5067 VSS 0.281047f
C15352 DVDD.n5068 VSS 0.281047f
C15353 DVDD.n5069 VSS 0.281047f
C15354 DVDD.n5070 VSS 0.268182f
C15355 DVDD.n5071 VSS 0.281047f
C15356 DVDD.n5072 VSS 0.281047f
C15357 DVDD.n5073 VSS 0.281047f
C15358 DVDD.n5074 VSS 0.281047f
C15359 DVDD.n5075 VSS 0.281047f
C15360 DVDD.n5076 VSS 0.281047f
C15361 DVDD.n5077 VSS 0.281047f
C15362 DVDD.n5078 VSS 0.281047f
C15363 DVDD.n5079 VSS 0.281047f
C15364 DVDD.n5080 VSS 0.281047f
C15365 DVDD.n5081 VSS 0.281047f
C15366 DVDD.n5082 VSS 0.281047f
C15367 DVDD.n5083 VSS 0.281047f
C15368 DVDD.n5084 VSS 0.216723f
C15369 DVDD.n5085 VSS 0.281047f
C15370 DVDD.n5086 VSS 0.24938f
C15371 DVDD.n5087 VSS 0.140524f
C15372 DVDD.n5088 VSS 0.00998f
C15373 DVDD.n5089 VSS 0.00586f
C15374 DVDD.n5090 VSS 0.019961f
C15375 DVDD.n5091 VSS 0.011429f
C15376 DVDD.n5092 VSS 0.019961f
C15377 DVDD.n5093 VSS 0.063742f
C15378 DVDD.n5094 VSS 0.011429f
C15379 DVDD.n5095 VSS 0.017326f
C15380 DVDD.n5096 VSS 0.108856f
C15381 DVDD.n5097 VSS 0.00998f
C15382 DVDD.n5098 VSS 0.01312f
C15383 DVDD.n5099 VSS 0.019961f
C15384 DVDD.n5100 VSS 0.019961f
C15385 DVDD.n5101 VSS 0.019961f
C15386 DVDD.n5102 VSS -0.294669f
C15387 DVDD.n5103 VSS 0.019961f
C15388 DVDD.n5104 VSS 0.00998f
C15389 DVDD.n5105 VSS 0.061904f
C15390 DVDD.n5106 VSS 0.140524f
C15391 DVDD.n5107 VSS 0.281047f
C15392 DVDD.n5108 VSS 0.24938f
C15393 DVDD.n5109 VSS 0.24938f
C15394 DVDD.n5110 VSS 0.281047f
C15395 DVDD.n5111 VSS 0.281047f
C15396 DVDD.n5112 VSS 0.281047f
C15397 DVDD.n5113 VSS 0.281047f
C15398 DVDD.n5114 VSS 0.281047f
C15399 DVDD.n5115 VSS 0.281047f
C15400 DVDD.n5116 VSS 0.281047f
C15401 DVDD.n5117 VSS 0.281047f
C15402 DVDD.n5118 VSS 0.281047f
C15403 DVDD.n5119 VSS 0.281047f
C15404 DVDD.n5120 VSS 0.281047f
C15405 DVDD.n5121 VSS 0.281047f
C15406 DVDD.n5122 VSS 0.281047f
C15407 DVDD.n5123 VSS 0.281047f
C15408 DVDD.n5124 VSS 0.281047f
C15409 DVDD.n5125 VSS 0.281047f
C15410 DVDD.n5126 VSS 0.281047f
C15411 DVDD.n5127 VSS 0.281047f
C15412 DVDD.n5128 VSS 0.281047f
C15413 DVDD.n5129 VSS 0.281047f
C15414 DVDD.n5130 VSS 0.281047f
C15415 DVDD.n5131 VSS 0.281047f
C15416 DVDD.n5132 VSS 0.281047f
C15417 DVDD.n5133 VSS 0.281047f
C15418 DVDD.n5134 VSS 0.281047f
C15419 DVDD.n5135 VSS 0.216723f
C15420 DVDD.n5136 VSS 0.140524f
C15421 DVDD.n5137 VSS 0.025252f
C15422 DVDD.n5138 VSS 0.005232f
C15423 DVDD.n5139 VSS 0.017881f
C15424 DVDD.n5140 VSS 0.011429f
C15425 DVDD.n5141 VSS 0.00998f
C15426 DVDD.n5142 VSS 0.011429f
C15427 DVDD.n5143 VSS 0.019961f
C15428 DVDD.n5144 VSS 0.019961f
C15429 DVDD.n5145 VSS 0.014971f
C15430 DVDD.n5146 VSS 0.019961f
C15431 DVDD.n5147 VSS 0.015051f
C15432 DVDD.n5148 VSS 0.019961f
C15433 DVDD.n5149 VSS 0.019961f
C15434 DVDD.n5150 VSS 0.019961f
C15435 DVDD.n5151 VSS 0.011429f
C15436 DVDD.n5152 VSS 0.019961f
C15437 DVDD.n5153 VSS 0.019961f
C15438 DVDD.n5154 VSS 0.010544f
C15439 DVDD.n5155 VSS 0.010866f
C15440 DVDD.n5156 VSS 0.019961f
C15441 DVDD.n5157 VSS 0.011429f
C15442 DVDD.n5158 VSS 0.019961f
C15443 DVDD.n5159 VSS 0.011429f
C15444 DVDD.n5160 VSS 0.019961f
C15445 DVDD.n5161 VSS 0.011429f
C15446 DVDD.n5162 VSS 0.019961f
C15447 DVDD.n5163 VSS 0.011429f
C15448 DVDD.n5164 VSS 0.019961f
C15449 DVDD.n5165 VSS 0.011429f
C15450 DVDD.n5166 VSS 0.019961f
C15451 DVDD.n5167 VSS 0.011429f
C15452 DVDD.n5168 VSS 0.019961f
C15453 DVDD.n5169 VSS 0.019961f
C15454 DVDD.n5170 VSS 0.010383f
C15455 DVDD.n5171 VSS 0.011027f
C15456 DVDD.n5172 VSS 0.019961f
C15457 DVDD.n5173 VSS 0.011429f
C15458 DVDD.n5174 VSS 0.019961f
C15459 DVDD.n5175 VSS 0.011429f
C15460 DVDD.n5176 VSS 0.019961f
C15461 DVDD.n5177 VSS 0.011429f
C15462 DVDD.n5178 VSS 0.019961f
C15463 DVDD.n5179 VSS 0.011429f
C15464 DVDD.n5180 VSS 0.019961f
C15465 DVDD.n5181 VSS 0.011429f
C15466 DVDD.n5182 VSS 0.019961f
C15467 DVDD.n5183 VSS 0.011429f
C15468 DVDD.n5184 VSS 0.019961f
C15469 DVDD.n5185 VSS 0.019961f
C15470 DVDD.n5186 VSS 0.010222f
C15471 DVDD.n5187 VSS 0.011188f
C15472 DVDD.n5188 VSS 0.019961f
C15473 DVDD.n5189 VSS 0.011429f
C15474 DVDD.n5190 VSS 0.019961f
C15475 DVDD.n5191 VSS 0.011429f
C15476 DVDD.n5192 VSS 0.019961f
C15477 DVDD.n5193 VSS 0.019961f
C15478 DVDD.n5194 VSS 0.015856f
C15479 DVDD.n5195 VSS 0.019961f
C15480 DVDD.n5196 VSS 0.012073f
C15481 DVDD.n5197 VSS -0.36209f
C15482 DVDD.n5198 VSS 0.011429f
C15483 DVDD.n5199 VSS 0.019961f
C15484 DVDD.n5200 VSS 0.011429f
C15485 DVDD.n5201 VSS 0.019961f
C15486 DVDD.n5202 VSS 0.011429f
C15487 DVDD.n5203 VSS 0.019961f
C15488 DVDD.n5204 VSS 0.011429f
C15489 DVDD.n5205 VSS 0.019961f
C15490 DVDD.n5206 VSS 0.011429f
C15491 DVDD.n5207 VSS 0.019961f
C15492 DVDD.n5208 VSS 0.019961f
C15493 DVDD.n5209 VSS 0.010624f
C15494 DVDD.n5210 VSS 0.010785f
C15495 DVDD.n5211 VSS 0.019961f
C15496 DVDD.n5212 VSS 0.011429f
C15497 DVDD.n5213 VSS 0.019961f
C15498 DVDD.n5214 VSS 0.011429f
C15499 DVDD.n5215 VSS 0.019961f
C15500 DVDD.n5216 VSS 0.011429f
C15501 DVDD.n5217 VSS 0.019961f
C15502 DVDD.n5218 VSS 0.011429f
C15503 DVDD.n5219 VSS 0.019961f
C15504 DVDD.n5220 VSS 0.011429f
C15505 DVDD.n5221 VSS 0.019961f
C15506 DVDD.n5222 VSS 0.011429f
C15507 DVDD.n5223 VSS 0.019961f
C15508 DVDD.n5224 VSS 0.019961f
C15509 DVDD.n5225 VSS 0.010463f
C15510 DVDD.n5226 VSS 0.010946f
C15511 DVDD.n5227 VSS 0.019961f
C15512 DVDD.n5228 VSS 0.011429f
C15513 DVDD.n5229 VSS 0.019961f
C15514 DVDD.n5230 VSS 0.011429f
C15515 DVDD.n5231 VSS 0.019961f
C15516 DVDD.n5232 VSS 0.011429f
C15517 DVDD.n5233 VSS 0.019961f
C15518 DVDD.n5234 VSS 0.011429f
C15519 DVDD.n5235 VSS 0.019961f
C15520 DVDD.n5236 VSS 0.011429f
C15521 DVDD.n5237 VSS 0.019961f
C15522 DVDD.n5238 VSS 0.011429f
C15523 DVDD.n5239 VSS 0.019961f
C15524 DVDD.n5240 VSS 0.019961f
C15525 DVDD.n5241 VSS 0.019961f
C15526 DVDD.n5242 VSS 0.011107f
C15527 DVDD.n5243 VSS 0.00998f
C15528 DVDD.n5244 VSS 0.140524f
C15529 DVDD.n5245 VSS 0.140524f
C15530 DVDD.n5246 VSS 0.24938f
C15531 DVDD.n5247 VSS 0.536365f
C15532 DVDD.n5248 VSS 0.536365f
C15533 DVDD.n5249 VSS 0.172191f
C15534 DVDD.n5250 VSS 0.172191f
C15535 DVDD.n5251 VSS 0.536365f
C15536 DVDD.n5252 VSS 0.24938f
C15537 DVDD.n5253 VSS 0.281047f
C15538 DVDD.n5254 VSS 0.281047f
C15539 DVDD.n5255 VSS 0.281047f
C15540 DVDD.n5256 VSS 0.281047f
C15541 DVDD.n5257 VSS 0.281047f
C15542 DVDD.n5258 VSS 0.281047f
C15543 DVDD.n5259 VSS 0.281047f
C15544 DVDD.n5260 VSS 0.281047f
C15545 DVDD.n5261 VSS 0.281047f
C15546 DVDD.n5262 VSS 0.281047f
C15547 DVDD.n5263 VSS 0.281047f
C15548 DVDD.n5264 VSS 0.281047f
C15549 DVDD.n5265 VSS 0.281047f
C15550 DVDD.n5266 VSS 0.281047f
C15551 DVDD.n5267 VSS 0.281047f
C15552 DVDD.n5268 VSS 0.281047f
C15553 DVDD.n5269 VSS 0.281047f
C15554 DVDD.n5270 VSS 0.281047f
C15555 DVDD.n5271 VSS 0.281047f
C15556 DVDD.n5272 VSS 0.281047f
C15557 DVDD.n5273 VSS 0.281047f
C15558 DVDD.n5274 VSS 0.281047f
C15559 DVDD.n5275 VSS 0.281047f
C15560 DVDD.n5276 VSS 0.281047f
C15561 DVDD.n5277 VSS 0.281047f
C15562 DVDD.n5278 VSS 0.281047f
C15563 DVDD.n5279 VSS 0.281047f
C15564 DVDD.n5280 VSS 0.281047f
C15565 DVDD.n5281 VSS 0.281047f
C15566 DVDD.n5282 VSS 0.281047f
C15567 DVDD.n5283 VSS 0.164274f
C15568 DVDD.n5284 VSS 0.164274f
C15569 DVDD.n5285 VSS 0.281047f
C15570 DVDD.n5286 VSS 0.281047f
C15571 DVDD.n5287 VSS 0.281047f
C15572 DVDD.n5288 VSS 0.281047f
C15573 DVDD.n5289 VSS 0.281047f
C15574 DVDD.n5290 VSS 0.281047f
C15575 DVDD.n5291 VSS 0.281047f
C15576 DVDD.n5292 VSS 0.281047f
C15577 DVDD.n5293 VSS 0.281047f
C15578 DVDD.n5294 VSS 0.281047f
C15579 DVDD.n5295 VSS 0.281047f
C15580 DVDD.n5296 VSS 0.281047f
C15581 DVDD.n5297 VSS 0.281047f
C15582 DVDD.n5298 VSS 0.281047f
C15583 DVDD.n5299 VSS 0.281047f
C15584 DVDD.n5300 VSS 0.281047f
C15585 DVDD.n5301 VSS 0.268182f
C15586 DVDD.n5302 VSS 0.281047f
C15587 DVDD.n5303 VSS 0.281047f
C15588 DVDD.n5304 VSS 0.281047f
C15589 DVDD.n5305 VSS 0.281047f
C15590 DVDD.n5306 VSS 0.281047f
C15591 DVDD.n5307 VSS 0.281047f
C15592 DVDD.n5308 VSS 0.281047f
C15593 DVDD.n5309 VSS 0.281047f
C15594 DVDD.n5310 VSS 0.281047f
C15595 DVDD.n5311 VSS 0.281047f
C15596 DVDD.n5312 VSS 0.281047f
C15597 DVDD.n5313 VSS 0.281047f
C15598 DVDD.n5314 VSS 0.281047f
C15599 DVDD.n5315 VSS 0.281047f
C15600 DVDD.n5316 VSS 0.281047f
C15601 DVDD.n5317 VSS 0.216723f
C15602 DVDD.n5318 VSS 0.140524f
C15603 DVDD.n5319 VSS 0.00998f
C15604 DVDD.n5320 VSS 0.108856f
C15605 DVDD.n5321 VSS 0.460165f
C15606 DVDD.n5322 VSS 0.262245f
C15607 DVDD.n5323 VSS 0.172191f
C15608 DVDD.n5324 VSS 0.172191f
C15609 DVDD.n5325 VSS 0.281047f
C15610 DVDD.n5326 VSS 0.281047f
C15611 DVDD.n5327 VSS 0.281047f
C15612 DVDD.n5328 VSS 0.281047f
C15613 DVDD.n5329 VSS 0.281047f
C15614 DVDD.n5330 VSS 0.281047f
C15615 DVDD.n5331 VSS 0.281047f
C15616 DVDD.n5332 VSS 0.281047f
C15617 DVDD.n5333 VSS 0.281047f
C15618 DVDD.n5334 VSS 0.281047f
C15619 DVDD.n5335 VSS 0.281047f
C15620 DVDD.n5336 VSS 0.281047f
C15621 DVDD.n5337 VSS 0.281047f
C15622 DVDD.n5338 VSS 0.281047f
C15623 DVDD.n5339 VSS 0.280058f
C15624 DVDD.n5340 VSS 0.140524f
C15625 DVDD.n5341 VSS 0.025252f
C15626 DVDD.n5342 VSS 0.140524f
C15627 DVDD.n5343 VSS 0.141513f
C15628 DVDD.n5344 VSS 0.281047f
C15629 DVDD.n5345 VSS 0.281047f
C15630 DVDD.n5346 VSS 0.281047f
C15631 DVDD.n5347 VSS 0.281047f
C15632 DVDD.n5348 VSS 0.281047f
C15633 DVDD.n5349 VSS 0.281047f
C15634 DVDD.n5350 VSS 0.281047f
C15635 DVDD.n5351 VSS 0.281047f
C15636 DVDD.n5352 VSS 0.281047f
C15637 DVDD.n5353 VSS 0.281047f
C15638 DVDD.n5354 VSS 0.281047f
C15639 DVDD.n5355 VSS 0.281047f
C15640 DVDD.n5356 VSS 0.281047f
C15641 DVDD.n5357 VSS 0.281047f
C15642 DVDD.n5358 VSS 0.281047f
C15643 DVDD.n5359 VSS 0.241463f
C15644 DVDD.n5360 VSS 0.202869f
C15645 DVDD.n5361 VSS 0.10094f
C15646 DVDD.n5362 VSS 0.025252f
C15647 DVDD.n5363 VSS 0.140524f
C15648 DVDD.n5364 VSS 0.218702f
C15649 DVDD.n5365 VSS 0.281047f
C15650 DVDD.n5366 VSS 0.281047f
C15651 DVDD.n5367 VSS 0.281047f
C15652 DVDD.n5368 VSS 0.281047f
C15653 DVDD.n5369 VSS 0.281047f
C15654 DVDD.n5370 VSS 0.281047f
C15655 DVDD.n5371 VSS 0.281047f
C15656 DVDD.n5372 VSS 0.281047f
C15657 DVDD.n5373 VSS 0.281047f
C15658 DVDD.n5374 VSS 0.281047f
C15659 DVDD.n5375 VSS 0.281047f
C15660 DVDD.n5376 VSS 0.281047f
C15661 DVDD.n5377 VSS 0.281047f
C15662 DVDD.n5378 VSS 0.281047f
C15663 DVDD.n5379 VSS 0.281047f
C15664 DVDD.n5380 VSS 0.266203f
C15665 DVDD.n5381 VSS 0.140524f
C15666 DVDD.n5382 VSS 0.025252f
C15667 DVDD.n5383 VSS 0.140524f
C15668 DVDD.n5384 VSS 0.155368f
C15669 DVDD.n5385 VSS 0.281047f
C15670 DVDD.n5386 VSS 0.281047f
C15671 DVDD.n5387 VSS 0.281047f
C15672 DVDD.n5388 VSS 0.281047f
C15673 DVDD.n5389 VSS 0.281047f
C15674 DVDD.n5390 VSS 0.281047f
C15675 DVDD.n5391 VSS 0.281047f
C15676 DVDD.n5392 VSS 0.281047f
C15677 DVDD.n5393 VSS 0.281047f
C15678 DVDD.n5394 VSS 0.281047f
C15679 DVDD.n5395 VSS 0.281047f
C15680 DVDD.n5396 VSS 0.281047f
C15681 DVDD.n5397 VSS 0.281047f
C15682 DVDD.n5398 VSS 0.281047f
C15683 DVDD.n5399 VSS 0.233546f
C15684 DVDD.n5400 VSS 0.233546f
C15685 DVDD.n5401 VSS 0.338444f
C15686 DVDD.n5402 VSS 0.095991f
C15687 DVDD.n5403 VSS 0.188025f
C15688 DVDD.n5404 VSS 0.140524f
C15689 DVDD.n5405 VSS 0.281047f
C15690 DVDD.n5406 VSS 0.281047f
C15691 DVDD.n5407 VSS 0.130628f
C15692 DVDD.n5408 VSS 0.015871f
C15693 DVDD.n5409 VSS 0.015871f
C15694 DVDD.n5410 VSS 0.015871f
C15695 DVDD.n5411 VSS 0.015871f
C15696 DVDD.n5412 VSS 0.015871f
C15697 DVDD.n5413 VSS 0.015871f
C15698 DVDD.n5414 VSS 0.015871f
C15699 DVDD.n5415 VSS 0.015871f
C15700 DVDD.n5416 VSS 0.015871f
C15701 DVDD.n5417 VSS 0.092033f
C15702 DVDD.n5418 VSS 0.015871f
C15703 DVDD.n5419 VSS 0.018174f
C15704 DVDD.n5420 VSS 3.87861f
C15705 DVDD.n5422 VSS 3.95424f
C15706 DVDD.n5423 VSS 0.015999f
C15707 DVDD.n5424 VSS 0.614473f
C15708 DVDD.n5425 VSS 0.148702f
C15709 DVDD.n5426 VSS 0.060206f
C15710 DVDD.n5427 VSS 0.027215f
C15711 DVDD.n5428 VSS 0.016673f
C15712 DVDD.n5429 VSS 0.091044f
C15713 DVDD.n5430 VSS 0.023765f
C15714 DVDD.n5431 VSS 0.029828f
C15715 DVDD.n5432 VSS 0.018512f
C15716 DVDD.n5433 VSS 0.070763f
C15717 DVDD.n5434 VSS 0.070763f
C15718 DVDD.n5435 VSS 0.070763f
C15719 DVDD.n5436 VSS 0.026256f
C15720 DVDD.n5437 VSS 0.070763f
C15721 DVDD.n5438 VSS 0.026256f
C15722 DVDD.n5439 VSS 0.070763f
C15723 DVDD.n5440 VSS 0.070763f
C15724 DVDD.n5441 VSS 0.024148f
C15725 DVDD.n5442 VSS 0.025873f
C15726 DVDD.n5443 VSS 0.070763f
C15727 DVDD.n5444 VSS 0.026256f
C15728 DVDD.n5445 VSS 0.070763f
C15729 DVDD.n5446 VSS 0.026256f
C15730 DVDD.n5447 VSS 0.070763f
C15731 DVDD.n5448 VSS 0.026256f
C15732 DVDD.n5449 VSS 0.070763f
C15733 DVDD.n5450 VSS 0.026256f
C15734 DVDD.n5451 VSS 0.070763f
C15735 DVDD.n5452 VSS 0.026256f
C15736 DVDD.n5453 VSS 0.070763f
C15737 DVDD.n5454 VSS 0.026256f
C15738 DVDD.n5455 VSS 0.070763f
C15739 DVDD.n5456 VSS 0.038806f
C15740 DVDD.n5457 VSS 0.035382f
C15741 DVDD.n5458 VSS 0.023765f
C15742 DVDD.n5459 VSS 0.023956f
C15743 DVDD.n5460 VSS 0.067339f
C15744 DVDD.n5461 VSS 0.026256f
C15745 DVDD.n5462 VSS 0.070763f
C15746 DVDD.n5463 VSS 0.026256f
C15747 DVDD.n5464 VSS 0.070763f
C15748 DVDD.n5465 VSS 0.026256f
C15749 DVDD.n5466 VSS 0.070763f
C15750 DVDD.n5467 VSS 0.026256f
C15751 DVDD.n5468 VSS 0.070763f
C15752 DVDD.n5469 VSS 0.026256f
C15753 DVDD.n5470 VSS 0.070763f
C15754 DVDD.n5471 VSS 0.070763f
C15755 DVDD.n5472 VSS 0.026256f
C15756 DVDD.n5473 VSS 0.023764f
C15757 DVDD.n5474 VSS 0.140524f
C15758 DVDD.n5475 VSS 0.013032f
C15759 DVDD.n5476 VSS 0.011691f
C15760 DVDD.n5477 VSS 0.140524f
C15761 DVDD.n5478 VSS 0.01744f
C15762 DVDD.n5479 VSS 0.026256f
C15763 DVDD.n5480 VSS 0.070763f
C15764 DVDD.n5481 VSS 0.070763f
C15765 DVDD.n5482 VSS 0.025129f
C15766 DVDD.n5483 VSS 0.018808f
C15767 DVDD.n5484 VSS 0.024672f
C15768 DVDD.n5485 VSS -0.254989f
C15769 DVDD.n5486 VSS 0.035381f
C15770 DVDD.n5487 VSS 5.3752f
C15771 DVDD.n5488 VSS 2.06325f
C15772 DVDD.n5489 VSS 2.68118f
C15773 DVDD.n5490 VSS 0.881825f
C15774 DVDD.n5491 VSS 0.528763f
C15775 DVDD.n5492 VSS 6.16644f
C15776 DVDD.t176 VSS 4.705029f
C15777 DVDD.t64 VSS 4.80305f
C15778 DVDD.n5493 VSS 6.16644f
C15779 DVDD.t199 VSS 4.78523f
C15780 DVDD.t103 VSS 4.72285f
C15781 DVDD.t100 VSS 3.92977f
C15782 DVDD.n5494 VSS 6.16644f
C15783 DVDD.n5495 VSS 1.02061f
C15784 DVDD.t106 VSS 4.78523f
C15785 DVDD.n5496 VSS 6.16644f
C15786 DVDD.t79 VSS 4.705029f
C15787 DVDD.t195 VSS 4.80305f
C15788 DVDD.n5497 VSS 6.16644f
C15789 DVDD.n5498 VSS 0.888222f
C15790 DVDD.n5499 VSS 1.02588f
C15791 DVDD.n5500 VSS 6.16644f
C15792 DVDD.t85 VSS 4.00997f
C15793 DVDD.n5501 VSS 0.93566f
C15794 DVDD.n5502 VSS 8.47284f
C15795 DVDD.n5503 VSS 0.070927f
C15796 DVDD.n5504 VSS 0.027214f
C15797 DVDD.n5505 VSS 0.049477f
C15798 DVDD.n5506 VSS 0.035463f
C15799 DVDD.n5507 VSS 0.027214f
C15800 DVDD.n5508 VSS 0.056913f
C15801 DVDD.n5509 VSS 0.027214f
C15802 DVDD.n5510 VSS 0.070927f
C15803 DVDD.n5511 VSS 0.070927f
C15804 DVDD.n5512 VSS 0.031546f
C15805 DVDD.n5513 VSS 0.020098f
C15806 DVDD.n5514 VSS 0.070927f
C15807 DVDD.n5515 VSS 0.070927f
C15808 DVDD.n5516 VSS 0.070927f
C15809 DVDD.n5517 VSS 0.024532f
C15810 DVDD.n5518 VSS 0.070927f
C15811 DVDD.n5519 VSS 0.027215f
C15812 DVDD.n5520 VSS 0.070927f
C15813 DVDD.n5521 VSS 0.027215f
C15814 DVDD.n5522 VSS 0.070927f
C15815 DVDD.n5523 VSS 0.027215f
C15816 DVDD.n5524 VSS 0.070927f
C15817 DVDD.n5525 VSS 0.027215f
C15818 DVDD.n5526 VSS 0.070927f
C15819 DVDD.n5527 VSS 0.027215f
C15820 DVDD.n5528 VSS 0.070927f
C15821 DVDD.n5529 VSS 0.027215f
C15822 DVDD.n5530 VSS 0.070927f
C15823 DVDD.n5531 VSS 0.070927f
C15824 DVDD.n5532 VSS 0.026065f
C15825 DVDD.n5533 VSS 0.024915f
C15826 DVDD.n5534 VSS 0.070927f
C15827 DVDD.n5535 VSS 0.027215f
C15828 DVDD.n5536 VSS 0.070927f
C15829 DVDD.n5537 VSS 0.027215f
C15830 DVDD.n5538 VSS 0.047475f
C15831 DVDD.n5539 VSS 0.035463f
C15832 DVDD.n5540 VSS 0.027215f
C15833 DVDD.n5541 VSS 0.058915f
C15834 DVDD.n5542 VSS 0.027215f
C15835 DVDD.n5543 VSS 0.070927f
C15836 DVDD.n5544 VSS 0.027215f
C15837 DVDD.n5545 VSS 0.070927f
C15838 DVDD.n5546 VSS 0.027215f
C15839 DVDD.n5547 VSS 0.070927f
C15840 DVDD.n5548 VSS 0.070927f
C15841 DVDD.n5549 VSS 0.025681f
C15842 DVDD.n5550 VSS 0.025298f
C15843 DVDD.n5551 VSS 0.070927f
C15844 DVDD.n5552 VSS 0.027215f
C15845 DVDD.n5553 VSS 0.070927f
C15846 DVDD.n5554 VSS 0.027215f
C15847 DVDD.n5555 VSS 0.070927f
C15848 DVDD.n5556 VSS 0.027215f
C15849 DVDD.n5557 VSS 0.070927f
C15850 DVDD.n5558 VSS 0.027215f
C15851 DVDD.n5559 VSS 0.070927f
C15852 DVDD.n5560 VSS 0.027215f
C15853 DVDD.n5561 VSS 0.066065f
C15854 DVDD.n5562 VSS -0.172196f
C15855 DVDD.n5563 VSS 0.01399f
C15856 DVDD.n5564 VSS 0.070927f
C15857 DVDD.n5565 VSS 0.140524f
C15858 DVDD.n5566 VSS 0.140524f
C15859 DVDD.n5567 VSS 0.026256f
C15860 DVDD.n5568 VSS 0.02089f
C15861 DVDD.n5569 VSS 0.004024f
C15862 DVDD.n5570 VSS 0.010924f
C15863 DVDD.n5571 VSS 0.017823f
C15864 DVDD.n5572 VSS 0.003258f
C15865 DVDD.n5573 VSS 0.007857f
C15866 DVDD.n5574 VSS 0.014757f
C15867 DVDD.n5575 VSS 0.021657f
C15868 DVDD.n5576 VSS 0.004791f
C15869 DVDD.n5577 VSS 0.281047f
C15870 DVDD.n5578 VSS 0.281047f
C15871 DVDD.n5579 VSS 0.281047f
C15872 DVDD.n5580 VSS 0.281047f
C15873 DVDD.n5581 VSS 0.281047f
C15874 DVDD.n5582 VSS 0.281047f
C15875 DVDD.n5583 VSS 0.281047f
C15876 DVDD.n5584 VSS 0.281047f
C15877 DVDD.n5585 VSS 0.281047f
C15878 DVDD.n5586 VSS 0.281047f
C15879 DVDD.n5587 VSS 0.281047f
C15880 DVDD.n5588 VSS 0.281047f
C15881 DVDD.n5589 VSS 0.253338f
C15882 DVDD.n5590 VSS 0.031667f
C15883 DVDD.n5591 VSS 0.399293f
C15884 DVDD.n5592 VSS 1.29492f
C15885 DVDD.n5593 VSS 0.253338f
C15886 DVDD.n5594 VSS 0.253338f
C15887 DVDD.n5595 VSS 0.281047f
C15888 DVDD.n5596 VSS 0.281047f
C15889 DVDD.n5597 VSS 0.281047f
C15890 DVDD.n5598 VSS 0.281047f
C15891 DVDD.n5599 VSS 0.281047f
C15892 DVDD.n5600 VSS 0.281047f
C15893 DVDD.n5601 VSS 0.281047f
C15894 DVDD.n5602 VSS 0.281047f
C15895 DVDD.n5603 VSS 0.197921f
C15896 DVDD.n5604 VSS 0.001341f
C15897 DVDD.n5605 VSS 0.018207f
C15898 DVDD.n5606 VSS 0.011307f
C15899 DVDD.n5607 VSS 0.004408f
C15900 DVDD.n5608 VSS 0.021273f
C15901 DVDD.n5609 VSS 0.014374f
C15902 DVDD.n5610 VSS 0.007474f
C15903 DVDD.n5611 VSS 0.026256f
C15904 DVDD.n5612 VSS 0.070927f
C15905 DVDD.n5613 VSS 0.026256f
C15906 DVDD.n5614 VSS 0.070927f
C15907 DVDD.n5615 VSS 0.070927f
C15908 DVDD.n5616 VSS 0.024148f
C15909 DVDD.n5617 VSS 0.025873f
C15910 DVDD.n5618 VSS 0.070927f
C15911 DVDD.n5619 VSS 0.026256f
C15912 DVDD.n5620 VSS 0.070927f
C15913 DVDD.n5621 VSS 0.026256f
C15914 DVDD.n5622 VSS 0.070927f
C15915 DVDD.n5623 VSS 0.026256f
C15916 DVDD.n5624 VSS 0.070927f
C15917 DVDD.n5625 VSS 0.026256f
C15918 DVDD.n5626 VSS 0.070927f
C15919 DVDD.n5627 VSS 0.026256f
C15920 DVDD.n5628 VSS 0.070927f
C15921 DVDD.n5629 VSS 0.026256f
C15922 DVDD.n5630 VSS 0.070927f
C15923 DVDD.n5631 VSS 0.038895f
C15924 DVDD.n5632 VSS 0.035463f
C15925 DVDD.n5633 VSS 0.023765f
C15926 DVDD.n5634 VSS 0.023956f
C15927 DVDD.n5635 VSS 0.067495f
C15928 DVDD.n5636 VSS 0.026256f
C15929 DVDD.n5637 VSS 0.070927f
C15930 DVDD.n5638 VSS 0.026256f
C15931 DVDD.n5639 VSS 0.070927f
C15932 DVDD.n5640 VSS 0.026256f
C15933 DVDD.n5641 VSS 0.070927f
C15934 DVDD.n5642 VSS 0.026256f
C15935 DVDD.n5643 VSS 0.070927f
C15936 DVDD.n5644 VSS 0.026256f
C15937 DVDD.n5645 VSS 0.070927f
C15938 DVDD.n5646 VSS 0.026256f
C15939 DVDD.n5647 VSS 0.070927f
C15940 DVDD.n5648 VSS 0.070927f
C15941 DVDD.n5649 VSS 9.58e-19
C15942 DVDD.n5650 VSS 0.023765f
C15943 DVDD.n5651 VSS 0.140524f
C15944 DVDD.n5652 VSS 0.01744f
C15945 DVDD.n5653 VSS 0.026256f
C15946 DVDD.n5654 VSS 0.070927f
C15947 DVDD.n5655 VSS 0.070927f
C15948 DVDD.n5656 VSS 0.025129f
C15949 DVDD.n5657 VSS 0.018808f
C15950 DVDD.n5658 VSS 0.024672f
C15951 DVDD.n5659 VSS -0.254896f
C15952 DVDD.n5660 VSS 0.035463f
C15953 DVDD.n5661 VSS 5.39089f
C15954 DVDD.n5662 VSS 2.07216f
C15955 DVDD.n5663 VSS 2.6901f
C15956 DVDD.n5664 VSS 0.883168f
C15957 DVDD.n5665 VSS 0.030555f
C15958 DVDD.n5666 VSS 0.018174f
C15959 DVDD.n5667 VSS 0.045832f
C15960 DVDD.n5668 VSS 0.018174f
C15961 DVDD.n5669 VSS 0.06111f
C15962 DVDD.n5670 VSS 0.018174f
C15963 DVDD.n5671 VSS 0.06111f
C15964 DVDD.n5672 VSS 0.06111f
C15965 DVDD.n5673 VSS 0.06111f
C15966 DVDD.n5674 VSS 0.015999f
C15967 DVDD.n5675 VSS 0.281047f
C15968 DVDD.n5676 VSS 0.281047f
C15969 DVDD.n5677 VSS 0.281047f
C15970 DVDD.n5678 VSS 0.281047f
C15971 DVDD.n5679 VSS 0.281047f
C15972 DVDD.n5680 VSS 0.281047f
C15973 DVDD.n5681 VSS 0.281047f
C15974 DVDD.n5682 VSS 0.281047f
C15975 DVDD.n5683 VSS 0.281047f
C15976 DVDD.n5684 VSS 0.281047f
C15977 DVDD.n5685 VSS 0.281047f
C15978 DVDD.n5686 VSS 0.253338f
C15979 DVDD.n5687 VSS 0.281047f
C15980 DVDD.n5688 VSS 0.144482f
C15981 DVDD.n5689 VSS 0.399293f
C15982 DVDD.n5690 VSS 1.29492f
C15983 DVDD.n5691 VSS 0.253338f
C15984 DVDD.n5692 VSS 0.281047f
C15985 DVDD.n5693 VSS 0.281047f
C15986 DVDD.n5694 VSS 0.281047f
C15987 DVDD.n5695 VSS 0.281047f
C15988 DVDD.n5696 VSS 0.281047f
C15989 DVDD.n5697 VSS 0.281047f
C15990 DVDD.n5698 VSS 0.281047f
C15991 DVDD.n5699 VSS 0.281047f
C15992 DVDD.n5700 VSS 0.281047f
C15993 DVDD.n5701 VSS 0.281047f
C15994 DVDD.n5702 VSS 0.281047f
C15995 DVDD.n5703 VSS 0.121721f
C15996 DVDD.n5704 VSS 0.090054f
C15997 DVDD.n5705 VSS 0.015871f
C15998 DVDD.n5706 VSS 0.057397f
C15999 DVDD.n5707 VSS 0.101929f
C16000 DVDD.n5708 VSS 0.06455f
C16001 DVDD.n5709 VSS 0.140524f
C16002 DVDD.n5710 VSS 0.167243f
C16003 DVDD.n5711 VSS 0.257297f
C16004 DVDD.n5712 VSS 0.338444f
C16005 DVDD.n5713 VSS 0.164274f
C16006 DVDD.n5714 VSS 0.164274f
C16007 DVDD.n5715 VSS 0.281047f
C16008 DVDD.n5716 VSS 0.281047f
C16009 DVDD.n5717 VSS 0.281047f
C16010 DVDD.n5718 VSS 0.281047f
C16011 DVDD.n5719 VSS 0.281047f
C16012 DVDD.n5720 VSS 0.281047f
C16013 DVDD.n5721 VSS 0.281047f
C16014 DVDD.n5722 VSS 0.281047f
C16015 DVDD.n5723 VSS 0.281047f
C16016 DVDD.n5724 VSS 0.281047f
C16017 DVDD.n5725 VSS 0.281047f
C16018 DVDD.n5726 VSS 0.281047f
C16019 DVDD.n5727 VSS 0.281047f
C16020 DVDD.n5728 VSS 0.281047f
C16021 DVDD.n5729 VSS 0.153388f
C16022 DVDD.n5730 VSS 0.00998f
C16023 DVDD.n5731 VSS 0.011429f
C16024 DVDD.n5732 VSS 0.063742f
C16025 DVDD.n5733 VSS 0.00586f
C16026 DVDD.n5734 VSS 0.027607f
C16027 DVDD.n5735 VSS 0.140524f
C16028 DVDD.n5736 VSS 0.00998f
C16029 DVDD.n5737 VSS 0.011429f
C16030 DVDD.n5738 VSS 0.019961f
C16031 DVDD.n5739 VSS 0.019961f
C16032 DVDD.n5740 VSS 0.01312f
C16033 DVDD.n5741 VSS 0.019961f
C16034 DVDD.n5742 VSS 0.018834f
C16035 DVDD.n5743 VSS 0.019961f
C16036 DVDD.n5744 VSS 0.019961f
C16037 DVDD.n5745 VSS 0.011107f
C16038 DVDD.n5746 VSS 0.010302f
C16039 DVDD.n5747 VSS 0.019961f
C16040 DVDD.n5748 VSS 0.011429f
C16041 DVDD.n5749 VSS 0.019961f
C16042 DVDD.n5750 VSS 0.011429f
C16043 DVDD.n5751 VSS 0.019961f
C16044 DVDD.n5752 VSS 0.011429f
C16045 DVDD.n5753 VSS 0.019961f
C16046 DVDD.n5754 VSS 0.011429f
C16047 DVDD.n5755 VSS 0.019961f
C16048 DVDD.n5756 VSS 0.011429f
C16049 DVDD.n5757 VSS 0.019961f
C16050 DVDD.n5758 VSS 0.011429f
C16051 DVDD.n5759 VSS 0.019961f
C16052 DVDD.n5760 VSS 0.019961f
C16053 DVDD.n5761 VSS 0.010946f
C16054 DVDD.n5762 VSS 0.010463f
C16055 DVDD.n5763 VSS 0.019961f
C16056 DVDD.n5764 VSS 0.011429f
C16057 DVDD.n5765 VSS 0.019961f
C16058 DVDD.n5766 VSS 0.011429f
C16059 DVDD.n5767 VSS 0.019961f
C16060 DVDD.n5768 VSS 0.011429f
C16061 DVDD.n5769 VSS 0.019961f
C16062 DVDD.n5770 VSS 0.011429f
C16063 DVDD.n5771 VSS 0.019961f
C16064 DVDD.n5772 VSS 0.011429f
C16065 DVDD.n5773 VSS 0.019961f
C16066 DVDD.n5774 VSS 0.019961f
C16067 DVDD.n5775 VSS 0.011429f
C16068 DVDD.n5776 VSS 0.019961f
C16069 DVDD.n5777 VSS 0.011429f
C16070 DVDD.n5778 VSS 0.019961f
C16071 DVDD.n5779 VSS 0.011429f
C16072 DVDD.n5780 VSS 0.019961f
C16073 DVDD.n5781 VSS 0.019961f
C16074 DVDD.n5782 VSS 0.019961f
C16075 DVDD.n5783 VSS 0.010785f
C16076 DVDD.n5784 VSS 0.00998f
C16077 DVDD.n5785 VSS 0.140524f
C16078 DVDD.n5786 VSS 0.00998f
C16079 DVDD.n5787 VSS 0.011429f
C16080 DVDD.n5788 VSS 0.019961f
C16081 DVDD.n5789 VSS -0.36209f
C16082 DVDD.n5790 VSS 0.012073f
C16083 DVDD.n5791 VSS 0.019961f
C16084 DVDD.n5792 VSS 0.015856f
C16085 DVDD.n5793 VSS 0.019961f
C16086 DVDD.n5794 VSS 0.019961f
C16087 DVDD.n5795 VSS 0.011429f
C16088 DVDD.n5796 VSS 0.019961f
C16089 DVDD.n5797 VSS 0.019961f
C16090 DVDD.n5798 VSS 0.010544f
C16091 DVDD.n5799 VSS 0.010866f
C16092 DVDD.n5800 VSS 0.019961f
C16093 DVDD.n5801 VSS 0.011429f
C16094 DVDD.n5802 VSS 0.019961f
C16095 DVDD.n5803 VSS 0.011429f
C16096 DVDD.n5804 VSS 0.019961f
C16097 DVDD.n5805 VSS 0.011429f
C16098 DVDD.n5806 VSS 0.019961f
C16099 DVDD.n5807 VSS 0.011429f
C16100 DVDD.n5808 VSS 0.019961f
C16101 DVDD.n5809 VSS 0.011429f
C16102 DVDD.n5810 VSS 0.019961f
C16103 DVDD.n5811 VSS 0.011429f
C16104 DVDD.n5812 VSS 0.019961f
C16105 DVDD.n5813 VSS 0.019961f
C16106 DVDD.n5814 VSS 0.010383f
C16107 DVDD.n5815 VSS 0.011027f
C16108 DVDD.n5816 VSS 0.019961f
C16109 DVDD.n5817 VSS 0.011429f
C16110 DVDD.n5818 VSS 0.019961f
C16111 DVDD.n5819 VSS 0.011429f
C16112 DVDD.n5820 VSS 0.019961f
C16113 DVDD.n5821 VSS 0.011429f
C16114 DVDD.n5822 VSS 0.019961f
C16115 DVDD.n5823 VSS 0.011429f
C16116 DVDD.n5824 VSS 0.019961f
C16117 DVDD.n5825 VSS 0.011429f
C16118 DVDD.n5826 VSS 0.019961f
C16119 DVDD.n5827 VSS 0.011429f
C16120 DVDD.n5828 VSS 0.019961f
C16121 DVDD.n5829 VSS 0.019961f
C16122 DVDD.n5830 VSS 0.010222f
C16123 DVDD.n5831 VSS 0.011188f
C16124 DVDD.n5832 VSS 0.019961f
C16125 DVDD.n5833 VSS 0.019961f
C16126 DVDD.n5834 VSS 0.011429f
C16127 DVDD.n5835 VSS 0.00998f
C16128 DVDD.n5836 VSS 0.140524f
C16129 DVDD.n5837 VSS 0.00998f
C16130 DVDD.n5838 VSS 0.011429f
C16131 DVDD.n5839 VSS 0.019961f
C16132 DVDD.n5840 VSS 0.019961f
C16133 DVDD.n5841 VSS 0.015051f
C16134 DVDD.n5842 VSS 0.019961f
C16135 DVDD.n5843 VSS 0.014971f
C16136 DVDD.n5844 VSS 0.019961f
C16137 DVDD.n5845 VSS 0.011429f
C16138 DVDD.n5846 VSS 0.019961f
C16139 DVDD.n5847 VSS 0.011429f
C16140 DVDD.n5848 VSS 0.061904f
C16141 DVDD.n5849 VSS 0.005232f
C16142 DVDD.n5850 VSS 0.025252f
C16143 DVDD.n5851 VSS 0.140524f
C16144 DVDD.n5852 VSS 0.268182f
C16145 DVDD.n5853 VSS 0.281047f
C16146 DVDD.n5854 VSS 0.281047f
C16147 DVDD.n5855 VSS 0.281047f
C16148 DVDD.n5856 VSS 0.281047f
C16149 DVDD.n5857 VSS 0.281047f
C16150 DVDD.n5858 VSS 0.153388f
C16151 DVDD.n5859 VSS 0.281047f
C16152 DVDD.n5860 VSS 0.281047f
C16153 DVDD.n5861 VSS 0.281047f
C16154 DVDD.n5862 VSS 0.281047f
C16155 DVDD.n5863 VSS 0.281047f
C16156 DVDD.n5864 VSS 0.281047f
C16157 DVDD.n5865 VSS 0.281047f
C16158 DVDD.n5866 VSS 0.281047f
C16159 DVDD.n5867 VSS 0.281047f
C16160 DVDD.n5868 VSS 0.281047f
C16161 DVDD.n5869 VSS 0.281047f
C16162 DVDD.n5870 VSS 0.281047f
C16163 DVDD.n5871 VSS 0.281047f
C16164 DVDD.n5872 VSS 0.281047f
C16165 DVDD.n5873 VSS 0.281047f
C16166 DVDD.n5874 VSS 0.281047f
C16167 DVDD.n5875 VSS 0.281047f
C16168 DVDD.n5876 VSS 0.164274f
C16169 DVDD.n5877 VSS 0.164274f
C16170 DVDD.n5878 VSS 0.164274f
C16171 DVDD.n5879 VSS 0.338444f
C16172 DVDD.n5880 VSS 0.257297f
C16173 DVDD.n5881 VSS 0.257297f
C16174 DVDD.n5882 VSS 0.281047f
C16175 DVDD.n5883 VSS 0.121721f
C16176 DVDD.n5884 VSS 0.281047f
C16177 DVDD.n5885 VSS 0.281047f
C16178 DVDD.n5886 VSS 0.281047f
C16179 DVDD.n5887 VSS 0.281047f
C16180 DVDD.n5888 VSS 0.281047f
C16181 DVDD.n5889 VSS 0.281047f
C16182 DVDD.n5890 VSS 0.281047f
C16183 DVDD.n5891 VSS 0.281047f
C16184 DVDD.n5892 VSS 0.281047f
C16185 DVDD.n5893 VSS 0.281047f
C16186 DVDD.n5894 VSS 0.281047f
C16187 DVDD.n5895 VSS 0.253338f
C16188 DVDD.n5896 VSS 0.031667f
C16189 DVDD.n5897 VSS 0.399293f
C16190 DVDD.n5898 VSS 1.29492f
C16191 DVDD.n5899 VSS 0.253338f
C16192 DVDD.n5900 VSS 0.253338f
C16193 DVDD.n5901 VSS 0.281047f
C16194 DVDD.n5902 VSS 0.281047f
C16195 DVDD.n5903 VSS 0.281047f
C16196 DVDD.n5904 VSS 0.281047f
C16197 DVDD.n5905 VSS 0.281047f
C16198 DVDD.n5906 VSS 0.281047f
C16199 DVDD.n5907 VSS 0.281047f
C16200 DVDD.n5908 VSS 0.281047f
C16201 DVDD.n5909 VSS 0.179118f
C16202 DVDD.n5910 VSS 0.015871f
C16203 DVDD.n5911 VSS 0.015871f
C16204 DVDD.n5912 VSS 0.015871f
C16205 DVDD.n5913 VSS 0.015871f
C16206 DVDD.n5914 VSS 0.057397f
C16207 DVDD.n5915 VSS 0.015871f
C16208 DVDD.n5916 VSS 0.020862f
C16209 DVDD.n5917 VSS 3.9735f
C16210 DVDD.n5918 VSS 0.015999f
C16211 DVDD.n5919 VSS 0.605223f
C16212 DVDD.n5920 VSS 0.148162f
C16213 DVDD.n5921 VSS 0.05901f
C16214 DVDD.n5922 VSS 0.140524f
C16215 DVDD.n5923 VSS 0.023765f
C16216 DVDD.n5924 VSS 0.027215f
C16217 DVDD.n5925 VSS 0.070927f
C16218 DVDD.n5926 VSS 0.070927f
C16219 DVDD.n5927 VSS 0.029828f
C16220 DVDD.n5928 VSS 0.018512f
C16221 DVDD.n5929 VSS 0.026211f
C16222 DVDD.n5930 VSS 0.070927f
C16223 DVDD.n5931 VSS 0.070927f
C16224 DVDD.n5932 VSS 0.026256f
C16225 DVDD.n5933 VSS 0.016482f
C16226 DVDD.n5934 VSS 0.140524f
C16227 DVDD.n5935 VSS 0.140524f
C16228 DVDD.n5936 VSS 0.281047f
C16229 DVDD.n5937 VSS 0.257297f
C16230 DVDD.n5938 VSS 0.167243f
C16231 DVDD.n5939 VSS 0.536365f
C16232 DVDD.n5940 VSS 0.536365f
C16233 DVDD.n5941 VSS 0.164274f
C16234 DVDD.n5942 VSS 0.164274f
C16235 DVDD.n5943 VSS 0.164274f
C16236 DVDD.n5944 VSS 0.536365f
C16237 DVDD.n5945 VSS 0.257297f
C16238 DVDD.n5946 VSS 0.281047f
C16239 DVDD.n5947 VSS 0.281047f
C16240 DVDD.n5948 VSS 0.281047f
C16241 DVDD.n5949 VSS 0.281047f
C16242 DVDD.n5950 VSS 0.173181f
C16243 DVDD.n5951 VSS 0.281047f
C16244 DVDD.n5952 VSS 0.281047f
C16245 DVDD.n5953 VSS 0.140524f
C16246 DVDD.n5954 VSS 0.140524f
C16247 DVDD.n5955 VSS 0.026266f
C16248 DVDD.n5956 VSS 0.140524f
C16249 DVDD.n5957 VSS 0.197921f
C16250 DVDD.n5958 VSS 0.281047f
C16251 DVDD.n5959 VSS 0.281047f
C16252 DVDD.n5960 VSS 0.281047f
C16253 DVDD.n5961 VSS 0.281047f
C16254 DVDD.n5962 VSS 0.281047f
C16255 DVDD.n5963 VSS 0.281047f
C16256 DVDD.n5964 VSS 0.281047f
C16257 DVDD.n5965 VSS 0.281047f
C16258 DVDD.n5966 VSS 0.281047f
C16259 DVDD.n5967 VSS 0.281047f
C16260 DVDD.n5968 VSS 0.281047f
C16261 DVDD.n5969 VSS 0.253338f
C16262 DVDD.n5970 VSS 0.253338f
C16263 DVDD.n5971 VSS 0.031667f
C16264 DVDD.n5972 VSS 0.399293f
C16265 DVDD.n5973 VSS 1.29492f
C16266 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n0 VSS 1.82434f
C16267 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t0 VSS 0.228818f
C16268 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t8 VSS 0.308392f
C16269 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t3 VSS 0.302472f
C16270 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n1 VSS 1.36191f
C16271 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t4 VSS 0.325049f
C16272 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t1 VSS 0.321259f
C16273 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t11 VSS 0.404429f
C16274 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t12 VSS 0.76375f
C16275 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n2 VSS 0.644041f
C16276 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t6 VSS 0.404429f
C16277 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t7 VSS 0.76375f
C16278 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n3 VSS 0.646847f
C16279 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t2 VSS 0.631504f
C16280 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t10 VSS 0.358296f
C16281 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t9 VSS 0.631504f
C16282 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t5 VSS 0.358296f
C16283 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n4 VSS 0.915343f
C16284 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n5 VSS 0.909193f
C16285 DVSS.n0 VSS 0.125986f
C16286 DVSS.n1 VSS 0.167293f
C16287 DVSS.n2 VSS 0.195519f
C16288 DVSS.n3 VSS 0.195519f
C16289 DVSS.n4 VSS 0.195519f
C16290 DVSS.n5 VSS 0.110151f
C16291 DVSS.n6 VSS 0.097759f
C16292 DVSS.n7 VSS 0.014208f
C16293 DVSS.n8 VSS 0.014208f
C16294 DVSS.n9 VSS 0.014208f
C16295 DVSS.n10 VSS 0.014208f
C16296 DVSS.n11 VSS 0.014208f
C16297 DVSS.n12 VSS 0.014208f
C16298 DVSS.n13 VSS 0.014208f
C16299 DVSS.n14 VSS 0.014208f
C16300 DVSS.n15 VSS 0.014208f
C16301 DVSS.n16 VSS 0.014208f
C16302 DVSS.n17 VSS 0.014208f
C16303 DVSS.n18 VSS 0.014208f
C16304 DVSS.n19 VSS 0.014208f
C16305 DVSS.n20 VSS 0.014208f
C16306 DVSS.n21 VSS 0.014208f
C16307 DVSS.n22 VSS 0.014208f
C16308 DVSS.n23 VSS 0.014208f
C16309 DVSS.n24 VSS 0.014208f
C16310 DVSS.n25 VSS 0.007104f
C16311 DVSS.n26 VSS 0.245123f
C16312 DVSS.n27 VSS 0.195519f
C16313 DVSS.n28 VSS 0.177619f
C16314 DVSS.n29 VSS 0.195519f
C16315 DVSS.n30 VSS 0.195519f
C16316 DVSS.n31 VSS 0.195519f
C16317 DVSS.n32 VSS 0.195519f
C16318 DVSS.n33 VSS 0.195519f
C16319 DVSS.n34 VSS 0.195519f
C16320 DVSS.n35 VSS 0.195519f
C16321 DVSS.n36 VSS 0.195519f
C16322 DVSS.n37 VSS 0.195519f
C16323 DVSS.n38 VSS 0.195519f
C16324 DVSS.n39 VSS 0.195519f
C16325 DVSS.n40 VSS 0.235449f
C16326 DVSS.n41 VSS 0.235449f
C16327 DVSS.n42 VSS 0.114282f
C16328 DVSS.n43 VSS 0.235449f
C16329 DVSS.n44 VSS 0.114282f
C16330 DVSS.n45 VSS 0.195519f
C16331 DVSS.n46 VSS 0.373138f
C16332 DVSS.n47 VSS 0.235449f
C16333 DVSS.n48 VSS 0.097759f
C16334 DVSS.n49 VSS 0.195519f
C16335 DVSS.n50 VSS 0.140443f
C16336 DVSS.n51 VSS 0.195519f
C16337 DVSS.n52 VSS 0.195519f
C16338 DVSS.n53 VSS 0.195519f
C16339 DVSS.n54 VSS 0.124609f
C16340 DVSS.n55 VSS 0.001932f
C16341 DVSS.n56 VSS 0.022822f
C16342 DVSS.n57 VSS 0.025524f
C16343 DVSS.n58 VSS 0.044051f
C16344 DVSS.t141 VSS 4.56431f
C16345 DVSS.n60 VSS 0.81856f
C16346 DVSS.n61 VSS 0.22488f
C16347 DVSS.n62 VSS 0.05105f
C16348 DVSS.n63 VSS 0.022822f
C16349 DVSS.n64 VSS 0.05105f
C16350 DVSS.n65 VSS 0.022822f
C16351 DVSS.n66 VSS 0.05105f
C16352 DVSS.n67 VSS 0.022822f
C16353 DVSS.n68 VSS 0.05105f
C16354 DVSS.n69 VSS 0.022822f
C16355 DVSS.n70 VSS 0.05105f
C16356 DVSS.n71 VSS 0.022822f
C16357 DVSS.n72 VSS 0.022822f
C16358 DVSS.n73 VSS 0.022822f
C16359 DVSS.n74 VSS 0.05105f
C16360 DVSS.n75 VSS 0.05105f
C16361 DVSS.n76 VSS 0.05105f
C16362 DVSS.n77 VSS 0.022822f
C16363 DVSS.n78 VSS 0.022822f
C16364 DVSS.n79 VSS 0.022822f
C16365 DVSS.n80 VSS 0.05105f
C16366 DVSS.n81 VSS 0.05105f
C16367 DVSS.n82 VSS 0.05105f
C16368 DVSS.n83 VSS 0.022822f
C16369 DVSS.n84 VSS 0.022822f
C16370 DVSS.n85 VSS 0.022822f
C16371 DVSS.n86 VSS 0.05105f
C16372 DVSS.n87 VSS 0.05105f
C16373 DVSS.n88 VSS 0.05105f
C16374 DVSS.n89 VSS 0.022822f
C16375 DVSS.n90 VSS 0.022822f
C16376 DVSS.n91 VSS 0.022822f
C16377 DVSS.n92 VSS 0.05105f
C16378 DVSS.n93 VSS 0.05105f
C16379 DVSS.n94 VSS 0.05105f
C16380 DVSS.n95 VSS 0.022822f
C16381 DVSS.n96 VSS 0.022822f
C16382 DVSS.n97 VSS 0.022822f
C16383 DVSS.n98 VSS 0.05105f
C16384 DVSS.n99 VSS 0.05105f
C16385 DVSS.n100 VSS 0.05105f
C16386 DVSS.n101 VSS 0.012791f
C16387 DVSS.n102 VSS 0.168669f
C16388 DVSS.n103 VSS 0.140443f
C16389 DVSS.n104 VSS 0.195519f
C16390 DVSS.n105 VSS 0.097759f
C16391 DVSS.n106 VSS 0.071599f
C16392 DVSS.n107 VSS 0.114282f
C16393 DVSS.n108 VSS 0.195519f
C16394 DVSS.n109 VSS 0.195519f
C16395 DVSS.n110 VSS 0.195519f
C16396 DVSS.n111 VSS 0.195519f
C16397 DVSS.n112 VSS 0.195519f
C16398 DVSS.n113 VSS 0.195519f
C16399 DVSS.n114 VSS 0.195519f
C16400 DVSS.n115 VSS 0.195519f
C16401 DVSS.n116 VSS 0.195519f
C16402 DVSS.n117 VSS 0.195519f
C16403 DVSS.n118 VSS 0.195519f
C16404 DVSS.n119 VSS 0.195519f
C16405 DVSS.n120 VSS 0.195519f
C16406 DVSS.n121 VSS 0.195519f
C16407 DVSS.n122 VSS 0.195519f
C16408 DVSS.n123 VSS 0.427345f
C16409 DVSS.n124 VSS 0.195519f
C16410 DVSS.n125 VSS 0.195519f
C16411 DVSS.n126 VSS 0.195519f
C16412 DVSS.n127 VSS 0.173489f
C16413 DVSS.n128 VSS 0.173489f
C16414 DVSS.n129 VSS 0.373138f
C16415 DVSS.n130 VSS 0.195519f
C16416 DVSS.n131 VSS 0.195519f
C16417 DVSS.n132 VSS 0.11979f
C16418 DVSS.n133 VSS 0.235449f
C16419 DVSS.n134 VSS 0.11979f
C16420 DVSS.n135 VSS 0.173489f
C16421 DVSS.n136 VSS 0.195519f
C16422 DVSS.n137 VSS 0.195519f
C16423 DVSS.n138 VSS 0.195519f
C16424 DVSS.n139 VSS 0.195519f
C16425 DVSS.n140 VSS 0.195519f
C16426 DVSS.n141 VSS 0.116347f
C16427 DVSS.n142 VSS 0.195519f
C16428 DVSS.n143 VSS 0.195519f
C16429 DVSS.n144 VSS 0.116347f
C16430 DVSS.n145 VSS 0.195519f
C16431 DVSS.n146 VSS 0.195519f
C16432 DVSS.n147 VSS 0.195519f
C16433 DVSS.n148 VSS 0.195519f
C16434 DVSS.n149 VSS 0.195519f
C16435 DVSS.n150 VSS 0.173489f
C16436 DVSS.n151 VSS 0.173489f
C16437 DVSS.n152 VSS 0.195519f
C16438 DVSS.n153 VSS 0.195519f
C16439 DVSS.n154 VSS 0.195519f
C16440 DVSS.n155 VSS 0.235449f
C16441 DVSS.n156 VSS 0.195519f
C16442 DVSS.n157 VSS 0.195519f
C16443 DVSS.n158 VSS 0.195519f
C16444 DVSS.n159 VSS 0.195519f
C16445 DVSS.n160 VSS 0.195519f
C16446 DVSS.n161 VSS 0.195519f
C16447 DVSS.n162 VSS 0.195519f
C16448 DVSS.n163 VSS 0.195519f
C16449 DVSS.n164 VSS 0.195519f
C16450 DVSS.n165 VSS 0.195519f
C16451 DVSS.n166 VSS 0.195519f
C16452 DVSS.n167 VSS 0.195519f
C16453 DVSS.n168 VSS 0.161785f
C16454 DVSS.n169 VSS 0.480814f
C16455 DVSS.n170 VSS 0.161785f
C16456 DVSS.n171 VSS 0.195519f
C16457 DVSS.n172 VSS 0.195519f
C16458 DVSS.n173 VSS 0.195519f
C16459 DVSS.n174 VSS 0.195519f
C16460 DVSS.n175 VSS 0.195519f
C16461 DVSS.n176 VSS 0.195519f
C16462 DVSS.n177 VSS 0.195519f
C16463 DVSS.n178 VSS 0.195519f
C16464 DVSS.n179 VSS 0.195519f
C16465 DVSS.n180 VSS 0.195519f
C16466 DVSS.n181 VSS 0.195519f
C16467 DVSS.n182 VSS 0.195519f
C16468 DVSS.n183 VSS 0.195519f
C16469 DVSS.n184 VSS 0.235449f
C16470 DVSS.n185 VSS 0.235449f
C16471 DVSS.n186 VSS 0.373138f
C16472 DVSS.n187 VSS 0.195519f
C16473 DVSS.n188 VSS 0.195519f
C16474 DVSS.n189 VSS 0.183815f
C16475 DVSS.n190 VSS 0.195519f
C16476 DVSS.n191 VSS 0.195519f
C16477 DVSS.n192 VSS 0.195519f
C16478 DVSS.n193 VSS 0.195519f
C16479 DVSS.n194 VSS 0.480814f
C16480 DVSS.n195 VSS 0.109463f
C16481 DVSS.n196 VSS 0.195519f
C16482 DVSS.n197 VSS 0.195519f
C16483 DVSS.n198 VSS 0.195519f
C16484 DVSS.n199 VSS 0.195519f
C16485 DVSS.n200 VSS 0.125297f
C16486 DVSS.n201 VSS 0.195519f
C16487 DVSS.n202 VSS 0.125297f
C16488 DVSS.n203 VSS 0.235449f
C16489 DVSS.n204 VSS 0.125297f
C16490 DVSS.n205 VSS 0.195519f
C16491 DVSS.n206 VSS 0.195519f
C16492 DVSS.n207 VSS 0.195519f
C16493 DVSS.n208 VSS 0.195519f
C16494 DVSS.n209 VSS 0.195519f
C16495 DVSS.n210 VSS 0.195519f
C16496 DVSS.n211 VSS 0.195519f
C16497 DVSS.n212 VSS 0.195519f
C16498 DVSS.n213 VSS 0.195519f
C16499 DVSS.n214 VSS 0.195519f
C16500 DVSS.n215 VSS 0.195519f
C16501 DVSS.n216 VSS 0.195519f
C16502 DVSS.n217 VSS 0.195519f
C16503 DVSS.n218 VSS 0.195519f
C16504 DVSS.n219 VSS 0.195519f
C16505 DVSS.n220 VSS 0.195519f
C16506 DVSS.n221 VSS 0.195519f
C16507 DVSS.n222 VSS 0.195519f
C16508 DVSS.n223 VSS 0.195519f
C16509 DVSS.n224 VSS 0.135624f
C16510 DVSS.n225 VSS 0.195519f
C16511 DVSS.n226 VSS 0.195519f
C16512 DVSS.n227 VSS 0.195519f
C16513 DVSS.n228 VSS 0.107398f
C16514 DVSS.n229 VSS 0.255315f
C16515 DVSS.n230 VSS 0.025155f
C16516 DVSS.n231 VSS 0.053611f
C16517 DVSS.n232 VSS 0.025155f
C16518 DVSS.n233 VSS 0.053611f
C16519 DVSS.n234 VSS 0.025155f
C16520 DVSS.n235 VSS 0.053611f
C16521 DVSS.n236 VSS 0.025155f
C16522 DVSS.n237 VSS 0.053611f
C16523 DVSS.n238 VSS 0.025155f
C16524 DVSS.n239 VSS 0.053611f
C16525 DVSS.n240 VSS 0.025155f
C16526 DVSS.n241 VSS 0.026805f
C16527 DVSS.n242 VSS 0.003246f
C16528 DVSS.n243 VSS 0.152835f
C16529 DVSS.n244 VSS 0.157654f
C16530 DVSS.n245 VSS 0.162473f
C16531 DVSS.n246 VSS 0.195519f
C16532 DVSS.n247 VSS 3.341f
C16533 DVSS.n248 VSS 3.56769f
C16534 DVSS.n249 VSS 1.78032f
C16535 DVSS.n250 VSS 0.955224f
C16536 DVSS.n251 VSS 3.56769f
C16537 DVSS.n252 VSS 0.097759f
C16538 DVSS.n253 VSS 0.897965f
C16539 DVSS.n254 VSS 0.760275f
C16540 DVSS.n255 VSS 0.195519f
C16541 DVSS.n256 VSS 0.195519f
C16542 DVSS.n257 VSS 0.107398f
C16543 DVSS.n258 VSS 0.157654f
C16544 DVSS.n259 VSS 0.014099f
C16545 DVSS.n260 VSS 0.250596f
C16546 DVSS.n261 VSS 0.024648f
C16547 DVSS.n262 VSS 0.053611f
C16548 DVSS.n263 VSS 0.025155f
C16549 DVSS.n264 VSS 0.053611f
C16550 DVSS.n265 VSS 0.025155f
C16551 DVSS.n266 VSS 0.053611f
C16552 DVSS.n267 VSS 0.025155f
C16553 DVSS.n268 VSS 0.053611f
C16554 DVSS.n269 VSS 0.025155f
C16555 DVSS.n270 VSS 0.053611f
C16556 DVSS.n271 VSS 0.025155f
C16557 DVSS.n272 VSS 0.014606f
C16558 DVSS.n273 VSS 0.035668f
C16559 DVSS.n274 VSS 0.034155f
C16560 DVSS.t87 VSS 5.1253f
C16561 DVSS.t185 VSS 5.1253f
C16562 DVSS.t50 VSS 5.99639f
C16563 DVSS.n275 VSS 6.33094f
C16564 DVSS.n276 VSS 0.026805f
C16565 DVSS.n277 VSS 0.046261f
C16566 DVSS.n278 VSS 0.025155f
C16567 DVSS.n279 VSS 0.025155f
C16568 DVSS.n280 VSS 0.025155f
C16569 DVSS.n281 VSS 0.053611f
C16570 DVSS.n282 VSS 0.053611f
C16571 DVSS.n283 VSS 0.053611f
C16572 DVSS.n284 VSS 0.025155f
C16573 DVSS.n285 VSS 0.025155f
C16574 DVSS.n286 VSS 0.025155f
C16575 DVSS.n287 VSS 0.053611f
C16576 DVSS.n288 VSS 0.053611f
C16577 DVSS.n289 VSS 0.053611f
C16578 DVSS.n290 VSS 0.025155f
C16579 DVSS.n291 VSS 0.025155f
C16580 DVSS.n292 VSS 0.025155f
C16581 DVSS.n293 VSS 0.053611f
C16582 DVSS.n294 VSS 0.053611f
C16583 DVSS.n295 VSS 0.053611f
C16584 DVSS.n296 VSS 0.025155f
C16585 DVSS.n297 VSS 0.025155f
C16586 DVSS.n298 VSS 0.025155f
C16587 DVSS.n299 VSS 0.053611f
C16588 DVSS.n300 VSS 0.053611f
C16589 DVSS.n301 VSS 0.053611f
C16590 DVSS.n302 VSS 0.025155f
C16591 DVSS.n303 VSS 0.025155f
C16592 DVSS.n304 VSS 0.025155f
C16593 DVSS.n305 VSS 0.053611f
C16594 DVSS.n306 VSS 0.053611f
C16595 DVSS.n307 VSS 0.094343f
C16596 DVSS.n308 VSS 0.053611f
C16597 DVSS.n309 VSS 0.023634f
C16598 DVSS.n310 VSS 0.012578f
C16599 DVSS.n311 VSS 0.097759f
C16600 DVSS.n312 VSS 0.135624f
C16601 DVSS.n313 VSS 0.195519f
C16602 DVSS.n314 VSS 0.195519f
C16603 DVSS.n315 VSS 0.195519f
C16604 DVSS.n316 VSS 0.195519f
C16605 DVSS.n317 VSS 0.195519f
C16606 DVSS.n318 VSS 0.195519f
C16607 DVSS.n319 VSS 0.195519f
C16608 DVSS.n320 VSS 0.195519f
C16609 DVSS.n321 VSS 0.195519f
C16610 DVSS.n322 VSS 0.195519f
C16611 DVSS.n323 VSS 0.195519f
C16612 DVSS.n324 VSS 0.195519f
C16613 DVSS.n325 VSS 0.195519f
C16614 DVSS.n326 VSS 0.195519f
C16615 DVSS.n327 VSS 0.195519f
C16616 DVSS.n328 VSS 0.195519f
C16617 DVSS.n329 VSS 0.195519f
C16618 DVSS.n330 VSS 0.195519f
C16619 DVSS.n331 VSS 0.195519f
C16620 DVSS.n332 VSS 0.195519f
C16621 DVSS.n333 VSS 0.195519f
C16622 DVSS.n334 VSS 0.195519f
C16623 DVSS.n335 VSS 0.195519f
C16624 DVSS.n336 VSS 0.195519f
C16625 DVSS.n337 VSS 0.195519f
C16626 DVSS.n338 VSS 0.195519f
C16627 DVSS.n339 VSS 0.195519f
C16628 DVSS.n340 VSS 0.195519f
C16629 DVSS.n341 VSS 0.195519f
C16630 DVSS.n342 VSS 0.195519f
C16631 DVSS.n343 VSS 0.195519f
C16632 DVSS.n344 VSS 0.195519f
C16633 DVSS.n345 VSS 0.195519f
C16634 DVSS.n346 VSS 0.195519f
C16635 DVSS.n347 VSS 0.195519f
C16636 DVSS.n348 VSS 0.195519f
C16637 DVSS.n349 VSS 0.195519f
C16638 DVSS.n350 VSS 0.195519f
C16639 DVSS.n351 VSS 0.195519f
C16640 DVSS.n352 VSS 0.195519f
C16641 DVSS.n353 VSS 0.195519f
C16642 DVSS.n354 VSS 0.195519f
C16643 DVSS.n355 VSS 0.195519f
C16644 DVSS.n356 VSS 0.195519f
C16645 DVSS.n357 VSS 0.195519f
C16646 DVSS.n358 VSS 0.195519f
C16647 DVSS.n359 VSS 0.162473f
C16648 DVSS.n360 VSS 0.162473f
C16649 DVSS.n361 VSS 0.152835f
C16650 DVSS.n362 VSS 2.69904f
C16651 DVSS.n363 VSS 2.83673f
C16652 DVSS.n364 VSS 4.24508f
C16653 DVSS.n365 VSS 0.097759f
C16654 DVSS.n366 VSS 0.152835f
C16655 DVSS.n367 VSS 0.162473f
C16656 DVSS.n368 VSS 0.162473f
C16657 DVSS.n369 VSS 3.38739f
C16658 DVSS.n370 VSS 3.47869f
C16659 DVSS.n371 VSS 0.162473f
C16660 DVSS.n372 VSS 0.195519f
C16661 DVSS.n373 VSS 0.097759f
C16662 DVSS.n374 VSS 0.135624f
C16663 DVSS.n375 VSS 0.195519f
C16664 DVSS.n376 VSS 0.195519f
C16665 DVSS.n377 VSS 0.195519f
C16666 DVSS.n378 VSS 0.195519f
C16667 DVSS.n379 VSS 0.195519f
C16668 DVSS.n380 VSS 0.195519f
C16669 DVSS.n381 VSS 0.195519f
C16670 DVSS.n382 VSS 0.195519f
C16671 DVSS.n383 VSS 0.195519f
C16672 DVSS.n384 VSS 0.195519f
C16673 DVSS.n385 VSS 0.195519f
C16674 DVSS.n386 VSS 0.195519f
C16675 DVSS.n387 VSS 0.195519f
C16676 DVSS.n388 VSS 0.195519f
C16677 DVSS.n389 VSS 0.195519f
C16678 DVSS.n390 VSS 0.195519f
C16679 DVSS.n391 VSS 0.195519f
C16680 DVSS.n392 VSS 0.195519f
C16681 DVSS.n393 VSS 0.195519f
C16682 DVSS.n394 VSS 0.195519f
C16683 DVSS.n395 VSS 0.195519f
C16684 DVSS.n396 VSS 0.195519f
C16685 DVSS.n397 VSS 0.195519f
C16686 DVSS.n398 VSS 0.195519f
C16687 DVSS.n399 VSS 0.195519f
C16688 DVSS.n400 VSS 0.195519f
C16689 DVSS.n401 VSS 0.195519f
C16690 DVSS.n402 VSS 0.195519f
C16691 DVSS.n403 VSS 0.195519f
C16692 DVSS.n404 VSS 0.195519f
C16693 DVSS.n405 VSS 0.195519f
C16694 DVSS.n406 VSS 0.195519f
C16695 DVSS.n407 VSS 0.195519f
C16696 DVSS.n408 VSS 0.195519f
C16697 DVSS.n409 VSS 0.195519f
C16698 DVSS.n410 VSS 0.195519f
C16699 DVSS.n411 VSS 0.195519f
C16700 DVSS.n412 VSS 0.195519f
C16701 DVSS.n413 VSS 0.195519f
C16702 DVSS.n414 VSS 0.195519f
C16703 DVSS.n415 VSS 0.195519f
C16704 DVSS.n416 VSS 0.195519f
C16705 DVSS.n417 VSS 0.195519f
C16706 DVSS.n418 VSS 0.195519f
C16707 DVSS.n419 VSS 0.195519f
C16708 DVSS.n420 VSS 0.195519f
C16709 DVSS.n421 VSS 0.195519f
C16710 DVSS.n422 VSS 0.195519f
C16711 DVSS.n423 VSS 0.195519f
C16712 DVSS.n424 VSS 0.107398f
C16713 DVSS.n425 VSS 0.097759f
C16714 DVSS.n426 VSS 0.00213f
C16715 DVSS.n427 VSS 0.009332f
C16716 DVSS.n428 VSS 0.020996f
C16717 DVSS.n429 VSS 0.030401f
C16718 DVSS.n430 VSS -0.287832f
C16719 DVSS.n431 VSS 0.053611f
C16720 DVSS.n432 VSS 0.025155f
C16721 DVSS.n433 VSS 0.025155f
C16722 DVSS.n434 VSS 0.025155f
C16723 DVSS.n435 VSS 0.053611f
C16724 DVSS.n436 VSS 0.053611f
C16725 DVSS.n437 VSS 0.053611f
C16726 DVSS.n438 VSS 0.025155f
C16727 DVSS.n439 VSS 0.025155f
C16728 DVSS.n440 VSS 0.025155f
C16729 DVSS.n441 VSS 0.053611f
C16730 DVSS.n442 VSS 0.053611f
C16731 DVSS.n443 VSS 0.053611f
C16732 DVSS.n444 VSS 0.025155f
C16733 DVSS.n445 VSS 0.025155f
C16734 DVSS.n446 VSS 0.025155f
C16735 DVSS.n447 VSS 0.053611f
C16736 DVSS.n448 VSS 0.053611f
C16737 DVSS.n449 VSS 0.053611f
C16738 DVSS.n450 VSS 0.025155f
C16739 DVSS.n451 VSS 0.025155f
C16740 DVSS.n452 VSS 0.025155f
C16741 DVSS.n453 VSS 0.053611f
C16742 DVSS.n454 VSS 0.053611f
C16743 DVSS.n455 VSS 0.053611f
C16744 DVSS.n456 VSS 0.025155f
C16745 DVSS.n457 VSS 0.025155f
C16746 DVSS.n458 VSS 0.025155f
C16747 DVSS.n459 VSS 0.053611f
C16748 DVSS.n460 VSS 0.053611f
C16749 DVSS.n461 VSS 0.531994f
C16750 DVSS.n462 VSS 0.015519f
C16751 DVSS.n463 VSS 0.00426f
C16752 DVSS.n464 VSS 0.097759f
C16753 DVSS.n465 VSS 0.157654f
C16754 DVSS.n466 VSS 0.195519f
C16755 DVSS.n467 VSS 0.195519f
C16756 DVSS.n468 VSS 0.195519f
C16757 DVSS.n469 VSS 0.195519f
C16758 DVSS.n470 VSS 0.195519f
C16759 DVSS.n471 VSS 0.195519f
C16760 DVSS.n472 VSS 0.195519f
C16761 DVSS.n473 VSS 0.195519f
C16762 DVSS.n474 VSS 0.195519f
C16763 DVSS.n475 VSS 0.195519f
C16764 DVSS.n476 VSS 0.195519f
C16765 DVSS.n477 VSS 0.195519f
C16766 DVSS.n478 VSS 0.195519f
C16767 DVSS.n479 VSS 0.195519f
C16768 DVSS.n480 VSS 0.195519f
C16769 DVSS.n481 VSS 0.195519f
C16770 DVSS.n482 VSS 0.195519f
C16771 DVSS.n483 VSS 0.195519f
C16772 DVSS.n484 VSS 0.195519f
C16773 DVSS.n485 VSS 0.195519f
C16774 DVSS.n486 VSS 0.195519f
C16775 DVSS.n487 VSS 0.195519f
C16776 DVSS.n488 VSS 0.195519f
C16777 DVSS.n489 VSS 0.195519f
C16778 DVSS.n490 VSS 0.195519f
C16779 DVSS.n491 VSS 0.195519f
C16780 DVSS.n492 VSS 0.195519f
C16781 DVSS.n493 VSS 0.195519f
C16782 DVSS.n494 VSS 0.195519f
C16783 DVSS.n495 VSS 0.195519f
C16784 DVSS.n496 VSS 0.195519f
C16785 DVSS.n497 VSS 0.109463f
C16786 DVSS.n498 VSS 0.195519f
C16787 DVSS.n499 VSS 0.195519f
C16788 DVSS.n500 VSS 0.195519f
C16789 DVSS.n501 VSS 0.195519f
C16790 DVSS.n502 VSS 0.195519f
C16791 DVSS.n503 VSS 0.195519f
C16792 DVSS.n504 VSS 0.195519f
C16793 DVSS.n505 VSS 0.183815f
C16794 DVSS.n506 VSS 0.195519f
C16795 DVSS.n507 VSS 0.195519f
C16796 DVSS.n508 VSS 0.195519f
C16797 DVSS.n509 VSS 0.125297f
C16798 DVSS.n510 VSS 0.125297f
C16799 DVSS.n511 VSS 0.235449f
C16800 DVSS.n512 VSS 0.195519f
C16801 DVSS.n513 VSS 0.195519f
C16802 DVSS.n514 VSS 0.195519f
C16803 DVSS.n515 VSS 0.195519f
C16804 DVSS.n516 VSS 0.195519f
C16805 DVSS.n517 VSS 0.195519f
C16806 DVSS.n518 VSS 0.195519f
C16807 DVSS.n519 VSS 0.195519f
C16808 DVSS.n520 VSS 0.195519f
C16809 DVSS.n521 VSS 0.195519f
C16810 DVSS.n522 VSS 0.195519f
C16811 DVSS.n523 VSS 0.195519f
C16812 DVSS.n524 VSS 0.195519f
C16813 DVSS.n525 VSS 0.195519f
C16814 DVSS.n526 VSS 0.161785f
C16815 DVSS.n527 VSS 0.131493f
C16816 DVSS.n528 VSS 0.195519f
C16817 DVSS.n529 VSS 0.195519f
C16818 DVSS.n530 VSS 0.195519f
C16819 DVSS.n531 VSS 0.195519f
C16820 DVSS.n532 VSS 0.195519f
C16821 DVSS.n533 VSS 0.195519f
C16822 DVSS.n534 VSS 0.195519f
C16823 DVSS.n535 VSS 0.195519f
C16824 DVSS.n536 VSS 0.195519f
C16825 DVSS.n537 VSS 0.195519f
C16826 DVSS.n538 VSS 0.195519f
C16827 DVSS.n539 VSS 0.195519f
C16828 DVSS.n540 VSS 0.195519f
C16829 DVSS.n541 VSS 0.195519f
C16830 DVSS.n542 VSS 0.195519f
C16831 DVSS.n543 VSS 0.195519f
C16832 DVSS.n544 VSS 0.195519f
C16833 DVSS.n545 VSS 0.195519f
C16834 DVSS.n546 VSS 0.195519f
C16835 DVSS.n547 VSS 0.195519f
C16836 DVSS.n548 VSS 0.195519f
C16837 DVSS.n549 VSS 0.195519f
C16838 DVSS.n550 VSS 0.195519f
C16839 DVSS.n551 VSS 0.195519f
C16840 DVSS.n552 VSS 0.195519f
C16841 DVSS.n553 VSS 0.195519f
C16842 DVSS.n554 VSS 0.195519f
C16843 DVSS.n555 VSS 0.195519f
C16844 DVSS.n556 VSS 0.195519f
C16845 DVSS.n557 VSS 0.195519f
C16846 DVSS.n558 VSS 0.195519f
C16847 DVSS.n559 VSS 0.195519f
C16848 DVSS.n560 VSS 0.195519f
C16849 DVSS.n561 VSS 0.195519f
C16850 DVSS.n562 VSS 0.195519f
C16851 DVSS.n563 VSS 0.195519f
C16852 DVSS.n564 VSS 0.195519f
C16853 DVSS.n565 VSS 0.195519f
C16854 DVSS.n566 VSS 0.195519f
C16855 DVSS.n567 VSS 0.195519f
C16856 DVSS.n568 VSS 0.195519f
C16857 DVSS.n569 VSS 0.195519f
C16858 DVSS.n570 VSS 0.195519f
C16859 DVSS.n571 VSS 0.195519f
C16860 DVSS.n572 VSS 0.195519f
C16861 DVSS.n573 VSS 0.167981f
C16862 DVSS.n574 VSS 0.167981f
C16863 DVSS.n575 VSS 0.167981f
C16864 DVSS.n576 VSS 0.235449f
C16865 DVSS.n577 VSS 0.373138f
C16866 DVSS.n578 VSS 0.167981f
C16867 DVSS.n579 VSS 0.195519f
C16868 DVSS.n580 VSS 0.195519f
C16869 DVSS.n581 VSS 0.195519f
C16870 DVSS.n582 VSS 0.195519f
C16871 DVSS.n583 VSS 0.195519f
C16872 DVSS.n584 VSS 0.195519f
C16873 DVSS.n585 VSS 0.195519f
C16874 DVSS.n586 VSS 0.195519f
C16875 DVSS.n587 VSS 0.195519f
C16876 DVSS.n588 VSS 0.195519f
C16877 DVSS.n589 VSS 0.195519f
C16878 DVSS.n590 VSS 0.195519f
C16879 DVSS.n591 VSS 0.195519f
C16880 DVSS.n592 VSS 0.195519f
C16881 DVSS.n593 VSS 0.195519f
C16882 DVSS.n594 VSS 0.195519f
C16883 DVSS.n595 VSS 0.195519f
C16884 DVSS.n596 VSS 0.195519f
C16885 DVSS.n597 VSS 0.195519f
C16886 DVSS.n598 VSS 0.195519f
C16887 DVSS.n599 VSS 0.195519f
C16888 DVSS.n600 VSS 0.195519f
C16889 DVSS.n601 VSS 0.195519f
C16890 DVSS.n602 VSS 0.195519f
C16891 DVSS.n603 VSS 0.195519f
C16892 DVSS.n604 VSS 0.195519f
C16893 DVSS.n605 VSS 0.195519f
C16894 DVSS.n606 VSS 0.195519f
C16895 DVSS.n607 VSS 0.195519f
C16896 DVSS.n608 VSS 0.195519f
C16897 DVSS.n609 VSS 0.167981f
C16898 DVSS.n610 VSS 0.167981f
C16899 DVSS.n611 VSS 0.373138f
C16900 DVSS.n612 VSS 0.125297f
C16901 DVSS.n613 VSS 0.195519f
C16902 DVSS.n614 VSS 0.195519f
C16903 DVSS.n615 VSS 0.195519f
C16904 DVSS.n616 VSS 0.195519f
C16905 DVSS.n617 VSS 0.195519f
C16906 DVSS.n618 VSS 0.183815f
C16907 DVSS.n619 VSS 0.143051f
C16908 DVSS.n620 VSS 0.483842f
C16909 DVSS.n621 VSS 0.427345f
C16910 DVSS.n622 VSS 0.109463f
C16911 DVSS.n623 VSS 0.195519f
C16912 DVSS.n624 VSS 0.195519f
C16913 DVSS.n625 VSS 0.195519f
C16914 DVSS.n626 VSS 0.195519f
C16915 DVSS.n627 VSS 0.195519f
C16916 DVSS.n628 VSS 0.195519f
C16917 DVSS.n629 VSS 0.195519f
C16918 DVSS.n630 VSS 0.125297f
C16919 DVSS.n631 VSS 0.125297f
C16920 DVSS.n632 VSS 0.125297f
C16921 DVSS.n633 VSS 0.235449f
C16922 DVSS.n634 VSS 0.167981f
C16923 DVSS.n635 VSS 0.167981f
C16924 DVSS.n636 VSS 0.167981f
C16925 DVSS.n637 VSS 0.195519f
C16926 DVSS.n638 VSS 0.195519f
C16927 DVSS.n639 VSS 0.195519f
C16928 DVSS.n640 VSS 0.195519f
C16929 DVSS.n641 VSS 0.195519f
C16930 DVSS.n642 VSS 0.195519f
C16931 DVSS.n643 VSS 0.195519f
C16932 DVSS.n644 VSS 0.195519f
C16933 DVSS.n645 VSS 0.195519f
C16934 DVSS.n646 VSS 0.195519f
C16935 DVSS.n647 VSS 0.195519f
C16936 DVSS.n648 VSS 0.195519f
C16937 DVSS.n649 VSS 0.195519f
C16938 DVSS.n650 VSS 0.195519f
C16939 DVSS.n651 VSS 0.195519f
C16940 DVSS.n652 VSS 0.195519f
C16941 DVSS.n653 VSS 0.195519f
C16942 DVSS.n654 VSS 0.195519f
C16943 DVSS.n655 VSS 0.195519f
C16944 DVSS.n656 VSS 0.195519f
C16945 DVSS.n657 VSS 0.195519f
C16946 DVSS.n658 VSS 0.195519f
C16947 DVSS.n659 VSS 0.195519f
C16948 DVSS.n660 VSS 0.195519f
C16949 DVSS.n661 VSS 0.195519f
C16950 DVSS.n662 VSS 0.195519f
C16951 DVSS.n663 VSS 0.195519f
C16952 DVSS.n664 VSS 0.195519f
C16953 DVSS.n665 VSS 0.195519f
C16954 DVSS.n666 VSS 0.195519f
C16955 DVSS.n667 VSS 0.195519f
C16956 DVSS.n668 VSS 0.195519f
C16957 DVSS.n669 VSS 0.195519f
C16958 DVSS.n670 VSS 0.195519f
C16959 DVSS.n671 VSS 0.195519f
C16960 DVSS.n672 VSS 0.195519f
C16961 DVSS.n673 VSS 0.195519f
C16962 DVSS.n674 VSS 0.195519f
C16963 DVSS.n675 VSS 0.195519f
C16964 DVSS.n676 VSS 0.195519f
C16965 DVSS.n677 VSS 0.195519f
C16966 DVSS.n678 VSS 0.195519f
C16967 DVSS.n679 VSS 0.195519f
C16968 DVSS.n680 VSS 0.195519f
C16969 DVSS.n681 VSS 0.195519f
C16970 DVSS.n682 VSS 0.195519f
C16971 DVSS.n683 VSS 0.195519f
C16972 DVSS.n684 VSS 0.195519f
C16973 DVSS.n685 VSS 0.195519f
C16974 DVSS.n686 VSS 0.131493f
C16975 DVSS.n687 VSS 0.427345f
C16976 DVSS.n688 VSS 0.483842f
C16977 DVSS.n689 VSS 0.143051f
C16978 DVSS.n690 VSS 0.131493f
C16979 DVSS.n691 VSS 0.195519f
C16980 DVSS.n692 VSS 0.195519f
C16981 DVSS.n693 VSS 0.195519f
C16982 DVSS.n694 VSS 0.195519f
C16983 DVSS.n695 VSS 0.195519f
C16984 DVSS.n696 VSS 0.195519f
C16985 DVSS.n697 VSS 0.195519f
C16986 DVSS.n698 VSS 0.195519f
C16987 DVSS.n699 VSS 0.195519f
C16988 DVSS.n700 VSS 0.195519f
C16989 DVSS.n701 VSS 0.195519f
C16990 DVSS.n702 VSS 0.195519f
C16991 DVSS.n703 VSS 0.195519f
C16992 DVSS.n704 VSS 0.195519f
C16993 DVSS.n705 VSS 0.195519f
C16994 DVSS.n706 VSS 0.195519f
C16995 DVSS.n707 VSS 0.195519f
C16996 DVSS.n708 VSS 0.195519f
C16997 DVSS.n709 VSS 0.195519f
C16998 DVSS.n710 VSS 0.11979f
C16999 DVSS.n711 VSS 0.195519f
C17000 DVSS.n712 VSS 0.195519f
C17001 DVSS.n713 VSS 0.195519f
C17002 DVSS.n714 VSS 0.11979f
C17003 DVSS.n715 VSS 0.373138f
C17004 DVSS.n716 VSS 0.235449f
C17005 DVSS.n717 VSS 0.11979f
C17006 DVSS.n718 VSS 0.11979f
C17007 DVSS.n719 VSS 0.11979f
C17008 DVSS.n720 VSS 0.235449f
C17009 DVSS.n721 VSS 0.173489f
C17010 DVSS.n722 VSS 0.195519f
C17011 DVSS.n723 VSS 0.195519f
C17012 DVSS.n724 VSS 0.195519f
C17013 DVSS.n725 VSS 0.195519f
C17014 DVSS.n726 VSS 0.195519f
C17015 DVSS.n727 VSS 0.195519f
C17016 DVSS.n728 VSS 0.195519f
C17017 DVSS.n729 VSS 0.195519f
C17018 DVSS.n730 VSS 0.195519f
C17019 DVSS.n731 VSS 0.195519f
C17020 DVSS.n732 VSS 0.195519f
C17021 DVSS.n733 VSS 0.195519f
C17022 DVSS.n734 VSS 0.195519f
C17023 DVSS.n735 VSS 0.195519f
C17024 DVSS.n736 VSS 0.195519f
C17025 DVSS.n737 VSS 0.195519f
C17026 DVSS.n738 VSS 0.195519f
C17027 DVSS.n739 VSS 0.195519f
C17028 DVSS.n740 VSS 0.195519f
C17029 DVSS.n741 VSS 0.195519f
C17030 DVSS.n742 VSS 0.195519f
C17031 DVSS.n743 VSS 0.195519f
C17032 DVSS.n744 VSS 0.195519f
C17033 DVSS.n745 VSS 0.195519f
C17034 DVSS.n746 VSS 0.195519f
C17035 DVSS.n747 VSS 0.195519f
C17036 DVSS.n748 VSS 0.195519f
C17037 DVSS.n749 VSS 0.195519f
C17038 DVSS.n750 VSS 0.168669f
C17039 DVSS.n751 VSS 0.124609f
C17040 DVSS.n752 VSS 0.195519f
C17041 DVSS.n753 VSS 0.140443f
C17042 DVSS.n754 VSS 0.508225f
C17043 DVSS.n755 VSS 0.022822f
C17044 DVSS.n756 VSS 0.05105f
C17045 DVSS.n757 VSS 0.022822f
C17046 DVSS.n758 VSS 0.05105f
C17047 DVSS.n759 VSS 0.022822f
C17048 DVSS.n760 VSS 0.05105f
C17049 DVSS.n761 VSS 0.022822f
C17050 DVSS.n762 VSS 0.05105f
C17051 DVSS.n763 VSS 0.022822f
C17052 DVSS.n764 VSS 0.05105f
C17053 DVSS.n765 VSS 0.008466f
C17054 DVSS.n766 VSS 0.019048f
C17055 DVSS.n767 VSS 0.028263f
C17056 DVSS.n768 VSS -0.290394f
C17057 DVSS.n769 VSS 0.022822f
C17058 DVSS.n770 VSS 0.022822f
C17059 DVSS.n771 VSS 0.022822f
C17060 DVSS.n772 VSS 0.05105f
C17061 DVSS.n773 VSS 0.05105f
C17062 DVSS.n774 VSS 0.05105f
C17063 DVSS.n775 VSS 0.022822f
C17064 DVSS.n776 VSS 0.022822f
C17065 DVSS.n777 VSS 0.022822f
C17066 DVSS.n778 VSS 0.05105f
C17067 DVSS.n779 VSS 0.05105f
C17068 DVSS.n780 VSS 0.05105f
C17069 DVSS.n781 VSS 0.022822f
C17070 DVSS.n782 VSS 0.022822f
C17071 DVSS.n783 VSS 0.022822f
C17072 DVSS.n784 VSS 0.05105f
C17073 DVSS.n785 VSS 0.05105f
C17074 DVSS.n786 VSS 0.05105f
C17075 DVSS.n787 VSS 0.022822f
C17076 DVSS.n788 VSS 0.022822f
C17077 DVSS.n789 VSS 0.022822f
C17078 DVSS.n790 VSS 0.05105f
C17079 DVSS.n791 VSS 0.05105f
C17080 DVSS.n792 VSS 0.05105f
C17081 DVSS.n793 VSS 0.022822f
C17082 DVSS.n794 VSS 0.022822f
C17083 DVSS.n795 VSS 0.022822f
C17084 DVSS.n796 VSS 0.05105f
C17085 DVSS.n797 VSS 0.05105f
C17086 DVSS.n798 VSS 0.05105f
C17087 DVSS.n799 VSS 0.022822f
C17088 DVSS.n800 VSS 0.014079f
C17089 DVSS.n801 VSS 0.097759f
C17090 DVSS.n802 VSS 0.003864f
C17091 DVSS.n803 VSS 0.231009f
C17092 DVSS.n804 VSS 0.097759f
C17093 DVSS.n805 VSS 0.071599f
C17094 DVSS.n806 VSS 0.178996f
C17095 DVSS.n807 VSS 0.195519f
C17096 DVSS.n808 VSS 0.195519f
C17097 DVSS.n809 VSS 0.195519f
C17098 DVSS.n810 VSS 0.195519f
C17099 DVSS.n811 VSS 0.195519f
C17100 DVSS.n812 VSS 0.195519f
C17101 DVSS.n813 VSS 0.195519f
C17102 DVSS.n814 VSS 0.195519f
C17103 DVSS.n815 VSS 0.195519f
C17104 DVSS.n816 VSS 0.195519f
C17105 DVSS.n817 VSS 0.195519f
C17106 DVSS.n818 VSS 0.195519f
C17107 DVSS.n819 VSS 0.195519f
C17108 DVSS.n820 VSS 0.100513f
C17109 DVSS.n821 VSS 0.195519f
C17110 DVSS.n822 VSS 0.176242f
C17111 DVSS.n823 VSS 0.117036f
C17112 DVSS.n824 VSS 0.195519f
C17113 DVSS.n825 VSS 0.195519f
C17114 DVSS.n826 VSS 0.195519f
C17115 DVSS.n827 VSS 0.195519f
C17116 DVSS.n828 VSS 0.110151f
C17117 DVSS.n829 VSS 0.097759f
C17118 DVSS.n830 VSS 0.014208f
C17119 DVSS.n831 VSS 0.014208f
C17120 DVSS.n832 VSS 0.014208f
C17121 DVSS.n833 VSS 0.014208f
C17122 DVSS.n834 VSS 0.014208f
C17123 DVSS.n835 VSS 0.014208f
C17124 DVSS.n836 VSS 0.014208f
C17125 DVSS.n837 VSS 0.014208f
C17126 DVSS.n838 VSS 0.014208f
C17127 DVSS.n839 VSS 0.014208f
C17128 DVSS.n840 VSS 0.014208f
C17129 DVSS.n841 VSS 0.014208f
C17130 DVSS.n842 VSS 0.014208f
C17131 DVSS.n843 VSS 0.014208f
C17132 DVSS.n844 VSS 0.014208f
C17133 DVSS.n845 VSS 0.014208f
C17134 DVSS.n846 VSS 0.014208f
C17135 DVSS.n847 VSS 0.014208f
C17136 DVSS.n848 VSS 0.022973f
C17137 DVSS.n849 VSS 0.045947f
C17138 DVSS.n850 VSS 0.022973f
C17139 DVSS.n851 VSS 0.045947f
C17140 DVSS.n852 VSS 0.022973f
C17141 DVSS.n853 VSS 0.045947f
C17142 DVSS.n854 VSS 0.045947f
C17143 DVSS.n855 VSS 0.425519f
C17144 DVSS.n856 VSS 0.418209f
C17145 DVSS.n857 VSS 0.091242f
C17146 DVSS.n858 VSS 0.091242f
C17147 DVSS.n859 VSS 0.091242f
C17148 DVSS.n860 VSS 0.091242f
C17149 DVSS.n861 VSS 0.091242f
C17150 DVSS.n862 VSS 0.091242f
C17151 DVSS.n863 VSS 0.091242f
C17152 DVSS.n864 VSS 0.091242f
C17153 DVSS.n865 VSS 0.091242f
C17154 DVSS.n866 VSS 0.091242f
C17155 DVSS.n867 VSS 0.091242f
C17156 DVSS.n868 VSS 0.091242f
C17157 DVSS.n869 VSS 0.091242f
C17158 DVSS.n870 VSS 0.091242f
C17159 DVSS.n871 VSS 0.091242f
C17160 DVSS.n872 VSS 0.091242f
C17161 DVSS.n873 VSS 0.091242f
C17162 DVSS.n874 VSS 0.091242f
C17163 DVSS.n875 VSS 0.091242f
C17164 DVSS.n876 VSS 0.091242f
C17165 DVSS.n877 VSS 0.091242f
C17166 DVSS.n878 VSS 0.091242f
C17167 DVSS.n879 VSS 0.091242f
C17168 DVSS.n880 VSS 0.091242f
C17169 DVSS.n881 VSS 0.091242f
C17170 DVSS.n882 VSS 0.091242f
C17171 DVSS.n883 VSS 0.091242f
C17172 DVSS.n884 VSS 0.091242f
C17173 DVSS.n885 VSS 0.091242f
C17174 DVSS.n886 VSS 0.091242f
C17175 DVSS.n887 VSS 0.091242f
C17176 DVSS.n888 VSS 0.091242f
C17177 DVSS.n889 VSS 0.091242f
C17178 DVSS.n890 VSS 0.091242f
C17179 DVSS.n891 VSS 0.091242f
C17180 DVSS.n892 VSS 0.091242f
C17181 DVSS.n893 VSS 0.091242f
C17182 DVSS.n894 VSS 0.091242f
C17183 DVSS.n895 VSS 0.091242f
C17184 DVSS.n896 VSS 0.091242f
C17185 DVSS.n897 VSS 0.091242f
C17186 DVSS.n898 VSS 0.091242f
C17187 DVSS.n899 VSS 0.091242f
C17188 DVSS.n900 VSS 0.091242f
C17189 DVSS.n901 VSS 0.091242f
C17190 DVSS.n902 VSS 0.091242f
C17191 DVSS.n903 VSS 0.091242f
C17192 DVSS.n904 VSS 0.091242f
C17193 DVSS.n905 VSS 0.091242f
C17194 DVSS.n906 VSS 0.091242f
C17195 DVSS.n907 VSS 0.091242f
C17196 DVSS.n908 VSS 0.091242f
C17197 DVSS.n909 VSS 0.091242f
C17198 DVSS.n910 VSS 0.091242f
C17199 DVSS.n911 VSS 0.091242f
C17200 DVSS.n912 VSS 0.091242f
C17201 DVSS.n913 VSS 0.091242f
C17202 DVSS.n914 VSS 0.091242f
C17203 DVSS.n915 VSS 0.091242f
C17204 DVSS.n916 VSS 0.091242f
C17205 DVSS.n917 VSS 0.091242f
C17206 DVSS.n918 VSS 0.091242f
C17207 DVSS.n919 VSS 0.091242f
C17208 DVSS.n920 VSS 0.091242f
C17209 DVSS.n921 VSS 0.091242f
C17210 DVSS.n922 VSS 0.091242f
C17211 DVSS.n923 VSS 0.091242f
C17212 DVSS.n924 VSS 0.091242f
C17213 DVSS.n925 VSS 0.091242f
C17214 DVSS.n926 VSS 0.091242f
C17215 DVSS.n927 VSS 0.091242f
C17216 DVSS.n928 VSS 0.091242f
C17217 DVSS.n929 VSS 0.091242f
C17218 DVSS.n930 VSS 0.091242f
C17219 DVSS.n931 VSS 0.091242f
C17220 DVSS.n932 VSS 0.091242f
C17221 DVSS.n933 VSS 0.091242f
C17222 DVSS.n934 VSS 0.091242f
C17223 DVSS.n935 VSS 0.091242f
C17224 DVSS.n936 VSS 0.091242f
C17225 DVSS.n937 VSS 0.091242f
C17226 DVSS.n938 VSS 0.091242f
C17227 DVSS.n939 VSS 0.091242f
C17228 DVSS.n940 VSS 0.091242f
C17229 DVSS.n941 VSS 0.091242f
C17230 DVSS.n942 VSS 0.091242f
C17231 DVSS.n943 VSS 0.091242f
C17232 DVSS.n944 VSS 0.091242f
C17233 DVSS.n945 VSS 0.091242f
C17234 DVSS.n946 VSS 0.091242f
C17235 DVSS.n947 VSS 0.091242f
C17236 DVSS.n948 VSS 0.091242f
C17237 DVSS.n949 VSS 0.564419f
C17238 DVSS.n950 VSS 0.091242f
C17239 DVSS.n951 VSS 0.045069f
C17240 DVSS.n952 VSS 0.046852f
C17241 DVSS.n953 VSS 0.156736f
C17242 DVSS.n954 VSS 0.438797f
C17243 DVSS.n955 VSS 0.443963f
C17244 DVSS.n956 VSS 2.38486f
C17245 DVSS.n957 VSS 2.04954f
C17246 DVSS.n958 VSS 3.42614f
C17247 DVSS.n959 VSS 4.34598f
C17248 DVSS.n960 VSS 6.0154f
C17249 DVSS.n961 VSS 4.153491f
C17250 DVSS.n962 VSS 1.52773f
C17251 DVSS.n963 VSS 0.828695f
C17252 DVSS.n964 VSS 0.030675f
C17253 DVSS.n965 VSS 0.012179f
C17254 DVSS.n966 VSS 0.784185f
C17255 DVSS.n967 VSS 0.012179f
C17256 DVSS.n968 VSS 0.030675f
C17257 DVSS.n969 VSS 0.012179f
C17258 DVSS.n970 VSS 0.784185f
C17259 DVSS.n971 VSS 0.012179f
C17260 DVSS.n972 VSS 0.030675f
C17261 DVSS.n973 VSS 0.012179f
C17262 DVSS.n974 VSS 0.784185f
C17263 DVSS.n975 VSS 0.012179f
C17264 DVSS.n976 VSS 0.030675f
C17265 DVSS.n977 VSS 0.012179f
C17266 DVSS.n978 VSS 0.784185f
C17267 DVSS.n979 VSS 0.012179f
C17268 DVSS.n980 VSS 0.030675f
C17269 DVSS.n981 VSS 0.012179f
C17270 DVSS.n982 VSS 0.784185f
C17271 DVSS.n983 VSS 0.012179f
C17272 DVSS.n984 VSS 0.030675f
C17273 DVSS.n985 VSS 0.012179f
C17274 DVSS.n986 VSS 0.784185f
C17275 DVSS.n987 VSS 0.012179f
C17276 DVSS.n988 VSS 0.030675f
C17277 DVSS.n989 VSS 0.012179f
C17278 DVSS.n990 VSS 0.784185f
C17279 DVSS.n991 VSS 0.012179f
C17280 DVSS.n992 VSS 0.030675f
C17281 DVSS.n993 VSS 0.012179f
C17282 DVSS.n994 VSS 0.784185f
C17283 DVSS.n995 VSS 0.012179f
C17284 DVSS.n996 VSS 0.030675f
C17285 DVSS.n997 VSS 0.012179f
C17286 DVSS.n998 VSS 0.784185f
C17287 DVSS.n999 VSS 0.012179f
C17288 DVSS.n1000 VSS 0.030675f
C17289 DVSS.n1001 VSS 0.012179f
C17290 DVSS.n1002 VSS 0.784185f
C17291 DVSS.n1003 VSS 0.012179f
C17292 DVSS.n1004 VSS 0.030675f
C17293 DVSS.n1005 VSS 0.012179f
C17294 DVSS.n1006 VSS 0.784185f
C17295 DVSS.n1007 VSS 0.012179f
C17296 DVSS.n1008 VSS 0.030675f
C17297 DVSS.n1009 VSS 0.012179f
C17298 DVSS.n1010 VSS 0.784185f
C17299 DVSS.n1011 VSS 0.012179f
C17300 DVSS.n1012 VSS 0.030675f
C17301 DVSS.n1013 VSS 0.012179f
C17302 DVSS.n1014 VSS 0.784185f
C17303 DVSS.n1015 VSS 0.012179f
C17304 DVSS.n1016 VSS 0.030675f
C17305 DVSS.n1017 VSS 0.012179f
C17306 DVSS.n1018 VSS 0.784185f
C17307 DVSS.n1019 VSS 0.012179f
C17308 DVSS.n1020 VSS 0.02313f
C17309 DVSS.n1021 VSS 0.012179f
C17310 DVSS.n1022 VSS 0.584976f
C17311 DVSS.n1023 VSS 1.57833f
C17312 DVSS.n1024 VSS 1.58068f
C17313 DVSS.n1025 VSS 0.030675f
C17314 DVSS.n1026 VSS 0.012179f
C17315 DVSS.n1027 VSS 0.784185f
C17316 DVSS.n1028 VSS 0.012179f
C17317 DVSS.n1029 VSS 0.030675f
C17318 DVSS.n1030 VSS 0.012179f
C17319 DVSS.n1031 VSS 0.784185f
C17320 DVSS.n1032 VSS 0.012179f
C17321 DVSS.n1033 VSS 0.030675f
C17322 DVSS.n1034 VSS 0.012179f
C17323 DVSS.n1035 VSS 0.784185f
C17324 DVSS.n1036 VSS 0.012179f
C17325 DVSS.n1037 VSS 0.030675f
C17326 DVSS.n1038 VSS 0.012179f
C17327 DVSS.n1039 VSS 0.784185f
C17328 DVSS.n1040 VSS 0.012179f
C17329 DVSS.n1041 VSS 0.030675f
C17330 DVSS.n1042 VSS 0.012179f
C17331 DVSS.n1043 VSS 0.784185f
C17332 DVSS.n1044 VSS 0.012179f
C17333 DVSS.n1045 VSS 0.030675f
C17334 DVSS.n1046 VSS 0.012179f
C17335 DVSS.n1047 VSS 0.784185f
C17336 DVSS.n1048 VSS 0.012179f
C17337 DVSS.n1049 VSS 0.030675f
C17338 DVSS.n1050 VSS 0.012179f
C17339 DVSS.n1051 VSS 0.784185f
C17340 DVSS.n1052 VSS 0.012179f
C17341 DVSS.n1053 VSS 0.030675f
C17342 DVSS.n1054 VSS 0.012179f
C17343 DVSS.n1055 VSS 0.784185f
C17344 DVSS.n1056 VSS 0.012179f
C17345 DVSS.n1057 VSS 0.030675f
C17346 DVSS.n1058 VSS 0.012179f
C17347 DVSS.n1059 VSS 0.784185f
C17348 DVSS.n1060 VSS 0.012179f
C17349 DVSS.n1061 VSS 0.030675f
C17350 DVSS.n1062 VSS 0.012179f
C17351 DVSS.n1063 VSS 0.784185f
C17352 DVSS.n1064 VSS 0.012179f
C17353 DVSS.n1065 VSS 0.030675f
C17354 DVSS.n1066 VSS 0.012179f
C17355 DVSS.n1067 VSS 0.784185f
C17356 DVSS.n1068 VSS 0.012179f
C17357 DVSS.n1069 VSS 0.030675f
C17358 DVSS.n1070 VSS 0.012179f
C17359 DVSS.n1071 VSS 0.784185f
C17360 DVSS.n1072 VSS 0.012179f
C17361 DVSS.n1073 VSS 0.030675f
C17362 DVSS.n1074 VSS 0.012179f
C17363 DVSS.n1075 VSS 0.784185f
C17364 DVSS.n1076 VSS 0.012179f
C17365 DVSS.n1077 VSS 0.030675f
C17366 DVSS.n1078 VSS 0.012179f
C17367 DVSS.n1079 VSS 0.686161f
C17368 DVSS.n1080 VSS 0.012179f
C17369 DVSS.n1081 VSS 0.806668f
C17370 DVSS.n1082 VSS 0.171522f
C17371 DVSS.n1083 VSS 0.091242f
C17372 DVSS.n1084 VSS 0.091242f
C17373 DVSS.n1085 VSS 0.091242f
C17374 DVSS.n1086 VSS 0.091242f
C17375 DVSS.n1087 VSS 0.091242f
C17376 DVSS.n1088 VSS 0.091242f
C17377 DVSS.n1089 VSS 0.091242f
C17378 DVSS.n1090 VSS 0.091242f
C17379 DVSS.n1091 VSS 0.091242f
C17380 DVSS.n1092 VSS 0.091242f
C17381 DVSS.n1093 VSS 0.091242f
C17382 DVSS.n1094 VSS 0.091242f
C17383 DVSS.n1095 VSS 0.091242f
C17384 DVSS.n1096 VSS 0.087708f
C17385 DVSS.n1097 VSS 0.091242f
C17386 DVSS.n1098 VSS 0.091242f
C17387 DVSS.n1099 VSS 0.091242f
C17388 DVSS.n1100 VSS 0.057822f
C17389 DVSS.n1101 VSS 0.53332f
C17390 DVSS.n1102 VSS 0.091242f
C17391 DVSS.n1103 VSS 0.091242f
C17392 DVSS.n1104 VSS 0.091242f
C17393 DVSS.n1105 VSS 0.091242f
C17394 DVSS.n1106 VSS 0.085459f
C17395 DVSS.n1107 VSS 0.091242f
C17396 DVSS.n1108 VSS 0.091242f
C17397 DVSS.n1109 VSS 0.091242f
C17398 DVSS.n1110 VSS 0.045828f
C17399 DVSS.n1111 VSS 0.045621f
C17400 DVSS.n1112 VSS 0.004046f
C17401 DVSS.n1113 VSS 0.045621f
C17402 DVSS.n1114 VSS 0.091242f
C17403 DVSS.n1115 VSS 0.091242f
C17404 DVSS.n1116 VSS 0.091242f
C17405 DVSS.n1117 VSS 0.045621f
C17406 DVSS.n1118 VSS 0.045621f
C17407 DVSS.n1119 VSS 0.045621f
C17408 DVSS.n1120 VSS 0.003383f
C17409 DVSS.n1121 VSS 0.045876f
C17410 DVSS.n1122 VSS 0.091242f
C17411 DVSS.n1123 VSS 0.091242f
C17412 DVSS.n1124 VSS 0.091242f
C17413 DVSS.n1125 VSS 0.051404f
C17414 DVSS.n1126 VSS 0.091242f
C17415 DVSS.n1127 VSS 0.091242f
C17416 DVSS.n1128 VSS 0.091242f
C17417 DVSS.n1129 VSS 0.091242f
C17418 DVSS.n1130 VSS 0.091242f
C17419 DVSS.n1131 VSS 0.091242f
C17420 DVSS.n1132 VSS 0.091242f
C17421 DVSS.n1133 VSS 0.091242f
C17422 DVSS.n1134 VSS 0.091242f
C17423 DVSS.n1135 VSS 0.091242f
C17424 DVSS.n1136 VSS 0.091242f
C17425 DVSS.n1137 VSS 0.091242f
C17426 DVSS.n1138 VSS 0.091242f
C17427 DVSS.n1139 VSS 0.091242f
C17428 DVSS.n1140 VSS 0.091242f
C17429 DVSS.n1141 VSS 0.091242f
C17430 DVSS.n1142 VSS 0.091242f
C17431 DVSS.n1143 VSS 0.091242f
C17432 DVSS.n1144 VSS 0.091242f
C17433 DVSS.n1145 VSS 0.091242f
C17434 DVSS.n1146 VSS 0.091242f
C17435 DVSS.n1147 VSS 0.091242f
C17436 DVSS.n1148 VSS 0.091242f
C17437 DVSS.n1149 VSS 0.091242f
C17438 DVSS.n1150 VSS 0.091242f
C17439 DVSS.n1151 VSS 0.091242f
C17440 DVSS.n1152 VSS 0.091242f
C17441 DVSS.n1153 VSS 0.091242f
C17442 DVSS.n1154 VSS 0.059757f
C17443 DVSS.n1155 VSS 0.014782f
C17444 DVSS.n1156 VSS 0.314661f
C17445 DVSS.n1157 VSS 0.294016f
C17446 DVSS.n1158 VSS 0.459612f
C17447 DVSS.n1159 VSS 0.32107f
C17448 DVSS.t96 VSS 0.169789f
C17449 DVSS.t97 VSS 0.00716f
C17450 DVSS.t137 VSS 0.00716f
C17451 DVSS.n1160 VSS 0.014896f
C17452 DVSS.n1161 VSS 0.006708f
C17453 DVSS.n1162 VSS 0.010442f
C17454 DVSS.n1163 VSS 0.306906f
C17455 DVSS.t81 VSS 0.169789f
C17456 DVSS.n1164 VSS 0.076172f
C17457 DVSS.n1165 VSS 0.157624f
C17458 DVSS.n1166 VSS 0.474643f
C17459 DVSS.n1167 VSS 0.950214f
C17460 DVSS.n1168 VSS 0.017012f
C17461 DVSS.t148 VSS 0.264594f
C17462 DVSS.n1169 VSS 0.706847f
C17463 DVSS.t80 VSS 0.207656f
C17464 DVSS.t200 VSS 0.318062f
C17465 DVSS.t120 VSS 0.33572f
C17466 DVSS.t192 VSS 0.245168f
C17467 DVSS.t139 VSS 0.245168f
C17468 DVSS.n1170 VSS 0.163446f
C17469 DVSS.n1171 VSS 0.069635f
C17470 DVSS.n1172 VSS 0.026127f
C17471 DVSS.n1173 VSS 0.16385f
C17472 DVSS.n1174 VSS 0.245014f
C17473 DVSS.n1175 VSS 0.195519f
C17474 DVSS.n1176 VSS 0.730195f
C17475 DVSS.n1177 VSS 0.045403f
C17476 DVSS.n1178 VSS 0.045322f
C17477 DVSS.n1179 VSS 0.024049f
C17478 DVSS.n1180 VSS 0.115659f
C17479 DVSS.n1181 VSS 0.078712f
C17480 DVSS.n1182 VSS 0.018291f
C17481 DVSS.n1183 VSS 0.018291f
C17482 DVSS.n1184 VSS 0.018291f
C17483 DVSS.n1185 VSS 0.018291f
C17484 DVSS.n1186 VSS 0.018291f
C17485 DVSS.n1187 VSS 0.018291f
C17486 DVSS.n1188 VSS 0.018291f
C17487 DVSS.n1189 VSS 0.018291f
C17488 DVSS.n1190 VSS 0.034301f
C17489 DVSS.n1191 VSS 0.022973f
C17490 DVSS.n1192 VSS 0.056274f
C17491 DVSS.n1193 VSS 3.32663f
C17492 DVSS.n1194 VSS 1.29489f
C17493 DVSS.n1195 VSS 0.020154f
C17494 DVSS.n1196 VSS 0.022186f
C17495 DVSS.n1197 VSS 0.034301f
C17496 DVSS.n1198 VSS 0.024049f
C17497 DVSS.n1199 VSS 0.034301f
C17498 DVSS.n1200 VSS 0.024049f
C17499 DVSS.n1201 VSS 0.034301f
C17500 DVSS.n1202 VSS 0.034301f
C17501 DVSS.n1203 VSS 0.02117f
C17502 DVSS.n1204 VSS 0.02117f
C17503 DVSS.n1205 VSS 0.034301f
C17504 DVSS.n1206 VSS 0.024049f
C17505 DVSS.n1207 VSS 0.034301f
C17506 DVSS.n1208 VSS 0.024049f
C17507 DVSS.n1209 VSS 0.034301f
C17508 DVSS.n1210 VSS 0.034301f
C17509 DVSS.n1211 VSS 0.022186f
C17510 DVSS.n1212 VSS 0.020154f
C17511 DVSS.n1213 VSS 0.034301f
C17512 DVSS.n1214 VSS 0.118001f
C17513 DVSS.n1215 VSS 0.186547f
C17514 DVSS.n1216 VSS 2.04288f
C17515 DVSS.n1217 VSS 1.32029f
C17516 DVSS.n1218 VSS 0.068367f
C17517 DVSS.n1219 VSS 0.257333f
C17518 DVSS.n1220 VSS 0.023334f
C17519 DVSS.n1221 VSS 0.026721f
C17520 DVSS.n1222 VSS 0.045621f
C17521 DVSS.n1223 VSS 0.045621f
C17522 DVSS.n1224 VSS 0.091242f
C17523 DVSS.n1225 VSS 0.091242f
C17524 DVSS.n1226 VSS 0.091242f
C17525 DVSS.n1227 VSS 0.091242f
C17526 DVSS.n1228 VSS 0.045621f
C17527 DVSS.n1229 VSS 0.042127f
C17528 DVSS.n1230 VSS 0.051083f
C17529 DVSS.n1231 VSS 0.045621f
C17530 DVSS.n1232 VSS 0.091242f
C17531 DVSS.n1233 VSS 0.091242f
C17532 DVSS.n1234 VSS 0.091242f
C17533 DVSS.n1235 VSS 0.091242f
C17534 DVSS.n1236 VSS 0.091242f
C17535 DVSS.n1237 VSS 0.091242f
C17536 DVSS.n1238 VSS 0.091242f
C17537 DVSS.n1239 VSS 0.045621f
C17538 DVSS.n1240 VSS 0.042127f
C17539 DVSS.n1241 VSS 0.065489f
C17540 DVSS.n1242 VSS 0.026721f
C17541 DVSS.n1243 VSS 0.045621f
C17542 DVSS.n1244 VSS 0.045621f
C17543 DVSS.n1245 VSS 0.091242f
C17544 DVSS.n1246 VSS 0.091242f
C17545 DVSS.n1247 VSS 0.091242f
C17546 DVSS.n1248 VSS 0.091242f
C17547 DVSS.n1249 VSS 0.045621f
C17548 DVSS.n1250 VSS 0.023334f
C17549 DVSS.n1251 VSS 0.051321f
C17550 DVSS.n1252 VSS 0.045803f
C17551 DVSS.n1253 VSS 0.091242f
C17552 DVSS.n1254 VSS 0.091242f
C17553 DVSS.n1255 VSS 0.091242f
C17554 DVSS.n1256 VSS 0.091242f
C17555 DVSS.n1257 VSS 0.091242f
C17556 DVSS.n1258 VSS 0.091242f
C17557 DVSS.n1259 VSS 0.091242f
C17558 DVSS.n1260 VSS 0.045621f
C17559 DVSS.n1261 VSS 0.042127f
C17560 DVSS.n1262 VSS 0.065489f
C17561 DVSS.n1263 VSS 0.026721f
C17562 DVSS.n1264 VSS 0.045621f
C17563 DVSS.n1265 VSS 0.045621f
C17564 DVSS.n1266 VSS 0.091242f
C17565 DVSS.n1267 VSS 0.091242f
C17566 DVSS.n1268 VSS 0.091242f
C17567 DVSS.n1269 VSS 0.045621f
C17568 DVSS.n1270 VSS 0.023334f
C17569 DVSS.n1271 VSS 0.251763f
C17570 DVSS.n1272 VSS 1.32067f
C17571 DVSS.n1273 VSS 4.153491f
C17572 DVSS.n1274 VSS 1.44834f
C17573 DVSS.t161 VSS 0.652381f
C17574 DVSS.n1275 VSS 0.069635f
C17575 DVSS.t162 VSS 0.01432f
C17576 DVSS.n1276 VSS 0.038163f
C17577 DVSS.n1277 VSS 0.0119f
C17578 DVSS.n1278 VSS 0.136562f
C17579 DVSS.t131 VSS 0.01432f
C17580 DVSS.t207 VSS 0.014215f
C17581 DVSS.n1279 VSS 0.026627f
C17582 DVSS.n1280 VSS 0.018226f
C17583 DVSS.t160 VSS 0.01432f
C17584 DVSS.n1281 VSS 0.028639f
C17585 DVSS.n1282 VSS 0.011953f
C17586 DVSS.t164 VSS 0.01432f
C17587 DVSS.t102 VSS 0.01432f
C17588 DVSS.n1283 VSS 0.032655f
C17589 DVSS.n1284 VSS 0.011953f
C17590 DVSS.n1285 VSS 0.035564f
C17591 DVSS.t175 VSS 0.191157f
C17592 DVSS.n1286 VSS 0.853894f
C17593 DVSS.t64 VSS 0.255618f
C17594 DVSS.n1287 VSS 0.677268f
C17595 DVSS.t168 VSS 0.01432f
C17596 DVSS.t203 VSS 0.01432f
C17597 DVSS.n1288 VSS 0.032399f
C17598 DVSS.n1289 VSS 0.020154f
C17599 DVSS.n1290 VSS 0.02385f
C17600 DVSS.n1291 VSS 0.023355f
C17601 DVSS.n1292 VSS 0.02385f
C17602 DVSS.t67 VSS 0.01432f
C17603 DVSS.t174 VSS 0.01432f
C17604 DVSS.n1293 VSS 0.032399f
C17605 DVSS.n1294 VSS 0.020154f
C17606 DVSS.n1295 VSS 0.677268f
C17607 DVSS.n1296 VSS 0.049341f
C17608 DVSS.t68 VSS 0.162261f
C17609 DVSS.t173 VSS 0.522349f
C17610 DVSS.t145 VSS 0.00716f
C17611 DVSS.t166 VSS 0.00716f
C17612 DVSS.n1297 VSS 0.014896f
C17613 DVSS.n1298 VSS 0.006708f
C17614 DVSS.n1299 VSS 0.011206f
C17615 DVSS.t144 VSS 0.271177f
C17616 DVSS.n1300 VSS -0.001185f
C17617 DVSS.t76 VSS 0.365645f
C17618 DVSS.n1301 VSS 0.074006f
C17619 DVSS.n1302 VSS 0.209286f
C17620 DVSS.t72 VSS 0.298962f
C17621 DVSS.t90 VSS 0.135588f
C17622 DVSS.n1303 VSS 0.195603f
C17623 DVSS.t181 VSS 0.143259f
C17624 DVSS.n1304 VSS 0.283557f
C17625 DVSS.n1305 VSS 0.049238f
C17626 DVSS.t71 VSS 0.01432f
C17627 DVSS.n1306 VSS 0.038163f
C17628 DVSS.n1307 VSS 0.0119f
C17629 DVSS.n1308 VSS 0.010771f
C17630 DVSS.t110 VSS 0.01432f
C17631 DVSS.t84 VSS 0.01432f
C17632 DVSS.n1309 VSS 0.032655f
C17633 DVSS.n1310 VSS 0.011953f
C17634 DVSS.n1311 VSS 0.025288f
C17635 DVSS.t112 VSS 0.01432f
C17636 DVSS.t209 VSS 0.014215f
C17637 DVSS.n1312 VSS 0.677268f
C17638 DVSS.t172 VSS 0.01432f
C17639 DVSS.t153 VSS 0.01432f
C17640 DVSS.n1313 VSS 0.032399f
C17641 DVSS.n1314 VSS 0.020154f
C17642 DVSS.n1315 VSS 0.020849f
C17643 DVSS.t156 VSS 0.205646f
C17644 DVSS.n1316 VSS 0.048972f
C17645 DVSS.n1317 VSS 0.182438f
C17646 DVSS.n1318 VSS 0.195519f
C17647 DVSS.n1319 VSS 0.195519f
C17648 DVSS.n1320 VSS 0.195519f
C17649 DVSS.n1321 VSS 0.195519f
C17650 DVSS.n1322 VSS 0.195519f
C17651 DVSS.n1323 VSS 0.195519f
C17652 DVSS.n1324 VSS 0.195519f
C17653 DVSS.n1325 VSS 0.195519f
C17654 DVSS.n1326 VSS 0.195519f
C17655 DVSS.n1327 VSS 0.195519f
C17656 DVSS.n1328 VSS 0.195519f
C17657 DVSS.n1329 VSS 0.195519f
C17658 DVSS.n1330 VSS 0.195519f
C17659 DVSS.n1331 VSS 0.195519f
C17660 DVSS.n1332 VSS 0.195519f
C17661 DVSS.n1333 VSS 0.195519f
C17662 DVSS.n1334 VSS 0.195519f
C17663 DVSS.n1335 VSS 0.195519f
C17664 DVSS.n1336 VSS 0.195519f
C17665 DVSS.n1337 VSS 0.195519f
C17666 DVSS.n1338 VSS 0.195519f
C17667 DVSS.n1339 VSS 0.195519f
C17668 DVSS.n1340 VSS 0.195519f
C17669 DVSS.n1341 VSS 0.195519f
C17670 DVSS.n1342 VSS 0.195519f
C17671 DVSS.n1343 VSS 0.195519f
C17672 DVSS.n1344 VSS 0.195519f
C17673 DVSS.n1345 VSS 0.195519f
C17674 DVSS.n1346 VSS 0.195519f
C17675 DVSS.n1347 VSS 0.195519f
C17676 DVSS.n1348 VSS 0.195519f
C17677 DVSS.n1349 VSS 0.195519f
C17678 DVSS.n1350 VSS 0.195519f
C17679 DVSS.n1351 VSS 0.195519f
C17680 DVSS.n1352 VSS 0.195519f
C17681 DVSS.n1353 VSS 0.195519f
C17682 DVSS.n1354 VSS 0.125268f
C17683 DVSS.n1355 VSS 0.195519f
C17684 DVSS.n1356 VSS 0.195519f
C17685 DVSS.n1357 VSS 0.195519f
C17686 DVSS.n1358 VSS 0.195519f
C17687 DVSS.n1359 VSS 0.195519f
C17688 DVSS.n1360 VSS 0.195519f
C17689 DVSS.n1361 VSS 0.195519f
C17690 DVSS.n1362 VSS 0.195519f
C17691 DVSS.n1363 VSS 0.195519f
C17692 DVSS.n1364 VSS 0.195519f
C17693 DVSS.n1365 VSS 0.195519f
C17694 DVSS.n1366 VSS 0.145262f
C17695 DVSS.n1367 VSS 0.693874f
C17696 DVSS.n1368 VSS 0.073369f
C17697 DVSS.n1369 VSS 0.045621f
C17698 DVSS.n1370 VSS 3.59239f
C17699 DVSS.n1371 VSS 0.091242f
C17700 DVSS.n1372 VSS 2.16852f
C17701 DVSS.n1373 VSS 0.051083f
C17702 DVSS.n1374 VSS 0.091242f
C17703 DVSS.n1375 VSS 0.091242f
C17704 DVSS.n1376 VSS 0.091242f
C17705 DVSS.n1377 VSS 0.091242f
C17706 DVSS.n1378 VSS 0.045621f
C17707 DVSS.n1379 VSS 0.018761f
C17708 DVSS.n1380 VSS 0.018761f
C17709 DVSS.n1381 VSS 0.018761f
C17710 DVSS.n1382 VSS 0.018761f
C17711 DVSS.n1383 VSS 0.018761f
C17712 DVSS.n1384 VSS 0.045621f
C17713 DVSS.n1385 VSS 0.018761f
C17714 DVSS.n1386 VSS 0.018761f
C17715 DVSS.n1387 VSS 0.018761f
C17716 DVSS.n1388 VSS 0.018761f
C17717 DVSS.n1389 VSS 0.024667f
C17718 DVSS.n1390 VSS 0.023913f
C17719 DVSS.n1391 VSS 0.091242f
C17720 DVSS.n1392 VSS 0.091242f
C17721 DVSS.n1393 VSS 0.091242f
C17722 DVSS.n1394 VSS 0.091242f
C17723 DVSS.n1395 VSS 0.091242f
C17724 DVSS.n1396 VSS 0.091242f
C17725 DVSS.n1397 VSS 0.091242f
C17726 DVSS.n1398 VSS 0.091242f
C17727 DVSS.n1399 VSS 0.091242f
C17728 DVSS.n1400 VSS 0.091242f
C17729 DVSS.n1401 VSS 0.091242f
C17730 DVSS.n1402 VSS 0.091242f
C17731 DVSS.n1403 VSS 0.091242f
C17732 DVSS.n1404 VSS 0.091242f
C17733 DVSS.n1405 VSS 0.091242f
C17734 DVSS.n1406 VSS 0.091242f
C17735 DVSS.n1407 VSS 0.091242f
C17736 DVSS.n1408 VSS 0.091242f
C17737 DVSS.n1409 VSS 0.091242f
C17738 DVSS.n1410 VSS 0.091242f
C17739 DVSS.n1411 VSS 0.091242f
C17740 DVSS.n1412 VSS 0.091242f
C17741 DVSS.n1413 VSS 0.091242f
C17742 DVSS.n1414 VSS 0.091242f
C17743 DVSS.n1415 VSS 0.091242f
C17744 DVSS.n1416 VSS 0.091242f
C17745 DVSS.n1417 VSS 0.091242f
C17746 DVSS.n1418 VSS 0.091242f
C17747 DVSS.n1419 VSS 0.091242f
C17748 DVSS.n1420 VSS 0.091242f
C17749 DVSS.n1421 VSS 0.091242f
C17750 DVSS.n1422 VSS 0.091242f
C17751 DVSS.n1423 VSS 0.091242f
C17752 DVSS.n1424 VSS 0.091242f
C17753 DVSS.n1425 VSS 0.091242f
C17754 DVSS.n1426 VSS 0.091242f
C17755 DVSS.n1427 VSS 0.01157f
C17756 DVSS.n1428 VSS 0.009121f
C17757 DVSS.n1429 VSS 0.009121f
C17758 DVSS.n1430 VSS 0.009121f
C17759 DVSS.n1431 VSS 0.045621f
C17760 DVSS.n1432 VSS 0.009121f
C17761 DVSS.n1433 VSS 0.009121f
C17762 DVSS.n1434 VSS 0.01157f
C17763 DVSS.n1435 VSS 0.011063f
C17764 DVSS.n1436 VSS 0.045621f
C17765 DVSS.n1437 VSS 0.031324f
C17766 DVSS.n1438 VSS 1.41454f
C17767 DVSS.n1439 VSS 0.690269f
C17768 DVSS.n1440 VSS -0.174112f
C17769 DVSS.n1441 VSS 0.051275f
C17770 DVSS.n1442 VSS 0.052427f
C17771 DVSS.t100 VSS 0.34564f
C17772 DVSS.n1443 VSS 0.002477f
C17773 DVSS.n1444 VSS 0.003802f
C17774 DVSS.t44 VSS 0.579651f
C17775 DVSS.n1445 VSS 0.018622f
C17776 DVSS.t95 VSS 0.380092f
C17777 DVSS.n1446 VSS 0.431805f
C17778 DVSS.n1447 VSS 0.5005f
C17779 DVSS.n1448 VSS 0.016227f
C17780 DVSS.n1449 VSS 0.024049f
C17781 DVSS.n1450 VSS 0.014219f
C17782 DVSS.n1451 VSS 0.033502f
C17783 DVSS.n1452 VSS 0.032717f
C17784 DVSS.n1453 VSS 0.271177f
C17785 DVSS.t40 VSS 0.549643f
C17786 DVSS.n1454 VSS 0.123308f
C17787 DVSS.n1455 VSS 0.031885f
C17788 DVSS.n1456 VSS 0.123308f
C17789 DVSS.n1457 VSS 0.031885f
C17790 DVSS.n1458 VSS 0.059647f
C17791 DVSS.t86 VSS 0.01432f
C17792 DVSS.t77 VSS 0.01432f
C17793 DVSS.n1459 VSS 0.032655f
C17794 DVSS.n1460 VSS 0.011123f
C17795 DVSS.t73 VSS 0.01432f
C17796 DVSS.t208 VSS 0.014215f
C17797 DVSS.n1461 VSS 0.026627f
C17798 DVSS.n1462 VSS 0.018226f
C17799 DVSS.t75 VSS 0.01432f
C17800 DVSS.n1463 VSS 0.028639f
C17801 DVSS.n1464 VSS 0.011953f
C17802 DVSS.n1465 VSS 0.023043f
C17803 DVSS.n1466 VSS 0.007635f
C17804 DVSS.n1467 VSS 0.019376f
C17805 DVSS.n1468 VSS -0.046792f
C17806 DVSS.n1469 VSS 0.031738f
C17807 DVSS.n1470 VSS 0.002529f
C17808 DVSS.t69 VSS 0.01432f
C17809 DVSS.n1471 VSS 0.038163f
C17810 DVSS.n1472 VSS 0.009513f
C17811 DVSS.n1473 VSS 0.035564f
C17812 DVSS.n1474 VSS 0.048972f
C17813 DVSS.n1475 VSS 0.078155f
C17814 DVSS.n1476 VSS 0.081457f
C17815 DVSS.n1477 VSS 0.639876f
C17816 DVSS.n1478 VSS 0.055297f
C17817 DVSS.n1479 VSS 0.33949f
C17818 DVSS.n1480 VSS 0.390526f
C17819 DVSS.n1481 VSS 0.520357f
C17820 DVSS.n1482 VSS 0.137875f
C17821 DVSS.n1483 VSS 0.017012f
C17822 DVSS.n1484 VSS -0.005939f
C17823 DVSS.n1485 VSS 0.00423f
C17824 DVSS.n1486 VSS 0.00423f
C17825 DVSS.n1487 VSS 0.068858f
C17826 DVSS.n1488 VSS 0.019182f
C17827 DVSS.n1489 VSS 0.231512f
C17828 DVSS.n1490 VSS 0.248134f
C17829 DVSS.n1491 VSS 0.734187f
C17830 DVSS.n1492 VSS 0.50453f
C17831 DVSS.n1493 VSS 0.457939f
C17832 DVSS.n1494 VSS 0.19052f
C17833 DVSS.n1495 VSS 0.052427f
C17834 DVSS.n1496 VSS 0.051275f
C17835 DVSS.n1497 VSS 0.052427f
C17836 DVSS.n1498 VSS 0.096181f
C17837 DVSS.n1499 VSS 0.052427f
C17838 DVSS.n1500 VSS 0.033284f
C17839 DVSS.n1501 VSS 0.046908f
C17840 DVSS.n1502 VSS 0.284843f
C17841 DVSS.n1503 VSS 0.017199f
C17842 DVSS.n1504 VSS 0.683543f
C17843 DVSS.t42 VSS 0.036785f
C17844 DVSS.n1505 VSS 0.070728f
C17845 DVSS.n1506 VSS 0.057728f
C17846 DVSS.t43 VSS 0.036785f
C17847 DVSS.n1507 VSS 0.182719f
C17848 DVSS.t41 VSS 0.036785f
C17849 DVSS.n1508 VSS 0.070728f
C17850 DVSS.n1509 VSS 0.072998f
C17851 DVSS.n1510 VSS 0.08164f
C17852 DVSS.n1511 VSS 0.419404f
C17853 DVSS.n1512 VSS 0.01307f
C17854 DVSS.n1513 VSS 0.057822f
C17855 DVSS.n1514 VSS 0.182934f
C17856 DVSS.n1515 VSS 0.793092f
C17857 DVSS.n1516 VSS 0.680665f
C17858 DVSS.n1517 VSS 0.418135f
C17859 DVSS.n1518 VSS 0.035618f
C17860 DVSS.n1519 VSS 0.00728f
C17861 DVSS.n1520 VSS 0.067789f
C17862 DVSS.n1521 VSS 0.091242f
C17863 DVSS.n1522 VSS 0.091242f
C17864 DVSS.n1523 VSS 0.091242f
C17865 DVSS.n1524 VSS 0.091242f
C17866 DVSS.n1525 VSS 0.091242f
C17867 DVSS.n1526 VSS 0.091242f
C17868 DVSS.n1527 VSS 0.091242f
C17869 DVSS.n1528 VSS 0.091242f
C17870 DVSS.n1529 VSS 0.091242f
C17871 DVSS.n1530 VSS 0.091242f
C17872 DVSS.n1531 VSS 0.091242f
C17873 DVSS.n1532 VSS 0.338098f
C17874 DVSS.n1533 VSS 0.091242f
C17875 DVSS.n1534 VSS 0.194467f
C17876 DVSS.n1535 VSS 0.171522f
C17877 DVSS.n1536 VSS 0.091242f
C17878 DVSS.n1537 VSS 0.091242f
C17879 DVSS.n1538 VSS 0.091242f
C17880 DVSS.n1539 VSS 0.091242f
C17881 DVSS.n1540 VSS 0.091242f
C17882 DVSS.n1541 VSS 0.091242f
C17883 DVSS.n1542 VSS 0.091242f
C17884 DVSS.n1543 VSS 0.091242f
C17885 DVSS.n1544 VSS 0.091242f
C17886 DVSS.n1545 VSS 0.091242f
C17887 DVSS.n1546 VSS 0.091242f
C17888 DVSS.n1547 VSS 0.091242f
C17889 DVSS.n1548 VSS 0.091242f
C17890 DVSS.n1549 VSS 0.091242f
C17891 DVSS.n1550 VSS 0.091242f
C17892 DVSS.n1551 VSS 0.091242f
C17893 DVSS.n1552 VSS 0.091242f
C17894 DVSS.n1553 VSS 0.091242f
C17895 DVSS.n1554 VSS 0.091242f
C17896 DVSS.n1555 VSS 0.091242f
C17897 DVSS.n1556 VSS 0.091242f
C17898 DVSS.n1557 VSS 0.091242f
C17899 DVSS.n1558 VSS 0.091242f
C17900 DVSS.n1559 VSS 0.091242f
C17901 DVSS.n1560 VSS 0.091242f
C17902 DVSS.n1561 VSS 0.091242f
C17903 DVSS.n1562 VSS 0.091242f
C17904 DVSS.n1563 VSS 0.091242f
C17905 DVSS.n1564 VSS 0.091242f
C17906 DVSS.n1565 VSS 0.091242f
C17907 DVSS.n1566 VSS 0.091242f
C17908 DVSS.n1567 VSS 0.091242f
C17909 DVSS.n1568 VSS 0.091242f
C17910 DVSS.n1569 VSS 0.091242f
C17911 DVSS.n1570 VSS 0.091242f
C17912 DVSS.n1571 VSS 0.091242f
C17913 DVSS.n1572 VSS 0.091242f
C17914 DVSS.n1573 VSS 0.059115f
C17915 DVSS.t179 VSS 0.347421f
C17916 DVSS.t154 VSS 0.270381f
C17917 DVSS.n1574 VSS 0.021765f
C17918 DVSS.t79 VSS 0.00358f
C17919 DVSS.t155 VSS 0.00358f
C17920 DVSS.n1575 VSS 0.007228f
C17921 DVSS.n1576 VSS 8.04e-19
C17922 DVSS.n1577 VSS 0.020878f
C17923 DVSS.t180 VSS 0.009228f
C17924 DVSS.n1578 VSS 0.003762f
C17925 DVSS.n1579 VSS 0.020878f
C17926 DVSS.n1580 VSS 0.018089f
C17927 DVSS.t125 VSS 0.009228f
C17928 DVSS.n1581 VSS 0.003762f
C17929 DVSS.n1582 VSS 0.020878f
C17930 DVSS.t135 VSS 0.00358f
C17931 DVSS.t123 VSS 0.00358f
C17932 DVSS.n1583 VSS 0.007228f
C17933 DVSS.n1584 VSS 8.04e-19
C17934 DVSS.n1585 VSS 0.020878f
C17935 DVSS.n1586 VSS 0.428559f
C17936 DVSS.t124 VSS 0.405941f
C17937 DVSS.t122 VSS 0.271862f
C17938 DVSS.n1587 VSS 0.157533f
C17939 DVSS.n1588 VSS 0.016769f
C17940 DVSS.t133 VSS 0.009228f
C17941 DVSS.n1589 VSS 0.003762f
C17942 DVSS.n1590 VSS 0.058151f
C17943 DVSS.n1591 VSS 0.091242f
C17944 DVSS.n1592 VSS 0.091242f
C17945 DVSS.n1593 VSS 0.091242f
C17946 DVSS.n1594 VSS 1.12525f
C17947 DVSS.n1595 VSS 0.04787f
C17948 DVSS.n1596 VSS 0.289187f
C17949 DVSS.n1597 VSS 1.96044f
C17950 DVSS.n1598 VSS 1.28426f
C17951 DVSS.n1599 VSS 0.091242f
C17952 DVSS.n1600 VSS 0.091242f
C17953 DVSS.n1601 VSS 0.091242f
C17954 DVSS.n1602 VSS 0.091242f
C17955 DVSS.n1603 VSS 0.091242f
C17956 DVSS.n1604 VSS 0.091242f
C17957 DVSS.n1605 VSS 0.059954f
C17958 DVSS.n1606 VSS 0.091242f
C17959 DVSS.n1607 VSS 0.091242f
C17960 DVSS.n1608 VSS 0.091242f
C17961 DVSS.n1609 VSS 0.058793f
C17962 DVSS.n1610 VSS 0.059954f
C17963 DVSS.n1611 VSS 0.091242f
C17964 DVSS.n1612 VSS 0.091242f
C17965 DVSS.n1613 VSS 0.091242f
C17966 DVSS.n1614 VSS 0.084495f
C17967 DVSS.n1615 VSS 0.062018f
C17968 DVSS.n1616 VSS 0.091242f
C17969 DVSS.n1617 VSS 0.091242f
C17970 DVSS.n1618 VSS 0.091242f
C17971 DVSS.n1619 VSS 0.049798f
C17972 DVSS.n1620 VSS 0.045621f
C17973 DVSS.n1621 VSS 0.091242f
C17974 DVSS.n1622 VSS 0.091242f
C17975 DVSS.n1623 VSS 0.091242f
C17976 DVSS.n1624 VSS 0.045621f
C17977 DVSS.n1625 VSS 0.045621f
C17978 DVSS.n1626 VSS 0.026069f
C17979 DVSS.n1627 VSS 0.026069f
C17980 DVSS.n1628 VSS 0.026069f
C17981 DVSS.n1629 VSS 0.026069f
C17982 DVSS.n1631 VSS 0.026069f
C17983 DVSS.n1633 VSS 0.091242f
C17984 DVSS.n1634 VSS 0.091242f
C17985 DVSS.n1635 VSS 0.091242f
C17986 DVSS.n1636 VSS 0.091242f
C17987 DVSS.n1637 VSS 0.091242f
C17988 DVSS.n1638 VSS 0.091242f
C17989 DVSS.n1639 VSS 0.091242f
C17990 DVSS.n1640 VSS 0.091242f
C17991 DVSS.n1641 VSS 0.091242f
C17992 DVSS.n1642 VSS 0.091242f
C17993 DVSS.n1643 VSS 0.085781f
C17994 DVSS.n1644 VSS 0.091242f
C17995 DVSS.n1645 VSS 0.091242f
C17996 DVSS.n1646 VSS 0.091242f
C17997 DVSS.n1647 VSS 0.062018f
C17998 DVSS.n1648 VSS 0.044886f
C17999 DVSS.n1649 VSS 0.091242f
C18000 DVSS.n1650 VSS 0.091242f
C18001 DVSS.n1651 VSS 0.091242f
C18002 DVSS.n1652 VSS 0.091242f
C18003 DVSS.n1653 VSS 0.062006f
C18004 DVSS.n1654 VSS 0.043216f
C18005 DVSS.t184 VSS 0.00358f
C18006 DVSS.t14 VSS 0.00358f
C18007 DVSS.n1655 VSS 0.007228f
C18008 DVSS.n1656 VSS 8.04e-19
C18009 DVSS.t198 VSS 0.009228f
C18010 DVSS.n1657 VSS 0.003762f
C18011 DVSS.n1658 VSS 0.010233f
C18012 DVSS.n1659 VSS 0.021765f
C18013 DVSS.t183 VSS 0.157043f
C18014 DVSS.t5 VSS 0.225194f
C18015 DVSS.n1660 VSS 0.011819f
C18016 DVSS.n1661 VSS 0.058472f
C18017 DVSS.n1662 VSS 0.059954f
C18018 DVSS.n1663 VSS 0.091242f
C18019 DVSS.n1664 VSS 0.091242f
C18020 DVSS.n1665 VSS 0.091242f
C18021 DVSS.n1666 VSS 0.091242f
C18022 DVSS.n1667 VSS 0.091242f
C18023 DVSS.n1668 VSS 0.091242f
C18024 DVSS.n1669 VSS 0.091242f
C18025 DVSS.n1670 VSS 0.091242f
C18026 DVSS.t7 VSS 0.009228f
C18027 DVSS.n1671 VSS 0.003762f
C18028 DVSS.n1672 VSS 0.009949f
C18029 DVSS.n1673 VSS 0.020878f
C18030 DVSS.n1674 VSS 0.059954f
C18031 DVSS.n1675 VSS 0.049155f
C18032 DVSS.n1676 VSS 0.091242f
C18033 DVSS.n1677 VSS 0.091242f
C18034 DVSS.n1678 VSS 0.091242f
C18035 DVSS.n1679 VSS 0.091242f
C18036 DVSS.n1680 VSS 0.091242f
C18037 DVSS.n1681 VSS 0.062006f
C18038 DVSS.n1682 VSS 0.059954f
C18039 DVSS.n1683 VSS 0.091242f
C18040 DVSS.n1684 VSS 0.091242f
C18041 DVSS.n1685 VSS 0.091242f
C18042 DVSS.n1686 VSS 0.087708f
C18043 DVSS.n1687 VSS 0.0604f
C18044 DVSS.n1688 VSS 0.047359f
C18045 DVSS.t129 VSS 0.009228f
C18046 DVSS.n1689 VSS 0.003762f
C18047 DVSS.n1690 VSS 0.016769f
C18048 DVSS.t24 VSS 0.00358f
C18049 DVSS.t127 VSS 0.00358f
C18050 DVSS.n1691 VSS 0.007228f
C18051 DVSS.n1692 VSS 8.04e-19
C18052 DVSS.n1693 VSS 0.020878f
C18053 DVSS.t23 VSS 0.140746f
C18054 DVSS.n1694 VSS 1.75893f
C18055 DVSS.n1695 VSS 0.426683f
C18056 DVSS.n1696 VSS 0.032717f
C18057 DVSS.n1697 VSS 0.012545f
C18058 DVSS.n1698 VSS 0.119454f
C18059 DVSS.n1699 VSS 0.137921f
C18060 DVSS.t157 VSS 0.253343f
C18061 DVSS.t9 VSS 0.386001f
C18062 DVSS.n1700 VSS 1.11727f
C18063 DVSS.n1701 VSS 0.281396f
C18064 DVSS.n1702 VSS 0.169688f
C18065 DVSS.n1703 VSS 0.06847f
C18066 DVSS.n1704 VSS 0.018261f
C18067 DVSS.n1705 VSS 0.056389f
C18068 DVSS.n1706 VSS 0.041956f
C18069 DVSS.t39 VSS 0.061308f
C18070 DVSS.n1707 VSS 0.078791f
C18071 DVSS.n1708 VSS 0.060846f
C18072 DVSS.n1709 VSS 0.017188f
C18073 DVSS.n1715 VSS 0.044009f
C18074 DVSS.n1717 VSS 0.113603f
C18075 DVSS.n1718 VSS 0.113603f
C18076 DVSS.n1719 VSS 0.113603f
C18077 DVSS.n1721 VSS 0.07264f
C18078 DVSS.n1722 VSS 0.113603f
C18079 DVSS.n1723 VSS 0.113603f
C18080 DVSS.n1724 VSS 0.044405f
C18081 DVSS.n1726 VSS 0.044009f
C18082 DVSS.n1727 VSS 0.044009f
C18083 DVSS.n1728 VSS 0.044009f
C18084 DVSS.n1729 VSS 0.044009f
C18085 DVSS.n1730 VSS 0.121884f
C18086 DVSS.n1731 VSS 0.033742f
C18087 DVSS.t108 VSS 0.00358f
C18088 DVSS.n1732 VSS 0.008605f
C18089 DVSS.n1733 VSS 0.00654f
C18090 DVSS.n1734 VSS 3.77592f
C18091 DVSS.n1735 VSS 0.069074f
C18092 DVSS.n1736 VSS 0.091242f
C18093 DVSS.n1737 VSS 0.091242f
C18094 DVSS.n1738 VSS 0.091242f
C18095 DVSS.n1739 VSS 0.067789f
C18096 DVSS.n1740 VSS 0.045621f
C18097 DVSS.n1741 VSS 0.091242f
C18098 DVSS.n1742 VSS 0.091242f
C18099 DVSS.n1743 VSS 0.091242f
C18100 DVSS.n1744 VSS 0.044979f
C18101 DVSS.n1745 VSS 0.045621f
C18102 DVSS.n1746 VSS 0.004452f
C18103 DVSS.n1747 VSS 0.004452f
C18104 DVSS.n1748 VSS 0.009374f
C18105 DVSS.n1749 VSS 0.006517f
C18106 DVSS.n1750 VSS 0.006517f
C18107 DVSS.n1751 VSS 0.011004f
C18108 DVSS.n1752 VSS 0.014566f
C18109 DVSS.n1753 VSS 0.006253f
C18110 DVSS.n1754 VSS 0.007267f
C18111 DVSS.n1755 VSS 0.005502f
C18112 DVSS.n1756 VSS 0.011004f
C18113 DVSS.n1757 VSS 0.005502f
C18114 DVSS.n1758 VSS 0.025702f
C18115 DVSS.n1759 VSS 0.025702f
C18116 DVSS.n1760 VSS 0.035515f
C18117 DVSS.n1761 VSS 0.025702f
C18118 DVSS.n1762 VSS 0.020562f
C18119 DVSS.n1763 VSS 0.045621f
C18120 DVSS.n1764 VSS 0.091242f
C18121 DVSS.n1765 VSS 0.091242f
C18122 DVSS.n1766 VSS 0.091242f
C18123 DVSS.n1767 VSS 0.091242f
C18124 DVSS.n1768 VSS 0.091242f
C18125 DVSS.n1769 VSS 0.045621f
C18126 DVSS.n1770 VSS 0.045621f
C18127 DVSS.n1771 VSS 0.045621f
C18128 DVSS.n1772 VSS 0.007104f
C18129 DVSS.n1773 VSS 0.005403f
C18130 DVSS.n1774 VSS 0.011004f
C18131 DVSS.n1775 VSS 0.011004f
C18132 DVSS.n1776 VSS 0.011004f
C18133 DVSS.n1777 VSS 0.005403f
C18134 DVSS.n1778 VSS 0.005653f
C18135 DVSS.n1779 VSS 0.005403f
C18136 DVSS.n1780 VSS 0.006854f
C18137 DVSS.n1781 VSS 0.011004f
C18138 DVSS.n1782 VSS 0.011004f
C18139 DVSS.n1783 VSS 0.011004f
C18140 DVSS.n1784 VSS 0.00391f
C18141 DVSS.n1786 VSS 0.019257f
C18142 DVSS.n1787 VSS 0.035983f
C18143 DVSS.n1788 VSS 0.019111f
C18144 DVSS.n1789 VSS 0.010281f
C18145 DVSS.n1790 VSS 0.091242f
C18146 DVSS.n1791 VSS 0.091242f
C18147 DVSS.n1792 VSS 0.091242f
C18148 DVSS.n1793 VSS 0.091242f
C18149 DVSS.n1794 VSS 0.091242f
C18150 DVSS.n1795 VSS 0.091242f
C18151 DVSS.n1796 VSS 0.012227f
C18152 DVSS.n1797 VSS 0.044979f
C18153 DVSS.n1798 VSS 0.035661f
C18154 DVSS.n1799 VSS 0.010602f
C18155 DVSS.n1801 VSS 0.003102f
C18156 DVSS.n1802 VSS 0.011004f
C18157 DVSS.n1803 VSS 0.170455f
C18158 DVSS.t19 VSS 2.17764f
C18159 DVSS.n1804 VSS 0.2462f
C18160 DVSS.n1805 VSS 0.005502f
C18161 DVSS.n1806 VSS 0.170484f
C18162 DVSS.n1807 VSS 0.027506f
C18163 DVSS.n1808 VSS 0.007234f
C18164 DVSS.n1809 VSS 0.044979f
C18165 DVSS.n1810 VSS 0.044979f
C18166 DVSS.n1811 VSS 0.109669f
C18167 DVSS.n1812 VSS 0.030398f
C18168 DVSS.n1813 VSS 0.077955f
C18169 DVSS.n1814 VSS 0.2462f
C18170 DVSS.n1815 VSS 0.08924f
C18171 DVSS.n1816 VSS 0.027506f
C18172 DVSS.n1817 VSS 0.005403f
C18173 DVSS.n1818 VSS 0.005502f
C18174 DVSS.n1819 VSS 0.005403f
C18175 DVSS.n1820 VSS 0.0081f
C18176 DVSS.n1821 VSS 0.016578f
C18177 DVSS.n1822 VSS 0.005783f
C18178 DVSS.n1823 VSS 0.040481f
C18179 DVSS.n1824 VSS 0.008336f
C18180 DVSS.n1825 VSS 0.008004f
C18181 DVSS.n1826 VSS 0.008054f
C18182 DVSS.n1827 VSS 0.005703f
C18183 DVSS.n1828 VSS 0.011004f
C18184 DVSS.n1829 VSS 0.006266f
C18185 DVSS.n1830 VSS 0.007104f
C18186 DVSS.n1831 VSS 0.005403f
C18187 DVSS.n1832 VSS 0.007104f
C18188 DVSS.n1833 VSS 0.01024f
C18189 DVSS.n1834 VSS 0.009323f
C18190 DVSS.n1835 VSS 0.007104f
C18191 DVSS.n1836 VSS 0.018241f
C18192 DVSS.n1837 VSS 0.024667f
C18193 DVSS.n1838 VSS 0.018241f
C18194 DVSS.n1839 VSS 0.018241f
C18195 DVSS.n1840 VSS 0.024147f
C18196 DVSS.n1841 VSS 0.019282f
C18197 DVSS.n1842 VSS 0.018241f
C18198 DVSS.n1843 VSS 0.024667f
C18199 DVSS.n1844 VSS 0.018241f
C18200 DVSS.n1845 VSS 0.024667f
C18201 DVSS.n1846 VSS 0.018241f
C18202 DVSS.n1847 VSS 0.024667f
C18203 DVSS.n1848 VSS 0.018241f
C18204 DVSS.n1849 VSS 0.018241f
C18205 DVSS.n1850 VSS 0.019282f
C18206 DVSS.n1851 VSS 0.024147f
C18207 DVSS.n1852 VSS 0.010725f
C18208 DVSS.n1853 VSS 0.019846f
C18209 DVSS.n1854 VSS 0.021957f
C18210 DVSS.n1855 VSS 0.024667f
C18211 DVSS.n1858 VSS 0.024667f
C18212 DVSS.n1859 VSS 0.010178f
C18213 DVSS.n1860 VSS 0.261647f
C18214 DVSS.n1861 VSS -0.078269f
C18215 DVSS.n1862 VSS 0.849155f
C18216 DVSS.n1863 VSS 0.215798f
C18217 DVSS.n1864 VSS 0.006839f
C18218 DVSS.n1865 VSS 0.232574f
C18219 DVSS.n1866 VSS 0.112316f
C18220 DVSS.n1867 VSS 0.418309f
C18221 DVSS.n1868 VSS 0.054446f
C18222 DVSS.n1869 VSS 0.007821f
C18223 DVSS.n1870 VSS 0.035983f
C18224 DVSS.n1871 VSS 0.091242f
C18225 DVSS.n1872 VSS 0.091242f
C18226 DVSS.n1873 VSS 0.010281f
C18227 DVSS.n1874 VSS 0.044979f
C18228 DVSS.n1875 VSS 0.007821f
C18229 DVSS.n1876 VSS 0.015642f
C18230 DVSS.n1877 VSS 0.044979f
C18231 DVSS.n1878 VSS 0.016358f
C18232 DVSS.n1879 VSS 0.101959f
C18233 DVSS.n1880 VSS 0.109669f
C18234 DVSS.n1882 VSS 0.044979f
C18235 DVSS.n1883 VSS 0.029067f
C18236 DVSS.n1884 VSS 0.020562f
C18237 DVSS.n1885 VSS 0.091242f
C18238 DVSS.n1886 VSS 0.091242f
C18239 DVSS.n1887 VSS 0.091242f
C18240 DVSS.n1888 VSS 0.045621f
C18241 DVSS.n1889 VSS 0.008537f
C18242 DVSS.n1890 VSS 0.285584f
C18243 DVSS.n1891 VSS 0.045621f
C18244 DVSS.n1892 VSS 0.045621f
C18245 DVSS.n1893 VSS 0.045621f
C18246 DVSS.n1894 VSS 0.091242f
C18247 DVSS.n1895 VSS 0.091242f
C18248 DVSS.n1896 VSS 0.091242f
C18249 DVSS.n1897 VSS 0.091242f
C18250 DVSS.n1898 VSS 0.045621f
C18251 DVSS.n1899 VSS 0.045621f
C18252 DVSS.n1900 VSS 0.379506f
C18253 DVSS.n1901 VSS 0.045621f
C18254 DVSS.n1902 VSS 0.045621f
C18255 DVSS.n1903 VSS 0.091242f
C18256 DVSS.n1904 VSS 0.091242f
C18257 DVSS.n1905 VSS 0.091242f
C18258 DVSS.n1906 VSS 0.091242f
C18259 DVSS.n1907 VSS 0.091242f
C18260 DVSS.n1908 VSS 0.020562f
C18261 DVSS.n1909 VSS 0.044979f
C18262 DVSS.n1912 VSS 0.029067f
C18263 DVSS.n1913 VSS 0.044979f
C18264 DVSS.n1914 VSS 0.030398f
C18265 DVSS.n1915 VSS 0.143005f
C18266 DVSS.n1916 VSS 0.188043f
C18267 DVSS.n1917 VSS 0.16584f
C18268 DVSS.n1918 VSS 0.087925f
C18269 DVSS.n1919 VSS 0.099719f
C18270 DVSS.n1920 VSS 0.014357f
C18271 DVSS.n1921 VSS 0.19818f
C18272 DVSS.n1922 VSS 1.16483f
C18273 DVSS.n1923 VSS 0.170484f
C18274 DVSS.n1924 VSS 0.288962f
C18275 DVSS.n1925 VSS 0.032146f
C18276 DVSS.n1926 VSS 0.045621f
C18277 DVSS.n1927 VSS 0.091242f
C18278 DVSS.n1928 VSS 0.091242f
C18279 DVSS.n1929 VSS 0.091242f
C18280 DVSS.n1930 VSS 0.045621f
C18281 DVSS.n1931 VSS 0.045621f
C18282 DVSS.n1932 VSS 0.045621f
C18283 DVSS.n1933 VSS 0.007104f
C18284 DVSS.n1934 VSS 0.005653f
C18285 DVSS.n1935 VSS 0.011004f
C18286 DVSS.n1936 VSS 0.005403f
C18287 DVSS.n1937 VSS 0.005403f
C18288 DVSS.n1938 VSS 0.007104f
C18289 DVSS.n1939 VSS 0.011004f
C18290 DVSS.n1940 VSS 0.011004f
C18291 DVSS.n1941 VSS 0.011004f
C18292 DVSS.n1942 VSS 0.005403f
C18293 DVSS.n1943 VSS 0.007267f
C18294 DVSS.n1944 VSS 0.007267f
C18295 DVSS.n1945 VSS 0.005403f
C18296 DVSS.n1946 VSS 0.005502f
C18297 DVSS.n1947 VSS 0.011004f
C18298 DVSS.n1948 VSS 0.005502f
C18299 DVSS.n1949 VSS 0.011004f
C18300 DVSS.n1950 VSS 0.011004f
C18301 DVSS.n1951 VSS 0.005753f
C18302 DVSS.n1952 VSS 0.045621f
C18303 DVSS.n1953 VSS 0.045621f
C18304 DVSS.n1954 VSS 0.091242f
C18305 DVSS.n1955 VSS 0.091242f
C18306 DVSS.n1956 VSS 0.091242f
C18307 DVSS.n1957 VSS 0.091242f
C18308 DVSS.n1958 VSS 0.025059f
C18309 DVSS.n1959 VSS 0.022721f
C18310 DVSS.n1960 VSS 0.021204f
C18311 DVSS.n1961 VSS 0.021204f
C18312 DVSS.n1962 VSS 0.045621f
C18313 DVSS.n1963 VSS 0.045621f
C18314 DVSS.n1964 VSS 0.029067f
C18315 DVSS.n1965 VSS 0.035515f
C18316 DVSS.n1966 VSS 0.025059f
C18317 DVSS.n1967 VSS 0.091242f
C18318 DVSS.n1968 VSS 0.091242f
C18319 DVSS.n1969 VSS 0.091242f
C18320 DVSS.n1970 VSS 0.091242f
C18321 DVSS.n1971 VSS 0.091242f
C18322 DVSS.n1972 VSS 0.091242f
C18323 DVSS.n1973 VSS 0.025059f
C18324 DVSS.n1975 VSS 0.044979f
C18325 DVSS.n1977 VSS 0.044979f
C18326 DVSS.n1979 VSS 0.029067f
C18327 DVSS.n1980 VSS 0.044979f
C18328 DVSS.n1981 VSS 0.021204f
C18329 DVSS.n1982 VSS 0.009518f
C18330 DVSS.n1983 VSS 0.045621f
C18331 DVSS.n1984 VSS 0.045621f
C18332 DVSS.n1985 VSS 0.045621f
C18333 DVSS.n1986 VSS 0.091242f
C18334 DVSS.n1987 VSS 0.091242f
C18335 DVSS.n1988 VSS 0.091242f
C18336 DVSS.n1989 VSS 0.091242f
C18337 DVSS.n1990 VSS 0.091242f
C18338 DVSS.n1991 VSS 0.091242f
C18339 DVSS.n1992 VSS 0.091242f
C18340 DVSS.n1993 VSS 0.091242f
C18341 DVSS.n1994 VSS 0.091242f
C18342 DVSS.n1995 VSS 0.091242f
C18343 DVSS.n1996 VSS 0.091242f
C18344 DVSS.n1997 VSS 0.091242f
C18345 DVSS.n1998 VSS 0.091242f
C18346 DVSS.n1999 VSS 0.091242f
C18347 DVSS.n2000 VSS 0.091242f
C18348 DVSS.n2001 VSS 0.091242f
C18349 DVSS.n2002 VSS 0.091242f
C18350 DVSS.n2003 VSS 0.091242f
C18351 DVSS.n2004 VSS 0.091242f
C18352 DVSS.n2005 VSS 0.091242f
C18353 DVSS.n2006 VSS 0.091242f
C18354 DVSS.n2007 VSS 0.091242f
C18355 DVSS.n2008 VSS 0.091242f
C18356 DVSS.n2009 VSS 0.091242f
C18357 DVSS.n2010 VSS 0.091242f
C18358 DVSS.n2011 VSS 0.091242f
C18359 DVSS.n2012 VSS 0.091242f
C18360 DVSS.n2013 VSS 0.091242f
C18361 DVSS.n2014 VSS 0.091242f
C18362 DVSS.n2015 VSS 0.091242f
C18363 DVSS.n2016 VSS 0.091242f
C18364 DVSS.n2017 VSS 0.091242f
C18365 DVSS.n2018 VSS 0.091242f
C18366 DVSS.n2019 VSS 0.091242f
C18367 DVSS.n2020 VSS 0.082246f
C18368 DVSS.n2021 VSS 0.046906f
C18369 DVSS.n2022 VSS 0.120102f
C18370 DVSS.n2023 VSS 0.439756f
C18371 DVSS.n2024 VSS 0.082246f
C18372 DVSS.n2025 VSS 0.091242f
C18373 DVSS.n2026 VSS 0.091242f
C18374 DVSS.n2027 VSS 0.091242f
C18375 DVSS.n2028 VSS 0.091242f
C18376 DVSS.n2029 VSS 0.091242f
C18377 DVSS.n2030 VSS 0.091242f
C18378 DVSS.n2031 VSS 0.091242f
C18379 DVSS.n2032 VSS 0.091242f
C18380 DVSS.n2033 VSS 0.091242f
C18381 DVSS.n2034 VSS 0.091242f
C18382 DVSS.n2035 VSS 0.091242f
C18383 DVSS.n2036 VSS 0.091242f
C18384 DVSS.n2037 VSS 0.091242f
C18385 DVSS.n2038 VSS 0.091242f
C18386 DVSS.n2039 VSS 0.091242f
C18387 DVSS.n2040 VSS 0.091242f
C18388 DVSS.n2041 VSS 0.091242f
C18389 DVSS.n2042 VSS 0.091242f
C18390 DVSS.n2043 VSS 0.091242f
C18391 DVSS.n2044 VSS 0.091242f
C18392 DVSS.n2045 VSS 0.091242f
C18393 DVSS.n2046 VSS 0.091242f
C18394 DVSS.n2047 VSS 0.091242f
C18395 DVSS.n2048 VSS 0.091242f
C18396 DVSS.n2049 VSS 0.091242f
C18397 DVSS.n2050 VSS 0.091242f
C18398 DVSS.n2051 VSS 0.091242f
C18399 DVSS.n2052 VSS 0.091242f
C18400 DVSS.n2053 VSS 0.091242f
C18401 DVSS.n2054 VSS 0.091242f
C18402 DVSS.n2055 VSS 0.091242f
C18403 DVSS.n2056 VSS 0.091242f
C18404 DVSS.n2057 VSS 0.091242f
C18405 DVSS.n2058 VSS 0.091242f
C18406 DVSS.n2059 VSS 0.091242f
C18407 DVSS.n2060 VSS 0.091242f
C18408 DVSS.n2061 VSS 0.091242f
C18409 DVSS.n2062 VSS 0.091242f
C18410 DVSS.n2063 VSS 0.091242f
C18411 DVSS.n2064 VSS 0.091242f
C18412 DVSS.n2065 VSS 0.091242f
C18413 DVSS.n2066 VSS 0.091242f
C18414 DVSS.n2067 VSS 0.091242f
C18415 DVSS.n2068 VSS 0.091242f
C18416 DVSS.n2069 VSS 0.091242f
C18417 DVSS.n2070 VSS 0.091242f
C18418 DVSS.n2071 VSS 0.091242f
C18419 DVSS.n2072 VSS 0.091242f
C18420 DVSS.n2073 VSS 0.091242f
C18421 DVSS.n2074 VSS 0.091242f
C18422 DVSS.n2075 VSS 0.091242f
C18423 DVSS.n2076 VSS 0.091242f
C18424 DVSS.n2077 VSS 0.091242f
C18425 DVSS.n2078 VSS 0.091242f
C18426 DVSS.n2079 VSS 0.091242f
C18427 DVSS.n2080 VSS 0.091242f
C18428 DVSS.n2081 VSS 0.084817f
C18429 DVSS.n2082 VSS 0.091242f
C18430 DVSS.n2083 VSS 0.091242f
C18431 DVSS.n2084 VSS 0.045621f
C18432 DVSS.n2085 VSS 0.045621f
C18433 DVSS.n2086 VSS 0.005502f
C18434 DVSS.n2087 VSS 0.039838f
C18435 DVSS.n2088 VSS 0.006425f
C18436 DVSS.n2089 VSS 0.009374f
C18437 DVSS.n2090 VSS 0.005403f
C18438 DVSS.n2091 VSS 0.011004f
C18439 DVSS.n2092 VSS 0.006754f
C18440 DVSS.n2093 VSS 0.005403f
C18441 DVSS.n2094 VSS 0.007104f
C18442 DVSS.n2095 VSS 0.011004f
C18443 DVSS.n2096 VSS 0.012125f
C18444 DVSS.n2097 VSS 0.006003f
C18445 DVSS.n2098 VSS 0.009154f
C18446 DVSS.n2099 VSS 0.010138f
C18447 DVSS.n2100 VSS 0.006266f
C18448 DVSS.n2101 VSS 0.005502f
C18449 DVSS.n2102 VSS 0.009323f
C18450 DVSS.n2103 VSS 0.01024f
C18451 DVSS.n2104 VSS 0.007234f
C18452 DVSS.n2105 VSS 0.005502f
C18453 DVSS.n2106 VSS 0.007234f
C18454 DVSS.n2107 VSS 0.005502f
C18455 DVSS.n2108 VSS 0.005808f
C18456 DVSS.n2109 VSS 0.011004f
C18457 DVSS.n2110 VSS 0.0081f
C18458 DVSS.n2111 VSS 0.0081f
C18459 DVSS.n2112 VSS 0.003617f
C18460 DVSS.n2113 VSS 0.008559f
C18461 DVSS.n2114 VSS 0.003617f
C18462 DVSS.n2115 VSS 0.004738f
C18463 DVSS.n2116 VSS 0.006425f
C18464 DVSS.n2117 VSS 0.045621f
C18465 DVSS.n2118 VSS 0.091242f
C18466 DVSS.n2119 VSS 0.091242f
C18467 DVSS.n2120 VSS 0.091242f
C18468 DVSS.n2121 VSS 0.091242f
C18469 DVSS.n2122 VSS 0.091242f
C18470 DVSS.n2123 VSS 0.045621f
C18471 DVSS.n2124 VSS 0.045621f
C18472 DVSS.n2125 VSS 0.005403f
C18473 DVSS.n2126 VSS 0.007104f
C18474 DVSS.n2127 VSS 0.011004f
C18475 DVSS.n2128 VSS 0.011004f
C18476 DVSS.n2129 VSS 0.006954f
C18477 DVSS.n2130 VSS 0.015756f
C18478 DVSS.n2131 VSS 0.006253f
C18479 DVSS.n2132 VSS 0.011004f
C18480 DVSS.n2133 VSS 0.011004f
C18481 DVSS.n2134 VSS 0.011004f
C18482 DVSS.n2135 VSS 0.006854f
C18483 DVSS.n2136 VSS 0.005403f
C18484 DVSS.n2137 VSS 0.045621f
C18485 DVSS.n2138 VSS 0.045621f
C18486 DVSS.n2139 VSS 0.091242f
C18487 DVSS.n2140 VSS 0.091242f
C18488 DVSS.n2141 VSS 0.091242f
C18489 DVSS.n2142 VSS 0.091242f
C18490 DVSS.n2143 VSS 0.091242f
C18491 DVSS.n2144 VSS 0.035661f
C18492 DVSS.n2145 VSS 0.044979f
C18493 DVSS.n2146 VSS 0.019111f
C18494 DVSS.n2147 VSS 0.007821f
C18495 DVSS.n2148 VSS 0.015642f
C18496 DVSS.n2149 VSS 0.007821f
C18497 DVSS.n2150 VSS 0.016358f
C18498 DVSS.n2151 VSS 0.101959f
C18499 DVSS.n2152 VSS 0.077955f
C18500 DVSS.n2153 VSS 0.08924f
C18501 DVSS.n2154 VSS 0.143056f
C18502 DVSS.n2155 VSS 0.188043f
C18503 DVSS.n2156 VSS 0.165582f
C18504 DVSS.n2157 VSS 0.087925f
C18505 DVSS.n2158 VSS 0.009374f
C18506 DVSS.n2159 VSS 0.014357f
C18507 DVSS.n2160 VSS 0.19818f
C18508 DVSS.n2161 VSS 1.16483f
C18509 DVSS.n2162 VSS 0.170455f
C18510 DVSS.n2163 VSS 0.289691f
C18511 DVSS.n2164 VSS 0.02751f
C18512 DVSS.n2165 VSS 0.019257f
C18513 DVSS.n2166 VSS 0.00391f
C18514 DVSS.n2167 VSS 0.006498f
C18515 DVSS.n2168 VSS 0.00391f
C18516 DVSS.n2169 VSS 0.005122f
C18517 DVSS.n2170 VSS 0.010602f
C18518 DVSS.n2171 VSS 0.046264f
C18519 DVSS.n2172 VSS 0.091242f
C18520 DVSS.n2173 VSS 0.091242f
C18521 DVSS.n2174 VSS 0.091242f
C18522 DVSS.n2175 VSS 0.091242f
C18523 DVSS.n2176 VSS 0.091242f
C18524 DVSS.n2177 VSS 0.0906f
C18525 DVSS.n2178 VSS 0.005122f
C18526 DVSS.n2179 VSS 0.045621f
C18527 DVSS.n2180 VSS 0.012227f
C18528 DVSS.n2181 VSS 0.00391f
C18529 DVSS.n2182 VSS 0.006348f
C18530 DVSS.n2183 VSS 0.003052f
C18531 DVSS.n2184 VSS 0.011004f
C18532 DVSS.n2185 VSS 0.011004f
C18533 DVSS.n2186 VSS 0.007104f
C18534 DVSS.n2187 VSS 0.005403f
C18535 DVSS.n2188 VSS 0.045621f
C18536 DVSS.n2189 VSS 0.045621f
C18537 DVSS.n2190 VSS 0.091242f
C18538 DVSS.n2191 VSS 0.091242f
C18539 DVSS.n2192 VSS 0.091242f
C18540 DVSS.n2193 VSS 0.091242f
C18541 DVSS.n2194 VSS 0.091242f
C18542 DVSS.n2195 VSS 0.045621f
C18543 DVSS.n2196 VSS 0.009518f
C18544 DVSS.n2197 VSS 0.045621f
C18545 DVSS.n2198 VSS 0.022721f
C18546 DVSS.n2199 VSS 0.007267f
C18547 DVSS.n2200 VSS 0.015756f
C18548 DVSS.n2201 VSS 0.006153f
C18549 DVSS.n2202 VSS 0.011004f
C18550 DVSS.n2203 VSS 0.011004f
C18551 DVSS.n2204 VSS 0.005502f
C18552 DVSS.n2205 VSS 0.011004f
C18553 DVSS.n2206 VSS 0.005502f
C18554 DVSS.n2207 VSS 0.011004f
C18555 DVSS.n2208 VSS 0.012125f
C18556 DVSS.n2209 VSS 0.007104f
C18557 DVSS.n2210 VSS 0.006504f
C18558 DVSS.n2211 VSS 0.045621f
C18559 DVSS.n2212 VSS 0.005783f
C18560 DVSS.n2213 VSS 0.091242f
C18561 DVSS.n2214 VSS 0.091242f
C18562 DVSS.n2215 VSS 0.091242f
C18563 DVSS.n2216 VSS 0.091242f
C18564 DVSS.n2217 VSS 0.091242f
C18565 DVSS.n2218 VSS 0.086102f
C18566 DVSS.n2219 VSS 0.091242f
C18567 DVSS.n2220 VSS 0.091242f
C18568 DVSS.n2221 VSS 0.091242f
C18569 DVSS.n2222 VSS 0.091242f
C18570 DVSS.n2223 VSS 0.091242f
C18571 DVSS.n2224 VSS 2.33046f
C18572 DVSS.n2225 VSS 0.091242f
C18573 DVSS.n2226 VSS 0.30967f
C18574 DVSS.n2227 VSS 0.074857f
C18575 DVSS.n2228 VSS 2.05044f
C18576 DVSS.n2229 VSS 0.024405f
C18577 DVSS.t107 VSS 0.111457f
C18578 DVSS.n2230 VSS 0.315346f
C18579 DVSS.n2231 VSS 0.047698f
C18580 DVSS.n2232 VSS 0.032881f
C18581 DVSS.n2233 VSS 0.303522f
C18582 DVSS.n2234 VSS 0.40817f
C18583 DVSS.n2235 VSS 1.19026f
C18584 DVSS.n2236 VSS 0.016769f
C18585 DVSS.n2237 VSS 0.200105f
C18586 DVSS.n2238 VSS 0.170595f
C18587 DVSS.t104 VSS 0.009546f
C18588 DVSS.t106 VSS 0.009546f
C18589 DVSS.n2239 VSS 0.02024f
C18590 DVSS.n2240 VSS 0.006738f
C18591 DVSS.t146 VSS 0.20223f
C18592 DVSS.n2241 VSS 0.207323f
C18593 DVSS.n2242 VSS 0.029237f
C18594 DVSS.n2243 VSS 0.209693f
C18595 DVSS.n2244 VSS 0.31779f
C18596 DVSS.n2245 VSS 0.022905f
C18597 DVSS.t105 VSS 0.220749f
C18598 DVSS.n2246 VSS 0.316694f
C18599 DVSS.n2247 VSS 0.036157f
C18600 DVSS.n2248 VSS 0.054201f
C18601 DVSS.n2249 VSS 0.280751f
C18602 DVSS.n2250 VSS 0.017496f
C18603 DVSS.n2251 VSS 0.030214f
C18604 DVSS.n2252 VSS 0.423272f
C18605 DVSS.n2253 VSS 2.06599f
C18606 DVSS.n2254 VSS 0.906259f
C18607 DVSS.t8 VSS 0.253343f
C18608 DVSS.t15 VSS 0.253343f
C18609 DVSS.n2255 VSS 0.287418f
C18610 DVSS.n2256 VSS 0.02291f
C18611 DVSS.n2257 VSS 0.012545f
C18612 DVSS.n2258 VSS 0.040306f
C18613 DVSS.n2259 VSS 0.036157f
C18614 DVSS.n2260 VSS 0.287418f
C18615 DVSS.t196 VSS 0.220749f
C18616 DVSS.t63 VSS 0.180748f
C18617 DVSS.t197 VSS 0.180748f
C18618 DVSS.t18 VSS 0.226675f
C18619 DVSS.n2261 VSS 0.016769f
C18620 DVSS.n2262 VSS 0.160844f
C18621 DVSS.t62 VSS 0.220749f
C18622 DVSS.n2263 VSS 0.388381f
C18623 DVSS.n2264 VSS 0.667402f
C18624 DVSS.n2265 VSS 0.091242f
C18625 DVSS.n2266 VSS 0.091242f
C18626 DVSS.n2267 VSS 0.089957f
C18627 DVSS.n2268 VSS 0.091242f
C18628 DVSS.n2269 VSS 0.01767f
C18629 DVSS.n2275 VSS 0.045621f
C18630 DVSS.n2276 VSS 0.008073f
C18631 DVSS.n2277 VSS 0.013127f
C18632 DVSS.n2278 VSS 0.036625f
C18633 DVSS.n2279 VSS 0.01767f
C18634 DVSS.n2280 VSS 0.026069f
C18635 DVSS.n2281 VSS 0.026069f
C18636 DVSS.n2282 VSS 0.091242f
C18637 DVSS.n2283 VSS 0.054617f
C18638 DVSS.n2284 VSS 0.091242f
C18639 DVSS.n2285 VSS 0.091242f
C18640 DVSS.n2286 VSS 0.091242f
C18641 DVSS.n2287 VSS 0.091242f
C18642 DVSS.n2288 VSS 0.091242f
C18643 DVSS.n2289 VSS 0.091242f
C18644 DVSS.n2290 VSS 0.091242f
C18645 DVSS.n2291 VSS 0.091242f
C18646 DVSS.n2292 VSS 0.091242f
C18647 DVSS.n2293 VSS 0.091242f
C18648 DVSS.n2294 VSS 0.091242f
C18649 DVSS.n2295 VSS 0.091242f
C18650 DVSS.n2296 VSS 0.091242f
C18651 DVSS.n2297 VSS 0.091242f
C18652 DVSS.n2298 VSS 0.091242f
C18653 DVSS.n2299 VSS 0.091242f
C18654 DVSS.n2300 VSS 0.091242f
C18655 DVSS.n2301 VSS 0.091242f
C18656 DVSS.n2302 VSS 0.091242f
C18657 DVSS.n2303 VSS 0.091242f
C18658 DVSS.n2304 VSS 0.091242f
C18659 DVSS.n2305 VSS 0.091242f
C18660 DVSS.n2306 VSS 0.091242f
C18661 DVSS.n2307 VSS 0.091242f
C18662 DVSS.n2308 VSS 0.091242f
C18663 DVSS.n2309 VSS 0.091242f
C18664 DVSS.n2310 VSS 0.091242f
C18665 DVSS.n2311 VSS 0.091242f
C18666 DVSS.n2312 VSS 0.091242f
C18667 DVSS.n2313 VSS 0.091242f
C18668 DVSS.n2314 VSS 0.091242f
C18669 DVSS.n2315 VSS 0.091242f
C18670 DVSS.n2316 VSS 0.091242f
C18671 DVSS.n2317 VSS 0.091242f
C18672 DVSS.n2318 VSS 0.091242f
C18673 DVSS.n2319 VSS 0.091242f
C18674 DVSS.n2320 VSS 0.091242f
C18675 DVSS.n2321 VSS 0.091242f
C18676 DVSS.n2322 VSS 0.091242f
C18677 DVSS.n2323 VSS 0.091242f
C18678 DVSS.n2324 VSS 0.091242f
C18679 DVSS.n2325 VSS 0.091242f
C18680 DVSS.n2326 VSS 0.091242f
C18681 DVSS.n2327 VSS 0.091242f
C18682 DVSS.n2328 VSS 0.091242f
C18683 DVSS.n2329 VSS 0.091242f
C18684 DVSS.n2330 VSS 0.091242f
C18685 DVSS.n2331 VSS 0.091242f
C18686 DVSS.n2332 VSS 0.091242f
C18687 DVSS.n2333 VSS 0.091242f
C18688 DVSS.n2334 VSS 0.091242f
C18689 DVSS.n2335 VSS 0.091242f
C18690 DVSS.n2336 VSS 0.091242f
C18691 DVSS.n2337 VSS 0.091242f
C18692 DVSS.n2338 VSS 0.091242f
C18693 DVSS.n2339 VSS 0.091242f
C18694 DVSS.n2340 VSS 0.091242f
C18695 DVSS.n2341 VSS 0.091242f
C18696 DVSS.n2342 VSS 0.091242f
C18697 DVSS.n2343 VSS 0.091242f
C18698 DVSS.n2344 VSS 0.091242f
C18699 DVSS.n2345 VSS 0.091242f
C18700 DVSS.n2346 VSS 0.091242f
C18701 DVSS.n2347 VSS 0.091242f
C18702 DVSS.n2348 VSS 0.091242f
C18703 DVSS.n2349 VSS 0.091242f
C18704 DVSS.n2350 VSS 0.091242f
C18705 DVSS.n2351 VSS 0.091242f
C18706 DVSS.n2352 VSS 0.091242f
C18707 DVSS.n2353 VSS 0.091242f
C18708 DVSS.n2354 VSS 0.091242f
C18709 DVSS.n2355 VSS 0.091242f
C18710 DVSS.n2356 VSS 0.091242f
C18711 DVSS.n2357 VSS 0.091242f
C18712 DVSS.n2358 VSS 0.091242f
C18713 DVSS.n2359 VSS 0.091242f
C18714 DVSS.n2360 VSS 0.091242f
C18715 DVSS.n2361 VSS 0.091242f
C18716 DVSS.n2362 VSS 0.091242f
C18717 DVSS.n2363 VSS 0.091242f
C18718 DVSS.n2364 VSS 0.091242f
C18719 DVSS.n2365 VSS 0.091242f
C18720 DVSS.n2366 VSS 0.091242f
C18721 DVSS.n2367 VSS 0.091242f
C18722 DVSS.n2368 VSS 0.091242f
C18723 DVSS.n2369 VSS 0.091242f
C18724 DVSS.n2370 VSS 0.091242f
C18725 DVSS.n2371 VSS 0.091242f
C18726 DVSS.n2372 VSS 0.091242f
C18727 DVSS.n2373 VSS 0.091242f
C18728 DVSS.n2374 VSS 0.091242f
C18729 DVSS.n2375 VSS 0.091242f
C18730 DVSS.n2376 VSS 0.091242f
C18731 DVSS.n2377 VSS 0.091242f
C18732 DVSS.n2378 VSS 0.091242f
C18733 DVSS.n2379 VSS 0.091242f
C18734 DVSS.n2380 VSS 0.091242f
C18735 DVSS.n2381 VSS 0.091242f
C18736 DVSS.n2382 VSS 0.091242f
C18737 DVSS.n2383 VSS 0.091242f
C18738 DVSS.n2384 VSS 0.091242f
C18739 DVSS.n2385 VSS 0.091242f
C18740 DVSS.n2386 VSS 0.091242f
C18741 DVSS.n2387 VSS 0.091242f
C18742 DVSS.n2388 VSS 0.091242f
C18743 DVSS.n2389 VSS 0.091242f
C18744 DVSS.n2390 VSS 0.054295f
C18745 DVSS.n2391 VSS 0.091242f
C18746 DVSS.n2392 VSS 0.045621f
C18747 DVSS.n2393 VSS 0.082246f
C18748 DVSS.n2394 VSS 0.082246f
C18749 DVSS.n2395 VSS 0.010281f
C18750 DVSS.n2396 VSS 0.197025f
C18751 DVSS.n2397 VSS 0.091242f
C18752 DVSS.n2398 VSS 0.091242f
C18753 DVSS.n2399 VSS 0.174165f
C18754 DVSS.n2400 VSS 0.340567f
C18755 DVSS.n2401 VSS 0.089957f
C18756 DVSS.n2402 VSS 0.091242f
C18757 DVSS.n2403 VSS 0.082568f
C18758 DVSS.n2406 VSS 0.026069f
C18759 DVSS.n2408 VSS 0.015605f
C18760 DVSS.n2410 VSS 0.026069f
C18761 DVSS.n2412 VSS 0.026069f
C18762 DVSS.n2414 VSS 0.026069f
C18763 DVSS.n2416 VSS 0.026069f
C18764 DVSS.n2418 VSS 0.022948f
C18765 DVSS.n2419 VSS 0.045621f
C18766 DVSS.n2420 VSS 1.21497f
C18767 DVSS.n2421 VSS 0.054295f
C18768 DVSS.n2422 VSS 0.026069f
C18769 DVSS.n2423 VSS 0.026069f
C18770 DVSS.n2424 VSS 0.026069f
C18771 DVSS.n2425 VSS 0.026069f
C18772 DVSS.n2426 VSS 0.091242f
C18773 DVSS.n2427 VSS 0.091242f
C18774 DVSS.n2428 VSS 0.091242f
C18775 DVSS.n2429 VSS 0.091242f
C18776 DVSS.n2430 VSS 0.091242f
C18777 DVSS.n2431 VSS 0.091242f
C18778 DVSS.n2432 VSS 0.091242f
C18779 DVSS.n2433 VSS 0.091242f
C18780 DVSS.n2434 VSS 0.091242f
C18781 DVSS.n2435 VSS 0.091242f
C18782 DVSS.n2436 VSS 0.091242f
C18783 DVSS.n2437 VSS 0.091242f
C18784 DVSS.n2438 VSS 0.091242f
C18785 DVSS.n2439 VSS 0.091242f
C18786 DVSS.n2440 VSS 0.091242f
C18787 DVSS.n2441 VSS 0.091242f
C18788 DVSS.n2442 VSS 0.091242f
C18789 DVSS.n2443 VSS 0.091242f
C18790 DVSS.n2444 VSS 0.091242f
C18791 DVSS.n2445 VSS 0.091242f
C18792 DVSS.n2446 VSS 0.091242f
C18793 DVSS.n2447 VSS 0.091242f
C18794 DVSS.n2448 VSS 0.091242f
C18795 DVSS.n2449 VSS 0.091242f
C18796 DVSS.n2450 VSS 0.091242f
C18797 DVSS.n2451 VSS 0.091242f
C18798 DVSS.n2452 VSS 0.091242f
C18799 DVSS.n2453 VSS 0.091242f
C18800 DVSS.n2454 VSS 0.091242f
C18801 DVSS.n2455 VSS 0.091242f
C18802 DVSS.n2456 VSS 0.091242f
C18803 DVSS.n2457 VSS 0.091242f
C18804 DVSS.n2458 VSS 0.091242f
C18805 DVSS.n2459 VSS 0.091242f
C18806 DVSS.n2460 VSS 0.091242f
C18807 DVSS.n2461 VSS 0.091242f
C18808 DVSS.n2462 VSS 0.091242f
C18809 DVSS.n2463 VSS 0.091242f
C18810 DVSS.n2464 VSS 0.091242f
C18811 DVSS.n2465 VSS 0.091242f
C18812 DVSS.n2466 VSS 0.091242f
C18813 DVSS.n2467 VSS 0.091242f
C18814 DVSS.n2468 VSS 0.091242f
C18815 DVSS.n2469 VSS 0.091242f
C18816 DVSS.n2470 VSS 0.091242f
C18817 DVSS.n2471 VSS 0.091242f
C18818 DVSS.n2472 VSS 0.091242f
C18819 DVSS.n2473 VSS 0.091242f
C18820 DVSS.n2474 VSS 0.091242f
C18821 DVSS.n2475 VSS 0.091242f
C18822 DVSS.n2476 VSS 0.091242f
C18823 DVSS.n2477 VSS 0.091242f
C18824 DVSS.n2478 VSS 0.091242f
C18825 DVSS.n2479 VSS 0.091242f
C18826 DVSS.n2480 VSS 0.091242f
C18827 DVSS.n2481 VSS 0.091242f
C18828 DVSS.n2482 VSS 0.091242f
C18829 DVSS.n2483 VSS 0.091242f
C18830 DVSS.n2484 VSS 0.091242f
C18831 DVSS.n2485 VSS 0.091242f
C18832 DVSS.n2486 VSS 0.091242f
C18833 DVSS.n2487 VSS 0.091242f
C18834 DVSS.n2488 VSS 0.091242f
C18835 DVSS.n2489 VSS 0.091242f
C18836 DVSS.n2490 VSS 0.091242f
C18837 DVSS.n2491 VSS 0.091242f
C18838 DVSS.n2492 VSS 0.091242f
C18839 DVSS.n2493 VSS 0.091242f
C18840 DVSS.n2494 VSS 0.091242f
C18841 DVSS.n2495 VSS 0.091242f
C18842 DVSS.n2496 VSS 0.091242f
C18843 DVSS.n2497 VSS 0.091242f
C18844 DVSS.n2498 VSS 0.091242f
C18845 DVSS.n2499 VSS 0.091242f
C18846 DVSS.n2500 VSS 0.091242f
C18847 DVSS.n2501 VSS 0.091242f
C18848 DVSS.n2502 VSS 0.091242f
C18849 DVSS.n2503 VSS 0.091242f
C18850 DVSS.n2504 VSS 0.091242f
C18851 DVSS.n2505 VSS 0.091242f
C18852 DVSS.n2506 VSS 0.091242f
C18853 DVSS.n2507 VSS 0.091242f
C18854 DVSS.n2508 VSS 0.091242f
C18855 DVSS.n2509 VSS 0.091242f
C18856 DVSS.n2510 VSS 0.091242f
C18857 DVSS.n2511 VSS 0.091242f
C18858 DVSS.n2512 VSS 0.091242f
C18859 DVSS.n2513 VSS 0.091242f
C18860 DVSS.n2514 VSS 0.091242f
C18861 DVSS.n2515 VSS 0.091242f
C18862 DVSS.n2516 VSS 0.091242f
C18863 DVSS.n2517 VSS 0.091242f
C18864 DVSS.n2518 VSS 0.091242f
C18865 DVSS.n2519 VSS 0.091242f
C18866 DVSS.n2520 VSS 0.091242f
C18867 DVSS.n2521 VSS 0.091242f
C18868 DVSS.n2522 VSS 0.091242f
C18869 DVSS.n2523 VSS 0.091242f
C18870 DVSS.n2524 VSS 0.091242f
C18871 DVSS.n2525 VSS 0.091242f
C18872 DVSS.n2526 VSS 0.091242f
C18873 DVSS.n2527 VSS 0.091242f
C18874 DVSS.n2528 VSS 0.091242f
C18875 DVSS.n2529 VSS 0.091242f
C18876 DVSS.n2530 VSS 0.091242f
C18877 DVSS.n2531 VSS 0.091242f
C18878 DVSS.n2532 VSS 0.091242f
C18879 DVSS.n2533 VSS 0.091242f
C18880 DVSS.n2534 VSS 0.091242f
C18881 DVSS.n2535 VSS 0.091242f
C18882 DVSS.n2536 VSS 0.091242f
C18883 DVSS.n2537 VSS 0.091242f
C18884 DVSS.n2538 VSS 0.091242f
C18885 DVSS.n2539 VSS 0.091242f
C18886 DVSS.n2540 VSS 0.091242f
C18887 DVSS.n2541 VSS 0.091242f
C18888 DVSS.n2542 VSS 0.091242f
C18889 DVSS.n2543 VSS 0.091242f
C18890 DVSS.n2544 VSS 0.091242f
C18891 DVSS.n2545 VSS 0.091242f
C18892 DVSS.n2546 VSS 0.091242f
C18893 DVSS.n2547 VSS 0.091242f
C18894 DVSS.n2548 VSS 0.091242f
C18895 DVSS.n2549 VSS 0.091242f
C18896 DVSS.n2550 VSS 0.091242f
C18897 DVSS.n2551 VSS 0.091242f
C18898 DVSS.n2552 VSS 0.091242f
C18899 DVSS.n2553 VSS 0.091242f
C18900 DVSS.n2554 VSS 0.091242f
C18901 DVSS.n2555 VSS 0.091242f
C18902 DVSS.n2556 VSS 0.091242f
C18903 DVSS.n2557 VSS 0.091242f
C18904 DVSS.n2558 VSS 0.091242f
C18905 DVSS.n2559 VSS 0.091242f
C18906 DVSS.n2560 VSS 0.091242f
C18907 DVSS.n2561 VSS 0.091242f
C18908 DVSS.n2562 VSS 0.091242f
C18909 DVSS.n2563 VSS 0.091242f
C18910 DVSS.n2564 VSS 0.091242f
C18911 DVSS.n2565 VSS 0.091242f
C18912 DVSS.n2566 VSS 0.091242f
C18913 DVSS.n2567 VSS 0.091242f
C18914 DVSS.n2568 VSS 0.091242f
C18915 DVSS.n2569 VSS 0.091242f
C18916 DVSS.n2570 VSS 0.091242f
C18917 DVSS.n2571 VSS 0.091242f
C18918 DVSS.n2572 VSS 0.091242f
C18919 DVSS.n2573 VSS 0.091242f
C18920 DVSS.n2574 VSS 0.091242f
C18921 DVSS.n2575 VSS 0.091242f
C18922 DVSS.n2576 VSS 0.091242f
C18923 DVSS.n2577 VSS 0.091242f
C18924 DVSS.n2578 VSS 0.091242f
C18925 DVSS.n2579 VSS 0.091242f
C18926 DVSS.n2580 VSS 0.091242f
C18927 DVSS.n2581 VSS 0.091242f
C18928 DVSS.n2582 VSS 0.091242f
C18929 DVSS.n2583 VSS 0.091242f
C18930 DVSS.n2584 VSS 0.091242f
C18931 DVSS.n2585 VSS 0.091242f
C18932 DVSS.n2586 VSS 0.091242f
C18933 DVSS.n2587 VSS 0.091242f
C18934 DVSS.n2588 VSS 0.091242f
C18935 DVSS.n2589 VSS 0.091242f
C18936 DVSS.n2590 VSS 0.091242f
C18937 DVSS.n2591 VSS 0.091242f
C18938 DVSS.n2592 VSS 0.091242f
C18939 DVSS.n2593 VSS 0.091242f
C18940 DVSS.n2594 VSS 0.091242f
C18941 DVSS.n2595 VSS 0.091242f
C18942 DVSS.n2596 VSS 0.091242f
C18943 DVSS.n2597 VSS 0.091242f
C18944 DVSS.n2598 VSS 0.091242f
C18945 DVSS.n2599 VSS 0.091242f
C18946 DVSS.n2600 VSS 0.091242f
C18947 DVSS.n2601 VSS 0.091242f
C18948 DVSS.n2602 VSS 0.091242f
C18949 DVSS.n2603 VSS 0.091242f
C18950 DVSS.n2604 VSS 0.091242f
C18951 DVSS.n2605 VSS 0.091242f
C18952 DVSS.n2606 VSS 0.091242f
C18953 DVSS.n2607 VSS 0.091242f
C18954 DVSS.n2608 VSS 0.091242f
C18955 DVSS.n2609 VSS 0.091242f
C18956 DVSS.n2610 VSS 0.091242f
C18957 DVSS.n2611 VSS 0.091242f
C18958 DVSS.n2612 VSS 0.091242f
C18959 DVSS.n2613 VSS 0.091242f
C18960 DVSS.n2614 VSS 0.091242f
C18961 DVSS.n2615 VSS 0.091242f
C18962 DVSS.n2616 VSS 0.091242f
C18963 DVSS.n2617 VSS 0.091242f
C18964 DVSS.n2618 VSS 0.091242f
C18965 DVSS.n2619 VSS 0.091242f
C18966 DVSS.n2620 VSS 0.091242f
C18967 DVSS.n2621 VSS 0.091242f
C18968 DVSS.n2622 VSS 0.091242f
C18969 DVSS.n2623 VSS 0.091242f
C18970 DVSS.n2624 VSS 0.091242f
C18971 DVSS.n2625 VSS 0.091242f
C18972 DVSS.n2626 VSS 0.091242f
C18973 DVSS.n2627 VSS 0.091242f
C18974 DVSS.n2628 VSS 0.091242f
C18975 DVSS.n2629 VSS 0.091242f
C18976 DVSS.n2630 VSS 0.091242f
C18977 DVSS.n2631 VSS 0.091242f
C18978 DVSS.n2632 VSS 0.054617f
C18979 DVSS.n2633 VSS 0.046906f
C18980 DVSS.n2634 VSS 0.091242f
C18981 DVSS.n2635 VSS 0.082246f
C18982 DVSS.n2636 VSS 0.045621f
C18983 DVSS.n2637 VSS 0.026069f
C18984 DVSS.n2638 VSS 0.026069f
C18985 DVSS.n2639 VSS 0.026069f
C18986 DVSS.n2643 VSS 0.036625f
C18987 DVSS.n2645 VSS 0.026069f
C18988 DVSS.n2646 VSS 0.045621f
C18989 DVSS.n2647 VSS 1.21754f
C18990 DVSS.n2648 VSS 0.045621f
C18991 DVSS.n2649 VSS 0.082568f
C18992 DVSS.n2650 VSS 0.091242f
C18993 DVSS.n2651 VSS 0.091242f
C18994 DVSS.n2652 VSS 0.340567f
C18995 DVSS.n2653 VSS 0.174165f
C18996 DVSS.n2654 VSS 0.19702f
C18997 DVSS.n2655 VSS 0.808965f
C18998 DVSS.n2656 VSS 1.02507f
C18999 DVSS.n2657 VSS 2.30086f
C19000 DVSS.n2658 VSS 1.18039f
C19001 DVSS.n2659 VSS 0.078417f
C19002 DVSS.n2660 VSS 0.436019f
C19003 DVSS.n2661 VSS 0.611621f
C19004 DVSS.n2662 VSS 0.020032f
C19005 DVSS.n2663 VSS 0.023106f
C19006 DVSS.n2664 VSS 0.01107f
C19007 DVSS.n2665 VSS 0.011731f
C19008 DVSS.n2666 VSS 0.041646f
C19009 DVSS.n2667 VSS 0.041646f
C19010 DVSS.n2668 VSS 0.010905f
C19011 DVSS.n2669 VSS 0.010244f
C19012 DVSS.n2670 VSS 0.012485f
C19013 DVSS.n2671 VSS 0.023106f
C19014 DVSS.n2672 VSS 0.011731f
C19015 DVSS.n2673 VSS 0.041646f
C19016 DVSS.n2674 VSS 0.010244f
C19017 DVSS.n2675 VSS 0.041646f
C19018 DVSS.n2676 VSS 0.083291f
C19019 DVSS.n2677 VSS 0.083291f
C19020 DVSS.n2678 VSS 0.083291f
C19021 DVSS.n2679 VSS 0.083291f
C19022 DVSS.n2680 VSS 0.041646f
C19023 DVSS.n2681 VSS 0.010244f
C19024 DVSS.n2682 VSS 0.011731f
C19025 DVSS.n2683 VSS 0.019845f
C19026 DVSS.n2684 VSS 0.011731f
C19027 DVSS.n2685 VSS 0.041646f
C19028 DVSS.n2686 VSS 0.011731f
C19029 DVSS.n2687 VSS 0.010244f
C19030 DVSS.n2688 VSS 0.013044f
C19031 DVSS.n2689 VSS 0.010244f
C19032 DVSS.n2690 VSS 0.041646f
C19033 DVSS.n2691 VSS 0.010244f
C19034 DVSS.t45 VSS 0.061308f
C19035 DVSS.n2692 VSS 0.021288f
C19036 DVSS.n2693 VSS 0.011731f
C19037 DVSS.n2694 VSS 0.041646f
C19038 DVSS.n2695 VSS 0.011731f
C19039 DVSS.n2696 VSS 0.010244f
C19040 DVSS.n2697 VSS 0.041646f
C19041 DVSS.n2698 VSS 0.083291f
C19042 DVSS.n2699 VSS 0.083291f
C19043 DVSS.n2700 VSS 0.083291f
C19044 DVSS.n2701 VSS 0.041646f
C19045 DVSS.n2702 VSS 0.010244f
C19046 DVSS.n2703 VSS 0.011235f
C19047 DVSS.n2704 VSS 0.023106f
C19048 DVSS.n2705 VSS 0.011731f
C19049 DVSS.n2706 VSS 0.041646f
C19050 DVSS.n2707 VSS 0.011731f
C19051 DVSS.n2708 VSS 0.010244f
C19052 DVSS.n2709 VSS 0.019264f
C19053 DVSS.n2710 VSS 0.010244f
C19054 DVSS.n2711 VSS 0.041646f
C19055 DVSS.n2712 VSS 0.010244f
C19056 DVSS.n2713 VSS 0.023106f
C19057 DVSS.n2714 VSS 0.011731f
C19058 DVSS.n2715 VSS 0.041646f
C19059 DVSS.n2716 VSS 0.010244f
C19060 DVSS.n2717 VSS 0.041646f
C19061 DVSS.n2718 VSS 0.083291f
C19062 DVSS.n2719 VSS 0.083291f
C19063 DVSS.n2720 VSS 0.083291f
C19064 DVSS.n2721 VSS 0.041646f
C19065 DVSS.n2722 VSS 0.010244f
C19066 DVSS.n2723 VSS 0.010244f
C19067 DVSS.n2724 VSS 0.010244f
C19068 DVSS.t38 VSS 0.061308f
C19069 DVSS.n2725 VSS 0.021288f
C19070 DVSS.n2726 VSS 0.011731f
C19071 DVSS.n2727 VSS 0.041646f
C19072 DVSS.n2728 VSS 0.010244f
C19073 DVSS.n2729 VSS 0.041646f
C19074 DVSS.n2730 VSS 0.041646f
C19075 DVSS.n2731 VSS 0.083291f
C19076 DVSS.n2732 VSS 0.083291f
C19077 DVSS.n2733 VSS 0.083291f
C19078 DVSS.n2734 VSS 0.041646f
C19079 DVSS.n2735 VSS 0.010244f
C19080 DVSS.n2736 VSS 0.010244f
C19081 DVSS.n2737 VSS 0.023106f
C19082 DVSS.n2738 VSS 0.011731f
C19083 DVSS.n2739 VSS 0.041646f
C19084 DVSS.n2740 VSS 0.011731f
C19085 DVSS.n2741 VSS 0.010244f
C19086 DVSS.n2742 VSS 0.014721f
C19087 DVSS.n2743 VSS 0.010244f
C19088 DVSS.n2744 VSS 0.041646f
C19089 DVSS.n2745 VSS 0.010244f
C19090 DVSS.n2746 VSS 0.019264f
C19091 DVSS.n2747 VSS 0.010244f
C19092 DVSS.n2748 VSS 0.023106f
C19093 DVSS.n2749 VSS 0.011731f
C19094 DVSS.n2750 VSS 0.041646f
C19095 DVSS.n2751 VSS 0.010244f
C19096 DVSS.n2752 VSS 0.041646f
C19097 DVSS.n2753 VSS 0.083291f
C19098 DVSS.n2754 VSS 0.083291f
C19099 DVSS.n2755 VSS 0.083291f
C19100 DVSS.n2756 VSS 0.041646f
C19101 DVSS.n2757 VSS 0.010244f
C19102 DVSS.n2758 VSS 0.010244f
C19103 DVSS.n2759 VSS 0.01528f
C19104 DVSS.n2760 VSS 0.011731f
C19105 DVSS.n2761 VSS 0.041646f
C19106 DVSS.n2762 VSS 0.011731f
C19107 DVSS.n2763 VSS 0.010244f
C19108 DVSS.n2764 VSS 0.023106f
C19109 DVSS.n2765 VSS 0.020488f
C19110 DVSS.n2766 VSS 0.041646f
C19111 DVSS.n2767 VSS 0.020488f
C19112 DVSS.n2768 VSS 0.023106f
C19113 DVSS.n2769 VSS 0.011731f
C19114 DVSS.n2770 VSS 0.041646f
C19115 DVSS.n2771 VSS 0.010244f
C19116 DVSS.n2772 VSS 0.041646f
C19117 DVSS.n2773 VSS 0.083291f
C19118 DVSS.n2774 VSS 0.083291f
C19119 DVSS.n2775 VSS 0.083291f
C19120 DVSS.n2776 VSS 0.041646f
C19121 DVSS.n2777 VSS 0.010244f
C19122 DVSS.n2778 VSS 0.010244f
C19123 DVSS.n2779 VSS 0.019264f
C19124 DVSS.n2780 VSS 0.011731f
C19125 DVSS.n2781 VSS 0.041646f
C19126 DVSS.n2782 VSS 0.011731f
C19127 DVSS.n2783 VSS 0.010244f
C19128 DVSS.n2784 VSS 0.023106f
C19129 DVSS.n2785 VSS 0.010244f
C19130 DVSS.n2786 VSS 0.041646f
C19131 DVSS.n2787 VSS 0.010244f
C19132 DVSS.n2788 VSS 0.023106f
C19133 DVSS.n2789 VSS 0.019636f
C19134 DVSS.n2790 VSS 0.041646f
C19135 DVSS.n2791 VSS 0.010244f
C19136 DVSS.n2792 VSS 0.041646f
C19137 DVSS.n2793 VSS 0.218779f
C19138 DVSS.n2794 VSS 0.011646f
C19139 DVSS.t35 VSS 0.061308f
C19140 DVSS.n2795 VSS 0.162297f
C19141 DVSS.n2796 VSS 0.097235f
C19142 DVSS.n2797 VSS 0.162297f
C19143 DVSS.n2798 VSS 0.011566f
C19144 DVSS.n2799 VSS 0.010409f
C19145 DVSS.n2800 VSS 0.023106f
C19146 DVSS.n2801 VSS 0.011646f
C19147 DVSS.n2802 VSS 0.019636f
C19148 DVSS.n2803 VSS 0.7102f
C19149 DVSS.n2804 VSS 0.996095f
C19150 DVSS.n2805 VSS 0.805693f
C19151 DVSS.n2806 VSS 0.083291f
C19152 DVSS.n2807 VSS 0.083291f
C19153 DVSS.n2808 VSS 0.083291f
C19154 DVSS.n2809 VSS 0.083291f
C19155 DVSS.n2810 VSS 0.083291f
C19156 DVSS.n2811 VSS 0.041646f
C19157 DVSS.n2812 VSS 0.041646f
C19158 DVSS.n2813 VSS 0.010244f
C19159 DVSS.n2814 VSS 0.010409f
C19160 DVSS.n2815 VSS 0.011566f
C19161 DVSS.n2816 VSS 0.023106f
C19162 DVSS.n2817 VSS 0.01882f
C19163 DVSS.n2818 VSS 0.023106f
C19164 DVSS.n2819 VSS 0.011731f
C19165 DVSS.n2820 VSS 0.010244f
C19166 DVSS.n2821 VSS 0.041646f
C19167 DVSS.n2822 VSS 0.010244f
C19168 DVSS.n2823 VSS 0.011731f
C19169 DVSS.n2824 VSS 0.023106f
C19170 DVSS.n2825 VSS 0.01882f
C19171 DVSS.n2826 VSS 0.019264f
C19172 DVSS.n2827 VSS 0.011731f
C19173 DVSS.n2828 VSS 0.023106f
C19174 DVSS.n2829 VSS 0.011731f
C19175 DVSS.n2830 VSS 0.023106f
C19176 DVSS.n2831 VSS 0.011731f
C19177 DVSS.n2832 VSS 0.023106f
C19178 DVSS.n2833 VSS 0.015839f
C19179 DVSS.n2834 VSS 0.011731f
C19180 DVSS.n2835 VSS 0.010244f
C19181 DVSS.n2836 VSS 0.041646f
C19182 DVSS.n2837 VSS 0.041646f
C19183 DVSS.n2838 VSS 0.010244f
C19184 DVSS.n2839 VSS 0.011731f
C19185 DVSS.n2840 VSS 0.015839f
C19186 DVSS.n2841 VSS 0.023106f
C19187 DVSS.n2842 VSS 0.011731f
C19188 DVSS.n2843 VSS 0.010244f
C19189 DVSS.n2844 VSS 0.041646f
C19190 DVSS.n2845 VSS 0.041646f
C19191 DVSS.n2846 VSS 0.083291f
C19192 DVSS.n2847 VSS 0.083291f
C19193 DVSS.n2848 VSS 0.083291f
C19194 DVSS.n2849 VSS 0.083291f
C19195 DVSS.n2850 VSS 0.083291f
C19196 DVSS.n2851 VSS 0.083291f
C19197 DVSS.n2852 VSS 0.083291f
C19198 DVSS.n2853 VSS 0.083291f
C19199 DVSS.n2854 VSS 0.083291f
C19200 DVSS.n2855 VSS 0.041646f
C19201 DVSS.n2856 VSS 0.041646f
C19202 DVSS.n2857 VSS 0.010244f
C19203 DVSS.n2858 VSS 0.011731f
C19204 DVSS.n2859 VSS 0.023106f
C19205 DVSS.n2860 VSS 0.023106f
C19206 DVSS.t48 VSS 0.061308f
C19207 DVSS.n2861 VSS 0.021288f
C19208 DVSS.n2862 VSS 0.019379f
C19209 DVSS.n2863 VSS 0.011731f
C19210 DVSS.n2864 VSS 0.010244f
C19211 DVSS.n2865 VSS 0.041646f
C19212 DVSS.n2866 VSS 0.010244f
C19213 DVSS.n2867 VSS 0.011731f
C19214 DVSS.n2868 VSS 0.019379f
C19215 DVSS.n2869 VSS 0.021288f
C19216 DVSS.n2870 VSS 0.01528f
C19217 DVSS.n2871 VSS 0.019264f
C19218 DVSS.n2872 VSS 0.019938f
C19219 DVSS.n2873 VSS 0.010409f
C19220 DVSS.n2874 VSS 0.011566f
C19221 DVSS.n2875 VSS 0.010244f
C19222 DVSS.n2876 VSS 0.011731f
C19223 DVSS.n2877 VSS 0.023106f
C19224 DVSS.n2878 VSS 0.011731f
C19225 DVSS.n2879 VSS 0.023106f
C19226 DVSS.n2880 VSS 0.011731f
C19227 DVSS.n2881 VSS 0.022081f
C19228 DVSS.n2882 VSS 0.012578f
C19229 DVSS.n2883 VSS 0.011731f
C19230 DVSS.n2884 VSS 0.010244f
C19231 DVSS.n2885 VSS 0.041646f
C19232 DVSS.n2886 VSS 0.041646f
C19233 DVSS.n2887 VSS 0.010244f
C19234 DVSS.n2888 VSS 0.011731f
C19235 DVSS.n2889 VSS 0.012578f
C19236 DVSS.n2890 VSS 0.022081f
C19237 DVSS.n2891 VSS 0.011731f
C19238 DVSS.n2892 VSS 0.010244f
C19239 DVSS.n2893 VSS 0.041646f
C19240 DVSS.n2894 VSS 0.041646f
C19241 DVSS.n2895 VSS 0.083291f
C19242 DVSS.n2896 VSS 0.083291f
C19243 DVSS.n2897 VSS 0.083291f
C19244 DVSS.n2898 VSS 0.083291f
C19245 DVSS.n2899 VSS 0.083291f
C19246 DVSS.n2900 VSS 0.083291f
C19247 DVSS.n2901 VSS 0.083291f
C19248 DVSS.n2902 VSS 0.083291f
C19249 DVSS.n2903 VSS 0.083291f
C19250 DVSS.n2904 VSS 0.041646f
C19251 DVSS.n2905 VSS 0.041646f
C19252 DVSS.n2906 VSS 0.083291f
C19253 DVSS.n2907 VSS 0.083291f
C19254 DVSS.n2908 VSS 0.041646f
C19255 DVSS.n2909 VSS 0.041646f
C19256 DVSS.n2910 VSS 0.010244f
C19257 DVSS.n2911 VSS 0.011731f
C19258 DVSS.n2912 VSS 0.023106f
C19259 DVSS.n2913 VSS 0.019938f
C19260 DVSS.n2914 VSS 0.011566f
C19261 DVSS.n2915 VSS 0.010409f
C19262 DVSS.n2916 VSS 0.014721f
C19263 DVSS.n2917 VSS 0.023106f
C19264 DVSS.n2918 VSS 0.011731f
C19265 DVSS.n2919 VSS 0.010244f
C19266 DVSS.n2920 VSS 0.041646f
C19267 DVSS.n2921 VSS 0.010244f
C19268 DVSS.n2922 VSS 0.011731f
C19269 DVSS.n2923 VSS 0.023106f
C19270 DVSS.n2924 VSS 0.023106f
C19271 DVSS.n2925 VSS 0.013696f
C19272 DVSS.n2926 VSS 0.010244f
C19273 DVSS.n2927 VSS 0.011731f
C19274 DVSS.n2928 VSS 0.021056f
C19275 DVSS.n2929 VSS 0.011731f
C19276 DVSS.n2930 VSS 0.023106f
C19277 DVSS.n2931 VSS 0.011731f
C19278 DVSS.n2932 VSS 0.023106f
C19279 DVSS.n2933 VSS 0.020963f
C19280 DVSS.n2934 VSS 0.010575f
C19281 DVSS.n2935 VSS 0.011401f
C19282 DVSS.n2936 VSS 0.010244f
C19283 DVSS.n2937 VSS 0.011731f
C19284 DVSS.n2938 VSS 0.014162f
C19285 DVSS.n2939 VSS 0.021288f
C19286 DVSS.n2940 VSS 0.011731f
C19287 DVSS.n2941 VSS 0.020497f
C19288 DVSS.n2942 VSS 0.011731f
C19289 DVSS.n2943 VSS 0.023106f
C19290 DVSS.n2944 VSS 0.023106f
C19291 DVSS.n2945 VSS 0.011731f
C19292 DVSS.n2946 VSS 0.010244f
C19293 DVSS.n2947 VSS 0.041646f
C19294 DVSS.n2948 VSS 0.041646f
C19295 DVSS.n2949 VSS 0.010244f
C19296 DVSS.n2950 VSS 0.011731f
C19297 DVSS.n2951 VSS 0.023106f
C19298 DVSS.n2952 VSS 0.020497f
C19299 DVSS.n2953 VSS 0.023106f
C19300 DVSS.n2954 VSS 0.011731f
C19301 DVSS.n2955 VSS 0.010244f
C19302 DVSS.n2956 VSS 0.041646f
C19303 DVSS.n2957 VSS 0.041646f
C19304 DVSS.n2958 VSS 0.083291f
C19305 DVSS.n2959 VSS 0.083291f
C19306 DVSS.n2960 VSS 0.083291f
C19307 DVSS.n2961 VSS 0.083291f
C19308 DVSS.n2962 VSS 0.083291f
C19309 DVSS.n2963 VSS 0.041646f
C19310 DVSS.n2964 VSS 0.041646f
C19311 DVSS.n2965 VSS 0.010244f
C19312 DVSS.n2966 VSS 0.011731f
C19313 DVSS.n2967 VSS 0.014162f
C19314 DVSS.n2968 VSS 0.013696f
C19315 DVSS.n2969 VSS 0.011401f
C19316 DVSS.n2970 VSS 0.010575f
C19317 DVSS.n2971 VSS 0.020963f
C19318 DVSS.n2972 VSS 0.023106f
C19319 DVSS.n2973 VSS 0.011731f
C19320 DVSS.n2974 VSS 0.010244f
C19321 DVSS.n2975 VSS 0.041646f
C19322 DVSS.n2976 VSS 0.041646f
C19323 DVSS.n2977 VSS 0.083291f
C19324 DVSS.n2978 VSS 0.083291f
C19325 DVSS.n2979 VSS 0.083291f
C19326 DVSS.n2980 VSS 0.083291f
C19327 DVSS.n2981 VSS 0.083291f
C19328 DVSS.n2982 VSS 0.083291f
C19329 DVSS.n2983 VSS 0.083291f
C19330 DVSS.n2984 VSS 0.083291f
C19331 DVSS.n2985 VSS 0.083291f
C19332 DVSS.n2986 VSS 0.041646f
C19333 DVSS.n2987 VSS 0.041646f
C19334 DVSS.n2988 VSS 0.010244f
C19335 DVSS.n2989 VSS 0.011731f
C19336 DVSS.n2990 VSS 0.021056f
C19337 DVSS.n2991 VSS 0.019264f
C19338 DVSS.n2992 VSS 0.013603f
C19339 DVSS.n2993 VSS 0.011731f
C19340 DVSS.n2994 VSS 0.010244f
C19341 DVSS.n2995 VSS 0.041646f
C19342 DVSS.n2996 VSS 0.010244f
C19343 DVSS.n2997 VSS 0.011731f
C19344 DVSS.n2998 VSS 0.013603f
C19345 DVSS.n2999 VSS 0.023106f
C19346 DVSS.n3000 VSS 0.021288f
C19347 DVSS.n3001 VSS 0.011731f
C19348 DVSS.n3002 VSS 0.021615f
C19349 DVSS.n3003 VSS 0.023106f
C19350 DVSS.n3004 VSS 0.01074f
C19351 DVSS.n3005 VSS 0.011235f
C19352 DVSS.n3006 VSS 0.023106f
C19353 DVSS.n3007 VSS 0.023106f
C19354 DVSS.n3008 VSS 0.011731f
C19355 DVSS.n3009 VSS 0.010244f
C19356 DVSS.n3010 VSS 0.041646f
C19357 DVSS.n3011 VSS 0.041646f
C19358 DVSS.n3012 VSS 0.010244f
C19359 DVSS.n3013 VSS 0.010244f
C19360 DVSS.n3014 VSS 0.011731f
C19361 DVSS.n3015 VSS 0.023106f
C19362 DVSS.n3016 VSS 0.023106f
C19363 DVSS.n3017 VSS 0.021615f
C19364 DVSS.n3018 VSS 0.023106f
C19365 DVSS.n3019 VSS 0.01074f
C19366 DVSS.n3020 VSS 0.010244f
C19367 DVSS.n3021 VSS 0.041646f
C19368 DVSS.n3022 VSS 0.041646f
C19369 DVSS.n3023 VSS 0.083291f
C19370 DVSS.n3024 VSS 0.083291f
C19371 DVSS.n3025 VSS 0.083291f
C19372 DVSS.n3026 VSS 0.083291f
C19373 DVSS.n3027 VSS 0.083291f
C19374 DVSS.n3028 VSS 0.083291f
C19375 DVSS.n3029 VSS 0.083291f
C19376 DVSS.n3030 VSS 0.083291f
C19377 DVSS.n3031 VSS 0.083291f
C19378 DVSS.n3032 VSS 0.083291f
C19379 DVSS.n3033 VSS 0.041646f
C19380 DVSS.n3034 VSS 0.041646f
C19381 DVSS.n3035 VSS 0.010244f
C19382 DVSS.n3036 VSS 0.011731f
C19383 DVSS.n3037 VSS 0.013044f
C19384 DVSS.n3038 VSS 0.014814f
C19385 DVSS.n3039 VSS 0.011731f
C19386 DVSS.n3040 VSS 0.010244f
C19387 DVSS.n3041 VSS 0.041646f
C19388 DVSS.n3042 VSS 0.010244f
C19389 DVSS.n3043 VSS 0.011731f
C19390 DVSS.n3044 VSS 0.014814f
C19391 DVSS.n3045 VSS 0.019845f
C19392 DVSS.n3046 VSS 0.011731f
C19393 DVSS.n3047 VSS 0.023106f
C19394 DVSS.n3048 VSS 0.023106f
C19395 DVSS.n3049 VSS 0.011731f
C19396 DVSS.n3050 VSS 0.010244f
C19397 DVSS.n3051 VSS 0.041646f
C19398 DVSS.n3052 VSS 0.041646f
C19399 DVSS.n3053 VSS 0.010244f
C19400 DVSS.n3054 VSS 0.010244f
C19401 DVSS.n3055 VSS 0.011731f
C19402 DVSS.n3056 VSS 0.023106f
C19403 DVSS.n3057 VSS 0.023106f
C19404 DVSS.n3058 VSS 0.019264f
C19405 DVSS.n3059 VSS 0.022174f
C19406 DVSS.n3060 VSS 0.01107f
C19407 DVSS.n3061 VSS 0.010244f
C19408 DVSS.n3062 VSS 0.041646f
C19409 DVSS.n3063 VSS 0.041646f
C19410 DVSS.n3064 VSS 0.083291f
C19411 DVSS.n3065 VSS 0.083291f
C19412 DVSS.n3066 VSS 0.083291f
C19413 DVSS.n3067 VSS 0.083291f
C19414 DVSS.n3068 VSS 0.083291f
C19415 DVSS.n3069 VSS 0.083291f
C19416 DVSS.n3070 VSS 0.083291f
C19417 DVSS.n3071 VSS 0.083291f
C19418 DVSS.n3072 VSS 0.010244f
C19419 DVSS.n3073 VSS 0.041646f
C19420 DVSS.n3074 VSS 0.010244f
C19421 DVSS.n3075 VSS 0.011731f
C19422 DVSS.n3076 VSS 0.010244f
C19423 DVSS.n3077 VSS 0.023106f
C19424 DVSS.n3078 VSS 0.011553f
C19425 DVSS.n3079 VSS 0.010905f
C19426 DVSS.n3080 VSS 0.041646f
C19427 DVSS.n3081 VSS 0.010244f
C19428 DVSS.n3082 VSS 0.041646f
C19429 DVSS.n3083 VSS 0.083291f
C19430 DVSS.n3084 VSS 0.083291f
C19431 DVSS.n3085 VSS 0.083291f
C19432 DVSS.n3086 VSS 0.083291f
C19433 DVSS.n3087 VSS 0.083291f
C19434 DVSS.n3088 VSS 0.083291f
C19435 DVSS.n3089 VSS 0.010244f
C19436 DVSS.n3090 VSS 0.041646f
C19437 DVSS.n3091 VSS 0.011731f
C19438 DVSS.n3092 VSS 0.010244f
C19439 DVSS.n3093 VSS 0.005124f
C19440 DVSS.n3094 VSS 0.010244f
C19441 DVSS.n3095 VSS 0.01107f
C19442 DVSS.n3096 VSS 0.018727f
C19443 DVSS.n3097 VSS 0.023106f
C19444 DVSS.n3098 VSS 0.011739f
C19445 DVSS.n3099 VSS 0.011731f
C19446 DVSS.n3100 VSS 0.041646f
C19447 DVSS.n3101 VSS 0.010244f
C19448 DVSS.n3102 VSS 0.041646f
C19449 DVSS.n3103 VSS 0.083291f
C19450 DVSS.n3104 VSS 0.083291f
C19451 DVSS.n3105 VSS 0.083291f
C19452 DVSS.n3106 VSS 0.083291f
C19453 DVSS.n3107 VSS 0.083291f
C19454 DVSS.n3108 VSS 0.083291f
C19455 DVSS.n3109 VSS 0.010244f
C19456 DVSS.n3110 VSS 0.041646f
C19457 DVSS.n3111 VSS 0.010244f
C19458 DVSS.n3112 VSS 0.011731f
C19459 DVSS.n3113 VSS 0.010244f
C19460 DVSS.n3114 VSS 0.02292f
C19461 DVSS.n3115 VSS 0.023106f
C19462 DVSS.n3116 VSS 0.011731f
C19463 DVSS.n3117 VSS 0.041646f
C19464 DVSS.n3118 VSS 0.010244f
C19465 DVSS.n3119 VSS 0.041646f
C19466 DVSS.n3120 VSS 0.083291f
C19467 DVSS.n3121 VSS 0.083291f
C19468 DVSS.n3122 VSS 0.083291f
C19469 DVSS.n3123 VSS 0.083291f
C19470 DVSS.n3124 VSS 0.083291f
C19471 DVSS.n3125 VSS 0.083291f
C19472 DVSS.n3126 VSS 0.010244f
C19473 DVSS.n3127 VSS 0.041646f
C19474 DVSS.n3128 VSS 0.010244f
C19475 DVSS.n3129 VSS 0.011731f
C19476 DVSS.n3130 VSS 0.010244f
C19477 DVSS.n3131 VSS 0.023106f
C19478 DVSS.n3132 VSS 0.012298f
C19479 DVSS.t46 VSS 0.061308f
C19480 DVSS.n3133 VSS 0.021288f
C19481 DVSS.n3134 VSS 0.023106f
C19482 DVSS.n3135 VSS 0.011731f
C19483 DVSS.n3136 VSS 0.041646f
C19484 DVSS.n3137 VSS 0.010244f
C19485 DVSS.n3138 VSS 0.041646f
C19486 DVSS.n3139 VSS 0.083291f
C19487 DVSS.n3140 VSS 0.083291f
C19488 DVSS.n3141 VSS 0.083291f
C19489 DVSS.n3142 VSS 0.083291f
C19490 DVSS.n3143 VSS 0.083291f
C19491 DVSS.n3144 VSS 0.083291f
C19492 DVSS.n3145 VSS 0.010244f
C19493 DVSS.n3146 VSS 0.041646f
C19494 DVSS.n3147 VSS 0.010244f
C19495 DVSS.n3148 VSS 0.011731f
C19496 DVSS.n3149 VSS 0.011401f
C19497 DVSS.n3150 VSS 0.023106f
C19498 DVSS.n3151 VSS 0.023106f
C19499 DVSS.n3152 VSS 0.010244f
C19500 DVSS.n3153 VSS 0.011731f
C19501 DVSS.n3154 VSS 0.041646f
C19502 DVSS.n3155 VSS 0.010244f
C19503 DVSS.n3156 VSS 0.041646f
C19504 DVSS.n3157 VSS 0.083291f
C19505 DVSS.n3158 VSS 0.083291f
C19506 DVSS.n3159 VSS 0.083291f
C19507 DVSS.n3160 VSS 0.083291f
C19508 DVSS.n3161 VSS 0.083291f
C19509 DVSS.n3162 VSS 0.083291f
C19510 DVSS.n3163 VSS 0.010244f
C19511 DVSS.n3164 VSS 0.041646f
C19512 DVSS.n3165 VSS 0.010244f
C19513 DVSS.n3166 VSS 0.011731f
C19514 DVSS.n3167 VSS 0.010244f
C19515 DVSS.n3168 VSS 0.023106f
C19516 DVSS.n3169 VSS 0.013416f
C19517 DVSS.n3170 VSS 0.011731f
C19518 DVSS.n3171 VSS 0.041646f
C19519 DVSS.n3172 VSS 0.010244f
C19520 DVSS.n3173 VSS 0.041646f
C19521 DVSS.n3174 VSS 0.083291f
C19522 DVSS.n3175 VSS 0.083291f
C19523 DVSS.n3176 VSS 0.083291f
C19524 DVSS.n3177 VSS 0.083291f
C19525 DVSS.n3178 VSS 0.083291f
C19526 DVSS.n3179 VSS 0.083291f
C19527 DVSS.n3180 VSS 0.010244f
C19528 DVSS.n3181 VSS 0.041646f
C19529 DVSS.n3182 VSS 0.011566f
C19530 DVSS.n3183 VSS 0.010244f
C19531 DVSS.t36 VSS 0.061308f
C19532 DVSS.n3184 VSS 0.021288f
C19533 DVSS.n3185 VSS 0.010244f
C19534 DVSS.n3186 VSS 0.010409f
C19535 DVSS.n3187 VSS 0.016305f
C19536 DVSS.n3188 VSS 0.016491f
C19537 DVSS.n3189 VSS 0.023106f
C19538 DVSS.n3190 VSS 0.011731f
C19539 DVSS.n3191 VSS 0.041646f
C19540 DVSS.n3192 VSS 0.010244f
C19541 DVSS.n3193 VSS 0.041646f
C19542 DVSS.n3194 VSS 0.083291f
C19543 DVSS.n3195 VSS 0.083291f
C19544 DVSS.n3196 VSS 0.083291f
C19545 DVSS.n3197 VSS 0.083291f
C19546 DVSS.n3198 VSS 0.083291f
C19547 DVSS.n3199 VSS 0.083291f
C19548 DVSS.n3200 VSS 0.010244f
C19549 DVSS.n3201 VSS 0.041646f
C19550 DVSS.n3202 VSS 0.010244f
C19551 DVSS.n3203 VSS 0.011731f
C19552 DVSS.n3204 VSS 0.010244f
C19553 DVSS.n3205 VSS 0.013975f
C19554 DVSS.n3206 VSS 0.019264f
C19555 DVSS.n3207 VSS 0.023106f
C19556 DVSS.n3208 VSS 0.011731f
C19557 DVSS.n3209 VSS 0.041646f
C19558 DVSS.n3210 VSS 0.020488f
C19559 DVSS.n3211 VSS 0.041646f
C19560 DVSS.n3212 VSS 0.083291f
C19561 DVSS.n3213 VSS 0.083291f
C19562 DVSS.n3214 VSS 0.083291f
C19563 DVSS.n3215 VSS 0.083291f
C19564 DVSS.n3216 VSS 0.083291f
C19565 DVSS.n3217 VSS 0.083291f
C19566 DVSS.n3218 VSS 0.010244f
C19567 DVSS.n3219 VSS 0.041646f
C19568 DVSS.n3220 VSS 0.010244f
C19569 DVSS.n3221 VSS 0.011731f
C19570 DVSS.n3222 VSS 0.010244f
C19571 DVSS.n3223 VSS 0.023106f
C19572 DVSS.n3224 VSS 0.023106f
C19573 DVSS.n3225 VSS 0.011731f
C19574 DVSS.n3226 VSS 0.041646f
C19575 DVSS.n3227 VSS 0.010244f
C19576 DVSS.n3228 VSS 0.041646f
C19577 DVSS.n3229 VSS 0.083291f
C19578 DVSS.n3230 VSS 0.083291f
C19579 DVSS.n3231 VSS 0.083291f
C19580 DVSS.n3232 VSS 0.083291f
C19581 DVSS.n3233 VSS 0.083291f
C19582 DVSS.n3234 VSS 0.083291f
C19583 DVSS.n3235 VSS 0.010244f
C19584 DVSS.n3236 VSS 0.041646f
C19585 DVSS.n3237 VSS 0.010244f
C19586 DVSS.n3238 VSS 0.011731f
C19587 DVSS.n3239 VSS 0.010409f
C19588 DVSS.n3240 VSS 0.015373f
C19589 DVSS.n3241 VSS 0.023106f
C19590 DVSS.n3242 VSS 0.010244f
C19591 DVSS.n3243 VSS 0.041646f
C19592 DVSS.n3244 VSS 0.011566f
C19593 DVSS.n3245 VSS 0.021288f
C19594 DVSS.n3246 VSS 0.010244f
C19595 DVSS.n3247 VSS 0.019264f
C19596 DVSS.n3248 VSS 0.010575f
C19597 DVSS.n3249 VSS 0.023106f
C19598 DVSS.n3250 VSS 0.019264f
C19599 DVSS.n3251 VSS 0.019264f
C19600 DVSS.n3252 VSS 0.018727f
C19601 DVSS.n3253 VSS 0.021288f
C19602 DVSS.n3254 VSS 0.041646f
C19603 DVSS.n3255 VSS 0.010244f
C19604 DVSS.n3256 VSS 0.011731f
C19605 DVSS.n3257 VSS 0.023106f
C19606 DVSS.n3258 VSS 0.023106f
C19607 DVSS.n3259 VSS 0.011731f
C19608 DVSS.n3260 VSS 0.010244f
C19609 DVSS.n3261 VSS 0.011731f
C19610 DVSS.n3262 VSS 0.023106f
C19611 DVSS.n3263 VSS 0.022733f
C19612 DVSS.n3264 VSS 0.011731f
C19613 DVSS.n3265 VSS 0.041646f
C19614 DVSS.n3266 VSS 0.010244f
C19615 DVSS.n3267 VSS 0.011731f
C19616 DVSS.n3268 VSS 0.011926f
C19617 DVSS.n3269 VSS 0.015932f
C19618 DVSS.n3270 VSS 0.010905f
C19619 DVSS.n3271 VSS 0.01107f
C19620 DVSS.n3272 VSS 0.010244f
C19621 DVSS.n3273 VSS 0.011731f
C19622 DVSS.n3274 VSS 0.023106f
C19623 DVSS.n3275 VSS 0.023106f
C19624 DVSS.n3276 VSS 0.011731f
C19625 DVSS.n3277 VSS 0.041646f
C19626 DVSS.n3278 VSS 0.010244f
C19627 DVSS.n3279 VSS 0.011731f
C19628 DVSS.n3280 VSS 0.023106f
C19629 DVSS.n3281 VSS 0.011739f
C19630 DVSS.n3282 VSS 0.011731f
C19631 DVSS.n3283 VSS 0.010244f
C19632 DVSS.n3284 VSS 0.011731f
C19633 DVSS.n3285 VSS 0.02292f
C19634 DVSS.n3286 VSS 0.023106f
C19635 DVSS.n3287 VSS 0.011731f
C19636 DVSS.n3288 VSS 0.041646f
C19637 DVSS.n3289 VSS 0.010244f
C19638 DVSS.n3290 VSS 0.01074f
C19639 DVSS.n3291 VSS 0.011235f
C19640 DVSS.n3292 VSS 0.023106f
C19641 DVSS.n3293 VSS 0.023106f
C19642 DVSS.n3294 VSS 0.011731f
C19643 DVSS.n3295 VSS 0.010244f
C19644 DVSS.n3296 VSS 0.011731f
C19645 DVSS.n3297 VSS 0.012298f
C19646 DVSS.n3298 VSS 0.021288f
C19647 DVSS.n3299 VSS 0.016305f
C19648 DVSS.n3300 VSS 0.011731f
C19649 DVSS.n3301 VSS 0.041646f
C19650 DVSS.n3302 VSS 0.010244f
C19651 DVSS.n3303 VSS 0.011731f
C19652 DVSS.n3304 VSS 0.017609f
C19653 DVSS.n3305 VSS 0.023106f
C19654 DVSS.n3306 VSS 0.011731f
C19655 DVSS.n3307 VSS 0.010244f
C19656 DVSS.n3308 VSS 0.011731f
C19657 DVSS.n3309 VSS 0.023106f
C19658 DVSS.n3310 VSS 0.023106f
C19659 DVSS.n3311 VSS 0.012857f
C19660 DVSS.n3312 VSS 0.011401f
C19661 DVSS.n3313 VSS 0.041646f
C19662 DVSS.n3314 VSS 0.010244f
C19663 DVSS.n3315 VSS 0.011731f
C19664 DVSS.n3316 VSS 0.021802f
C19665 DVSS.n3317 VSS 0.023106f
C19666 DVSS.n3318 VSS 0.011731f
C19667 DVSS.n3319 VSS 0.010244f
C19668 DVSS.n3320 VSS 0.011731f
C19669 DVSS.n3321 VSS 0.023106f
C19670 DVSS.n3322 VSS 0.023106f
C19671 DVSS.n3323 VSS 0.011731f
C19672 DVSS.n3324 VSS 0.041646f
C19673 DVSS.n3325 VSS 0.010244f
C19674 DVSS.n3326 VSS 0.011731f
C19675 DVSS.n3327 VSS 0.023106f
C19676 DVSS.n3328 VSS 0.011731f
C19677 DVSS.n3329 VSS 0.013416f
C19678 DVSS.n3330 VSS 0.021288f
C19679 DVSS.n3331 VSS 0.016305f
C19680 DVSS.n3332 VSS 0.010409f
C19681 DVSS.n3333 VSS 0.011566f
C19682 DVSS.n3334 VSS 0.016491f
C19683 DVSS.n3335 VSS 0.023106f
C19684 DVSS.n3336 VSS 0.011731f
C19685 DVSS.n3337 VSS 0.041646f
C19686 DVSS.n3338 VSS 0.010244f
C19687 DVSS.n3339 VSS 0.011731f
C19688 DVSS.n3340 VSS 0.023106f
C19689 DVSS.n3341 VSS 0.023106f
C19690 DVSS.n3342 VSS 0.011731f
C19691 DVSS.n3343 VSS 0.010244f
C19692 DVSS.n3344 VSS 0.011731f
C19693 DVSS.n3345 VSS 0.013975f
C19694 DVSS.n3346 VSS 0.019264f
C19695 DVSS.n3347 VSS 0.020684f
C19696 DVSS.n3348 VSS 0.011731f
C19697 DVSS.n3349 VSS 0.041646f
C19698 DVSS.n3350 VSS 0.010244f
C19699 DVSS.n3351 VSS 0.011731f
C19700 DVSS.n3352 VSS 0.023106f
C19701 DVSS.n3353 VSS 0.023106f
C19702 DVSS.n3354 VSS 0.023106f
C19703 DVSS.n3355 VSS 0.011731f
C19704 DVSS.n3356 VSS 0.010244f
C19705 DVSS.n3357 VSS 0.011731f
C19706 DVSS.n3358 VSS 0.023106f
C19707 DVSS.n3359 VSS 0.014534f
C19708 DVSS.n3360 VSS 0.011731f
C19709 DVSS.n3361 VSS 0.041646f
C19710 DVSS.n3362 VSS 0.010244f
C19711 DVSS.n3363 VSS 0.011731f
C19712 DVSS.n3364 VSS 0.016305f
C19713 DVSS.n3365 VSS 0.015373f
C19714 DVSS.n3366 VSS 0.011731f
C19715 DVSS.n3367 VSS 0.010244f
C19716 DVSS.n3368 VSS 0.011731f
C19717 DVSS.n3369 VSS 0.023106f
C19718 DVSS.n3370 VSS 0.023106f
C19719 DVSS.n3371 VSS 0.023106f
C19720 DVSS.n3372 VSS 0.010409f
C19721 DVSS.n3373 VSS 0.041646f
C19722 DVSS.n3374 VSS 0.010244f
C19723 DVSS.n3375 VSS 0.019636f
C19724 DVSS.n3376 VSS 0.083291f
C19725 DVSS.n3377 VSS 0.083291f
C19726 DVSS.n3378 VSS 0.083291f
C19727 DVSS.n3379 VSS 0.083291f
C19728 DVSS.n3380 VSS 0.083291f
C19729 DVSS.n3381 VSS 0.083291f
C19730 DVSS.n3382 VSS 0.083291f
C19731 DVSS.n3383 VSS 0.083291f
C19732 DVSS.n3384 VSS 0.083291f
C19733 DVSS.n3385 VSS 0.083291f
C19734 DVSS.n3386 VSS 0.083291f
C19735 DVSS.n3387 VSS 0.083291f
C19736 DVSS.n3388 VSS 0.083291f
C19737 DVSS.n3389 VSS 0.083291f
C19738 DVSS.n3390 VSS 0.083291f
C19739 DVSS.n3391 VSS 0.083291f
C19740 DVSS.n3392 VSS 0.083291f
C19741 DVSS.n3393 VSS 0.083291f
C19742 DVSS.n3394 VSS 0.083291f
C19743 DVSS.n3395 VSS 0.075079f
C19744 DVSS.n3396 VSS 0.009385f
C19745 DVSS.n3397 VSS 0.402052f
C19746 DVSS.n3398 VSS 0.109006f
C19747 DVSS.n3399 VSS 0.075079f
C19748 DVSS.n3400 VSS 0.075079f
C19749 DVSS.n3401 VSS 0.083291f
C19750 DVSS.n3402 VSS 0.083291f
C19751 DVSS.n3403 VSS 0.083291f
C19752 DVSS.n3404 VSS 0.083291f
C19753 DVSS.n3405 VSS 0.083291f
C19754 DVSS.n3406 VSS 0.083291f
C19755 DVSS.n3407 VSS 0.083291f
C19756 DVSS.n3408 VSS 0.082998f
C19757 DVSS.n3409 VSS 0.083291f
C19758 DVSS.n3410 VSS 0.083291f
C19759 DVSS.n3411 VSS 0.041939f
C19760 DVSS.n3412 VSS 0.083291f
C19761 DVSS.n3413 VSS 0.083291f
C19762 DVSS.n3414 VSS 0.083291f
C19763 DVSS.n3415 VSS 0.083291f
C19764 DVSS.n3416 VSS 0.083291f
C19765 DVSS.n3417 VSS 0.05191f
C19766 DVSS.n3418 VSS 0.041698f
C19767 DVSS.n3419 VSS 0.019636f
C19768 DVSS.n3420 VSS 0.018261f
C19769 DVSS.n3421 VSS 0.023106f
C19770 DVSS.n3422 VSS 0.023106f
C19771 DVSS.n3423 VSS 0.011566f
C19772 DVSS.n3424 VSS 0.010244f
C19773 DVSS.n3425 VSS 0.041646f
C19774 DVSS.n3426 VSS 0.041646f
C19775 DVSS.n3427 VSS 0.083291f
C19776 DVSS.n3428 VSS 0.083291f
C19777 DVSS.n3429 VSS 0.041646f
C19778 DVSS.n3430 VSS 0.041646f
C19779 DVSS.n3431 VSS 0.010244f
C19780 DVSS.n3432 VSS 0.011731f
C19781 DVSS.n3433 VSS 0.016305f
C19782 DVSS.t49 VSS 0.061308f
C19783 DVSS.n3434 VSS 0.021288f
C19784 DVSS.n3435 VSS 0.014534f
C19785 DVSS.n3436 VSS 0.011731f
C19786 DVSS.n3437 VSS 0.010244f
C19787 DVSS.n3438 VSS 0.041646f
C19788 DVSS.n3439 VSS 0.041646f
C19789 DVSS.n3440 VSS 0.083291f
C19790 DVSS.n3441 VSS 0.083291f
C19791 DVSS.n3442 VSS 0.041646f
C19792 DVSS.n3443 VSS 0.041646f
C19793 DVSS.n3444 VSS 0.020488f
C19794 DVSS.n3445 VSS 0.011731f
C19795 DVSS.n3446 VSS 0.023106f
C19796 DVSS.n3447 VSS 0.020684f
C19797 DVSS.n3448 VSS 0.011731f
C19798 DVSS.n3449 VSS 0.010244f
C19799 DVSS.n3450 VSS 0.041646f
C19800 DVSS.n3451 VSS 0.041646f
C19801 DVSS.n3452 VSS 0.083291f
C19802 DVSS.n3453 VSS 0.083291f
C19803 DVSS.n3454 VSS 0.041646f
C19804 DVSS.n3455 VSS 0.041646f
C19805 DVSS.n3456 VSS 0.010244f
C19806 DVSS.n3457 VSS 0.011731f
C19807 DVSS.n3458 VSS 0.023106f
C19808 DVSS.n3459 VSS 0.023106f
C19809 DVSS.n3460 VSS 0.011731f
C19810 DVSS.n3461 VSS 0.010244f
C19811 DVSS.n3462 VSS 0.041646f
C19812 DVSS.n3463 VSS 0.041646f
C19813 DVSS.n3464 VSS 0.083291f
C19814 DVSS.n3465 VSS 0.083291f
C19815 DVSS.n3466 VSS 0.041646f
C19816 DVSS.n3467 VSS 0.041646f
C19817 DVSS.n3468 VSS 0.010244f
C19818 DVSS.n3469 VSS 0.011731f
C19819 DVSS.n3470 VSS 0.023106f
C19820 DVSS.n3471 VSS 0.023106f
C19821 DVSS.n3472 VSS 0.011731f
C19822 DVSS.n3473 VSS 0.010244f
C19823 DVSS.n3474 VSS 0.041646f
C19824 DVSS.n3475 VSS 0.041646f
C19825 DVSS.n3476 VSS 0.083291f
C19826 DVSS.n3477 VSS 0.083291f
C19827 DVSS.n3478 VSS 0.041646f
C19828 DVSS.n3479 VSS 0.041646f
C19829 DVSS.n3480 VSS 0.010244f
C19830 DVSS.n3481 VSS 0.011731f
C19831 DVSS.n3482 VSS 0.021802f
C19832 DVSS.n3483 VSS 0.019264f
C19833 DVSS.n3484 VSS 0.012857f
C19834 DVSS.n3485 VSS 0.023106f
C19835 DVSS.n3486 VSS 0.010575f
C19836 DVSS.n3487 VSS 0.010244f
C19837 DVSS.n3488 VSS 0.041646f
C19838 DVSS.n3489 VSS 0.041646f
C19839 DVSS.n3490 VSS 0.083291f
C19840 DVSS.n3491 VSS 0.083291f
C19841 DVSS.n3492 VSS 0.041646f
C19842 DVSS.n3493 VSS 0.041646f
C19843 DVSS.n3494 VSS 0.010244f
C19844 DVSS.n3495 VSS 0.011731f
C19845 DVSS.n3496 VSS 0.017609f
C19846 DVSS.n3497 VSS 0.016305f
C19847 DVSS.n3498 VSS 0.011731f
C19848 DVSS.n3499 VSS 0.010244f
C19849 DVSS.n3500 VSS 0.041646f
C19850 DVSS.n3501 VSS 0.041646f
C19851 DVSS.n3502 VSS 0.083291f
C19852 DVSS.n3503 VSS 0.083291f
C19853 DVSS.n3504 VSS 0.041646f
C19854 DVSS.n3505 VSS 0.041646f
C19855 DVSS.n3506 VSS 0.010244f
C19856 DVSS.n3507 VSS 0.011235f
C19857 DVSS.n3508 VSS 0.01074f
C19858 DVSS.n3509 VSS 0.023106f
C19859 DVSS.n3510 VSS 0.023106f
C19860 DVSS.n3511 VSS 0.011731f
C19861 DVSS.n3512 VSS 0.010244f
C19862 DVSS.n3513 VSS 0.041646f
C19863 DVSS.n3514 VSS 0.041646f
C19864 DVSS.n3515 VSS 0.083291f
C19865 DVSS.n3516 VSS 0.083291f
C19866 DVSS.n3517 VSS 0.041646f
C19867 DVSS.n3518 VSS 0.041646f
C19868 DVSS.n3519 VSS 0.010244f
C19869 DVSS.n3520 VSS 0.011731f
C19870 DVSS.n3521 VSS 0.023106f
C19871 DVSS.n3522 VSS 0.023106f
C19872 DVSS.n3523 VSS 0.011731f
C19873 DVSS.n3524 VSS 0.010244f
C19874 DVSS.n3525 VSS 0.041646f
C19875 DVSS.n3526 VSS 0.041646f
C19876 DVSS.n3527 VSS 0.083291f
C19877 DVSS.n3528 VSS 0.083291f
C19878 DVSS.n3529 VSS 0.041646f
C19879 DVSS.n3530 VSS 0.041646f
C19880 DVSS.n3531 VSS 0.010244f
C19881 DVSS.n3532 VSS 0.011731f
C19882 DVSS.n3533 VSS 0.01118f
C19883 DVSS.t34 VSS 0.061308f
C19884 DVSS.n3534 VSS 0.021288f
C19885 DVSS.n3535 VSS 0.022733f
C19886 DVSS.n3536 VSS 0.011731f
C19887 DVSS.n3537 VSS 0.010244f
C19888 DVSS.n3538 VSS 0.041646f
C19889 DVSS.n3539 VSS 0.041646f
C19890 DVSS.n3540 VSS 0.083291f
C19891 DVSS.n3541 VSS 0.083291f
C19892 DVSS.n3542 VSS 0.041646f
C19893 DVSS.n3543 VSS 0.041646f
C19894 DVSS.n3544 VSS 0.010244f
C19895 DVSS.n3545 VSS 0.011731f
C19896 DVSS.n3546 VSS 0.023106f
C19897 DVSS.n3547 VSS 0.023106f
C19898 DVSS.n3548 VSS 0.011731f
C19899 DVSS.n3549 VSS 0.010244f
C19900 DVSS.n3550 VSS 0.041646f
C19901 DVSS.n3551 VSS 0.010244f
C19902 DVSS.n3552 VSS 0.010905f
C19903 DVSS.n3553 VSS 0.012485f
C19904 DVSS.n3554 VSS 0.010785f
C19905 DVSS.n3555 VSS 0.010621f
C19906 DVSS.n3556 VSS 0.264688f
C19907 DVSS.n3557 VSS 0.736899f
C19908 DVSS.n3558 VSS 1.78375f
C19909 DVSS.n3559 VSS 1.9237f
C19910 DVSS.t134 VSS 0.270381f
C19911 DVSS.t132 VSS 0.224453f
C19912 DVSS.n3560 VSS 0.017292f
C19913 DVSS.n3561 VSS 0.016314f
C19914 DVSS.n3562 VSS 0.020324f
C19915 DVSS.n3563 VSS 0.017051f
C19916 DVSS.n3564 VSS -0.053672f
C19917 DVSS.n3565 VSS 0.166574f
C19918 DVSS.n3566 VSS 0.383816f
C19919 DVSS.n3567 VSS 0.542461f
C19920 DVSS.n3568 VSS 0.474092f
C19921 DVSS.n3569 VSS 0.506686f
C19922 DVSS.n3570 VSS 0.032717f
C19923 DVSS.n3571 VSS 0.012545f
C19924 DVSS.n3572 VSS 0.122398f
C19925 DVSS.n3573 VSS 0.144857f
C19926 DVSS.n3574 VSS 0.030051f
C19927 DVSS.n3575 VSS 0.058251f
C19928 DVSS.n3576 VSS 0.013846f
C19929 DVSS.n3577 VSS 0.032049f
C19930 DVSS.n3578 VSS 0.02291f
C19931 DVSS.n3579 VSS 0.272603f
C19932 DVSS.n3580 VSS 0.165826f
C19933 DVSS.n3581 VSS 0.042514f
C19934 DVSS.t59 VSS 0.004535f
C19935 DVSS.t58 VSS 0.004535f
C19936 DVSS.n3582 VSS 0.081701f
C19937 DVSS.n3583 VSS 0.097495f
C19938 DVSS.n3584 VSS 0.014888f
C19939 DVSS.n3585 VSS 0.021171f
C19940 DVSS.n3586 VSS -0.009054f
C19941 DVSS.n3587 VSS 0.154468f
C19942 DVSS.t103 VSS 0.145191f
C19943 DVSS.n3588 VSS 0.277025f
C19944 DVSS.n3589 VSS 1.30727f
C19945 DVSS.n3590 VSS 1.87801f
C19946 DVSS.n3591 VSS 2.21408f
C19947 DVSS.n3592 VSS 2.50959f
C19948 DVSS.n3594 VSS 0.044009f
C19949 DVSS.n3595 VSS 0.044009f
C19950 DVSS.n3596 VSS 0.044009f
C19951 DVSS.n3597 VSS 0.044009f
C19952 DVSS.n3602 VSS 0.026238f
C19953 DVSS.t60 VSS 0.056298f
C19954 DVSS.t17 VSS 0.174081f
C19955 DVSS.n3603 VSS 0.131116f
C19956 DVSS.n3604 VSS 0.209348f
C19957 DVSS.t10 VSS 0.007546f
C19958 DVSS.n3605 VSS 0.006791f
C19959 DVSS.t12 VSS 0.007546f
C19960 DVSS.n3606 VSS 0.006791f
C19961 DVSS.t158 VSS 0.00358f
C19962 DVSS.n3607 VSS 0.008604f
C19963 DVSS.n3608 VSS 0.007294f
C19964 DVSS.t28 VSS 0.008049f
C19965 DVSS.t116 VSS 0.007637f
C19966 DVSS.t26 VSS 0.007637f
C19967 DVSS.n3609 VSS 0.016105f
C19968 DVSS.n3610 VSS 0.009806f
C19969 DVSS.t4 VSS 0.007637f
C19970 DVSS.t30 VSS 0.007637f
C19971 DVSS.n3611 VSS 0.016105f
C19972 DVSS.n3612 VSS 0.00752f
C19973 DVSS.n3613 VSS 0.082476f
C19974 DVSS.n3614 VSS 0.018914f
C19975 DVSS.n3615 VSS 0.011754f
C19976 DVSS.n3616 VSS 0.025512f
C19977 DVSS.n3617 VSS 0.018575f
C19978 DVSS.n3618 VSS 0.01972f
C19979 DVSS.n3619 VSS 0.01379f
C19980 DVSS.n3620 VSS 0.063597f
C19981 DVSS.n3621 VSS 0.10033f
C19982 DVSS.n3622 VSS 0.221503f
C19983 DVSS.n3623 VSS 0.112582f
C19984 DVSS.n3624 VSS 0.097764f
C19985 DVSS.n3628 VSS 0.044009f
C19986 DVSS.n3629 VSS 0.042959f
C19987 DVSS.n3633 VSS 0.041675f
C19988 DVSS.n3634 VSS 0.077855f
C19989 DVSS.n3635 VSS 0.042959f
C19990 DVSS.n3636 VSS 0.042959f
C19991 DVSS.n3637 VSS 0.042959f
C19992 DVSS.n3638 VSS 0.042959f
C19993 DVSS.n3639 VSS 0.042959f
C19994 DVSS.n3640 VSS 0.042959f
C19995 DVSS.n3641 VSS 0.042959f
C19996 DVSS.n3642 VSS 0.042959f
C19997 DVSS.n3643 VSS 0.042959f
C19998 DVSS.n3644 VSS 0.044009f
C19999 DVSS.n3645 VSS 0.847436f
C20000 DVSS.n3646 VSS 0.041047f
C20001 DVSS.n3647 VSS 1.12056f
C20002 DVSS.n3648 VSS 1.63488f
C20003 DVSS.n3649 VSS -0.015824f
C20004 DVSS.n3650 VSS 0.04649f
C20005 DVSS.t33 VSS 0.061308f
C20006 DVSS.n3651 VSS 0.067966f
C20007 DVSS.n3652 VSS 0.097137f
C20008 DVSS.n3653 VSS 0.032215f
C20009 DVSS.n3654 VSS 0.045942f
C20010 DVSS.n3655 VSS 0.091242f
C20011 DVSS.n3656 VSS 0.091242f
C20012 DVSS.n3657 VSS 0.091242f
C20013 DVSS.n3658 VSS 0.091242f
C20014 DVSS.n3659 VSS 0.091242f
C20015 DVSS.n3660 VSS 0.091242f
C20016 DVSS.n3661 VSS 0.091242f
C20017 DVSS.n3662 VSS 0.091242f
C20018 DVSS.n3663 VSS 0.091242f
C20019 DVSS.n3664 VSS 0.091242f
C20020 DVSS.n3665 VSS 0.091242f
C20021 DVSS.n3666 VSS 0.091242f
C20022 DVSS.n3667 VSS 0.091242f
C20023 DVSS.n3668 VSS 0.091242f
C20024 DVSS.n3669 VSS 0.091242f
C20025 DVSS.n3670 VSS 0.091242f
C20026 DVSS.n3671 VSS 0.091242f
C20027 DVSS.n3672 VSS 0.091242f
C20028 DVSS.n3673 VSS 0.091242f
C20029 DVSS.n3674 VSS 0.091242f
C20030 DVSS.n3675 VSS 0.091242f
C20031 DVSS.n3676 VSS 0.062018f
C20032 DVSS.n3677 VSS 0.05301f
C20033 DVSS.n3678 VSS 0.091242f
C20034 DVSS.n3679 VSS 0.091242f
C20035 DVSS.n3680 VSS 0.091242f
C20036 DVSS.n3681 VSS 0.091242f
C20037 DVSS.n3682 VSS 0.091242f
C20038 DVSS.n3683 VSS 0.091242f
C20039 DVSS.n3684 VSS 0.091242f
C20040 DVSS.n3685 VSS 0.091242f
C20041 DVSS.n3686 VSS 0.091242f
C20042 DVSS.n3687 VSS 0.091242f
C20043 DVSS.n3688 VSS 0.091242f
C20044 DVSS.n3689 VSS 0.091242f
C20045 DVSS.n3690 VSS 0.091242f
C20046 DVSS.n3691 VSS 0.091242f
C20047 DVSS.n3692 VSS 0.091242f
C20048 DVSS.n3693 VSS 0.091242f
C20049 DVSS.n3694 VSS 0.091242f
C20050 DVSS.n3695 VSS 0.091242f
C20051 DVSS.n3696 VSS 0.091242f
C20052 DVSS.n3697 VSS 0.091242f
C20053 DVSS.n3698 VSS 0.091242f
C20054 DVSS.n3699 VSS 0.091242f
C20055 DVSS.n3700 VSS 0.091242f
C20056 DVSS.n3701 VSS 0.091242f
C20057 DVSS.n3702 VSS 0.091242f
C20058 DVSS.n3703 VSS 0.091242f
C20059 DVSS.n3704 VSS 0.091242f
C20060 DVSS.n3705 VSS 0.091242f
C20061 DVSS.n3706 VSS 0.091242f
C20062 DVSS.n3707 VSS 0.091242f
C20063 DVSS.n3708 VSS 0.091242f
C20064 DVSS.n3709 VSS 0.091242f
C20065 DVSS.n3710 VSS 0.091242f
C20066 DVSS.n3711 VSS 0.091242f
C20067 DVSS.n3712 VSS 0.091242f
C20068 DVSS.n3713 VSS 0.091242f
C20069 DVSS.n3714 VSS 0.091242f
C20070 DVSS.n3715 VSS 0.091242f
C20071 DVSS.n3716 VSS 0.091242f
C20072 DVSS.n3717 VSS 0.091242f
C20073 DVSS.n3718 VSS 0.091242f
C20074 DVSS.n3719 VSS 0.091242f
C20075 DVSS.n3720 VSS 0.091242f
C20076 DVSS.n3721 VSS 0.091242f
C20077 DVSS.n3722 VSS 0.091242f
C20078 DVSS.n3723 VSS 0.091242f
C20079 DVSS.n3724 VSS 0.091242f
C20080 DVSS.n3725 VSS 0.091242f
C20081 DVSS.n3726 VSS 0.046906f
C20082 DVSS.n3727 VSS 0.12011f
C20083 DVSS.n3728 VSS 0.439641f
C20084 DVSS.n3729 VSS 0.082246f
C20085 DVSS.n3730 VSS 0.082246f
C20086 DVSS.n3731 VSS 0.091242f
C20087 DVSS.n3732 VSS 0.091242f
C20088 DVSS.n3733 VSS 0.091242f
C20089 DVSS.n3734 VSS 0.091242f
C20090 DVSS.n3735 VSS 0.091242f
C20091 DVSS.n3736 VSS 0.091242f
C20092 DVSS.n3737 VSS 0.091242f
C20093 DVSS.n3738 VSS 0.091242f
C20094 DVSS.n3739 VSS 0.091242f
C20095 DVSS.n3740 VSS 0.091242f
C20096 DVSS.n3741 VSS 0.091242f
C20097 DVSS.n3742 VSS 0.091242f
C20098 DVSS.n3743 VSS 0.090921f
C20099 DVSS.n3744 VSS 0.104004f
C20100 DVSS.n3745 VSS 0.059799f
C20101 DVSS.n3746 VSS 0.127192f
C20102 DVSS.n3747 VSS 0.059166f
C20103 DVSS.n3748 VSS 0.198298f
C20104 DVSS.n3749 VSS 1.01342f
C20105 DVSS.n3750 VSS 1.18421f
C20106 DVSS.n3751 VSS 0.2064f
C20107 DVSS.t11 VSS 0.320788f
C20108 DVSS.n3752 VSS 0.343618f
C20109 DVSS.n3753 VSS 0.037943f
C20110 DVSS.n3754 VSS 0.070566f
C20111 DVSS.n3755 VSS 0.093424f
C20112 DVSS.n3756 VSS 0.122064f
C20113 DVSS.n3757 VSS 0.021934f
C20114 DVSS.n3758 VSS 0.036157f
C20115 DVSS.n3759 VSS 0.254084f
C20116 DVSS.t27 VSS 0.181488f
C20117 DVSS.t29 VSS 0.220008f
C20118 DVSS.n3760 VSS 0.281711f
C20119 DVSS.t3 VSS 0.220749f
C20120 DVSS.n3761 VSS 0.160844f
C20121 DVSS.t25 VSS 0.226675f
C20122 DVSS.t128 VSS 0.180748f
C20123 DVSS.t115 VSS 0.180748f
C20124 DVSS.t126 VSS 0.214823f
C20125 DVSS.n3762 VSS 0.157533f
C20126 DVSS.t61 VSS 0.009228f
C20127 DVSS.n3763 VSS 0.003762f
C20128 DVSS.n3764 VSS 0.020878f
C20129 DVSS.n3765 VSS 0.009949f
C20130 DVSS.n3766 VSS -0.005431f
C20131 DVSS.n3767 VSS 0.021765f
C20132 DVSS.n3768 VSS 0.01024f
C20133 DVSS.n3769 VSS 0.044918f
C20134 DVSS.n3770 VSS 0.046937f
C20135 DVSS.n3771 VSS 0.069074f
C20136 DVSS.n3772 VSS 0.091242f
C20137 DVSS.n3773 VSS 0.091242f
C20138 DVSS.n3774 VSS 0.091242f
C20139 DVSS.n3775 VSS 0.091242f
C20140 DVSS.n3776 VSS 0.091242f
C20141 DVSS.n3777 VSS 0.091242f
C20142 DVSS.n3778 VSS 0.049155f
C20143 DVSS.n3779 VSS 0.091242f
C20144 DVSS.n3780 VSS 0.091242f
C20145 DVSS.n3781 VSS 0.091242f
C20146 DVSS.n3782 VSS 0.091242f
C20147 DVSS.n3783 VSS 0.091242f
C20148 DVSS.n3784 VSS 0.091242f
C20149 DVSS.n3785 VSS 0.091242f
C20150 DVSS.n3786 VSS 0.058472f
C20151 DVSS.n3787 VSS 0.063027f
C20152 DVSS.n3788 VSS 0.018089f
C20153 DVSS.n3789 VSS 0.158919f
C20154 DVSS.t0 VSS 0.185933f
C20155 DVSS.t16 VSS 0.220008f
C20156 DVSS.t6 VSS 0.220008f
C20157 DVSS.t13 VSS 0.248158f
C20158 DVSS.t31 VSS 0.091114f
C20159 DVSS.n3790 VSS 0.090123f
C20160 DVSS.n3791 VSS -0.005431f
C20161 DVSS.n3792 VSS 0.01024f
C20162 DVSS.n3793 VSS 0.045393f
C20163 DVSS.n3794 VSS 0.046937f
C20164 DVSS.n3795 VSS 0.074857f
C20165 DVSS.n3796 VSS 0.091242f
C20166 DVSS.n3797 VSS 0.091242f
C20167 DVSS.n3798 VSS 0.091242f
C20168 DVSS.n3799 VSS 0.091242f
C20169 DVSS.n3800 VSS 0.091242f
C20170 DVSS.n3801 VSS 0.081925f
C20171 DVSS.n3802 VSS 0.04694f
C20172 DVSS.n3803 VSS 0.054938f
C20173 DVSS.n3804 VSS 0.051083f
C20174 DVSS.n3805 VSS 0.091242f
C20175 DVSS.n3806 VSS 0.091242f
C20176 DVSS.n3807 VSS 0.091242f
C20177 DVSS.n3808 VSS 0.091242f
C20178 DVSS.n3809 VSS 0.091242f
C20179 DVSS.n3810 VSS 0.091242f
C20180 DVSS.n3811 VSS 0.091242f
C20181 DVSS.n3812 VSS 0.091242f
C20182 DVSS.n3813 VSS 0.091242f
C20183 DVSS.n3814 VSS 0.091242f
C20184 DVSS.n3815 VSS 0.091242f
C20185 DVSS.n3816 VSS 0.091242f
C20186 DVSS.n3817 VSS 0.091242f
C20187 DVSS.n3818 VSS 0.091242f
C20188 DVSS.n3819 VSS 0.091242f
C20189 DVSS.n3820 VSS 0.091242f
C20190 DVSS.n3821 VSS 0.091242f
C20191 DVSS.n3822 VSS 0.091242f
C20192 DVSS.n3823 VSS 0.091242f
C20193 DVSS.n3824 VSS 0.091242f
C20194 DVSS.n3825 VSS 0.091242f
C20195 DVSS.n3826 VSS 0.091242f
C20196 DVSS.n3827 VSS 0.091242f
C20197 DVSS.n3828 VSS 0.058472f
C20198 DVSS.n3831 VSS 0.026069f
C20199 DVSS.n3834 VSS 0.026069f
C20200 DVSS.n3837 VSS 0.026069f
C20201 DVSS.n3839 VSS 0.025518f
C20202 DVSS.n3840 VSS 0.045621f
C20203 DVSS.n3841 VSS 0.045621f
C20204 DVSS.n3842 VSS 0.091242f
C20205 DVSS.n3843 VSS 0.091242f
C20206 DVSS.n3844 VSS 0.091242f
C20207 DVSS.n3845 VSS 0.091242f
C20208 DVSS.n3846 VSS 0.091242f
C20209 DVSS.n3847 VSS 0.078391f
C20210 DVSS.n3848 VSS 0.091242f
C20211 DVSS.n3849 VSS 0.091242f
C20212 DVSS.n3850 VSS 0.091242f
C20213 DVSS.n3851 VSS 0.091242f
C20214 DVSS.n3852 VSS 0.091242f
C20215 DVSS.n3853 VSS 0.091242f
C20216 DVSS.n3854 VSS 0.091242f
C20217 DVSS.n3855 VSS 0.0604f
C20218 DVSS.t147 VSS 0.009228f
C20219 DVSS.n3856 VSS 0.003762f
C20220 DVSS.n3857 VSS 0.020878f
C20221 DVSS.n3858 VSS 0.059954f
C20222 DVSS.n3859 VSS 0.072287f
C20223 DVSS.n3860 VSS 0.091242f
C20224 DVSS.n3861 VSS 0.091242f
C20225 DVSS.n3862 VSS 0.091242f
C20226 DVSS.n3863 VSS 0.091242f
C20227 DVSS.n3864 VSS 0.091242f
C20228 DVSS.n3865 VSS 0.091242f
C20229 DVSS.n3866 VSS 0.052368f
C20230 DVSS.n3867 VSS 0.091242f
C20231 DVSS.n3868 VSS 0.091242f
C20232 DVSS.n3869 VSS 0.091242f
C20233 DVSS.n3870 VSS 0.091242f
C20234 DVSS.n3871 VSS 0.091242f
C20235 DVSS.n3872 VSS 0.091242f
C20236 DVSS.n3873 VSS 0.091242f
C20237 DVSS.n3874 VSS 0.058472f
C20238 DVSS.n3875 VSS 0.063027f
C20239 DVSS.n3876 VSS 0.058472f
C20240 DVSS.n3877 VSS 0.059954f
C20241 DVSS.n3878 VSS 0.052368f
C20242 DVSS.n3879 VSS 0.091242f
C20243 DVSS.n3880 VSS 0.091242f
C20244 DVSS.n3881 VSS 0.091242f
C20245 DVSS.n3882 VSS 0.091242f
C20246 DVSS.n3883 VSS 0.091242f
C20247 DVSS.n3884 VSS 0.091242f
C20248 DVSS.n3885 VSS 0.058793f
C20249 DVSS.n3886 VSS 0.059954f
C20250 DVSS.n3887 VSS 0.07807f
C20251 DVSS.n3888 VSS 0.091242f
C20252 DVSS.n3889 VSS 0.091242f
C20253 DVSS.n3890 VSS 0.091242f
C20254 DVSS.n3891 VSS 0.091242f
C20255 DVSS.n3892 VSS 0.091242f
C20256 DVSS.n3893 VSS 0.078712f
C20257 DVSS.n3894 VSS 0.059954f
C20258 DVSS.n3895 VSS 0.020878f
C20259 DVSS.n3896 VSS 0.021765f
C20260 DVSS.n3897 VSS -0.005431f
C20261 DVSS.n3898 VSS 0.009949f
C20262 DVSS.n3899 VSS 0.011819f
C20263 DVSS.n3900 VSS 0.009949f
C20264 DVSS.n3901 VSS -0.005431f
C20265 DVSS.n3902 VSS 0.157533f
C20266 DVSS.t78 VSS 0.149635f
C20267 DVSS.n3903 VSS 0.159475f
C20268 DVSS.n3904 VSS 0.01413f
C20269 DVSS.n3905 VSS 0.057522f
C20270 DVSS.n3906 VSS 0.077749f
C20271 DVSS.n3907 VSS 0.091242f
C20272 DVSS.n3908 VSS 0.091242f
C20273 DVSS.n3909 VSS 0.091242f
C20274 DVSS.n3910 VSS 0.091242f
C20275 DVSS.n3911 VSS 0.091242f
C20276 DVSS.n3912 VSS 0.091242f
C20277 DVSS.n3913 VSS 0.091242f
C20278 DVSS.n3914 VSS 0.091242f
C20279 DVSS.n3915 VSS 0.091242f
C20280 DVSS.n3916 VSS 0.091242f
C20281 DVSS.n3917 VSS 0.091242f
C20282 DVSS.n3918 VSS 0.091242f
C20283 DVSS.n3919 VSS 0.091242f
C20284 DVSS.n3920 VSS 0.091242f
C20285 DVSS.n3921 VSS 0.091242f
C20286 DVSS.n3922 VSS 0.091242f
C20287 DVSS.n3923 VSS 0.091242f
C20288 DVSS.n3924 VSS 0.091242f
C20289 DVSS.n3925 VSS 0.091242f
C20290 DVSS.n3926 VSS 0.091242f
C20291 DVSS.n3927 VSS 0.091242f
C20292 DVSS.n3928 VSS 0.091242f
C20293 DVSS.n3929 VSS 0.091242f
C20294 DVSS.n3930 VSS 0.091242f
C20295 DVSS.n3931 VSS 0.091242f
C20296 DVSS.n3932 VSS 0.091242f
C20297 DVSS.n3933 VSS 0.091242f
C20298 DVSS.n3934 VSS 0.091242f
C20299 DVSS.n3935 VSS 0.091242f
C20300 DVSS.n3936 VSS 0.069074f
C20301 DVSS.n3937 VSS 0.045621f
C20302 DVSS.n3938 VSS 0.222421f
C20303 DVSS.n3939 VSS 0.067217f
C20304 DVSS.n3940 VSS -0.028752f
C20305 DVSS.n3941 VSS 0.02291f
C20306 DVSS.n3942 VSS 1.01501f
C20307 DVSS.n3943 VSS 0.94857f
C20308 DVSS.n3944 VSS 1.26149f
C20309 DVSS.n3945 VSS 0.641625f
C20310 DVSS.n3946 VSS 0.017199f
C20311 DVSS.n3947 VSS 0.172721f
C20312 DVSS.n3948 VSS 0.016261f
C20313 DVSS.n3949 VSS -0.004747f
C20314 DVSS.n3950 VSS 0.551277f
C20315 DVSS.n3951 VSS 0.261545f
C20316 DVSS.n3952 VSS 0.013016f
C20317 DVSS.t47 VSS 0.036785f
C20318 DVSS.n3953 VSS 0.081479f
C20319 DVSS.n3954 VSS 0.126681f
C20320 DVSS.n3955 VSS 0.040888f
C20321 DVSS.n3956 VSS 0.302413f
C20322 DVSS.n3957 VSS 0.195409f
C20323 DVSS.n3958 VSS 0.006702f
C20324 DVSS.n3959 VSS 0.068334f
C20325 DVSS.n3960 VSS 0.156848f
C20326 DVSS.n3961 VSS 0.052427f
C20327 DVSS.n3962 VSS 0.051275f
C20328 DVSS.n3963 VSS 0.051275f
C20329 DVSS.n3964 VSS 0.051275f
C20330 DVSS.n3965 VSS 0.052427f
C20331 DVSS.n3966 VSS 0.168686f
C20332 DVSS.n3967 VSS 0.168686f
C20333 DVSS.n3968 VSS 0.166466f
C20334 DVSS.n3969 VSS 0.168686f
C20335 DVSS.n3970 VSS 0.052427f
C20336 DVSS.n3971 VSS 0.051275f
C20337 DVSS.n3972 VSS 0.051275f
C20338 DVSS.n3973 VSS 0.051275f
C20339 DVSS.n3974 VSS 0.052427f
C20340 DVSS.n3975 VSS 0.085083f
C20341 DVSS.n3976 VSS 0.296566f
C20342 DVSS.n3977 VSS 0.085823f
C20343 DVSS.n3978 VSS 0.24933f
C20344 DVSS.n3979 VSS 0.046908f
C20345 DVSS.n3980 VSS 0.091925f
C20346 DVSS.n3981 VSS 0.389893f
C20347 DVSS.n3982 VSS -0.010233f
C20348 DVSS.n3983 VSS 0.301402f
C20349 DVSS.n3984 VSS 0.741875f
C20350 DVSS.n3985 VSS 1.23012f
C20351 DVSS.n3986 VSS 0.497603f
C20352 DVSS.n3987 VSS -0.129851f
C20353 DVSS.n3988 VSS 0.025757f
C20354 DVSS.n3989 VSS 0.01005f
C20355 DVSS.n3990 VSS 0.011063f
C20356 DVSS.n3991 VSS 0.018241f
C20357 DVSS.n3992 VSS 0.011992f
C20358 DVSS.n3993 VSS 0.018241f
C20359 DVSS.n3994 VSS 0.011992f
C20360 DVSS.n3995 VSS 0.018241f
C20361 DVSS.n3996 VSS 0.018241f
C20362 DVSS.n3997 VSS 0.010556f
C20363 DVSS.n3998 VSS 0.010556f
C20364 DVSS.n3999 VSS 0.018241f
C20365 DVSS.n4000 VSS 0.011992f
C20366 DVSS.n4001 VSS 0.018241f
C20367 DVSS.n4002 VSS 0.018241f
C20368 DVSS.n4003 VSS 0.011992f
C20369 DVSS.n4004 VSS 0.045621f
C20370 DVSS.n4005 VSS 0.091242f
C20371 DVSS.n4006 VSS 0.091242f
C20372 DVSS.n4007 VSS 0.091242f
C20373 DVSS.n4008 VSS 0.091242f
C20374 DVSS.n4009 VSS 0.091242f
C20375 DVSS.n4010 VSS 0.091242f
C20376 DVSS.n4011 VSS 0.091242f
C20377 DVSS.n4012 VSS 0.091242f
C20378 DVSS.n4013 VSS 0.091242f
C20379 DVSS.n4014 VSS 0.091242f
C20380 DVSS.n4015 VSS 0.091242f
C20381 DVSS.n4016 VSS 0.091242f
C20382 DVSS.n4017 VSS 0.091242f
C20383 DVSS.n4018 VSS 0.091242f
C20384 DVSS.n4019 VSS 0.091242f
C20385 DVSS.n4020 VSS 0.091242f
C20386 DVSS.n4021 VSS 0.091242f
C20387 DVSS.n4022 VSS 0.091242f
C20388 DVSS.n4023 VSS 0.091242f
C20389 DVSS.n4024 VSS 0.091242f
C20390 DVSS.n4025 VSS 0.091242f
C20391 DVSS.n4026 VSS 0.091242f
C20392 DVSS.n4027 VSS 0.091242f
C20393 DVSS.n4028 VSS 0.091242f
C20394 DVSS.n4029 VSS 0.091242f
C20395 DVSS.n4030 VSS 0.091242f
C20396 DVSS.n4031 VSS 0.091242f
C20397 DVSS.n4032 VSS 0.091242f
C20398 DVSS.n4033 VSS 0.091242f
C20399 DVSS.n4034 VSS 0.091242f
C20400 DVSS.n4035 VSS 0.046906f
C20401 DVSS.n4036 VSS 0.12011f
C20402 DVSS.n4037 VSS 0.439641f
C20403 DVSS.n4038 VSS 0.082246f
C20404 DVSS.n4039 VSS 0.082246f
C20405 DVSS.n4040 VSS 0.091242f
C20406 DVSS.n4041 VSS 0.091242f
C20407 DVSS.n4042 VSS 0.091242f
C20408 DVSS.n4043 VSS 0.091242f
C20409 DVSS.n4044 VSS 0.091242f
C20410 DVSS.n4045 VSS 0.091242f
C20411 DVSS.n4046 VSS 0.091242f
C20412 DVSS.n4047 VSS 0.091242f
C20413 DVSS.n4048 VSS 0.091242f
C20414 DVSS.n4049 VSS 0.091242f
C20415 DVSS.n4050 VSS 0.091242f
C20416 DVSS.n4051 VSS 0.091242f
C20417 DVSS.n4052 VSS 0.091242f
C20418 DVSS.n4053 VSS 0.091242f
C20419 DVSS.n4054 VSS 0.091242f
C20420 DVSS.n4055 VSS 0.091242f
C20421 DVSS.n4056 VSS 0.091242f
C20422 DVSS.n4057 VSS 0.091242f
C20423 DVSS.n4058 VSS 0.091242f
C20424 DVSS.n4059 VSS 0.091242f
C20425 DVSS.n4060 VSS 0.091242f
C20426 DVSS.n4061 VSS 0.091242f
C20427 DVSS.n4062 VSS 0.091242f
C20428 DVSS.n4063 VSS 0.091242f
C20429 DVSS.n4064 VSS 0.091242f
C20430 DVSS.n4065 VSS 0.091242f
C20431 DVSS.n4066 VSS 0.091242f
C20432 DVSS.n4067 VSS 0.091242f
C20433 DVSS.n4068 VSS 0.091242f
C20434 DVSS.n4069 VSS 0.091242f
C20435 DVSS.n4070 VSS 0.091242f
C20436 DVSS.n4071 VSS 0.091242f
C20437 DVSS.n4072 VSS 0.091242f
C20438 DVSS.n4073 VSS 0.091242f
C20439 DVSS.n4074 VSS 0.091242f
C20440 DVSS.n4075 VSS 0.091242f
C20441 DVSS.n4076 VSS 0.091242f
C20442 DVSS.n4077 VSS 0.091242f
C20443 DVSS.n4078 VSS 0.091242f
C20444 DVSS.n4079 VSS 0.091242f
C20445 DVSS.n4080 VSS 0.091242f
C20446 DVSS.n4081 VSS 0.091242f
C20447 DVSS.n4082 VSS 0.091242f
C20448 DVSS.n4083 VSS 0.091242f
C20449 DVSS.n4084 VSS 0.091242f
C20450 DVSS.n4085 VSS 0.091242f
C20451 DVSS.n4086 VSS 0.091242f
C20452 DVSS.n4087 VSS 0.091242f
C20453 DVSS.n4088 VSS 0.091242f
C20454 DVSS.n4089 VSS 0.091242f
C20455 DVSS.n4090 VSS 0.091242f
C20456 DVSS.n4091 VSS 0.091242f
C20457 DVSS.n4092 VSS 0.049798f
C20458 DVSS.n4093 VSS 0.045621f
C20459 DVSS.n4094 VSS 0.009121f
C20460 DVSS.n4095 VSS 0.045621f
C20461 DVSS.n4096 VSS 0.087066f
C20462 DVSS.n4097 VSS 0.091242f
C20463 DVSS.n4098 VSS 0.091242f
C20464 DVSS.n4099 VSS 0.091242f
C20465 DVSS.n4100 VSS 0.091242f
C20466 DVSS.n4101 VSS 0.091242f
C20467 DVSS.n4102 VSS 0.091242f
C20468 DVSS.n4103 VSS 0.091242f
C20469 DVSS.n4104 VSS 0.091242f
C20470 DVSS.n4105 VSS 0.091242f
C20471 DVSS.n4106 VSS 0.091242f
C20472 DVSS.n4107 VSS 0.091242f
C20473 DVSS.n4108 VSS 0.091242f
C20474 DVSS.n4109 VSS 0.091242f
C20475 DVSS.n4110 VSS 0.091242f
C20476 DVSS.n4111 VSS 0.091242f
C20477 DVSS.n4112 VSS 0.091242f
C20478 DVSS.n4113 VSS 0.091242f
C20479 DVSS.n4114 VSS 0.091242f
C20480 DVSS.n4115 VSS 0.091242f
C20481 DVSS.n4116 VSS 0.091242f
C20482 DVSS.n4117 VSS 0.091242f
C20483 DVSS.n4118 VSS 0.091242f
C20484 DVSS.n4119 VSS 0.091242f
C20485 DVSS.n4120 VSS 0.091242f
C20486 DVSS.n4121 VSS 0.091242f
C20487 DVSS.n4122 VSS 0.091242f
C20488 DVSS.n4123 VSS 0.091242f
C20489 DVSS.n4124 VSS 0.091242f
C20490 DVSS.n4125 VSS 0.091242f
C20491 DVSS.n4126 VSS 0.091242f
C20492 DVSS.n4127 VSS 0.091242f
C20493 DVSS.n4128 VSS 0.091242f
C20494 DVSS.n4129 VSS 0.091242f
C20495 DVSS.n4130 VSS 0.091242f
C20496 DVSS.n4131 VSS 0.091242f
C20497 DVSS.n4132 VSS 0.091242f
C20498 DVSS.n4133 VSS 0.091242f
C20499 DVSS.n4134 VSS 0.091242f
C20500 DVSS.n4135 VSS 0.091242f
C20501 DVSS.n4136 VSS 0.091242f
C20502 DVSS.n4137 VSS 0.091242f
C20503 DVSS.n4138 VSS 0.091242f
C20504 DVSS.n4139 VSS 0.091242f
C20505 DVSS.n4140 VSS 0.091242f
C20506 DVSS.n4141 VSS 0.091242f
C20507 DVSS.n4142 VSS 0.091242f
C20508 DVSS.n4143 VSS 0.091242f
C20509 DVSS.n4144 VSS 0.091242f
C20510 DVSS.n4145 VSS 0.091242f
C20511 DVSS.n4146 VSS 0.091242f
C20512 DVSS.n4147 VSS 0.091242f
C20513 DVSS.n4148 VSS 0.091242f
C20514 DVSS.n4149 VSS 0.091242f
C20515 DVSS.n4150 VSS 0.091242f
C20516 DVSS.n4151 VSS 0.091242f
C20517 DVSS.n4152 VSS 0.091242f
C20518 DVSS.n4153 VSS 0.091242f
C20519 DVSS.n4154 VSS 0.091242f
C20520 DVSS.n4155 VSS 0.091242f
C20521 DVSS.n4156 VSS 0.091242f
C20522 DVSS.n4157 VSS 0.091242f
C20523 DVSS.n4158 VSS 0.091242f
C20524 DVSS.n4159 VSS 0.091242f
C20525 DVSS.n4160 VSS 0.091242f
C20526 DVSS.n4161 VSS 0.091242f
C20527 DVSS.n4162 VSS 0.091242f
C20528 DVSS.n4163 VSS 0.091242f
C20529 DVSS.n4164 VSS 0.091242f
C20530 DVSS.n4165 VSS 0.091242f
C20531 DVSS.n4166 VSS 0.091242f
C20532 DVSS.n4167 VSS 0.085781f
C20533 DVSS.n4168 VSS 0.045621f
C20534 DVSS.n4169 VSS 0.038377f
C20535 DVSS.n4170 VSS 0.044465f
C20536 DVSS.n4171 VSS 0.045621f
C20537 DVSS.n4172 VSS 0.091242f
C20538 DVSS.n4173 VSS 0.091242f
C20539 DVSS.n4174 VSS 0.091242f
C20540 DVSS.n4175 VSS 0.091242f
C20541 DVSS.n4176 VSS 0.091242f
C20542 DVSS.n4177 VSS 0.091242f
C20543 DVSS.n4178 VSS 0.091242f
C20544 DVSS.n4179 VSS 0.063291f
C20545 DVSS.n4180 VSS 0.091242f
C20546 DVSS.n4181 VSS 0.309288f
C20547 DVSS.n4182 VSS 0.041445f
C20548 DVSS.n4183 VSS 1.84602f
C20549 DVSS.n4184 VSS 0.359812f
C20550 DVSS.n4185 VSS 0.009513f
C20551 DVSS.t65 VSS 0.01432f
C20552 DVSS.n4186 VSS 0.038163f
C20553 DVSS.n4187 VSS 0.002529f
C20554 DVSS.n4188 VSS 0.024717f
C20555 DVSS.n4189 VSS 0.584991f
C20556 DVSS.n4190 VSS 3.49018f
C20557 DVSS.n4191 VSS 5.2878f
C20558 DVSS.n4192 VSS 3.96165f
C20559 DVSS.n4193 VSS 0.195519f
C20560 DVSS.n4194 VSS 0.195519f
C20561 DVSS.n4195 VSS 0.195519f
C20562 DVSS.n4196 VSS 0.195519f
C20563 DVSS.n4197 VSS 0.195519f
C20564 DVSS.n4198 VSS 0.195519f
C20565 DVSS.n4199 VSS 0.195519f
C20566 DVSS.n4200 VSS 0.195519f
C20567 DVSS.n4201 VSS 0.195519f
C20568 DVSS.n4202 VSS 0.179685f
C20569 DVSS.n4203 VSS 0.127955f
C20570 DVSS.n4204 VSS 0.113594f
C20571 DVSS.n4205 VSS 0.195519f
C20572 DVSS.n4206 VSS 0.195519f
C20573 DVSS.n4207 VSS 0.195519f
C20574 DVSS.n4208 VSS 0.195519f
C20575 DVSS.n4209 VSS 0.195519f
C20576 DVSS.n4210 VSS 0.195519f
C20577 DVSS.n4211 VSS 0.195519f
C20578 DVSS.n4212 VSS 0.195519f
C20579 DVSS.n4213 VSS 0.113594f
C20580 DVSS.n4214 VSS 0.195519f
C20581 DVSS.n4215 VSS 0.195519f
C20582 DVSS.n4216 VSS 0.195519f
C20583 DVSS.n4217 VSS 0.195519f
C20584 DVSS.n4218 VSS 0.195519f
C20585 DVSS.n4219 VSS 0.195519f
C20586 DVSS.n4220 VSS 0.179685f
C20587 DVSS.n4221 VSS 0.195519f
C20588 DVSS.n4222 VSS 0.195519f
C20589 DVSS.n4223 VSS 0.195519f
C20590 DVSS.n4224 VSS 0.195519f
C20591 DVSS.n4225 VSS 0.195519f
C20592 DVSS.n4226 VSS 0.195519f
C20593 DVSS.n4227 VSS 0.195519f
C20594 DVSS.n4228 VSS 0.195519f
C20595 DVSS.n4229 VSS 0.195519f
C20596 DVSS.n4230 VSS 0.195519f
C20597 DVSS.n4231 VSS 0.195519f
C20598 DVSS.n4232 VSS 0.195519f
C20599 DVSS.n4233 VSS 0.195519f
C20600 DVSS.n4234 VSS 0.195519f
C20601 DVSS.n4235 VSS 0.195519f
C20602 DVSS.n4236 VSS 0.195519f
C20603 DVSS.n4237 VSS 0.11979f
C20604 DVSS.n4238 VSS 0.122398f
C20605 DVSS.n4239 VSS 0.173489f
C20606 DVSS.n4240 VSS 0.195519f
C20607 DVSS.n4241 VSS 0.195519f
C20608 DVSS.n4242 VSS 0.195519f
C20609 DVSS.n4243 VSS 0.195519f
C20610 DVSS.n4244 VSS 0.195519f
C20611 DVSS.n4245 VSS 0.195519f
C20612 DVSS.n4246 VSS 0.195519f
C20613 DVSS.n4247 VSS 0.195519f
C20614 DVSS.n4248 VSS 0.195519f
C20615 DVSS.n4249 VSS 0.195519f
C20616 DVSS.n4250 VSS 0.195519f
C20617 DVSS.n4251 VSS 0.195519f
C20618 DVSS.n4252 VSS 0.195519f
C20619 DVSS.n4253 VSS 0.195519f
C20620 DVSS.n4254 VSS 0.195519f
C20621 DVSS.n4255 VSS 0.195519f
C20622 DVSS.n4256 VSS 0.195519f
C20623 DVSS.n4257 VSS 0.195519f
C20624 DVSS.n4258 VSS 0.195519f
C20625 DVSS.n4259 VSS 0.195519f
C20626 DVSS.n4260 VSS 0.195519f
C20627 DVSS.n4261 VSS 0.195519f
C20628 DVSS.n4262 VSS 0.195519f
C20629 DVSS.n4263 VSS 0.195519f
C20630 DVSS.n4264 VSS 0.195519f
C20631 DVSS.n4265 VSS 0.195519f
C20632 DVSS.n4266 VSS 0.195519f
C20633 DVSS.n4267 VSS 0.195519f
C20634 DVSS.n4268 VSS 0.195519f
C20635 DVSS.n4269 VSS 0.195519f
C20636 DVSS.n4270 VSS 0.195519f
C20637 DVSS.n4271 VSS 0.195519f
C20638 DVSS.n4272 VSS 0.195519f
C20639 DVSS.n4273 VSS 0.195519f
C20640 DVSS.n4274 VSS 0.195519f
C20641 DVSS.n4275 VSS 0.195519f
C20642 DVSS.n4276 VSS 0.195519f
C20643 DVSS.n4277 VSS 0.195519f
C20644 DVSS.n4278 VSS 0.195519f
C20645 DVSS.n4279 VSS 0.195519f
C20646 DVSS.n4280 VSS 0.195519f
C20647 DVSS.n4281 VSS 0.195519f
C20648 DVSS.n4282 VSS 0.195519f
C20649 DVSS.n4283 VSS 0.195519f
C20650 DVSS.n4284 VSS 0.195519f
C20651 DVSS.n4285 VSS 0.195519f
C20652 DVSS.n4286 VSS 0.195519f
C20653 DVSS.n4287 VSS 0.195519f
C20654 DVSS.n4288 VSS 0.195519f
C20655 DVSS.n4289 VSS 0.195519f
C20656 DVSS.n4290 VSS 0.195519f
C20657 DVSS.n4291 VSS 0.195519f
C20658 DVSS.n4292 VSS 0.195519f
C20659 DVSS.n4293 VSS 0.195519f
C20660 DVSS.n4294 VSS 0.195519f
C20661 DVSS.n4295 VSS 0.195519f
C20662 DVSS.n4296 VSS 0.195519f
C20663 DVSS.n4297 VSS 0.195519f
C20664 DVSS.n4298 VSS 0.195519f
C20665 DVSS.n4299 VSS 0.195519f
C20666 DVSS.n4300 VSS 0.195519f
C20667 DVSS.n4301 VSS 0.195519f
C20668 DVSS.n4302 VSS 0.195519f
C20669 DVSS.n4303 VSS 0.195519f
C20670 DVSS.n4304 VSS 0.195519f
C20671 DVSS.n4305 VSS 0.195519f
C20672 DVSS.n4306 VSS 0.195519f
C20673 DVSS.n4307 VSS 0.104332f
C20674 DVSS.n4308 VSS 0.195519f
C20675 DVSS.n4309 VSS 0.195519f
C20676 DVSS.n4310 VSS 0.195519f
C20677 DVSS.n4311 VSS 0.195519f
C20678 DVSS.n4312 VSS 0.195519f
C20679 DVSS.n4313 VSS 0.195519f
C20680 DVSS.n4314 VSS 0.195519f
C20681 DVSS.n4315 VSS 0.195519f
C20682 DVSS.n4316 VSS 0.195519f
C20683 DVSS.n4317 VSS 0.195519f
C20684 DVSS.n4318 VSS 0.195519f
C20685 DVSS.n4319 VSS 0.195519f
C20686 DVSS.n4320 VSS 0.195519f
C20687 DVSS.n4321 VSS 0.195519f
C20688 DVSS.n4322 VSS 0.195519f
C20689 DVSS.n4323 VSS 0.195519f
C20690 DVSS.n4324 VSS 0.195519f
C20691 DVSS.n4325 VSS 0.195519f
C20692 DVSS.n4326 VSS 0.195519f
C20693 DVSS.n4327 VSS 0.195519f
C20694 DVSS.n4328 VSS 0.195519f
C20695 DVSS.n4329 VSS 0.195519f
C20696 DVSS.n4330 VSS 0.176242f
C20697 DVSS.n4331 VSS 0.195519f
C20698 DVSS.n4332 VSS 0.195519f
C20699 DVSS.n4333 VSS 0.176242f
C20700 DVSS.n4334 VSS 0.192765f
C20701 DVSS.n4335 VSS 0.02203f
C20702 DVSS.n4336 VSS 0.009474f
C20703 DVSS.t149 VSS 0.01432f
C20704 DVSS.n4337 VSS 0.038163f
C20705 DVSS.n4338 VSS 0.002529f
C20706 DVSS.n4339 VSS 0.031738f
C20707 DVSS.n4340 VSS 0.125268f
C20708 DVSS.n4341 VSS 0.037865f
C20709 DVSS.n4342 VSS 0.117036f
C20710 DVSS.n4343 VSS 0.176242f
C20711 DVSS.n4344 VSS 0.195519f
C20712 DVSS.n4345 VSS 0.195519f
C20713 DVSS.n4346 VSS 0.195519f
C20714 DVSS.n4347 VSS 0.195519f
C20715 DVSS.n4348 VSS 0.195519f
C20716 DVSS.n4349 VSS 0.195519f
C20717 DVSS.n4350 VSS 0.195519f
C20718 DVSS.n4351 VSS 0.195519f
C20719 DVSS.n4352 VSS 0.195519f
C20720 DVSS.n4353 VSS 0.195519f
C20721 DVSS.n4354 VSS 0.195519f
C20722 DVSS.n4355 VSS 0.195519f
C20723 DVSS.n4356 VSS 0.195519f
C20724 DVSS.n4357 VSS 0.195519f
C20725 DVSS.n4358 VSS 0.195519f
C20726 DVSS.n4359 VSS 0.195519f
C20727 DVSS.n4360 VSS 0.195519f
C20728 DVSS.n4361 VSS 0.195519f
C20729 DVSS.n4362 VSS 0.195519f
C20730 DVSS.n4363 VSS 0.195519f
C20731 DVSS.n4364 VSS 0.195519f
C20732 DVSS.n4365 VSS 0.145262f
C20733 DVSS.n4366 VSS 0.195519f
C20734 DVSS.n4367 VSS 0.195519f
C20735 DVSS.n4368 VSS 0.148016f
C20736 DVSS.n4369 VSS 0.195519f
C20737 DVSS.n4370 VSS 0.195519f
C20738 DVSS.n4371 VSS 0.195519f
C20739 DVSS.n4372 VSS 0.195519f
C20740 DVSS.n4373 VSS 0.195519f
C20741 DVSS.n4374 VSS 0.195519f
C20742 DVSS.n4375 VSS 0.176931f
C20743 DVSS.n4376 VSS 0.078155f
C20744 DVSS.n4377 VSS 0.024973f
C20745 DVSS.n4378 VSS 0.02385f
C20746 DVSS.t191 VSS 0.01432f
C20747 DVSS.t170 VSS 0.01432f
C20748 DVSS.n4379 VSS 0.032399f
C20749 DVSS.n4380 VSS 0.020154f
C20750 DVSS.t37 VSS 0.546681f
C20751 DVSS.n4381 VSS 0.081457f
C20752 DVSS.n4382 VSS 0.02385f
C20753 DVSS.t99 VSS 0.249187f
C20754 DVSS.n4383 VSS 0.637612f
C20755 DVSS.t32 VSS 0.574145f
C20756 DVSS.n4384 VSS 0.123308f
C20757 DVSS.n4385 VSS 0.031885f
C20758 DVSS.n4386 VSS 0.059647f
C20759 DVSS.n4387 VSS 0.031885f
C20760 DVSS.n4388 VSS 0.123308f
C20761 DVSS.n4389 VSS 0.677268f
C20762 DVSS.t98 VSS 0.306125f
C20763 DVSS.t188 VSS 0.342298f
C20764 DVSS.n4390 VSS 0.018264f
C20765 DVSS.n4391 VSS 0.002529f
C20766 DVSS.t189 VSS 0.01432f
C20767 DVSS.n4392 VSS 0.038163f
C20768 DVSS.n4393 VSS 0.009513f
C20769 DVSS.n4394 VSS 0.035564f
C20770 DVSS.t201 VSS 0.01432f
C20771 DVSS.t121 VSS 0.01432f
C20772 DVSS.n4395 VSS 0.032655f
C20773 DVSS.n4396 VSS 0.011953f
C20774 DVSS.t193 VSS 0.01432f
C20775 DVSS.t206 VSS 0.014215f
C20776 DVSS.n4397 VSS 0.026627f
C20777 DVSS.n4398 VSS 0.018226f
C20778 DVSS.t140 VSS 0.01432f
C20779 DVSS.n4399 VSS 0.028639f
C20780 DVSS.n4400 VSS 0.011953f
C20781 DVSS.n4401 VSS 0.023915f
C20782 DVSS.n4402 VSS 0.025288f
C20783 DVSS.n4403 VSS -0.047331f
C20784 DVSS.n4404 VSS 0.166583f
C20785 DVSS.t169 VSS 0.326891f
C20786 DVSS.t190 VSS 0.263254f
C20787 DVSS.n4405 VSS 0.163445f
C20788 DVSS.n4406 VSS 0.046383f
C20789 DVSS.n4407 VSS 0.020849f
C20790 DVSS.n4408 VSS 0.024973f
C20791 DVSS.n4409 VSS 0.092382f
C20792 DVSS.n4410 VSS 0.023355f
C20793 DVSS.n4411 VSS 0.127955f
C20794 DVSS.n4412 VSS 0.116347f
C20795 DVSS.n4413 VSS 0.195519f
C20796 DVSS.n4414 VSS 0.195519f
C20797 DVSS.n4415 VSS 0.195519f
C20798 DVSS.n4416 VSS 0.195519f
C20799 DVSS.n4417 VSS 0.195519f
C20800 DVSS.n4418 VSS 0.195519f
C20801 DVSS.n4419 VSS 0.195519f
C20802 DVSS.n4420 VSS 0.195519f
C20803 DVSS.n4421 VSS 0.195519f
C20804 DVSS.n4422 VSS 0.11084f
C20805 DVSS.n4423 VSS 0.125268f
C20806 DVSS.n4424 VSS 0.031738f
C20807 DVSS.t151 VSS 0.01432f
C20808 DVSS.n4425 VSS 0.002529f
C20809 DVSS.n4426 VSS 0.038163f
C20810 DVSS.n4427 VSS 0.009513f
C20811 DVSS.n4428 VSS 0.035564f
C20812 DVSS.n4429 VSS -0.047331f
C20813 DVSS.n4430 VSS 0.210794f
C20814 DVSS.t171 VSS 0.326891f
C20815 DVSS.t152 VSS 0.263254f
C20816 DVSS.t150 VSS 0.256556f
C20817 DVSS.n4431 VSS 0.163445f
C20818 DVSS.n4432 VSS 0.046383f
C20819 DVSS.t204 VSS 0.325551f
C20820 DVSS.t111 VSS 0.245168f
C20821 DVSS.t83 VSS 0.23646f
C20822 DVSS.t109 VSS 0.326891f
C20823 DVSS.t113 VSS 0.245168f
C20824 DVSS.n4433 VSS 0.163446f
C20825 DVSS.n4434 VSS 0.049341f
C20826 DVSS.n4435 VSS 0.026627f
C20827 DVSS.n4436 VSS 0.018226f
C20828 DVSS.t114 VSS 0.01432f
C20829 DVSS.n4437 VSS 0.028639f
C20830 DVSS.n4438 VSS 0.011953f
C20831 DVSS.n4439 VSS 0.023915f
C20832 DVSS.t205 VSS 0.01432f
C20833 DVSS.n4440 VSS 0.038163f
C20834 DVSS.n4441 VSS 0.0119f
C20835 DVSS.n4442 VSS 0.010771f
C20836 DVSS.n4443 VSS 0.027526f
C20837 DVSS.n4444 VSS 0.092451f
C20838 DVSS.n4445 VSS 0.320192f
C20839 DVSS.t70 VSS 0.391867f
C20840 DVSS.n4446 VSS 0.193152f
C20841 DVSS.t74 VSS 0.056178f
C20842 DVSS.n4447 VSS 0.118198f
C20843 DVSS.n4448 VSS 0.002205f
C20844 DVSS.t91 VSS 0.00716f
C20845 DVSS.t182 VSS 0.00716f
C20846 DVSS.n4449 VSS 0.014896f
C20847 DVSS.n4450 VSS 0.006708f
C20848 DVSS.n4451 VSS 0.010442f
C20849 DVSS.n4452 VSS 0.019198f
C20850 DVSS.n4453 VSS 0.050086f
C20851 DVSS.n4454 VSS 0.249904f
C20852 DVSS.t85 VSS 0.384538f
C20853 DVSS.t165 VSS 0.271177f
C20854 DVSS.t138 VSS 0.204494f
C20855 DVSS.n4455 VSS 0.173767f
C20856 DVSS.n4456 VSS 0.00233f
C20857 DVSS.n4457 VSS 0.257173f
C20858 DVSS.t66 VSS 0.16893f
C20859 DVSS.n4458 VSS 0.271177f
C20860 DVSS.n4459 VSS 0.046383f
C20861 DVSS.n4460 VSS 0.020849f
C20862 DVSS.n4461 VSS 0.024973f
C20863 DVSS.n4462 VSS 0.092382f
C20864 DVSS.n4463 VSS 0.024973f
C20865 DVSS.n4464 VSS 0.020849f
C20866 DVSS.n4465 VSS 0.046383f
C20867 DVSS.n4466 VSS 0.181155f
C20868 DVSS.n4467 VSS 0.29808f
C20869 DVSS.t202 VSS 0.331191f
C20870 DVSS.t176 VSS 0.009228f
C20871 DVSS.n4468 VSS 0.009531f
C20872 DVSS.t2 VSS 0.00358f
C20873 DVSS.t178 VSS 0.00358f
C20874 DVSS.n4469 VSS 0.007228f
C20875 DVSS.n4470 VSS 0.006574f
C20876 DVSS.n4471 VSS 0.258416f
C20877 DVSS.t130 VSS 0.154482f
C20878 DVSS.n4472 VSS 0.271177f
C20879 DVSS.t159 VSS 0.238947f
C20880 DVSS.t56 VSS 0.271177f
C20881 DVSS.t163 VSS 0.271177f
C20882 DVSS.t1 VSS 0.236724f
C20883 DVSS.t199 VSS 0.271177f
C20884 DVSS.t177 VSS 0.271177f
C20885 DVSS.t101 VSS 0.137811f
C20886 DVSS.n4473 VSS 0.142663f
C20887 DVSS.t57 VSS 0.009228f
C20888 DVSS.n4474 VSS 0.009531f
C20889 DVSS.n4475 VSS 0.012036f
C20890 DVSS.n4476 VSS -0.004569f
C20891 DVSS.n4477 VSS 0.027295f
C20892 DVSS.n4478 VSS 0.253676f
C20893 DVSS.t167 VSS 0.301184f
C20894 DVSS.n4479 VSS 0.291109f
C20895 DVSS.n4480 VSS -0.047331f
C20896 DVSS.n4481 VSS 0.025288f
C20897 DVSS.n4482 VSS 0.018531f
C20898 DVSS.n4483 VSS 0.080873f
C20899 DVSS.n4484 VSS 0.028014f
C20900 DVSS.n4485 VSS 0.112316f
C20901 DVSS.n4486 VSS 0.435662f
C20902 DVSS.n4487 VSS 2.18931f
C20903 DVSS.n4488 VSS 0.704323f
C20904 DVSS.n4489 VSS 2.80051f
C20905 DVSS.n4490 VSS 1.4099f
C20906 DVSS.n4491 VSS 2.33847f
C20907 DVSS.n4492 VSS 0.068367f
C20908 DVSS.n4493 VSS 0.257333f
C20909 DVSS.n4494 VSS 0.023334f
C20910 DVSS.n4495 VSS 0.026721f
C20911 DVSS.n4496 VSS 0.045621f
C20912 DVSS.n4497 VSS 0.045621f
C20913 DVSS.n4498 VSS 0.091242f
C20914 DVSS.n4499 VSS 0.091242f
C20915 DVSS.n4500 VSS 0.091242f
C20916 DVSS.n4501 VSS 0.091242f
C20917 DVSS.n4502 VSS 0.045621f
C20918 DVSS.n4503 VSS 0.042127f
C20919 DVSS.n4504 VSS 0.061042f
C20920 DVSS.n4505 VSS 0.045621f
C20921 DVSS.n4506 VSS 0.091242f
C20922 DVSS.n4507 VSS 0.091242f
C20923 DVSS.n4508 VSS 0.091242f
C20924 DVSS.n4509 VSS 0.045621f
C20925 DVSS.n4510 VSS 0.091242f
C20926 DVSS.n4511 VSS 0.978121f
C20927 DVSS.n4513 VSS 0.026069f
C20928 DVSS.n4515 VSS 0.026069f
C20929 DVSS.n4517 VSS 0.026069f
C20930 DVSS.n4519 VSS 0.026069f
C20931 DVSS.n4521 VSS 0.026069f
C20932 DVSS.n4523 VSS 0.026069f
C20933 DVSS.n4525 VSS 0.016706f
C20934 DVSS.n4527 VSS 0.020011f
C20935 DVSS.n4528 VSS 1.47754f
C20936 DVSS.n4529 VSS 0.038017f
C20937 DVSS.n4532 VSS 0.022765f
C20938 DVSS.n4534 VSS 0.022765f
C20939 DVSS.n4535 VSS 0.065916f
C20940 DVSS.n4536 VSS 0.028456f
C20941 DVSS.n4537 VSS 0.085385f
C20942 DVSS.n4538 VSS 0.013035f
C20943 DVSS.n4539 VSS 0.011382f
C20944 DVSS.n4540 VSS 0.045621f
C20945 DVSS.n4541 VSS 0.026069f
C20946 DVSS.n4543 VSS 0.024233f
C20947 DVSS.n4544 VSS 0.044465f
C20948 DVSS.n4545 VSS 0.045621f
C20949 DVSS.n4546 VSS 0.271007f
C20950 DVSS.n4547 VSS 1.46646f
C20951 DVSS.n4548 VSS 1.0806f
C20952 DVSS.n4549 VSS 0.091242f
C20953 DVSS.n4550 VSS 0.091242f
C20954 DVSS.n4551 VSS 0.073251f
C20955 DVSS.n4552 VSS 0.091242f
C20956 DVSS.n4553 VSS 0.091242f
C20957 DVSS.n4554 VSS 0.091242f
C20958 DVSS.n4555 VSS 0.091242f
C20959 DVSS.n4556 VSS 0.091242f
C20960 DVSS.n4557 VSS 0.091242f
C20961 DVSS.n4558 VSS 0.091242f
C20962 DVSS.n4559 VSS 0.045621f
C20963 DVSS.n4560 VSS 0.045803f
C20964 DVSS.n4561 VSS 0.051321f
C20965 DVSS.n4562 VSS 0.251763f
C20966 DVSS.n4563 VSS 0.026721f
C20967 DVSS.n4564 VSS 0.026721f
C20968 DVSS.n4565 VSS 0.023334f
C20969 DVSS.n4566 VSS 0.045621f
C20970 DVSS.n4567 VSS 0.045621f
C20971 DVSS.n4568 VSS 0.045621f
C20972 DVSS.n4569 VSS 0.091242f
C20973 DVSS.n4570 VSS 0.091242f
C20974 DVSS.n4571 VSS 0.091242f
C20975 DVSS.n4572 VSS 0.091242f
C20976 DVSS.n4573 VSS 0.091242f
C20977 DVSS.n4574 VSS 0.045621f
C20978 DVSS.n4575 VSS 0.042127f
C20979 DVSS.n4576 VSS 0.051508f
C20980 DVSS.n4577 VSS 0.045803f
C20981 DVSS.n4578 VSS 0.091242f
C20982 DVSS.n4579 VSS 0.091242f
C20983 DVSS.n4580 VSS 0.091242f
C20984 DVSS.n4581 VSS 0.091242f
C20985 DVSS.n4582 VSS 0.045621f
C20986 DVSS.n4583 VSS 0.251763f
C20987 DVSS.n4584 VSS 0.026721f
C20988 DVSS.n4585 VSS 0.045621f
C20989 DVSS.n4586 VSS 0.091242f
C20990 DVSS.n4587 VSS 0.091242f
C20991 DVSS.n4588 VSS 0.091242f
C20992 DVSS.n4589 VSS 0.091242f
C20993 DVSS.n4590 VSS 0.091242f
C20994 DVSS.n4591 VSS 0.045621f
C20995 DVSS.n4592 VSS 0.045621f
C20996 DVSS.n4593 VSS 0.045621f
C20997 DVSS.n4594 VSS 0.026721f
C20998 DVSS.n4595 VSS 0.042127f
C20999 DVSS.n4596 VSS 0.023334f
C21000 DVSS.n4597 VSS 0.023334f
C21001 DVSS.n4598 VSS 0.026721f
C21002 DVSS.n4599 VSS 0.068367f
C21003 DVSS.n4600 VSS 0.044619f
C21004 DVSS.n4601 VSS 0.065489f
C21005 DVSS.n4602 VSS 0.045621f
C21006 DVSS.n4603 VSS 0.045621f
C21007 DVSS.n4604 VSS 0.091242f
C21008 DVSS.n4605 VSS 0.091242f
C21009 DVSS.n4606 VSS 0.091242f
C21010 DVSS.n4607 VSS 0.091242f
C21011 DVSS.n4608 VSS 0.091242f
C21012 DVSS.n4609 VSS 0.091242f
C21013 DVSS.n4610 VSS 0.091242f
C21014 DVSS.n4611 VSS 0.091242f
C21015 DVSS.n4612 VSS 0.091242f
C21016 DVSS.n4613 VSS 0.091242f
C21017 DVSS.n4614 VSS 0.045621f
C21018 DVSS.n4615 VSS 0.026721f
C21019 DVSS.n4616 VSS 0.045621f
C21020 DVSS.n4617 VSS 0.045621f
C21021 DVSS.n4618 VSS 0.042127f
C21022 DVSS.n4619 VSS 0.051321f
C21023 DVSS.n4620 VSS 0.045803f
C21024 DVSS.n4621 VSS 0.056223f
C21025 DVSS.n4622 VSS 0.091242f
C21026 DVSS.n4623 VSS 0.091242f
C21027 DVSS.n4624 VSS 0.091242f
C21028 DVSS.n4625 VSS 0.091242f
C21029 DVSS.n4626 VSS 0.091242f
C21030 DVSS.n4627 VSS 0.091242f
C21031 DVSS.n4628 VSS 0.091242f
C21032 DVSS.n4629 VSS 0.091242f
C21033 DVSS.n4630 VSS 0.091242f
C21034 DVSS.n4631 VSS 0.091242f
C21035 DVSS.n4632 VSS 0.091242f
C21036 DVSS.n4633 VSS 0.091242f
C21037 DVSS.n4634 VSS 0.091242f
C21038 DVSS.n4635 VSS 0.055902f
C21039 DVSS.n4636 VSS 0.045803f
C21040 DVSS.n4637 VSS 0.051508f
C21041 DVSS.n4638 VSS 0.257333f
C21042 DVSS.n4639 VSS 0.026721f
C21043 DVSS.n4640 VSS 0.023334f
C21044 DVSS.n4641 VSS 0.045621f
C21045 DVSS.n4642 VSS 0.045621f
C21046 DVSS.n4643 VSS 0.091242f
C21047 DVSS.n4644 VSS 0.091242f
C21048 DVSS.n4645 VSS 0.091242f
C21049 DVSS.n4646 VSS 0.091242f
C21050 DVSS.n4647 VSS 0.091242f
C21051 DVSS.n4648 VSS 0.045621f
C21052 DVSS.n4649 VSS 0.045621f
C21053 DVSS.n4650 VSS 0.042127f
C21054 DVSS.n4651 VSS 0.051321f
C21055 DVSS.n4652 VSS 0.045803f
C21056 DVSS.n4653 VSS 0.080961f
C21057 DVSS.n4654 VSS 0.091242f
C21058 DVSS.n4655 VSS 0.091242f
C21059 DVSS.n4656 VSS 0.091242f
C21060 DVSS.n4657 VSS 0.091242f
C21061 DVSS.n4658 VSS 0.091242f
C21062 DVSS.n4659 VSS 0.091242f
C21063 DVSS.n4660 VSS 0.091242f
C21064 DVSS.n4661 VSS 0.091242f
C21065 DVSS.n4662 VSS 0.075821f
C21066 DVSS.n4663 VSS 0.091242f
C21067 DVSS.n4664 VSS 0.091242f
C21068 DVSS.n4665 VSS 0.091242f
C21069 DVSS.n4666 VSS 0.091242f
C21070 DVSS.n4667 VSS 0.091242f
C21071 DVSS.n4668 VSS 0.045621f
C21072 DVSS.n4669 VSS 0.045621f
C21073 DVSS.n4670 VSS 0.023334f
C21074 DVSS.n4671 VSS 0.026721f
C21075 DVSS.n4672 VSS 0.065489f
C21076 DVSS.n4673 VSS 0.044619f
C21077 DVSS.n4674 VSS 1.29078f
C21078 DVSS.n4675 VSS 1.99722f
C21079 DVSS.n4676 VSS 2.04346f
C21080 DVSS.n4677 VSS 2.0452f
C21081 DVSS.n4678 VSS 1.32179f
C21082 DVSS.n4679 VSS 0.044619f
C21083 DVSS.n4680 VSS 0.068367f
C21084 DVSS.n4681 VSS 0.026721f
C21085 DVSS.n4682 VSS 0.023334f
C21086 DVSS.n4683 VSS 0.045621f
C21087 DVSS.n4684 VSS 0.045621f
C21088 DVSS.n4685 VSS 0.091242f
C21089 DVSS.n4686 VSS 0.091242f
C21090 DVSS.n4687 VSS 0.091242f
C21091 DVSS.n4688 VSS 0.091242f
C21092 DVSS.n4689 VSS 0.091242f
C21093 DVSS.n4690 VSS 0.045621f
C21094 DVSS.n4691 VSS 0.045621f
C21095 DVSS.n4692 VSS 0.023334f
C21096 DVSS.n4693 VSS 0.026721f
C21097 DVSS.n4694 VSS 0.257333f
C21098 DVSS.n4695 VSS 0.051508f
C21099 DVSS.n4696 VSS 0.045803f
C21100 DVSS.n4697 VSS 0.08064f
C21101 DVSS.n4698 VSS 0.091242f
C21102 DVSS.n4699 VSS 0.091242f
C21103 DVSS.n4700 VSS 0.091242f
C21104 DVSS.n4701 VSS 0.091242f
C21105 DVSS.n4702 VSS 0.091242f
C21106 DVSS.n4703 VSS 0.091242f
C21107 DVSS.n4704 VSS 0.091242f
C21108 DVSS.n4705 VSS 0.077106f
C21109 DVSS.n4706 VSS 0.091242f
C21110 DVSS.n4707 VSS 0.091242f
C21111 DVSS.n4708 VSS 0.091242f
C21112 DVSS.n4709 VSS 0.091242f
C21113 DVSS.n4710 VSS 0.091242f
C21114 DVSS.n4711 VSS 0.091242f
C21115 DVSS.n4712 VSS 0.045621f
C21116 DVSS.n4713 VSS 0.045621f
C21117 DVSS.n4714 VSS 0.045621f
C21118 DVSS.n4715 VSS 0.042127f
C21119 DVSS.n4716 VSS 0.026721f
C21120 DVSS.n4717 VSS 0.251763f
C21121 DVSS.n4718 VSS 0.044619f
C21122 DVSS.n4719 VSS 0.068367f
C21123 DVSS.n4720 VSS 0.026721f
C21124 DVSS.n4721 VSS 0.023334f
C21125 DVSS.n4722 VSS 0.045621f
C21126 DVSS.n4723 VSS 0.045621f
C21127 DVSS.n4724 VSS 0.091242f
C21128 DVSS.n4725 VSS 0.091242f
C21129 DVSS.n4726 VSS 0.091242f
C21130 DVSS.n4727 VSS 0.091242f
C21131 DVSS.n4728 VSS 0.091242f
C21132 DVSS.n4729 VSS 0.091242f
C21133 DVSS.n4730 VSS 0.045621f
C21134 DVSS.n4731 VSS 0.045621f
C21135 DVSS.n4732 VSS 0.023334f
C21136 DVSS.n4733 VSS 0.026721f
C21137 DVSS.n4734 VSS 0.257333f
C21138 DVSS.n4735 VSS 0.051508f
C21139 DVSS.n4736 VSS 0.045803f
C21140 DVSS.n4737 VSS 0.059757f
C21141 DVSS.n4738 VSS 0.091242f
C21142 DVSS.n4739 VSS 0.091242f
C21143 DVSS.n4740 VSS 0.091242f
C21144 DVSS.n4741 VSS 0.091242f
C21145 DVSS.n4742 VSS 0.091242f
C21146 DVSS.n4743 VSS 0.091242f
C21147 DVSS.n4744 VSS 0.091242f
C21148 DVSS.n4745 VSS 0.091242f
C21149 DVSS.n4746 VSS 0.091242f
C21150 DVSS.n4747 VSS 0.091242f
C21151 DVSS.n4748 VSS 0.091242f
C21152 DVSS.n4749 VSS 0.091242f
C21153 DVSS.n4750 VSS 0.091242f
C21154 DVSS.n4751 VSS 0.091242f
C21155 DVSS.n4752 VSS 0.045621f
C21156 DVSS.n4753 VSS 0.045803f
C21157 DVSS.n4754 VSS 0.051321f
C21158 DVSS.n4755 VSS 0.251763f
C21159 DVSS.n4756 VSS 0.026721f
C21160 DVSS.n4757 VSS 0.026721f
C21161 DVSS.n4758 VSS 0.023334f
C21162 DVSS.n4759 VSS 0.045621f
C21163 DVSS.n4760 VSS 0.045621f
C21164 DVSS.n4761 VSS 0.045621f
C21165 DVSS.n4762 VSS 0.091242f
C21166 DVSS.n4763 VSS 0.091242f
C21167 DVSS.n4764 VSS 0.091242f
C21168 DVSS.n4765 VSS 0.091242f
C21169 DVSS.n4766 VSS 0.091242f
C21170 DVSS.n4767 VSS 0.045621f
C21171 DVSS.n4768 VSS 0.042127f
C21172 DVSS.n4769 VSS 0.051508f
C21173 DVSS.n4770 VSS 0.045803f
C21174 DVSS.n4771 VSS 0.091242f
C21175 DVSS.n4772 VSS 0.091242f
C21176 DVSS.n4773 VSS 0.091242f
C21177 DVSS.n4774 VSS 0.091242f
C21178 DVSS.n4775 VSS 0.045621f
C21179 DVSS.n4776 VSS 0.251763f
C21180 DVSS.n4777 VSS 0.026721f
C21181 DVSS.n4778 VSS 0.045621f
C21182 DVSS.n4779 VSS 0.091242f
C21183 DVSS.n4780 VSS 0.091242f
C21184 DVSS.n4781 VSS 0.091242f
C21185 DVSS.n4782 VSS 0.091242f
C21186 DVSS.n4783 VSS 0.091242f
C21187 DVSS.n4784 VSS 0.045621f
C21188 DVSS.n4785 VSS 0.045621f
C21189 DVSS.n4786 VSS 0.045621f
C21190 DVSS.n4787 VSS 0.026721f
C21191 DVSS.n4788 VSS 0.042127f
C21192 DVSS.n4789 VSS 0.023334f
C21193 DVSS.n4790 VSS 0.023334f
C21194 DVSS.n4791 VSS 0.026721f
C21195 DVSS.n4792 VSS 0.068367f
C21196 DVSS.n4793 VSS 0.044619f
C21197 DVSS.n4794 VSS 0.065489f
C21198 DVSS.n4795 VSS 0.045621f
C21199 DVSS.n4796 VSS 0.045621f
C21200 DVSS.n4797 VSS 0.091242f
C21201 DVSS.n4798 VSS 0.091242f
C21202 DVSS.n4799 VSS 0.091242f
C21203 DVSS.n4800 VSS 0.091242f
C21204 DVSS.n4801 VSS 0.091242f
C21205 DVSS.n4802 VSS 0.091242f
C21206 DVSS.n4803 VSS 0.026069f
C21207 DVSS.n4804 VSS 0.026069f
C21208 DVSS.n4805 VSS 0.026069f
C21209 DVSS.n4806 VSS 0.026069f
C21210 DVSS.n4807 VSS 0.011382f
C21211 DVSS.n4808 VSS 0.045621f
C21212 DVSS.n4810 VSS 0.022765f
C21213 DVSS.n4812 VSS 0.022765f
C21214 DVSS.n4814 VSS 0.038017f
C21215 DVSS.n4815 VSS 0.016706f
C21216 DVSS.n4817 VSS 0.071742f
C21217 DVSS.n4819 VSS 0.028456f
C21218 DVSS.n4820 VSS 0.082472f
C21219 DVSS.n4821 VSS 0.013035f
C21220 DVSS.n4822 VSS 0.020011f
C21221 DVSS.n4823 VSS 0.026069f
C21222 DVSS.n4824 VSS 0.026069f
C21223 DVSS.n4825 VSS 0.026069f
C21224 DVSS.n4830 VSS 0.044465f
C21225 DVSS.n4831 VSS 0.045621f
C21226 DVSS.n4835 VSS 0.091242f
C21227 DVSS.n4836 VSS 0.091242f
C21228 DVSS.n4837 VSS 0.091242f
C21229 DVSS.n4838 VSS 0.091242f
C21230 DVSS.n4839 VSS 0.091242f
C21231 DVSS.n4840 VSS 0.091242f
C21232 DVSS.n4841 VSS 0.091242f
C21233 DVSS.n4842 VSS 0.091242f
C21234 DVSS.n4843 VSS 0.091242f
C21235 DVSS.n4844 VSS 0.091242f
C21236 DVSS.n4845 VSS 0.046906f
C21237 DVSS.n4846 VSS 0.091242f
C21238 DVSS.n4847 VSS 0.089957f
C21239 DVSS.n4848 VSS 0.047098f
C21240 DVSS.n4849 VSS 0.340567f
C21241 DVSS.n4850 VSS 0.174165f
C21242 DVSS.n4851 VSS 0.091242f
C21243 DVSS.n4852 VSS 0.051404f
C21244 DVSS.n4853 VSS 0.091242f
C21245 DVSS.n4854 VSS 0.058151f
C21246 DVSS.n4855 VSS 0.091242f
C21247 DVSS.n4856 VSS 0.041604f
C21248 DVSS.n4857 VSS 0.054617f
C21249 DVSS.n4858 VSS 0.082246f
C21250 DVSS.n4859 VSS 0.091242f
C21251 DVSS.n4860 VSS 0.091242f
C21252 DVSS.n4861 VSS 0.091242f
C21253 DVSS.n4862 VSS 0.091242f
C21254 DVSS.n4863 VSS 0.091242f
C21255 DVSS.n4864 VSS 0.091242f
C21256 DVSS.n4865 VSS 0.091242f
C21257 DVSS.n4866 VSS 0.091242f
C21258 DVSS.n4867 VSS 0.091242f
C21259 DVSS.n4868 VSS 0.091242f
C21260 DVSS.n4869 VSS 0.091242f
C21261 DVSS.n4870 VSS 0.091242f
C21262 DVSS.n4871 VSS 0.056223f
C21263 DVSS.n4872 VSS 0.045621f
C21264 DVSS.n4874 VSS 0.024233f
C21265 DVSS.n4875 VSS 0.045621f
C21266 DVSS.n4876 VSS 0.08064f
C21267 DVSS.n4877 VSS 0.091242f
C21268 DVSS.n4878 VSS 0.091242f
C21269 DVSS.n4879 VSS 0.091242f
C21270 DVSS.n4880 VSS 0.091242f
C21271 DVSS.n4881 VSS 0.091242f
C21272 DVSS.n4882 VSS 0.091242f
C21273 DVSS.n4883 VSS 0.063934f
C21274 DVSS.n4884 VSS 0.045803f
C21275 DVSS.n4885 VSS 0.051508f
C21276 DVSS.n4886 VSS 0.257333f
C21277 DVSS.n4887 VSS 0.026721f
C21278 DVSS.n4888 VSS 0.023334f
C21279 DVSS.n4889 VSS 0.045621f
C21280 DVSS.n4890 VSS 0.045621f
C21281 DVSS.n4891 VSS 0.091242f
C21282 DVSS.n4892 VSS 0.091242f
C21283 DVSS.n4893 VSS 0.091242f
C21284 DVSS.n4894 VSS 0.091242f
C21285 DVSS.n4895 VSS 0.091242f
C21286 DVSS.n4896 VSS 0.045621f
C21287 DVSS.n4897 VSS 0.045621f
C21288 DVSS.n4898 VSS 0.042127f
C21289 DVSS.n4899 VSS 0.051321f
C21290 DVSS.n4900 VSS 0.045803f
C21291 DVSS.n4901 VSS 0.072929f
C21292 DVSS.n4902 VSS 0.091242f
C21293 DVSS.n4903 VSS 0.091242f
C21294 DVSS.n4904 VSS 0.091242f
C21295 DVSS.n4905 VSS 0.091242f
C21296 DVSS.n4906 VSS 0.091242f
C21297 DVSS.n4907 VSS 0.091242f
C21298 DVSS.n4908 VSS 0.091242f
C21299 DVSS.n4909 VSS 0.091242f
C21300 DVSS.n4910 VSS 0.085781f
C21301 DVSS.n4911 VSS 0.091242f
C21302 DVSS.n4912 VSS 0.091242f
C21303 DVSS.n4913 VSS 0.091242f
C21304 DVSS.n4914 VSS 0.091242f
C21305 DVSS.n4915 VSS 0.091242f
C21306 DVSS.n4916 VSS 0.045621f
C21307 DVSS.n4917 VSS 0.045621f
C21308 DVSS.n4918 VSS 0.023334f
C21309 DVSS.n4919 VSS 0.026721f
C21310 DVSS.n4920 VSS 0.065489f
C21311 DVSS.n4921 VSS 0.044619f
C21312 DVSS.n4922 VSS 1.32141f
C21313 DVSS.n4923 VSS 2.04462f
C21314 DVSS.n4924 VSS 2.00358f
C21315 DVSS.n4925 VSS 2.80051f
C21316 DVSS.n4926 VSS 1.41279f
C21317 DVSS.n4927 VSS 2.34034f
C21318 DVSS.n4928 VSS 3.42636f
C21319 DVSS.n4929 VSS 2.13461f
C21320 DVSS.n4930 VSS 1.0789f
C21321 DVSS.n4931 VSS 0.024049f
C21322 DVSS.n4932 VSS 0.69228f
C21323 DVSS.n4933 VSS 0.676387f
C21324 DVSS.n4934 VSS 0.036625f
C21325 DVSS.n4935 VSS 0.338051f
C21326 DVSS.n4936 VSS 0.806716f
C21327 DVSS.n4937 VSS 0.376911f
C21328 DVSS.n4938 VSS 0.195519f
C21329 DVSS.n4939 VSS 0.195519f
C21330 DVSS.n4940 VSS 0.11084f
C21331 DVSS.n4941 VSS 0.135658f
C21332 DVSS.n4942 VSS 0.079024f
C21333 DVSS.n4943 VSS 0.07451f
C21334 DVSS.n4944 VSS 1.18906f
C21335 DVSS.n4945 VSS 0.495656f
C21336 DVSS.n4946 VSS 0.397285f
C21337 DVSS.n4947 VSS -0.005939f
C21338 DVSS.n4948 VSS 0.00423f
C21339 DVSS.n4949 VSS 0.00423f
C21340 DVSS.n4950 VSS 0.068858f
C21341 DVSS.n4951 VSS 0.019182f
C21342 DVSS.n4952 VSS 0.186341f
C21343 DVSS.n4953 VSS 0.248134f
C21344 DVSS.n4954 VSS 0.137875f
C21345 DVSS.n4955 VSS 0.209286f
C21346 DVSS.t194 VSS 0.169789f
C21347 DVSS.n4956 VSS 0.060777f
C21348 DVSS.n4957 VSS 0.002205f
C21349 DVSS.t82 VSS 0.00716f
C21350 DVSS.t195 VSS 0.00716f
C21351 DVSS.n4958 VSS 0.014896f
C21352 DVSS.n4959 VSS 0.006708f
C21353 DVSS.n4960 VSS 0.010442f
C21354 DVSS.n4961 VSS 0.019963f
C21355 DVSS.n4962 VSS 0.062886f
C21356 DVSS.n4963 VSS 0.349001f
C21357 DVSS.t136 VSS 0.169789f
C21358 DVSS.n4964 VSS 0.060777f
C21359 DVSS.n4965 VSS 0.002205f
C21360 DVSS.n4966 VSS 0.209286f
C21361 DVSS.n4967 VSS 0.137875f
C21362 DVSS.n4968 VSS 0.248134f
C21363 DVSS.n4969 VSS 0.231512f
C21364 DVSS.n4970 VSS 0.017012f
C21365 DVSS.n4971 VSS 0.00423f
C21366 DVSS.n4972 VSS 0.00423f
C21367 DVSS.n4973 VSS 0.068858f
C21368 DVSS.n4974 VSS 0.019182f
C21369 DVSS.n4975 VSS -0.005939f
C21370 DVSS.n4976 VSS 0.294016f
C21371 DVSS.n4977 VSS 0.439408f
C21372 DVSS.n4978 VSS 0.029922f
C21373 DVSS.n4979 VSS 0.07992f
C21374 DVSS.n4980 VSS 0.077106f
C21375 DVSS.n4981 VSS 0.091242f
C21376 DVSS.n4982 VSS 0.091242f
C21377 DVSS.n4983 VSS 0.091242f
C21378 DVSS.n4984 VSS 0.091242f
C21379 DVSS.n4985 VSS 0.091242f
C21380 DVSS.n4986 VSS 0.091242f
C21381 DVSS.n4987 VSS 0.091242f
C21382 DVSS.n4988 VSS 0.091242f
C21383 DVSS.n4989 VSS 0.091242f
C21384 DVSS.n4990 VSS 0.091242f
C21385 DVSS.n4991 VSS 0.091242f
C21386 DVSS.n4992 VSS 0.091242f
C21387 DVSS.n4993 VSS 0.091242f
C21388 DVSS.n4994 VSS 0.091242f
C21389 DVSS.n4995 VSS 0.091242f
C21390 DVSS.n4996 VSS 0.091242f
C21391 DVSS.n4997 VSS 0.091242f
C21392 DVSS.n4998 VSS 0.091242f
C21393 DVSS.n4999 VSS 0.091242f
C21394 DVSS.n5000 VSS 0.091242f
C21395 DVSS.n5001 VSS 0.091242f
C21396 DVSS.n5002 VSS 0.091242f
C21397 DVSS.n5003 VSS 0.091242f
C21398 DVSS.n5004 VSS 0.091242f
C21399 DVSS.n5005 VSS 0.091242f
C21400 DVSS.n5006 VSS 0.091242f
C21401 DVSS.n5007 VSS 0.091242f
C21402 DVSS.n5008 VSS 0.091242f
C21403 DVSS.n5009 VSS 0.091242f
C21404 DVSS.n5010 VSS 0.091242f
C21405 DVSS.n5011 VSS 0.091242f
C21406 DVSS.n5012 VSS 0.091242f
C21407 DVSS.n5013 VSS 0.091242f
C21408 DVSS.n5014 VSS 0.091242f
C21409 DVSS.n5015 VSS 0.091242f
C21410 DVSS.n5016 VSS 0.091242f
C21411 DVSS.n5017 VSS 0.091242f
C21412 DVSS.n5018 VSS 0.091242f
C21413 DVSS.n5019 VSS 0.091242f
C21414 DVSS.n5020 VSS 0.091242f
C21415 DVSS.n5021 VSS 0.091242f
C21416 DVSS.n5022 VSS 0.091242f
C21417 DVSS.n5023 VSS 0.091242f
C21418 DVSS.n5024 VSS 0.091242f
C21419 DVSS.n5025 VSS 0.091242f
C21420 DVSS.n5026 VSS 0.091242f
C21421 DVSS.n5027 VSS 0.091242f
C21422 DVSS.n5028 VSS 0.091242f
C21423 DVSS.n5029 VSS 0.091242f
C21424 DVSS.n5030 VSS 0.091242f
C21425 DVSS.n5031 VSS 0.091242f
C21426 DVSS.n5032 VSS 0.091242f
C21427 DVSS.n5033 VSS 0.091242f
C21428 DVSS.n5034 VSS 0.091242f
C21429 DVSS.n5035 VSS 0.091242f
C21430 DVSS.n5036 VSS 0.091242f
C21431 DVSS.n5037 VSS 0.091242f
C21432 DVSS.n5038 VSS 0.091242f
C21433 DVSS.n5039 VSS 0.091242f
C21434 DVSS.n5040 VSS 0.091242f
C21435 DVSS.n5041 VSS 0.091242f
C21436 DVSS.n5042 VSS 0.091242f
C21437 DVSS.n5043 VSS 0.045621f
C21438 DVSS.n5044 VSS 0.045621f
C21439 DVSS.n5045 VSS 0.011779f
C21440 DVSS.n5046 VSS 0.004953f
C21441 DVSS.n5047 VSS 0.045621f
C21442 DVSS.n5048 VSS 0.045621f
C21443 DVSS.n5049 VSS 0.091242f
C21444 DVSS.n5050 VSS 0.091242f
C21445 DVSS.n5051 VSS 0.091242f
C21446 DVSS.n5052 VSS 0.091242f
C21447 DVSS.n5053 VSS 0.091242f
C21448 DVSS.n5054 VSS 0.045621f
C21449 DVSS.n5055 VSS 0.045621f
C21450 DVSS.n5056 VSS 0.004953f
C21451 DVSS.n5057 VSS 0.010501f
C21452 DVSS.n5058 VSS 0.045621f
C21453 DVSS.n5059 VSS 0.045621f
C21454 DVSS.n5060 VSS 0.091242f
C21455 DVSS.n5061 VSS 0.091242f
C21456 DVSS.n5062 VSS 0.091242f
C21457 DVSS.n5063 VSS 0.091242f
C21458 DVSS.n5064 VSS 0.091242f
C21459 DVSS.n5065 VSS 0.091242f
C21460 DVSS.n5066 VSS 0.091242f
C21461 DVSS.n5067 VSS 0.091242f
C21462 DVSS.n5068 VSS 0.091242f
C21463 DVSS.n5069 VSS 0.091242f
C21464 DVSS.n5070 VSS 0.091242f
C21465 DVSS.n5071 VSS 0.091242f
C21466 DVSS.n5072 VSS 0.091242f
C21467 DVSS.n5073 VSS 0.091242f
C21468 DVSS.n5074 VSS 0.049155f
C21469 DVSS.n5075 VSS 0.057771f
C21470 DVSS.n5076 VSS 0.045621f
C21471 DVSS.n5077 VSS 0.091242f
C21472 DVSS.n5078 VSS 0.091242f
C21473 DVSS.n5079 VSS 0.091242f
C21474 DVSS.n5080 VSS 0.091242f
C21475 DVSS.n5081 VSS 0.091242f
C21476 DVSS.n5082 VSS 0.091242f
C21477 DVSS.n5083 VSS 0.091242f
C21478 DVSS.n5084 VSS 0.091242f
C21479 DVSS.n5085 VSS 0.091242f
C21480 DVSS.n5086 VSS 0.091242f
C21481 DVSS.n5087 VSS 0.091242f
C21482 DVSS.n5088 VSS 0.091242f
C21483 DVSS.n5089 VSS 0.091242f
C21484 DVSS.n5090 VSS 0.091242f
C21485 DVSS.n5091 VSS 0.091242f
C21486 DVSS.n5092 VSS 0.091242f
C21487 DVSS.n5093 VSS 0.091242f
C21488 DVSS.n5094 VSS 0.091242f
C21489 DVSS.n5095 VSS 0.091242f
C21490 DVSS.n5096 VSS 0.091242f
C21491 DVSS.n5097 VSS 0.091242f
C21492 DVSS.n5098 VSS 0.091242f
C21493 DVSS.n5099 VSS 0.091242f
C21494 DVSS.n5100 VSS 0.091242f
C21495 DVSS.n5101 VSS 0.091242f
C21496 DVSS.n5102 VSS 0.091242f
C21497 DVSS.n5103 VSS 0.091242f
C21498 DVSS.n5104 VSS 0.338098f
C21499 DVSS.n5105 VSS 0.091242f
C21500 DVSS.n5106 VSS 0.091242f
C21501 DVSS.n5107 VSS 0.091242f
C21502 DVSS.n5108 VSS 0.194467f
C21503 DVSS.n5109 VSS 0.667361f
C21504 DVSS.n5110 VSS 0.81998f
C21505 DVSS.n5111 VSS 1.34585f
C21506 DVSS.n5112 VSS 1.8704f
C21507 DVSS.n5113 VSS 1.91961f
C21508 DVSS.n5114 VSS 1.80894f
C21509 DVSS.n5115 VSS 0.471354f
C21510 DVSS.n5116 VSS 0.030675f
C21511 DVSS.n5117 VSS 0.030675f
C21512 DVSS.n5118 VSS 0.012179f
C21513 DVSS.n5119 VSS 0.784185f
C21514 DVSS.n5120 VSS 0.784185f
C21515 DVSS.n5121 VSS 0.784185f
C21516 DVSS.n5122 VSS 0.012179f
C21517 DVSS.n5123 VSS 0.030675f
C21518 DVSS.n5124 VSS 0.030675f
C21519 DVSS.n5125 VSS 0.030675f
C21520 DVSS.n5126 VSS 0.012179f
C21521 DVSS.n5127 VSS 0.784185f
C21522 DVSS.n5128 VSS 0.784185f
C21523 DVSS.n5129 VSS 0.784185f
C21524 DVSS.n5130 VSS 0.012179f
C21525 DVSS.n5131 VSS 0.030675f
C21526 DVSS.n5132 VSS 0.030675f
C21527 DVSS.n5133 VSS 0.030675f
C21528 DVSS.n5134 VSS 0.012179f
C21529 DVSS.n5135 VSS 0.784185f
C21530 DVSS.n5136 VSS 0.784185f
C21531 DVSS.n5137 VSS 0.784185f
C21532 DVSS.n5138 VSS 0.012179f
C21533 DVSS.n5139 VSS 0.030675f
C21534 DVSS.n5140 VSS 0.030675f
C21535 DVSS.n5141 VSS 0.030675f
C21536 DVSS.n5142 VSS 0.012179f
C21537 DVSS.n5143 VSS 0.784185f
C21538 DVSS.n5144 VSS 0.784185f
C21539 DVSS.n5145 VSS 0.784185f
C21540 DVSS.n5146 VSS 0.012179f
C21541 DVSS.n5147 VSS 0.030675f
C21542 DVSS.n5148 VSS 0.030675f
C21543 DVSS.n5149 VSS 0.030675f
C21544 DVSS.n5150 VSS 0.012179f
C21545 DVSS.n5151 VSS 0.784185f
C21546 DVSS.n5152 VSS 0.784185f
C21547 DVSS.n5153 VSS 0.784185f
C21548 DVSS.n5154 VSS 0.012179f
C21549 DVSS.n5155 VSS 0.030675f
C21550 DVSS.n5156 VSS 0.030675f
C21551 DVSS.n5157 VSS 0.030675f
C21552 DVSS.n5158 VSS 0.012179f
C21553 DVSS.n5159 VSS 0.784185f
C21554 DVSS.n5160 VSS 0.784185f
C21555 DVSS.n5161 VSS 0.784185f
C21556 DVSS.n5162 VSS 0.012179f
C21557 DVSS.n5163 VSS 0.030675f
C21558 DVSS.n5164 VSS 0.030675f
C21559 DVSS.n5165 VSS 0.030675f
C21560 DVSS.n5166 VSS 0.012179f
C21561 DVSS.n5167 VSS 0.784185f
C21562 DVSS.n5168 VSS 0.784185f
C21563 DVSS.n5169 VSS 0.784185f
C21564 DVSS.n5170 VSS 0.012179f
C21565 DVSS.n5171 VSS 0.030675f
C21566 DVSS.n5172 VSS 0.030675f
C21567 DVSS.n5173 VSS 0.030675f
C21568 DVSS.n5174 VSS 0.012179f
C21569 DVSS.n5175 VSS 0.784185f
C21570 DVSS.n5176 VSS 0.784185f
C21571 DVSS.n5177 VSS 0.784185f
C21572 DVSS.n5178 VSS 0.012179f
C21573 DVSS.n5179 VSS 0.030675f
C21574 DVSS.n5180 VSS 0.030675f
C21575 DVSS.n5181 VSS 0.030675f
C21576 DVSS.n5182 VSS 0.012179f
C21577 DVSS.n5183 VSS 0.784185f
C21578 DVSS.n5184 VSS 0.784185f
C21579 DVSS.n5185 VSS 0.784185f
C21580 DVSS.n5186 VSS 0.012179f
C21581 DVSS.n5187 VSS 0.030675f
C21582 DVSS.n5188 VSS 0.030675f
C21583 DVSS.n5189 VSS 0.030675f
C21584 DVSS.n5190 VSS 0.012179f
C21585 DVSS.n5191 VSS 0.784185f
C21586 DVSS.n5192 VSS 0.784185f
C21587 DVSS.n5193 VSS 0.784185f
C21588 DVSS.n5194 VSS 0.012179f
C21589 DVSS.n5195 VSS 0.030675f
C21590 DVSS.n5196 VSS 0.030675f
C21591 DVSS.n5197 VSS 0.030675f
C21592 DVSS.n5198 VSS 0.012179f
C21593 DVSS.n5199 VSS 0.784185f
C21594 DVSS.n5200 VSS 0.784185f
C21595 DVSS.n5201 VSS 0.784185f
C21596 DVSS.n5202 VSS 0.012179f
C21597 DVSS.n5203 VSS 0.030675f
C21598 DVSS.n5204 VSS 0.030675f
C21599 DVSS.n5205 VSS 0.030675f
C21600 DVSS.n5206 VSS 0.012179f
C21601 DVSS.n5207 VSS 0.784185f
C21602 DVSS.n5208 VSS 0.784185f
C21603 DVSS.n5209 VSS 0.784185f
C21604 DVSS.n5210 VSS 0.012179f
C21605 DVSS.n5211 VSS 0.030675f
C21606 DVSS.n5212 VSS 0.030675f
C21607 DVSS.n5213 VSS 0.030675f
C21608 DVSS.n5214 VSS 0.012179f
C21609 DVSS.n5215 VSS 0.784185f
C21610 DVSS.n5216 VSS 0.784185f
C21611 DVSS.n5217 VSS 0.784185f
C21612 DVSS.n5218 VSS 0.012179f
C21613 DVSS.n5219 VSS 0.030675f
C21614 DVSS.n5220 VSS 0.030675f
C21615 DVSS.n5221 VSS 0.030675f
C21616 DVSS.n5222 VSS 0.030675f
C21617 DVSS.n5223 VSS 0.012179f
C21618 DVSS.n5224 VSS 0.784185f
C21619 DVSS.n5225 VSS 0.784185f
C21620 DVSS.n5226 VSS 0.784185f
C21621 DVSS.n5227 VSS 0.012179f
C21622 DVSS.n5228 VSS 0.012179f
C21623 DVSS.n5229 VSS 0.022883f
C21624 DVSS.n5230 VSS 0.015337f
C21625 DVSS.n5231 VSS 2.30011f
C21626 DVSS.n5232 VSS 0.392092f
C21627 DVSS.n5233 VSS 0.5913f
C21628 DVSS.n5234 VSS 0.784185f
C21629 DVSS.n5235 VSS 0.012179f
C21630 DVSS.n5236 VSS 0.030675f
C21631 DVSS.n5237 VSS 0.030675f
C21632 DVSS.n5238 VSS 0.030675f
C21633 DVSS.n5239 VSS 0.012179f
C21634 DVSS.n5240 VSS 0.784185f
C21635 DVSS.n5241 VSS 0.784185f
C21636 DVSS.n5242 VSS 0.784185f
C21637 DVSS.n5243 VSS 0.012179f
C21638 DVSS.n5244 VSS 0.030675f
C21639 DVSS.n5245 VSS 0.030675f
C21640 DVSS.n5246 VSS 0.030675f
C21641 DVSS.n5247 VSS 0.012179f
C21642 DVSS.n5248 VSS 0.784185f
C21643 DVSS.n5249 VSS 0.784185f
C21644 DVSS.n5250 VSS 0.784185f
C21645 DVSS.n5251 VSS 0.012179f
C21646 DVSS.n5252 VSS 0.030675f
C21647 DVSS.n5253 VSS 0.030675f
C21648 DVSS.n5254 VSS 0.030675f
C21649 DVSS.n5255 VSS 0.012179f
C21650 DVSS.n5256 VSS 0.784185f
C21651 DVSS.n5257 VSS 0.784185f
C21652 DVSS.n5258 VSS 0.784185f
C21653 DVSS.n5259 VSS 0.012179f
C21654 DVSS.n5260 VSS 0.030675f
C21655 DVSS.n5261 VSS 0.030675f
C21656 DVSS.n5262 VSS 0.030675f
C21657 DVSS.n5263 VSS 0.012179f
C21658 DVSS.n5264 VSS 0.784185f
C21659 DVSS.n5265 VSS 0.784185f
C21660 DVSS.n5266 VSS 0.784185f
C21661 DVSS.n5267 VSS 0.012179f
C21662 DVSS.n5268 VSS 0.030675f
C21663 DVSS.n5269 VSS 0.030675f
C21664 DVSS.n5270 VSS 0.030675f
C21665 DVSS.n5271 VSS 0.012179f
C21666 DVSS.n5272 VSS 0.784185f
C21667 DVSS.n5273 VSS 0.784185f
C21668 DVSS.n5274 VSS 0.784185f
C21669 DVSS.n5275 VSS 0.012179f
C21670 DVSS.n5276 VSS 0.030675f
C21671 DVSS.n5277 VSS 0.030675f
C21672 DVSS.n5278 VSS 0.030675f
C21673 DVSS.n5279 VSS 0.012179f
C21674 DVSS.n5280 VSS 0.784185f
C21675 DVSS.n5281 VSS 0.784185f
C21676 DVSS.n5282 VSS 0.784185f
C21677 DVSS.n5283 VSS 0.012179f
C21678 DVSS.n5284 VSS 0.030675f
C21679 DVSS.n5285 VSS 0.030675f
C21680 DVSS.n5286 VSS 0.030675f
C21681 DVSS.n5287 VSS 0.012179f
C21682 DVSS.n5288 VSS 0.784185f
C21683 DVSS.n5289 VSS 0.784185f
C21684 DVSS.n5290 VSS 0.784185f
C21685 DVSS.n5291 VSS 0.012179f
C21686 DVSS.n5292 VSS 0.030675f
C21687 DVSS.n5293 VSS 0.030675f
C21688 DVSS.n5294 VSS 0.030675f
C21689 DVSS.n5295 VSS 0.012179f
C21690 DVSS.n5296 VSS 0.784185f
C21691 DVSS.n5297 VSS 0.784185f
C21692 DVSS.n5298 VSS 0.784185f
C21693 DVSS.n5299 VSS 0.012179f
C21694 DVSS.n5300 VSS 0.030675f
C21695 DVSS.n5301 VSS 0.030675f
C21696 DVSS.n5302 VSS 0.030675f
C21697 DVSS.n5303 VSS 0.012179f
C21698 DVSS.n5304 VSS 0.784185f
C21699 DVSS.n5305 VSS 0.784185f
C21700 DVSS.n5306 VSS 0.784185f
C21701 DVSS.n5307 VSS 0.012179f
C21702 DVSS.n5308 VSS 0.030675f
C21703 DVSS.n5309 VSS 0.030675f
C21704 DVSS.n5310 VSS 0.030675f
C21705 DVSS.n5311 VSS 0.012179f
C21706 DVSS.n5312 VSS 0.784185f
C21707 DVSS.n5313 VSS 0.784185f
C21708 DVSS.n5314 VSS 0.784185f
C21709 DVSS.n5315 VSS 0.012179f
C21710 DVSS.n5316 VSS 0.030675f
C21711 DVSS.n5317 VSS 0.030675f
C21712 DVSS.n5318 VSS 0.030675f
C21713 DVSS.n5319 VSS 0.012179f
C21714 DVSS.n5320 VSS 0.784185f
C21715 DVSS.n5321 VSS 0.784185f
C21716 DVSS.n5322 VSS 0.784185f
C21717 DVSS.n5323 VSS 0.012179f
C21718 DVSS.n5324 VSS 0.030675f
C21719 DVSS.n5325 VSS 0.030675f
C21720 DVSS.n5326 VSS 0.030675f
C21721 DVSS.n5327 VSS 0.012179f
C21722 DVSS.n5328 VSS 0.784185f
C21723 DVSS.n5329 VSS 0.784185f
C21724 DVSS.n5330 VSS 0.784185f
C21725 DVSS.n5331 VSS 0.012179f
C21726 DVSS.n5332 VSS 0.030675f
C21727 DVSS.n5333 VSS 0.030675f
C21728 DVSS.n5334 VSS 0.030675f
C21729 DVSS.n5335 VSS 0.012179f
C21730 DVSS.n5336 VSS 0.784185f
C21731 DVSS.n5337 VSS 0.784185f
C21732 DVSS.n5338 VSS 0.784185f
C21733 DVSS.n5339 VSS 0.012179f
C21734 DVSS.n5340 VSS 0.030675f
C21735 DVSS.n5341 VSS 0.030675f
C21736 DVSS.n5342 VSS 0.030675f
C21737 DVSS.n5343 VSS 0.030675f
C21738 DVSS.n5344 VSS 0.012179f
C21739 DVSS.n5345 VSS 0.784185f
C21740 DVSS.n5346 VSS 0.784185f
C21741 DVSS.n5347 VSS 0.553356f
C21742 DVSS.n5348 VSS 0.012179f
C21743 DVSS.n5349 VSS 1.91432f
C21744 DVSS.n5350 VSS 0.390646f
C21745 DVSS.n5351 VSS 1.12456f
C21746 DVSS.n5352 VSS 1.77831f
C21747 DVSS.n5353 VSS 5.96489f
C21748 DVSS.n5354 VSS 2.37815f
C21749 DVSS.n5355 VSS 2.37781f
C21750 DVSS.n5356 VSS 4.34557f
C21751 DVSS.n5357 VSS 2.04923f
C21752 DVSS.n5358 VSS 3.32639f
C21753 DVSS.n5359 VSS 0.045445f
C21754 DVSS.n5360 VSS 0.046912f
C21755 DVSS.n5361 VSS 0.04889f
C21756 DVSS.n5362 VSS 0.078712f
C21757 DVSS.n5363 VSS 0.091242f
C21758 DVSS.n5364 VSS 0.091242f
C21759 DVSS.n5365 VSS 0.091242f
C21760 DVSS.n5366 VSS 0.091242f
C21761 DVSS.n5367 VSS 0.091242f
C21762 DVSS.n5368 VSS 0.091242f
C21763 DVSS.n5369 VSS 0.091242f
C21764 DVSS.n5370 VSS 0.091242f
C21765 DVSS.n5371 VSS 0.091242f
C21766 DVSS.n5372 VSS 0.091242f
C21767 DVSS.n5373 VSS 0.091242f
C21768 DVSS.n5374 VSS 0.091242f
C21769 DVSS.n5375 VSS 0.091242f
C21770 DVSS.n5376 VSS 0.091242f
C21771 DVSS.n5377 VSS 0.091242f
C21772 DVSS.n5378 VSS 0.091242f
C21773 DVSS.n5379 VSS 0.091242f
C21774 DVSS.n5380 VSS 0.091242f
C21775 DVSS.n5381 VSS 0.091242f
C21776 DVSS.n5382 VSS 0.091242f
C21777 DVSS.n5383 VSS 0.091242f
C21778 DVSS.n5384 VSS 0.091242f
C21779 DVSS.n5385 VSS 0.091242f
C21780 DVSS.n5386 VSS 0.091242f
C21781 DVSS.n5387 VSS 0.091242f
C21782 DVSS.n5388 VSS 0.091242f
C21783 DVSS.n5389 VSS 0.091242f
C21784 DVSS.n5390 VSS 0.091242f
C21785 DVSS.n5391 VSS 0.091242f
C21786 DVSS.n5392 VSS 0.091242f
C21787 DVSS.n5393 VSS 0.091242f
C21788 DVSS.n5394 VSS 0.091242f
C21789 DVSS.n5395 VSS 0.091242f
C21790 DVSS.n5396 VSS 0.091242f
C21791 DVSS.n5397 VSS 0.091242f
C21792 DVSS.n5398 VSS 0.091242f
C21793 DVSS.n5399 VSS 0.091242f
C21794 DVSS.n5400 VSS 0.091242f
C21795 DVSS.n5401 VSS 0.091242f
C21796 DVSS.n5402 VSS 0.091242f
C21797 DVSS.n5403 VSS 0.091242f
C21798 DVSS.n5404 VSS 0.091242f
C21799 DVSS.n5405 VSS 0.091242f
C21800 DVSS.n5406 VSS 0.091242f
C21801 DVSS.n5407 VSS 0.091242f
C21802 DVSS.n5408 VSS 0.091242f
C21803 DVSS.n5409 VSS 0.091242f
C21804 DVSS.n5410 VSS 0.091242f
C21805 DVSS.n5411 VSS 0.091242f
C21806 DVSS.n5412 VSS 0.091242f
C21807 DVSS.n5413 VSS 0.091242f
C21808 DVSS.n5414 VSS 0.091242f
C21809 DVSS.n5415 VSS 0.091242f
C21810 DVSS.n5416 VSS 0.091242f
C21811 DVSS.n5417 VSS 0.091242f
C21812 DVSS.n5418 VSS 0.091242f
C21813 DVSS.n5419 VSS 0.091242f
C21814 DVSS.n5420 VSS 0.091242f
C21815 DVSS.n5421 VSS 0.091242f
C21816 DVSS.n5422 VSS 0.091242f
C21817 DVSS.n5423 VSS 0.091242f
C21818 DVSS.n5424 VSS 0.091242f
C21819 DVSS.n5425 VSS 0.091242f
C21820 DVSS.n5426 VSS 0.091242f
C21821 DVSS.n5427 VSS 0.091242f
C21822 DVSS.n5428 VSS 0.091242f
C21823 DVSS.n5429 VSS 0.091242f
C21824 DVSS.n5430 VSS 0.091242f
C21825 DVSS.n5431 VSS 0.091242f
C21826 DVSS.n5432 VSS 0.091242f
C21827 DVSS.n5433 VSS 0.091242f
C21828 DVSS.n5434 VSS 0.091242f
C21829 DVSS.n5435 VSS 0.091242f
C21830 DVSS.n5436 VSS 0.091242f
C21831 DVSS.n5437 VSS 0.091242f
C21832 DVSS.n5438 VSS 0.091242f
C21833 DVSS.n5439 VSS 0.091242f
C21834 DVSS.n5440 VSS 0.091242f
C21835 DVSS.n5441 VSS 0.091242f
C21836 DVSS.n5442 VSS 0.091242f
C21837 DVSS.n5443 VSS 0.091242f
C21838 DVSS.n5444 VSS 0.091242f
C21839 DVSS.n5445 VSS 0.091242f
C21840 DVSS.n5446 VSS 0.091242f
C21841 DVSS.n5447 VSS 0.091242f
C21842 DVSS.n5448 VSS 0.091242f
C21843 DVSS.n5449 VSS 0.091242f
C21844 DVSS.n5450 VSS 0.091242f
C21845 DVSS.n5451 VSS 0.091242f
C21846 DVSS.n5452 VSS 0.091242f
C21847 DVSS.n5453 VSS 0.091242f
C21848 DVSS.n5454 VSS 0.091242f
C21849 DVSS.n5455 VSS 0.091242f
C21850 DVSS.n5456 VSS 0.091242f
C21851 DVSS.n5457 VSS 0.091242f
C21852 DVSS.n5458 VSS 0.091242f
C21853 DVSS.n5459 VSS 0.091242f
C21854 DVSS.n5460 VSS 0.091242f
C21855 DVSS.n5461 VSS 0.091242f
C21856 DVSS.n5462 VSS 0.091242f
C21857 DVSS.n5463 VSS 0.091242f
C21858 DVSS.n5464 VSS 0.091242f
C21859 DVSS.n5465 VSS 0.091242f
C21860 DVSS.n5466 VSS 0.091242f
C21861 DVSS.n5467 VSS 0.091242f
C21862 DVSS.n5468 VSS 0.091242f
C21863 DVSS.n5469 VSS 0.091242f
C21864 DVSS.n5470 VSS 0.091242f
C21865 DVSS.n5471 VSS 0.091242f
C21866 DVSS.n5472 VSS 0.091242f
C21867 DVSS.n5473 VSS 0.091242f
C21868 DVSS.n5474 VSS 0.091242f
C21869 DVSS.n5475 VSS 0.091242f
C21870 DVSS.n5476 VSS 0.091242f
C21871 DVSS.n5477 VSS 0.091242f
C21872 DVSS.n5478 VSS 0.091242f
C21873 DVSS.n5479 VSS 0.091242f
C21874 DVSS.n5480 VSS 0.091242f
C21875 DVSS.n5481 VSS 0.091242f
C21876 DVSS.n5482 VSS 0.091242f
C21877 DVSS.n5483 VSS 0.091242f
C21878 DVSS.n5484 VSS 0.091242f
C21879 DVSS.n5485 VSS 0.091242f
C21880 DVSS.n5486 VSS 0.091242f
C21881 DVSS.n5487 VSS 0.091242f
C21882 DVSS.n5488 VSS 0.091242f
C21883 DVSS.n5489 VSS 0.091242f
C21884 DVSS.n5490 VSS 0.091242f
C21885 DVSS.n5491 VSS 0.091242f
C21886 DVSS.n5492 VSS 0.091242f
C21887 DVSS.n5493 VSS 0.091242f
C21888 DVSS.n5494 VSS 0.091242f
C21889 DVSS.n5495 VSS 0.091242f
C21890 DVSS.n5496 VSS 0.091242f
C21891 DVSS.n5497 VSS 0.091242f
C21892 DVSS.n5498 VSS 0.091242f
C21893 DVSS.n5499 VSS 0.091242f
C21894 DVSS.n5500 VSS 0.091242f
C21895 DVSS.n5501 VSS 0.091242f
C21896 DVSS.n5502 VSS 0.091242f
C21897 DVSS.n5503 VSS 0.091242f
C21898 DVSS.n5504 VSS 0.091242f
C21899 DVSS.n5505 VSS 0.091242f
C21900 DVSS.n5506 VSS 0.091242f
C21901 DVSS.n5507 VSS 0.091242f
C21902 DVSS.n5508 VSS 0.091242f
C21903 DVSS.n5509 VSS 0.091242f
C21904 DVSS.n5510 VSS 0.091242f
C21905 DVSS.n5511 VSS 0.091242f
C21906 DVSS.n5512 VSS 0.091242f
C21907 DVSS.n5513 VSS 0.091242f
C21908 DVSS.n5514 VSS 0.091242f
C21909 DVSS.n5515 VSS 0.091242f
C21910 DVSS.n5516 VSS 0.091242f
C21911 DVSS.n5517 VSS 0.091242f
C21912 DVSS.n5518 VSS 0.091242f
C21913 DVSS.n5519 VSS 0.091242f
C21914 DVSS.n5520 VSS 0.091242f
C21915 DVSS.n5521 VSS 0.091242f
C21916 DVSS.n5522 VSS 0.091242f
C21917 DVSS.n5523 VSS 0.091242f
C21918 DVSS.n5524 VSS 0.091242f
C21919 DVSS.n5525 VSS 0.091242f
C21920 DVSS.n5526 VSS 0.091242f
C21921 DVSS.n5527 VSS 0.091242f
C21922 DVSS.n5528 VSS 0.091242f
C21923 DVSS.n5529 VSS 0.091242f
C21924 DVSS.n5530 VSS 0.091242f
C21925 DVSS.n5531 VSS 0.091242f
C21926 DVSS.n5532 VSS 0.091242f
C21927 DVSS.n5533 VSS 0.091242f
C21928 DVSS.n5534 VSS 0.091242f
C21929 DVSS.n5535 VSS 0.091242f
C21930 DVSS.n5536 VSS 0.091242f
C21931 DVSS.n5537 VSS 0.091242f
C21932 DVSS.n5538 VSS 0.091242f
C21933 DVSS.n5539 VSS 0.091242f
C21934 DVSS.n5540 VSS 0.091242f
C21935 DVSS.n5541 VSS 0.091242f
C21936 DVSS.n5542 VSS 0.091242f
C21937 DVSS.n5543 VSS 0.091242f
C21938 DVSS.n5544 VSS 0.091242f
C21939 DVSS.n5545 VSS 0.091242f
C21940 DVSS.n5546 VSS 0.091242f
C21941 DVSS.n5547 VSS 0.082246f
C21942 DVSS.n5548 VSS 0.082246f
C21943 DVSS.n5549 VSS 0.091242f
C21944 DVSS.n5550 VSS 0.046906f
C21945 DVSS.n5551 VSS 0.12011f
C21946 DVSS.n5552 VSS 0.045621f
C21947 DVSS.n5553 VSS 0.008996f
C21948 DVSS.n5554 VSS 0.134627f
C21949 DVSS.n5555 VSS 0.106547f
C21950 DVSS.n5556 VSS 0.007104f
C21951 DVSS.n5557 VSS 0.025114f
C21952 DVSS.n5558 VSS 0.007104f
C21953 DVSS.n5559 VSS 0.025114f
C21954 DVSS.n5560 VSS 0.247841f
C21955 DVSS.n5561 VSS 0.12174f
C21956 DVSS.n5562 VSS 0.352343f
C21957 DVSS.n5563 VSS 0.730699f
C21958 DVSS.n5564 VSS 0.192765f
C21959 DVSS.n5565 VSS 0.195519f
C21960 DVSS.n5566 VSS 0.117036f
C21961 DVSS.n5567 VSS 0.176242f
C21962 DVSS.n5568 VSS 0.195519f
C21963 DVSS.n5569 VSS 0.195519f
C21964 DVSS.n5570 VSS 0.195519f
C21965 DVSS.n5571 VSS 0.195519f
C21966 DVSS.n5572 VSS 0.195519f
C21967 DVSS.n5573 VSS 0.195519f
C21968 DVSS.n5574 VSS 0.195519f
C21969 DVSS.n5575 VSS 0.195519f
C21970 DVSS.n5576 VSS 0.195519f
C21971 DVSS.n5577 VSS 0.195519f
C21972 DVSS.n5578 VSS 0.195519f
C21973 DVSS.n5579 VSS 0.195519f
C21974 DVSS.n5580 VSS 0.195519f
C21975 DVSS.n5581 VSS 0.195519f
C21976 DVSS.n5582 VSS 0.178996f
C21977 DVSS.n5583 VSS 0.178996f
C21978 DVSS.n5584 VSS 0.235449f
C21979 DVSS.n5585 VSS 0.114282f
C21980 DVSS.n5586 VSS 0.114282f
C21981 DVSS.n5587 VSS 0.195519f
C21982 DVSS.n5588 VSS 0.195519f
C21983 DVSS.n5589 VSS 0.195519f
C21984 DVSS.n5590 VSS 0.195519f
C21985 DVSS.n5591 VSS 0.195519f
C21986 DVSS.n5592 VSS 0.195519f
C21987 DVSS.n5593 VSS 0.195519f
C21988 DVSS.n5594 VSS 0.195519f
C21989 DVSS.n5595 VSS 0.195519f
C21990 DVSS.n5596 VSS 0.195519f
C21991 DVSS.n5597 VSS 0.195519f
C21992 DVSS.n5598 VSS 0.195519f
C21993 DVSS.n5599 VSS 0.195519f
C21994 DVSS.n5600 VSS 0.195519f
C21995 DVSS.n5601 VSS 0.195519f
C21996 DVSS.n5602 VSS 0.195519f
C21997 DVSS.n5603 VSS 0.195519f
C21998 DVSS.n5604 VSS 0.195519f
C21999 DVSS.n5605 VSS 0.195519f
C22000 DVSS.n5606 VSS 0.195519f
C22001 DVSS.n5607 VSS 0.195519f
C22002 DVSS.n5608 VSS 0.195519f
C22003 DVSS.n5609 VSS 0.195519f
C22004 DVSS.n5610 VSS 0.195519f
C22005 DVSS.n5611 VSS 0.195519f
C22006 DVSS.n5612 VSS 0.195519f
C22007 DVSS.n5613 VSS 0.195519f
C22008 DVSS.n5614 VSS 0.176931f
C22009 DVSS.n5615 VSS 0.480814f
C22010 DVSS.n5616 VSS 0.483842f
C22011 DVSS.n5617 VSS 0.143051f
C22012 DVSS.n5618 VSS 0.176931f
C22013 DVSS.n5619 VSS 0.195519f
C22014 DVSS.n5620 VSS 0.195519f
C22015 DVSS.n5621 VSS 0.195519f
C22016 DVSS.n5622 VSS 0.195519f
C22017 DVSS.n5623 VSS 0.195519f
C22018 DVSS.n5624 VSS 0.195519f
C22019 DVSS.n5625 VSS 0.195519f
C22020 DVSS.n5626 VSS 0.195519f
C22021 DVSS.n5627 VSS 0.195519f
C22022 DVSS.n5628 VSS 0.195519f
C22023 DVSS.n5629 VSS 0.195519f
C22024 DVSS.n5630 VSS 0.195519f
C22025 DVSS.n5631 VSS 0.195519f
C22026 DVSS.n5632 VSS 0.195519f
C22027 DVSS.n5633 VSS 0.195519f
C22028 DVSS.n5634 VSS 0.195519f
C22029 DVSS.n5635 VSS 0.195519f
C22030 DVSS.n5636 VSS 0.195519f
C22031 DVSS.n5637 VSS 0.195519f
C22032 DVSS.n5638 VSS 0.195519f
C22033 DVSS.n5639 VSS 0.195519f
C22034 DVSS.n5640 VSS 0.195519f
C22035 DVSS.n5641 VSS 0.195519f
C22036 DVSS.n5642 VSS 0.195519f
C22037 DVSS.n5643 VSS 0.195519f
C22038 DVSS.n5644 VSS 0.195519f
C22039 DVSS.n5645 VSS 0.195519f
C22040 DVSS.n5646 VSS 0.195519f
C22041 DVSS.n5647 VSS 0.195519f
C22042 DVSS.n5648 VSS 0.195519f
C22043 DVSS.n5649 VSS 0.195519f
C22044 DVSS.n5650 VSS 0.195519f
C22045 DVSS.n5651 VSS 0.195519f
C22046 DVSS.n5652 VSS 0.195519f
C22047 DVSS.n5653 VSS 0.195519f
C22048 DVSS.n5654 VSS 0.195519f
C22049 DVSS.n5655 VSS 0.195519f
C22050 DVSS.n5656 VSS 0.195519f
C22051 DVSS.n5657 VSS 0.195519f
C22052 DVSS.n5658 VSS 0.195519f
C22053 DVSS.n5659 VSS 0.195519f
C22054 DVSS.n5660 VSS 0.195519f
C22055 DVSS.n5661 VSS 0.195519f
C22056 DVSS.n5662 VSS 0.195519f
C22057 DVSS.n5663 VSS 0.195519f
C22058 DVSS.n5664 VSS 0.173489f
C22059 DVSS.n5665 VSS 0.173489f
C22060 DVSS.n5666 VSS 0.373138f
C22061 DVSS.n5667 VSS 0.235449f
C22062 DVSS.n5668 VSS 0.11979f
C22063 DVSS.n5669 VSS 0.11979f
C22064 DVSS.n5670 VSS 0.235449f
C22065 DVSS.n5671 VSS 0.173489f
C22066 DVSS.n5672 VSS 0.195519f
C22067 DVSS.n5673 VSS 0.195519f
C22068 DVSS.n5674 VSS 0.195519f
C22069 DVSS.n5675 VSS 0.195519f
C22070 DVSS.n5676 VSS 0.116347f
C22071 DVSS.n5677 VSS 0.195519f
C22072 DVSS.n5678 VSS 0.195519f
C22073 DVSS.n5679 VSS 0.195519f
C22074 DVSS.n5680 VSS 0.195519f
C22075 DVSS.n5681 VSS 0.195519f
C22076 DVSS.n5682 VSS 0.195519f
C22077 DVSS.n5683 VSS 0.176931f
C22078 DVSS.n5684 VSS 0.195519f
C22079 DVSS.n5685 VSS 0.195519f
C22080 DVSS.n5686 VSS 0.195519f
C22081 DVSS.n5687 VSS 0.195519f
C22082 DVSS.n5688 VSS 0.195519f
C22083 DVSS.n5689 VSS 0.195519f
C22084 DVSS.n5690 VSS 0.195519f
C22085 DVSS.n5691 VSS 0.195519f
C22086 DVSS.n5692 VSS 0.195519f
C22087 DVSS.n5693 VSS 0.195519f
C22088 DVSS.n5694 VSS 0.195519f
C22089 DVSS.n5695 VSS 0.195519f
C22090 DVSS.n5696 VSS 0.195519f
C22091 DVSS.n5697 VSS 0.195519f
C22092 DVSS.n5698 VSS 0.195519f
C22093 DVSS.n5699 VSS 0.195519f
C22094 DVSS.n5700 VSS 0.195519f
C22095 DVSS.n5701 VSS 0.195519f
C22096 DVSS.n5702 VSS 0.195519f
C22097 DVSS.n5703 VSS 0.195519f
C22098 DVSS.n5704 VSS 0.195519f
C22099 DVSS.n5705 VSS 0.195519f
C22100 DVSS.n5706 VSS 0.195519f
C22101 DVSS.n5707 VSS 0.195519f
C22102 DVSS.n5708 VSS 0.195519f
C22103 DVSS.n5709 VSS 0.195519f
C22104 DVSS.n5710 VSS 0.195519f
C22105 DVSS.n5711 VSS 0.195519f
C22106 DVSS.n5712 VSS 0.195519f
C22107 DVSS.n5713 VSS 0.195519f
C22108 DVSS.n5714 VSS 0.195519f
C22109 DVSS.n5715 VSS 0.195519f
C22110 DVSS.n5716 VSS 0.124609f
C22111 DVSS.n5717 VSS 0.097759f
C22112 DVSS.n5718 VSS 0.01141f
C22113 DVSS.n5719 VSS 0.021441f
C22114 DVSS.n5720 VSS 0.022361f
C22115 DVSS.n5721 VSS 0.089424f
C22116 DVSS.n5722 VSS 0.797033f
C22117 DVSS.n5723 VSS 0.643507f
C22118 DVSS.n5724 VSS 1.21903f
C22119 DVSS.n5725 VSS 1.03466f
C22120 DVSS.t92 VSS 4.65162f
C22121 DVSS.t117 VSS 5.1253f
C22122 DVSS.t20 VSS 5.1253f
C22123 DVSS.t53 VSS 5.89821f
C22124 DVSS.n5726 VSS 5.8537f
C22125 DVSS.n5727 VSS 0.025525f
C22126 DVSS.n5728 VSS 0.032524f
C22127 DVSS.n5729 VSS 0.033964f
C22128 DVSS.n5730 VSS 0.013251f
C22129 DVSS.n5731 VSS 0.002945f
C22130 DVSS.n5732 VSS 0.097759f
C22131 DVSS.n5733 VSS 0.168669f
C22132 DVSS.n5734 VSS 0.195519f
C22133 DVSS.n5735 VSS 0.195519f
C22134 DVSS.n5736 VSS 0.195519f
C22135 DVSS.n5737 VSS 0.195519f
C22136 DVSS.n5738 VSS 0.195519f
C22137 DVSS.n5739 VSS 0.114282f
C22138 DVSS.n5740 VSS 0.071599f
C22139 DVSS.n5741 VSS 0.373138f
C22140 DVSS.n5742 VSS 0.178996f
C22141 DVSS.n5743 VSS 0.195519f
C22142 DVSS.n5744 VSS 0.195519f
C22143 DVSS.n5745 VSS 0.195519f
C22144 DVSS.n5746 VSS 0.195519f
C22145 DVSS.n5747 VSS 0.195519f
C22146 DVSS.n5748 VSS 0.195519f
C22147 DVSS.n5749 VSS 0.195519f
C22148 DVSS.n5750 VSS 0.195519f
C22149 DVSS.n5751 VSS 0.195519f
C22150 DVSS.n5752 VSS 0.195519f
C22151 DVSS.n5753 VSS 0.195519f
C22152 DVSS.n5754 VSS 0.195519f
C22153 DVSS.n5755 VSS 0.195519f
C22154 DVSS.n5756 VSS 0.125986f
C22155 DVSS.n5757 VSS 0.195519f
C22156 DVSS.n5758 VSS 0.148016f
C22157 DVSS.n5759 VSS 0.195519f
C22158 DVSS.n5760 VSS 0.195519f
C22159 DVSS.n5761 VSS 0.195519f
C22160 DVSS.n5762 VSS 0.195519f
C22161 DVSS.n5763 VSS 0.195519f
C22162 DVSS.n5764 VSS 0.195519f
C22163 DVSS.n5765 VSS 0.195519f
C22164 DVSS.n5766 VSS 0.195519f
C22165 DVSS.n5767 VSS 0.195519f
C22166 DVSS.n5768 VSS 0.195519f
C22167 DVSS.n5769 VSS 0.195519f
C22168 DVSS.n5770 VSS 0.195519f
C22169 DVSS.n5771 VSS 0.195519f
C22170 DVSS.n5772 VSS 0.195519f
C22171 DVSS.n5773 VSS 0.195519f
C22172 DVSS.n5774 VSS 0.178996f
C22173 DVSS.n5775 VSS 0.178996f
C22174 DVSS.n5776 VSS 0.373138f
C22175 DVSS.n5777 VSS 0.235449f
C22176 DVSS.n5778 VSS 0.178996f
C22177 DVSS.n5779 VSS 0.178996f
C22178 DVSS.n5780 VSS 0.178996f
C22179 DVSS.n5781 VSS 0.195519f
C22180 DVSS.n5782 VSS 0.195519f
C22181 DVSS.n5783 VSS 0.195519f
C22182 DVSS.n5784 VSS 0.195519f
C22183 DVSS.n5785 VSS 0.195519f
C22184 DVSS.n5786 VSS 0.195519f
C22185 DVSS.n5787 VSS 0.195519f
C22186 DVSS.n5788 VSS 0.195519f
C22187 DVSS.n5789 VSS 0.195519f
C22188 DVSS.n5790 VSS 0.195519f
C22189 DVSS.n5791 VSS 0.195519f
C22190 DVSS.n5792 VSS 0.195519f
C22191 DVSS.n5793 VSS 0.195519f
C22192 DVSS.n5794 VSS 0.195519f
C22193 DVSS.n5795 VSS 0.195519f
C22194 DVSS.n5796 VSS 0.195519f
C22195 DVSS.n5797 VSS 0.195519f
C22196 DVSS.n5798 VSS 0.191388f
C22197 DVSS.n5799 VSS 0.191388f
C22198 DVSS.n5800 VSS 0.195519f
C22199 DVSS.n5801 VSS 0.115659f
C22200 DVSS.n5802 VSS 0.10189f
C22201 DVSS.n5803 VSS 0.10189f
C22202 DVSS.n5804 VSS 0.195519f
C22203 DVSS.n5805 VSS 0.195519f
C22204 DVSS.n5806 VSS 0.195519f
C22205 DVSS.n5807 VSS 0.730699f
C22206 DVSS.n5808 VSS 0.356766f
C22207 DVSS.n5809 VSS 0.564545f
C22208 DVSS.n5810 VSS 0.007104f
C22209 DVSS.n5811 VSS 0.098683f
C22210 DVSS.n5812 VSS 0.247841f
C22211 DVSS.n5813 VSS 0.12174f
C22212 DVSS.n5814 VSS 0.352343f
C22213 DVSS.n5815 VSS 0.730699f
C22214 DVSS.n5816 VSS 0.145262f
C22215 DVSS.n5817 VSS 0.167293f
C22216 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t2 VSS 1.55629f
C22217 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t0 VSS 1.49904f
C22218 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t8 VSS 1.23679f
C22219 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t7 VSS 1.35457f
C22220 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n0 VSS 0.969197f
C22221 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t3 VSS 1.23679f
C22222 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t6 VSS 1.35457f
C22223 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n1 VSS 0.969197f
C22224 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n2 VSS 0.255239f
C22225 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t1 VSS 1.87506f
C22226 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n3 VSS 1.17912f
C22227 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t5 VSS 0.624028f
C22228 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t4 VSS 0.718195f
C22229 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n4 VSS 0.810212f
C22230 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t0 VSS 0.227858f
C22231 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t1 VSS 0.789415f
C22232 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t7 VSS 0.785268f
C22233 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t9 VSS 1.58711f
C22234 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t6 VSS 0.785268f
C22235 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t8 VSS 1.58711f
C22236 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t4 VSS 0.785268f
C22237 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t5 VSS 1.58711f
C22238 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.n0 VSS 2.81472f
C22239 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.n1 VSS 2.35462f
C22240 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.n2 VSS 1.65739f
C22241 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t2 VSS 0.785268f
C22242 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A.t3 VSS 1.58711f
C22243 VDD.n0 VSS 0.017489f
C22244 VDD.t59 VSS 0.038343f
C22245 VDD.t53 VSS 0.038343f
C22246 VDD.n1 VSS 0.072898f
C22247 VDD.t58 VSS 0.292125f
C22248 VDD.n2 VSS 0.105718f
C22249 VDD.n3 VSS 0.141622f
C22250 VDD.n4 VSS 0.141622f
C22251 VDD.n5 VSS 0.141622f
C22252 VDD.n6 VSS 0.141622f
C22253 VDD.n7 VSS 0.141622f
C22254 VDD.n8 VSS 0.141622f
C22255 VDD.n9 VSS 0.141622f
C22256 VDD.n10 VSS 0.141622f
C22257 VDD.n11 VSS 0.141622f
C22258 VDD.n12 VSS 0.119681f
C22259 VDD.t22 VSS 0.293345f
C22260 VDD.n13 VSS 0.133643f
C22261 VDD.n14 VSS 0.141622f
C22262 VDD.n15 VSS 0.141622f
C22263 VDD.n16 VSS 0.141622f
C22264 VDD.n17 VSS 0.141622f
C22265 VDD.n18 VSS 0.141622f
C22266 VDD.n19 VSS 0.141622f
C22267 VDD.n20 VSS 0.141622f
C22268 VDD.n21 VSS 0.141622f
C22269 VDD.n22 VSS 0.141622f
C22270 VDD.n23 VSS 0.141622f
C22271 VDD.n24 VSS 0.141622f
C22272 VDD.n25 VSS 0.141622f
C22273 VDD.n26 VSS 0.141622f
C22274 VDD.n27 VSS 0.141622f
C22275 VDD.n28 VSS 0.141622f
C22276 VDD.n29 VSS 0.141622f
C22277 VDD.n30 VSS 0.141622f
C22278 VDD.n31 VSS 0.141622f
C22279 VDD.n32 VSS 0.141622f
C22280 VDD.n33 VSS 0.141622f
C22281 VDD.n34 VSS 0.141622f
C22282 VDD.n35 VSS 0.141622f
C22283 VDD.n36 VSS 0.141622f
C22284 VDD.n37 VSS 0.141622f
C22285 VDD.n38 VSS 0.141622f
C22286 VDD.n39 VSS 0.110705f
C22287 VDD.t48 VSS 0.038343f
C22288 VDD.n40 VSS 0.071805f
C22289 VDD.t54 VSS 0.263699f
C22290 VDD.n41 VSS 0.004753f
C22291 VDD.n42 VSS 0.005027f
C22292 VDD.n43 VSS 0.00595f
C22293 VDD.n44 VSS 0.005027f
C22294 VDD.n45 VSS 0.09057f
C22295 VDD.n48 VSS 0.00595f
C22296 VDD.n49 VSS 0.005027f
C22297 VDD.n50 VSS 0.00595f
C22298 VDD.n51 VSS 0.005027f
C22299 VDD.n52 VSS 0.00595f
C22300 VDD.n53 VSS 0.00595f
C22301 VDD.n54 VSS 0.09057f
C22302 VDD.n55 VSS 0.00595f
C22303 VDD.n56 VSS 0.00595f
C22304 VDD.n57 VSS 0.00595f
C22305 VDD.n58 VSS 0.005027f
C22306 VDD.n59 VSS 0.005027f
C22307 VDD.n60 VSS 0.005027f
C22308 VDD.n61 VSS 0.005027f
C22309 VDD.n63 VSS 0.005027f
C22310 VDD.n64 VSS 0.00595f
C22311 VDD.n65 VSS 0.00595f
C22312 VDD.n66 VSS 0.005027f
C22313 VDD.n67 VSS 0.00595f
C22314 VDD.n68 VSS 0.006873f
C22315 VDD.n69 VSS 0.006873f
C22316 VDD.n71 VSS 0.00595f
C22317 VDD.n72 VSS 0.005027f
C22318 VDD.n73 VSS 0.005027f
C22319 VDD.n74 VSS 0.006873f
C22320 VDD.n75 VSS 0.006873f
C22321 VDD.n77 VSS 0.11087f
C22322 VDD.n79 VSS 0.008925f
C22323 VDD.n80 VSS 0.008925f
C22324 VDD.n81 VSS 0.00595f
C22325 VDD.n82 VSS 0.005027f
C22326 VDD.n83 VSS 0.005027f
C22327 VDD.n84 VSS 0.008925f
C22328 VDD.n85 VSS 0.00595f
C22329 VDD.n86 VSS 0.005027f
C22330 VDD.n87 VSS 0.005027f
C22331 VDD.n88 VSS 0.008925f
C22332 VDD.n89 VSS 0.00595f
C22333 VDD.n90 VSS 0.00595f
C22334 VDD.t19 VSS 0.09057f
C22335 VDD.n91 VSS 0.00595f
C22336 VDD.n92 VSS 0.00595f
C22337 VDD.n93 VSS 0.006873f
C22338 VDD.n94 VSS 0.006873f
C22339 VDD.n96 VSS 0.11087f
C22340 VDD.n98 VSS 0.006873f
C22341 VDD.n99 VSS 0.005463f
C22342 VDD.n100 VSS 0.031332f
C22343 VDD.n101 VSS 5.25574f
C22344 VDD.n102 VSS 0.141622f
C22345 VDD.n103 VSS 0.141622f
C22346 VDD.n104 VSS 0.141622f
C22347 VDD.n105 VSS 0.141622f
C22348 VDD.n106 VSS 0.141622f
C22349 VDD.n107 VSS 0.141622f
C22350 VDD.n108 VSS 0.141622f
C22351 VDD.n109 VSS 0.141622f
C22352 VDD.n110 VSS 0.141622f
C22353 VDD.n111 VSS 0.141622f
C22354 VDD.n112 VSS 0.141622f
C22355 VDD.n113 VSS 0.141622f
C22356 VDD.n114 VSS 3.26028f
C22357 VDD.n115 VSS 0.141622f
C22358 VDD.n116 VSS 0.479377f
C22359 VDD.n117 VSS 0.112201f
C22360 VDD.n118 VSS 2.85234f
C22361 VDD.n119 VSS 0.118742f
C22362 VDD.n120 VSS 0.052788f
C22363 VDD.t21 VSS 0.047284f
C22364 VDD.n121 VSS 0.0812f
C22365 VDD.n122 VSS 0.394944f
C22366 VDD.t20 VSS 0.4184f
C22367 VDD.n123 VSS 0.099804f
C22368 VDD.n124 VSS 0.060576f
C22369 VDD.n125 VSS 0.0216f
C22370 VDD.t55 VSS 0.038343f
C22371 VDD.n126 VSS 0.053359f
C22372 VDD.n127 VSS -0.010986f
C22373 VDD.n128 VSS 0.126609f
C22374 VDD.t47 VSS 0.264953f
C22375 VDD.n129 VSS 0.328885f
C22376 VDD.n130 VSS 0.115346f
C22377 VDD.n131 VSS 0.101728f
C22378 VDD.n132 VSS 0.141622f
C22379 VDD.n133 VSS 0.141622f
C22380 VDD.n134 VSS 0.141622f
C22381 VDD.n135 VSS 0.141622f
C22382 VDD.n136 VSS 0.141622f
C22383 VDD.n137 VSS 0.141622f
C22384 VDD.n138 VSS 0.141622f
C22385 VDD.n139 VSS 0.141622f
C22386 VDD.n140 VSS 0.141622f
C22387 VDD.n141 VSS 0.141622f
C22388 VDD.n142 VSS 0.141622f
C22389 VDD.n143 VSS 0.141622f
C22390 VDD.n144 VSS 0.141622f
C22391 VDD.n145 VSS 0.141622f
C22392 VDD.n146 VSS 0.141622f
C22393 VDD.n147 VSS 0.141622f
C22394 VDD.n148 VSS 0.141622f
C22395 VDD.n149 VSS 0.141622f
C22396 VDD.n150 VSS 0.141622f
C22397 VDD.n151 VSS 0.141622f
C22398 VDD.n152 VSS 0.141622f
C22399 VDD.n153 VSS 0.141622f
C22400 VDD.n154 VSS 0.141622f
C22401 VDD.n155 VSS 0.141622f
C22402 VDD.n156 VSS 0.141622f
C22403 VDD.n157 VSS 0.141622f
C22404 VDD.n158 VSS 0.141622f
C22405 VDD.n159 VSS 0.141622f
C22406 VDD.n160 VSS 0.141622f
C22407 VDD.n161 VSS 0.141622f
C22408 VDD.n162 VSS 0.141622f
C22409 VDD.n163 VSS 0.141622f
C22410 VDD.n164 VSS 0.141622f
C22411 VDD.n165 VSS 0.141622f
C22412 VDD.n166 VSS 0.141622f
C22413 VDD.n167 VSS 0.141622f
C22414 VDD.n168 VSS 0.141622f
C22415 VDD.n169 VSS 0.141622f
C22416 VDD.n170 VSS 0.141622f
C22417 VDD.n171 VSS 0.141622f
C22418 VDD.n172 VSS 0.141622f
C22419 VDD.n173 VSS 0.141622f
C22420 VDD.n174 VSS 0.141622f
C22421 VDD.n175 VSS 0.141622f
C22422 VDD.n176 VSS 0.141622f
C22423 VDD.n177 VSS 0.141622f
C22424 VDD.n178 VSS 0.141622f
C22425 VDD.n179 VSS 0.141622f
C22426 VDD.n180 VSS 0.141622f
C22427 VDD.n181 VSS 0.141622f
C22428 VDD.n182 VSS 0.141622f
C22429 VDD.n183 VSS 0.141622f
C22430 VDD.n184 VSS 0.141622f
C22431 VDD.n185 VSS 0.141622f
C22432 VDD.n186 VSS 0.141622f
C22433 VDD.n187 VSS 0.141622f
C22434 VDD.n188 VSS 0.141622f
C22435 VDD.n189 VSS 0.141622f
C22436 VDD.n190 VSS 0.141622f
C22437 VDD.n191 VSS 0.141622f
C22438 VDD.n192 VSS 0.141622f
C22439 VDD.n193 VSS 0.07879f
C22440 VDD.n194 VSS 0.088781f
C22441 VDD.n195 VSS 0.309947f
C22442 VDD.t23 VSS 0.038343f
C22443 VDD.n196 VSS 0.072898f
C22444 VDD.t51 VSS 0.025824f
C22445 VDD.t49 VSS 0.064977f
C22446 VDD.t65 VSS 0.070262f
C22447 VDD.n197 VSS 0.084175f
C22448 VDD.n198 VSS 0.004346f
C22449 VDD.n199 VSS 0.002342f
C22450 VDD.n200 VSS 0.006155f
C22451 VDD.n201 VSS 0.033853f
C22452 VDD.n202 VSS 0.005232f
C22453 VDD.n203 VSS 0.006155f
C22454 VDD.n204 VSS 0.003693f
C22455 VDD.n205 VSS 0.007078f
C22456 VDD.n206 VSS 0.007078f
C22457 VDD.n207 VSS 0.054164f
C22458 VDD.t60 VSS 0.022568f
C22459 VDD.n208 VSS 0.007078f
C22460 VDD.n211 VSS 0.003693f
C22461 VDD.n212 VSS 0.005232f
C22462 VDD.n213 VSS 0.005232f
C22463 VDD.n214 VSS 0.003693f
C22464 VDD.n215 VSS 0.007078f
C22465 VDD.n216 VSS 0.004616f
C22466 VDD.n217 VSS 0.006155f
C22467 VDD.n218 VSS 0.033853f
C22468 VDD.n219 VSS 0.006155f
C22469 VDD.n220 VSS 0.004616f
C22470 VDD.n221 VSS 0.004616f
C22471 VDD.n222 VSS 0.007078f
C22472 VDD.n223 VSS 0.007078f
C22473 VDD.n224 VSS 0.054164f
C22474 VDD.n225 VSS 0.007078f
C22475 VDD.n226 VSS 0.00289f
C22476 VDD.n227 VSS 0.105427f
C22477 VDD.n228 VSS 0.060235f
C22478 VDD.n229 VSS 0.04516f
C22479 VDD.n230 VSS 0.026432f
C22480 VDD.n231 VSS -0.014f
C22481 VDD.n232 VSS 0.123596f
C22482 VDD.t50 VSS 0.292125f
C22483 VDD.n233 VSS 0.410363f
C22484 VDD.n234 VSS 0.027116f
C22485 VDD.n235 VSS 0.115872f
C22486 VDD.n236 VSS 0.092752f
C22487 VDD.n237 VSS 0.141622f
C22488 VDD.n238 VSS 0.141622f
C22489 VDD.n239 VSS 0.141622f
C22490 VDD.n240 VSS 0.141622f
C22491 VDD.n241 VSS 0.141622f
C22492 VDD.n242 VSS 0.141622f
C22493 VDD.n243 VSS 0.141622f
C22494 VDD.n244 VSS 0.141622f
C22495 VDD.n245 VSS 0.141622f
C22496 VDD.n246 VSS 0.141622f
C22497 VDD.n247 VSS 0.141622f
C22498 VDD.n248 VSS 0.141622f
C22499 VDD.n249 VSS 0.141622f
C22500 VDD.n250 VSS 0.141622f
C22501 VDD.n251 VSS 0.141622f
C22502 VDD.n252 VSS 0.141622f
C22503 VDD.n253 VSS 0.141622f
C22504 VDD.n254 VSS 0.141622f
C22505 VDD.n255 VSS 0.141622f
C22506 VDD.n256 VSS 0.141622f
C22507 VDD.n257 VSS 0.141622f
C22508 VDD.n258 VSS 0.141622f
C22509 VDD.n259 VSS 0.141622f
C22510 VDD.n260 VSS 0.141622f
C22511 VDD.n261 VSS 0.141622f
C22512 VDD.n262 VSS 0.141622f
C22513 VDD.n263 VSS 0.141622f
C22514 VDD.n264 VSS 0.141622f
C22515 VDD.n265 VSS 0.141622f
C22516 VDD.n266 VSS 0.141622f
C22517 VDD.n267 VSS 0.141622f
C22518 VDD.n268 VSS 0.141622f
C22519 VDD.n269 VSS 0.141622f
C22520 VDD.n270 VSS 0.141622f
C22521 VDD.n271 VSS 0.083776f
C22522 VDD.t25 VSS 0.038343f
C22523 VDD.n272 VSS 0.072893f
C22524 VDD.t6 VSS 0.294644f
C22525 VDD.n274 VSS 0.070811f
C22526 VDD.n275 VSS 0.13115f
C22527 VDD.n276 VSS 0.040463f
C22528 VDD.n277 VSS 0.040463f
C22529 VDD.n278 VSS 0.040463f
C22530 VDD.n279 VSS 0.040463f
C22531 VDD.n281 VSS 0.043747f
C22532 VDD.n282 VSS 0.039309f
C22533 VDD.n284 VSS 0.071053f
C22534 VDD.n285 VSS 0.035334f
C22535 VDD.n286 VSS 0.005027f
C22536 VDD.n287 VSS 0.036773f
C22537 VDD.n288 VSS 0.00595f
C22538 VDD.n289 VSS 0.154975f
C22539 VDD.n290 VSS 0.006873f
C22540 VDD.n291 VSS 0.175684f
C22541 VDD.n292 VSS 0.003056f
C22542 VDD.n294 VSS 0.00595f
C22543 VDD.n295 VSS 0.491663f
C22544 VDD.n297 VSS 0.003817f
C22545 VDD.n299 VSS 0.006873f
C22546 VDD.n300 VSS 0.126599f
C22547 VDD.n301 VSS 0.005027f
C22548 VDD.n302 VSS 0.036773f
C22549 VDD.n304 VSS 0.00595f
C22550 VDD.t36 VSS 0.126599f
C22551 VDD.n305 VSS 0.00595f
C22552 VDD.n306 VSS 0.00595f
C22553 VDD.n307 VSS 0.00595f
C22554 VDD.n308 VSS 0.00595f
C22555 VDD.n309 VSS 0.010976f
C22556 VDD.n310 VSS 0.00595f
C22557 VDD.n311 VSS 0.006873f
C22558 VDD.n312 VSS 0.154975f
C22559 VDD.n313 VSS 0.00595f
C22560 VDD.n314 VSS 0.00595f
C22561 VDD.n315 VSS 0.006873f
C22562 VDD.n317 VSS 0.005027f
C22563 VDD.n318 VSS 0.005027f
C22564 VDD.n319 VSS 0.005027f
C22565 VDD.n320 VSS 0.005027f
C22566 VDD.n322 VSS 0.006873f
C22567 VDD.n324 VSS 0.00595f
C22568 VDD.n325 VSS 0.006873f
C22569 VDD.n326 VSS 0.003817f
C22570 VDD.n327 VSS 0.003056f
C22571 VDD.n328 VSS 0.00595f
C22572 VDD.n329 VSS 0.005027f
C22573 VDD.n330 VSS 0.00595f
C22574 VDD.n331 VSS 0.003056f
C22575 VDD.n332 VSS 0.003817f
C22576 VDD.n333 VSS 0.005027f
C22577 VDD.n334 VSS 0.005027f
C22578 VDD.n335 VSS 0.010976f
C22579 VDD.n336 VSS 0.005027f
C22580 VDD.n337 VSS 0.005027f
C22581 VDD.n338 VSS 0.00595f
C22582 VDD.n340 VSS 0.005027f
C22583 VDD.n341 VSS 0.005027f
C22584 VDD.n342 VSS 0.012777f
C22585 VDD.n343 VSS 0.402851f
C22586 VDD.t64 VSS 0.030006f
C22587 VDD.n344 VSS 0.071094f
C22588 VDD.n345 VSS 0.063863f
C22589 VDD.t14 VSS 0.030006f
C22590 VDD.n346 VSS 0.071094f
C22591 VDD.n347 VSS 0.022232f
C22592 VDD.n348 VSS 0.03715f
C22593 VDD.t63 VSS 0.248821f
C22594 VDD.n349 VSS 0.071746f
C22595 VDD.n350 VSS 0.019893f
C22596 VDD.n351 VSS 0.019786f
C22597 VDD.n352 VSS 0.019699f
C22598 VDD.n353 VSS 0.022232f
C22599 VDD.n354 VSS 0.03715f
C22600 VDD.n355 VSS 0.035551f
C22601 VDD.n356 VSS 0.046643f
C22602 VDD.n357 VSS 0.314342f
C22603 VDD.t13 VSS 0.248821f
C22604 VDD.n358 VSS 0.071746f
C22605 VDD.n359 VSS 0.402851f
C22606 VDD.n360 VSS 0.021826f
C22607 VDD.n361 VSS 0.052373f
C22608 VDD.t1 VSS 0.041955f
C22609 VDD.n362 VSS 0.055972f
C22610 VDD.n363 VSS 0.032754f
C22611 VDD.n364 VSS 0.351015f
C22612 VDD.t0 VSS 0.249418f
C22613 VDD.n365 VSS 0.071746f
C22614 VDD.n366 VSS 0.510776f
C22615 VDD.n367 VSS 0.178825f
C22616 VDD.n368 VSS 0.050987f
C22617 VDD.n369 VSS 0.043444f
C22618 VDD.n370 VSS 0.050771f
C22619 VDD.n371 VSS 0.148993f
C22620 VDD.n372 VSS 0.148993f
C22621 VDD.n373 VSS 0.402851f
C22622 VDD.n374 VSS 0.333462f
C22623 VDD.t45 VSS 0.249418f
C22624 VDD.n375 VSS 0.071746f
C22625 VDD.n376 VSS 0.052373f
C22626 VDD.n377 VSS 0.022232f
C22627 VDD.n378 VSS 0.016419f
C22628 VDD.n379 VSS 0.019893f
C22629 VDD.t46 VSS 0.030006f
C22630 VDD.n380 VSS 0.071094f
C22631 VDD.n381 VSS 0.082655f
C22632 VDD.n382 VSS 0.099469f
C22633 VDD.n383 VSS 0.196277f
C22634 VDD.n384 VSS 0.036773f
C22635 VDD.n385 VSS 0.00595f
C22636 VDD.n386 VSS 0.126599f
C22637 VDD.n387 VSS 0.00595f
C22638 VDD.n388 VSS 0.00595f
C22639 VDD.n389 VSS 0.00595f
C22640 VDD.n390 VSS 0.006873f
C22641 VDD.n391 VSS 0.006873f
C22642 VDD.n393 VSS 0.005027f
C22643 VDD.n394 VSS 0.005027f
C22644 VDD.n395 VSS 0.005027f
C22645 VDD.n396 VSS 0.005027f
C22646 VDD.n397 VSS 0.003817f
C22647 VDD.n398 VSS 0.003056f
C22648 VDD.n399 VSS 0.00595f
C22649 VDD.n400 VSS 0.126599f
C22650 VDD.n401 VSS 0.00595f
C22651 VDD.n402 VSS 0.006873f
C22652 VDD.n403 VSS 0.126579f
C22653 VDD.n404 VSS 0.126579f
C22654 VDD.n405 VSS 0.00595f
C22655 VDD.n406 VSS 0.00595f
C22656 VDD.n407 VSS 0.00595f
C22657 VDD.n408 VSS 0.00595f
C22658 VDD.n411 VSS 0.005027f
C22659 VDD.n412 VSS 0.005027f
C22660 VDD.n413 VSS 0.006873f
C22661 VDD.n414 VSS 0.00595f
C22662 VDD.n415 VSS 0.00595f
C22663 VDD.n416 VSS 0.00595f
C22664 VDD.n417 VSS 0.006873f
C22665 VDD.n418 VSS 0.006873f
C22666 VDD.n419 VSS 0.005027f
C22667 VDD.n420 VSS 0.005027f
C22668 VDD.n421 VSS 0.00595f
C22669 VDD.n422 VSS 0.005027f
C22670 VDD.n423 VSS 0.00595f
C22671 VDD.n424 VSS 0.007514f
C22672 VDD.n425 VSS 0.006873f
C22673 VDD.n426 VSS 0.00595f
C22674 VDD.n427 VSS 0.126599f
C22675 VDD.n428 VSS 0.003056f
C22676 VDD.n429 VSS 0.00595f
C22677 VDD.n430 VSS 0.00595f
C22678 VDD.n432 VSS 0.00595f
C22679 VDD.t12 VSS 0.126599f
C22680 VDD.n433 VSS 0.00595f
C22681 VDD.n434 VSS 0.036773f
C22682 VDD.n435 VSS 0.00595f
C22683 VDD.n436 VSS 0.005549f
C22684 VDD.n437 VSS 0.005027f
C22685 VDD.n438 VSS 0.00595f
C22686 VDD.n439 VSS 0.005027f
C22687 VDD.n440 VSS 0.005027f
C22688 VDD.n441 VSS 0.006873f
C22689 VDD.n442 VSS 0.491663f
C22690 VDD.n443 VSS 0.003817f
C22691 VDD.n444 VSS 0.005027f
C22692 VDD.n445 VSS 0.005549f
C22693 VDD.n446 VSS 0.171145f
C22694 VDD.n447 VSS 0.008566f
C22695 VDD.n448 VSS 0.00595f
C22696 VDD.n449 VSS 0.005027f
C22697 VDD.n451 VSS 0.00595f
C22698 VDD.n452 VSS 0.005027f
C22699 VDD.n454 VSS 0.006873f
C22700 VDD.n455 VSS 0.091607f
C22701 VDD.n456 VSS 0.090823f
C22702 VDD.n458 VSS 0.039309f
C22703 VDD.n459 VSS 0.046162f
C22704 VDD.n460 VSS 2.52e-19
C22705 VDD.n461 VSS 0.043495f
C22706 VDD.n462 VSS 0.111844f
C22707 VDD.n463 VSS 0.111844f
C22708 VDD.n464 VSS 0.085117f
C22709 VDD.n465 VSS 0.035334f
C22710 VDD.n467 VSS 0.442248f
C22711 VDD.n468 VSS 0.444813f
C22712 VDD.n469 VSS 0.070811f
C22713 VDD.n471 VSS 0.040463f
C22714 VDD.n473 VSS 0.040463f
C22715 VDD.n475 VSS 0.040463f
C22716 VDD.n476 VSS 0.070811f
C22717 VDD.n480 VSS 0.141622f
C22718 VDD.n481 VSS 0.139627f
C22719 VDD.n482 VSS 0.015957f
C22720 VDD.n483 VSS 0.141622f
C22721 VDD.n484 VSS 0.141622f
C22722 VDD.n485 VSS 0.141622f
C22723 VDD.n486 VSS 0.141622f
C22724 VDD.n487 VSS 0.141622f
C22725 VDD.n488 VSS 0.141622f
C22726 VDD.n489 VSS 0.141622f
C22727 VDD.n490 VSS 0.141622f
C22728 VDD.n491 VSS 0.141622f
C22729 VDD.n492 VSS 0.141622f
C22730 VDD.n493 VSS 0.141622f
C22731 VDD.n494 VSS 0.141622f
C22732 VDD.n495 VSS 0.141622f
C22733 VDD.n496 VSS 0.141622f
C22734 VDD.n497 VSS 0.141622f
C22735 VDD.n498 VSS 0.141622f
C22736 VDD.n499 VSS 0.141622f
C22737 VDD.n500 VSS 0.141622f
C22738 VDD.n501 VSS 0.141622f
C22739 VDD.n502 VSS 0.141622f
C22740 VDD.n503 VSS 0.141622f
C22741 VDD.n504 VSS 0.141622f
C22742 VDD.n505 VSS 0.141622f
C22743 VDD.n506 VSS 0.141622f
C22744 VDD.n507 VSS 0.141622f
C22745 VDD.n508 VSS 0.141622f
C22746 VDD.n509 VSS 0.141622f
C22747 VDD.n510 VSS 0.141622f
C22748 VDD.n511 VSS 0.141622f
C22749 VDD.n512 VSS 0.141622f
C22750 VDD.n513 VSS 0.141622f
C22751 VDD.n514 VSS 0.141622f
C22752 VDD.n515 VSS 0.141622f
C22753 VDD.n516 VSS 0.141622f
C22754 VDD.n517 VSS 0.141622f
C22755 VDD.n518 VSS 0.141622f
C22756 VDD.n519 VSS 0.141622f
C22757 VDD.n520 VSS 0.141622f
C22758 VDD.n521 VSS 0.141622f
C22759 VDD.n522 VSS 0.141622f
C22760 VDD.n523 VSS 0.141622f
C22761 VDD.n524 VSS 0.141622f
C22762 VDD.n525 VSS 0.141622f
C22763 VDD.n526 VSS 0.141622f
C22764 VDD.n527 VSS 0.141622f
C22765 VDD.n528 VSS 0.141622f
C22766 VDD.n529 VSS 0.141622f
C22767 VDD.n530 VSS 0.141622f
C22768 VDD.n531 VSS 0.141622f
C22769 VDD.n532 VSS 0.141622f
C22770 VDD.n533 VSS 0.141622f
C22771 VDD.n534 VSS 0.141622f
C22772 VDD.n535 VSS 0.141622f
C22773 VDD.n536 VSS 0.141622f
C22774 VDD.n537 VSS 0.141622f
C22775 VDD.n538 VSS 0.141622f
C22776 VDD.n539 VSS 0.141622f
C22777 VDD.n540 VSS 0.141622f
C22778 VDD.n541 VSS 0.141622f
C22779 VDD.n542 VSS 0.141622f
C22780 VDD.n543 VSS 0.141622f
C22781 VDD.n544 VSS 0.141622f
C22782 VDD.n545 VSS 0.141622f
C22783 VDD.n546 VSS 0.141622f
C22784 VDD.n547 VSS 0.141622f
C22785 VDD.n548 VSS 0.141622f
C22786 VDD.n549 VSS 0.141622f
C22787 VDD.n550 VSS 0.141622f
C22788 VDD.n551 VSS 0.141622f
C22789 VDD.n552 VSS 0.141622f
C22790 VDD.n553 VSS 0.141622f
C22791 VDD.n554 VSS 0.141622f
C22792 VDD.n555 VSS 0.120678f
C22793 VDD.t42 VSS 0.034774f
C22794 VDD.n556 VSS 0.073966f
C22795 VDD.t26 VSS 0.195427f
C22796 VDD.n557 VSS 0.838056f
C22797 VDD.n558 VSS 0.141622f
C22798 VDD.n559 VSS 0.141622f
C22799 VDD.n560 VSS 0.141622f
C22800 VDD.n561 VSS 0.141622f
C22801 VDD.n562 VSS 0.141622f
C22802 VDD.n563 VSS 0.141622f
C22803 VDD.n564 VSS 0.141622f
C22804 VDD.n565 VSS 0.141622f
C22805 VDD.n566 VSS 0.141622f
C22806 VDD.n567 VSS 0.141622f
C22807 VDD.n568 VSS 0.141622f
C22808 VDD.n569 VSS 0.141622f
C22809 VDD.n570 VSS 0.141622f
C22810 VDD.n571 VSS 0.141622f
C22811 VDD.n572 VSS 0.141622f
C22812 VDD.n573 VSS 0.141622f
C22813 VDD.n574 VSS 0.141622f
C22814 VDD.t62 VSS 0.038343f
C22815 VDD.n575 VSS 0.054086f
C22816 VDD.t2 VSS 0.222621f
C22817 VDD.t56 VSS 0.402215f
C22818 VDD.t3 VSS 0.037442f
C22819 VDD.n576 VSS 0.057572f
C22820 VDD.n577 VSS 0.010691f
C22821 VDD.n578 VSS 0.300415f
C22822 VDD.t5 VSS 0.037442f
C22823 VDD.n579 VSS -0.011615f
C22824 VDD.t32 VSS 0.295445f
C22825 VDD.n580 VSS 0.128587f
C22826 VDD.t33 VSS 0.279774f
C22827 VDD.t8 VSS 0.417875f
C22828 VDD.t9 VSS 0.041947f
C22829 VDD.n581 VSS 0.058362f
C22830 VDD.t11 VSS 0.037442f
C22831 VDD.n582 VSS 0.121783f
C22832 VDD.n583 VSS 0.288985f
C22833 VDD.t10 VSS 0.224167f
C22834 VDD.t4 VSS 0.222621f
C22835 VDD.n584 VSS 0.088484f
C22836 VDD.n585 VSS 0.044457f
C22837 VDD.n586 VSS 0.133401f
C22838 VDD.n587 VSS 0.050619f
C22839 VDD.n588 VSS 0.029815f
C22840 VDD.n589 VSS 0.02767f
C22841 VDD.t57 VSS 0.041049f
C22842 VDD.n590 VSS 0.063229f
C22843 VDD.n591 VSS 0.031049f
C22844 VDD.n592 VSS 0.010691f
C22845 VDD.n593 VSS 0.018514f
C22846 VDD.n594 VSS 0.332023f
C22847 VDD.n595 VSS -0.015187f
C22848 VDD.n596 VSS 0.088484f
C22849 VDD.t61 VSS 0.224247f
C22850 VDD.n597 VSS 0.443879f
C22851 VDD.n598 VSS 0.228379f
C22852 VDD.n599 VSS 0.071136f
C22853 VDD.n600 VSS 0.141622f
C22854 VDD.n601 VSS 0.141622f
C22855 VDD.n602 VSS 0.141622f
C22856 VDD.n603 VSS 0.08627f
C22857 VDD.n604 VSS 0.141622f
C22858 VDD.n605 VSS 0.141622f
C22859 VDD.n606 VSS 0.141622f
C22860 VDD.n607 VSS 0.141622f
C22861 VDD.n608 VSS 0.141622f
C22862 VDD.n609 VSS 0.141622f
C22863 VDD.n610 VSS 0.141622f
C22864 VDD.n611 VSS 0.141622f
C22865 VDD.n612 VSS 0.141622f
C22866 VDD.n613 VSS 0.141622f
C22867 VDD.n614 VSS 0.055851f
C22868 VDD.n615 VSS 0.071133f
C22869 VDD.n616 VSS 0.141123f
C22870 VDD.n617 VSS 0.141622f
C22871 VDD.n618 VSS 0.141622f
C22872 VDD.n619 VSS 0.141622f
C22873 VDD.n620 VSS 0.141622f
C22874 VDD.n621 VSS 0.141622f
C22875 VDD.n622 VSS 0.141622f
C22876 VDD.n623 VSS 0.141622f
C22877 VDD.n624 VSS 0.141622f
C22878 VDD.n625 VSS 0.141622f
C22879 VDD.n626 VSS 0.141622f
C22880 VDD.n627 VSS 0.141622f
C22881 VDD.n628 VSS 0.141622f
C22882 VDD.n629 VSS 0.141622f
C22883 VDD.n630 VSS 0.141622f
C22884 VDD.n631 VSS 0.141622f
C22885 VDD.n632 VSS 0.141622f
C22886 VDD.n633 VSS 0.141622f
C22887 VDD.n634 VSS 0.141622f
C22888 VDD.n635 VSS 0.141622f
C22889 VDD.n636 VSS 0.141622f
C22890 VDD.n637 VSS 0.141622f
C22891 VDD.n638 VSS 0.141622f
C22892 VDD.n639 VSS 0.141622f
C22893 VDD.n640 VSS 0.141622f
C22894 VDD.n641 VSS 0.141622f
C22895 VDD.n642 VSS 0.141622f
C22896 VDD.n643 VSS 0.141622f
C22897 VDD.n644 VSS 0.141622f
C22898 VDD.n645 VSS 0.981831f
C22899 VDD.n646 VSS 0.141622f
C22900 VDD.n647 VSS 0.274251f
C22901 VDD.n648 VSS 0.133145f
C22902 VDD.n649 VSS 0.818007f
C22903 VDD.t17 VSS 0.224925f
C22904 VDD.t30 VSS 0.224925f
C22905 VDD.t34 VSS 0.224925f
C22906 VDD.t15 VSS 0.300754f
C22907 VDD.n650 VSS 0.409718f
C22908 VDD.t16 VSS 0.046856f
C22909 VDD.n651 VSS 0.074363f
C22910 VDD.t35 VSS 0.012965f
C22911 VDD.t31 VSS 0.012965f
C22912 VDD.n652 VSS 0.042855f
C22913 VDD.n653 VSS 0.054956f
C22914 VDD.t18 VSS 0.012965f
C22915 VDD.t27 VSS 0.012965f
C22916 VDD.n654 VSS 0.042855f
C22917 VDD.n655 VSS 0.049119f
C22918 VDD.t29 VSS 0.046856f
C22919 VDD.t44 VSS 0.034774f
C22920 VDD.t38 VSS 0.009261f
C22921 VDD.t40 VSS 0.009261f
C22922 VDD.n656 VSS 0.032673f
C22923 VDD.n657 VSS 0.056023f
C22924 VDD.n658 VSS 0.060796f
C22925 VDD.n659 VSS 0.054858f
C22926 VDD.n660 VSS -0.087449f
C22927 VDD.n661 VSS 0.019176f
C22928 VDD.t28 VSS 0.221238f
C22929 VDD.t43 VSS 0.304202f
C22930 VDD.t37 VSS 0.224925f
C22931 VDD.t39 VSS 0.224925f
C22932 VDD.t41 VSS 0.261027f
C22933 VDD.n662 VSS 0.229552f
C22934 VDD.n663 VSS 0.084197f
C22935 VDD.n664 VSS 0.091755f
C22936 VDD.n665 VSS 0.141622f
C22937 VDD.n666 VSS 0.141622f
C22938 VDD.n667 VSS 0.141622f
C22939 VDD.n668 VSS 0.141622f
C22940 VDD.n669 VSS 0.141622f
C22941 VDD.n670 VSS 0.141622f
C22942 VDD.n671 VSS 0.141622f
C22943 VDD.n672 VSS 0.141622f
C22944 VDD.n673 VSS 0.141622f
C22945 VDD.n674 VSS 0.141622f
C22946 VDD.n675 VSS 0.141622f
C22947 VDD.n676 VSS 0.141622f
C22948 VDD.n677 VSS 0.141622f
C22949 VDD.n678 VSS 0.141622f
C22950 VDD.n679 VSS 0.141622f
C22951 VDD.n680 VSS 0.141622f
C22952 VDD.n681 VSS 0.141622f
C22953 VDD.n682 VSS 0.141622f
C22954 VDD.n683 VSS 0.141622f
C22955 VDD.n684 VSS 0.141622f
C22956 VDD.n685 VSS 0.141622f
C22957 VDD.n686 VSS 0.141622f
C22958 VDD.n687 VSS 0.141622f
C22959 VDD.n688 VSS 0.141622f
C22960 VDD.n689 VSS 0.141622f
C22961 VDD.n690 VSS 0.141622f
C22962 VDD.n691 VSS 0.141622f
C22963 VDD.n692 VSS 0.141622f
C22964 VDD.n693 VSS 0.141622f
C22965 VDD.n694 VSS 0.141622f
C22966 VDD.n695 VSS 0.141622f
C22967 VDD.n696 VSS 0.141622f
C22968 VDD.n697 VSS 0.141622f
C22969 VDD.n698 VSS 0.141622f
C22970 VDD.n699 VSS 0.141622f
C22971 VDD.n700 VSS 0.141622f
C22972 VDD.n701 VSS 0.141622f
C22973 VDD.n702 VSS 0.141622f
C22974 VDD.n703 VSS 0.141622f
C22975 VDD.n704 VSS 0.141622f
C22976 VDD.n705 VSS 0.141622f
C22977 VDD.n706 VSS 0.141622f
C22978 VDD.n707 VSS 0.141622f
C22979 VDD.n708 VSS 0.141622f
C22980 VDD.n709 VSS 0.141622f
C22981 VDD.n710 VSS 0.141622f
C22982 VDD.n711 VSS 0.141622f
C22983 VDD.n712 VSS 0.141622f
C22984 VDD.n713 VSS 0.141622f
C22985 VDD.n714 VSS 0.141622f
C22986 VDD.n715 VSS 0.141622f
C22987 VDD.n716 VSS 0.141622f
C22988 VDD.n717 VSS 0.141622f
C22989 VDD.n718 VSS 0.141622f
C22990 VDD.n719 VSS 0.141622f
C22991 VDD.n720 VSS 0.141622f
C22992 VDD.n721 VSS 0.141622f
C22993 VDD.n722 VSS 0.141622f
C22994 VDD.n723 VSS 0.141622f
C22995 VDD.n724 VSS 0.141622f
C22996 VDD.n725 VSS 0.141622f
C22997 VDD.n726 VSS 0.141622f
C22998 VDD.n727 VSS 0.141622f
C22999 VDD.n728 VSS 0.141622f
C23000 VDD.n729 VSS 0.141622f
C23001 VDD.n730 VSS 0.141622f
C23002 VDD.n731 VSS 0.141622f
C23003 VDD.n732 VSS 0.141622f
C23004 VDD.n733 VSS 0.141622f
C23005 VDD.n734 VSS 0.141622f
C23006 VDD.n735 VSS 0.141622f
C23007 VDD.n736 VSS 0.141622f
C23008 VDD.n737 VSS 0.141622f
C23009 VDD.n738 VSS 0.141622f
C23010 VDD.n739 VSS 0.141622f
C23011 VDD.n740 VSS 0.141622f
C23012 VDD.n741 VSS 0.141622f
C23013 VDD.n742 VSS 0.141622f
C23014 VDD.n743 VSS 0.141622f
C23015 VDD.n744 VSS 0.141622f
C23016 VDD.n745 VSS 0.141622f
C23017 VDD.n746 VSS 0.141622f
C23018 VDD.n747 VSS 0.141622f
C23019 VDD.n748 VSS 0.141622f
C23020 VDD.n749 VSS 0.141622f
C23021 VDD.n750 VSS 0.141622f
C23022 VDD.n751 VSS 0.141622f
C23023 VDD.n752 VSS 0.141622f
C23024 VDD.n753 VSS 0.141622f
C23025 VDD.n754 VSS 0.141622f
C23026 VDD.n755 VSS 0.141622f
C23027 VDD.n756 VSS 0.141622f
C23028 VDD.n757 VSS 0.141622f
C23029 VDD.n758 VSS 0.141622f
C23030 VDD.n759 VSS 0.141622f
C23031 VDD.n760 VSS 0.141622f
C23032 VDD.n761 VSS 0.141622f
C23033 VDD.n762 VSS 0.141622f
C23034 VDD.n763 VSS 0.141622f
C23035 VDD.n764 VSS 0.141622f
C23036 VDD.n765 VSS 0.141622f
C23037 VDD.n766 VSS 0.141622f
C23038 VDD.n767 VSS 0.141622f
C23039 VDD.n768 VSS 0.141622f
C23040 VDD.n769 VSS 0.141622f
C23041 VDD.n770 VSS 0.141622f
C23042 VDD.n771 VSS 0.141622f
C23043 VDD.n772 VSS 0.141622f
C23044 VDD.n773 VSS 0.141622f
C23045 VDD.n774 VSS 0.141622f
C23046 VDD.n775 VSS 0.141622f
C23047 VDD.n776 VSS 0.141622f
C23048 VDD.n777 VSS 0.141622f
C23049 VDD.n778 VSS 0.141622f
C23050 VDD.n779 VSS 0.141622f
C23051 VDD.n780 VSS 0.141622f
C23052 VDD.n781 VSS 0.141622f
C23053 VDD.n782 VSS 0.141622f
C23054 VDD.n783 VSS 0.141622f
C23055 VDD.n784 VSS 0.141622f
C23056 VDD.n785 VSS 0.141622f
C23057 VDD.n786 VSS 0.141622f
C23058 VDD.n787 VSS 0.141622f
C23059 VDD.n788 VSS 0.141622f
C23060 VDD.n789 VSS 0.141622f
C23061 VDD.n790 VSS 0.141622f
C23062 VDD.n791 VSS 0.141622f
C23063 VDD.n792 VSS 0.141622f
C23064 VDD.n793 VSS 0.141622f
C23065 VDD.n794 VSS 0.141622f
C23066 VDD.n795 VSS 0.141622f
C23067 VDD.n796 VSS 0.141622f
C23068 VDD.n797 VSS 0.141622f
C23069 VDD.n798 VSS 0.141622f
C23070 VDD.n799 VSS 0.141622f
C23071 VDD.n800 VSS 0.141622f
C23072 VDD.n801 VSS 0.141622f
C23073 VDD.n802 VSS 0.141622f
C23074 VDD.n803 VSS 0.141622f
C23075 VDD.n804 VSS 0.127659f
C23076 VDD.n805 VSS 0.127659f
C23077 VDD.n806 VSS 0.127659f
C23078 VDD.n807 VSS 0.084774f
C23079 VDD.n808 VSS 0.084774f
C23080 VDD.n809 VSS 0.141622f
C23081 VDD.n810 VSS 0.141622f
C23082 VDD.n811 VSS 0.528613f
C23083 VDD.n812 VSS 0.270928f
C23084 VDD.n813 VSS 0.272098f
C23085 VDD.n816 VSS 0.040463f
C23086 VDD.n817 VSS 0.070811f
C23087 VDD.n818 VSS 1.35581f
C23088 VDD.n820 VSS 0.272098f
C23089 VDD.n821 VSS 0.13115f
C23090 VDD.n822 VSS 0.040463f
C23091 VDD.n823 VSS 0.040463f
C23092 VDD.n824 VSS 0.040463f
C23093 VDD.n825 VSS 0.040463f
C23094 VDD.n826 VSS 0.070811f
C23095 VDD.n828 VSS 0.040463f
C23096 VDD.n830 VSS 0.040463f
C23097 VDD.n832 VSS 0.040463f
C23098 VDD.n834 VSS 0.040463f
C23099 VDD.n835 VSS 0.141622f
C23100 VDD.n836 VSS 0.072806f
C23101 VDD.n837 VSS 0.141622f
C23102 VDD.n838 VSS 0.141622f
C23103 VDD.n839 VSS 0.141622f
C23104 VDD.n840 VSS 0.141622f
C23105 VDD.n841 VSS 0.141622f
C23106 VDD.n842 VSS 0.141622f
C23107 VDD.n843 VSS 0.141622f
C23108 VDD.n844 VSS 0.141622f
C23109 VDD.n845 VSS 0.141622f
C23110 VDD.n846 VSS 0.141622f
C23111 VDD.n847 VSS 0.141622f
C23112 VDD.n848 VSS 0.141622f
C23113 VDD.n849 VSS 0.141622f
C23114 VDD.n850 VSS 0.141622f
C23115 VDD.n851 VSS 0.141622f
C23116 VDD.n852 VSS 0.141622f
C23117 VDD.n853 VSS 0.127659f
C23118 VDD.n854 VSS 0.127659f
C23119 VDD.n855 VSS 0.084774f
C23120 VDD.n856 VSS 0.084774f
C23121 VDD.n857 VSS 0.141622f
C23122 VDD.n858 VSS 0.139627f
C23123 VDD.n859 VSS 0.528613f
C23124 VDD.n860 VSS 0.270928f
C23125 VDD.n861 VSS 0.141622f
C23126 VDD.n862 VSS 0.070811f
C23127 VDD.n866 VSS 0.070811f
C23128 VDD.n868 VSS 0.035619f
C23129 VDD.n869 VSS 0.070811f
C23130 VDD.n870 VSS 0.098309f
C23131 VDD.n871 VSS 1.42132f
C23132 VDD.n872 VSS 0.380286f
C23133 VDD.t7 VSS 0.038343f
C23134 VDD.n873 VSS 0.054909f
C23135 VDD.n874 VSS -0.014f
C23136 VDD.n875 VSS 0.123596f
C23137 VDD.t24 VSS 0.293345f
C23138 VDD.n876 VSS 0.308315f
C23139 VDD.n877 VSS 0.089135f
C23140 VDD.n878 VSS 0.128657f
C23141 VDD.n879 VSS 0.141622f
C23142 VDD.n880 VSS 0.141622f
C23143 VDD.n881 VSS 0.141622f
C23144 VDD.n882 VSS 0.141622f
C23145 VDD.n883 VSS 0.141622f
C23146 VDD.n884 VSS 0.141622f
C23147 VDD.n885 VSS 0.141622f
C23148 VDD.n886 VSS 0.141622f
C23149 VDD.n887 VSS 0.141622f
C23150 VDD.n888 VSS 0.141622f
C23151 VDD.n889 VSS 0.141622f
C23152 VDD.n890 VSS 0.141622f
C23153 VDD.n891 VSS 0.141622f
C23154 VDD.n892 VSS 0.141622f
C23155 VDD.n893 VSS 0.141622f
C23156 VDD.n894 VSS 0.141622f
C23157 VDD.n895 VSS 0.141622f
C23158 VDD.n896 VSS 0.141622f
C23159 VDD.n897 VSS 0.141622f
C23160 VDD.n898 VSS 0.141622f
C23161 VDD.n899 VSS 0.141622f
C23162 VDD.n900 VSS 0.141622f
C23163 VDD.n901 VSS 0.141622f
C23164 VDD.n902 VSS 0.141622f
C23165 VDD.n903 VSS 0.141622f
C23166 VDD.n904 VSS 0.141622f
C23167 VDD.n905 VSS 0.141622f
C23168 VDD.n906 VSS 0.141622f
C23169 VDD.n907 VSS 0.141622f
C23170 VDD.n908 VSS 0.141622f
C23171 VDD.n909 VSS 0.141622f
C23172 VDD.n910 VSS 0.141622f
C23173 VDD.n911 VSS 0.141622f
C23174 VDD.n912 VSS 0.141622f
C23175 VDD.n913 VSS 0.141622f
C23176 VDD.n914 VSS 0.141622f
C23177 VDD.n915 VSS 0.141622f
C23178 VDD.n916 VSS 0.141622f
C23179 VDD.n917 VSS 0.141622f
C23180 VDD.n918 VSS 0.141622f
C23181 VDD.n919 VSS 0.141622f
C23182 VDD.n920 VSS 0.141622f
C23183 VDD.n921 VSS 0.141622f
C23184 VDD.n922 VSS 0.141622f
C23185 VDD.n923 VSS 0.141622f
C23186 VDD.n924 VSS 0.106715f
C23187 VDD.n925 VSS 0.088781f
C23188 VDD.n926 VSS 0.309947f
C23189 VDD.t52 VSS 0.293345f
C23190 VDD.n927 VSS 0.123596f
C23191 VDD.n928 VSS -0.014f
C23192 VDD.n929 VSS 0.054909f
C23193 CS.t1 VSS 0.699042f
C23194 CS.t2 VSS 0.46855f
C23195 CS.n0 VSS 0.746188f
C23196 CS.t0 VSS 0.33386f
C23197 CS.n1 VSS 0.141089f
C23198 CS.n2 VSS 4.58968f
C23199 SL.t2 VSS 0.410577f
C23200 SL.n0 VSS 0.46338f
C23201 SL.n1 VSS 8.832179f
C23202 SL.t1 VSS 0.956628f
C23203 SL.t0 VSS 0.57598f
C23204 SL.n2 VSS 1.0146f
.ends

